module Benchmark_testing25000(I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1863,I1871,I1879,I1887,I1895,I1903,I1911,I1919,I1927,I1935,I1943,I1951,I1959,I1967,I1975,I1983,I1991,I1999,I2007,I2015,I2023,I2031,I2039,I2047,I2055,I2063,I2071,I2079,I2087,I2095,I2103,I2111,I2119,I2127,I2135,I2143,I2151,I2159,I2167,I2175,I2183,I2191,I2199,I2207,I2215,I2223,I2231,I2239,I2247,I2255,I2263,I2271,I2279,I2287,I2295,I2303,I2311,I2319,I2327,I2335,I2343,I2351,I2359,I2367,I2375,I2383,I2391,I2399,I2407,I2415,I2423,I2431,I2439,I2447,I2455,I2463,I2471,I2479,I2487,I2495,I2503,I2511,I2519,I2527,I2535,I2543,I2551,I2559,I2567,I2575,I2583,I2591,I2599,I2607,I2615,I2623,I2631,I2639,I2647,I2655,I2663,I2671,I2679,I2687,I2695,I2703,I2711,I2719,I2727,I2735,I2743,I2751,I2759,I2767,I2775,I2783,I2791,I2799,I2807,I2815,I2823,I2831,I2839,I2847,I2855,I2863,I2871,I2879,I2887,I2895,I2903,I2911,I2919,I2927,I2935,I2943,I2951,I2959,I2967,I2975,I2983,I2991,I2999,I3007,I3015,I3023,I3031,I3039,I3047,I3055,I3063,I3071,I3079,I3087,I3095,I3103,I3111,I3119,I3127,I3135,I3143,I3151,I3159,I3167,I3175,I3183,I3191,I3199,I3207,I3215,I3223,I3231,I3239,I3247,I3255,I3263,I3271,I3279,I3287,I3295,I3303,I3311,I3319,I3327,I3335,I3343,I3351,I3359,I3367,I3375,I3383,I3391,I3399,I3407,I3415,I3423,I3431,I3439,I3447,I3455,I3463,I3471,I3479,I3487,I3495,I3503,I3511,I3519,I3527,I3535,I3543,I3551,I3559,I3567,I3575,I3583,I3591,I3599,I3607,I3615,I3623,I3631,I3639,I3647,I3655,I3663,I3671,I3679,I3687,I3695,I3703,I3711,I3719,I3727,I3735,I3743,I3751,I3759,I3767,I3775,I3783,I3791,I3799,I3807,I3815,I3823,I3831,I3839,I3847,I3855,I3863,I3871,I3879,I3887,I3895,I3903,I3911,I3919,I3927,I3935,I3943,I3951,I3959,I3967,I3975,I3983,I3991,I3999,I4007,I4015,I4023,I4031,I4039,I4047,I4055,I4063,I4071,I4079,I4087,I4095,I4103,I4111,I4119,I4127,I4135,I4143,I4151,I4159,I4167,I4175,I4183,I4191,I4199,I4207,I4215,I4223,I4231,I4239,I4247,I4255,I4263,I4271,I4279,I4287,I4295,I4303,I4311,I4319,I4327,I4335,I4343,I4351,I4359,I4367,I4375,I4383,I4391,I4399,I4407,I4415,I4423,I4431,I4439,I4447,I4455,I4463,I4471,I4479,I4487,I4495,I4503,I4511,I4519,I4527,I4535,I4543,I4551,I4559,I4567,I4575,I4583,I4591,I4599,I4607,I4615,I4623,I4631,I4639,I4647,I4655,I4663,I4671,I4679,I4687,I4695,I4703,I4711,I4719,I4727,I4735,I4743,I4751,I4759,I4767,I4775,I4783,I4791,I4799,I4807,I4815,I4823,I4831,I4839,I4847,I4855,I4863,I4871,I4879,I4887,I4895,I4903,I4911,I4919,I4927,I4935,I4943,I4951,I4959,I4967,I4975,I4983,I4991,I4999,I5007,I5015,I5023,I5031,I5039,I5047,I5055,I5063,I5071,I5079,I5087,I5095,I5103,I5111,I5119,I5127,I5135,I5143,I5151,I5159,I5167,I5175,I5183,I5191,I5199,I5207,I5215,I5223,I5231,I5239,I5247,I5255,I5263,I5271,I5279,I5287,I5295,I5303,I5311,I5319,I5327,I5335,I5343,I5351,I5359,I5367,I5375,I5383,I5391,I5399,I5407,I5415,I5423,I5431,I5439,I5447,I5455,I5463,I5471,I5479,I5487,I5495,I5503,I5511,I5519,I5527,I5535,I5543,I5551,I5559,I5567,I5575,I5583,I5591,I5599,I5607,I5615,I5623,I5631,I5639,I5647,I5655,I5663,I5671,I5679,I5687,I5694_clk,I5701,I260625,I260628,I260622,I260631,I260637,I260640,I260619,I260649,I260646,I260634,I260643,I270568,I270571,I270553,I270574,I270565,I270556,I270547,I270577,I270562,I270559,I270550,I273543,I273546,I273528,I273549,I273540,I273531,I273522,I273552,I273537,I273534,I273525,I282049,I282022,I282043,I282028,I282025,I282031,I282037,I282052,I282040,I282046,I282034,I289829,I289817,I289826,I289835,I289814,I289832,I289823,I289838,I289811,I289820,I289808,I295039,I295054,I295036,I295051,I295033,I295030,I295045,I295042,I295048,I295057,I295027,I304763,I304757,I304754,I304766,I304751,I304772,I304781,I304775,I304778,I304769,I304760,I305358,I305352,I305349,I305361,I305346,I305367,I305376,I305370,I305373,I305364,I305355,I306548,I306542,I306539,I306551,I306536,I306557,I306566,I306560,I306563,I306554,I306545,I307747,I307726,I307753,I307756,I307741,I307744,I307738,I307732,I307750,I307735,I307729,I310932,I310917,I310914,I310911,I310929,I310926,I310905,I310908,I310935,I310920,I310923,I318802,I318799,I318793,I318823,I318796,I318820,I318817,I318814,I318808,I318811,I318805,I324817,I324820,I324814,I324823,I324829,I324832,I324811,I324841,I324838,I324826,I324835,I325395,I325398,I325392,I325401,I325407,I325410,I325389,I325419,I325416,I325404,I325413,I330153,I330156,I330138,I330159,I330150,I330141,I330132,I330162,I330147,I330144,I330135,I331331,I331328,I331322,I331349,I331340,I331334,I331337,I331352,I331346,I331343,I331325,I333797,I333770,I333791,I333776,I333773,I333779,I333785,I333800,I333788,I333794,I333782,I340421,I340409,I340418,I340427,I340406,I340424,I340415,I340430,I340403,I340412,I340400,I340982,I340970,I340979,I340988,I340967,I340985,I340976,I340991,I340964,I340973,I340961,I346617,I346632,I346614,I346629,I346611,I346608,I346623,I346620,I346626,I346635,I346605,I347909,I347924,I347906,I347921,I347903,I347900,I347915,I347912,I347918,I347927,I347897,I349198,I349213,I349210,I349195,I349192,I349219,I349207,I349201,I349216,I349204,I349189,I350524,I350539,I350536,I350521,I350518,I350545,I350533,I350527,I350542,I350530,I350515,I352380,I352374,I352371,I352383,I352368,I352389,I352398,I352392,I352395,I352386,I352377,I353653,I353638,I353635,I353632,I353650,I353647,I353626,I353629,I353656,I353641,I353644,I354979,I354964,I354961,I354958,I354976,I354973,I354952,I354955,I354982,I354967,I354970,I356305,I356290,I356287,I356284,I356302,I356299,I356278,I356281,I356308,I356293,I356296,I357631,I357616,I357613,I357610,I357628,I357625,I357604,I357607,I357634,I357619,I357622,I360283,I360268,I360265,I360262,I360280,I360277,I360256,I360259,I360286,I360271,I360274,I360946,I360931,I360928,I360925,I360943,I360940,I360919,I360922,I360949,I360934,I360937,I362237,I362234,I362228,I362258,I362231,I362255,I362252,I362249,I362243,I362246,I362240,I362883,I362880,I362874,I362904,I362877,I362901,I362898,I362895,I362889,I362892,I362886,I364784,I364787,I364781,I364790,I364796,I364799,I364778,I364808,I364805,I364793,I364802,I365940,I365946,I365937,I365961,I365949,I365955,I365943,I365934,I365964,I365958,I365952,I366573,I366558,I366555,I366567,I366561,I366576,I366546,I366564,I366570,I366549,I366552,I367145,I367148,I367130,I367151,I367142,I367133,I367124,I367154,I367139,I367136,I367127,I368335,I368338,I368320,I368341,I368332,I368323,I368314,I368344,I368329,I368326,I368317,I369525,I369528,I369510,I369531,I369522,I369513,I369504,I369534,I369519,I369516,I369507,I371316,I371289,I371310,I371295,I371292,I371298,I371304,I371319,I371307,I371313,I371301,I373781,I373769,I373772,I373757,I373763,I373775,I373784,I373754,I373778,I373766,I373760,I374914,I374902,I374911,I374920,I374899,I374917,I374908,I374923,I374896,I374905,I374893,I375475,I375463,I375472,I375481,I375460,I375478,I375469,I375484,I375457,I375466,I375454,I376027,I376042,I376024,I376039,I376021,I376018,I376033,I376030,I376036,I376045,I376015,I376670,I376685,I376682,I376667,I376664,I376691,I376679,I376673,I376688,I376676,I376661,I379136,I379121,I379118,I379115,I379133,I379130,I379109,I379112,I379139,I379124,I379127,I380441,I380444,I380438,I380447,I380453,I380456,I380435,I380465,I380462,I380450,I380459,I381019,I381022,I381016,I381025,I381031,I381034,I381013,I381043,I381040,I381028,I381037,I381597,I381600,I381594,I381603,I381609,I381612,I381591,I381621,I381618,I381606,I381615,I382190,I382193,I382175,I382196,I382187,I382178,I382169,I382199,I382184,I382181,I382172,I383422,I383437,I383419,I383434,I383416,I383413,I383428,I383425,I383431,I383440,I383410,I384083,I384068,I384065,I384062,I384080,I384077,I384056,I384059,I384086,I384071,I384074);
input I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1863,I1871,I1879,I1887,I1895,I1903,I1911,I1919,I1927,I1935,I1943,I1951,I1959,I1967,I1975,I1983,I1991,I1999,I2007,I2015,I2023,I2031,I2039,I2047,I2055,I2063,I2071,I2079,I2087,I2095,I2103,I2111,I2119,I2127,I2135,I2143,I2151,I2159,I2167,I2175,I2183,I2191,I2199,I2207,I2215,I2223,I2231,I2239,I2247,I2255,I2263,I2271,I2279,I2287,I2295,I2303,I2311,I2319,I2327,I2335,I2343,I2351,I2359,I2367,I2375,I2383,I2391,I2399,I2407,I2415,I2423,I2431,I2439,I2447,I2455,I2463,I2471,I2479,I2487,I2495,I2503,I2511,I2519,I2527,I2535,I2543,I2551,I2559,I2567,I2575,I2583,I2591,I2599,I2607,I2615,I2623,I2631,I2639,I2647,I2655,I2663,I2671,I2679,I2687,I2695,I2703,I2711,I2719,I2727,I2735,I2743,I2751,I2759,I2767,I2775,I2783,I2791,I2799,I2807,I2815,I2823,I2831,I2839,I2847,I2855,I2863,I2871,I2879,I2887,I2895,I2903,I2911,I2919,I2927,I2935,I2943,I2951,I2959,I2967,I2975,I2983,I2991,I2999,I3007,I3015,I3023,I3031,I3039,I3047,I3055,I3063,I3071,I3079,I3087,I3095,I3103,I3111,I3119,I3127,I3135,I3143,I3151,I3159,I3167,I3175,I3183,I3191,I3199,I3207,I3215,I3223,I3231,I3239,I3247,I3255,I3263,I3271,I3279,I3287,I3295,I3303,I3311,I3319,I3327,I3335,I3343,I3351,I3359,I3367,I3375,I3383,I3391,I3399,I3407,I3415,I3423,I3431,I3439,I3447,I3455,I3463,I3471,I3479,I3487,I3495,I3503,I3511,I3519,I3527,I3535,I3543,I3551,I3559,I3567,I3575,I3583,I3591,I3599,I3607,I3615,I3623,I3631,I3639,I3647,I3655,I3663,I3671,I3679,I3687,I3695,I3703,I3711,I3719,I3727,I3735,I3743,I3751,I3759,I3767,I3775,I3783,I3791,I3799,I3807,I3815,I3823,I3831,I3839,I3847,I3855,I3863,I3871,I3879,I3887,I3895,I3903,I3911,I3919,I3927,I3935,I3943,I3951,I3959,I3967,I3975,I3983,I3991,I3999,I4007,I4015,I4023,I4031,I4039,I4047,I4055,I4063,I4071,I4079,I4087,I4095,I4103,I4111,I4119,I4127,I4135,I4143,I4151,I4159,I4167,I4175,I4183,I4191,I4199,I4207,I4215,I4223,I4231,I4239,I4247,I4255,I4263,I4271,I4279,I4287,I4295,I4303,I4311,I4319,I4327,I4335,I4343,I4351,I4359,I4367,I4375,I4383,I4391,I4399,I4407,I4415,I4423,I4431,I4439,I4447,I4455,I4463,I4471,I4479,I4487,I4495,I4503,I4511,I4519,I4527,I4535,I4543,I4551,I4559,I4567,I4575,I4583,I4591,I4599,I4607,I4615,I4623,I4631,I4639,I4647,I4655,I4663,I4671,I4679,I4687,I4695,I4703,I4711,I4719,I4727,I4735,I4743,I4751,I4759,I4767,I4775,I4783,I4791,I4799,I4807,I4815,I4823,I4831,I4839,I4847,I4855,I4863,I4871,I4879,I4887,I4895,I4903,I4911,I4919,I4927,I4935,I4943,I4951,I4959,I4967,I4975,I4983,I4991,I4999,I5007,I5015,I5023,I5031,I5039,I5047,I5055,I5063,I5071,I5079,I5087,I5095,I5103,I5111,I5119,I5127,I5135,I5143,I5151,I5159,I5167,I5175,I5183,I5191,I5199,I5207,I5215,I5223,I5231,I5239,I5247,I5255,I5263,I5271,I5279,I5287,I5295,I5303,I5311,I5319,I5327,I5335,I5343,I5351,I5359,I5367,I5375,I5383,I5391,I5399,I5407,I5415,I5423,I5431,I5439,I5447,I5455,I5463,I5471,I5479,I5487,I5495,I5503,I5511,I5519,I5527,I5535,I5543,I5551,I5559,I5567,I5575,I5583,I5591,I5599,I5607,I5615,I5623,I5631,I5639,I5647,I5655,I5663,I5671,I5679,I5687,I5694_clk,I5701;
output I260625,I260628,I260622,I260631,I260637,I260640,I260619,I260649,I260646,I260634,I260643,I270568,I270571,I270553,I270574,I270565,I270556,I270547,I270577,I270562,I270559,I270550,I273543,I273546,I273528,I273549,I273540,I273531,I273522,I273552,I273537,I273534,I273525,I282049,I282022,I282043,I282028,I282025,I282031,I282037,I282052,I282040,I282046,I282034,I289829,I289817,I289826,I289835,I289814,I289832,I289823,I289838,I289811,I289820,I289808,I295039,I295054,I295036,I295051,I295033,I295030,I295045,I295042,I295048,I295057,I295027,I304763,I304757,I304754,I304766,I304751,I304772,I304781,I304775,I304778,I304769,I304760,I305358,I305352,I305349,I305361,I305346,I305367,I305376,I305370,I305373,I305364,I305355,I306548,I306542,I306539,I306551,I306536,I306557,I306566,I306560,I306563,I306554,I306545,I307747,I307726,I307753,I307756,I307741,I307744,I307738,I307732,I307750,I307735,I307729,I310932,I310917,I310914,I310911,I310929,I310926,I310905,I310908,I310935,I310920,I310923,I318802,I318799,I318793,I318823,I318796,I318820,I318817,I318814,I318808,I318811,I318805,I324817,I324820,I324814,I324823,I324829,I324832,I324811,I324841,I324838,I324826,I324835,I325395,I325398,I325392,I325401,I325407,I325410,I325389,I325419,I325416,I325404,I325413,I330153,I330156,I330138,I330159,I330150,I330141,I330132,I330162,I330147,I330144,I330135,I331331,I331328,I331322,I331349,I331340,I331334,I331337,I331352,I331346,I331343,I331325,I333797,I333770,I333791,I333776,I333773,I333779,I333785,I333800,I333788,I333794,I333782,I340421,I340409,I340418,I340427,I340406,I340424,I340415,I340430,I340403,I340412,I340400,I340982,I340970,I340979,I340988,I340967,I340985,I340976,I340991,I340964,I340973,I340961,I346617,I346632,I346614,I346629,I346611,I346608,I346623,I346620,I346626,I346635,I346605,I347909,I347924,I347906,I347921,I347903,I347900,I347915,I347912,I347918,I347927,I347897,I349198,I349213,I349210,I349195,I349192,I349219,I349207,I349201,I349216,I349204,I349189,I350524,I350539,I350536,I350521,I350518,I350545,I350533,I350527,I350542,I350530,I350515,I352380,I352374,I352371,I352383,I352368,I352389,I352398,I352392,I352395,I352386,I352377,I353653,I353638,I353635,I353632,I353650,I353647,I353626,I353629,I353656,I353641,I353644,I354979,I354964,I354961,I354958,I354976,I354973,I354952,I354955,I354982,I354967,I354970,I356305,I356290,I356287,I356284,I356302,I356299,I356278,I356281,I356308,I356293,I356296,I357631,I357616,I357613,I357610,I357628,I357625,I357604,I357607,I357634,I357619,I357622,I360283,I360268,I360265,I360262,I360280,I360277,I360256,I360259,I360286,I360271,I360274,I360946,I360931,I360928,I360925,I360943,I360940,I360919,I360922,I360949,I360934,I360937,I362237,I362234,I362228,I362258,I362231,I362255,I362252,I362249,I362243,I362246,I362240,I362883,I362880,I362874,I362904,I362877,I362901,I362898,I362895,I362889,I362892,I362886,I364784,I364787,I364781,I364790,I364796,I364799,I364778,I364808,I364805,I364793,I364802,I365940,I365946,I365937,I365961,I365949,I365955,I365943,I365934,I365964,I365958,I365952,I366573,I366558,I366555,I366567,I366561,I366576,I366546,I366564,I366570,I366549,I366552,I367145,I367148,I367130,I367151,I367142,I367133,I367124,I367154,I367139,I367136,I367127,I368335,I368338,I368320,I368341,I368332,I368323,I368314,I368344,I368329,I368326,I368317,I369525,I369528,I369510,I369531,I369522,I369513,I369504,I369534,I369519,I369516,I369507,I371316,I371289,I371310,I371295,I371292,I371298,I371304,I371319,I371307,I371313,I371301,I373781,I373769,I373772,I373757,I373763,I373775,I373784,I373754,I373778,I373766,I373760,I374914,I374902,I374911,I374920,I374899,I374917,I374908,I374923,I374896,I374905,I374893,I375475,I375463,I375472,I375481,I375460,I375478,I375469,I375484,I375457,I375466,I375454,I376027,I376042,I376024,I376039,I376021,I376018,I376033,I376030,I376036,I376045,I376015,I376670,I376685,I376682,I376667,I376664,I376691,I376679,I376673,I376688,I376676,I376661,I379136,I379121,I379118,I379115,I379133,I379130,I379109,I379112,I379139,I379124,I379127,I380441,I380444,I380438,I380447,I380453,I380456,I380435,I380465,I380462,I380450,I380459,I381019,I381022,I381016,I381025,I381031,I381034,I381013,I381043,I381040,I381028,I381037,I381597,I381600,I381594,I381603,I381609,I381612,I381591,I381621,I381618,I381606,I381615,I382190,I382193,I382175,I382196,I382187,I382178,I382169,I382199,I382184,I382181,I382172,I383422,I383437,I383419,I383434,I383416,I383413,I383428,I383425,I383431,I383440,I383410,I384083,I384068,I384065,I384062,I384080,I384077,I384056,I384059,I384086,I384071,I384074;
wire I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1863,I1871,I1879,I1887,I1895,I1903,I1911,I1919,I1927,I1935,I1943,I1951,I1959,I1967,I1975,I1983,I1991,I1999,I2007,I2015,I2023,I2031,I2039,I2047,I2055,I2063,I2071,I2079,I2087,I2095,I2103,I2111,I2119,I2127,I2135,I2143,I2151,I2159,I2167,I2175,I2183,I2191,I2199,I2207,I2215,I2223,I2231,I2239,I2247,I2255,I2263,I2271,I2279,I2287,I2295,I2303,I2311,I2319,I2327,I2335,I2343,I2351,I2359,I2367,I2375,I2383,I2391,I2399,I2407,I2415,I2423,I2431,I2439,I2447,I2455,I2463,I2471,I2479,I2487,I2495,I2503,I2511,I2519,I2527,I2535,I2543,I2551,I2559,I2567,I2575,I2583,I2591,I2599,I2607,I2615,I2623,I2631,I2639,I2647,I2655,I2663,I2671,I2679,I2687,I2695,I2703,I2711,I2719,I2727,I2735,I2743,I2751,I2759,I2767,I2775,I2783,I2791,I2799,I2807,I2815,I2823,I2831,I2839,I2847,I2855,I2863,I2871,I2879,I2887,I2895,I2903,I2911,I2919,I2927,I2935,I2943,I2951,I2959,I2967,I2975,I2983,I2991,I2999,I3007,I3015,I3023,I3031,I3039,I3047,I3055,I3063,I3071,I3079,I3087,I3095,I3103,I3111,I3119,I3127,I3135,I3143,I3151,I3159,I3167,I3175,I3183,I3191,I3199,I3207,I3215,I3223,I3231,I3239,I3247,I3255,I3263,I3271,I3279,I3287,I3295,I3303,I3311,I3319,I3327,I3335,I3343,I3351,I3359,I3367,I3375,I3383,I3391,I3399,I3407,I3415,I3423,I3431,I3439,I3447,I3455,I3463,I3471,I3479,I3487,I3495,I3503,I3511,I3519,I3527,I3535,I3543,I3551,I3559,I3567,I3575,I3583,I3591,I3599,I3607,I3615,I3623,I3631,I3639,I3647,I3655,I3663,I3671,I3679,I3687,I3695,I3703,I3711,I3719,I3727,I3735,I3743,I3751,I3759,I3767,I3775,I3783,I3791,I3799,I3807,I3815,I3823,I3831,I3839,I3847,I3855,I3863,I3871,I3879,I3887,I3895,I3903,I3911,I3919,I3927,I3935,I3943,I3951,I3959,I3967,I3975,I3983,I3991,I3999,I4007,I4015,I4023,I4031,I4039,I4047,I4055,I4063,I4071,I4079,I4087,I4095,I4103,I4111,I4119,I4127,I4135,I4143,I4151,I4159,I4167,I4175,I4183,I4191,I4199,I4207,I4215,I4223,I4231,I4239,I4247,I4255,I4263,I4271,I4279,I4287,I4295,I4303,I4311,I4319,I4327,I4335,I4343,I4351,I4359,I4367,I4375,I4383,I4391,I4399,I4407,I4415,I4423,I4431,I4439,I4447,I4455,I4463,I4471,I4479,I4487,I4495,I4503,I4511,I4519,I4527,I4535,I4543,I4551,I4559,I4567,I4575,I4583,I4591,I4599,I4607,I4615,I4623,I4631,I4639,I4647,I4655,I4663,I4671,I4679,I4687,I4695,I4703,I4711,I4719,I4727,I4735,I4743,I4751,I4759,I4767,I4775,I4783,I4791,I4799,I4807,I4815,I4823,I4831,I4839,I4847,I4855,I4863,I4871,I4879,I4887,I4895,I4903,I4911,I4919,I4927,I4935,I4943,I4951,I4959,I4967,I4975,I4983,I4991,I4999,I5007,I5015,I5023,I5031,I5039,I5047,I5055,I5063,I5071,I5079,I5087,I5095,I5103,I5111,I5119,I5127,I5135,I5143,I5151,I5159,I5167,I5175,I5183,I5191,I5199,I5207,I5215,I5223,I5231,I5239,I5247,I5255,I5263,I5271,I5279,I5287,I5295,I5303,I5311,I5319,I5327,I5335,I5343,I5351,I5359,I5367,I5375,I5383,I5391,I5399,I5407,I5415,I5423,I5431,I5439,I5447,I5455,I5463,I5471,I5479,I5487,I5495,I5503,I5511,I5519,I5527,I5535,I5543,I5551,I5559,I5567,I5575,I5583,I5591,I5599,I5607,I5615,I5623,I5631,I5639,I5647,I5655,I5663,I5671,I5679,I5687,I5694_clk,I5701,I5742_rst,I5759,I5776,I5793,I5810,I5827,I5725,I5713,I5872,I5889,I5906,I5923,I5940,I5722,I5971,I5988,I6005,I6022,I5731,I5710,I6067,I6084,I5728,I6115,I5719,I5734,I6160,I6177,I6194,I6211,I5707,I5716,I5704,I6303_rst,I6320,I6337,I6354,I6371,I6388,I6286,I6274,I6433,I6450,I6467,I6484,I6501,I6283,I6532,I6549,I6566,I6583,I6292,I6271,I6628,I6645,I6289,I6676,I6280,I6295,I6721,I6738,I6755,I6772,I6268,I6277,I6265,I6864_rst,I6881,I6898,I6915,I6838,I6946,I6963,I6853,I6835,I7008,I7025,I7042,I7059,I7076,I7093,I7110,I7127,I7144,I6850,I7175,I7192,I7209,I6832,I7240,I6829,I7271,I7288,I7305,I7322,I6844,I7353,I6841,I7384,I7401,I7418,I6847,I6856,I6826,I7510_rst,I7527,I7544,I7561,I7481,I7592,I7609,I7626,I7643,I7660,I7677,I7694,I7711,I7728,I7745,I7496,I7493,I7790,I7478,I7821,I7475,I7852,I7869,I7886,I7903,I7920,I7937,I7502,I7968,I7490,I7484,I8013,I8030,I7499,I8061,I8078,I8095,I7487,I7472,I8173_rst,I8190,I8207,I8224,I8144,I8255,I8272,I8289,I8306,I8323,I8340,I8357,I8374,I8391,I8408,I8159,I8156,I8453,I8141,I8484,I8138,I8515,I8532,I8549,I8566,I8583,I8600,I8165,I8631,I8153,I8147,I8676,I8693,I8162,I8724,I8741,I8758,I8150,I8135,I8836_rst,I8853,I8870,I8887,I8807,I8918,I8935,I8952,I8969,I8986,I9003,I9020,I9037,I9054,I9071,I8822,I8819,I9116,I8804,I9147,I8801,I9178,I9195,I9212,I9229,I9246,I9263,I8828,I9294,I8816,I8810,I9339,I9356,I8825,I9387,I9404,I9421,I8813,I8798,I9499_rst,I9516,I9533,I9550,I9470,I9581,I9598,I9615,I9632,I9649,I9666,I9683,I9700,I9717,I9734,I9485,I9482,I9779,I9467,I9810,I9464,I9841,I9858,I9875,I9892,I9909,I9926,I9491,I9957,I9479,I9473,I10002,I10019,I9488,I10050,I10067,I10084,I9476,I9461,I10162_rst,I10179,I10196,I10213,I10133,I10244,I10261,I10278,I10295,I10312,I10329,I10346,I10363,I10380,I10397,I10148,I10145,I10442,I10130,I10473,I10127,I10504,I10521,I10538,I10555,I10572,I10589,I10154,I10620,I10142,I10136,I10665,I10682,I10151,I10713,I10730,I10747,I10139,I10124,I10825_rst,I10842,I10859,I10876,I10796,I10907,I10924,I10941,I10958,I10975,I10992,I11009,I11026,I11043,I11060,I10811,I10808,I11105,I10793,I11136,I10790,I11167,I11184,I11201,I11218,I11235,I11252,I10817,I11283,I10805,I10799,I11328,I11345,I10814,I11376,I11393,I11410,I10802,I10787,I11488_rst,I11505,I11522,I11462,I11553,I11570,I11587,I11604,I11621,I11638,I11655,I11672,I11689,I11456,I11720,I11737,I11453,I11768,I11785,I11802,I11465,I11450,I11847,I11864,I11881,I11898,I11915,I11471,I11946,I11480,I11977,I11474,I11477,I11468,I11459,I12083_rst,I12100,I12117,I12057,I12148,I12165,I12182,I12199,I12216,I12233,I12250,I12267,I12284,I12051,I12315,I12332,I12048,I12363,I12380,I12397,I12060,I12045,I12442,I12459,I12476,I12493,I12510,I12066,I12541,I12075,I12572,I12069,I12072,I12063,I12054,I12678_rst,I12695,I12712,I12729,I12746,I12763,I12780,I12797,I12667,I12828,I12652,I12859,I12876,I12893,I12910,I12927,I12944,I12961,I12649,I12992,I13009,I12646,I13040,I13057,I12664,I13088,I12661,I13119,I13136,I12640,I12643,I13181,I13198,I13215,I13232,I12670,I13263,I12655,I12658,I13341_rst,I13358,I13375,I13392,I13409,I13426,I13443,I13460,I13330,I13491,I13315,I13522,I13539,I13556,I13573,I13590,I13607,I13624,I13312,I13655,I13672,I13309,I13703,I13720,I13327,I13751,I13324,I13782,I13799,I13303,I13306,I13844,I13861,I13878,I13895,I13333,I13926,I13318,I13321,I14004_rst,I14021,I14038,I14055,I14072,I14089,I14106,I14123,I13993,I14154,I13978,I14185,I14202,I14219,I14236,I14253,I14270,I14287,I13975,I14318,I14335,I13972,I14366,I14383,I13990,I14414,I13987,I14445,I14462,I13966,I13969,I14507,I14524,I14541,I14558,I13996,I14589,I13981,I13984,I14667_rst,I14684,I14701,I14718,I14735,I14752,I14769,I14786,I14656,I14817,I14641,I14848,I14865,I14882,I14899,I14916,I14933,I14950,I14638,I14981,I14998,I14635,I15029,I15046,I14653,I15077,I14650,I15108,I15125,I14629,I14632,I15170,I15187,I15204,I15221,I14659,I15252,I14644,I14647,I15330_rst,I15347,I15364,I15381,I15398,I15415,I15432,I15449,I15319,I15480,I15304,I15511,I15528,I15545,I15562,I15579,I15596,I15613,I15301,I15644,I15661,I15298,I15692,I15709,I15316,I15740,I15313,I15771,I15788,I15292,I15295,I15833,I15850,I15867,I15884,I15322,I15915,I15307,I15310,I15993_rst,I16010,I16027,I16044,I16061,I16078,I16095,I16112,I15982,I16143,I15967,I16174,I16191,I16208,I16225,I16242,I16259,I16276,I15964,I16307,I16324,I15961,I16355,I16372,I15979,I16403,I15976,I16434,I16451,I15955,I15958,I16496,I16513,I16530,I16547,I15985,I16578,I15970,I15973,I16656_rst,I16673,I16690,I16707,I16724,I16741,I16758,I16775,I16645,I16806,I16630,I16837,I16854,I16871,I16888,I16905,I16922,I16939,I16627,I16970,I16987,I16624,I17018,I17035,I16642,I17066,I16639,I17097,I17114,I16618,I16621,I17159,I17176,I17193,I17210,I16648,I17241,I16633,I16636,I17319_rst,I17336,I17353,I17370,I17387,I17404,I17421,I17438,I17308,I17469,I17293,I17500,I17517,I17534,I17551,I17568,I17585,I17602,I17290,I17633,I17650,I17287,I17681,I17698,I17305,I17729,I17302,I17760,I17777,I17281,I17284,I17822,I17839,I17856,I17873,I17311,I17904,I17296,I17299,I17982_rst,I17999,I18016,I18033,I18050,I18067,I18084,I17953,I18115,I18132,I18149,I18166,I18183,I18200,I18217,I17950,I18248,I17944,I18279,I18296,I18313,I17974,I17947,I18358,I17971,I18389,I17968,I17965,I18434,I18451,I18468,I18485,I18502,I17959,I18533,I18550,I17962,I17956,I18628_rst,I18645,I18662,I18679,I18696,I18713,I18730,I18599,I18761,I18778,I18795,I18812,I18829,I18846,I18863,I18596,I18894,I18590,I18925,I18942,I18959,I18620,I18593,I19004,I18617,I19035,I18614,I18611,I19080,I19097,I19114,I19131,I19148,I18605,I19179,I19196,I18608,I18602,I19274_rst,I19291,I19308,I19325,I19342,I19359,I19376,I19245,I19407,I19424,I19441,I19458,I19475,I19492,I19509,I19242,I19540,I19236,I19571,I19588,I19605,I19266,I19239,I19650,I19263,I19681,I19260,I19257,I19726,I19743,I19760,I19777,I19794,I19251,I19825,I19842,I19254,I19248,I19920_rst,I19937,I19954,I19971,I19988,I20005,I20022,I19891,I20053,I20070,I20087,I20104,I20121,I20138,I20155,I19888,I20186,I19882,I20217,I20234,I20251,I19912,I19885,I20296,I19909,I20327,I19906,I19903,I20372,I20389,I20406,I20423,I20440,I19897,I20471,I20488,I19900,I19894,I20566_rst,I20583,I20600,I20617,I20634,I20651,I20668,I20537,I20699,I20716,I20733,I20750,I20767,I20784,I20801,I20534,I20832,I20528,I20863,I20880,I20897,I20558,I20531,I20942,I20555,I20973,I20552,I20549,I21018,I21035,I21052,I21069,I21086,I20543,I21117,I21134,I20546,I20540,I21212_rst,I21229,I21246,I21263,I21280,I21174,I21311,I21328,I21345,I21362,I21379,I21396,I21183,I21427,I21177,I21458,I21475,I21492,I21509,I21204,I21201,I21554,I21571,I21588,I21198,I21619,I21195,I21186,I21664,I21681,I21698,I21189,I21192,I21743,I21760,I21180,I21824_rst,I21841,I21858,I21875,I21892,I21786,I21923,I21940,I21957,I21974,I21991,I22008,I21795,I22039,I21789,I22070,I22087,I22104,I22121,I21816,I21813,I22166,I22183,I22200,I21810,I22231,I21807,I21798,I22276,I22293,I22310,I21801,I21804,I22355,I22372,I21792,I22436_rst,I22453,I22470,I22487,I22504,I22398,I22535,I22552,I22569,I22586,I22603,I22620,I22407,I22651,I22401,I22682,I22699,I22716,I22733,I22428,I22425,I22778,I22795,I22812,I22422,I22843,I22419,I22410,I22888,I22905,I22922,I22413,I22416,I22967,I22984,I22404,I23048_rst,I23065,I23082,I23099,I23116,I23016,I23147,I23164,I23181,I23019,I23212,I23013,I23243,I23260,I23277,I23294,I23311,I23022,I23342,I23359,I23376,I23393,I23028,I23031,I23010,I23452,I23469,I23486,I23040,I23037,I23531,I23548,I23025,I23034,I23626_rst,I23643,I23660,I23677,I23694,I23594,I23725,I23742,I23759,I23597,I23790,I23591,I23821,I23838,I23855,I23872,I23889,I23600,I23920,I23937,I23954,I23971,I23606,I23609,I23588,I24030,I24047,I24064,I23618,I23615,I24109,I24126,I23603,I23612,I24204_rst,I24221,I24238,I24255,I24272,I24172,I24303,I24320,I24337,I24175,I24368,I24169,I24399,I24416,I24433,I24450,I24467,I24178,I24498,I24515,I24532,I24549,I24184,I24187,I24166,I24608,I24625,I24642,I24196,I24193,I24687,I24704,I24181,I24190,I24782_rst,I24799,I24816,I24833,I24850,I24750,I24881,I24898,I24915,I24753,I24946,I24747,I24977,I24994,I25011,I25028,I25045,I24756,I25076,I25093,I25110,I25127,I24762,I24765,I24744,I25186,I25203,I25220,I24774,I24771,I25265,I25282,I24759,I24768,I25360_rst,I25377,I25394,I25411,I25428,I25328,I25459,I25476,I25493,I25510,I25527,I25544,I25561,I25578,I25334,I25325,I25623,I25640,I25349,I25671,I25688,I25337,I25719,I25736,I25343,I25767,I25331,I25798,I25322,I25829,I25846,I25352,I25877,I25346,I25908,I25340,I25972_rst,I25989,I26006,I26023,I26040,I25940,I26071,I26088,I26105,I26122,I26139,I26156,I26173,I26190,I25946,I25937,I26235,I26252,I25961,I26283,I26300,I25949,I26331,I26348,I25955,I26379,I25943,I26410,I25934,I26441,I26458,I25964,I26489,I25958,I26520,I25952,I26584_rst,I26601,I26618,I26635,I26573,I26666,I26683,I26700,I26717,I26734,I26751,I26768,I26558,I26799,I26555,I26830,I26567,I26861,I26878,I26895,I26561,I26576,I26940,I26957,I26546,I26988,I26564,I27019,I27036,I26570,I27067,I27084,I26549,I26552,I27162_rst,I27179,I27196,I27213,I27230,I27247,I27145,I27278,I27295,I27312,I27148,I27130,I27357,I27374,I27391,I27151,I27142,I27436,I27453,I27470,I27133,I27501,I27518,I27124,I27549,I27566,I27583,I27154,I27614,I27631,I27648,I27665,I27139,I27136,I27127,I27757_rst,I27774,I27791,I27808,I27825,I27842,I27740,I27873,I27890,I27907,I27743,I27725,I27952,I27969,I27986,I27746,I27737,I28031,I28048,I28065,I27728,I28096,I28113,I27719,I28144,I28161,I28178,I27749,I28209,I28226,I28243,I28260,I27734,I27731,I27722,I28352_rst,I28369,I28386,I28403,I28420,I28437,I28454,I28323,I28485,I28502,I28519,I28536,I28553,I28570,I28587,I28320,I28314,I28632,I28649,I28666,I28341,I28697,I28714,I28332,I28326,I28759,I28329,I28790,I28807,I28344,I28838,I28338,I28335,I28883,I28317,I28947_rst,I28964,I28981,I28998,I29015,I29032,I29049,I28918,I29080,I29097,I29114,I29131,I29148,I29165,I29182,I28915,I28909,I29227,I29244,I29261,I28936,I29292,I29309,I28927,I28921,I29354,I28924,I29385,I29402,I28939,I29433,I28933,I28930,I29478,I28912,I29542_rst,I29559,I29576,I29593,I29610,I29627,I29644,I29513,I29675,I29692,I29709,I29726,I29743,I29760,I29777,I29510,I29504,I29822,I29839,I29856,I29531,I29887,I29904,I29522,I29516,I29949,I29519,I29980,I29997,I29534,I30028,I29528,I29525,I30073,I29507,I30137_rst,I30154,I30171,I30188,I30205,I30222,I30239,I30108,I30270,I30287,I30304,I30321,I30338,I30355,I30372,I30105,I30099,I30417,I30434,I30451,I30126,I30482,I30499,I30117,I30111,I30544,I30114,I30575,I30592,I30129,I30623,I30123,I30120,I30668,I30102,I30732_rst,I30749,I30766,I30783,I30800,I30817,I30834,I30851,I30868,I30885,I30902,I30919,I30936,I30953,I30721,I30984,I31001,I31018,I30694,I31049,I30715,I31080,I31097,I30700,I31128,I30697,I30703,I31173,I31190,I31207,I30709,I30724,I30712,I31266,I31283,I30718,I30706,I31361_rst,I31378,I31395,I31412,I31429,I31446,I31463,I31480,I31497,I31514,I31531,I31548,I31565,I31582,I31350,I31613,I31630,I31647,I31323,I31678,I31344,I31709,I31726,I31329,I31757,I31326,I31332,I31802,I31819,I31836,I31338,I31353,I31341,I31895,I31912,I31347,I31335,I31990_rst,I32007,I32024,I32041,I32058,I32075,I32092,I32109,I32126,I32143,I32160,I32177,I32194,I32211,I31979,I32242,I32259,I32276,I31952,I32307,I31973,I32338,I32355,I31958,I32386,I31955,I31961,I32431,I32448,I32465,I31967,I31982,I31970,I32524,I32541,I31976,I31964,I32619_rst,I32636,I32653,I32670,I32687,I32704,I32721,I32738,I32755,I32772,I32789,I32806,I32823,I32840,I32608,I32871,I32888,I32905,I32581,I32936,I32602,I32967,I32984,I32587,I33015,I32584,I32590,I33060,I33077,I33094,I32596,I32611,I32599,I33153,I33170,I32605,I32593,I33248_rst,I33265,I33282,I33299,I33316,I33333,I33350,I33367,I33384,I33401,I33418,I33435,I33452,I33469,I33237,I33500,I33517,I33534,I33210,I33565,I33231,I33596,I33613,I33216,I33644,I33213,I33219,I33689,I33706,I33723,I33225,I33240,I33228,I33782,I33799,I33234,I33222,I33877_rst,I33894,I33911,I33928,I33866,I33959,I33854,I33990,I34007,I34024,I34041,I34058,I33857,I34089,I33842,I34120,I34137,I34154,I34171,I34188,I34205,I33848,I34236,I34253,I34270,I33860,I33869,I33839,I34329,I33863,I33851,I34374,I34391,I33845,I34455_rst,I34472,I34489,I34506,I34444,I34537,I34432,I34568,I34585,I34602,I34619,I34636,I34435,I34667,I34420,I34698,I34715,I34732,I34749,I34766,I34783,I34426,I34814,I34831,I34848,I34438,I34447,I34417,I34907,I34441,I34429,I34952,I34969,I34423,I35033_rst,I35050,I35067,I35084,I35022,I35115,I35010,I35146,I35163,I35180,I35197,I35214,I35013,I35245,I34998,I35276,I35293,I35310,I35327,I35344,I35361,I35004,I35392,I35409,I35426,I35016,I35025,I34995,I35485,I35019,I35007,I35530,I35547,I35001,I35611_rst,I35628,I35645,I35662,I35600,I35693,I35588,I35724,I35741,I35758,I35775,I35792,I35591,I35823,I35576,I35854,I35871,I35888,I35905,I35922,I35939,I35582,I35970,I35987,I36004,I35594,I35603,I35573,I36063,I35597,I35585,I36108,I36125,I35579,I36189_rst,I36206,I36223,I36240,I36178,I36271,I36166,I36302,I36319,I36336,I36353,I36370,I36169,I36401,I36154,I36432,I36449,I36466,I36483,I36500,I36517,I36160,I36548,I36565,I36582,I36172,I36181,I36151,I36641,I36175,I36163,I36686,I36703,I36157,I36767_rst,I36784,I36801,I36818,I36756,I36849,I36744,I36880,I36897,I36914,I36931,I36948,I36747,I36979,I36732,I37010,I37027,I37044,I37061,I37078,I37095,I36738,I37126,I37143,I37160,I36750,I36759,I36729,I37219,I36753,I36741,I37264,I37281,I36735,I37345_rst,I37362,I37379,I37396,I37413,I37430,I37328,I37316,I37475,I37492,I37509,I37526,I37543,I37325,I37574,I37591,I37608,I37625,I37334,I37313,I37670,I37687,I37331,I37718,I37322,I37337,I37763,I37780,I37797,I37814,I37310,I37319,I37307,I37906_rst,I37923,I37940,I37957,I37974,I37991,I37889,I37877,I38036,I38053,I38070,I38087,I38104,I37886,I38135,I38152,I38169,I38186,I37895,I37874,I38231,I38248,I37892,I38279,I37883,I37898,I38324,I38341,I38358,I38375,I37871,I37880,I37868,I38467_rst,I38484,I38501,I38518,I38535,I38552,I38450,I38438,I38597,I38614,I38631,I38648,I38665,I38447,I38696,I38713,I38730,I38747,I38456,I38435,I38792,I38809,I38453,I38840,I38444,I38459,I38885,I38902,I38919,I38936,I38432,I38441,I38429,I39028_rst,I39045,I39062,I39079,I39096,I39113,I39011,I38999,I39158,I39175,I39192,I39209,I39226,I39008,I39257,I39274,I39291,I39308,I39017,I38996,I39353,I39370,I39014,I39401,I39005,I39020,I39446,I39463,I39480,I39497,I38993,I39002,I38990,I39589_rst,I39606,I39623,I39640,I39563,I39671,I39688,I39578,I39560,I39733,I39750,I39767,I39784,I39801,I39818,I39835,I39852,I39869,I39575,I39900,I39917,I39934,I39557,I39965,I39554,I39996,I40013,I40030,I40047,I39569,I40078,I39566,I40109,I40126,I40143,I39572,I39581,I39551,I40235_rst,I40252,I40269,I40286,I40209,I40317,I40334,I40224,I40206,I40379,I40396,I40413,I40430,I40447,I40464,I40481,I40498,I40515,I40221,I40546,I40563,I40580,I40203,I40611,I40200,I40642,I40659,I40676,I40693,I40215,I40724,I40212,I40755,I40772,I40789,I40218,I40227,I40197,I40881_rst,I40898,I40915,I40932,I40855,I40963,I40980,I40870,I40852,I41025,I41042,I41059,I41076,I41093,I41110,I41127,I41144,I41161,I40867,I41192,I41209,I41226,I40849,I41257,I40846,I41288,I41305,I41322,I41339,I40861,I41370,I40858,I41401,I41418,I41435,I40864,I40873,I40843,I41527_rst,I41544,I41561,I41578,I41501,I41609,I41626,I41516,I41498,I41671,I41688,I41705,I41722,I41739,I41756,I41773,I41790,I41807,I41513,I41838,I41855,I41872,I41495,I41903,I41492,I41934,I41951,I41968,I41985,I41507,I42016,I41504,I42047,I42064,I42081,I41510,I41519,I41489,I42173_rst,I42190,I42207,I42224,I42147,I42255,I42272,I42162,I42144,I42317,I42334,I42351,I42368,I42385,I42402,I42419,I42436,I42453,I42159,I42484,I42501,I42518,I42141,I42549,I42138,I42580,I42597,I42614,I42631,I42153,I42662,I42150,I42693,I42710,I42727,I42156,I42165,I42135,I42819_rst,I42836,I42853,I42870,I42793,I42901,I42918,I42808,I42790,I42963,I42980,I42997,I43014,I43031,I43048,I43065,I43082,I43099,I42805,I43130,I43147,I43164,I42787,I43195,I42784,I43226,I43243,I43260,I43277,I42799,I43308,I42796,I43339,I43356,I43373,I42802,I42811,I42781,I43465_rst,I43482,I43499,I43516,I43439,I43547,I43564,I43454,I43436,I43609,I43626,I43643,I43660,I43677,I43694,I43711,I43728,I43745,I43451,I43776,I43793,I43810,I43433,I43841,I43430,I43872,I43889,I43906,I43923,I43445,I43954,I43442,I43985,I44002,I44019,I43448,I43457,I43427,I44111_rst,I44128,I44145,I44162,I44085,I44193,I44210,I44100,I44082,I44255,I44272,I44289,I44306,I44323,I44340,I44357,I44374,I44391,I44097,I44422,I44439,I44456,I44079,I44487,I44076,I44518,I44535,I44552,I44569,I44091,I44600,I44088,I44631,I44648,I44665,I44094,I44103,I44073,I44757_rst,I44774,I44791,I44808,I44728,I44839,I44856,I44873,I44890,I44907,I44924,I44941,I44958,I44975,I44992,I44743,I44740,I45037,I44725,I45068,I44722,I45099,I45116,I45133,I45150,I45167,I45184,I44749,I45215,I44737,I44731,I45260,I45277,I44746,I45308,I45325,I45342,I44734,I44719,I45420_rst,I45437,I45454,I45471,I45391,I45502,I45519,I45536,I45553,I45570,I45587,I45604,I45621,I45638,I45655,I45406,I45403,I45700,I45388,I45731,I45385,I45762,I45779,I45796,I45813,I45830,I45847,I45412,I45878,I45400,I45394,I45923,I45940,I45409,I45971,I45988,I46005,I45397,I45382,I46083_rst,I46100,I46117,I46134,I46054,I46165,I46182,I46199,I46216,I46233,I46250,I46267,I46284,I46301,I46318,I46069,I46066,I46363,I46051,I46394,I46048,I46425,I46442,I46459,I46476,I46493,I46510,I46075,I46541,I46063,I46057,I46586,I46603,I46072,I46634,I46651,I46668,I46060,I46045,I46746_rst,I46763,I46780,I46720,I46811,I46828,I46845,I46862,I46879,I46896,I46913,I46930,I46947,I46714,I46978,I46995,I46711,I47026,I47043,I47060,I46723,I46708,I47105,I47122,I47139,I47156,I47173,I46729,I47204,I46738,I47235,I46732,I46735,I46726,I46717,I47341_rst,I47358,I47375,I47315,I47406,I47423,I47440,I47457,I47474,I47491,I47508,I47525,I47542,I47309,I47573,I47590,I47306,I47621,I47638,I47655,I47318,I47303,I47700,I47717,I47734,I47751,I47768,I47324,I47799,I47333,I47830,I47327,I47330,I47321,I47312,I47936_rst,I47953,I47970,I47910,I48001,I48018,I48035,I48052,I48069,I48086,I48103,I48120,I48137,I47904,I48168,I48185,I47901,I48216,I48233,I48250,I47913,I47898,I48295,I48312,I48329,I48346,I48363,I47919,I48394,I47928,I48425,I47922,I47925,I47916,I47907,I48531_rst,I48548,I48565,I48505,I48596,I48613,I48630,I48647,I48664,I48681,I48698,I48715,I48732,I48499,I48763,I48780,I48496,I48811,I48828,I48845,I48508,I48493,I48890,I48907,I48924,I48941,I48958,I48514,I48989,I48523,I49020,I48517,I48520,I48511,I48502,I49126_rst,I49143,I49109,I49088,I49188,I49205,I49222,I49239,I49256,I49273,I49290,I49307,I49324,I49115,I49355,I49372,I49389,I49406,I49118,I49437,I49454,I49471,I49488,I49505,I49103,I49536,I49553,I49106,I49100,I49094,I49612,I49112,I49643,I49097,I49091,I49721_rst,I49738,I49755,I49772,I49789,I49806,I49823,I49840,I49710,I49871,I49695,I49902,I49919,I49936,I49953,I49970,I49987,I50004,I49692,I50035,I50052,I49689,I50083,I50100,I49707,I50131,I49704,I50162,I50179,I49683,I49686,I50224,I50241,I50258,I50275,I49713,I50306,I49698,I49701,I50384_rst,I50401,I50418,I50435,I50452,I50469,I50486,I50503,I50373,I50534,I50358,I50565,I50582,I50599,I50616,I50633,I50650,I50667,I50355,I50698,I50715,I50352,I50746,I50763,I50370,I50794,I50367,I50825,I50842,I50346,I50349,I50887,I50904,I50921,I50938,I50376,I50969,I50361,I50364,I51047_rst,I51064,I51081,I51098,I51115,I51132,I51149,I51166,I51036,I51197,I51021,I51228,I51245,I51262,I51279,I51296,I51313,I51330,I51018,I51361,I51378,I51015,I51409,I51426,I51033,I51457,I51030,I51488,I51505,I51009,I51012,I51550,I51567,I51584,I51601,I51039,I51632,I51024,I51027,I51710_rst,I51727,I51744,I51761,I51778,I51795,I51812,I51829,I51699,I51860,I51684,I51891,I51908,I51925,I51942,I51959,I51976,I51993,I51681,I52024,I52041,I51678,I52072,I52089,I51696,I52120,I51693,I52151,I52168,I51672,I51675,I52213,I52230,I52247,I52264,I51702,I52295,I51687,I51690,I52373_rst,I52390,I52407,I52424,I52441,I52458,I52475,I52492,I52362,I52523,I52347,I52554,I52571,I52588,I52605,I52622,I52639,I52656,I52344,I52687,I52704,I52341,I52735,I52752,I52359,I52783,I52356,I52814,I52831,I52335,I52338,I52876,I52893,I52910,I52927,I52365,I52958,I52350,I52353,I53036_rst,I53053,I53070,I53087,I53104,I53121,I53138,I53155,I53025,I53186,I53010,I53217,I53234,I53251,I53268,I53285,I53302,I53319,I53007,I53350,I53367,I53004,I53398,I53415,I53022,I53446,I53019,I53477,I53494,I52998,I53001,I53539,I53556,I53573,I53590,I53028,I53621,I53013,I53016,I53699_rst,I53716,I53733,I53750,I53767,I53784,I53801,I53818,I53688,I53849,I53673,I53880,I53897,I53914,I53931,I53948,I53965,I53982,I53670,I54013,I54030,I53667,I54061,I54078,I53685,I54109,I53682,I54140,I54157,I53661,I53664,I54202,I54219,I54236,I54253,I53691,I54284,I53676,I53679,I54362_rst,I54379,I54396,I54413,I54430,I54447,I54464,I54481,I54351,I54512,I54336,I54543,I54560,I54577,I54594,I54611,I54628,I54645,I54333,I54676,I54693,I54330,I54724,I54741,I54348,I54772,I54345,I54803,I54820,I54324,I54327,I54865,I54882,I54899,I54916,I54354,I54947,I54339,I54342,I55025_rst,I55042,I55059,I55076,I55093,I55110,I55127,I55144,I55014,I55175,I54999,I55206,I55223,I55240,I55257,I55274,I55291,I55308,I54996,I55339,I55356,I54993,I55387,I55404,I55011,I55435,I55008,I55466,I55483,I54987,I54990,I55528,I55545,I55562,I55579,I55017,I55610,I55002,I55005,I55688_rst,I55705,I55722,I55739,I55756,I55773,I55790,I55807,I55677,I55838,I55662,I55869,I55886,I55903,I55920,I55937,I55954,I55971,I55659,I56002,I56019,I55656,I56050,I56067,I55674,I56098,I55671,I56129,I56146,I55650,I55653,I56191,I56208,I56225,I56242,I55680,I56273,I55665,I55668,I56351_rst,I56368,I56385,I56402,I56419,I56436,I56453,I56322,I56484,I56501,I56518,I56535,I56552,I56569,I56586,I56319,I56617,I56313,I56648,I56665,I56682,I56343,I56316,I56727,I56340,I56758,I56337,I56334,I56803,I56820,I56837,I56854,I56871,I56328,I56902,I56919,I56331,I56325,I56997_rst,I57014,I57031,I57048,I57065,I57082,I57099,I56968,I57130,I57147,I57164,I57181,I57198,I57215,I57232,I56965,I57263,I56959,I57294,I57311,I57328,I56989,I56962,I57373,I56986,I57404,I56983,I56980,I57449,I57466,I57483,I57500,I57517,I56974,I57548,I57565,I56977,I56971,I57643_rst,I57660,I57677,I57694,I57711,I57728,I57745,I57614,I57776,I57793,I57810,I57827,I57844,I57861,I57878,I57611,I57909,I57605,I57940,I57957,I57974,I57635,I57608,I58019,I57632,I58050,I57629,I57626,I58095,I58112,I58129,I58146,I58163,I57620,I58194,I58211,I57623,I57617,I58289_rst,I58306,I58323,I58340,I58357,I58374,I58391,I58260,I58422,I58439,I58456,I58473,I58490,I58507,I58524,I58257,I58555,I58251,I58586,I58603,I58620,I58281,I58254,I58665,I58278,I58696,I58275,I58272,I58741,I58758,I58775,I58792,I58809,I58266,I58840,I58857,I58269,I58263,I58935_rst,I58952,I58969,I58986,I59003,I59020,I59037,I58906,I59068,I59085,I59102,I59119,I59136,I59153,I59170,I58903,I59201,I58897,I59232,I59249,I59266,I58927,I58900,I59311,I58924,I59342,I58921,I58918,I59387,I59404,I59421,I59438,I59455,I58912,I59486,I59503,I58915,I58909,I59581_rst,I59598,I59615,I59632,I59649,I59666,I59683,I59552,I59714,I59731,I59748,I59765,I59782,I59799,I59816,I59549,I59847,I59543,I59878,I59895,I59912,I59573,I59546,I59957,I59570,I59988,I59567,I59564,I60033,I60050,I60067,I60084,I60101,I59558,I60132,I60149,I59561,I59555,I60227_rst,I60244,I60261,I60278,I60295,I60312,I60329,I60198,I60360,I60377,I60394,I60411,I60428,I60445,I60462,I60195,I60493,I60189,I60524,I60541,I60558,I60219,I60192,I60603,I60216,I60634,I60213,I60210,I60679,I60696,I60713,I60730,I60747,I60204,I60778,I60795,I60207,I60201,I60873_rst,I60890,I60907,I60924,I60941,I60958,I60975,I60844,I61006,I61023,I61040,I61057,I61074,I61091,I61108,I60841,I61139,I60835,I61170,I61187,I61204,I60865,I60838,I61249,I60862,I61280,I60859,I60856,I61325,I61342,I61359,I61376,I61393,I60850,I61424,I61441,I60853,I60847,I61519_rst,I61536,I61553,I61570,I61587,I61604,I61621,I61490,I61652,I61669,I61686,I61703,I61720,I61737,I61754,I61487,I61785,I61481,I61816,I61833,I61850,I61511,I61484,I61895,I61508,I61926,I61505,I61502,I61971,I61988,I62005,I62022,I62039,I61496,I62070,I62087,I61499,I61493,I62165_rst,I62182,I62199,I62216,I62233,I62250,I62267,I62136,I62298,I62315,I62332,I62349,I62366,I62383,I62400,I62133,I62431,I62127,I62462,I62479,I62496,I62157,I62130,I62541,I62154,I62572,I62151,I62148,I62617,I62634,I62651,I62668,I62685,I62142,I62716,I62733,I62145,I62139,I62811_rst,I62828,I62845,I62862,I62879,I62896,I62913,I62782,I62944,I62961,I62978,I62995,I63012,I63029,I63046,I62779,I63077,I62773,I63108,I63125,I63142,I62803,I62776,I63187,I62800,I63218,I62797,I62794,I63263,I63280,I63297,I63314,I63331,I62788,I63362,I63379,I62791,I62785,I63457_rst,I63474,I63491,I63508,I63525,I63542,I63559,I63428,I63590,I63607,I63624,I63641,I63658,I63675,I63692,I63425,I63723,I63419,I63754,I63771,I63788,I63449,I63422,I63833,I63446,I63864,I63443,I63440,I63909,I63926,I63943,I63960,I63977,I63434,I64008,I64025,I63437,I63431,I64103_rst,I64120,I64137,I64154,I64171,I64188,I64205,I64074,I64236,I64253,I64270,I64287,I64304,I64321,I64338,I64071,I64369,I64065,I64400,I64417,I64434,I64095,I64068,I64479,I64092,I64510,I64089,I64086,I64555,I64572,I64589,I64606,I64623,I64080,I64654,I64671,I64083,I64077,I64749_rst,I64766,I64783,I64800,I64817,I64834,I64851,I64720,I64882,I64899,I64916,I64933,I64950,I64967,I64984,I64717,I65015,I64711,I65046,I65063,I65080,I64741,I64714,I65125,I64738,I65156,I64735,I64732,I65201,I65218,I65235,I65252,I65269,I64726,I65300,I65317,I64729,I64723,I65395_rst,I65412,I65429,I65446,I65463,I65357,I65494,I65511,I65528,I65545,I65562,I65579,I65366,I65610,I65360,I65641,I65658,I65675,I65692,I65387,I65384,I65737,I65754,I65771,I65381,I65802,I65378,I65369,I65847,I65864,I65881,I65372,I65375,I65926,I65943,I65363,I66007_rst,I66024,I66041,I66058,I66075,I65969,I66106,I66123,I66140,I66157,I66174,I66191,I65978,I66222,I65972,I66253,I66270,I66287,I66304,I65999,I65996,I66349,I66366,I66383,I65993,I66414,I65990,I65981,I66459,I66476,I66493,I65984,I65987,I66538,I66555,I65975,I66619_rst,I66636,I66653,I66670,I66687,I66587,I66718,I66735,I66752,I66590,I66783,I66584,I66814,I66831,I66848,I66865,I66882,I66593,I66913,I66930,I66947,I66964,I66599,I66602,I66581,I67023,I67040,I67057,I66611,I66608,I67102,I67119,I66596,I66605,I67197_rst,I67214,I67231,I67248,I67265,I67165,I67296,I67313,I67330,I67168,I67361,I67162,I67392,I67409,I67426,I67443,I67460,I67171,I67491,I67508,I67525,I67542,I67177,I67180,I67159,I67601,I67618,I67635,I67189,I67186,I67680,I67697,I67174,I67183,I67775_rst,I67792,I67809,I67826,I67843,I67743,I67874,I67891,I67908,I67746,I67939,I67740,I67970,I67987,I68004,I68021,I68038,I67749,I68069,I68086,I68103,I68120,I67755,I67758,I67737,I68179,I68196,I68213,I67767,I67764,I68258,I68275,I67752,I67761,I68353_rst,I68370,I68387,I68404,I68421,I68321,I68452,I68469,I68486,I68324,I68517,I68318,I68548,I68565,I68582,I68599,I68616,I68327,I6864_rst7,I68664,I68681,I68698,I68333,I68336,I68315,I68757,I68774,I68791,I68345,I68342,I68836,I68853,I68330,I68339,I68931_rst,I68948,I68965,I68982,I68999,I68899,I69030,I69047,I69064,I68902,I69095,I68896,I69126,I69143,I69160,I69177,I69194,I68905,I69225,I69242,I69259,I69276,I68911,I68914,I68893,I69335,I69352,I69369,I68923,I68920,I69414,I69431,I68908,I68917,I69509_rst,I69526,I69543,I69560,I69577,I69477,I69608,I69625,I69642,I69480,I69673,I69474,I69704,I69721,I69738,I69755,I69772,I69483,I69803,I69820,I69837,I69854,I69489,I69492,I69471,I69913,I69930,I69947,I69501,I69498,I69992,I70009,I69486,I69495,I70087_rst,I70104,I70121,I70138,I70155,I70055,I70186,I70203,I70220,I70058,I70251,I70052,I70282,I70299,I70316,I70333,I70350,I70061,I70381,I70398,I70415,I70432,I70067,I70070,I70049,I70491,I70508,I70525,I70079,I70076,I70570,I70587,I70064,I70073,I70665_rst,I70682,I70699,I70716,I70733,I70633,I70764,I70781,I70798,I70636,I70829,I70630,I70860,I70877,I70894,I70911,I70928,I70639,I70959,I70976,I70993,I71010,I70645,I70648,I70627,I71069,I71086,I71103,I70657,I70654,I71148,I71165,I70642,I70651,I71243_rst,I71260,I71277,I71294,I71311,I71211,I71342,I71359,I71376,I71214,I71407,I71208,I71438,I71455,I71472,I71489,I71506,I71217,I71537,I71554,I71571,I71588,I71223,I71226,I71205,I71647,I71664,I71681,I71235,I71232,I71726,I71743,I71220,I71229,I71821_rst,I71838,I71855,I71872,I71889,I71789,I71920,I71937,I71954,I71971,I71988,I72005,I72022,I72039,I71795,I71786,I72084,I72101,I71810,I72132,I72149,I71798,I72180,I72197,I71804,I72228,I71792,I72259,I71783,I72290,I72307,I71813,I72338,I71807,I72369,I71801,I72433_rst,I72450,I72467,I72484,I72501,I72518,I72416,I72549,I72566,I72583,I72419,I72401,I72628,I72645,I72662,I72422,I72413,I72707,I72724,I72741,I72404,I72772,I72789,I72395,I72820,I72837,I72854,I72425,I72885,I72902,I72919,I72936,I72410,I72407,I72398,I73028_rst,I73045,I73062,I73079,I73096,I73113,I73011,I73144,I73161,I73178,I73014,I72996,I73223,I73240,I73257,I73017,I73008,I73302,I73319,I73336,I72999,I73367,I73384,I72990,I73415,I73432,I73449,I73020,I73480,I73497,I73514,I73531,I73005,I73002,I72993,I73623_rst,I73640,I73657,I73674,I73691,I73708,I73606,I73739,I73756,I73773,I73609,I73591,I73818,I73835,I73852,I73612,I73603,I73897,I73914,I73931,I73594,I73962,I73979,I73585,I74010,I74027,I74044,I73615,I74075,I74092,I74109,I74126,I73600,I73597,I73588,I74218_rst,I74235,I74252,I74269,I74286,I74303,I74201,I74334,I74351,I74368,I74204,I74186,I74413,I74430,I74447,I74207,I74198,I74492,I74509,I74526,I74189,I74557,I74574,I74180,I74605,I74622,I74639,I74210,I74670,I74687,I74704,I74721,I74195,I74192,I74183,I74813_rst,I74830,I74847,I74864,I74881,I74898,I74796,I74929,I74946,I74963,I74799,I74781,I75008,I75025,I75042,I74802,I74793,I75087,I7510_rst4,I75121,I74784,I75152,I75169,I74775,I75200,I75217,I75234,I74805,I75265,I75282,I75299,I75316,I74790,I74787,I74778,I75408_rst,I75425,I75442,I75459,I75476,I75493,I75391,I75524,I75541,I75558,I75394,I75376,I75603,I75620,I75637,I75397,I75388,I75682,I75699,I75716,I75379,I75747,I75764,I75370,I75795,I75812,I75829,I75400,I75860,I75877,I75894,I75911,I75385,I75382,I75373,I76003_rst,I76020,I76037,I76054,I76071,I76088,I75986,I76119,I76136,I76153,I75989,I75971,I76198,I76215,I76232,I75992,I75983,I76277,I76294,I76311,I75974,I76342,I76359,I75965,I76390,I76407,I76424,I75995,I76455,I76472,I76489,I76506,I75980,I75977,I75968,I76598_rst,I76615,I76632,I76649,I76666,I76683,I76581,I76714,I76731,I76748,I76584,I76566,I76793,I76810,I76827,I76587,I76578,I76872,I76889,I76906,I76569,I76937,I76954,I76560,I76985,I77002,I77019,I76590,I77050,I77067,I77084,I77101,I76575,I76572,I76563,I77193_rst,I77210,I77227,I77244,I77261,I77278,I77295,I77164,I77326,I77343,I77360,I77377,I77394,I77411,I77428,I77161,I77155,I77473,I77490,I77507,I77182,I77538,I77555,I77173,I77167,I77600,I77170,I77631,I77648,I77185,I77679,I77179,I77176,I77724,I77158,I77788_rst,I77805,I77822,I77839,I77856,I77873,I77890,I77759,I77921,I77938,I77955,I77972,I77989,I78006,I78023,I77756,I77750,I78068,I78085,I78102,I77777,I78133,I78150,I77768,I77762,I78195,I77765,I78226,I78243,I77780,I78274,I77774,I77771,I78319,I77753,I78383_rst,I78400,I78417,I78434,I78451,I78468,I78485,I78354,I78516,I78533,I78550,I78567,I78584,I78601,I78618,I78351,I78345,I78663,I78680,I78697,I78372,I78728,I78745,I78363,I78357,I78790,I78360,I78821,I78838,I78375,I78869,I78369,I78366,I78914,I78348,I78978_rst,I78995,I79012,I79029,I79046,I79063,I79080,I78949,I79111,I79128,I79145,I79162,I79179,I79196,I79213,I78946,I78940,I79258,I79275,I79292,I78967,I79323,I79340,I78958,I78952,I79385,I78955,I79416,I79433,I78970,I79464,I78964,I78961,I79509,I78943,I79573_rst,I79590,I79607,I79624,I79641,I79658,I79675,I79544,I79706,I79723,I79740,I79757,I79774,I79791,I79808,I79541,I79535,I79853,I79870,I79887,I79562,I79918,I79935,I79553,I79547,I79980,I79550,I80011,I80028,I79565,I80059,I79559,I79556,I80104,I79538,I80168_rst,I80185,I80202,I80219,I80236,I80253,I80270,I80139,I80301,I80318,I80335,I80352,I80369,I80386,I80403,I80136,I80130,I80448,I80465,I80482,I80157,I80513,I80530,I80148,I80142,I80575,I80145,I80606,I80623,I80160,I80654,I80154,I80151,I80699,I80133,I80763_rst,I80780,I80797,I80814,I80831,I80848,I80865,I80734,I80896,I80913,I80930,I80947,I80964,I80981,I80998,I80731,I80725,I81043,I81060,I81077,I80752,I81108,I81125,I80743,I80737,I81170,I80740,I81201,I81218,I80755,I81249,I80749,I80746,I81294,I80728,I81358_rst,I81375,I81392,I81409,I81426,I81443,I81460,I81329,I81491,I81508,I81525,I81542,I81559,I81576,I81593,I81326,I81320,I81638,I81655,I81672,I81347,I81703,I81720,I81338,I81332,I81765,I81335,I81796,I81813,I81350,I81844,I81344,I81341,I81889,I81323,I81953_rst,I81970,I81987,I82004,I82021,I82038,I82055,I81924,I82086,I82103,I82120,I82137,I82154,I82171,I82188,I81921,I81915,I82233,I82250,I82267,I81942,I82298,I82315,I81933,I81927,I82360,I81930,I82391,I82408,I81945,I82439,I81939,I81936,I82484,I81918,I82548_rst,I82565,I82582,I82599,I82616,I82633,I82650,I82667,I82684,I82701,I82718,I82735,I82752,I82769,I82537,I82800,I82817,I82834,I82510,I82865,I82531,I82896,I82913,I82516,I82944,I82513,I82519,I82989,I83006,I83023,I82525,I82540,I82528,I83082,I83099,I82534,I82522,I83177_rst,I83194,I83211,I83228,I83245,I83262,I83279,I83296,I83313,I83330,I83347,I83364,I83381,I83398,I83166,I83429,I83446,I83463,I83139,I83494,I83160,I83525,I83542,I83145,I83573,I83142,I83148,I83618,I83635,I83652,I83154,I83169,I83157,I83711,I83728,I83163,I83151,I83806_rst,I83823,I83840,I83857,I83874,I83891,I83908,I83925,I83942,I83959,I83976,I83993,I84010,I84027,I83795,I84058,I84075,I84092,I83768,I84123,I83789,I84154,I84171,I83774,I84202,I83771,I83777,I84247,I84264,I84281,I83783,I83798,I83786,I84340,I84357,I83792,I83780,I84435_rst,I84452,I84469,I84486,I84503,I84520,I84537,I84554,I84571,I84588,I84605,I84622,I84639,I84656,I84424,I84687,I84704,I84721,I84397,I84752,I84418,I84783,I84800,I84403,I84831,I84400,I84406,I84876,I84893,I84910,I84412,I84427,I84415,I84969,I84986,I84421,I84409,I85064_rst,I85081,I85098,I85115,I85132,I85149,I85166,I85183,I85200,I85217,I85234,I85251,I85268,I85285,I85053,I85316,I85333,I85350,I85026,I85381,I85047,I85412,I85429,I85032,I85460,I85029,I85035,I85505,I85522,I85539,I85041,I85056,I85044,I85598,I85615,I85050,I85038,I85693_rst,I85710,I85727,I85744,I85761,I85778,I85795,I85812,I85829,I85846,I85863,I85880,I85897,I85914,I85682,I85945,I85962,I85979,I85655,I86010,I85676,I86041,I86058,I85661,I86089,I85658,I85664,I86134,I86151,I86168,I85670,I85685,I85673,I86227,I86244,I85679,I85667,I86322_rst,I86339,I86356,I86373,I86390,I86407,I86424,I86441,I86458,I86475,I86492,I86509,I86526,I86543,I86311,I86574,I86591,I86608,I86284,I86639,I86305,I86670,I86687,I86290,I86718,I86287,I86293,I86763,I86780,I86797,I86299,I86314,I86302,I86856,I86873,I86308,I86296,I86951_rst,I86968,I86985,I87002,I87019,I87036,I87053,I87070,I87087,I87104,I87121,I87138,I87155,I87172,I86940,I87203,I87220,I87237,I86913,I87268,I86934,I87299,I87316,I86919,I87347,I86916,I86922,I87392,I87409,I87426,I86928,I86943,I86931,I87485,I87502,I86937,I86925,I87580_rst,I87597,I87614,I87631,I87648,I87665,I87682,I87699,I87716,I87733,I87750,I87767,I87784,I87801,I87569,I87832,I87849,I87866,I87542,I87897,I87563,I87928,I87945,I87548,I87976,I87545,I87551,I88021,I88038,I88055,I87557,I87572,I87560,I88114,I88131,I87566,I87554,I88209_rst,I88226,I88243,I88260,I88277,I88294,I88311,I88328,I88345,I8836_rst2,I88379,I88396,I88413,I88430,I88198,I88461,I88478,I88495,I88171,I88526,I88192,I88557,I88574,I88177,I88605,I88174,I88180,I88650,I88667,I88684,I88186,I88201,I88189,I88743,I88760,I88195,I88183,I88838_rst,I88855,I88872,I88889,I88906,I88923,I88940,I88957,I88974,I88991,I89008,I89025,I89042,I89059,I88827,I89090,I89107,I89124,I88800,I89155,I88821,I89186,I89203,I88806,I89234,I88803,I88809,I89279,I89296,I89313,I88815,I88830,I88818,I89372,I89389,I88824,I88812,I89467_rst,I89484,I89501,I89518,I89535,I89552,I89569,I89586,I89603,I89620,I89637,I89654,I89671,I89688,I89456,I89719,I89736,I89753,I89429,I89784,I89450,I89815,I89832,I89435,I89863,I89432,I89438,I89908,I89925,I89942,I89444,I89459,I89447,I90001,I90018,I89453,I89441,I90096_rst,I90113,I90130,I90147,I90164,I90181,I90198,I90215,I90232,I90249,I90266,I90283,I90300,I90317,I90085,I90348,I90365,I90382,I90058,I90413,I90079,I90444,I90461,I90064,I90492,I90061,I90067,I90537,I90554,I90571,I90073,I90088,I90076,I90630,I90647,I90082,I90070,I90725_rst,I90742,I90759,I90776,I90714,I90807,I90702,I90838,I90855,I90872,I90889,I90906,I90705,I90937,I90690,I90968,I90985,I91002,I91019,I91036,I91053,I90696,I91084,I91101,I91118,I90708,I90717,I90687,I91177,I90711,I90699,I91222,I91239,I90693,I91303_rst,I91320,I91337,I91354,I91292,I91385,I91280,I91416,I91433,I91450,I91467,I91484,I91283,I91515,I91268,I91546,I91563,I91580,I91597,I91614,I91631,I91274,I91662,I91679,I91696,I91286,I91295,I91265,I91755,I91289,I91277,I91800,I91817,I91271,I91881_rst,I91898,I91915,I91932,I91870,I91963,I91858,I91994,I92011,I92028,I92045,I92062,I91861,I92093,I91846,I92124,I92141,I92158,I92175,I92192,I92209,I91852,I92240,I92257,I92274,I91864,I91873,I91843,I92333,I91867,I91855,I92378,I92395,I91849,I92459_rst,I92476,I92493,I92510,I92448,I92541,I92436,I92572,I92589,I92606,I92623,I92640,I92439,I92671,I92424,I92702,I92719,I92736,I92753,I92770,I92787,I92430,I92818,I92835,I92852,I92442,I92451,I92421,I92911,I92445,I92433,I92956,I92973,I92427,I93037_rst,I93054,I93071,I93088,I93026,I93119,I93014,I93150,I93167,I93184,I93201,I93218,I93017,I93249,I93002,I93280,I93297,I93314,I93331,I93348,I93365,I93008,I93396,I93413,I93430,I93020,I93029,I92999,I93489,I93023,I93011,I93534,I93551,I93005,I93615_rst,I93632,I93649,I93666,I93604,I93697,I93592,I93728,I93745,I93762,I93779,I93796,I93595,I93827,I93580,I93858,I93875,I93892,I93909,I93926,I93943,I93586,I93974,I93991,I94008,I93598,I93607,I93577,I94067,I93601,I93589,I94112,I94129,I93583,I94193_rst,I94210,I94227,I94244,I94182,I94275,I94170,I94306,I94323,I94340,I94357,I94374,I94173,I94405,I94158,I94436,I94453,I94470,I94487,I94504,I94521,I94164,I94552,I94569,I94586,I94176,I94185,I94155,I94645,I94179,I94167,I94690,I94707,I94161,I94771_rst,I94788,I94805,I94822,I94839,I94856,I94754,I94742,I94901,I94918,I94935,I94952,I94969,I94751,I95000,I95017,I95034,I95051,I94760,I94739,I95096,I95113,I94757,I95144,I94748,I94763,I95189,I95206,I95223,I95240,I94736,I94745,I94733,I95332_rst,I95349,I95366,I95383,I95400,I95417,I95315,I95303,I95462,I95479,I95496,I95513,I95530,I95312,I95561,I95578,I95595,I95612,I95321,I95300,I95657,I95674,I95318,I95705,I95309,I95324,I95750,I95767,I95784,I95801,I95297,I95306,I95294,I95893_rst,I95910,I95927,I95944,I95961,I95978,I95876,I95864,I96023,I96040,I96057,I96074,I96091,I95873,I96122,I96139,I96156,I96173,I95882,I95861,I96218,I96235,I95879,I96266,I95870,I95885,I96311,I96328,I96345,I96362,I95858,I95867,I95855,I96454_rst,I96471,I96488,I96505,I96522,I96539,I96437,I96425,I96584,I96601,I96618,I96635,I96652,I96434,I96683,I96700,I96717,I96734,I96443,I96422,I96779,I96796,I96440,I96827,I96431,I96446,I96872,I96889,I96906,I96923,I96419,I96428,I96416,I97015_rst,I97032,I97049,I97066,I97083,I97100,I96998,I96986,I97145,I97162,I97179,I97196,I97213,I96995,I97244,I97261,I97278,I97295,I97004,I96983,I97340,I97357,I97001,I97388,I96992,I97007,I97433,I97450,I97467,I97484,I96980,I96989,I96977,I97576_rst,I97593,I97610,I97627,I97644,I97661,I97559,I97547,I97706,I97723,I97740,I97757,I97774,I97556,I97805,I97822,I97839,I97856,I97565,I97544,I97901,I97918,I97562,I97949,I97553,I97568,I97994,I98011,I98028,I98045,I97541,I97550,I97538,I98137_rst,I98154,I98171,I98188,I98205,I98222,I98120,I98108,I98267,I98284,I98301,I98318,I98335,I98117,I98366,I98383,I98400,I98417,I98126,I98105,I98462,I98479,I98123,I98510,I98114,I98129,I98555,I98572,I98589,I98606,I98102,I98111,I98099,I98698_rst,I98715,I98732,I98749,I98672,I98780,I98797,I98687,I98669,I98842,I98859,I98876,I98893,I98910,I98927,I98944,I98961,I98978,I98684,I99009,I99026,I99043,I98666,I99074,I98663,I99105,I99122,I99139,I99156,I98678,I99187,I98675,I99218,I99235,I99252,I98681,I98690,I98660,I99344_rst,I99361,I99378,I99395,I99318,I99426,I99443,I99333,I99315,I99488,I99505,I99522,I99539,I99556,I99573,I99590,I99607,I99624,I99330,I99655,I99672,I99689,I99312,I99720,I99309,I99751,I99768,I99785,I99802,I99324,I99833,I99321,I99864,I99881,I99898,I99327,I99336,I99306,I99990_rst,I100007,I100024,I100041,I99964,I100072,I100089,I99979,I99961,I100134,I100151,I100168,I100185,I100202,I100219,I100236,I100253,I100270,I99976,I100301,I100318,I100335,I99958,I100366,I99955,I100397,I100414,I100431,I100448,I99970,I100479,I99967,I100510,I100527,I100544,I99973,I99982,I99952,I100636_rst,I100653,I100670,I100687,I100610,I100718,I100735,I100625,I100607,I100780,I100797,I100814,I100831,I100848,I100865,I100882,I100899,I100916,I100622,I100947,I100964,I100981,I100604,I101012,I100601,I101043,I101060,I101077,I101094,I100616,I101125,I100613,I101156,I101173,I101190,I100619,I100628,I100598,I101282_rst,I101299,I101316,I101333,I101256,I101364,I101381,I101271,I101253,I101426,I101443,I101460,I101477,I101494,I101511,I101528,I101545,I101562,I101268,I101593,I101610,I10162_rst7,I101250,I101658,I101247,I101689,I101706,I101723,I101740,I101262,I101771,I101259,I101802,I101819,I101836,I101265,I101274,I101244,I101928_rst,I101945,I101962,I101979,I101902,I102010,I102027,I101917,I101899,I102072,I102089,I102106,I102123,I102140,I102157,I102174,I102191,I102208,I101914,I102239,I102256,I102273,I101896,I102304,I101893,I102335,I102352,I102369,I102386,I101908,I102417,I101905,I102448,I102465,I102482,I101911,I101920,I101890,I102574_rst,I102591,I102608,I102625,I102548,I102656,I102673,I102563,I102545,I102718,I102735,I102752,I102769,I102786,I102803,I102820,I102837,I102854,I102560,I102885,I102902,I102919,I102542,I102950,I102539,I102981,I102998,I103015,I103032,I102554,I103063,I102551,I103094,I103111,I103128,I102557,I102566,I102536,I103220_rst,I103237,I103254,I103271,I103194,I103302,I103319,I103209,I103191,I103364,I103381,I103398,I103415,I103432,I103449,I103466,I103483,I103500,I103206,I103531,I103548,I103565,I103188,I103596,I103185,I103627,I103644,I103661,I103678,I103200,I103709,I103197,I103740,I103757,I103774,I103203,I103212,I103182,I103866_rst,I103883,I103900,I103917,I103840,I103948,I103965,I103855,I103837,I104010,I104027,I104044,I104061,I104078,I104095,I104112,I104129,I104146,I103852,I104177,I104194,I104211,I103834,I104242,I103831,I104273,I104290,I104307,I104324,I103846,I104355,I103843,I104386,I104403,I104420,I103849,I103858,I103828,I104512_rst,I104529,I104546,I104563,I104486,I104594,I104611,I104501,I104483,I104656,I104673,I104690,I104707,I104724,I104741,I104758,I104775,I104792,I104498,I104823,I104840,I104857,I104480,I104888,I104477,I104919,I104936,I104953,I104970,I104492,I105001,I104489,I105032,I105049,I105066,I104495,I104504,I104474,I105158_rst,I105175,I105192,I105209,I105132,I105240,I105257,I105147,I105129,I105302,I105319,I105336,I105353,I105370,I105387,I105404,I105421,I105438,I105144,I105469,I105486,I105503,I105126,I105534,I105123,I105565,I105582,I105599,I105616,I105138,I105647,I105135,I105678,I105695,I105712,I105141,I105150,I105120,I105804_rst,I105821,I105838,I105855,I105778,I105886,I105903,I105793,I105775,I105948,I105965,I105982,I105999,I106016,I106033,I106050,I106067,I106084,I105790,I106115,I106132,I106149,I105772,I106180,I105769,I106211,I106228,I106245,I106262,I105784,I106293,I105781,I106324,I106341,I106358,I105787,I105796,I105766,I106450_rst,I106467,I106484,I106501,I106424,I106532,I106549,I106439,I106421,I106594,I106611,I106628,I106645,I106662,I106679,I106696,I106713,I106730,I106436,I106761,I106778,I106795,I106418,I106826,I106415,I106857,I106874,I106891,I106908,I106430,I106939,I106427,I106970,I106987,I107004,I106433,I106442,I106412,I107096_rst,I107113,I107130,I107147,I107070,I107178,I107195,I107085,I107067,I107240,I107257,I107274,I107291,I107308,I107325,I107342,I107359,I107376,I107082,I107407,I107424,I107441,I107064,I107472,I107061,I107503,I107520,I107537,I107554,I107076,I107585,I107073,I107616,I107633,I107650,I107079,I107088,I107058,I107742_rst,I107759,I107776,I107793,I107713,I107824,I107841,I107858,I107875,I107892,I107909,I107926,I107943,I107960,I107977,I107728,I107725,I108022,I107710,I108053,I107707,I108084,I108101,I108118,I108135,I108152,I108169,I107734,I108200,I107722,I107716,I108245,I108262,I107731,I108293,I108310,I108327,I107719,I107704,I108405_rst,I108422,I108439,I108456,I108376,I108487,I108504,I108521,I108538,I108555,I108572,I108589,I108606,I108623,I108640,I108391,I108388,I108685,I108373,I108716,I108370,I108747,I108764,I108781,I108798,I108815,I108832,I108397,I108863,I108385,I108379,I108908,I108925,I108394,I108956,I108973,I108990,I108382,I108367,I109068_rst,I109085,I109102,I109119,I109039,I109150,I109167,I109184,I109201,I109218,I109235,I109252,I109269,I109286,I109303,I109054,I109051,I109348,I109036,I109379,I109033,I109410,I109427,I109444,I109461,I109478,I109495,I109060,I109526,I109048,I109042,I109571,I109588,I109057,I109619,I109636,I109653,I109045,I109030,I109731_rst,I109748,I109765,I109782,I109702,I109813,I109830,I109847,I109864,I109881,I109898,I109915,I109932,I109949,I109966,I109717,I109714,I110011,I109699,I110042,I109696,I110073,I110090,I110107,I110124,I110141,I110158,I109723,I110189,I109711,I109705,I110234,I110251,I109720,I110282,I110299,I110316,I109708,I109693,I110394_rst,I110411,I110428,I110445,I110365,I110476,I110493,I110510,I110527,I110544,I110561,I110578,I110595,I110612,I110629,I110380,I110377,I110674,I110362,I110705,I110359,I110736,I110753,I110770,I110787,I110804,I110821,I110386,I110852,I110374,I110368,I110897,I110914,I110383,I110945,I110962,I110979,I110371,I110356,I111057_rst,I111074,I111091,I111108,I111028,I111139,I111156,I111173,I111190,I111207,I111224,I111241,I111258,I111275,I111292,I111043,I111040,I111337,I111025,I111368,I111022,I111399,I111416,I111433,I111450,I111467,I111484,I111049,I111515,I111037,I111031,I111560,I111577,I111046,I111608,I111625,I111642,I111034,I111019,I111720_rst,I111737,I111754,I111771,I111691,I111802,I111819,I111836,I111853,I111870,I111887,I111904,I111921,I111938,I111955,I111706,I111703,I112000,I111688,I112031,I111685,I112062,I112079,I112096,I112113,I112130,I112147,I111712,I112178,I111700,I111694,I112223,I112240,I111709,I112271,I112288,I112305,I111697,I111682,I112383_rst,I112400,I112417,I112434,I112354,I112465,I112482,I112499,I112516,I112533,I112550,I112567,I112584,I112601,I112618,I112369,I112366,I112663,I112351,I112694,I112348,I112725,I112742,I112759,I112776,I112793,I112810,I112375,I112841,I112363,I112357,I112886,I112903,I112372,I112934,I112951,I112968,I112360,I112345,I113046_rst,I113063,I113080,I113097,I113017,I113128,I113145,I113162,I113179,I113196,I113213,I113230,I113247,I113264,I113281,I113032,I113029,I113326,I113014,I113357,I113011,I113388,I113405,I113422,I113439,I113456,I113473,I113038,I113504,I113026,I113020,I113549,I113566,I113035,I113597,I113614,I113631,I113023,I113008,I113709_rst,I113726,I113743,I113683,I113774,I113791,I113808,I113825,I113842,I113859,I113876,I113893,I113910,I113677,I113941,I113958,I113674,I113989,I114006,I114023,I113686,I113671,I114068,I114085,I114102,I114119,I114136,I113692,I114167,I113701,I114198,I113695,I113698,I113689,I113680,I114304_rst,I114321,I114338,I114278,I114369,I114386,I114403,I114420,I114437,I114454,I114471,I114488,I114505,I114272,I114536,I114553,I114269,I114584,I114601,I114618,I114281,I114266,I114663,I114680,I114697,I114714,I114731,I114287,I114762,I114296,I114793,I114290,I114293,I114284,I114275,I114899_rst,I114916,I114933,I114873,I114964,I114981,I114998,I115015,I115032,I115049,I115066,I115083,I115100,I114867,I115131,I115148,I114864,I115179,I115196,I115213,I114876,I114861,I115258,I115275,I115292,I115309,I115326,I11488_rst2,I115357,I114891,I115388,I11488_rst5,I11488_rst8,I114879,I114870,I115494_rst,I115511,I115528,I115468,I115559,I115576,I115593,I115610,I115627,I115644,I115661,I115678,I115695,I115462,I115726,I115743,I115459,I115774,I115791,I115808,I115471,I115456,I115853,I115870,I115887,I115904,I115921,I115477,I115952,I115486,I115983,I115480,I115483,I115474,I115465,I116089_rst,I116106,I116123,I116063,I116154,I116171,I116188,I116205,I116222,I116239,I116256,I116273,I116290,I116057,I116321,I116338,I116054,I116369,I116386,I116403,I116066,I116051,I116448,I116465,I116482,I116499,I116516,I116072,I116547,I116081,I116578,I116075,I116078,I116069,I116060,I116684_rst,I116701,I116718,I116658,I116749,I116766,I116783,I116800,I116817,I116834,I116851,I116868,I116885,I116652,I116916,I116933,I116649,I116964,I116981,I116998,I116661,I116646,I117043,I117060,I117077,I117094,I117111,I116667,I117142,I116676,I117173,I116670,I116673,I116664,I116655,I117279_rst,I117296,I117313,I117253,I117344,I117361,I117378,I117395,I117412,I117429,I117446,I117463,I117480,I117247,I117511,I117528,I117244,I117559,I117576,I117593,I117256,I117241,I117638,I117655,I117672,I117689,I117706,I117262,I117737,I117271,I117768,I117265,I117268,I117259,I117250,I117874_rst,I117891,I117908,I117848,I117939,I117956,I117973,I117990,I118007,I118024,I118041,I118058,I118075,I117842,I118106,I118123,I117839,I118154,I118171,I118188,I117851,I117836,I118233,I118250,I118267,I118284,I118301,I117857,I118332,I117866,I118363,I117860,I117863,I117854,I117845,I118469_rst,I118486,I118452,I118431,I118531,I118548,I118565,I118582,I118599,I118616,I118633,I118650,I118667,I118458,I118698,I118715,I118732,I118749,I118461,I118780,I118797,I118814,I118831,I118848,I118446,I118879,I118896,I118449,I118443,I118437,I118955,I118455,I118986,I118440,I118434,I119064_rst,I119081,I119098,I119115,I119132,I119149,I119166,I119183,I119053,I119214,I119038,I119245,I119262,I119279,I119296,I119313,I119330,I119347,I119035,I119378,I119395,I119032,I119426,I119443,I119050,I119474,I119047,I119505,I119522,I119026,I119029,I119567,I119584,I119601,I119618,I119056,I119649,I119041,I119044,I119727_rst,I119744,I119761,I119778,I119795,I119812,I119829,I119846,I119716,I119877,I119701,I119908,I119925,I119942,I119959,I119976,I119993,I120010,I119698,I120041,I120058,I119695,I120089,I120106,I119713,I120137,I119710,I120168,I120185,I119689,I119692,I120230,I120247,I120264,I120281,I119719,I120312,I119704,I119707,I120390_rst,I120407,I120424,I120441,I120458,I120475,I120492,I120509,I120379,I120540,I120364,I120571,I120588,I120605,I120622,I120639,I120656,I120673,I120361,I120704,I120721,I120358,I120752,I120769,I120376,I120800,I120373,I12083_rst1,I120848,I120352,I120355,I120893,I120910,I120927,I120944,I120382,I120975,I120367,I120370,I121053_rst,I121070,I121087,I121104,I121121,I121138,I121155,I121172,I121042,I121203,I121027,I121234,I121251,I121268,I121285,I121302,I121319,I121336,I121024,I121367,I121384,I121021,I121415,I121432,I121039,I121463,I121036,I121494,I121511,I121015,I121018,I121556,I121573,I121590,I121607,I121045,I121638,I121030,I121033,I121716_rst,I121733,I121750,I121767,I121784,I121801,I121818,I121835,I121705,I121866,I121690,I121897,I121914,I121931,I121948,I121965,I121982,I121999,I121687,I122030,I122047,I121684,I122078,I122095,I121702,I122126,I121699,I122157,I122174,I121678,I121681,I122219,I122236,I122253,I122270,I121708,I122301,I121693,I121696,I122379_rst,I122396,I122413,I122430,I122447,I122464,I122481,I122498,I122368,I122529,I122353,I122560,I122577,I122594,I122611,I122628,I122645,I122662,I122350,I122693,I122710,I122347,I122741,I122758,I122365,I122789,I122362,I122820,I122837,I122341,I122344,I122882,I122899,I122916,I122933,I122371,I122964,I122356,I122359,I123042_rst,I123059,I123076,I123093,I123110,I123127,I123144,I123161,I123031,I123192,I123016,I123223,I123240,I123257,I123274,I123291,I123308,I123325,I123013,I123356,I123373,I123010,I123404,I123421,I123028,I123452,I123025,I123483,I123500,I123004,I123007,I123545,I123562,I123579,I123596,I123034,I123627,I123019,I123022,I123705_rst,I123722,I123739,I123756,I123773,I123790,I123807,I123824,I123694,I123855,I123679,I123886,I123903,I123920,I123937,I123954,I123971,I123988,I123676,I124019,I124036,I123673,I124067,I124084,I123691,I124115,I123688,I124146,I124163,I123667,I123670,I124208,I124225,I124242,I124259,I123697,I124290,I123682,I123685,I124368_rst,I124385,I124402,I124419,I124436,I124453,I124470,I124487,I124357,I124518,I124342,I124549,I124566,I124583,I124600,I124617,I124634,I124651,I124339,I124682,I124699,I124336,I124730,I124747,I124354,I124778,I124351,I124809,I124826,I124330,I124333,I124871,I124888,I124905,I124922,I124360,I124953,I124345,I124348,I125031_rst,I125048,I125065,I125082,I125099,I125116,I125133,I125150,I125020,I125181,I125005,I125212,I125229,I125246,I125263,I125280,I125297,I125314,I125002,I125345,I125362,I124999,I125393,I125410,I125017,I125441,I125014,I125472,I125489,I124993,I124996,I125534,I125551,I125568,I125585,I125023,I125616,I125008,I125011,I125694_rst,I125711,I125728,I125745,I125762,I125779,I125796,I125813,I125683,I125844,I125668,I125875,I125892,I125909,I125926,I125943,I125960,I125977,I125665,I126008,I126025,I125662,I126056,I126073,I125680,I126104,I125677,I126135,I126152,I125656,I125659,I126197,I126214,I126231,I126248,I125686,I126279,I125671,I125674,I126357_rst,I126374,I126391,I126408,I126425,I126442,I126459,I126476,I126346,I126507,I126331,I126538,I126555,I126572,I126589,I126606,I126623,I126640,I126328,I126671,I126688,I126325,I126719,I126736,I126343,I126767,I126340,I126798,I126815,I126319,I126322,I126860,I126877,I126894,I126911,I126349,I126942,I126334,I126337,I127020_rst,I127037,I127054,I127071,I127088,I127105,I127122,I127139,I127009,I127170,I126994,I127201,I127218,I127235,I127252,I127269,I127286,I127303,I126991,I127334,I127351,I126988,I127382,I127399,I127006,I127430,I127003,I127461,I127478,I126982,I126985,I127523,I127540,I127557,I127574,I127012,I127605,I126997,I127000,I127683_rst,I127700,I127717,I127734,I127751,I127768,I127785,I127654,I127816,I127833,I127850,I127867,I127884,I127901,I127918,I127651,I127949,I127645,I127980,I127997,I128014,I127675,I127648,I128059,I127672,I128090,I127669,I127666,I128135,I128152,I128169,I128186,I128203,I127660,I128234,I128251,I127663,I127657,I128329_rst,I128346,I128363,I128380,I128397,I128414,I128431,I128300,I128462,I128479,I128496,I128513,I128530,I128547,I128564,I128297,I128595,I128291,I128626,I128643,I128660,I128321,I128294,I128705,I128318,I128736,I128315,I128312,I128781,I128798,I128815,I128832,I128849,I128306,I128880,I128897,I128309,I128303,I128975_rst,I128992,I129009,I129026,I129043,I129060,I129077,I128946,I129108,I129125,I129142,I129159,I129176,I129193,I129210,I128943,I129241,I128937,I129272,I129289,I129306,I128967,I128940,I129351,I128964,I129382,I128961,I128958,I129427,I129444,I129461,I129478,I129495,I128952,I129526,I129543,I128955,I128949,I129621_rst,I129638,I129655,I129672,I129689,I129706,I129723,I129592,I129754,I129771,I129788,I129805,I129822,I129839,I129856,I129589,I129887,I129583,I129918,I129935,I129952,I129613,I129586,I129997,I129610,I130028,I129607,I129604,I130073,I130090,I130107,I130124,I130141,I129598,I130172,I130189,I129601,I129595,I130267_rst,I130284,I130301,I130318,I130335,I130352,I130369,I130238,I130400,I130417,I130434,I130451,I130468,I130485,I130502,I130235,I130533,I130229,I130564,I130581,I130598,I130259,I130232,I130643,I130256,I130674,I130253,I130250,I130719,I130736,I130753,I130770,I130787,I130244,I130818,I130835,I130247,I130241,I130913_rst,I130930,I130947,I130964,I130981,I130998,I131015,I130884,I131046,I131063,I131080,I131097,I131114,I131131,I131148,I130881,I131179,I130875,I131210,I131227,I131244,I130905,I130878,I131289,I130902,I131320,I130899,I130896,I131365,I131382,I131399,I131416,I131433,I130890,I131464,I131481,I130893,I130887,I131559_rst,I131576,I131593,I131610,I131627,I131644,I131661,I131530,I131692,I131709,I131726,I131743,I131760,I131777,I131794,I131527,I131825,I131521,I131856,I131873,I131890,I131551,I131524,I131935,I131548,I131966,I131545,I131542,I132011,I132028,I132045,I132062,I132079,I131536,I132110,I132127,I131539,I131533,I132205_rst,I132222,I132239,I132256,I132273,I132290,I132307,I132176,I132338,I132355,I132372,I132389,I132406,I132423,I132440,I132173,I132471,I132167,I132502,I132519,I132536,I132197,I132170,I132581,I132194,I132612,I132191,I132188,I132657,I132674,I132691,I132708,I132725,I132182,I132756,I132773,I132185,I132179,I132851_rst,I132868,I132885,I132902,I132919,I132936,I132953,I132822,I132984,I133001,I133018,I133035,I133052,I133069,I133086,I132819,I133117,I132813,I133148,I133165,I133182,I132843,I132816,I133227,I132840,I133258,I132837,I132834,I133303,I133320,I133337,I133354,I133371,I132828,I133402,I13341_rst9,I132831,I132825,I133497_rst,I133514,I133531,I133548,I133565,I133582,I133599,I133468,I133630,I133647,I133664,I133681,I133698,I133715,I133732,I133465,I133763,I133459,I133794,I133811,I133828,I133489,I133462,I133873,I133486,I133904,I133483,I133480,I133949,I133966,I133983,I134000,I134017,I133474,I134048,I134065,I133477,I133471,I134143_rst,I134160,I134177,I134194,I134211,I134228,I134245,I134114,I134276,I134293,I134310,I134327,I134344,I134361,I134378,I134111,I134409,I134105,I134440,I134457,I134474,I134135,I134108,I134519,I134132,I134550,I134129,I134126,I134595,I134612,I134629,I134646,I134663,I134120,I134694,I134711,I134123,I134117,I134789_rst,I134806,I134823,I134840,I134857,I134874,I134891,I134760,I134922,I134939,I134956,I134973,I134990,I135007,I135024,I134757,I135055,I134751,I135086,I135103,I135120,I134781,I134754,I135165,I134778,I135196,I134775,I134772,I135241,I135258,I135275,I135292,I135309,I134766,I135340,I135357,I134769,I134763,I135435_rst,I135452,I135469,I135486,I135503,I135520,I135537,I135406,I135568,I135585,I135602,I135619,I135636,I135653,I135670,I135403,I135701,I135397,I135732,I135749,I135766,I135427,I135400,I135811,I135424,I135842,I135421,I135418,I135887,I135904,I135921,I135938,I135955,I135412,I135986,I136003,I135415,I135409,I136081_rst,I136098,I136115,I136132,I136149,I136166,I136183,I136052,I136214,I136231,I136248,I136265,I136282,I136299,I136316,I136049,I136347,I136043,I136378,I136395,I136412,I136073,I136046,I136457,I136070,I136488,I136067,I136064,I136533,I136550,I136567,I136584,I136601,I136058,I136632,I136649,I136061,I136055,I136727_rst,I136744,I136761,I136778,I136795,I136689,I136826,I136843,I136860,I136877,I136894,I136911,I136698,I136942,I136692,I136973,I136990,I137007,I137024,I136719,I136716,I137069,I137086,I137103,I136713,I137134,I136710,I136701,I137179,I137196,I137213,I136704,I136707,I137258,I137275,I136695,I137339_rst,I137356,I137373,I137390,I137407,I137301,I137438,I137455,I137472,I137489,I137506,I137523,I137310,I137554,I137304,I137585,I137602,I137619,I137636,I137331,I137328,I137681,I137698,I137715,I137325,I137746,I137322,I137313,I137791,I137808,I137825,I137316,I137319,I137870,I137887,I137307,I137951_rst,I137968,I137985,I138002,I138019,I137919,I138050,I138067,I138084,I137922,I138115,I137916,I138146,I138163,I138180,I138197,I138214,I137925,I138245,I138262,I138279,I138296,I137931,I137934,I137913,I138355,I138372,I138389,I137943,I137940,I138434,I138451,I137928,I137937,I138529_rst,I138546,I138563,I138580,I138597,I138497,I138628,I138645,I138662,I138500,I138693,I138494,I138724,I138741,I138758,I138775,I138792,I138503,I138823,I138840,I138857,I138874,I138509,I138512,I138491,I138933,I138950,I138967,I138521,I138518,I139012,I139029,I138506,I138515,I139107_rst,I139124,I139141,I139158,I139175,I139075,I139206,I139223,I139240,I139078,I139271,I139072,I139302,I139319,I139336,I139353,I139370,I139081,I139401,I139418,I139435,I139452,I139087,I139090,I139069,I139511,I139528,I139545,I139099,I139096,I139590,I139607,I139084,I139093,I139685_rst,I139702,I139719,I139736,I139753,I139653,I139784,I139801,I139818,I139656,I139849,I139650,I139880,I139897,I139914,I139931,I139948,I139659,I139979,I139996,I140013,I140030,I139665,I139668,I139647,I140089,I140106,I140123,I139677,I139674,I140168,I140185,I139662,I139671,I140263_rst,I140280,I140297,I140314,I140331,I140231,I140362,I140379,I140396,I140413,I140430,I140447,I140464,I140481,I140237,I140228,I140526,I140543,I140252,I140574,I140591,I140240,I140622,I140639,I140246,I140670,I140234,I140701,I140225,I140732,I140749,I140255,I140780,I140249,I140811,I140243,I140875_rst,I140892,I140909,I140926,I140943,I140843,I140974,I140991,I141008,I141025,I141042,I141059,I141076,I141093,I140849,I140840,I141138,I141155,I140864,I141186,I141203,I140852,I141234,I141251,I140858,I141282,I140846,I141313,I140837,I141344,I141361,I140867,I141392,I140861,I141423,I140855,I141487_rst,I141504,I141521,I141538,I141555,I141455,I141586,I141603,I141620,I141637,I141654,I141671,I141688,I141705,I141461,I141452,I141750,I141767,I141476,I141798,I141815,I141464,I141846,I141863,I141470,I141894,I141458,I141925,I141449,I141956,I141973,I141479,I142004,I141473,I142035,I141467,I142099_rst,I142116,I142133,I142150,I142088,I142181,I142198,I142215,I142232,I142249,I142266,I142283,I142073,I142314,I142070,I142345,I142082,I142376,I142393,I142410,I142076,I142091,I142455,I142472,I142061,I142503,I142079,I142534,I142551,I142085,I142582,I142599,I142064,I142067,I142677_rst,I142694,I142711,I142728,I142666,I142759,I142776,I142793,I142810,I142827,I142844,I142861,I142651,I142892,I142648,I142923,I142660,I142954,I142971,I142988,I142654,I142669,I143033,I143050,I142639,I143081,I142657,I143112,I143129,I142663,I143160,I143177,I142642,I142645,I143255_rst,I143272,I143289,I143306,I143323,I143340,I143238,I143371,I143388,I143405,I143241,I143223,I143450,I143467,I143484,I143244,I143235,I143529,I143546,I143563,I143226,I143594,I143611,I143217,I143642,I143659,I143676,I143247,I143707,I143724,I143741,I143758,I143232,I143229,I143220,I143850_rst,I143867,I143884,I143901,I143918,I143935,I143833,I143966,I143983,I144000,I143836,I143818,I144045,I144062,I144079,I143839,I143830,I144124,I144141,I144158,I143821,I144189,I144206,I143812,I144237,I144254,I144271,I143842,I144302,I144319,I144336,I144353,I143827,I143824,I143815,I144445_rst,I144462,I144479,I144496,I144513,I144530,I144428,I144561,I144578,I144595,I144431,I144413,I144640,I144657,I144674,I144434,I144425,I144719,I144736,I144753,I144416,I144784,I144801,I144407,I144832,I144849,I144866,I144437,I144897,I144914,I144931,I144948,I144422,I144419,I144410,I145040_rst,I145057,I145074,I145091,I145108,I145125,I145023,I145156,I145173,I145190,I145026,I145008,I145235,I145252,I145269,I145029,I145020,I145314,I145331,I145348,I145011,I145379,I145396,I145002,I145427,I145444,I145461,I145032,I145492,I145509,I145526,I145543,I145017,I145014,I145005,I145635_rst,I145652,I145669,I145686,I145703,I145720,I145618,I145751,I145768,I145785,I145621,I145603,I145830,I145847,I145864,I145624,I145615,I145909,I145926,I145943,I145606,I145974,I145991,I145597,I146022,I146039,I146056,I145627,I146087,I146104,I146121,I146138,I145612,I145609,I145600,I146230_rst,I146247,I146264,I146281,I146298,I146315,I146213,I146346,I146363,I146380,I146216,I146198,I146425,I146442,I146459,I146219,I146210,I146504,I146521,I146538,I146201,I146569,I146586,I146192,I146617,I146634,I146651,I146222,I146682,I146699,I146716,I146733,I146207,I146204,I146195,I146825_rst,I146842,I146859,I146876,I146893,I146910,I146808,I146941,I146958,I146975,I146811,I146793,I147020,I147037,I147054,I146814,I146805,I147099,I147116,I147133,I146796,I147164,I147181,I146787,I147212,I147229,I147246,I146817,I147277,I147294,I147311,I147328,I146802,I146799,I146790,I147420_rst,I147437,I147454,I147471,I147488,I147505,I147403,I147536,I147553,I147570,I147406,I147388,I147615,I147632,I147649,I147409,I147400,I147694,I147711,I147728,I147391,I147759,I147776,I147382,I147807,I147824,I147841,I147412,I147872,I147889,I147906,I147923,I147397,I147394,I147385,I148015_rst,I148032,I148049,I148066,I148083,I148100,I147998,I148131,I148148,I148165,I148001,I147983,I148210,I148227,I148244,I148004,I147995,I148289,I148306,I148323,I147986,I148354,I148371,I147977,I148402,I148419,I148436,I148007,I148467,I148484,I148501,I148518,I147992,I147989,I147980,I148610_rst,I148627,I148644,I148661,I148678,I148695,I148593,I148726,I148743,I148760,I148596,I148578,I148805,I148822,I148839,I148599,I148590,I148884,I148901,I148918,I148581,I148949,I148966,I148572,I148997,I149014,I149031,I148602,I149062,I149079,I149096,I149113,I148587,I148584,I148575,I149205_rst,I149222,I149239,I149256,I149273,I149290,I149307,I149176,I149338,I149355,I149372,I149389,I149406,I149423,I149440,I149173,I149167,I149485,I149502,I149519,I149194,I149550,I149567,I149185,I149179,I149612,I149182,I149643,I149660,I149197,I149691,I149191,I149188,I149736,I149170,I149800_rst,I149817,I149834,I149851,I149868,I149885,I149902,I149771,I149933,I149950,I149967,I149984,I150001,I150018,I150035,I149768,I149762,I150080,I150097,I150114,I149789,I150145,I150162,I149780,I149774,I150207,I149777,I150238,I150255,I149792,I150286,I149786,I149783,I150331,I149765,I150395_rst,I150412,I150429,I150446,I150463,I150480,I150497,I150366,I150528,I150545,I150562,I150579,I150596,I150613,I150630,I150363,I150357,I150675,I150692,I150709,I150384,I150740,I150757,I150375,I150369,I150802,I150372,I150833,I150850,I150387,I150881,I150381,I150378,I150926,I150360,I150990_rst,I151007,I151024,I151041,I151058,I151075,I151092,I150961,I151123,I151140,I151157,I151174,I151191,I151208,I151225,I150958,I150952,I151270,I151287,I151304,I150979,I151335,I151352,I150970,I150964,I151397,I150967,I151428,I151445,I150982,I151476,I150976,I150973,I151521,I150955,I151585_rst,I151602,I151619,I151636,I151653,I151670,I151687,I151556,I151718,I151735,I151752,I151769,I151786,I151803,I151820,I151553,I151547,I151865,I151882,I151899,I151574,I151930,I151947,I151565,I151559,I151992,I151562,I152023,I152040,I151577,I152071,I151571,I151568,I152116,I151550,I152180_rst,I152197,I152214,I152231,I152248,I152265,I152282,I152151,I152313,I152330,I152347,I152364,I152381,I152398,I152415,I152148,I152142,I152460,I152477,I152494,I152169,I152525,I152542,I152160,I152154,I152587,I152157,I152618,I152635,I152172,I152666,I152166,I152163,I152711,I152145,I152775_rst,I152792,I152809,I152826,I152843,I152860,I152877,I152746,I152908,I152925,I152942,I152959,I152976,I152993,I153010,I152743,I152737,I153055,I153072,I153089,I152764,I153120,I153137,I152755,I152749,I153182,I152752,I153213,I153230,I152767,I153261,I152761,I152758,I15330_rst6,I152740,I153370_rst,I153387,I153404,I153421,I153438,I153455,I153472,I153489,I153506,I153523,I153540,I153557,I153574,I153591,I153359,I153622,I153639,I153656,I153332,I153687,I153353,I153718,I153735,I153338,I153766,I153335,I153341,I153811,I153828,I153845,I153347,I153362,I153350,I153904,I153921,I153356,I153344,I153999_rst,I154016,I154033,I154050,I154067,I154084,I154101,I154118,I154135,I154152,I154169,I154186,I154203,I154220,I153988,I154251,I154268,I154285,I153961,I154316,I153982,I154347,I154364,I153967,I154395,I153964,I153970,I154440,I154457,I154474,I153976,I153991,I153979,I154533,I154550,I153985,I153973,I154628_rst,I154645,I154662,I154679,I154696,I154713,I154730,I154747,I154764,I154781,I154798,I154815,I154832,I154849,I154617,I154880,I154897,I154914,I154590,I154945,I154611,I154976,I154993,I154596,I155024,I154593,I154599,I155069,I155086,I155103,I154605,I154620,I154608,I155162,I155179,I154614,I154602,I155257_rst,I155274,I155291,I155308,I155325,I155342,I155359,I155376,I155393,I155410,I155427,I155444,I155461,I155478,I155246,I155509,I155526,I155543,I155219,I155574,I155240,I155605,I155622,I155225,I155653,I155222,I155228,I155698,I155715,I155732,I155234,I155249,I155237,I155791,I155808,I155243,I155231,I155886_rst,I155903,I155920,I155937,I155954,I155971,I155988,I156005,I156022,I156039,I156056,I156073,I156090,I156107,I155875,I156138,I156155,I156172,I155848,I156203,I155869,I156234,I156251,I155854,I156282,I155851,I155857,I156327,I156344,I156361,I155863,I155878,I155866,I156420,I156437,I155872,I155860,I156515_rst,I156532,I156549,I156566,I156583,I156600,I156617,I156634,I156651,I156668,I156685,I156702,I156719,I156736,I156504,I156767,I156784,I156801,I156477,I156832,I156498,I156863,I156880,I156483,I156911,I156480,I156486,I156956,I156973,I156990,I156492,I156507,I156495,I157049,I157066,I156501,I156489,I157144_rst,I157161,I157178,I157195,I157212,I157229,I157246,I157263,I157280,I157297,I157314,I157331,I157348,I157365,I157133,I157396,I157413,I157430,I157106,I157461,I157127,I157492,I157509,I157112,I157540,I157109,I157115,I157585,I157602,I157619,I157121,I157136,I157124,I157678,I157695,I157130,I157118,I157773_rst,I157790,I157807,I157824,I157841,I157858,I157875,I157892,I157909,I157926,I157943,I157960,I157977,I157994,I157762,I158025,I158042,I158059,I157735,I158090,I157756,I158121,I158138,I157741,I158169,I157738,I157744,I158214,I158231,I158248,I157750,I157765,I157753,I158307,I158324,I157759,I157747,I158402_rst,I158419,I158436,I158453,I158470,I158487,I158504,I158521,I158538,I158555,I158572,I158589,I158606,I158623,I158391,I158654,I158671,I158688,I158364,I158719,I158385,I158750,I158767,I158370,I158798,I158367,I158373,I158843,I158860,I158877,I158379,I158394,I158382,I158936,I158953,I158388,I158376,I159031_rst,I159048,I159065,I159082,I159020,I159113,I159008,I159144,I159161,I159178,I159195,I159212,I159011,I159243,I158996,I159274,I159291,I159308,I159325,I159342,I159359,I159002,I159390,I159407,I159424,I159014,I159023,I158993,I159483,I159017,I159005,I159528,I159545,I158999,I159609_rst,I159626,I159643,I159660,I159598,I159691,I159586,I159722,I159739,I159756,I159773,I159790,I159589,I159821,I159574,I159852,I159869,I159886,I159903,I159920,I15993_rst7,I159580,I159968,I159985,I160002,I159592,I159601,I159571,I160061,I159595,I159583,I160106,I160123,I159577,I160187_rst,I160204,I160221,I160238,I160176,I160269,I160164,I160300,I160317,I160334,I160351,I160368,I160167,I160399,I160152,I160430,I160447,I160464,I160481,I160498,I160515,I160158,I160546,I160563,I160580,I160170,I160179,I160149,I160639,I160173,I160161,I160684,I160701,I160155,I160765_rst,I160782,I160799,I160816,I160754,I160847,I160742,I160878,I160895,I160912,I160929,I160946,I160745,I160977,I160730,I161008,I161025,I161042,I161059,I161076,I161093,I160736,I161124,I161141,I161158,I160748,I160757,I160727,I161217,I160751,I160739,I161262,I161279,I160733,I161343_rst,I161360,I161377,I161394,I161411,I161428,I161326,I161314,I161473,I161490,I161507,I161524,I161541,I161323,I161572,I161589,I161606,I161623,I161332,I161311,I161668,I161685,I161329,I161716,I161320,I161335,I161761,I161778,I161795,I161812,I161308,I161317,I161305,I161904_rst,I161921,I161938,I161955,I161972,I161989,I161887,I161875,I162034,I162051,I162068,I162085,I162102,I161884,I162133,I162150,I162167,I162184,I161893,I161872,I162229,I162246,I161890,I162277,I161881,I161896,I162322,I162339,I162356,I162373,I161869,I161878,I161866,I162465_rst,I162482,I162499,I162516,I162533,I162550,I162448,I162436,I162595,I162612,I162629,I162646,I162663,I162445,I162694,I162711,I162728,I162745,I162454,I162433,I162790,I162807,I162451,I162838,I162442,I162457,I162883,I162900,I162917,I162934,I162430,I162439,I162427,I163026_rst,I163043,I163060,I163077,I163094,I163111,I163009,I162997,I163156,I163173,I163190,I163207,I163224,I163006,I163255,I163272,I163289,I163306,I163015,I162994,I163351,I163368,I163012,I163399,I163003,I163018,I163444,I163461,I163478,I163495,I162991,I163000,I162988,I163587_rst,I163604,I163621,I163638,I163655,I163672,I163570,I163558,I163717,I163734,I163751,I163768,I163785,I163567,I163816,I163833,I163850,I163867,I163576,I163555,I163912,I163929,I163573,I163960,I163564,I163579,I164005,I164022,I164039,I164056,I163552,I163561,I163549,I164148_rst,I164165,I164182,I164199,I164216,I164233,I164131,I164119,I164278,I164295,I164312,I164329,I164346,I164128,I164377,I164394,I164411,I164428,I164137,I164116,I164473,I164490,I164134,I164521,I164125,I164140,I164566,I164583,I164600,I164617,I164113,I164122,I164110,I164709_rst,I164726,I164743,I164760,I164683,I164791,I164808,I164698,I164680,I164853,I164870,I164887,I164904,I164921,I164938,I164955,I164972,I164989,I164695,I165020,I165037,I165054,I164677,I165085,I164674,I165116,I165133,I165150,I165167,I164689,I165198,I164686,I165229,I165246,I165263,I164692,I164701,I164671,I165355_rst,I165372,I165389,I165406,I165329,I165437,I165454,I165344,I165326,I165499,I165516,I165533,I165550,I165567,I165584,I165601,I165618,I165635,I165341,I165666,I165683,I165700,I165323,I165731,I165320,I165762,I165779,I165796,I165813,I165335,I165844,I165332,I165875,I165892,I165909,I165338,I165347,I165317,I166001_rst,I166018,I166035,I166052,I165975,I166083,I166100,I165990,I165972,I166145,I166162,I166179,I166196,I166213,I166230,I166247,I166264,I166281,I165987,I166312,I166329,I166346,I165969,I166377,I165966,I166408,I166425,I166442,I166459,I165981,I166490,I165978,I166521,I166538,I166555,I165984,I165993,I165963,I166647_rst,I166664,I166681,I166698,I166621,I166729,I166746,I166636,I166618,I166791,I166808,I166825,I166842,I166859,I166876,I166893,I166910,I166927,I166633,I166958,I166975,I166992,I166615,I167023,I166612,I167054,I167071,I167088,I167105,I166627,I167136,I166624,I167167,I167184,I167201,I166630,I166639,I166609,I167293_rst,I167310,I167327,I167344,I167267,I167375,I167392,I167282,I167264,I167437,I167454,I167471,I167488,I167505,I167522,I167539,I167556,I167573,I167279,I167604,I167621,I167638,I167261,I167669,I167258,I167700,I167717,I167734,I167751,I167273,I167782,I167270,I167813,I167830,I167847,I167276,I167285,I167255,I167939_rst,I167956,I167973,I167990,I167913,I168021,I168038,I167928,I167910,I168083,I168100,I168117,I168134,I168151,I168168,I168185,I168202,I168219,I167925,I168250,I168267,I168284,I167907,I168315,I167904,I168346,I168363,I168380,I168397,I167919,I168428,I167916,I168459,I168476,I168493,I167922,I167931,I167901,I168585_rst,I168602,I168619,I168636,I168559,I168667,I168684,I168574,I168556,I168729,I168746,I168763,I168780,I168797,I168814,I168831,I168848,I168865,I168571,I168896,I168913,I168930,I168553,I168961,I168550,I168992,I169009,I169026,I169043,I168565,I169074,I168562,I169105,I169122,I169139,I168568,I168577,I168547,I169231_rst,I169248,I169265,I169282,I169205,I169313,I169330,I169220,I169202,I169375,I169392,I169409,I169426,I169443,I169460,I169477,I169494,I169511,I169217,I169542,I169559,I169576,I169199,I169607,I169196,I169638,I169655,I169672,I169689,I169211,I169720,I169208,I169751,I169768,I169785,I169214,I169223,I169193,I169877_rst,I169894,I169911,I169928,I169851,I169959,I169976,I169866,I169848,I170021,I170038,I170055,I170072,I170089,I170106,I170123,I170140,I170157,I169863,I170188,I170205,I170222,I169845,I170253,I169842,I170284,I170301,I170318,I170335,I169857,I170366,I169854,I170397,I170414,I170431,I169860,I169869,I169839,I170523_rst,I170540,I170557,I170574,I170497,I170605,I170622,I170512,I170494,I170667,I170684,I170701,I170718,I170735,I170752,I170769,I170786,I170803,I170509,I170834,I170851,I170868,I170491,I170899,I170488,I170930,I170947,I170964,I170981,I170503,I171012,I170500,I171043,I171060,I171077,I170506,I170515,I170485,I171169_rst,I171186,I171203,I171220,I171143,I171251,I171268,I171158,I171140,I171313,I171330,I171347,I171364,I171381,I171398,I171415,I171432,I171449,I171155,I171480,I171497,I171514,I171137,I171545,I171134,I171576,I171593,I171610,I171627,I171149,I171658,I171146,I171689,I171706,I171723,I171152,I171161,I171131,I171815_rst,I171832,I171849,I171866,I171789,I171897,I171914,I171804,I171786,I171959,I171976,I171993,I172010,I172027,I172044,I172061,I172078,I172095,I171801,I172126,I172143,I172160,I171783,I172191,I171780,I172222,I172239,I172256,I172273,I171795,I172304,I171792,I172335,I172352,I172369,I171798,I171807,I171777,I172461_rst,I172478,I172495,I172512,I172435,I172543,I172560,I172450,I172432,I172605,I172622,I172639,I172656,I172673,I172690,I172707,I172724,I172741,I172447,I172772,I172789,I172806,I172429,I172837,I172426,I172868,I172885,I172902,I172919,I172441,I172950,I172438,I172981,I172998,I173015,I172444,I172453,I172423,I173107_rst,I173124,I173141,I173158,I173081,I173189,I173206,I173096,I173078,I173251,I173268,I173285,I173302,I173319,I173336,I173353,I173370,I173387,I173093,I173418,I173435,I173452,I173075,I173483,I173072,I173514,I173531,I173548,I173565,I173087,I173596,I173084,I173627,I173644,I173661,I173090,I173099,I173069,I173753_rst,I173770,I173787,I173804,I173724,I173835,I173852,I173869,I173886,I173903,I173920,I173937,I173954,I173971,I173988,I173739,I173736,I174033,I173721,I174064,I173718,I174095,I174112,I174129,I174146,I174163,I174180,I173745,I174211,I173733,I173727,I174256,I174273,I173742,I174304,I174321,I174338,I173730,I173715,I174416_rst,I174433,I174450,I174467,I174387,I174498,I174515,I174532,I174549,I174566,I174583,I174600,I174617,I174634,I174651,I174402,I174399,I174696,I174384,I174727,I174381,I174758,I174775,I174792,I174809,I174826,I174843,I174408,I174874,I174396,I174390,I174919,I174936,I174405,I174967,I174984,I175001,I174393,I174378,I175079_rst,I175096,I175113,I175130,I175050,I175161,I175178,I175195,I175212,I175229,I175246,I175263,I175280,I175297,I175314,I175065,I175062,I175359,I175047,I175390,I175044,I175421,I175438,I175455,I175472,I175489,I175506,I175071,I175537,I175059,I175053,I175582,I175599,I175068,I175630,I175647,I175664,I175056,I175041,I175742_rst,I175759,I175776,I175793,I175713,I175824,I175841,I175858,I175875,I175892,I175909,I175926,I175943,I175960,I175977,I175728,I175725,I176022,I175710,I176053,I175707,I176084,I176101,I176118,I176135,I176152,I176169,I175734,I176200,I175722,I175716,I176245,I176262,I175731,I176293,I176310,I176327,I175719,I175704,I176405_rst,I176422,I176439,I176456,I176376,I176487,I176504,I176521,I176538,I176555,I176572,I176589,I176606,I176623,I176640,I176391,I176388,I176685,I176373,I176716,I176370,I176747,I176764,I176781,I176798,I176815,I176832,I176397,I176863,I176385,I176379,I176908,I176925,I176394,I176956,I176973,I176990,I176382,I176367,I177068_rst,I177085,I177102,I177119,I177039,I177150,I177167,I177184,I177201,I177218,I177235,I177252,I177269,I177286,I177303,I177054,I177051,I177348,I177036,I177379,I177033,I177410,I177427,I177444,I177461,I177478,I177495,I177060,I177526,I177048,I177042,I177571,I177588,I177057,I177619,I177636,I177653,I177045,I177030,I177731_rst,I177748,I177765,I177782,I177702,I177813,I177830,I177847,I177864,I177881,I177898,I177915,I177932,I177949,I177966,I177717,I177714,I178011,I177699,I178042,I177696,I178073,I178090,I178107,I178124,I178141,I178158,I177723,I178189,I177711,I177705,I178234,I178251,I177720,I178282,I178299,I178316,I177708,I177693,I178394_rst,I178411,I178428,I178445,I178365,I178476,I178493,I178510,I178527,I178544,I178561,I178578,I178595,I178612,I178629,I178380,I178377,I178674,I178362,I178705,I178359,I178736,I178753,I178770,I178787,I178804,I178821,I178386,I178852,I178374,I178368,I178897,I178914,I178383,I178945,I178962,I178979,I178371,I178356,I179057_rst,I179074,I179091,I179108,I179028,I179139,I179156,I179173,I179190,I179207,I179224,I179241,I179258,I179275,I179292,I179043,I179040,I179337,I179025,I179368,I179022,I179399,I179416,I179433,I179450,I179467,I179484,I179049,I179515,I179037,I179031,I179560,I179577,I179046,I179608,I179625,I179642,I179034,I179019,I179720_rst,I179737,I179754,I179694,I179785,I179802,I179819,I179836,I179853,I179870,I179887,I179904,I179921,I179688,I179952,I179969,I179685,I180000,I180017,I180034,I179697,I179682,I180079,I180096,I180113,I180130,I180147,I179703,I180178,I179712,I180209,I179706,I179709,I179700,I179691,I180315_rst,I180332,I180349,I180289,I180380,I180397,I180414,I180431,I180448,I180465,I180482,I180499,I180516,I180283,I180547,I180564,I180280,I180595,I180612,I180629,I180292,I180277,I180674,I180691,I180708,I180725,I180742,I180298,I180773,I180307,I180804,I180301,I180304,I180295,I180286,I180910_rst,I180927,I180944,I180884,I180975,I180992,I181009,I181026,I181043,I181060,I181077,I181094,I181111,I180878,I181142,I181159,I180875,I181190,I181207,I181224,I180887,I180872,I181269,I181286,I181303,I181320,I181337,I180893,I181368,I180902,I181399,I180896,I180899,I180890,I180881,I181505_rst,I181522,I181539,I181479,I181570,I181587,I181604,I181621,I181638,I181655,I181672,I181689,I181706,I181473,I181737,I181754,I181470,I181785,I181802,I181819,I181482,I181467,I181864,I181881,I181898,I181915,I181932,I181488,I181963,I181497,I181994,I181491,I181494,I181485,I181476,I182100_rst,I182117,I182083,I182062,I182162,I182179,I182196,I182213,I182230,I182247,I182264,I182281,I182298,I182089,I182329,I182346,I182363,I182380,I182092,I182411,I182428,I182445,I182462,I182479,I182077,I182510,I182527,I182080,I182074,I182068,I182586,I182086,I182617,I182071,I182065,I182695_rst,I182712,I182678,I182657,I182757,I182774,I182791,I182808,I182825,I182842,I182859,I182876,I182893,I182684,I182924,I182941,I182958,I182975,I182687,I183006,I183023,I183040,I183057,I183074,I182672,I183105,I183122,I182675,I182669,I182663,I183181,I182681,I183212,I182666,I182660,I183290_rst,I183307,I183324,I183341,I183358,I183375,I183392,I183409,I183279,I183440,I183264,I183471,I183488,I183505,I183522,I183539,I183556,I183573,I183261,I183604,I183621,I183258,I183652,I183669,I183276,I183700,I183273,I183731,I183748,I183252,I183255,I183793,I183810,I183827,I183844,I183282,I183875,I183267,I183270,I183953_rst,I183970,I183987,I184004,I184021,I184038,I184055,I184072,I183942,I184103,I183927,I184134,I184151,I184168,I184185,I184202,I184219,I184236,I183924,I184267,I184284,I183921,I184315,I184332,I183939,I184363,I183936,I184394,I184411,I183915,I183918,I184456,I184473,I184490,I184507,I183945,I184538,I183930,I183933,I184616_rst,I184633,I184650,I184667,I184684,I184701,I184718,I184735,I184605,I184766,I184590,I184797,I184814,I184831,I184848,I184865,I184882,I184899,I184587,I184930,I184947,I184584,I184978,I184995,I184602,I185026,I184599,I185057,I185074,I184578,I184581,I185119,I185136,I185153,I185170,I184608,I185201,I184593,I184596,I185279_rst,I185296,I185313,I185330,I185347,I185364,I185381,I185398,I185268,I185429,I185253,I185460,I185477,I185494,I185511,I185528,I185545,I185562,I185250,I185593,I185610,I185247,I185641,I185658,I185265,I185689,I185262,I185720,I185737,I185241,I185244,I185782,I185799,I185816,I185833,I185271,I185864,I185256,I185259,I185942_rst,I185959,I185976,I185993,I186010,I186027,I186044,I186061,I185931,I186092,I185916,I186123,I186140,I186157,I186174,I186191,I186208,I186225,I185913,I186256,I186273,I185910,I186304,I186321,I185928,I186352,I185925,I186383,I186400,I185904,I185907,I186445,I186462,I186479,I186496,I185934,I186527,I185919,I185922,I186605_rst,I186622,I186639,I186656,I186673,I186690,I186707,I186724,I186594,I186755,I186579,I186786,I186803,I186820,I186837,I186854,I186871,I186888,I186576,I186919,I186936,I186573,I186967,I186984,I186591,I187015,I186588,I187046,I187063,I186567,I186570,I187108,I187125,I187142,I187159,I186597,I187190,I186582,I186585,I187268_rst,I187285,I187302,I187319,I187336,I187353,I187370,I187387,I187257,I187418,I187242,I187449,I187466,I187483,I187500,I187517,I187534,I187551,I187239,I187582,I187599,I187236,I187630,I187647,I187254,I187678,I187251,I187709,I187726,I187230,I187233,I187771,I187788,I187805,I187822,I187260,I187853,I187245,I187248,I187931_rst,I187948,I187965,I187982,I187999,I188016,I188033,I188050,I187920,I188081,I187905,I188112,I188129,I188146,I188163,I188180,I188197,I188214,I187902,I188245,I188262,I187899,I188293,I188310,I187917,I188341,I187914,I188372,I188389,I187893,I187896,I188434,I188451,I188468,I188485,I187923,I188516,I187908,I187911,I188594_rst,I188611,I188628,I188645,I188662,I188679,I188696,I188713,I188583,I188744,I188568,I188775,I188792,I188809,I188826,I188843,I188860,I188877,I188565,I188908,I188925,I188562,I188956,I188973,I188580,I189004,I188577,I189035,I189052,I188556,I188559,I189097,I189114,I189131,I189148,I188586,I189179,I188571,I188574,I189257_rst,I189274,I189291,I189308,I189325,I189342,I189359,I189376,I189246,I189407,I189231,I189438,I189455,I189472,I189489,I189506,I189523,I189540,I189228,I189571,I189588,I189225,I189619,I189636,I189243,I189667,I189240,I189698,I189715,I189219,I189222,I189760,I189777,I189794,I189811,I189249,I189842,I189234,I189237,I189920_rst,I189937,I189954,I189971,I189988,I190005,I190022,I190039,I189909,I190070,I189894,I190101,I190118,I190135,I190152,I190169,I190186,I190203,I189891,I190234,I190251,I189888,I190282,I190299,I189906,I190330,I189903,I190361,I190378,I189882,I189885,I190423,I190440,I190457,I190474,I189912,I190505,I189897,I189900,I190583_rst,I190600,I190617,I190634,I190651,I190668,I190685,I190702,I190572,I190733,I190557,I190764,I190781,I190798,I190815,I190832,I190849,I190866,I190554,I190897,I190914,I190551,I190945,I190962,I190569,I190993,I190566,I191024,I191041,I190545,I190548,I191086,I191103,I191120,I191137,I190575,I191168,I190560,I190563,I191246_rst,I191263,I191280,I191297,I191314,I191331,I191348,I191365,I191235,I191396,I191220,I191427,I191444,I191461,I191478,I191495,I191512,I191529,I191217,I191560,I191577,I191214,I191608,I191625,I191232,I191656,I191229,I191687,I191704,I191208,I191211,I191749,I191766,I191783,I191800,I191238,I191831,I191223,I191226,I191909_rst,I191926,I191943,I191960,I191977,I191994,I192011,I192028,I191898,I192059,I191883,I192090,I192107,I192124,I192141,I192158,I192175,I192192,I191880,I192223,I192240,I191877,I192271,I192288,I191895,I192319,I191892,I192350,I192367,I191871,I191874,I192412,I192429,I192446,I192463,I191901,I192494,I191886,I191889,I192572_rst,I192589,I192606,I192623,I192640,I192657,I192674,I192691,I192561,I192722,I192546,I192753,I192770,I192787,I192804,I192821,I192838,I192855,I192543,I192886,I192903,I192540,I192934,I192951,I192558,I192982,I192555,I193013,I193030,I192534,I192537,I193075,I193092,I193109,I193126,I192564,I193157,I192549,I192552,I193235_rst,I193252,I193269,I193286,I193303,I193320,I193337,I193206,I193368,I193385,I193402,I193419,I193436,I193453,I193470,I193203,I193501,I193197,I193532,I193549,I193566,I193227,I193200,I193611,I193224,I193642,I193221,I193218,I193687,I193704,I193721,I193738,I193755,I193212,I193786,I193803,I193215,I193209,I193881_rst,I193898,I193915,I193932,I193949,I193966,I193983,I193852,I194014,I194031,I194048,I194065,I194082,I194099,I194116,I193849,I194147,I193843,I194178,I194195,I194212,I193873,I193846,I194257,I193870,I194288,I193867,I193864,I194333,I194350,I194367,I194384,I194401,I193858,I194432,I194449,I193861,I193855,I194527_rst,I194544,I194561,I194578,I194595,I194612,I194629,I194498,I194660,I194677,I194694,I194711,I194728,I194745,I194762,I194495,I194793,I194489,I194824,I194841,I194858,I194519,I194492,I194903,I194516,I194934,I194513,I194510,I194979,I194996,I195013,I195030,I195047,I194504,I195078,I195095,I194507,I194501,I195173_rst,I195190,I195207,I195224,I195241,I195258,I195275,I195144,I195306,I195323,I195340,I195357,I195374,I195391,I195408,I195141,I195439,I195135,I195470,I195487,I195504,I195165,I195138,I195549,I195162,I195580,I195159,I195156,I195625,I195642,I195659,I195676,I195693,I195150,I195724,I195741,I195153,I195147,I195819_rst,I195836,I195853,I195870,I195887,I195904,I195921,I195790,I195952,I195969,I195986,I196003,I196020,I196037,I196054,I195787,I196085,I195781,I196116,I196133,I196150,I195811,I195784,I196195,I195808,I196226,I195805,I195802,I196271,I196288,I196305,I196322,I196339,I195796,I196370,I196387,I195799,I195793,I196465_rst,I196482,I196499,I196516,I196533,I196550,I196567,I196436,I196598,I196615,I196632,I196649,I196666,I196683,I196700,I196433,I196731,I196427,I196762,I196779,I196796,I196457,I196430,I196841,I196454,I196872,I196451,I196448,I196917,I196934,I196951,I196968,I196985,I196442,I197016,I197033,I196445,I196439,I197111_rst,I197128,I197145,I197162,I197179,I197196,I197213,I197082,I197244,I197261,I197278,I197295,I197312,I197329,I197346,I197079,I197377,I197073,I197408,I197425,I197442,I197103,I197076,I197487,I197100,I197518,I197097,I197094,I197563,I197580,I197597,I197614,I197631,I197088,I197662,I197679,I197091,I197085,I197757_rst,I197774,I197791,I197808,I197825,I197719,I197856,I197873,I197890,I197907,I197924,I197941,I197728,I197972,I197722,I198003,I198020,I198037,I198054,I197749,I197746,I198099,I198116,I198133,I197743,I198164,I197740,I197731,I198209,I198226,I198243,I197734,I197737,I198288,I198305,I197725,I198369_rst,I198386,I198403,I198420,I198437,I198331,I198468,I198485,I198502,I198519,I198536,I198553,I198340,I198584,I198334,I198615,I198632,I198649,I198666,I198361,I198358,I198711,I198728,I198745,I198355,I198776,I198352,I198343,I198821,I198838,I198855,I198346,I198349,I198900,I198917,I198337,I198981_rst,I198998,I199015,I199032,I199049,I198943,I199080,I199097,I199114,I199131,I199148,I199165,I198952,I199196,I198946,I199227,I199244,I199261,I199278,I198973,I198970,I199323,I199340,I199357,I198967,I199388,I198964,I198955,I199433,I199450,I199467,I198958,I198961,I199512,I199529,I198949,I199593_rst,I199610,I199627,I199644,I199661,I199555,I199692,I199709,I199726,I199743,I199760,I199777,I199564,I199808,I199558,I199839,I199856,I199873,I199890,I199585,I199582,I199935,I199952,I199969,I199579,I200000,I199576,I199567,I200045,I200062,I200079,I199570,I199573,I200124,I200141,I199561,I200205_rst,I200222,I200239,I200256,I200273,I200173,I200304,I200321,I200338,I200176,I200369,I200170,I200400,I200417,I200434,I200451,I200468,I200179,I200499,I200516,I200533,I200550,I200185,I200188,I200167,I200609,I200626,I200643,I200197,I200194,I200688,I200705,I200182,I200191,I200783_rst,I200800,I200817,I200834,I200851,I200751,I200882,I200899,I200916,I200754,I200947,I200748,I200978,I200995,I201012,I201029,I201046,I200757,I201077,I201094,I201111,I201128,I200763,I200766,I200745,I201187,I201204,I201221,I200775,I200772,I201266,I201283,I200760,I200769,I201361_rst,I201378,I201395,I201412,I201429,I201329,I201460,I201477,I201494,I201332,I201525,I201326,I201556,I201573,I201590,I201607,I201624,I201335,I201655,I201672,I201689,I201706,I201341,I201344,I201323,I201765,I201782,I201799,I201353,I201350,I201844,I201861,I201338,I201347,I201939_rst,I201956,I201973,I201990,I202007,I201907,I202038,I202055,I202072,I201910,I202103,I201904,I202134,I202151,I202168,I202185,I202202,I201913,I202233,I202250,I202267,I202284,I201919,I201922,I201901,I202343,I202360,I202377,I201931,I201928,I202422,I202439,I201916,I201925,I202517_rst,I202534,I202551,I202568,I202585,I202485,I202616,I202633,I202650,I202488,I202681,I202482,I202712,I202729,I202746,I202763,I202780,I202491,I202811,I202828,I202845,I202862,I202497,I202500,I202479,I202921,I202938,I202955,I202509,I202506,I203000,I203017,I202494,I202503,I203095_rst,I203112,I203129,I203146,I203163,I203063,I203194,I203211,I203228,I203066,I203259,I203060,I203290,I203307,I203324,I203341,I203358,I203069,I203389,I203406,I203423,I203440,I203075,I203078,I203057,I203499,I203516,I203533,I203087,I203084,I203578,I203595,I203072,I203081,I203673_rst,I203690,I203707,I203724,I203741,I203641,I203772,I203789,I203806,I203644,I203837,I203638,I203868,I203885,I203902,I203919,I203936,I203647,I203967,I203984,I204001,I204018,I203653,I203656,I203635,I204077,I204094,I204111,I203665,I203662,I204156,I204173,I203650,I203659,I204251_rst,I204268,I204285,I204302,I204319,I204219,I204350,I204367,I204384,I204222,I204415,I204216,I204446,I204463,I204480,I204497,I204514,I204225,I204545,I204562,I204579,I204596,I204231,I204234,I204213,I204655,I204672,I204689,I204243,I204240,I204734,I204751,I204228,I204237,I204829_rst,I204846,I204863,I204880,I204897,I204797,I204928,I204945,I204962,I204800,I204993,I204794,I205024,I205041,I205058,I205075,I205092,I204803,I205123,I205140,I205157,I205174,I204809,I204812,I204791,I205233,I205250,I205267,I204821,I204818,I205312,I205329,I204806,I204815,I205407_rst,I205424,I205441,I205458,I205475,I205375,I205506,I205523,I205540,I205378,I205571,I205372,I205602,I205619,I205636,I205653,I205670,I205381,I205701,I205718,I205735,I205752,I205387,I205390,I205369,I205811,I205828,I205845,I205399,I205396,I205890,I205907,I205384,I205393,I205985_rst,I206002,I206019,I206036,I206053,I205953,I206084,I206101,I206118,I205956,I206149,I205950,I206180,I206197,I206214,I206231,I206248,I205959,I206279,I206296,I206313,I206330,I205965,I205968,I205947,I206389,I206406,I206423,I205977,I205974,I206468,I206485,I205962,I205971,I206563_rst,I206580,I206597,I206614,I206631,I206531,I206662,I206679,I206696,I206534,I206727,I206528,I206758,I206775,I206792,I206809,I206826,I206537,I206857,I206874,I206891,I206908,I206543,I206546,I206525,I206967,I206984,I207001,I206555,I206552,I207046,I207063,I206540,I206549,I207141_rst,I207158,I207175,I207192,I207209,I207109,I207240,I207257,I207274,I207291,I207308,I207325,I207342,I207359,I207115,I207106,I207404,I207421,I207130,I207452,I207469,I207118,I207500,I207517,I207124,I207548,I207112,I207579,I207103,I207610,I207627,I207133,I207658,I207127,I207689,I207121,I207753_rst,I207770,I207787,I207804,I207821,I207721,I207852,I207869,I207886,I207903,I207920,I207937,I207954,I207971,I207727,I207718,I208016,I208033,I207742,I208064,I208081,I207730,I208112,I208129,I207736,I208160,I207724,I208191,I207715,I208222,I208239,I207745,I208270,I207739,I208301,I207733,I208365_rst,I208382,I208399,I208416,I208433,I208333,I208464,I208481,I208498,I208515,I208532,I208549,I208566,I208583,I208339,I208330,I208628,I208645,I208354,I208676,I208693,I208342,I208724,I208741,I208348,I208772,I208336,I208803,I208327,I208834,I208851,I208357,I208882,I208351,I208913,I208345,I208977_rst,I208994,I209011,I209028,I208966,I209059,I209076,I209093,I209110,I209127,I209144,I209161,I208951,I209192,I208948,I209223,I208960,I209254,I209271,I209288,I208954,I208969,I209333,I209350,I208939,I209381,I208957,I209412,I209429,I208963,I209460,I209477,I208942,I208945,I209555_rst,I209572,I209589,I209606,I209623,I209640,I209538,I209671,I209688,I209705,I209541,I209523,I209750,I209767,I209784,I209544,I209535,I209829,I209846,I209863,I209526,I209894,I209911,I209517,I209942,I209959,I209976,I209547,I210007,I210024,I210041,I210058,I209532,I209529,I209520,I210150_rst,I210167,I210184,I210201,I210218,I210235,I210133,I210266,I210283,I210300,I210136,I210118,I210345,I210362,I210379,I210139,I210130,I210424,I210441,I210458,I210121,I210489,I210506,I210112,I210537,I210554,I210571,I210142,I210602,I210619,I210636,I210653,I210127,I210124,I210115,I210745_rst,I210762,I210779,I210796,I210813,I210830,I210728,I210861,I210878,I210895,I210731,I210713,I210940,I210957,I210974,I210734,I210725,I211019,I211036,I211053,I210716,I211084,I211101,I210707,I211132,I211149,I211166,I210737,I211197,I211214,I211231,I211248,I210722,I210719,I210710,I211340_rst,I211357,I211374,I211391,I211408,I211425,I211323,I211456,I211473,I211490,I211326,I211308,I211535,I211552,I211569,I211329,I211320,I211614,I211631,I211648,I211311,I211679,I211696,I211302,I211727,I211744,I211761,I211332,I211792,I211809,I211826,I211843,I211317,I211314,I211305,I211935_rst,I211952,I211969,I211986,I212003,I212020,I211918,I212051,I212068,I212085,I211921,I211903,I212130,I212147,I212164,I211924,I211915,I212209,I212226,I212243,I211906,I212274,I212291,I211897,I212322,I212339,I212356,I211927,I212387,I212404,I212421,I212438,I211912,I211909,I211900,I212530_rst,I212547,I212564,I212581,I212598,I212615,I212513,I212646,I212663,I212680,I212516,I212498,I212725,I212742,I212759,I212519,I212510,I212804,I212821,I212838,I212501,I212869,I212886,I212492,I212917,I212934,I212951,I212522,I212982,I212999,I213016,I213033,I212507,I212504,I212495,I213125_rst,I213142,I213159,I213176,I213193,I213210,I213108,I213241,I213258,I213275,I213111,I213093,I213320,I213337,I213354,I213114,I213105,I213399,I213416,I213433,I213096,I213464,I213481,I213087,I213512,I213529,I213546,I213117,I213577,I213594,I213611,I213628,I213102,I213099,I213090,I213720_rst,I213737,I213754,I213771,I213788,I213805,I213703,I213836,I213853,I213870,I213706,I213688,I213915,I213932,I213949,I213709,I213700,I213994,I214011,I214028,I213691,I214059,I214076,I213682,I214107,I214124,I214141,I213712,I214172,I214189,I214206,I214223,I213697,I213694,I213685,I214315_rst,I214332,I214349,I214366,I214383,I214400,I214417,I214286,I214448,I214465,I214482,I214499,I214516,I214533,I214550,I214283,I214277,I214595,I214612,I214629,I214304,I214660,I214677,I214295,I214289,I214722,I214292,I214753,I214770,I214307,I214801,I214301,I214298,I214846,I214280,I214910_rst,I214927,I214944,I214961,I214978,I214995,I215012,I214881,I215043,I215060,I215077,I215094,I215111,I215128,I215145,I214878,I214872,I215190,I215207,I215224,I214899,I215255,I215272,I214890,I214884,I215317,I214887,I215348,I215365,I214902,I215396,I214896,I214893,I215441,I214875,I215505_rst,I215522,I215539,I215556,I215573,I215590,I215607,I215476,I215638,I215655,I215672,I215689,I215706,I215723,I215740,I215473,I215467,I215785,I215802,I215819,I215494,I215850,I215867,I215485,I215479,I215912,I215482,I215943,I215960,I215497,I215991,I215491,I215488,I216036,I215470,I216100_rst,I216117,I216134,I216151,I216168,I216185,I216202,I216071,I216233,I216250,I216267,I216284,I216301,I216318,I216335,I216068,I216062,I216380,I216397,I216414,I216089,I216445,I216462,I216080,I216074,I216507,I216077,I216538,I216555,I216092,I216586,I216086,I216083,I216631,I216065,I216695_rst,I216712,I216729,I216746,I216763,I216780,I216797,I216666,I216828,I216845,I216862,I216879,I216896,I216913,I216930,I216663,I216657,I216975,I216992,I217009,I216684,I217040,I217057,I216675,I216669,I217102,I216672,I217133,I217150,I216687,I217181,I216681,I216678,I217226,I216660,I217290_rst,I217307,I217324,I217341,I217358,I217375,I217392,I217261,I217423,I217440,I217457,I217474,I217491,I217508,I217525,I217258,I217252,I217570,I217587,I217604,I217279,I217635,I217652,I217270,I217264,I217697,I217267,I217728,I217745,I217282,I217776,I217276,I217273,I217821,I217255,I217885_rst,I217902,I217919,I217936,I217953,I217970,I217987,I218004,I218021,I218038,I218055,I218072,I218089,I218106,I217874,I218137,I218154,I218171,I217847,I218202,I217868,I218233,I218250,I217853,I218281,I217850,I217856,I218326,I218343,I218360,I217862,I217877,I217865,I218419,I218436,I217871,I217859,I218514_rst,I218531,I218548,I218565,I218582,I218599,I218616,I218633,I218650,I218667,I218684,I218701,I218718,I218735,I218503,I218766,I218783,I218800,I218476,I218831,I218497,I218862,I218879,I218482,I218910,I218479,I218485,I218955,I218972,I218989,I218491,I218506,I218494,I219048,I219065,I218500,I218488,I219143_rst,I219160,I219177,I219194,I219211,I219228,I219245,I219262,I219279,I219296,I219313,I219330,I219347,I219364,I219132,I219395,I219412,I219429,I219105,I219460,I219126,I219491,I219508,I219111,I219539,I219108,I219114,I219584,I219601,I219618,I219120,I219135,I219123,I219677,I219694,I219129,I219117,I219772_rst,I219789,I219806,I219823,I219840,I219857,I219874,I219891,I219908,I219925,I219942,I219959,I219976,I219993,I219761,I220024,I220041,I220058,I219734,I220089,I219755,I220120,I220137,I219740,I220168,I219737,I219743,I220213,I220230,I220247,I219749,I219764,I219752,I220306,I220323,I219758,I219746,I220401_rst,I220418,I220435,I220452,I220469,I220486,I220503,I220520,I220537,I220554,I220571,I220588,I220605,I220622,I220390,I220653,I220670,I220687,I220363,I220718,I220384,I220749,I220766,I220369,I220797,I220366,I220372,I220842,I220859,I220876,I220378,I220393,I220381,I220935,I220952,I220387,I220375,I221030_rst,I221047,I221064,I221081,I221098,I221115,I221132,I221149,I221166,I221183,I221200,I221217,I221234,I221251,I221019,I221282,I221299,I221316,I220992,I221347,I221013,I221378,I221395,I220998,I221426,I220995,I221001,I221471,I221488,I221505,I221007,I221022,I221010,I221564,I221581,I221016,I221004,I221659_rst,I221676,I221693,I221710,I221648,I221741,I221636,I221772,I221789,I221806,I221823,I221840,I221639,I221871,I221624,I221902,I221919,I221936,I221953,I221970,I221987,I221630,I222018,I222035,I222052,I221642,I221651,I221621,I222111,I221645,I221633,I222156,I222173,I221627,I222237_rst,I222254,I222271,I222288,I222226,I222319,I222214,I222350,I222367,I222384,I222401,I222418,I222217,I222449,I222202,I222480,I222497,I222514,I222531,I222548,I222565,I222208,I222596,I222613,I222630,I222220,I222229,I222199,I222689,I222223,I222211,I222734,I222751,I222205,I222815_rst,I222832,I222849,I222866,I222804,I222897,I222792,I222928,I222945,I222962,I222979,I222996,I222795,I223027,I222780,I223058,I223075,I223092,I223109,I223126,I223143,I222786,I223174,I223191,I223208,I222798,I222807,I222777,I223267,I222801,I222789,I223312,I223329,I222783,I223393_rst,I223410,I223427,I223444,I223382,I223475,I223370,I223506,I223523,I223540,I223557,I223574,I223373,I223605,I223358,I223636,I223653,I223670,I223687,I223704,I223721,I223364,I223752,I223769,I223786,I223376,I223385,I223355,I223845,I223379,I223367,I223890,I223907,I223361,I223971_rst,I223988,I224005,I224022,I223960,I224053,I223948,I224084,I224101,I224118,I224135,I224152,I223951,I224183,I223936,I224214,I224231,I224248,I224265,I224282,I224299,I223942,I224330,I224347,I22436_rst4,I223954,I223963,I223933,I224423,I223957,I223945,I224468,I224485,I223939,I224549_rst,I224566,I224583,I224600,I224538,I224631,I224526,I224662,I224679,I224696,I224713,I224730,I224529,I224761,I224514,I224792,I224809,I224826,I224843,I224860,I224877,I224520,I224908,I224925,I224942,I224532,I224541,I224511,I225001,I224535,I224523,I225046,I225063,I224517,I225127_rst,I225144,I225161,I225178,I225116,I225209,I225104,I225240,I225257,I225274,I225291,I225308,I225107,I225339,I225092,I225370,I225387,I225404,I225421,I225438,I225455,I225098,I225486,I225503,I225520,I225110,I225119,I225089,I225579,I225113,I225101,I225624,I225641,I225095,I225705_rst,I225722,I225739,I225756,I225694,I225787,I225682,I225818,I225835,I225852,I225869,I225886,I225685,I225917,I225670,I225948,I225965,I225982,I225999,I226016,I226033,I225676,I226064,I226081,I226098,I225688,I225697,I225667,I226157,I225691,I225679,I226202,I226219,I225673,I226283_rst,I226300,I226317,I226334,I226351,I226368,I226266,I226254,I226413,I226430,I226447,I226464,I226481,I226263,I226512,I226529,I226546,I226563,I226272,I226251,I226608,I226625,I226269,I226656,I226260,I226275,I226701,I226718,I226735,I226752,I226248,I226257,I226245,I226844_rst,I226861,I226878,I226895,I226912,I226929,I226827,I226815,I226974,I226991,I227008,I227025,I227042,I226824,I227073,I227090,I227107,I227124,I226833,I226812,I227169,I227186,I226830,I227217,I226821,I226836,I227262,I227279,I227296,I227313,I226809,I226818,I226806,I227405_rst,I227422,I227439,I227456,I227473,I227490,I227388,I227376,I227535,I227552,I227569,I227586,I227603,I227385,I227634,I227651,I227668,I227685,I227394,I227373,I227730,I227747,I227391,I227778,I227382,I227397,I227823,I227840,I227857,I227874,I227370,I227379,I227367,I227966_rst,I227983,I228000,I228017,I228034,I228051,I227949,I227937,I228096,I228113,I228130,I228147,I228164,I227946,I228195,I228212,I228229,I228246,I227955,I227934,I228291,I228308,I227952,I228339,I227943,I227958,I228384,I228401,I228418,I228435,I227931,I227940,I227928,I228527_rst,I228544,I228561,I228578,I228501,I228609,I228626,I228516,I228498,I228671,I228688,I228705,I228722,I228739,I228756,I228773,I228790,I228807,I228513,I228838,I228855,I228872,I228495,I228903,I228492,I228934,I228951,I228968,I228985,I228507,I229016,I228504,I229047,I229064,I229081,I228510,I228519,I228489,I229173_rst,I229190,I229207,I229224,I229147,I229255,I229272,I229162,I229144,I229317,I229334,I229351,I229368,I229385,I229402,I229419,I229436,I229453,I229159,I229484,I229501,I229518,I229141,I229549,I229138,I229580,I229597,I229614,I229631,I229153,I229662,I229150,I229693,I229710,I229727,I229156,I229165,I229135,I229819_rst,I229836,I229853,I229870,I229793,I229901,I229918,I229808,I229790,I229963,I229980,I229997,I230014,I230031,I230048,I230065,I230082,I230099,I229805,I230130,I230147,I230164,I229787,I230195,I229784,I230226,I230243,I230260,I230277,I229799,I230308,I229796,I230339,I230356,I230373,I229802,I229811,I229781,I230465_rst,I23048_rst2,I230499,I230516,I230439,I230547,I230564,I230454,I230436,I230609,I230626,I230643,I230660,I230677,I230694,I230711,I230728,I230745,I230451,I230776,I230793,I230810,I230433,I230841,I230430,I230872,I230889,I230906,I230923,I230445,I230954,I230442,I230985,I231002,I231019,I230448,I230457,I230427,I231111_rst,I231128,I231145,I231162,I231085,I231193,I231210,I231100,I231082,I231255,I231272,I231289,I231306,I231323,I231340,I231357,I231374,I231391,I231097,I231422,I231439,I231456,I231079,I231487,I231076,I231518,I231535,I231552,I231569,I231091,I231600,I231088,I231631,I231648,I231665,I231094,I231103,I231073,I231757_rst,I231774,I231791,I231808,I231731,I231839,I231856,I231746,I231728,I231901,I231918,I231935,I231952,I231969,I231986,I232003,I232020,I232037,I231743,I232068,I232085,I232102,I231725,I232133,I231722,I232164,I232181,I232198,I232215,I231737,I232246,I231734,I232277,I232294,I232311,I231740,I231749,I231719,I232403_rst,I232420,I232437,I232454,I232377,I232485,I232502,I232392,I232374,I232547,I232564,I232581,I232598,I232615,I232632,I232649,I232666,I232683,I232389,I232714,I232731,I232748,I232371,I232779,I232368,I232810,I232827,I232844,I232861,I232383,I232892,I232380,I232923,I232940,I232957,I232386,I232395,I232365,I233049_rst,I233066,I233083,I233100,I233023,I233131,I233148,I233038,I233020,I233193,I233210,I233227,I233244,I233261,I233278,I233295,I233312,I233329,I233035,I233360,I233377,I233394,I233017,I233425,I233014,I233456,I233473,I233490,I233507,I233029,I233538,I233026,I233569,I233586,I233603,I233032,I233041,I233011,I233695_rst,I233712,I233729,I233746,I233669,I233777,I233794,I233684,I233666,I233839,I233856,I233873,I233890,I233907,I233924,I233941,I233958,I233975,I233681,I234006,I234023,I234040,I233663,I234071,I233660,I234102,I234119,I234136,I234153,I233675,I234184,I233672,I234215,I234232,I234249,I233678,I233687,I233657,I234341_rst,I234358,I234375,I234392,I234315,I234423,I234440,I234330,I234312,I234485,I234502,I234519,I234536,I234553,I234570,I234587,I234604,I234621,I234327,I234652,I234669,I234686,I234309,I234717,I234306,I234748,I234765,I234782,I234799,I234321,I234830,I234318,I234861,I234878,I234895,I234324,I234333,I234303,I234987_rst,I235004,I235021,I235038,I234961,I235069,I235086,I234976,I234958,I235131,I235148,I235165,I235182,I235199,I235216,I235233,I235250,I235267,I234973,I235298,I235315,I235332,I234955,I235363,I234952,I235394,I235411,I235428,I235445,I234967,I235476,I234964,I235507,I235524,I235541,I234970,I234979,I234949,I235633_rst,I235650,I235667,I235684,I235607,I235715,I235732,I235622,I235604,I235777,I235794,I235811,I235828,I235845,I235862,I235879,I235896,I235913,I235619,I235944,I235961,I235978,I235601,I236009,I235598,I236040,I236057,I236074,I236091,I235613,I236122,I235610,I236153,I236170,I236187,I235616,I235625,I235595,I236279_rst,I236296,I236313,I236330,I236253,I236361,I236378,I23626_rst8,I236250,I236423,I236440,I236457,I236474,I236491,I236508,I236525,I236542,I236559,I23626_rst5,I236590,I236607,I236624,I236247,I236655,I236244,I236686,I236703,I236720,I236737,I236259,I236768,I236256,I236799,I236816,I236833,I23626_rst2,I236271,I236241,I236925_rst,I236942,I236959,I236976,I236896,I237007,I237024,I237041,I237058,I237075,I237092,I237109,I237126,I237143,I237160,I236911,I236908,I237205,I236893,I237236,I236890,I237267,I237284,I237301,I237318,I237335,I237352,I236917,I237383,I236905,I236899,I237428,I237445,I236914,I237476,I237493,I237510,I236902,I236887,I237588_rst,I237605,I237622,I237639,I237559,I237670,I237687,I237704,I237721,I237738,I237755,I237772,I237789,I237806,I237823,I237574,I237571,I237868,I237556,I237899,I237553,I237930,I237947,I237964,I237981,I237998,I238015,I237580,I238046,I237568,I237562,I238091,I238108,I237577,I238139,I238156,I238173,I237565,I237550,I238251_rst,I238268,I238285,I238302,I238222,I238333,I238350,I238367,I238384,I238401,I238418,I238435,I238452,I238469,I238486,I238237,I238234,I238531,I238219,I238562,I238216,I238593,I238610,I238627,I238644,I238661,I238678,I238243,I238709,I238231,I238225,I238754,I238771,I238240,I238802,I238819,I238836,I238228,I238213,I238914_rst,I238931,I238948,I238965,I238885,I238996,I239013,I239030,I239047,I239064,I239081,I239098,I239115,I239132,I239149,I238900,I238897,I239194,I238882,I239225,I238879,I239256,I239273,I239290,I239307,I239324,I239341,I238906,I239372,I238894,I238888,I239417,I239434,I238903,I239465,I239482,I239499,I238891,I238876,I239577_rst,I239594,I239611,I239628,I239548,I239659,I239676,I239693,I239710,I239727,I239744,I239761,I239778,I239795,I239812,I239563,I239560,I239857,I239545,I239888,I239542,I239919,I239936,I239953,I239970,I239987,I240004,I239569,I240035,I239557,I239551,I240080,I240097,I239566,I240128,I240145,I240162,I239554,I239539,I240240_rst,I240257,I240274,I240214,I240305,I240322,I240339,I240356,I240373,I240390,I240407,I240424,I240441,I240208,I240472,I240489,I240205,I240520,I240537,I240554,I240217,I240202,I240599,I240616,I240633,I240650,I240667,I240223,I240698,I240232,I240729,I240226,I240229,I240220,I240211,I240835_rst,I240852,I240869,I240809,I240900,I240917,I240934,I240951,I240968,I240985,I241002,I241019,I241036,I240803,I241067,I241084,I240800,I241115,I241132,I241149,I240812,I240797,I241194,I241211,I241228,I241245,I241262,I240818,I241293,I240827,I241324,I240821,I240824,I240815,I240806,I241430_rst,I241447,I241464,I241404,I241495,I241512,I241529,I241546,I241563,I241580,I241597,I241614,I241631,I241398,I241662,I241679,I241395,I241710,I241727,I241744,I241407,I241392,I241789,I241806,I241823,I241840,I241857,I241413,I241888,I241422,I241919,I241416,I241419,I241410,I241401,I242025_rst,I24204_rst2,I242059,I241999,I242090,I242107,I242124,I242141,I242158,I242175,I242192,I242209,I242226,I241993,I242257,I242274,I241990,I242305,I242322,I242339,I242002,I241987,I242384,I242401,I242418,I242435,I242452,I242008,I242483,I242017,I242514,I242011,I242014,I242005,I241996,I242620_rst,I242637,I242603,I242582,I242682,I242699,I242716,I242733,I242750,I242767,I242784,I242801,I242818,I242609,I242849,I242866,I242883,I242900,I242612,I242931,I242948,I242965,I242982,I242999,I242597,I243030,I243047,I242600,I242594,I242588,I243106,I242606,I243137,I242591,I242585,I243215_rst,I243232,I243198,I243177,I243277,I243294,I243311,I243328,I243345,I243362,I243379,I243396,I243413,I243204,I243444,I243461,I243478,I243495,I243207,I243526,I243543,I243560,I243577,I243594,I243192,I243625,I243642,I243195,I243189,I243183,I243701,I243201,I243732,I243186,I243180,I243810_rst,I243827,I243844,I243861,I243878,I243895,I243912,I243929,I243799,I243960,I243784,I243991,I244008,I244025,I244042,I244059,I244076,I244093,I243781,I244124,I244141,I243778,I244172,I244189,I243796,I244220,I243793,I244251,I244268,I243772,I243775,I244313,I244330,I244347,I244364,I243802,I244395,I243787,I243790,I244473_rst,I244490,I244507,I244524,I244541,I244558,I244575,I244592,I244462,I244623,I244447,I244654,I244671,I244688,I244705,I244722,I244739,I244756,I244444,I244787,I244804,I244441,I244835,I244852,I244459,I244883,I244456,I244914,I244931,I244435,I244438,I244976,I244993,I245010,I245027,I244465,I245058,I244450,I244453,I245136_rst,I245153,I245170,I245187,I245204,I245221,I245238,I245255,I245125,I245286,I245110,I245317,I245334,I245351,I245368,I245385,I245402,I245419,I245107,I245450,I245467,I245104,I245498,I245515,I245122,I245546,I245119,I245577,I245594,I245098,I245101,I245639,I245656,I245673,I245690,I245128,I245721,I245113,I245116,I245799_rst,I245816,I245833,I245850,I245867,I245884,I245901,I245918,I245788,I245949,I245773,I245980,I245997,I246014,I246031,I246048,I246065,I246082,I245770,I246113,I246130,I245767,I246161,I246178,I245785,I246209,I245782,I246240,I246257,I245761,I245764,I246302,I246319,I246336,I246353,I245791,I246384,I245776,I245779,I246462_rst,I246479,I246496,I246513,I246530,I246547,I246564,I246581,I246451,I246612,I246436,I246643,I246660,I246677,I246694,I246711,I246728,I246745,I246433,I246776,I246793,I246430,I246824,I246841,I246448,I246872,I246445,I246903,I246920,I246424,I246427,I246965,I246982,I246999,I247016,I246454,I247047,I246439,I246442,I247125_rst,I247142,I247159,I247176,I247193,I247210,I247227,I247244,I247114,I247275,I247099,I247306,I247323,I247340,I247357,I247374,I247391,I247408,I247096,I247439,I247456,I247093,I247487,I247504,I247111,I247535,I247108,I247566,I247583,I247087,I247090,I247628,I247645,I247662,I247679,I247117,I247710,I247102,I247105,I247788_rst,I247805,I24782_rst2,I247839,I247856,I247873,I247890,I247907,I247777,I247938,I247762,I247969,I247986,I248003,I248020,I248037,I248054,I248071,I247759,I248102,I248119,I247756,I248150,I248167,I247774,I248198,I247771,I248229,I248246,I247750,I247753,I248291,I248308,I248325,I248342,I247780,I248373,I247765,I247768,I248451_rst,I248468,I248485,I248502,I248519,I248536,I248553,I248570,I248440,I248601,I248425,I248632,I248649,I248666,I248683,I248700,I248717,I248734,I248422,I248765,I248782,I248419,I248813,I248830,I248437,I248861,I248434,I248892,I248909,I248413,I248416,I248954,I248971,I248988,I249005,I248443,I249036,I248428,I248431,I249114_rst,I249131,I249148,I249165,I249182,I249199,I249216,I249233,I249103,I249264,I249088,I249295,I249312,I249329,I249346,I249363,I249380,I249397,I249085,I249428,I249445,I249082,I249476,I249493,I249100,I249524,I249097,I249555,I249572,I249076,I249079,I249617,I249634,I249651,I249668,I249106,I249699,I249091,I249094,I249777_rst,I249794,I249811,I249828,I249845,I249862,I249879,I249896,I249766,I249927,I249751,I249958,I249975,I249992,I250009,I250026,I250043,I250060,I249748,I250091,I250108,I249745,I250139,I250156,I249763,I250187,I249760,I250218,I250235,I249739,I249742,I250280,I250297,I250314,I250331,I249769,I250362,I249754,I249757,I250440_rst,I250457,I250474,I250491,I250508,I250525,I250542,I250559,I250429,I250590,I250414,I250621,I250638,I250655,I250672,I250689,I250706,I250723,I250411,I250754,I250771,I250408,I250802,I250819,I250426,I250850,I250423,I250881,I250898,I250402,I250405,I250943,I250960,I250977,I250994,I250432,I251025,I250417,I250420,I251103_rst,I251120,I251137,I251154,I251171,I251188,I251205,I251222,I251092,I251253,I251077,I251284,I251301,I251318,I251335,I251352,I251369,I251386,I251074,I251417,I251434,I251071,I251465,I251482,I251089,I251513,I251086,I251544,I251561,I251065,I251068,I251606,I251623,I251640,I251657,I251095,I251688,I251080,I251083,I251766_rst,I251783,I251800,I251817,I251834,I251851,I251868,I251885,I251755,I251916,I251740,I251947,I251964,I251981,I251998,I252015,I252032,I252049,I251737,I252080,I252097,I251734,I252128,I252145,I251752,I252176,I251749,I252207,I252224,I251728,I251731,I252269,I252286,I252303,I252320,I251758,I252351,I251743,I251746,I252429_rst,I252446,I252463,I252480,I252497,I252514,I252531,I252400,I252562,I252579,I252596,I252613,I252630,I252647,I252664,I252397,I252695,I252391,I252726,I252743,I252760,I252421,I252394,I252805,I252418,I252836,I252415,I252412,I252881,I252898,I252915,I252932,I252949,I252406,I252980,I252997,I252409,I252403,I253075_rst,I253092,I253109,I253126,I253143,I253160,I253177,I253046,I253208,I253225,I253242,I253259,I253276,I253293,I253310,I253043,I253341,I253037,I253372,I253389,I253406,I253067,I253040,I253451,I253064,I253482,I253061,I253058,I253527,I253544,I253561,I253578,I253595,I253052,I253626,I253643,I253055,I253049,I253721_rst,I253738,I253755,I253772,I253789,I253806,I253823,I253692,I253854,I253871,I253888,I253905,I253922,I253939,I253956,I253689,I253987,I253683,I254018,I254035,I254052,I253713,I253686,I254097,I253710,I254128,I253707,I253704,I254173,I254190,I254207,I254224,I254241,I253698,I254272,I254289,I253701,I253695,I254367_rst,I254384,I254401,I254418,I254435,I254452,I254469,I254338,I254500,I254517,I254534,I254551,I254568,I254585,I254602,I254335,I254633,I254329,I254664,I254681,I254698,I254359,I254332,I254743,I254356,I254774,I254353,I254350,I254819,I254836,I254853,I254870,I254887,I254344,I254918,I254935,I254347,I254341,I255013_rst,I255030,I255047,I255064,I255081,I255098,I255115,I254984,I255146,I255163,I255180,I255197,I255214,I255231,I255248,I254981,I255279,I254975,I255310,I255327,I255344,I255005,I254978,I255389,I255002,I255420,I254999,I254996,I255465,I255482,I255499,I255516,I255533,I254990,I255564,I255581,I254993,I254987,I255659_rst,I255676,I255693,I255710,I255727,I255744,I255761,I255630,I255792,I255809,I255826,I255843,I255860,I255877,I255894,I255627,I255925,I255621,I255956,I255973,I255990,I255651,I255624,I256035,I255648,I256066,I255645,I255642,I256111,I256128,I256145,I256162,I256179,I255636,I256210,I256227,I255639,I255633,I256305_rst,I256322,I256339,I256356,I256373,I256390,I256407,I256276,I256438,I256455,I256472,I256489,I256506,I256523,I256540,I256273,I256571,I256267,I256602,I256619,I256636,I256297,I256270,I256681,I256294,I256712,I256291,I256288,I256757,I256774,I256791,I256808,I256825,I256282,I256856,I256873,I256285,I256279,I256951_rst,I256968,I256985,I257002,I257019,I257036,I257053,I256922,I257084,I257101,I257118,I257135,I257152,I257169,I257186,I256919,I257217,I256913,I257248,I257265,I257282,I256943,I256916,I257327,I256940,I257358,I256937,I256934,I257403,I257420,I257437,I257454,I257471,I256928,I257502,I257519,I256931,I256925,I257597_rst,I257614,I257631,I257648,I257665,I257682,I257699,I257568,I257730,I257747,I257764,I257781,I257798,I257815,I257832,I257565,I257863,I257559,I257894,I257911,I257928,I257589,I257562,I257973,I257586,I258004,I257583,I257580,I258049,I258066,I258083,I258100,I258117,I257574,I258148,I258165,I257577,I257571,I258243_rst,I258260,I258277,I258294,I258311,I258328,I258345,I258214,I258376,I258393,I258410,I258427,I258444,I258461,I258478,I258211,I258509,I258205,I258540,I258557,I258574,I258235,I258208,I258619,I258232,I258650,I258229,I258226,I258695,I258712,I258729,I258746,I258763,I258220,I258794,I258811,I258223,I258217,I258889_rst,I258906,I258923,I258940,I258957,I258851,I258988,I259005,I259022,I259039,I259056,I259073,I258860,I259104,I258854,I259135,I259152,I259169,I259186,I258881,I258878,I259231,I259248,I259265,I258875,I259296,I258872,I258863,I259341,I259358,I259375,I258866,I258869,I259420,I259437,I258857,I259501_rst,I259518,I259535,I259552,I259569,I259469,I259600,I259617,I259634,I259472,I259665,I259466,I259696,I259713,I259730,I259747,I259764,I259475,I259795,I259812,I259829,I259846,I259481,I259484,I259463,I259905,I259922,I259939,I259493,I259490,I259984,I260001,I259478,I259487,I260079_rst,I260096,I260113,I260130,I260147,I260047,I260178,I260195,I260212,I260050,I260243,I260044,I260274,I260291,I260308,I260325,I260342,I260053,I260373,I260390,I260407,I260424,I260059,I260062,I260041,I260483,I260500,I260517,I260071,I260068,I260562,I260579,I260056,I260065,I260657_rst,I260674,I260691,I260708,I260725,I260756,I260773,I260790,I260821,I260852,I260869,I260886,I260903,I260920,I260951,I260968,I260985,I261002,I261061,I261078,I261095,I261140,I261157,I261235_rst,I261252,I261269,I261286,I261303,I261203,I261334,I261351,I261368,I261206,I261399,I261200,I261430,I261447,I261464,I261481,I261498,I261209,I261529,I261546,I261563,I261580,I261215,I261218,I261197,I261639,I261656,I261673,I261227,I261224,I261718,I261735,I261212,I261221,I261813_rst,I261830,I261847,I261864,I261881,I261781,I261912,I261929,I261946,I261784,I261977,I261778,I262008,I262025,I262042,I262059,I262076,I261787,I262107,I262124,I262141,I262158,I261793,I261796,I261775,I262217,I262234,I262251,I261805,I261802,I262296,I262313,I261790,I261799,I262391_rst,I262408,I262425,I262442,I262459,I262359,I262490,I262507,I262524,I262362,I262555,I262356,I262586,I262603,I262620,I262637,I262654,I262365,I262685,I262702,I262719,I262736,I262371,I262374,I262353,I262795,I262812,I262829,I262383,I262380,I262874,I262891,I262368,I262377,I262969_rst,I262986,I263003,I263020,I263037,I262937,I263068,I263085,I263102,I262940,I263133,I262934,I263164,I263181,I263198,I263215,I263232,I262943,I263263,I263280,I263297,I263314,I262949,I262952,I262931,I263373,I263390,I263407,I262961,I262958,I263452,I263469,I262946,I262955,I263547_rst,I263564,I263581,I263598,I263615,I263515,I263646,I263663,I263680,I263518,I263711,I263512,I263742,I263759,I263776,I263793,I263810,I263521,I263841,I263858,I263875,I263892,I263527,I263530,I263509,I263951,I263968,I263985,I263539,I263536,I264030,I264047,I263524,I263533,I264125_rst,I264142,I264159,I264176,I264193,I264093,I264224,I264241,I264258,I264096,I264289,I264090,I264320,I264337,I264354,I264371,I264388,I264099,I264419,I264436,I264453,I264470,I264105,I264108,I264087,I264529,I264546,I264563,I264117,I264114,I264608,I264625,I264102,I264111,I264703_rst,I264720,I264737,I264754,I264771,I264671,I264802,I264819,I264836,I264674,I264867,I264668,I264898,I264915,I264932,I264949,I264966,I264677,I264997,I265014,I265031,I265048,I264683,I264686,I264665,I265107,I265124,I265141,I264695,I264692,I265186,I265203,I264680,I264689,I265281_rst,I265298,I265315,I265332,I265349,I265249,I265380,I265397,I265414,I265252,I265445,I265246,I265476,I265493,I265510,I265527,I265544,I265255,I265575,I265592,I265609,I265626,I265261,I265264,I265243,I265685,I265702,I265719,I265273,I265270,I265764,I265781,I265258,I265267,I265859_rst,I265876,I265893,I265910,I265927,I265827,I265958,I265975,I265992,I265830,I266023,I265824,I266054,I266071,I266088,I266105,I266122,I265833,I266153,I266170,I266187,I266204,I265839,I26584_rst2,I265821,I266263,I266280,I266297,I265851,I26584_rst8,I266342,I266359,I265836,I26584_rst5,I266437_rst,I266454,I266471,I266488,I266505,I266405,I266536,I266553,I266570,I266408,I266601,I266402,I266632,I266649,I266666,I266683,I266700,I266411,I266731,I266748,I266765,I266782,I266417,I266420,I266399,I266841,I266858,I266875,I266429,I266426,I266920,I266937,I266414,I266423,I267015_rst,I267032,I267049,I267066,I267083,I267100,I266998,I267131,I267148,I267165,I267001,I266983,I267210,I267227,I267244,I267004,I266995,I267289,I267306,I267323,I266986,I267354,I267371,I266977,I267402,I267419,I267436,I267007,I267467,I267484,I267501,I267518,I266992,I266989,I266980,I267610_rst,I267627,I267644,I267661,I267678,I267695,I267593,I267726,I267743,I267760,I267596,I267578,I267805,I267822,I267839,I267599,I267590,I267884,I267901,I267918,I267581,I267949,I267966,I267572,I267997,I268014,I268031,I267602,I268062,I268079,I268096,I268113,I267587,I267584,I267575,I268205_rst,I268222,I268239,I268256,I268273,I268290,I268188,I268321,I268338,I268355,I268191,I268173,I268400,I268417,I268434,I268194,I268185,I268479,I268496,I268513,I268176,I268544,I268561,I268167,I268592,I268609,I268626,I268197,I268657,I268674,I268691,I268708,I268182,I268179,I268170,I268800_rst,I268817,I268834,I268851,I268868,I268885,I268783,I268916,I268933,I268950,I268786,I268768,I268995,I269012,I269029,I268789,I268780,I269074,I269091,I269108,I268771,I269139,I269156,I268762,I269187,I269204,I269221,I268792,I269252,I269269,I269286,I269303,I268777,I268774,I268765,I269395_rst,I269412,I269429,I269446,I269463,I269480,I269378,I269511,I269528,I269545,I269381,I269363,I269590,I269607,I269624,I269384,I269375,I269669,I269686,I269703,I269366,I269734,I269751,I269357,I269782,I269799,I269816,I269387,I269847,I269864,I269881,I269898,I269372,I269369,I269360,I269990_rst,I270007,I270024,I270041,I270058,I270075,I269973,I270106,I270123,I270140,I269976,I269958,I270185,I270202,I270219,I269979,I269970,I270264,I270281,I270298,I269961,I270329,I270346,I269952,I270377,I270394,I270411,I269982,I270442,I270459,I270476,I270493,I269967,I269964,I269955,I270585_rst,I270602,I270619,I270636,I270653,I270670,I270701,I270718,I270735,I270780,I270797,I270814,I270859,I270876,I270893,I270924,I270941,I270972,I270989,I271006,I271037,I271054,I271071,I271088,I271180_rst,I271197,I271214,I271231,I271248,I271265,I271163,I271296,I271313,I271330,I271166,I271148,I271375,I271392,I271409,I271169,I271160,I271454,I271471,I271488,I271151,I271519,I271536,I271142,I271567,I271584,I271601,I271172,I271632,I271649,I271666,I271683,I271157,I271154,I271145,I271775_rst,I271792,I271809,I271826,I271843,I271860,I271758,I271891,I271908,I271925,I271761,I271743,I271970,I271987,I272004,I271764,I271755,I272049,I272066,I272083,I271746,I272114,I272131,I271737,I272162,I272179,I272196,I271767,I272227,I272244,I272261,I272278,I271752,I271749,I271740,I272370_rst,I272387,I272404,I272421,I272438,I272455,I272353,I272486,I272503,I272520,I272356,I272338,I272565,I272582,I272599,I272359,I272350,I272644,I272661,I272678,I272341,I272709,I272726,I272332,I272757,I272774,I272791,I272362,I272822,I272839,I272856,I272873,I272347,I272344,I272335,I272965_rst,I272982,I272999,I273016,I273033,I273050,I272948,I273081,I273098,I273115,I272951,I272933,I273160,I273177,I273194,I272954,I272945,I273239,I273256,I273273,I272936,I273304,I273321,I272927,I273352,I273369,I273386,I272957,I273417,I273434,I273451,I273468,I272942,I272939,I272930,I273560_rst,I273577,I273594,I273611,I273628,I273645,I273676,I273693,I273710,I273755,I273772,I273789,I273834,I273851,I273868,I273899,I273916,I273947,I273964,I273981,I274012,I274029,I274046,I274063,I274155_rst,I274172,I274189,I274206,I274223,I274240,I274138,I274271,I274288,I274305,I274141,I274123,I274350,I274367,I274384,I274144,I274135,I274429,I274446,I274463,I274126,I274494,I274511,I274117,I274542,I274559,I274576,I274147,I274607,I274624,I274641,I274658,I274132,I274129,I274120,I274750_rst,I274767,I274784,I274801,I274818,I274835,I274733,I274866,I274883,I274900,I274736,I274718,I274945,I274962,I274979,I274739,I274730,I275024,I275041,I275058,I274721,I275089,I275106,I274712,I275137,I275154,I275171,I274742,I275202,I275219,I275236,I275253,I274727,I274724,I274715,I275345_rst,I275362,I275379,I275396,I275413,I275430,I275447,I275316,I275478,I275495,I275512,I275529,I275546,I275563,I275580,I275313,I275307,I275625,I275642,I275659,I275334,I275690,I275707,I275325,I275319,I275752,I275322,I275783,I275800,I275337,I275831,I275331,I275328,I275876,I275310,I275940_rst,I275957,I275974,I275991,I276008,I276025,I276042,I275911,I276073,I276090,I276107,I276124,I276141,I276158,I276175,I275908,I275902,I276220,I276237,I276254,I275929,I276285,I276302,I275920,I275914,I276347,I275917,I276378,I276395,I275932,I276426,I275926,I275923,I276471,I275905,I276535_rst,I276552,I276569,I276586,I276603,I276620,I276637,I276506,I276668,I276685,I276702,I276719,I276736,I276753,I276770,I276503,I276497,I276815,I276832,I276849,I276524,I276880,I276897,I276515,I276509,I276942,I276512,I276973,I276990,I276527,I277021,I276521,I276518,I277066,I276500,I277130_rst,I277147,I277164,I277181,I277198,I277215,I277232,I277101,I277263,I277280,I277297,I277314,I277331,I277348,I277365,I277098,I277092,I277410,I277427,I277444,I277119,I277475,I277492,I277110,I277104,I277537,I277107,I277568,I277585,I277122,I277616,I277116,I277113,I277661,I277095,I277725_rst,I277742,I277759,I277776,I277793,I277810,I277827,I277696,I277858,I277875,I277892,I277909,I277926,I277943,I277960,I277693,I277687,I278005,I278022,I278039,I277714,I278070,I278087,I277705,I277699,I278132,I277702,I278163,I278180,I277717,I278211,I277711,I277708,I278256,I277690,I278320_rst,I278337,I278354,I278371,I278388,I278405,I278422,I278291,I278453,I278470,I278487,I278504,I278521,I278538,I278555,I278288,I278282,I278600,I278617,I278634,I278309,I278665,I278682,I278300,I278294,I278727,I278297,I278758,I278775,I278312,I278806,I278306,I278303,I278851,I278285,I278915_rst,I278932,I278949,I278966,I278983,I279000,I279017,I279034,I279051,I279068,I279085,I279102,I279119,I279136,I278904,I279167,I279184,I279201,I278877,I279232,I278898,I279263,I279280,I278883,I279311,I278880,I278886,I279356,I279373,I279390,I278892,I278907,I278895,I279449,I279466,I278901,I278889,I279544_rst,I279561,I279578,I279595,I279612,I279629,I279646,I279663,I279680,I279697,I279714,I279731,I279748,I279765,I279533,I279796,I279813,I279830,I279506,I279861,I279527,I279892,I279909,I279512,I279940,I279509,I279515,I279985,I280002,I280019,I279521,I279536,I279524,I280078,I280095,I279530,I279518,I280173_rst,I280190,I280207,I280224,I280241,I280258,I280275,I280292,I280309,I280326,I280343,I280360,I280377,I280394,I280162,I280425,I280442,I280459,I280135,I280490,I280156,I280521,I280538,I280141,I280569,I280138,I280144,I280614,I280631,I280648,I280150,I280165,I280153,I280707,I280724,I280159,I280147,I280802_rst,I280819,I280836,I280853,I280870,I280887,I280904,I280921,I280938,I280955,I280972,I280989,I281006,I281023,I280791,I281054,I281071,I281088,I280764,I281119,I280785,I281150,I281167,I280770,I281198,I280767,I280773,I281243,I281260,I281277,I280779,I280794,I280782,I281336,I281353,I280788,I280776,I281431_rst,I281448,I281465,I281482,I281499,I281516,I281533,I281550,I281567,I281584,I281601,I281618,I281635,I281652,I281420,I281683,I281700,I281717,I281393,I281748,I281414,I281779,I281796,I281399,I281827,I281396,I281402,I281872,I281889,I281906,I281408,I281423,I281411,I281965,I281982,I281417,I281405,I282060_rst,I282077,I282094,I282111,I282128,I282145,I282162,I282179,I282196,I282213,I282230,I282247,I282264,I282281,I282312,I282329,I282346,I282377,I282408,I282425,I282456,I282501,I282518,I282535,I282594,I282611,I282689_rst,I282706,I282723,I282740,I282757,I282774,I282791,I282808,I282825,I282842,I282859,I282876,I282893,I282910,I282678,I282941,I282958,I282975,I282651,I283006,I282672,I283037,I283054,I282657,I283085,I282654,I282660,I283130,I283147,I283164,I282666,I282681,I282669,I283223,I283240,I282675,I282663,I283318_rst,I283335,I283352,I283369,I283386,I283403,I283420,I283437,I283454,I283471,I283488,I283505,I28352_rst2,I283539,I283307,I283570,I283587,I283604,I283280,I283635,I283301,I283666,I283683,I283286,I283714,I283283,I283289,I283759,I283776,I283793,I283295,I283310,I283298,I283852,I283869,I283304,I283292,I283947_rst,I283964,I283981,I283998,I284015,I284032,I284049,I284066,I284083,I284100,I284117,I284134,I284151,I284168,I283936,I284199,I284216,I284233,I283909,I284264,I283930,I284295,I284312,I283915,I284343,I283912,I283918,I284388,I284405,I284422,I283924,I283939,I283927,I284481,I284498,I283933,I283921,I284576_rst,I284593,I284610,I284627,I284644,I284661,I284678,I284695,I284712,I284729,I284746,I284763,I284780,I284797,I284565,I284828,I284845,I284862,I284538,I284893,I284559,I284924,I284941,I284544,I284972,I284541,I284547,I285017,I285034,I285051,I284553,I284568,I284556,I285110,I285127,I284562,I284550,I285205_rst,I285222,I285239,I285256,I285273,I285290,I285307,I285324,I285341,I285358,I285375,I285392,I285409,I285426,I285194,I285457,I285474,I285491,I285167,I285522,I285188,I285553,I285570,I285173,I285601,I285170,I285176,I285646,I285663,I285680,I285182,I285197,I285185,I285739,I285756,I285191,I285179,I285834_rst,I285851,I285868,I285885,I285823,I285916,I285811,I285947,I285964,I285981,I285998,I286015,I285814,I286046,I285799,I286077,I286094,I286111,I286128,I286145,I286162,I285805,I286193,I286210,I286227,I285817,I285826,I285796,I286286,I285820,I285808,I286331,I286348,I285802,I286412_rst,I286429,I286446,I286463,I286401,I286494,I286389,I286525,I286542,I286559,I286576,I286593,I286392,I286624,I286377,I286655,I286672,I286689,I286706,I286723,I286740,I286383,I286771,I286788,I286805,I286395,I286404,I286374,I286864,I286398,I286386,I286909,I286926,I286380,I286990_rst,I287007,I287024,I287041,I286979,I287072,I286967,I287103,I287120,I287137,I287154,I287171,I286970,I287202,I286955,I287233,I287250,I287267,I287284,I287301,I287318,I286961,I287349,I287366,I287383,I286973,I286982,I286952,I287442,I286976,I286964,I287487,I287504,I286958,I287568_rst,I287585,I287602,I287619,I287557,I287650,I287545,I287681,I287698,I287715,I287732,I287749,I287548,I287780,I287533,I287811,I287828,I287845,I287862,I287879,I287896,I287539,I287927,I287944,I287961,I287551,I287560,I287530,I288020,I287554,I287542,I288065,I288082,I287536,I288146_rst,I288163,I288180,I288197,I288135,I288228,I288123,I288259,I288276,I288293,I288310,I288327,I288126,I288358,I288111,I288389,I288406,I288423,I288440,I288457,I288474,I288117,I288505,I288522,I288539,I288129,I288138,I288108,I288598,I288132,I288120,I288643,I288660,I288114,I288724_rst,I288741,I288758,I288775,I288792,I288809,I288707,I288695,I288854,I288871,I288888,I288905,I288922,I288704,I288953,I288970,I288987,I289004,I288713,I288692,I289049,I289066,I288710,I289097,I288701,I288716,I289142,I289159,I289176,I289193,I288689,I288698,I288686,I289285_rst,I289302,I289319,I289336,I289353,I289370,I289268,I289256,I289415,I289432,I289449,I289466,I289483,I289265,I289514,I289531,I289548,I289565,I289274,I289253,I289610,I289627,I289271,I289658,I289262,I289277,I289703,I289720,I289737,I289754,I289250,I289259,I289247,I289846_rst,I289863,I289880,I289897,I289914,I289931,I289976,I289993,I290010,I290027,I290044,I290075,I290092,I290109,I290126,I290171,I290188,I290219,I290264,I290281,I290298,I290315,I290407_rst,I290424,I290441,I290458,I290475,I290492,I290390,I290378,I290537,I290554,I290571,I290588,I290605,I290387,I290636,I290653,I290670,I290687,I290396,I290375,I290732,I290749,I290393,I290780,I290384,I290399,I290825,I290842,I290859,I290876,I290372,I290381,I290369,I290968_rst,I290985,I291002,I291019,I291036,I291053,I290951,I290939,I291098,I291115,I291132,I291149,I291166,I290948,I291197,I291214,I291231,I291248,I290957,I290936,I291293,I291310,I290954,I291341,I290945,I290960,I291386,I291403,I291420,I291437,I290933,I290942,I290930,I291529_rst,I291546,I291563,I291580,I291597,I291614,I291512,I291500,I291659,I291676,I291693,I291710,I291727,I291509,I291758,I291775,I291792,I291809,I291518,I291497,I291854,I291871,I291515,I291902,I291506,I291521,I291947,I291964,I291981,I291998,I291494,I291503,I291491,I292090_rst,I292107,I292124,I292141,I292158,I292175,I292073,I292061,I292220,I292237,I292254,I292271,I292288,I292070,I292319,I292336,I292353,I292370,I292079,I292058,I292415,I292432,I292076,I292463,I292067,I292082,I292508,I292525,I292542,I292559,I292055,I292064,I292052,I292651_rst,I292668,I292685,I292702,I292719,I292736,I292634,I292622,I292781,I292798,I292815,I292832,I292849,I292631,I292880,I292897,I292914,I292931,I292640,I292619,I292976,I292993,I292637,I293024,I292628,I292643,I293069,I293086,I293103,I293120,I292616,I292625,I292613,I293212_rst,I293229,I293246,I293263,I293280,I293297,I293195,I293183,I293342,I293359,I293376,I293393,I293410,I293192,I293441,I293458,I293475,I293492,I293201,I293180,I293537,I293554,I293198,I293585,I293189,I293204,I293630,I293647,I293664,I293681,I293177,I293186,I293174,I293773_rst,I293790,I293807,I293824,I293747,I293855,I293872,I293762,I293744,I293917,I293934,I293951,I293968,I293985,I294002,I294019,I294036,I294053,I293759,I294084,I294101,I294118,I293741,I294149,I293738,I294180,I294197,I294214,I294231,I293753,I294262,I293750,I294293,I294310,I294327,I293756,I293765,I293735,I294419_rst,I294436,I294453,I294470,I294393,I294501,I294518,I294408,I294390,I294563,I294580,I294597,I294614,I294631,I294648,I294665,I294682,I294699,I294405,I294730,I294747,I294764,I294387,I294795,I294384,I294826,I294843,I294860,I294877,I294399,I294908,I294396,I294939,I294956,I294973,I294402,I294411,I294381,I295065_rst,I295082,I295099,I295116,I295147,I295164,I295209,I295226,I295243,I295260,I295277,I295294,I295311,I295328,I295345,I295376,I295393,I295410,I295441,I295472,I295489,I295506,I295523,I295554,I295585,I295602,I295619,I295711_rst,I295728,I295745,I295762,I295685,I295793,I295810,I295700,I295682,I295855,I295872,I295889,I295906,I295923,I295940,I295957,I295974,I295991,I295697,I296022,I296039,I296056,I295679,I296087,I295676,I296118,I296135,I296152,I296169,I295691,I296200,I295688,I296231,I296248,I296265,I295694,I295703,I295673,I296357_rst,I296374,I296391,I296408,I296331,I296439,I296456,I296346,I296328,I296501,I296518,I296535,I296552,I296569,I296586,I296603,I296620,I296637,I296343,I296668,I296685,I296702,I296325,I296733,I296322,I296764,I296781,I296798,I296815,I296337,I296846,I296334,I296877,I296894,I296911,I296340,I296349,I296319,I297003_rst,I297020,I297037,I297054,I296977,I297085,I297102,I296992,I296974,I297147,I297164,I297181,I297198,I297215,I297232,I297249,I297266,I297283,I296989,I297314,I297331,I297348,I296971,I297379,I296968,I297410,I297427,I297444,I297461,I296983,I297492,I296980,I297523,I297540,I297557,I296986,I296995,I296965,I297649_rst,I297666,I297683,I297700,I297623,I297731,I297748,I297638,I297620,I297793,I297810,I297827,I297844,I297861,I297878,I297895,I297912,I297929,I297635,I297960,I297977,I297994,I297617,I298025,I297614,I298056,I298073,I298090,I298107,I297629,I298138,I297626,I298169,I298186,I298203,I297632,I297641,I297611,I298295_rst,I298312,I298329,I298346,I298269,I298377,I298394,I298284,I298266,I298439,I298456,I298473,I298490,I298507,I298524,I298541,I298558,I298575,I298281,I298606,I298623,I298640,I298263,I298671,I298260,I298702,I298719,I298736,I298753,I298275,I298784,I298272,I298815,I298832,I298849,I298278,I298287,I298257,I298941_rst,I298958,I298975,I298992,I298915,I299023,I299040,I298930,I298912,I299085,I299102,I299119,I299136,I299153,I299170,I299187,I299204,I299221,I298927,I299252,I299269,I299286,I298909,I299317,I298906,I299348,I299365,I299382,I299399,I298921,I299430,I298918,I299461,I299478,I299495,I298924,I298933,I298903,I299587_rst,I299604,I299621,I299638,I299561,I299669,I299686,I299576,I299558,I299731,I299748,I299765,I299782,I299799,I299816,I299833,I299850,I299867,I299573,I299898,I299915,I299932,I299555,I299963,I299552,I299994,I300011,I300028,I300045,I299567,I300076,I299564,I300107,I300124,I300141,I299570,I299579,I299549,I300233_rst,I300250,I300267,I300284,I300207,I300315,I300332,I300222,I300204,I300377,I300394,I300411,I300428,I300445,I300462,I300479,I300496,I300513,I300219,I300544,I300561,I300578,I300201,I300609,I300198,I300640,I300657,I300674,I300691,I300213,I300722,I300210,I300753,I300770,I300787,I300216,I300225,I300195,I300879_rst,I300896,I300913,I300930,I300850,I300961,I300978,I300995,I301012,I301029,I301046,I301063,I301080,I301097,I301114,I300865,I300862,I301159,I300847,I301190,I300844,I301221,I301238,I301255,I301272,I301289,I301306,I300871,I301337,I300859,I300853,I301382,I301399,I300868,I301430,I301447,I301464,I300856,I300841,I301542_rst,I301559,I301576,I301593,I301513,I301624,I301641,I301658,I301675,I301692,I301709,I301726,I301743,I301760,I301777,I301528,I301525,I301822,I301510,I301853,I301507,I301884,I301901,I301918,I301935,I301952,I301969,I301534,I302000,I301522,I301516,I302045,I302062,I301531,I302093,I302110,I302127,I301519,I301504,I302205_rst,I302222,I302239,I302256,I302176,I302287,I302304,I302321,I302338,I302355,I302372,I302389,I302406,I302423,I302440,I302191,I302188,I302485,I302173,I302516,I302170,I302547,I302564,I302581,I302598,I302615,I302632,I302197,I302663,I302185,I302179,I302708,I302725,I302194,I302756,I302773,I302790,I302182,I302167,I302868_rst,I302885,I302902,I302919,I302839,I302950,I302967,I302984,I303001,I303018,I303035,I303052,I303069,I303086,I303103,I302854,I302851,I303148,I302836,I303179,I302833,I303210,I303227,I303244,I303261,I303278,I303295,I302860,I303326,I302848,I302842,I303371,I303388,I302857,I303419,I303436,I303453,I302845,I302830,I303531_rst,I303548,I303565,I303582,I303502,I303613,I303630,I303647,I303664,I303681,I303698,I303715,I303732,I303749,I303766,I303517,I303514,I303811,I303499,I303842,I303496,I303873,I303890,I303907,I303924,I303941,I303958,I303523,I303989,I303511,I303505,I304034,I304051,I303520,I304082,I304099,I304116,I303508,I303493,I304194_rst,I304211,I304228,I304168,I304259,I304276,I304293,I304310,I304327,I304344,I304361,I304378,I304395,I304162,I304426,I304443,I304159,I304474,I304491,I304508,I304171,I304156,I304553,I304570,I304587,I304604,I304621,I304177,I304652,I304186,I304683,I304180,I304183,I304174,I304165,I304789_rst,I304806,I304823,I304854,I304871,I304888,I304905,I304922,I304939,I304956,I304973,I304990,I305021,I305038,I305069,I305086,I305103,I305148,I305165,I305182,I305199,I305216,I305247,I305278,I305384_rst,I305401,I305418,I305449,I305466,I305483,I305500,I305517,I305534,I305551,I305568,I305585,I305616,I305633,I305664,I305681,I305698,I305743,I305760,I305777,I305794,I305811,I305842,I305873,I305979_rst,I305996,I306013,I305953,I306044,I306061,I306078,I306095,I306112,I306129,I306146,I306163,I306180,I305947,I306211,I306228,I305944,I306259,I306276,I306293,I305956,I305941,I306338,I306355,I306372,I306389,I306406,I305962,I306437,I305971,I306468,I305965,I305968,I305959,I305950,I306574_rst,I306591,I306608,I306639,I306656,I306673,I306690,I306707,I306724,I306741,I306758,I306775,I306806,I306823,I306854,I306871,I306888,I306933,I306950,I306967,I306984,I307001,I307032,I307063,I307169_rst,I307186,I307203,I307143,I307234,I307251,I307268,I307285,I307302,I307319,I307336,I307353,I307370,I307137,I307401,I307418,I307134,I307449,I307466,I307483,I307146,I307131,I307528,I307545,I307562,I307579,I307596,I307152,I307627,I307161,I307658,I307155,I307158,I307149,I307140,I307764_rst,I307781,I307826,I307843,I307860,I307877,I307894,I307911,I307928,I307945,I307962,I307993,I308010,I308027,I308044,I308075,I308092,I308109,I308126,I308143,I308174,I308191,I308250,I308281,I308359_rst,I308376,I308342,I308321,I308421,I308438,I308455,I308472,I308489,I308506,I308523,I308540,I308557,I308348,I308588,I308605,I308622,I308639,I308351,I308670,I308687,I308704,I308721,I308738,I308336,I308769,I308786,I308339,I308333,I308327,I308845,I308345,I308876,I308330,I308324,I308954_rst,I308971,I308988,I309005,I309022,I309039,I309056,I309073,I308943,I309104,I308928,I309135,I309152,I309169,I309186,I309203,I309220,I309237,I308925,I309268,I309285,I308922,I309316,I309333,I308940,I309364,I308937,I309395,I309412,I308916,I308919,I309457,I309474,I309491,I309508,I308946,I309539,I308931,I308934,I309617_rst,I309634,I309651,I309668,I309685,I309702,I309719,I309736,I309606,I309767,I309591,I309798,I309815,I309832,I309849,I309866,I309883,I309900,I309588,I309931,I309948,I309585,I309979,I309996,I309603,I310027,I309600,I310058,I310075,I309579,I309582,I310120,I310137,I310154,I310171,I309609,I310202,I309594,I309597,I310280_rst,I310297,I310314,I310331,I310348,I310365,I310382,I310399,I310269,I310430,I310254,I310461,I310478,I310495,I310512,I310529,I310546,I310563,I310251,I310594,I310611,I310248,I310642,I310659,I310266,I310690,I310263,I310721,I310738,I310242,I310245,I310783,I310800,I310817,I310834,I310272,I310865,I310257,I310260,I310943_rst,I310960,I310977,I310994,I311011,I311028,I311045,I311062,I311093,I311124,I311141,I311158,I311175,I311192,I311209,I311226,I311257,I311274,I311305,I311322,I311353,I311384,I311401,I311446,I311463,I311480,I311497,I311528,I311606_rst,I311623,I311640,I311657,I311674,I311691,I311708,I311725,I311595,I311756,I311580,I311787,I311804,I311821,I311838,I311855,I311872,I311889,I311577,I311920,I311937,I311574,I311968,I311985,I311592,I312016,I311589,I312047,I312064,I311568,I311571,I312109,I312126,I312143,I312160,I311598,I312191,I311583,I311586,I312269_rst,I312286,I312303,I312320,I312337,I312354,I312371,I312388,I312258,I312419,I312243,I312450,I312467,I312484,I312501,I312518,I312535,I312552,I312240,I312583,I312600,I312237,I312631,I312648,I312255,I312679,I312252,I312710,I312727,I312231,I312234,I312772,I312789,I312806,I312823,I312261,I312854,I312246,I312249,I312932_rst,I312949,I312966,I312983,I313000,I313017,I313034,I313051,I312921,I313082,I312906,I313113,I313130,I313147,I313164,I313181,I313198,I313215,I312903,I313246,I313263,I312900,I313294,I313311,I312918,I313342,I312915,I313373,I313390,I312894,I312897,I313435,I313452,I313469,I313486,I312924,I313517,I312909,I312912,I313595_rst,I31361_rst2,I313629,I313646,I313663,I313680,I313697,I313714,I313584,I313745,I313569,I313776,I313793,I313810,I313827,I313844,I313861,I313878,I313566,I313909,I313926,I313563,I313957,I313974,I313581,I314005,I313578,I314036,I314053,I313557,I313560,I314098,I314115,I314132,I314149,I313587,I314180,I313572,I313575,I314258_rst,I314275,I314292,I314309,I314326,I314343,I314360,I314377,I314247,I314408,I314232,I314439,I314456,I314473,I314490,I314507,I314524,I314541,I314229,I314572,I314589,I314226,I314620,I314637,I314244,I314668,I314241,I314699,I314716,I314220,I314223,I314761,I314778,I314795,I314812,I314250,I314843,I314235,I314238,I314921_rst,I314938,I314955,I314972,I314989,I315006,I315023,I315040,I314910,I315071,I314895,I315102,I315119,I315136,I315153,I315170,I315187,I315204,I314892,I315235,I315252,I314889,I315283,I315300,I314907,I315331,I314904,I315362,I315379,I314883,I314886,I315424,I315441,I315458,I315475,I314913,I315506,I314898,I314901,I315584_rst,I315601,I315618,I315635,I315652,I315669,I315686,I315703,I315573,I315734,I315558,I315765,I315782,I315799,I315816,I315833,I315850,I315867,I315555,I315898,I315915,I315552,I315946,I315963,I315570,I315994,I315567,I316025,I316042,I315546,I315549,I316087,I316104,I316121,I316138,I315576,I316169,I315561,I315564,I316247_rst,I316264,I316281,I316298,I316315,I316332,I316349,I316218,I316380,I316397,I316414,I316431,I316448,I316465,I316482,I316215,I316513,I316209,I316544,I316561,I316578,I316239,I316212,I316623,I316236,I316654,I316233,I316230,I316699,I316716,I316733,I316750,I316767,I316224,I316798,I316815,I316227,I316221,I316893_rst,I316910,I316927,I316944,I316961,I316978,I316995,I316864,I317026,I317043,I317060,I317077,I317094,I317111,I317128,I316861,I317159,I316855,I317190,I317207,I317224,I316885,I316858,I317269,I316882,I317300,I316879,I316876,I317345,I317362,I317379,I317396,I317413,I316870,I317444,I317461,I316873,I316867,I317539_rst,I317556,I317573,I317590,I317607,I317624,I317641,I317510,I317672,I317689,I317706,I317723,I317740,I317757,I317774,I317507,I317805,I317501,I317836,I317853,I317870,I317531,I317504,I317915,I317528,I317946,I317525,I317522,I317991,I318008,I318025,I318042,I318059,I317516,I318090,I318107,I317519,I317513,I318185_rst,I318202,I318219,I318236,I318253,I318270,I318287,I318156,I318318,I318335,I318352,I318369,I318386,I318403,I318420,I318153,I318451,I318147,I318482,I318499,I318516,I318177,I318150,I318561,I318174,I318592,I318171,I318168,I318637,I318654,I318671,I318688,I318705,I318162,I318736,I318753,I318165,I318159,I318831_rst,I318848,I318865,I318882,I318899,I318916,I318933,I318964,I318981,I318998,I319015,I319032,I319049,I319066,I319097,I319128,I319145,I319162,I319207,I319238,I319283,I319300,I319317,I319334,I319351,I319382,I319399,I319477_rst,I319494,I319511,I319528,I319545,I319562,I319579,I319448,I319610,I319627,I319644,I319661,I319678,I319695,I319712,I319445,I319743,I319439,I319774,I319791,I319808,I319469,I319442,I319853,I319466,I319884,I319463,I319460,I319929,I319946,I319963,I319980,I319997,I319454,I320028,I320045,I319457,I319451,I320123_rst,I320140,I320157,I320174,I320191,I320208,I320225,I320094,I320256,I320273,I320290,I320307,I320324,I320341,I320358,I320091,I320389,I320085,I320420,I320437,I320454,I320115,I320088,I320499,I320112,I320530,I320109,I320106,I320575,I320592,I320609,I320626,I320643,I320100,I320674,I320691,I320103,I320097,I320769_rst,I320786,I320803,I320820,I320837,I320731,I320868,I320885,I320902,I320919,I320936,I320953,I320740,I320984,I320734,I321015,I321032,I321049,I321066,I320761,I320758,I321111,I321128,I321145,I320755,I321176,I320752,I320743,I321221,I321238,I321255,I320746,I320749,I321300,I321317,I320737,I321381_rst,I321398,I321415,I321432,I321449,I321349,I321480,I321497,I321514,I321352,I321545,I321346,I321576,I321593,I321610,I321627,I321644,I321355,I321675,I321692,I321709,I321726,I321361,I321364,I321343,I321785,I321802,I321819,I321373,I321370,I321864,I321881,I321358,I321367,I321959_rst,I321976,I321993,I322010,I322027,I321927,I322058,I322075,I322092,I321930,I322123,I321924,I322154,I322171,I322188,I322205,I322222,I321933,I322253,I322270,I322287,I322304,I321939,I321942,I321921,I322363,I322380,I322397,I321951,I321948,I322442,I322459,I321936,I321945,I322537_rst,I322554,I322571,I322588,I322605,I322505,I322636,I322653,I322670,I322508,I322701,I322502,I322732,I322749,I322766,I322783,I322800,I322511,I322831,I322848,I322865,I322882,I322517,I322520,I322499,I322941,I322958,I322975,I322529,I322526,I323020,I323037,I322514,I322523,I323115_rst,I323132,I323149,I323166,I323183,I323083,I323214,I323231,I323248,I323086,I323279,I323080,I323310,I323327,I323344,I323361,I323378,I323089,I323409,I323426,I323443,I323460,I323095,I323098,I323077,I323519,I323536,I323553,I323107,I323104,I323598,I323615,I323092,I323101,I323693_rst,I323710,I323727,I323744,I323761,I323661,I323792,I323809,I323826,I323664,I323857,I323658,I323888,I323905,I323922,I323939,I323956,I323667,I323987,I324004,I324021,I324038,I323673,I323676,I323655,I324097,I324114,I324131,I323685,I323682,I324176,I324193,I323670,I323679,I324271_rst,I324288,I324305,I324322,I324339,I324239,I324370,I324387,I324404,I324242,I324435,I324236,I324466,I324483,I324500,I324517,I324534,I324245,I324565,I324582,I324599,I324616,I324251,I324254,I324233,I324675,I324692,I324709,I324263,I324260,I324754,I324771,I324248,I324257,I324849_rst,I324866,I324883,I324900,I324917,I324948,I324965,I324982,I325013,I325044,I325061,I325078,I325095,I325112,I325143,I325160,I325177,I325194,I325253,I325270,I325287,I325332,I325349,I325427_rst,I325444,I325461,I325478,I325495,I325526,I325543,I325560,I325591,I325622,I325639,I325656,I325673,I325690,I325721,I325738,I325755,I325772,I325831,I325848,I325865,I325910,I325927,I326005_rst,I326022,I326039,I326056,I326073,I326090,I325988,I326121,I326138,I326155,I325991,I325973,I326200,I326217,I326234,I325994,I325985,I326279,I326296,I326313,I325976,I326344,I326361,I325967,I326392,I326409,I326426,I325997,I326457,I326474,I326491,I326508,I325982,I325979,I325970,I326600_rst,I326617,I326634,I326651,I326668,I326685,I326583,I326716,I326733,I326750,I326586,I326568,I326795,I326812,I326829,I326589,I326580,I326874,I326891,I326908,I326571,I326939,I326956,I326562,I326987,I327004,I327021,I326592,I327052,I327069,I327086,I327103,I326577,I326574,I326565,I327195_rst,I327212,I327229,I327246,I327263,I327280,I327178,I327311,I327328,I327345,I327181,I327163,I327390,I327407,I327424,I327184,I327175,I327469,I327486,I327503,I327166,I327534,I327551,I327157,I327582,I327599,I327616,I327187,I327647,I327664,I327681,I327698,I327172,I327169,I327160,I327790_rst,I327807,I327824,I327841,I327858,I327875,I327773,I327906,I327923,I327940,I327776,I327758,I327985,I328002,I328019,I327779,I327770,I328064,I328081,I328098,I327761,I328129,I328146,I327752,I328177,I328194,I328211,I327782,I328242,I328259,I328276,I328293,I327767,I327764,I327755,I328385_rst,I328402,I328419,I328436,I328453,I328470,I328368,I328501,I328518,I328535,I328371,I328353,I328580,I328597,I328614,I328374,I328365,I328659,I328676,I328693,I328356,I328724,I328741,I328347,I328772,I328789,I328806,I328377,I328837,I328854,I328871,I328888,I328362,I328359,I328350,I328980_rst,I328997,I329014,I329031,I329048,I329065,I328963,I329096,I329113,I329130,I328966,I328948,I329175,I329192,I329209,I328969,I328960,I329254,I329271,I329288,I328951,I329319,I329336,I328942,I329367,I329384,I329401,I328972,I329432,I329449,I329466,I329483,I328957,I328954,I328945,I329575_rst,I329592,I329609,I329626,I329643,I329660,I329558,I329691,I329708,I329725,I329561,I329543,I329770,I329787,I329804,I329564,I329555,I329849,I329866,I329883,I329546,I329914,I329931,I329537,I329962,I329979,I329996,I329567,I330027,I330044,I330061,I330078,I329552,I329549,I329540,I330170_rst,I330187,I330204,I330221,I330238,I330255,I330286,I330303,I330320,I330365,I330382,I330399,I330444,I330461,I330478,I330509,I330526,I330557,I330574,I330591,I330622,I330639,I330656,I330673,I330765_rst,I330782,I330799,I330816,I330833,I330850,I330867,I330736,I330898,I330915,I330932,I330949,I330966,I330983,I331000,I330733,I330727,I331045,I331062,I331079,I330754,I331110,I331127,I330745,I330739,I331172,I330742,I331203,I331220,I330757,I331251,I330751,I330748,I331296,I330730,I331360_rst,I331377,I331394,I331411,I331428,I331445,I331462,I331493,I331510,I331527,I331544,I331561,I331578,I331595,I331640,I331657,I331674,I331705,I331722,I331767,I331798,I331815,I331846,I331891,I331955_rst,I331972,I331989,I332006,I332023,I332040,I332057,I331926,I332088,I332105,I332122,I332139,I332156,I332173,I332190,I331923,I331917,I332235,I332252,I332269,I331944,I332300,I332317,I331935,I331929,I332362,I331932,I332393,I332410,I331947,I332441,I331941,I331938,I33248_rst6,I331920,I332550_rst,I332567,I332584,I332601,I332618,I332635,I332652,I332669,I332686,I332703,I332720,I332737,I332754,I332771,I332539,I332802,I332819,I332836,I332512,I332867,I332533,I332898,I332915,I332518,I332946,I332515,I332521,I332991,I333008,I333025,I332527,I332542,I332530,I333084,I333101,I332536,I332524,I333179_rst,I333196,I333213,I333230,I333247,I333264,I333281,I333298,I333315,I333332,I333349,I333366,I333383,I333400,I333168,I333431,I333448,I333465,I333141,I333496,I333162,I333527,I333544,I333147,I333575,I333144,I333150,I333620,I333637,I333654,I333156,I333171,I333159,I333713,I333730,I333165,I333153,I333808_rst,I333825,I333842,I333859,I333876,I333893,I333910,I333927,I333944,I333961,I333978,I333995,I334012,I334029,I334060,I334077,I334094,I334125,I334156,I334173,I334204,I334249,I334266,I334283,I334342,I334359,I334437_rst,I334454,I334471,I334488,I334505,I334522,I334539,I334556,I334573,I334590,I334607,I334624,I334641,I334658,I334426,I334689,I334706,I334723,I334399,I334754,I334420,I334785,I334802,I334405,I334833,I334402,I334408,I334878,I334895,I334912,I334414,I334429,I334417,I334971,I334988,I334423,I334411,I335066_rst,I335083,I335100,I335117,I335134,I335151,I335168,I335185,I335202,I335219,I335236,I335253,I335270,I335287,I335055,I335318,I335335,I335352,I335028,I335383,I335049,I335414,I335431,I335034,I335462,I335031,I335037,I335507,I335524,I335541,I335043,I335058,I335046,I335600,I335617,I335052,I335040,I335695_rst,I335712,I335729,I335746,I335763,I335780,I335797,I335814,I335831,I335848,I335865,I335882,I335899,I335916,I335684,I335947,I335964,I335981,I335657,I336012,I335678,I336043,I336060,I335663,I336091,I335660,I335666,I336136,I336153,I336170,I335672,I335687,I335675,I336229,I336246,I335681,I335669,I336324_rst,I336341,I336358,I336375,I336392,I336409,I336426,I336443,I336460,I336477,I336494,I336511,I336528,I336545,I336313,I336576,I336593,I336610,I336286,I336641,I336307,I336672,I336689,I336292,I336720,I336289,I336295,I336765,I336782,I336799,I336301,I336316,I336304,I336858,I336875,I336310,I336298,I336953_rst,I336970,I336987,I337004,I337021,I337038,I337055,I337072,I337089,I337106,I337123,I337140,I337157,I337174,I336942,I337205,I337222,I337239,I336915,I337270,I336936,I337301,I337318,I336921,I337349,I336918,I336924,I337394,I337411,I337428,I336930,I336945,I336933,I337487,I337504,I336939,I336927,I337582_rst,I337599,I337616,I337633,I337571,I337664,I337559,I337695,I337712,I337729,I337746,I337763,I337562,I337794,I337547,I337825,I337842,I337859,I337876,I337893,I337910,I337553,I337941,I337958,I337975,I337565,I337574,I337544,I338034,I337568,I337556,I338079,I338096,I337550,I338160_rst,I338177,I338194,I338211,I338149,I338242,I338137,I338273,I338290,I338307,I338324,I338341,I338140,I338372,I338125,I338403,I338420,I338437,I338454,I338471,I338488,I338131,I338519,I338536,I338553,I338143,I338152,I338122,I338612,I338146,I338134,I338657,I338674,I338128,I338738_rst,I338755,I33877_rst2,I338789,I338727,I338820,I338715,I338851,I338868,I338885,I338902,I338919,I338718,I338950,I338703,I338981,I338998,I339015,I339032,I339049,I339066,I338709,I339097,I339114,I339131,I338721,I338730,I338700,I339190,I338724,I338712,I339235,I339252,I338706,I339316_rst,I339333,I339350,I339367,I339384,I339401,I339299,I339287,I339446,I339463,I339480,I339497,I339514,I339296,I339545,I339562,I339579,I339596,I339305,I339284,I339641,I339658,I339302,I339689,I339293,I339308,I339734,I339751,I339768,I339785,I339281,I339290,I339278,I339877_rst,I339894,I339911,I339928,I339945,I339962,I339860,I339848,I340007,I340024,I340041,I340058,I340075,I339857,I340106,I340123,I340140,I340157,I339866,I339845,I340202,I340219,I339863,I340250,I339854,I339869,I340295,I340312,I340329,I340346,I339842,I339851,I339839,I340438_rst,I340455,I340472,I340489,I340506,I340523,I340568,I340585,I340602,I340619,I340636,I340667,I340684,I340701,I340718,I340763,I340780,I340811,I340856,I340873,I340890,I340907,I340999_rst,I341016,I341033,I341050,I341067,I341084,I341129,I341146,I341163,I341180,I341197,I341228,I341245,I341262,I341279,I341324,I341341,I341372,I341417,I341434,I341451,I341468,I341560_rst,I341577,I341594,I341611,I341628,I341645,I341543,I341531,I341690,I341707,I341724,I341741,I341758,I341540,I341789,I341806,I341823,I341840,I341549,I341528,I341885,I341902,I341546,I341933,I341537,I341552,I341978,I341995,I342012,I342029,I341525,I341534,I341522,I342121_rst,I342138,I342155,I342172,I342095,I342203,I342220,I342110,I342092,I342265,I342282,I342299,I342316,I342333,I342350,I342367,I342384,I342401,I342107,I342432,I342449,I342466,I342089,I342497,I342086,I342528,I342545,I342562,I342579,I342101,I342610,I342098,I342641,I342658,I342675,I342104,I342113,I342083,I342767_rst,I342784,I342801,I342818,I342741,I342849,I342866,I342756,I342738,I342911,I342928,I342945,I342962,I342979,I342996,I343013,I343030,I343047,I342753,I343078,I343095,I343112,I342735,I343143,I342732,I343174,I343191,I343208,I343225,I342747,I343256,I342744,I343287,I343304,I343321,I342750,I342759,I342729,I343413_rst,I343430,I343447,I343464,I343387,I343495,I343512,I343402,I343384,I343557,I343574,I343591,I343608,I343625,I343642,I343659,I343676,I343693,I343399,I343724,I343741,I343758,I343381,I343789,I343378,I343820,I343837,I343854,I343871,I343393,I343902,I343390,I343933,I343950,I343967,I343396,I343405,I343375,I344059_rst,I344076,I344093,I344110,I344033,I344141,I344158,I344048,I344030,I344203,I344220,I344237,I344254,I344271,I344288,I344305,I344322,I344339,I344045,I344370,I344387,I344404,I344027,I344435,I344024,I344466,I344483,I344500,I344517,I344039,I344548,I344036,I344579,I344596,I344613,I344042,I344051,I344021,I344705_rst,I344722,I344739,I344756,I344679,I344787,I344804,I344694,I344676,I344849,I344866,I344883,I344900,I344917,I344934,I344951,I344968,I344985,I344691,I345016,I345033,I345050,I344673,I345081,I344670,I345112,I345129,I345146,I345163,I344685,I345194,I344682,I345225,I345242,I345259,I344688,I344697,I344667,I345351_rst,I345368,I345385,I345402,I345325,I345433,I345450,I345340,I345322,I345495,I345512,I345529,I345546,I345563,I345580,I345597,I345614,I345631,I345337,I345662,I345679,I345696,I345319,I345727,I345316,I345758,I345775,I345792,I345809,I345331,I345840,I345328,I345871,I345888,I345905,I345334,I345343,I345313,I345997_rst,I346014,I346031,I346048,I345971,I346079,I346096,I345986,I345968,I346141,I346158,I346175,I346192,I346209,I346226,I346243,I346260,I346277,I345983,I346308,I346325,I346342,I345965,I346373,I345962,I346404,I346421,I346438,I346455,I345977,I346486,I345974,I346517,I346534,I346551,I345980,I345989,I345959,I346643_rst,I346660,I346677,I346694,I346725,I346742,I346787,I346804,I346821,I346838,I346855,I346872,I346889,I346906,I346923,I346954,I346971,I346988,I347019,I347050,I347067,I347084,I347101,I347132,I347163,I347180,I347197,I347289_rst,I347306,I347323,I347340,I347263,I347371,I347388,I347278,I347260,I347433,I347450,I347467,I347484,I347501,I347518,I347535,I347552,I347569,I347275,I347600,I347617,I347634,I347257,I347665,I347254,I347696,I347713,I347730,I347747,I347269,I347778,I347266,I347809,I347826,I347843,I347272,I347281,I347251,I347935_rst,I347952,I347969,I347986,I348017,I348034,I348079,I348096,I348113,I348130,I348147,I348164,I348181,I348198,I348215,I348246,I348263,I348280,I348311,I348342,I348359,I348376,I348393,I348424,I348455,I348472,I348489,I348581_rst,I348598,I348615,I348632,I348555,I348663,I348680,I348570,I348552,I348725,I348742,I348759,I348776,I348793,I348810,I348827,I348844,I348861,I348567,I348892,I348909,I348926,I348549,I348957,I348546,I348988,I349005,I349022,I349039,I348561,I349070,I348558,I349101,I349118,I349135,I348564,I348573,I348543,I349227_rst,I349244,I349261,I349278,I349309,I349326,I349343,I349360,I349377,I349394,I349411,I349428,I349445,I349462,I349507,I349538,I349569,I349586,I349603,I349620,I349637,I349654,I349685,I349730,I349747,I349778,I349795,I349812,I349890_rst,I349907,I349924,I349941,I349861,I349972,I349989,I350006,I350023,I350040,I350057,I350074,I350091,I350108,I350125,I349876,I349873,I350170,I349858,I350201,I349855,I350232,I350249,I350266,I350283,I350300,I350317,I349882,I350348,I349870,I349864,I350393,I350410,I349879,I350441,I350458,I350475,I349867,I349852,I350553_rst,I350570,I350587,I350604,I350635,I350652,I350669,I350686,I350703,I350720,I350737,I350754,I350771,I350788,I350833,I350864,I350895,I350912,I350929,I350946,I350963,I350980,I351011,I351056,I351073,I351104,I351121,I351138,I351216_rst,I351233,I351250,I351190,I351281,I351298,I351315,I351332,I351349,I351366,I351383,I351400,I351417,I351184,I351448,I351465,I351181,I351496,I351513,I351530,I351193,I351178,I351575,I351592,I351609,I351626,I351643,I351199,I351674,I351208,I351705,I351202,I351205,I351196,I351187,I351811_rst,I351828,I351845,I351785,I351876,I351893,I351910,I351927,I351944,I351961,I351978,I351995,I352012,I351779,I352043,I352060,I351776,I352091,I352108,I352125,I351788,I351773,I352170,I352187,I352204,I352221,I352238,I351794,I352269,I351803,I352300,I351797,I351800,I351791,I351782,I352406_rst,I352423,I352440,I352471,I352488,I352505,I352522,I352539,I352556,I352573,I352590,I352607,I352638,I352655,I352686,I352703,I352720,I352765,I352782,I352799,I352816,I352833,I352864,I352895,I353001_rst,I353018,I353035,I353052,I353069,I353086,I353103,I353120,I352990,I353151,I352975,I353182,I353199,I353216,I353233,I353250,I353267,I353284,I352972,I353315,I353332,I352969,I353363,I353380,I352987,I353411,I352984,I353442,I353459,I352963,I352966,I353504,I353521,I353538,I353555,I352993,I353586,I352978,I352981,I353664_rst,I353681,I353698,I353715,I353732,I353749,I353766,I353783,I353814,I353845,I353862,I353879,I353896,I353913,I353930,I353947,I353978,I353995,I354026,I354043,I354074,I354105,I354122,I354167,I354184,I354201,I354218,I354249,I354327_rst,I354344,I354361,I354378,I354395,I354412,I354429,I354446,I354316,I354477,I354301,I354508,I354525,I354542,I354559,I354576,I354593,I354610,I354298,I354641,I354658,I354295,I354689,I354706,I354313,I354737,I354310,I354768,I354785,I354289,I354292,I354830,I354847,I354864,I354881,I354319,I354912,I354304,I354307,I354990_rst,I355007,I355024,I355041,I355058,I355075,I355092,I355109,I355140,I355171,I355188,I355205,I355222,I355239,I355256,I355273,I355304,I355321,I355352,I355369,I355400,I355431,I355448,I355493,I355510,I355527,I355544,I355575,I355653_rst,I355670,I355687,I355704,I355721,I355738,I355755,I355772,I355642,I355803,I355627,I355834,I355851,I355868,I355885,I355902,I355919,I355936,I355624,I355967,I355984,I355621,I356015,I356032,I355639,I356063,I355636,I356094,I35611_rst1,I355615,I355618,I356156,I356173,I356190,I356207,I355645,I356238,I355630,I355633,I356316_rst,I356333,I356350,I356367,I356384,I356401,I356418,I356435,I356466,I356497,I356514,I356531,I356548,I356565,I356582,I356599,I356630,I356647,I356678,I356695,I356726,I356757,I356774,I356819,I356836,I356853,I356870,I356901,I356979_rst,I356996,I357013,I357030,I357047,I357064,I357081,I357098,I356968,I357129,I356953,I357160,I357177,I357194,I357211,I357228,I357245,I357262,I356950,I357293,I357310,I356947,I357341,I357358,I356965,I357389,I356962,I357420,I357437,I356941,I356944,I357482,I357499,I357516,I357533,I356971,I357564,I356956,I356959,I357642_rst,I357659,I357676,I357693,I357710,I357727,I357744,I357761,I357792,I357823,I357840,I357857,I357874,I357891,I357908,I357925,I357956,I357973,I358004,I358021,I358052,I358083,I358100,I358145,I358162,I358179,I358196,I358227,I358305_rst,I358322,I358339,I358356,I358373,I358390,I358407,I358424,I358294,I358455,I358279,I358486,I358503,I358520,I358537,I358554,I358571,I358588,I358276,I358619,I358636,I358273,I358667,I358684,I358291,I358715,I358288,I358746,I358763,I358267,I358270,I358808,I358825,I358842,I358859,I358297,I358890,I358282,I358285,I358968_rst,I358985,I359002,I359019,I359036,I359053,I359070,I359087,I358957,I359118,I358942,I359149,I359166,I359183,I359200,I359217,I359234,I359251,I358939,I359282,I359299,I358936,I359330,I359347,I358954,I359378,I358951,I359409,I359426,I358930,I358933,I359471,I359488,I359505,I359522,I358960,I359553,I358945,I358948,I359631_rst,I359648,I359665,I359682,I359699,I359716,I359733,I359750,I359620,I359781,I359605,I359812,I359829,I359846,I359863,I359880,I359897,I359914,I359602,I359945,I359962,I359599,I359993,I360010,I359617,I360041,I359614,I360072,I360089,I359593,I359596,I360134,I360151,I360168,I360185,I359623,I360216,I359608,I359611,I360294_rst,I360311,I360328,I360345,I360362,I360379,I360396,I360413,I360444,I360475,I360492,I360509,I360526,I360543,I360560,I360577,I360608,I360625,I360656,I360673,I360704,I360735,I360752,I360797,I360814,I360831,I360848,I360879,I360957_rst,I360974,I360991,I361008,I361025,I361042,I361059,I361076,I361107,I361138,I361155,I361172,I361189,I361206,I361223,I361240,I361271,I361288,I361319,I361336,I361367,I361398,I361415,I361460,I361477,I361494,I361511,I361542,I361620_rst,I361637,I361654,I361671,I361688,I361705,I361722,I361591,I361753,I361770,I361787,I361804,I361821,I361838,I361855,I361588,I361886,I361582,I361917,I361934,I361951,I361612,I361585,I361996,I361609,I362027,I361606,I361603,I362072,I362089,I362106,I362123,I362140,I361597,I362171,I362188,I361600,I361594,I362266_rst,I362283,I362300,I362317,I362334,I362351,I362368,I362399,I362416,I362433,I362450,I362467,I362484,I362501,I362532,I362563,I362580,I362597,I362642,I362673,I362718,I362735,I362752,I362769,I362786,I362817,I362834,I362912_rst,I362929,I362946,I362963,I362980,I362997,I363014,I363045,I363062,I363079,I363096,I363113,I363130,I363147,I363178,I363209,I363226,I363243,I363288,I363319,I363364,I363381,I363398,I363415,I363432,I363463,I363480,I363558_rst,I363575,I363592,I363609,I363626,I363643,I363660,I363529,I363691,I363708,I363725,I363742,I363759,I363776,I363793,I363526,I363824,I363520,I363855,I363872,I363889,I363550,I363523,I363934,I363547,I363965,I363544,I363541,I364010,I364027,I364044,I364061,I364078,I363535,I364109,I364126,I363538,I363532,I364204_rst,I364221,I364238,I364255,I364272,I364166,I364303,I364320,I364337,I364354,I364371,I364388,I364175,I364419,I364169,I364450,I364467,I364484,I364501,I364196,I364193,I364546,I364563,I364580,I364190,I364611,I364187,I364178,I364656,I364673,I364690,I364181,I364184,I364735,I364752,I364172,I364816_rst,I364833,I364850,I364867,I364884,I364915,I364932,I364949,I364980,I365011,I365028,I365045,I365062,I365079,I365110,I365127,I365144,I365161,I365220,I365237,I365254,I365299,I365316,I365394_rst,I365411,I365428,I365445,I365462,I365362,I365493,I365510,I365527,I365365,I365558,I365359,I365589,I365606,I365623,I365640,I365657,I365368,I365688,I365705,I365722,I365739,I365374,I365377,I365356,I365798,I365815,I365832,I365386,I365383,I365877,I365894,I365371,I365380,I365972_rst,I365989,I366006,I366023,I366040,I366071,I366088,I366105,I366122,I366139,I366156,I366173,I366190,I366235,I366252,I366283,I366300,I366331,I366348,I366379,I366410,I366441,I366458,I366489,I366520,I366584_rst,I366601,I366618,I366635,I366666,I366683,I366700,I366717,I366734,I366751,I366768,I366799,I366830,I366861,I366878,I366895,I366940,I366957,I366988,I367019,I367036,I367067,I367084,I367162_rst,I367179,I367196,I367213,I367230,I367247,I367278,I367295,I367312,I367357,I367374,I367391,I367436,I367453,I367470,I367501,I367518,I367549,I367566,I367583,I367614,I367631,I367648,I367665,I367757_rst,I367774,I367791,I367808,I367825,I367842,I367740,I367873,I367890,I367907,I367743,I367725,I367952,I367969,I367986,I367746,I367737,I368031,I368048,I368065,I367728,I368096,I368113,I367719,I368144,I368161,I368178,I367749,I368209,I368226,I368243,I368260,I367734,I367731,I367722,I368352_rst,I368369,I368386,I368403,I368420,I368437,I368468,I368485,I368502,I368547,I368564,I368581,I368626,I368643,I368660,I368691,I368708,I368739,I368756,I368773,I368804,I368821,I368838,I368855,I368947_rst,I368964,I368981,I368998,I369015,I369032,I368930,I369063,I369080,I369097,I368933,I368915,I369142,I369159,I369176,I368936,I368927,I369221,I369238,I369255,I368918,I369286,I369303,I368909,I369334,I369351,I369368,I368939,I369399,I369416,I369433,I369450,I368924,I368921,I368912,I369542_rst,I369559,I369576,I369593,I369610,I369627,I369658,I369675,I369692,I369737,I369754,I369771,I369816,I369833,I369850,I369881,I369898,I369929,I369946,I369963,I369994,I370011,I370028,I370045,I370137_rst,I370154,I370171,I370188,I370205,I370222,I370239,I370108,I370270,I370287,I370304,I370321,I370338,I370355,I370372,I370105,I370099,I370417,I370434,I370451,I370126,I370482,I370499,I370117,I370111,I370544,I370114,I370575,I370592,I370129,I370623,I370123,I370120,I370668,I370102,I370732_rst,I370749,I370766,I370783,I370800,I370817,I370834,I370703,I370865,I370882,I370899,I370916,I370933,I370950,I370967,I370700,I370694,I371012,I371029,I371046,I370721,I371077,I371094,I370712,I370706,I371139,I370709,I371170,I371187,I370724,I371218,I370718,I370715,I371263,I370697,I371327_rst,I371344,I371361,I371378,I371395,I371412,I371429,I371446,I371463,I371480,I371497,I371514,I371531,I371548,I371579,I371596,I371613,I371644,I371675,I371692,I371723,I371768,I371785,I371802,I371861,I371878,I371956_rst,I371973,I371990,I372007,I372024,I372041,I372058,I372075,I372092,I372109,I372126,I372143,I372160,I372177,I371945,I372208,I372225,I372242,I371918,I372273,I371939,I372304,I372321,I371924,I372352,I371921,I371927,I372397,I372414,I372431,I371933,I371948,I371936,I372490,I372507,I371942,I371930,I372585_rst,I372602,I372619,I372636,I372653,I372670,I372687,I372704,I372721,I372738,I372755,I372772,I372789,I372806,I372574,I372837,I372854,I372871,I372547,I372902,I372568,I372933,I372950,I372553,I372981,I372550,I372556,I373026,I373043,I373060,I372562,I372577,I372565,I373119,I373136,I372571,I372559,I373214_rst,I373231,I373248,I373265,I373203,I373296,I373191,I373327,I373344,I373361,I373378,I373395,I373194,I373426,I373179,I37345_rst7,I373474,I373491,I373508,I373525,I373542,I373185,I373573,I373590,I373607,I373197,I373206,I373176,I373666,I373200,I373188,I373711,I373728,I373182,I373792_rst,I373809,I373826,I373843,I373874,I373905,I373922,I373939,I373956,I373973,I374004,I374035,I374052,I374069,I374086,I374103,I374120,I374151,I374168,I374185,I374244,I374289,I374306,I374370_rst,I374387,I374404,I374421,I374438,I374455,I374353,I374341,I374500,I374517,I374534,I374551,I374568,I374350,I374599,I374616,I374633,I374650,I374359,I374338,I374695,I374712,I374356,I374743,I374347,I374362,I374788,I374805,I374822,I374839,I374335,I374344,I374332,I374931_rst,I374948,I374965,I374982,I374999,I375016,I375061,I375078,I375095,I375112,I375129,I375160,I375177,I375194,I375211,I375256,I375273,I375304,I375349,I375366,I375383,I375400,I375492_rst,I375509,I375526,I375543,I375560,I375577,I375622,I375639,I375656,I375673,I375690,I375721,I375738,I375755,I375772,I375817,I375834,I375865,I375910,I375927,I375944,I375961,I376053_rst,I376070,I376087,I376104,I376135,I376152,I376197,I376214,I376231,I376248,I376265,I376282,I376299,I376316,I376333,I376364,I376381,I376398,I376429,I376460,I376477,I376494,I376511,I376542,I376573,I376590,I376607,I376699_rst,I376716,I376733,I376750,I376781,I376798,I376815,I376832,I376849,I376866,I376883,I376900,I376917,I376934,I376979,I377010,I377041,I377058,I377075,I377092,I377109,I377126,I377157,I377202,I377219,I377250,I377267,I377284,I377362_rst,I377379,I377396,I377336,I377427,I377444,I377461,I377478,I377495,I377512,I377529,I377546,I377563,I377330,I377594,I377611,I377327,I377642,I377659,I377676,I377339,I377324,I377721,I377738,I377755,I377772,I377789,I377345,I377820,I377354,I377851,I377348,I377351,I377342,I377333,I377957_rst,I377974,I377991,I377931,I378022,I378039,I378056,I378073,I378090,I378107,I378124,I378141,I378158,I377925,I378189,I378206,I377922,I378237,I378254,I378271,I377934,I377919,I378316,I378333,I378350,I378367,I378384,I377940,I378415,I377949,I378446,I377943,I377946,I377937,I377928,I378552_rst,I378569,I378535,I378514,I378614,I378631,I378648,I378665,I378682,I378699,I378716,I378733,I378750,I378541,I378781,I378798,I378815,I378832,I378544,I378863,I378880,I378897,I378914,I378931,I378529,I378962,I378979,I378532,I378526,I378520,I379038,I378538,I37906_rst9,I378523,I378517,I379147_rst,I379164,I379181,I379198,I379215,I379232,I379249,I379266,I379297,I379328,I379345,I379362,I379379,I379396,I379413,I379430,I379461,I379478,I379509,I379526,I379557,I379588,I379605,I379650,I379667,I379684,I379701,I379732,I379810_rst,I379827,I379844,I379861,I379878,I379895,I379912,I379929,I379799,I379960,I379784,I379991,I380008,I380025,I380042,I380059,I380076,I380093,I379781,I380124,I380141,I379778,I380172,I380189,I379796,I380220,I379793,I380251,I380268,I379772,I379775,I380313,I380330,I380347,I380364,I379802,I380395,I379787,I379790,I380473_rst,I380490,I380507,I380524,I380541,I380572,I380589,I380606,I380637,I380668,I380685,I380702,I380719,I380736,I380767,I380784,I380801,I380818,I380877,I380894,I380911,I380956,I380973,I381051_rst,I381068,I381085,I381102,I381119,I381150,I381167,I381184,I381215,I381246,I381263,I381280,I381297,I381314,I381345,I381362,I381379,I381396,I381455,I381472,I381489,I381534,I381551,I381629_rst,I381646,I381663,I381680,I381697,I381728,I381745,I381762,I381793,I381824,I381841,I381858,I381875,I381892,I381923,I381940,I381957,I381974,I382033,I382050,I382067,I382112,I382129,I382207_rst,I382224,I382241,I382258,I382275,I382292,I382323,I382340,I382357,I382402,I382419,I382436,I382481,I382498,I382515,I382546,I382563,I382594,I382611,I382628,I382659,I382676,I382693,I382710,I382802_rst,I382819,I382836,I382853,I382776,I382884,I382901,I382791,I382773,I382946,I382963,I382980,I382997,I383014,I383031,I383048,I383065,I383082,I382788,I383113,I383130,I383147,I382770,I383178,I382767,I383209,I383226,I383243,I383260,I382782,I383291,I382779,I383322,I383339,I383356,I382785,I382794,I382764,I383448_rst,I383465,I383482,I383499,I383530,I383547,I383592,I383609,I383626,I383643,I383660,I383677,I383694,I383711,I383728,I383759,I383776,I383793,I383824,I383855,I383872,I383889,I383906,I383937,I383968,I383985,I384002,I384094_rst,I384111,I384128,I384145,I384162,I384179,I384196,I384213,I384244,I384275,I384292,I384309,I384326,I384343,I384360,I384377,I384408,I384425,I384456,I384473,I384504,I384535,I384552,I384597,I384614,I384631,I384648,I38467_rst9;
not I_0 (I5742_rst,I5701);
nand I_1 (I5759,I1327,I4311);
and I_2 (I5776,I5759,I5543);
DFFARX1 I_3  ( .D(I5776), .CLK(I5694_clk), .RSTB(I5742_rst), .Q(I5793) );
not I_4 (I5810,I5793);
nor I_5 (I5827,I2279,I4311);
or I_6 (I5725,I5827,I5793);
not I_7 (I5713,I5827);
DFFARX1 I_8  ( .D(I2031), .CLK(I5694_clk), .RSTB(I5742_rst), .Q(I5872) );
nor I_9 (I5889,I5872,I5827);
nand I_10 (I5906,I4263,I2583);
and I_11 (I5923,I5906,I4319);
DFFARX1 I_12  ( .D(I5923), .CLK(I5694_clk), .RSTB(I5742_rst), .Q(I5940) );
nor I_13 (I5722,I5940,I5793);
not I_14 (I5971,I5940);
nor I_15 (I5988,I5872,I5971);
DFFARX1 I_16  ( .D(I1639), .CLK(I5694_clk), .RSTB(I5742_rst), .Q(I6005) );
and I_17 (I6022,I6005,I2111);
or I_18 (I5731,I6022,I5827);
nand I_19 (I5710,I6022,I5988);
DFFARX1 I_20  ( .D(I2951), .CLK(I5694_clk), .RSTB(I5742_rst), .Q(I6067) );
and I_21 (I6084,I6067,I5810);
nor I_22 (I5728,I6022,I6084);
nor I_23 (I6115,I6067,I5872);
DFFARX1 I_24  ( .D(I6115), .CLK(I5694_clk), .RSTB(I5742_rst), .Q(I5719) );
nor I_25 (I5734,I6067,I5793);
not I_26 (I6160,I6067);
nor I_27 (I6177,I5940,I6160);
and I_28 (I6194,I5827,I6177);
or I_29 (I6211,I6022,I6194);
DFFARX1 I_30  ( .D(I6211), .CLK(I5694_clk), .RSTB(I5742_rst), .Q(I5707) );
nand I_31 (I5716,I6067,I5889);
nand I_32 (I5704,I6067,I5971);
not I_33 (I6303_rst,I5701);
nand I_34 (I6320,I4759,I3511);
and I_35 (I6337,I6320,I2615);
DFFARX1 I_36  ( .D(I6337), .CLK(I5694_clk), .RSTB(I6303_rst), .Q(I6354) );
not I_37 (I6371,I6354);
nor I_38 (I6388,I4495,I3511);
or I_39 (I6286,I6388,I6354);
not I_40 (I6274,I6388);
DFFARX1 I_41  ( .D(I1695), .CLK(I5694_clk), .RSTB(I6303_rst), .Q(I6433) );
nor I_42 (I6450,I6433,I6388);
nand I_43 (I6467,I2263,I4999);
and I_44 (I6484,I6467,I3319);
DFFARX1 I_45  ( .D(I6484), .CLK(I5694_clk), .RSTB(I6303_rst), .Q(I6501) );
nor I_46 (I6283,I6501,I6354);
not I_47 (I6532,I6501);
nor I_48 (I6549,I6433,I6532);
DFFARX1 I_49  ( .D(I2543), .CLK(I5694_clk), .RSTB(I6303_rst), .Q(I6566) );
and I_50 (I6583,I6566,I2927);
or I_51 (I6292,I6583,I6388);
nand I_52 (I6271,I6583,I6549);
DFFARX1 I_53  ( .D(I3871), .CLK(I5694_clk), .RSTB(I6303_rst), .Q(I6628) );
and I_54 (I6645,I6628,I6371);
nor I_55 (I6289,I6583,I6645);
nor I_56 (I6676,I6628,I6433);
DFFARX1 I_57  ( .D(I6676), .CLK(I5694_clk), .RSTB(I6303_rst), .Q(I6280) );
nor I_58 (I6295,I6628,I6354);
not I_59 (I6721,I6628);
nor I_60 (I6738,I6501,I6721);
and I_61 (I6755,I6388,I6738);
or I_62 (I6772,I6583,I6755);
DFFARX1 I_63  ( .D(I6772), .CLK(I5694_clk), .RSTB(I6303_rst), .Q(I6268) );
nand I_64 (I6277,I6628,I6450);
nand I_65 (I6265,I6628,I6532);
not I_66 (I6864_rst,I5701);
not I_67 (I6881,I3055);
nor I_68 (I6898,I5111,I4271);
nand I_69 (I6915,I6898,I5663);
DFFARX1 I_70  ( .D(I6915), .CLK(I5694_clk), .RSTB(I6864_rst), .Q(I6838) );
nor I_71 (I6946,I6881,I5111);
nand I_72 (I6963,I6946,I5015);
not I_73 (I6853,I6963);
DFFARX1 I_74  ( .D(I6963), .CLK(I5694_clk), .RSTB(I6864_rst), .Q(I6835) );
not I_75 (I7008,I5111);
not I_76 (I7025,I7008);
not I_77 (I7042,I4223);
nor I_78 (I7059,I7042,I1615);
and I_79 (I7076,I7059,I4279);
or I_80 (I7093,I7076,I5471);
DFFARX1 I_81  ( .D(I7093), .CLK(I5694_clk), .RSTB(I6864_rst), .Q(I7110) );
nor I_82 (I7127,I7110,I6963);
nor I_83 (I7144,I7110,I7025);
nand I_84 (I6850,I6915,I7144);
nand I_85 (I7175,I6881,I4223);
nand I_86 (I7192,I7175,I7110);
and I_87 (I7209,I7175,I7192);
DFFARX1 I_88  ( .D(I7209), .CLK(I5694_clk), .RSTB(I6864_rst), .Q(I6832) );
DFFARX1 I_89  ( .D(I7175), .CLK(I5694_clk), .RSTB(I6864_rst), .Q(I7240) );
and I_90 (I6829,I7008,I7240);
DFFARX1 I_91  ( .D(I3031), .CLK(I5694_clk), .RSTB(I6864_rst), .Q(I7271) );
not I_92 (I7288,I7271);
nor I_93 (I7305,I6963,I7288);
and I_94 (I7322,I7271,I7305);
nand I_95 (I6844,I7271,I7025);
DFFARX1 I_96  ( .D(I7271), .CLK(I5694_clk), .RSTB(I6864_rst), .Q(I7353) );
not I_97 (I6841,I7353);
DFFARX1 I_98  ( .D(I3735), .CLK(I5694_clk), .RSTB(I6864_rst), .Q(I7384) );
not I_99 (I7401,I7384);
or I_100 (I7418,I7401,I7322);
DFFARX1 I_101  ( .D(I7418), .CLK(I5694_clk), .RSTB(I6864_rst), .Q(I6847) );
nand I_102 (I6856,I7401,I7127);
DFFARX1 I_103  ( .D(I7401), .CLK(I5694_clk), .RSTB(I6864_rst), .Q(I6826) );
not I_104 (I7510_rst,I5701);
not I_105 (I7527,I5431);
nor I_106 (I7544,I1463,I3927);
nand I_107 (I7561,I7544,I1687);
DFFARX1 I_108  ( .D(I7561), .CLK(I5694_clk), .RSTB(I7510_rst), .Q(I7481) );
nor I_109 (I7592,I7527,I1463);
nand I_110 (I7609,I7592,I5551);
nand I_111 (I7626,I7609,I7561);
not I_112 (I7643,I1463);
not I_113 (I7660,I1727);
nor I_114 (I7677,I7660,I5335);
and I_115 (I7694,I7677,I3951);
or I_116 (I7711,I7694,I3791);
DFFARX1 I_117  ( .D(I7711), .CLK(I5694_clk), .RSTB(I7510_rst), .Q(I7728) );
nor I_118 (I7745,I7728,I7609);
nand I_119 (I7496,I7643,I7745);
not I_120 (I7493,I7728);
and I_121 (I7790,I7728,I7626);
DFFARX1 I_122  ( .D(I7790), .CLK(I5694_clk), .RSTB(I7510_rst), .Q(I7478) );
DFFARX1 I_123  ( .D(I7728), .CLK(I5694_clk), .RSTB(I7510_rst), .Q(I7821) );
and I_124 (I7475,I7643,I7821);
nand I_125 (I7852,I7527,I1727);
not I_126 (I7869,I7852);
nor I_127 (I7886,I7728,I7869);
DFFARX1 I_128  ( .D(I1967), .CLK(I5694_clk), .RSTB(I7510_rst), .Q(I7903) );
nand I_129 (I7920,I7903,I7852);
and I_130 (I7937,I7643,I7920);
DFFARX1 I_131  ( .D(I7937), .CLK(I5694_clk), .RSTB(I7510_rst), .Q(I7502) );
not I_132 (I7968,I7903);
nand I_133 (I7490,I7903,I7886);
nand I_134 (I7484,I7903,I7869);
DFFARX1 I_135  ( .D(I4367), .CLK(I5694_clk), .RSTB(I7510_rst), .Q(I8013) );
not I_136 (I8030,I8013);
nor I_137 (I7499,I7903,I8030);
nor I_138 (I8061,I8030,I7968);
and I_139 (I8078,I7609,I8061);
or I_140 (I8095,I7852,I8078);
DFFARX1 I_141  ( .D(I8095), .CLK(I5694_clk), .RSTB(I7510_rst), .Q(I7487) );
DFFARX1 I_142  ( .D(I8030), .CLK(I5694_clk), .RSTB(I7510_rst), .Q(I7472) );
not I_143 (I8173_rst,I5701);
not I_144 (I8190,I1263);
nor I_145 (I8207,I4679,I2791);
nand I_146 (I8224,I8207,I2967);
DFFARX1 I_147  ( .D(I8224), .CLK(I5694_clk), .RSTB(I8173_rst), .Q(I8144) );
nor I_148 (I8255,I8190,I4679);
nand I_149 (I8272,I8255,I4447);
nand I_150 (I8289,I8272,I8224);
not I_151 (I8306,I4679);
not I_152 (I8323,I5583);
nor I_153 (I8340,I8323,I3287);
and I_154 (I8357,I8340,I5527);
or I_155 (I8374,I8357,I4519);
DFFARX1 I_156  ( .D(I8374), .CLK(I5694_clk), .RSTB(I8173_rst), .Q(I8391) );
nor I_157 (I8408,I8391,I8272);
nand I_158 (I8159,I8306,I8408);
not I_159 (I8156,I8391);
and I_160 (I8453,I8391,I8289);
DFFARX1 I_161  ( .D(I8453), .CLK(I5694_clk), .RSTB(I8173_rst), .Q(I8141) );
DFFARX1 I_162  ( .D(I8391), .CLK(I5694_clk), .RSTB(I8173_rst), .Q(I8484) );
and I_163 (I8138,I8306,I8484);
nand I_164 (I8515,I8190,I5583);
not I_165 (I8532,I8515);
nor I_166 (I8549,I8391,I8532);
DFFARX1 I_167  ( .D(I2231), .CLK(I5694_clk), .RSTB(I8173_rst), .Q(I8566) );
nand I_168 (I8583,I8566,I8515);
and I_169 (I8600,I8306,I8583);
DFFARX1 I_170  ( .D(I8600), .CLK(I5694_clk), .RSTB(I8173_rst), .Q(I8165) );
not I_171 (I8631,I8566);
nand I_172 (I8153,I8566,I8549);
nand I_173 (I8147,I8566,I8532);
DFFARX1 I_174  ( .D(I5047), .CLK(I5694_clk), .RSTB(I8173_rst), .Q(I8676) );
not I_175 (I8693,I8676);
nor I_176 (I8162,I8566,I8693);
nor I_177 (I8724,I8693,I8631);
and I_178 (I8741,I8272,I8724);
or I_179 (I8758,I8515,I8741);
DFFARX1 I_180  ( .D(I8758), .CLK(I5694_clk), .RSTB(I8173_rst), .Q(I8150) );
DFFARX1 I_181  ( .D(I8693), .CLK(I5694_clk), .RSTB(I8173_rst), .Q(I8135) );
not I_182 (I8836_rst,I5701);
not I_183 (I8853,I3279);
nor I_184 (I8870,I3983,I1311);
nand I_185 (I8887,I8870,I5311);
DFFARX1 I_186  ( .D(I8887), .CLK(I5694_clk), .RSTB(I8836_rst), .Q(I8807) );
nor I_187 (I8918,I8853,I3983);
nand I_188 (I8935,I8918,I5103);
nand I_189 (I8952,I8935,I8887);
not I_190 (I8969,I3983);
not I_191 (I8986,I1927);
nor I_192 (I9003,I8986,I1943);
and I_193 (I9020,I9003,I3991);
or I_194 (I9037,I9020,I3719);
DFFARX1 I_195  ( .D(I9037), .CLK(I5694_clk), .RSTB(I8836_rst), .Q(I9054) );
nor I_196 (I9071,I9054,I8935);
nand I_197 (I8822,I8969,I9071);
not I_198 (I8819,I9054);
and I_199 (I9116,I9054,I8952);
DFFARX1 I_200  ( .D(I9116), .CLK(I5694_clk), .RSTB(I8836_rst), .Q(I8804) );
DFFARX1 I_201  ( .D(I9054), .CLK(I5694_clk), .RSTB(I8836_rst), .Q(I9147) );
and I_202 (I8801,I8969,I9147);
nand I_203 (I9178,I8853,I1927);
not I_204 (I9195,I9178);
nor I_205 (I9212,I9054,I9195);
DFFARX1 I_206  ( .D(I2511), .CLK(I5694_clk), .RSTB(I8836_rst), .Q(I9229) );
nand I_207 (I9246,I9229,I9178);
and I_208 (I9263,I8969,I9246);
DFFARX1 I_209  ( .D(I9263), .CLK(I5694_clk), .RSTB(I8836_rst), .Q(I8828) );
not I_210 (I9294,I9229);
nand I_211 (I8816,I9229,I9212);
nand I_212 (I8810,I9229,I9195);
DFFARX1 I_213  ( .D(I4983), .CLK(I5694_clk), .RSTB(I8836_rst), .Q(I9339) );
not I_214 (I9356,I9339);
nor I_215 (I8825,I9229,I9356);
nor I_216 (I9387,I9356,I9294);
and I_217 (I9404,I8935,I9387);
or I_218 (I9421,I9178,I9404);
DFFARX1 I_219  ( .D(I9421), .CLK(I5694_clk), .RSTB(I8836_rst), .Q(I8813) );
DFFARX1 I_220  ( .D(I9356), .CLK(I5694_clk), .RSTB(I8836_rst), .Q(I8798) );
not I_221 (I9499_rst,I5701);
not I_222 (I9516,I3039);
nor I_223 (I9533,I4927,I1471);
nand I_224 (I9550,I9533,I1647);
DFFARX1 I_225  ( .D(I9550), .CLK(I5694_clk), .RSTB(I9499_rst), .Q(I9470) );
nor I_226 (I9581,I9516,I4927);
nand I_227 (I9598,I9581,I3207);
nand I_228 (I9615,I9598,I9550);
not I_229 (I9632,I4927);
not I_230 (I9649,I3151);
nor I_231 (I9666,I9649,I5055);
and I_232 (I9683,I9666,I1655);
or I_233 (I9700,I9683,I2207);
DFFARX1 I_234  ( .D(I9700), .CLK(I5694_clk), .RSTB(I9499_rst), .Q(I9717) );
nor I_235 (I9734,I9717,I9598);
nand I_236 (I9485,I9632,I9734);
not I_237 (I9482,I9717);
and I_238 (I9779,I9717,I9615);
DFFARX1 I_239  ( .D(I9779), .CLK(I5694_clk), .RSTB(I9499_rst), .Q(I9467) );
DFFARX1 I_240  ( .D(I9717), .CLK(I5694_clk), .RSTB(I9499_rst), .Q(I9810) );
and I_241 (I9464,I9632,I9810);
nand I_242 (I9841,I9516,I3151);
not I_243 (I9858,I9841);
nor I_244 (I9875,I9717,I9858);
DFFARX1 I_245  ( .D(I5399), .CLK(I5694_clk), .RSTB(I9499_rst), .Q(I9892) );
nand I_246 (I9909,I9892,I9841);
and I_247 (I9926,I9632,I9909);
DFFARX1 I_248  ( .D(I9926), .CLK(I5694_clk), .RSTB(I9499_rst), .Q(I9491) );
not I_249 (I9957,I9892);
nand I_250 (I9479,I9892,I9875);
nand I_251 (I9473,I9892,I9858);
DFFARX1 I_252  ( .D(I2567), .CLK(I5694_clk), .RSTB(I9499_rst), .Q(I10002) );
not I_253 (I10019,I10002);
nor I_254 (I9488,I9892,I10019);
nor I_255 (I10050,I10019,I9957);
and I_256 (I10067,I9598,I10050);
or I_257 (I10084,I9841,I10067);
DFFARX1 I_258  ( .D(I10084), .CLK(I5694_clk), .RSTB(I9499_rst), .Q(I9476) );
DFFARX1 I_259  ( .D(I10019), .CLK(I5694_clk), .RSTB(I9499_rst), .Q(I9461) );
not I_260 (I10162_rst,I5701);
not I_261 (I10179,I4695);
nor I_262 (I10196,I2319,I5631);
nand I_263 (I10213,I10196,I3751);
DFFARX1 I_264  ( .D(I10213), .CLK(I5694_clk), .RSTB(I10162_rst), .Q(I10133) );
nor I_265 (I10244,I10179,I2319);
nand I_266 (I10261,I10244,I2327);
nand I_267 (I10278,I10261,I10213);
not I_268 (I10295,I2319);
not I_269 (I10312,I1575);
nor I_270 (I10329,I10312,I2295);
and I_271 (I10346,I10329,I4631);
or I_272 (I10363,I10346,I4919);
DFFARX1 I_273  ( .D(I10363), .CLK(I5694_clk), .RSTB(I10162_rst), .Q(I10380) );
nor I_274 (I10397,I10380,I10261);
nand I_275 (I10148,I10295,I10397);
not I_276 (I10145,I10380);
and I_277 (I10442,I10380,I10278);
DFFARX1 I_278  ( .D(I10442), .CLK(I5694_clk), .RSTB(I10162_rst), .Q(I10130) );
DFFARX1 I_279  ( .D(I10380), .CLK(I5694_clk), .RSTB(I10162_rst), .Q(I10473) );
and I_280 (I10127,I10295,I10473);
nand I_281 (I10504,I10179,I1575);
not I_282 (I10521,I10504);
nor I_283 (I10538,I10380,I10521);
DFFARX1 I_284  ( .D(I1847), .CLK(I5694_clk), .RSTB(I10162_rst), .Q(I10555) );
nand I_285 (I10572,I10555,I10504);
and I_286 (I10589,I10295,I10572);
DFFARX1 I_287  ( .D(I10589), .CLK(I5694_clk), .RSTB(I10162_rst), .Q(I10154) );
not I_288 (I10620,I10555);
nand I_289 (I10142,I10555,I10538);
nand I_290 (I10136,I10555,I10521);
DFFARX1 I_291  ( .D(I2655), .CLK(I5694_clk), .RSTB(I10162_rst), .Q(I10665) );
not I_292 (I10682,I10665);
nor I_293 (I10151,I10555,I10682);
nor I_294 (I10713,I10682,I10620);
and I_295 (I10730,I10261,I10713);
or I_296 (I10747,I10504,I10730);
DFFARX1 I_297  ( .D(I10747), .CLK(I5694_clk), .RSTB(I10162_rst), .Q(I10139) );
DFFARX1 I_298  ( .D(I10682), .CLK(I5694_clk), .RSTB(I10162_rst), .Q(I10124) );
not I_299 (I10825_rst,I5701);
not I_300 (I10842,I4295);
nor I_301 (I10859,I4527,I1287);
nand I_302 (I10876,I10859,I5127);
DFFARX1 I_303  ( .D(I10876), .CLK(I5694_clk), .RSTB(I10825_rst), .Q(I10796) );
nor I_304 (I10907,I10842,I4527);
nand I_305 (I10924,I10907,I3743);
nand I_306 (I10941,I10924,I10876);
not I_307 (I10958,I4527);
not I_308 (I10975,I3007);
nor I_309 (I10992,I10975,I2831);
and I_310 (I11009,I10992,I5607);
or I_311 (I11026,I11009,I4663);
DFFARX1 I_312  ( .D(I11026), .CLK(I5694_clk), .RSTB(I10825_rst), .Q(I11043) );
nor I_313 (I11060,I11043,I10924);
nand I_314 (I10811,I10958,I11060);
not I_315 (I10808,I11043);
and I_316 (I11105,I11043,I10941);
DFFARX1 I_317  ( .D(I11105), .CLK(I5694_clk), .RSTB(I10825_rst), .Q(I10793) );
DFFARX1 I_318  ( .D(I11043), .CLK(I5694_clk), .RSTB(I10825_rst), .Q(I11136) );
and I_319 (I10790,I10958,I11136);
nand I_320 (I11167,I10842,I3007);
not I_321 (I11184,I11167);
nor I_322 (I11201,I11043,I11184);
DFFARX1 I_323  ( .D(I2023), .CLK(I5694_clk), .RSTB(I10825_rst), .Q(I11218) );
nand I_324 (I11235,I11218,I11167);
and I_325 (I11252,I10958,I11235);
DFFARX1 I_326  ( .D(I11252), .CLK(I5694_clk), .RSTB(I10825_rst), .Q(I10817) );
not I_327 (I11283,I11218);
nand I_328 (I10805,I11218,I11201);
nand I_329 (I10799,I11218,I11184);
DFFARX1 I_330  ( .D(I4903), .CLK(I5694_clk), .RSTB(I10825_rst), .Q(I11328) );
not I_331 (I11345,I11328);
nor I_332 (I10814,I11218,I11345);
nor I_333 (I11376,I11345,I11283);
and I_334 (I11393,I10924,I11376);
or I_335 (I11410,I11167,I11393);
DFFARX1 I_336  ( .D(I11410), .CLK(I5694_clk), .RSTB(I10825_rst), .Q(I10802) );
DFFARX1 I_337  ( .D(I11345), .CLK(I5694_clk), .RSTB(I10825_rst), .Q(I10787) );
not I_338 (I11488_rst,I5701);
or I_339 (I11505,I3895,I4079);
or I_340 (I11522,I3919,I3895);
DFFARX1 I_341  ( .D(I11522), .CLK(I5694_clk), .RSTB(I11488_rst), .Q(I11462) );
nor I_342 (I11553,I4791,I1503);
not I_343 (I11570,I11553);
not I_344 (I11587,I4791);
and I_345 (I11604,I11587,I3639);
nor I_346 (I11621,I11604,I4079);
nor I_347 (I11638,I5383,I4511);
DFFARX1 I_348  ( .D(I11638), .CLK(I5694_clk), .RSTB(I11488_rst), .Q(I11655) );
nand I_349 (I11672,I11655,I11505);
and I_350 (I11689,I11621,I11672);
DFFARX1 I_351  ( .D(I11689), .CLK(I5694_clk), .RSTB(I11488_rst), .Q(I11456) );
nor I_352 (I11720,I5383,I3919);
DFFARX1 I_353  ( .D(I11720), .CLK(I5694_clk), .RSTB(I11488_rst), .Q(I11737) );
and I_354 (I11453,I11553,I11737);
DFFARX1 I_355  ( .D(I4479), .CLK(I5694_clk), .RSTB(I11488_rst), .Q(I11768) );
and I_356 (I11785,I11768,I4055);
DFFARX1 I_357  ( .D(I11785), .CLK(I5694_clk), .RSTB(I11488_rst), .Q(I11802) );
not I_358 (I11465,I11802);
DFFARX1 I_359  ( .D(I11785), .CLK(I5694_clk), .RSTB(I11488_rst), .Q(I11450) );
DFFARX1 I_360  ( .D(I2879), .CLK(I5694_clk), .RSTB(I11488_rst), .Q(I11847) );
not I_361 (I11864,I11847);
nor I_362 (I11881,I11522,I11864);
and I_363 (I11898,I11785,I11881);
or I_364 (I11915,I11505,I11898);
DFFARX1 I_365  ( .D(I11915), .CLK(I5694_clk), .RSTB(I11488_rst), .Q(I11471) );
nor I_366 (I11946,I11847,I11655);
nand I_367 (I11480,I11621,I11946);
nor I_368 (I11977,I11847,I11570);
nand I_369 (I11474,I11720,I11977);
not I_370 (I11477,I11847);
nand I_371 (I11468,I11847,I11570);
DFFARX1 I_372  ( .D(I11847), .CLK(I5694_clk), .RSTB(I11488_rst), .Q(I11459) );
not I_373 (I12083_rst,I5701);
or I_374 (I12100,I3535,I1975);
or I_375 (I12117,I3375,I3535);
DFFARX1 I_376  ( .D(I12117), .CLK(I5694_clk), .RSTB(I12083_rst), .Q(I12057) );
nor I_377 (I12148,I2671,I4871);
not I_378 (I12165,I12148);
not I_379 (I12182,I2671);
and I_380 (I12199,I12182,I5655);
nor I_381 (I12216,I12199,I1975);
nor I_382 (I12233,I2455,I4831);
DFFARX1 I_383  ( .D(I12233), .CLK(I5694_clk), .RSTB(I12083_rst), .Q(I12250) );
nand I_384 (I12267,I12250,I12100);
and I_385 (I12284,I12216,I12267);
DFFARX1 I_386  ( .D(I12284), .CLK(I5694_clk), .RSTB(I12083_rst), .Q(I12051) );
nor I_387 (I12315,I2455,I3375);
DFFARX1 I_388  ( .D(I12315), .CLK(I5694_clk), .RSTB(I12083_rst), .Q(I12332) );
and I_389 (I12048,I12148,I12332);
DFFARX1 I_390  ( .D(I5575), .CLK(I5694_clk), .RSTB(I12083_rst), .Q(I12363) );
and I_391 (I12380,I12363,I3351);
DFFARX1 I_392  ( .D(I12380), .CLK(I5694_clk), .RSTB(I12083_rst), .Q(I12397) );
not I_393 (I12060,I12397);
DFFARX1 I_394  ( .D(I12380), .CLK(I5694_clk), .RSTB(I12083_rst), .Q(I12045) );
DFFARX1 I_395  ( .D(I4287), .CLK(I5694_clk), .RSTB(I12083_rst), .Q(I12442) );
not I_396 (I12459,I12442);
nor I_397 (I12476,I12117,I12459);
and I_398 (I12493,I12380,I12476);
or I_399 (I12510,I12100,I12493);
DFFARX1 I_400  ( .D(I12510), .CLK(I5694_clk), .RSTB(I12083_rst), .Q(I12066) );
nor I_401 (I12541,I12442,I12250);
nand I_402 (I12075,I12216,I12541);
nor I_403 (I12572,I12442,I12165);
nand I_404 (I12069,I12315,I12572);
not I_405 (I12072,I12442);
nand I_406 (I12063,I12442,I12165);
DFFARX1 I_407  ( .D(I12442), .CLK(I5694_clk), .RSTB(I12083_rst), .Q(I12054) );
not I_408 (I12678_rst,I5701);
not I_409 (I12695,I2799);
nor I_410 (I12712,I4031,I3431);
nand I_411 (I12729,I12712,I5039);
nor I_412 (I12746,I12695,I4031);
nand I_413 (I12763,I12746,I1439);
not I_414 (I12780,I12763);
not I_415 (I12797,I4031);
nor I_416 (I12667,I12763,I12797);
not I_417 (I12828,I12797);
nand I_418 (I12652,I12763,I12828);
not I_419 (I12859,I1447);
nor I_420 (I12876,I12859,I2175);
and I_421 (I12893,I12876,I1527);
or I_422 (I12910,I12893,I4503);
DFFARX1 I_423  ( .D(I12910), .CLK(I5694_clk), .RSTB(I12678_rst), .Q(I12927) );
nor I_424 (I12944,I12927,I12780);
DFFARX1 I_425  ( .D(I12927), .CLK(I5694_clk), .RSTB(I12678_rst), .Q(I12961) );
not I_426 (I12649,I12961);
nand I_427 (I12992,I12695,I1447);
and I_428 (I13009,I12992,I12944);
DFFARX1 I_429  ( .D(I12992), .CLK(I5694_clk), .RSTB(I12678_rst), .Q(I12646) );
DFFARX1 I_430  ( .D(I2447), .CLK(I5694_clk), .RSTB(I12678_rst), .Q(I13040) );
nor I_431 (I13057,I13040,I12763);
nand I_432 (I12664,I12927,I13057);
nor I_433 (I13088,I13040,I12828);
not I_434 (I12661,I13040);
nand I_435 (I13119,I13040,I12729);
and I_436 (I13136,I12797,I13119);
DFFARX1 I_437  ( .D(I13136), .CLK(I5694_clk), .RSTB(I12678_rst), .Q(I12640) );
DFFARX1 I_438  ( .D(I13040), .CLK(I5694_clk), .RSTB(I12678_rst), .Q(I12643) );
DFFARX1 I_439  ( .D(I3695), .CLK(I5694_clk), .RSTB(I12678_rst), .Q(I13181) );
not I_440 (I13198,I13181);
nand I_441 (I13215,I13198,I12763);
and I_442 (I13232,I12992,I13215);
DFFARX1 I_443  ( .D(I13232), .CLK(I5694_clk), .RSTB(I12678_rst), .Q(I12670) );
or I_444 (I13263,I13198,I13009);
DFFARX1 I_445  ( .D(I13263), .CLK(I5694_clk), .RSTB(I12678_rst), .Q(I12655) );
nand I_446 (I12658,I13198,I13088);
not I_447 (I13341_rst,I5701);
not I_448 (I13358,I1431);
nor I_449 (I13375,I2591,I2807);
nand I_450 (I13392,I13375,I2127);
nor I_451 (I13409,I13358,I2591);
nand I_452 (I13426,I13409,I4087);
not I_453 (I13443,I13426);
not I_454 (I13460,I2591);
nor I_455 (I13330,I13426,I13460);
not I_456 (I13491,I13460);
nand I_457 (I13315,I13426,I13491);
not I_458 (I13522,I4151);
nor I_459 (I13539,I13522,I5559);
and I_460 (I13556,I13539,I4255);
or I_461 (I13573,I13556,I4639);
DFFARX1 I_462  ( .D(I13573), .CLK(I5694_clk), .RSTB(I13341_rst), .Q(I13590) );
nor I_463 (I13607,I13590,I13443);
DFFARX1 I_464  ( .D(I13590), .CLK(I5694_clk), .RSTB(I13341_rst), .Q(I13624) );
not I_465 (I13312,I13624);
nand I_466 (I13655,I13358,I4151);
and I_467 (I13672,I13655,I13607);
DFFARX1 I_468  ( .D(I13655), .CLK(I5694_clk), .RSTB(I13341_rst), .Q(I13309) );
DFFARX1 I_469  ( .D(I1599), .CLK(I5694_clk), .RSTB(I13341_rst), .Q(I13703) );
nor I_470 (I13720,I13703,I13426);
nand I_471 (I13327,I13590,I13720);
nor I_472 (I13751,I13703,I13491);
not I_473 (I13324,I13703);
nand I_474 (I13782,I13703,I13392);
and I_475 (I13799,I13460,I13782);
DFFARX1 I_476  ( .D(I13799), .CLK(I5694_clk), .RSTB(I13341_rst), .Q(I13303) );
DFFARX1 I_477  ( .D(I13703), .CLK(I5694_clk), .RSTB(I13341_rst), .Q(I13306) );
DFFARX1 I_478  ( .D(I2423), .CLK(I5694_clk), .RSTB(I13341_rst), .Q(I13844) );
not I_479 (I13861,I13844);
nand I_480 (I13878,I13861,I13426);
and I_481 (I13895,I13655,I13878);
DFFARX1 I_482  ( .D(I13895), .CLK(I5694_clk), .RSTB(I13341_rst), .Q(I13333) );
or I_483 (I13926,I13861,I13672);
DFFARX1 I_484  ( .D(I13926), .CLK(I5694_clk), .RSTB(I13341_rst), .Q(I13318) );
nand I_485 (I13321,I13861,I13751);
not I_486 (I14004_rst,I5701);
not I_487 (I14021,I5263);
nor I_488 (I14038,I3191,I5175);
nand I_489 (I14055,I14038,I3399);
nor I_490 (I14072,I14021,I3191);
nand I_491 (I14089,I14072,I3799);
not I_492 (I14106,I14089);
not I_493 (I14123,I3191);
nor I_494 (I13993,I14089,I14123);
not I_495 (I14154,I14123);
nand I_496 (I13978,I14089,I14154);
not I_497 (I14185,I1887);
nor I_498 (I14202,I14185,I1791);
and I_499 (I14219,I14202,I3343);
or I_500 (I14236,I14219,I1607);
DFFARX1 I_501  ( .D(I14236), .CLK(I5694_clk), .RSTB(I14004_rst), .Q(I14253) );
nor I_502 (I14270,I14253,I14106);
DFFARX1 I_503  ( .D(I14253), .CLK(I5694_clk), .RSTB(I14004_rst), .Q(I14287) );
not I_504 (I13975,I14287);
nand I_505 (I14318,I14021,I1887);
and I_506 (I14335,I14318,I14270);
DFFARX1 I_507  ( .D(I14318), .CLK(I5694_clk), .RSTB(I14004_rst), .Q(I13972) );
DFFARX1 I_508  ( .D(I5503), .CLK(I5694_clk), .RSTB(I14004_rst), .Q(I14366) );
nor I_509 (I14383,I14366,I14089);
nand I_510 (I13990,I14253,I14383);
nor I_511 (I14414,I14366,I14154);
not I_512 (I13987,I14366);
nand I_513 (I14445,I14366,I14055);
and I_514 (I14462,I14123,I14445);
DFFARX1 I_515  ( .D(I14462), .CLK(I5694_clk), .RSTB(I14004_rst), .Q(I13966) );
DFFARX1 I_516  ( .D(I14366), .CLK(I5694_clk), .RSTB(I14004_rst), .Q(I13969) );
DFFARX1 I_517  ( .D(I4583), .CLK(I5694_clk), .RSTB(I14004_rst), .Q(I14507) );
not I_518 (I14524,I14507);
nand I_519 (I14541,I14524,I14089);
and I_520 (I14558,I14318,I14541);
DFFARX1 I_521  ( .D(I14558), .CLK(I5694_clk), .RSTB(I14004_rst), .Q(I13996) );
or I_522 (I14589,I14524,I14335);
DFFARX1 I_523  ( .D(I14589), .CLK(I5694_clk), .RSTB(I14004_rst), .Q(I13981) );
nand I_524 (I13984,I14524,I14414);
not I_525 (I14667_rst,I5701);
not I_526 (I14684,I5567);
nor I_527 (I14701,I5447,I5351);
nand I_528 (I14718,I14701,I5079);
nor I_529 (I14735,I14684,I5447);
nand I_530 (I14752,I14735,I4471);
not I_531 (I14769,I14752);
not I_532 (I14786,I5447);
nor I_533 (I14656,I14752,I14786);
not I_534 (I14817,I14786);
nand I_535 (I14641,I14752,I14817);
not I_536 (I14848,I1255);
nor I_537 (I14865,I14848,I4111);
and I_538 (I14882,I14865,I3615);
or I_539 (I14899,I14882,I5319);
DFFARX1 I_540  ( .D(I14899), .CLK(I5694_clk), .RSTB(I14667_rst), .Q(I14916) );
nor I_541 (I14933,I14916,I14769);
DFFARX1 I_542  ( .D(I14916), .CLK(I5694_clk), .RSTB(I14667_rst), .Q(I14950) );
not I_543 (I14638,I14950);
nand I_544 (I14981,I14684,I1255);
and I_545 (I14998,I14981,I14933);
DFFARX1 I_546  ( .D(I14981), .CLK(I5694_clk), .RSTB(I14667_rst), .Q(I14635) );
DFFARX1 I_547  ( .D(I4951), .CLK(I5694_clk), .RSTB(I14667_rst), .Q(I15029) );
nor I_548 (I15046,I15029,I14752);
nand I_549 (I14653,I14916,I15046);
nor I_550 (I15077,I15029,I14817);
not I_551 (I14650,I15029);
nand I_552 (I15108,I15029,I14718);
and I_553 (I15125,I14786,I15108);
DFFARX1 I_554  ( .D(I15125), .CLK(I5694_clk), .RSTB(I14667_rst), .Q(I14629) );
DFFARX1 I_555  ( .D(I15029), .CLK(I5694_clk), .RSTB(I14667_rst), .Q(I14632) );
DFFARX1 I_556  ( .D(I4911), .CLK(I5694_clk), .RSTB(I14667_rst), .Q(I15170) );
not I_557 (I15187,I15170);
nand I_558 (I15204,I15187,I14752);
and I_559 (I15221,I14981,I15204);
DFFARX1 I_560  ( .D(I15221), .CLK(I5694_clk), .RSTB(I14667_rst), .Q(I14659) );
or I_561 (I15252,I15187,I14998);
DFFARX1 I_562  ( .D(I15252), .CLK(I5694_clk), .RSTB(I14667_rst), .Q(I14644) );
nand I_563 (I14647,I15187,I15077);
not I_564 (I15330_rst,I5701);
not I_565 (I15347,I4863);
nor I_566 (I15364,I4775,I2367);
nand I_567 (I15381,I15364,I4591);
nor I_568 (I15398,I15347,I4775);
nand I_569 (I15415,I15398,I3135);
not I_570 (I15432,I15415);
not I_571 (I15449,I4775);
nor I_572 (I15319,I15415,I15449);
not I_573 (I15480,I15449);
nand I_574 (I15304,I15415,I15480);
not I_575 (I15511,I5287);
nor I_576 (I15528,I15511,I1951);
and I_577 (I15545,I15528,I5511);
or I_578 (I15562,I15545,I4623);
DFFARX1 I_579  ( .D(I15562), .CLK(I5694_clk), .RSTB(I15330_rst), .Q(I15579) );
nor I_580 (I15596,I15579,I15432);
DFFARX1 I_581  ( .D(I15579), .CLK(I5694_clk), .RSTB(I15330_rst), .Q(I15613) );
not I_582 (I15301,I15613);
nand I_583 (I15644,I15347,I5287);
and I_584 (I15661,I15644,I15596);
DFFARX1 I_585  ( .D(I15644), .CLK(I5694_clk), .RSTB(I15330_rst), .Q(I15298) );
DFFARX1 I_586  ( .D(I3447), .CLK(I5694_clk), .RSTB(I15330_rst), .Q(I15692) );
nor I_587 (I15709,I15692,I15415);
nand I_588 (I15316,I15579,I15709);
nor I_589 (I15740,I15692,I15480);
not I_590 (I15313,I15692);
nand I_591 (I15771,I15692,I15381);
and I_592 (I15788,I15449,I15771);
DFFARX1 I_593  ( .D(I15788), .CLK(I5694_clk), .RSTB(I15330_rst), .Q(I15292) );
DFFARX1 I_594  ( .D(I15692), .CLK(I5694_clk), .RSTB(I15330_rst), .Q(I15295) );
DFFARX1 I_595  ( .D(I3071), .CLK(I5694_clk), .RSTB(I15330_rst), .Q(I15833) );
not I_596 (I15850,I15833);
nand I_597 (I15867,I15850,I15415);
and I_598 (I15884,I15644,I15867);
DFFARX1 I_599  ( .D(I15884), .CLK(I5694_clk), .RSTB(I15330_rst), .Q(I15322) );
or I_600 (I15915,I15850,I15661);
DFFARX1 I_601  ( .D(I15915), .CLK(I5694_clk), .RSTB(I15330_rst), .Q(I15307) );
nand I_602 (I15310,I15850,I15740);
not I_603 (I15993_rst,I5701);
not I_604 (I16010,I2527);
nor I_605 (I16027,I5327,I1735);
nand I_606 (I16044,I16027,I4727);
nor I_607 (I16061,I16010,I5327);
nand I_608 (I16078,I16061,I1895);
not I_609 (I16095,I16078);
not I_610 (I16112,I5327);
nor I_611 (I15982,I16078,I16112);
not I_612 (I16143,I16112);
nand I_613 (I15967,I16078,I16143);
not I_614 (I16174,I4607);
nor I_615 (I16191,I16174,I3159);
and I_616 (I16208,I16191,I3215);
or I_617 (I16225,I16208,I3231);
DFFARX1 I_618  ( .D(I16225), .CLK(I5694_clk), .RSTB(I15993_rst), .Q(I16242) );
nor I_619 (I16259,I16242,I16095);
DFFARX1 I_620  ( .D(I16242), .CLK(I5694_clk), .RSTB(I15993_rst), .Q(I16276) );
not I_621 (I15964,I16276);
nand I_622 (I16307,I16010,I4607);
and I_623 (I16324,I16307,I16259);
DFFARX1 I_624  ( .D(I16307), .CLK(I5694_clk), .RSTB(I15993_rst), .Q(I15961) );
DFFARX1 I_625  ( .D(I4199), .CLK(I5694_clk), .RSTB(I15993_rst), .Q(I16355) );
nor I_626 (I16372,I16355,I16078);
nand I_627 (I15979,I16242,I16372);
nor I_628 (I16403,I16355,I16143);
not I_629 (I15976,I16355);
nand I_630 (I16434,I16355,I16044);
and I_631 (I16451,I16112,I16434);
DFFARX1 I_632  ( .D(I16451), .CLK(I5694_clk), .RSTB(I15993_rst), .Q(I15955) );
DFFARX1 I_633  ( .D(I16355), .CLK(I5694_clk), .RSTB(I15993_rst), .Q(I15958) );
DFFARX1 I_634  ( .D(I1215), .CLK(I5694_clk), .RSTB(I15993_rst), .Q(I16496) );
not I_635 (I16513,I16496);
nand I_636 (I16530,I16513,I16078);
and I_637 (I16547,I16307,I16530);
DFFARX1 I_638  ( .D(I16547), .CLK(I5694_clk), .RSTB(I15993_rst), .Q(I15985) );
or I_639 (I16578,I16513,I16324);
DFFARX1 I_640  ( .D(I16578), .CLK(I5694_clk), .RSTB(I15993_rst), .Q(I15970) );
nand I_641 (I15973,I16513,I16403);
not I_642 (I16656_rst,I5701);
not I_643 (I16673,I1959);
nor I_644 (I16690,I3295,I3807);
nand I_645 (I16707,I16690,I3255);
nor I_646 (I16724,I16673,I3295);
nand I_647 (I16741,I16724,I4127);
not I_648 (I16758,I16741);
not I_649 (I16775,I3295);
nor I_650 (I16645,I16741,I16775);
not I_651 (I16806,I16775);
nand I_652 (I16630,I16741,I16806);
not I_653 (I16837,I4191);
nor I_654 (I16854,I16837,I3487);
and I_655 (I16871,I16854,I4095);
or I_656 (I16888,I16871,I4439);
DFFARX1 I_657  ( .D(I16888), .CLK(I5694_clk), .RSTB(I16656_rst), .Q(I16905) );
nor I_658 (I16922,I16905,I16758);
DFFARX1 I_659  ( .D(I16905), .CLK(I5694_clk), .RSTB(I16656_rst), .Q(I16939) );
not I_660 (I16627,I16939);
nand I_661 (I16970,I16673,I4191);
and I_662 (I16987,I16970,I16922);
DFFARX1 I_663  ( .D(I16970), .CLK(I5694_clk), .RSTB(I16656_rst), .Q(I16624) );
DFFARX1 I_664  ( .D(I4103), .CLK(I5694_clk), .RSTB(I16656_rst), .Q(I17018) );
nor I_665 (I17035,I17018,I16741);
nand I_666 (I16642,I16905,I17035);
nor I_667 (I17066,I17018,I16806);
not I_668 (I16639,I17018);
nand I_669 (I17097,I17018,I16707);
and I_670 (I17114,I16775,I17097);
DFFARX1 I_671  ( .D(I17114), .CLK(I5694_clk), .RSTB(I16656_rst), .Q(I16618) );
DFFARX1 I_672  ( .D(I17018), .CLK(I5694_clk), .RSTB(I16656_rst), .Q(I16621) );
DFFARX1 I_673  ( .D(I4615), .CLK(I5694_clk), .RSTB(I16656_rst), .Q(I17159) );
not I_674 (I17176,I17159);
nand I_675 (I17193,I17176,I16741);
and I_676 (I17210,I16970,I17193);
DFFARX1 I_677  ( .D(I17210), .CLK(I5694_clk), .RSTB(I16656_rst), .Q(I16648) );
or I_678 (I17241,I17176,I16987);
DFFARX1 I_679  ( .D(I17241), .CLK(I5694_clk), .RSTB(I16656_rst), .Q(I16633) );
nand I_680 (I16636,I17176,I17066);
not I_681 (I17319_rst,I5701);
not I_682 (I17336,I3327);
nor I_683 (I17353,I3391,I1831);
nand I_684 (I17370,I17353,I4559);
nor I_685 (I17387,I17336,I3391);
nand I_686 (I17404,I17387,I4687);
not I_687 (I17421,I17404);
not I_688 (I17438,I3391);
nor I_689 (I17308,I17404,I17438);
not I_690 (I17469,I17438);
nand I_691 (I17293,I17404,I17469);
not I_692 (I17500,I3415);
nor I_693 (I17517,I17500,I1799);
and I_694 (I17534,I17517,I5007);
or I_695 (I17551,I17534,I5391);
DFFARX1 I_696  ( .D(I17551), .CLK(I5694_clk), .RSTB(I17319_rst), .Q(I17568) );
nor I_697 (I17585,I17568,I17421);
DFFARX1 I_698  ( .D(I17568), .CLK(I5694_clk), .RSTB(I17319_rst), .Q(I17602) );
not I_699 (I17290,I17602);
nand I_700 (I17633,I17336,I3415);
and I_701 (I17650,I17633,I17585);
DFFARX1 I_702  ( .D(I17633), .CLK(I5694_clk), .RSTB(I17319_rst), .Q(I17287) );
DFFARX1 I_703  ( .D(I2303), .CLK(I5694_clk), .RSTB(I17319_rst), .Q(I17681) );
nor I_704 (I17698,I17681,I17404);
nand I_705 (I17305,I17568,I17698);
nor I_706 (I17729,I17681,I17469);
not I_707 (I17302,I17681);
nand I_708 (I17760,I17681,I17370);
and I_709 (I17777,I17438,I17760);
DFFARX1 I_710  ( .D(I17777), .CLK(I5694_clk), .RSTB(I17319_rst), .Q(I17281) );
DFFARX1 I_711  ( .D(I17681), .CLK(I5694_clk), .RSTB(I17319_rst), .Q(I17284) );
DFFARX1 I_712  ( .D(I5671), .CLK(I5694_clk), .RSTB(I17319_rst), .Q(I17822) );
not I_713 (I17839,I17822);
nand I_714 (I17856,I17839,I17404);
and I_715 (I17873,I17633,I17856);
DFFARX1 I_716  ( .D(I17873), .CLK(I5694_clk), .RSTB(I17319_rst), .Q(I17311) );
or I_717 (I17904,I17839,I17650);
DFFARX1 I_718  ( .D(I17904), .CLK(I5694_clk), .RSTB(I17319_rst), .Q(I17296) );
nand I_719 (I17299,I17839,I17729);
not I_720 (I17982_rst,I5701);
not I_721 (I17999,I1479);
nor I_722 (I18016,I3887,I1231);
nand I_723 (I18033,I18016,I2399);
nor I_724 (I18050,I17999,I3887);
nand I_725 (I18067,I18050,I1455);
DFFARX1 I_726  ( .D(I18067), .CLK(I5694_clk), .RSTB(I17982_rst), .Q(I18084) );
not I_727 (I17953,I18084);
not I_728 (I18115,I3887);
not I_729 (I18132,I18115);
not I_730 (I18149,I1559);
nor I_731 (I18166,I18149,I4415);
and I_732 (I18183,I18166,I2391);
or I_733 (I18200,I18183,I2495);
DFFARX1 I_734  ( .D(I18200), .CLK(I5694_clk), .RSTB(I17982_rst), .Q(I18217) );
DFFARX1 I_735  ( .D(I18217), .CLK(I5694_clk), .RSTB(I17982_rst), .Q(I17950) );
DFFARX1 I_736  ( .D(I18217), .CLK(I5694_clk), .RSTB(I17982_rst), .Q(I18248) );
DFFARX1 I_737  ( .D(I18217), .CLK(I5694_clk), .RSTB(I17982_rst), .Q(I17944) );
nand I_738 (I18279,I17999,I1559);
nand I_739 (I18296,I18279,I18033);
and I_740 (I18313,I18115,I18296);
DFFARX1 I_741  ( .D(I18313), .CLK(I5694_clk), .RSTB(I17982_rst), .Q(I17974) );
and I_742 (I17947,I18279,I18248);
DFFARX1 I_743  ( .D(I1359), .CLK(I5694_clk), .RSTB(I17982_rst), .Q(I18358) );
nor I_744 (I17971,I18358,I18279);
nor I_745 (I18389,I18358,I18033);
nand I_746 (I17968,I18067,I18389);
not I_747 (I17965,I18358);
DFFARX1 I_748  ( .D(I5343), .CLK(I5694_clk), .RSTB(I17982_rst), .Q(I18434) );
not I_749 (I18451,I18434);
nor I_750 (I18468,I18451,I18132);
and I_751 (I18485,I18358,I18468);
or I_752 (I18502,I18279,I18485);
DFFARX1 I_753  ( .D(I18502), .CLK(I5694_clk), .RSTB(I17982_rst), .Q(I17959) );
not I_754 (I18533,I18451);
nor I_755 (I18550,I18358,I18533);
nand I_756 (I17962,I18451,I18550);
nand I_757 (I17956,I18115,I18533);
not I_758 (I18628_rst,I5701);
not I_759 (I18645,I3143);
nor I_760 (I18662,I5423,I2063);
nand I_761 (I18679,I18662,I3335);
nor I_762 (I18696,I18645,I5423);
nand I_763 (I18713,I18696,I4135);
DFFARX1 I_764  ( .D(I18713), .CLK(I5694_clk), .RSTB(I18628_rst), .Q(I18730) );
not I_765 (I18599,I18730);
not I_766 (I18761,I5423);
not I_767 (I18778,I18761);
not I_768 (I18795,I2239);
nor I_769 (I18812,I18795,I3383);
and I_770 (I18829,I18812,I2103);
or I_771 (I18846,I18829,I4167);
DFFARX1 I_772  ( .D(I18846), .CLK(I5694_clk), .RSTB(I18628_rst), .Q(I18863) );
DFFARX1 I_773  ( .D(I18863), .CLK(I5694_clk), .RSTB(I18628_rst), .Q(I18596) );
DFFARX1 I_774  ( .D(I18863), .CLK(I5694_clk), .RSTB(I18628_rst), .Q(I18894) );
DFFARX1 I_775  ( .D(I18863), .CLK(I5694_clk), .RSTB(I18628_rst), .Q(I18590) );
nand I_776 (I18925,I18645,I2239);
nand I_777 (I18942,I18925,I18679);
and I_778 (I18959,I18761,I18942);
DFFARX1 I_779  ( .D(I18959), .CLK(I5694_clk), .RSTB(I18628_rst), .Q(I18620) );
and I_780 (I18593,I18925,I18894);
DFFARX1 I_781  ( .D(I2271), .CLK(I5694_clk), .RSTB(I18628_rst), .Q(I19004) );
nor I_782 (I18617,I19004,I18925);
nor I_783 (I19035,I19004,I18679);
nand I_784 (I18614,I18713,I19035);
not I_785 (I18611,I19004);
DFFARX1 I_786  ( .D(I3999), .CLK(I5694_clk), .RSTB(I18628_rst), .Q(I19080) );
not I_787 (I19097,I19080);
nor I_788 (I19114,I19097,I18778);
and I_789 (I19131,I19004,I19114);
or I_790 (I19148,I18925,I19131);
DFFARX1 I_791  ( .D(I19148), .CLK(I5694_clk), .RSTB(I18628_rst), .Q(I18605) );
not I_792 (I19179,I19097);
nor I_793 (I19196,I19004,I19179);
nand I_794 (I18608,I19097,I19196);
nand I_795 (I18602,I18761,I19179);
not I_796 (I19274_rst,I5701);
not I_797 (I19291,I3583);
nor I_798 (I19308,I1591,I5639);
nand I_799 (I19325,I19308,I5591);
nor I_800 (I19342,I19291,I1591);
nand I_801 (I19359,I19342,I2199);
DFFARX1 I_802  ( .D(I19359), .CLK(I5694_clk), .RSTB(I19274_rst), .Q(I19376) );
not I_803 (I19245,I19376);
not I_804 (I19407,I1591);
not I_805 (I19424,I19407);
not I_806 (I19441,I3663);
nor I_807 (I19458,I19441,I2535);
and I_808 (I19475,I19458,I4383);
or I_809 (I19492,I19475,I2159);
DFFARX1 I_810  ( .D(I19492), .CLK(I5694_clk), .RSTB(I19274_rst), .Q(I19509) );
DFFARX1 I_811  ( .D(I19509), .CLK(I5694_clk), .RSTB(I19274_rst), .Q(I19242) );
DFFARX1 I_812  ( .D(I19509), .CLK(I5694_clk), .RSTB(I19274_rst), .Q(I19540) );
DFFARX1 I_813  ( .D(I19509), .CLK(I5694_clk), .RSTB(I19274_rst), .Q(I19236) );
nand I_814 (I19571,I19291,I3663);
nand I_815 (I19588,I19571,I19325);
and I_816 (I19605,I19407,I19588);
DFFARX1 I_817  ( .D(I19605), .CLK(I5694_clk), .RSTB(I19274_rst), .Q(I19266) );
and I_818 (I19239,I19571,I19540);
DFFARX1 I_819  ( .D(I5183), .CLK(I5694_clk), .RSTB(I19274_rst), .Q(I19650) );
nor I_820 (I19263,I19650,I19571);
nor I_821 (I19681,I19650,I19325);
nand I_822 (I19260,I19359,I19681);
not I_823 (I19257,I19650);
DFFARX1 I_824  ( .D(I5271), .CLK(I5694_clk), .RSTB(I19274_rst), .Q(I19726) );
not I_825 (I19743,I19726);
nor I_826 (I19760,I19743,I19424);
and I_827 (I19777,I19650,I19760);
or I_828 (I19794,I19571,I19777);
DFFARX1 I_829  ( .D(I19794), .CLK(I5694_clk), .RSTB(I19274_rst), .Q(I19251) );
not I_830 (I19825,I19743);
nor I_831 (I19842,I19650,I19825);
nand I_832 (I19254,I19743,I19842);
nand I_833 (I19248,I19407,I19825);
not I_834 (I19920_rst,I5701);
not I_835 (I19937,I5279);
nor I_836 (I19954,I2919,I4887);
nand I_837 (I19971,I19954,I1247);
nor I_838 (I19988,I19937,I2919);
nand I_839 (I20005,I19988,I2095);
DFFARX1 I_840  ( .D(I20005), .CLK(I5694_clk), .RSTB(I19920_rst), .Q(I20022) );
not I_841 (I19891,I20022);
not I_842 (I20053,I2919);
not I_843 (I20070,I20053);
not I_844 (I20087,I1863);
nor I_845 (I20104,I20087,I1711);
and I_846 (I20121,I20104,I3439);
or I_847 (I20138,I20121,I1671);
DFFARX1 I_848  ( .D(I20138), .CLK(I5694_clk), .RSTB(I19920_rst), .Q(I20155) );
DFFARX1 I_849  ( .D(I20155), .CLK(I5694_clk), .RSTB(I19920_rst), .Q(I19888) );
DFFARX1 I_850  ( .D(I20155), .CLK(I5694_clk), .RSTB(I19920_rst), .Q(I20186) );
DFFARX1 I_851  ( .D(I20155), .CLK(I5694_clk), .RSTB(I19920_rst), .Q(I19882) );
nand I_852 (I20217,I19937,I1863);
nand I_853 (I20234,I20217,I19971);
and I_854 (I20251,I20053,I20234);
DFFARX1 I_855  ( .D(I20251), .CLK(I5694_clk), .RSTB(I19920_rst), .Q(I19912) );
and I_856 (I19885,I20217,I20186);
DFFARX1 I_857  ( .D(I3479), .CLK(I5694_clk), .RSTB(I19920_rst), .Q(I20296) );
nor I_858 (I19909,I20296,I20217);
nor I_859 (I20327,I20296,I19971);
nand I_860 (I19906,I20005,I20327);
not I_861 (I19903,I20296);
DFFARX1 I_862  ( .D(I3111), .CLK(I5694_clk), .RSTB(I19920_rst), .Q(I20372) );
not I_863 (I20389,I20372);
nor I_864 (I20406,I20389,I20070);
and I_865 (I20423,I20296,I20406);
or I_866 (I20440,I20217,I20423);
DFFARX1 I_867  ( .D(I20440), .CLK(I5694_clk), .RSTB(I19920_rst), .Q(I19897) );
not I_868 (I20471,I20389);
nor I_869 (I20488,I20296,I20471);
nand I_870 (I19900,I20389,I20488);
nand I_871 (I19894,I20053,I20471);
not I_872 (I20566_rst,I5701);
not I_873 (I20583,I2079);
nor I_874 (I20600,I3847,I1551);
nand I_875 (I20617,I20600,I2375);
nor I_876 (I20634,I20583,I3847);
nand I_877 (I20651,I20634,I2991);
DFFARX1 I_878  ( .D(I20651), .CLK(I5694_clk), .RSTB(I20566_rst), .Q(I20668) );
not I_879 (I20537,I20668);
not I_880 (I20699,I3847);
not I_881 (I20716,I20699);
not I_882 (I20733,I2431);
nor I_883 (I20750,I20733,I2871);
and I_884 (I20767,I20750,I1703);
or I_885 (I20784,I20767,I2167);
DFFARX1 I_886  ( .D(I20784), .CLK(I5694_clk), .RSTB(I20566_rst), .Q(I20801) );
DFFARX1 I_887  ( .D(I20801), .CLK(I5694_clk), .RSTB(I20566_rst), .Q(I20534) );
DFFARX1 I_888  ( .D(I20801), .CLK(I5694_clk), .RSTB(I20566_rst), .Q(I20832) );
DFFARX1 I_889  ( .D(I20801), .CLK(I5694_clk), .RSTB(I20566_rst), .Q(I20528) );
nand I_890 (I20863,I20583,I2431);
nand I_891 (I20880,I20863,I20617);
and I_892 (I20897,I20699,I20880);
DFFARX1 I_893  ( .D(I20897), .CLK(I5694_clk), .RSTB(I20566_rst), .Q(I20558) );
and I_894 (I20531,I20863,I20832);
DFFARX1 I_895  ( .D(I1911), .CLK(I5694_clk), .RSTB(I20566_rst), .Q(I20942) );
nor I_896 (I20555,I20942,I20863);
nor I_897 (I20973,I20942,I20617);
nand I_898 (I20552,I20651,I20973);
not I_899 (I20549,I20942);
DFFARX1 I_900  ( .D(I4351), .CLK(I5694_clk), .RSTB(I20566_rst), .Q(I21018) );
not I_901 (I21035,I21018);
nor I_902 (I21052,I21035,I20716);
and I_903 (I21069,I20942,I21052);
or I_904 (I21086,I20863,I21069);
DFFARX1 I_905  ( .D(I21086), .CLK(I5694_clk), .RSTB(I20566_rst), .Q(I20543) );
not I_906 (I21117,I21035);
nor I_907 (I21134,I20942,I21117);
nand I_908 (I20546,I21035,I21134);
nand I_909 (I20540,I20699,I21117);
not I_910 (I21212_rst,I5701);
or I_911 (I21229,I1743,I4895);
or I_912 (I21246,I3911,I1743);
nor I_913 (I21263,I2575,I2407);
DFFARX1 I_914  ( .D(I21263), .CLK(I5694_clk), .RSTB(I21212_rst), .Q(I21280) );
DFFARX1 I_915  ( .D(I21263), .CLK(I5694_clk), .RSTB(I21212_rst), .Q(I21174) );
not I_916 (I21311,I2575);
and I_917 (I21328,I21311,I3175);
nor I_918 (I21345,I21328,I4895);
nor I_919 (I21362,I3263,I1855);
DFFARX1 I_920  ( .D(I21362), .CLK(I5694_clk), .RSTB(I21212_rst), .Q(I21379) );
not I_921 (I21396,I21379);
DFFARX1 I_922  ( .D(I21379), .CLK(I5694_clk), .RSTB(I21212_rst), .Q(I21183) );
nor I_923 (I21427,I3263,I3911);
and I_924 (I21177,I21427,I21280);
DFFARX1 I_925  ( .D(I1935), .CLK(I5694_clk), .RSTB(I21212_rst), .Q(I21458) );
and I_926 (I21475,I21458,I1823);
nand I_927 (I21492,I21475,I21246);
and I_928 (I21509,I21379,I21492);
DFFARX1 I_929  ( .D(I21509), .CLK(I5694_clk), .RSTB(I21212_rst), .Q(I21204) );
nor I_930 (I21201,I21475,I21345);
not I_931 (I21554,I21475);
nor I_932 (I21571,I21229,I21554);
nor I_933 (I21588,I21475,I21427);
nand I_934 (I21198,I21246,I21588);
nor I_935 (I21619,I21475,I21396);
not I_936 (I21195,I21475);
nand I_937 (I21186,I21475,I21396);
DFFARX1 I_938  ( .D(I3943), .CLK(I5694_clk), .RSTB(I21212_rst), .Q(I21664) );
and I_939 (I21681,I21664,I21571);
or I_940 (I21698,I21229,I21681);
DFFARX1 I_941  ( .D(I21698), .CLK(I5694_clk), .RSTB(I21212_rst), .Q(I21189) );
nand I_942 (I21192,I21664,I21619);
nand I_943 (I21743,I21664,I21345);
and I_944 (I21760,I21263,I21743);
DFFARX1 I_945  ( .D(I21760), .CLK(I5694_clk), .RSTB(I21212_rst), .Q(I21180) );
not I_946 (I21824_rst,I5701);
or I_947 (I21841,I4655,I5519);
or I_948 (I21858,I1375,I4655);
nor I_949 (I21875,I3831,I5135);
DFFARX1 I_950  ( .D(I21875), .CLK(I5694_clk), .RSTB(I21824_rst), .Q(I21892) );
DFFARX1 I_951  ( .D(I21875), .CLK(I5694_clk), .RSTB(I21824_rst), .Q(I21786) );
not I_952 (I21923,I3831);
and I_953 (I21940,I21923,I3679);
nor I_954 (I21957,I21940,I5519);
nor I_955 (I21974,I4247,I1415);
DFFARX1 I_956  ( .D(I21974), .CLK(I5694_clk), .RSTB(I21824_rst), .Q(I21991) );
not I_957 (I22008,I21991);
DFFARX1 I_958  ( .D(I21991), .CLK(I5694_clk), .RSTB(I21824_rst), .Q(I21795) );
nor I_959 (I22039,I4247,I1375);
and I_960 (I21789,I22039,I21892);
DFFARX1 I_961  ( .D(I5599), .CLK(I5694_clk), .RSTB(I21824_rst), .Q(I22070) );
and I_962 (I22087,I22070,I1271);
nand I_963 (I22104,I22087,I21858);
and I_964 (I22121,I21991,I22104);
DFFARX1 I_965  ( .D(I22121), .CLK(I5694_clk), .RSTB(I21824_rst), .Q(I21816) );
nor I_966 (I21813,I22087,I21957);
not I_967 (I22166,I22087);
nor I_968 (I22183,I21841,I22166);
nor I_969 (I22200,I22087,I22039);
nand I_970 (I21810,I21858,I22200);
nor I_971 (I22231,I22087,I22008);
not I_972 (I21807,I22087);
nand I_973 (I21798,I22087,I22008);
DFFARX1 I_974  ( .D(I4751), .CLK(I5694_clk), .RSTB(I21824_rst), .Q(I22276) );
and I_975 (I22293,I22276,I22183);
or I_976 (I22310,I21841,I22293);
DFFARX1 I_977  ( .D(I22310), .CLK(I5694_clk), .RSTB(I21824_rst), .Q(I21801) );
nand I_978 (I21804,I22276,I22231);
nand I_979 (I22355,I22276,I21957);
and I_980 (I22372,I21875,I22355);
DFFARX1 I_981  ( .D(I22372), .CLK(I5694_clk), .RSTB(I21824_rst), .Q(I21792) );
not I_982 (I22436_rst,I5701);
or I_983 (I22453,I4935,I2151);
or I_984 (I22470,I5359,I4935);
nor I_985 (I22487,I2823,I3367);
DFFARX1 I_986  ( .D(I22487), .CLK(I5694_clk), .RSTB(I22436_rst), .Q(I22504) );
DFFARX1 I_987  ( .D(I22487), .CLK(I5694_clk), .RSTB(I22436_rst), .Q(I22398) );
not I_988 (I22535,I2823);
and I_989 (I22552,I22535,I3063);
nor I_990 (I22569,I22552,I2151);
nor I_991 (I22586,I3495,I1335);
DFFARX1 I_992  ( .D(I22586), .CLK(I5694_clk), .RSTB(I22436_rst), .Q(I22603) );
not I_993 (I22620,I22603);
DFFARX1 I_994  ( .D(I22603), .CLK(I5694_clk), .RSTB(I22436_rst), .Q(I22407) );
nor I_995 (I22651,I3495,I5359);
and I_996 (I22401,I22651,I22504);
DFFARX1 I_997  ( .D(I2943), .CLK(I5694_clk), .RSTB(I22436_rst), .Q(I22682) );
and I_998 (I22699,I22682,I5031);
nand I_999 (I22716,I22699,I22470);
and I_1000 (I22733,I22603,I22716);
DFFARX1 I_1001  ( .D(I22733), .CLK(I5694_clk), .RSTB(I22436_rst), .Q(I22428) );
nor I_1002 (I22425,I22699,I22569);
not I_1003 (I22778,I22699);
nor I_1004 (I22795,I22453,I22778);
nor I_1005 (I22812,I22699,I22651);
nand I_1006 (I22422,I22470,I22812);
nor I_1007 (I22843,I22699,I22620);
not I_1008 (I22419,I22699);
nand I_1009 (I22410,I22699,I22620);
DFFARX1 I_1010  ( .D(I3703), .CLK(I5694_clk), .RSTB(I22436_rst), .Q(I22888) );
and I_1011 (I22905,I22888,I22795);
or I_1012 (I22922,I22453,I22905);
DFFARX1 I_1013  ( .D(I22922), .CLK(I5694_clk), .RSTB(I22436_rst), .Q(I22413) );
nand I_1014 (I22416,I22888,I22843);
nand I_1015 (I22967,I22888,I22569);
and I_1016 (I22984,I22487,I22967);
DFFARX1 I_1017  ( .D(I22984), .CLK(I5694_clk), .RSTB(I22436_rst), .Q(I22404) );
not I_1018 (I23048_rst,I5701);
nand I_1019 (I23065,I3607,I1623);
and I_1020 (I23082,I23065,I4343);
DFFARX1 I_1021  ( .D(I23082), .CLK(I5694_clk), .RSTB(I23048_rst), .Q(I23099) );
not I_1022 (I23116,I23099);
DFFARX1 I_1023  ( .D(I23099), .CLK(I5694_clk), .RSTB(I23048_rst), .Q(I23016) );
nor I_1024 (I23147,I4119,I1623);
DFFARX1 I_1025  ( .D(I5647), .CLK(I5694_clk), .RSTB(I23048_rst), .Q(I23164) );
DFFARX1 I_1026  ( .D(I23164), .CLK(I5694_clk), .RSTB(I23048_rst), .Q(I23181) );
not I_1027 (I23019,I23181);
DFFARX1 I_1028  ( .D(I23164), .CLK(I5694_clk), .RSTB(I23048_rst), .Q(I23212) );
and I_1029 (I23013,I23099,I23212);
nand I_1030 (I23243,I5295,I5415);
and I_1031 (I23260,I23243,I4543);
DFFARX1 I_1032  ( .D(I23260), .CLK(I5694_clk), .RSTB(I23048_rst), .Q(I23277) );
nor I_1033 (I23294,I23277,I23116);
not I_1034 (I23311,I23277);
nand I_1035 (I23022,I23099,I23311);
DFFARX1 I_1036  ( .D(I4975), .CLK(I5694_clk), .RSTB(I23048_rst), .Q(I23342) );
and I_1037 (I23359,I23342,I1871);
nor I_1038 (I23376,I23359,I23277);
nor I_1039 (I23393,I23359,I23311);
nand I_1040 (I23028,I23147,I23393);
not I_1041 (I23031,I23359);
DFFARX1 I_1042  ( .D(I23359), .CLK(I5694_clk), .RSTB(I23048_rst), .Q(I23010) );
DFFARX1 I_1043  ( .D(I3863), .CLK(I5694_clk), .RSTB(I23048_rst), .Q(I23452) );
nand I_1044 (I23469,I23452,I23164);
and I_1045 (I23486,I23147,I23469);
DFFARX1 I_1046  ( .D(I23486), .CLK(I5694_clk), .RSTB(I23048_rst), .Q(I23040) );
nor I_1047 (I23037,I23452,I23359);
and I_1048 (I23531,I23452,I23294);
or I_1049 (I23548,I23147,I23531);
DFFARX1 I_1050  ( .D(I23548), .CLK(I5694_clk), .RSTB(I23048_rst), .Q(I23025) );
nand I_1051 (I23034,I23452,I23376);
not I_1052 (I23626_rst,I5701);
nand I_1053 (I23643,I5119,I1279);
and I_1054 (I23660,I23643,I1783);
DFFARX1 I_1055  ( .D(I23660), .CLK(I5694_clk), .RSTB(I23626_rst), .Q(I23677) );
not I_1056 (I23694,I23677);
DFFARX1 I_1057  ( .D(I23677), .CLK(I5694_clk), .RSTB(I23626_rst), .Q(I23594) );
nor I_1058 (I23725,I2223,I1279);
DFFARX1 I_1059  ( .D(I2639), .CLK(I5694_clk), .RSTB(I23626_rst), .Q(I23742) );
DFFARX1 I_1060  ( .D(I23742), .CLK(I5694_clk), .RSTB(I23626_rst), .Q(I23759) );
not I_1061 (I23597,I23759);
DFFARX1 I_1062  ( .D(I23742), .CLK(I5694_clk), .RSTB(I23626_rst), .Q(I23790) );
and I_1063 (I23591,I23677,I23790);
nand I_1064 (I23821,I3183,I3023);
and I_1065 (I23838,I23821,I2735);
DFFARX1 I_1066  ( .D(I23838), .CLK(I5694_clk), .RSTB(I23626_rst), .Q(I23855) );
nor I_1067 (I23872,I23855,I23694);
not I_1068 (I23889,I23855);
nand I_1069 (I23600,I23677,I23889);
DFFARX1 I_1070  ( .D(I1999), .CLK(I5694_clk), .RSTB(I23626_rst), .Q(I23920) );
and I_1071 (I23937,I23920,I4071);
nor I_1072 (I23954,I23937,I23855);
nor I_1073 (I23971,I23937,I23889);
nand I_1074 (I23606,I23725,I23971);
not I_1075 (I23609,I23937);
DFFARX1 I_1076  ( .D(I23937), .CLK(I5694_clk), .RSTB(I23626_rst), .Q(I23588) );
DFFARX1 I_1077  ( .D(I5087), .CLK(I5694_clk), .RSTB(I23626_rst), .Q(I24030) );
nand I_1078 (I24047,I24030,I23742);
and I_1079 (I24064,I23725,I24047);
DFFARX1 I_1080  ( .D(I24064), .CLK(I5694_clk), .RSTB(I23626_rst), .Q(I23618) );
nor I_1081 (I23615,I24030,I23937);
and I_1082 (I24109,I24030,I23872);
or I_1083 (I24126,I23725,I24109);
DFFARX1 I_1084  ( .D(I24126), .CLK(I5694_clk), .RSTB(I23626_rst), .Q(I23603) );
nand I_1085 (I23612,I24030,I23954);
not I_1086 (I24204_rst,I5701);
nand I_1087 (I24221,I3119,I4943);
and I_1088 (I24238,I24221,I2855);
DFFARX1 I_1089  ( .D(I24238), .CLK(I5694_clk), .RSTB(I24204_rst), .Q(I24255) );
not I_1090 (I24272,I24255);
DFFARX1 I_1091  ( .D(I24255), .CLK(I5694_clk), .RSTB(I24204_rst), .Q(I24172) );
nor I_1092 (I24303,I2839,I4943);
DFFARX1 I_1093  ( .D(I5023), .CLK(I5694_clk), .RSTB(I24204_rst), .Q(I24320) );
DFFARX1 I_1094  ( .D(I24320), .CLK(I5694_clk), .RSTB(I24204_rst), .Q(I24337) );
not I_1095 (I24175,I24337);
DFFARX1 I_1096  ( .D(I24320), .CLK(I5694_clk), .RSTB(I24204_rst), .Q(I24368) );
and I_1097 (I24169,I24255,I24368);
nand I_1098 (I24399,I3575,I3687);
and I_1099 (I24416,I24399,I3839);
DFFARX1 I_1100  ( .D(I24416), .CLK(I5694_clk), .RSTB(I24204_rst), .Q(I24433) );
nor I_1101 (I24450,I24433,I24272);
not I_1102 (I24467,I24433);
nand I_1103 (I24178,I24255,I24467);
DFFARX1 I_1104  ( .D(I5367), .CLK(I5694_clk), .RSTB(I24204_rst), .Q(I24498) );
and I_1105 (I24515,I24498,I4175);
nor I_1106 (I24532,I24515,I24433);
nor I_1107 (I24549,I24515,I24467);
nand I_1108 (I24184,I24303,I24549);
not I_1109 (I24187,I24515);
DFFARX1 I_1110  ( .D(I24515), .CLK(I5694_clk), .RSTB(I24204_rst), .Q(I24166) );
DFFARX1 I_1111  ( .D(I3095), .CLK(I5694_clk), .RSTB(I24204_rst), .Q(I24608) );
nand I_1112 (I24625,I24608,I24320);
and I_1113 (I24642,I24303,I24625);
DFFARX1 I_1114  ( .D(I24642), .CLK(I5694_clk), .RSTB(I24204_rst), .Q(I24196) );
nor I_1115 (I24193,I24608,I24515);
and I_1116 (I24687,I24608,I24450);
or I_1117 (I24704,I24303,I24687);
DFFARX1 I_1118  ( .D(I24704), .CLK(I5694_clk), .RSTB(I24204_rst), .Q(I24181) );
nand I_1119 (I24190,I24608,I24532);
not I_1120 (I24782_rst,I5701);
nand I_1121 (I24799,I2903,I2887);
and I_1122 (I24816,I24799,I2647);
DFFARX1 I_1123  ( .D(I24816), .CLK(I5694_clk), .RSTB(I24782_rst), .Q(I24833) );
not I_1124 (I24850,I24833);
DFFARX1 I_1125  ( .D(I24833), .CLK(I5694_clk), .RSTB(I24782_rst), .Q(I24750) );
nor I_1126 (I24881,I2743,I2887);
DFFARX1 I_1127  ( .D(I3247), .CLK(I5694_clk), .RSTB(I24782_rst), .Q(I24898) );
DFFARX1 I_1128  ( .D(I24898), .CLK(I5694_clk), .RSTB(I24782_rst), .Q(I24915) );
not I_1129 (I24753,I24915);
DFFARX1 I_1130  ( .D(I24898), .CLK(I5694_clk), .RSTB(I24782_rst), .Q(I24946) );
and I_1131 (I24747,I24833,I24946);
nand I_1132 (I24977,I2439,I5615);
and I_1133 (I24994,I24977,I3975);
DFFARX1 I_1134  ( .D(I24994), .CLK(I5694_clk), .RSTB(I24782_rst), .Q(I25011) );
nor I_1135 (I25028,I25011,I24850);
not I_1136 (I25045,I25011);
nand I_1137 (I24756,I24833,I25045);
DFFARX1 I_1138  ( .D(I5215), .CLK(I5694_clk), .RSTB(I24782_rst), .Q(I25076) );
and I_1139 (I25093,I25076,I2623);
nor I_1140 (I25110,I25093,I25011);
nor I_1141 (I25127,I25093,I25045);
nand I_1142 (I24762,I24881,I25127);
not I_1143 (I24765,I25093);
DFFARX1 I_1144  ( .D(I25093), .CLK(I5694_clk), .RSTB(I24782_rst), .Q(I24744) );
DFFARX1 I_1145  ( .D(I1839), .CLK(I5694_clk), .RSTB(I24782_rst), .Q(I25186) );
nand I_1146 (I25203,I25186,I24898);
and I_1147 (I25220,I24881,I25203);
DFFARX1 I_1148  ( .D(I25220), .CLK(I5694_clk), .RSTB(I24782_rst), .Q(I24774) );
nor I_1149 (I24771,I25186,I25093);
and I_1150 (I25265,I25186,I25028);
or I_1151 (I25282,I24881,I25265);
DFFARX1 I_1152  ( .D(I25282), .CLK(I5694_clk), .RSTB(I24782_rst), .Q(I24759) );
nand I_1153 (I24768,I25186,I25110);
not I_1154 (I25360_rst,I5701);
or I_1155 (I25377,I3223,I2687);
or I_1156 (I25394,I5167,I3223);
nor I_1157 (I25411,I1879,I2055);
not I_1158 (I25428,I25411);
DFFARX1 I_1159  ( .D(I25411), .CLK(I5694_clk), .RSTB(I25360_rst), .Q(I25328) );
nand I_1160 (I25459,I25411,I25377);
not I_1161 (I25476,I1879);
and I_1162 (I25493,I25476,I2343);
nor I_1163 (I25510,I25493,I2687);
nor I_1164 (I25527,I2783,I1535);
DFFARX1 I_1165  ( .D(I25527), .CLK(I5694_clk), .RSTB(I25360_rst), .Q(I25544) );
nor I_1166 (I25561,I25544,I25428);
not I_1167 (I25578,I25544);
nand I_1168 (I25334,I25411,I25578);
DFFARX1 I_1169  ( .D(I25544), .CLK(I5694_clk), .RSTB(I25360_rst), .Q(I25325) );
nor I_1170 (I25623,I2783,I5167);
nand I_1171 (I25640,I25394,I25623);
nor I_1172 (I25349,I25377,I25623);
and I_1173 (I25671,I25623,I25561);
or I_1174 (I25688,I25510,I25671);
DFFARX1 I_1175  ( .D(I25688), .CLK(I5694_clk), .RSTB(I25360_rst), .Q(I25337) );
DFFARX1 I_1176  ( .D(I4375), .CLK(I5694_clk), .RSTB(I25360_rst), .Q(I25719) );
and I_1177 (I25736,I25719,I3519);
not I_1178 (I25343,I25736);
DFFARX1 I_1179  ( .D(I25736), .CLK(I5694_clk), .RSTB(I25360_rst), .Q(I25767) );
not I_1180 (I25331,I25767);
and I_1181 (I25798,I25736,I25459);
DFFARX1 I_1182  ( .D(I25798), .CLK(I5694_clk), .RSTB(I25360_rst), .Q(I25322) );
DFFARX1 I_1183  ( .D(I2503), .CLK(I5694_clk), .RSTB(I25360_rst), .Q(I25829) );
and I_1184 (I25846,I25829,I25640);
DFFARX1 I_1185  ( .D(I25846), .CLK(I5694_clk), .RSTB(I25360_rst), .Q(I25352) );
nor I_1186 (I25877,I25829,I25736);
nand I_1187 (I25346,I25510,I25877);
nor I_1188 (I25908,I25829,I25578);
nand I_1189 (I25340,I25394,I25908);
not I_1190 (I25972_rst,I5701);
or I_1191 (I25989,I3711,I4487);
or I_1192 (I26006,I2815,I3711);
nor I_1193 (I26023,I1759,I3103);
not I_1194 (I26040,I26023);
DFFARX1 I_1195  ( .D(I26023), .CLK(I5694_clk), .RSTB(I25972_rst), .Q(I25940) );
nand I_1196 (I26071,I26023,I25989);
not I_1197 (I26088,I1759);
and I_1198 (I26105,I26088,I4231);
nor I_1199 (I26122,I26105,I4487);
nor I_1200 (I26139,I3727,I3463);
DFFARX1 I_1201  ( .D(I26139), .CLK(I5694_clk), .RSTB(I25972_rst), .Q(I26156) );
nor I_1202 (I26173,I26156,I26040);
not I_1203 (I26190,I26156);
nand I_1204 (I25946,I26023,I26190);
DFFARX1 I_1205  ( .D(I26156), .CLK(I5694_clk), .RSTB(I25972_rst), .Q(I25937) );
nor I_1206 (I26235,I3727,I2815);
nand I_1207 (I26252,I26006,I26235);
nor I_1208 (I25961,I25989,I26235);
and I_1209 (I26283,I26235,I26173);
or I_1210 (I26300,I26122,I26283);
DFFARX1 I_1211  ( .D(I26300), .CLK(I5694_clk), .RSTB(I25972_rst), .Q(I25949) );
DFFARX1 I_1212  ( .D(I5479), .CLK(I5694_clk), .RSTB(I25972_rst), .Q(I26331) );
and I_1213 (I26348,I26331,I2479);
not I_1214 (I25955,I26348);
DFFARX1 I_1215  ( .D(I26348), .CLK(I5694_clk), .RSTB(I25972_rst), .Q(I26379) );
not I_1216 (I25943,I26379);
and I_1217 (I26410,I26348,I26071);
DFFARX1 I_1218  ( .D(I26410), .CLK(I5694_clk), .RSTB(I25972_rst), .Q(I25934) );
DFFARX1 I_1219  ( .D(I2351), .CLK(I5694_clk), .RSTB(I25972_rst), .Q(I26441) );
and I_1220 (I26458,I26441,I26252);
DFFARX1 I_1221  ( .D(I26458), .CLK(I5694_clk), .RSTB(I25972_rst), .Q(I25964) );
nor I_1222 (I26489,I26441,I26348);
nand I_1223 (I25958,I26122,I26489);
nor I_1224 (I26520,I26441,I26190);
nand I_1225 (I25952,I26006,I26520);
not I_1226 (I26584_rst,I5701);
or I_1227 (I26601,I5455,I2119);
or I_1228 (I26618,I5439,I5455);
nor I_1229 (I26635,I4967,I4335);
or I_1230 (I26573,I26635,I26601);
not I_1231 (I26666,I4967);
and I_1232 (I26683,I26666,I2679);
nor I_1233 (I26700,I26683,I2119);
not I_1234 (I26717,I26700);
nor I_1235 (I26734,I1495,I4159);
DFFARX1 I_1236  ( .D(I26734), .CLK(I5694_clk), .RSTB(I26584_rst), .Q(I26751) );
nor I_1237 (I26768,I26751,I26700);
nand I_1238 (I26558,I26601,I26768);
nor I_1239 (I26799,I26751,I26717);
not I_1240 (I26555,I26751);
nor I_1241 (I26830,I1495,I5439);
or I_1242 (I26567,I26601,I26830);
DFFARX1 I_1243  ( .D(I1207), .CLK(I5694_clk), .RSTB(I26584_rst), .Q(I26861) );
and I_1244 (I26878,I26861,I1423);
nor I_1245 (I26895,I26878,I26751);
DFFARX1 I_1246  ( .D(I26895), .CLK(I5694_clk), .RSTB(I26584_rst), .Q(I26561) );
nor I_1247 (I26576,I26878,I26830);
not I_1248 (I26940,I26878);
nor I_1249 (I26957,I26618,I26940);
nand I_1250 (I26546,I26878,I26717);
DFFARX1 I_1251  ( .D(I3455), .CLK(I5694_clk), .RSTB(I26584_rst), .Q(I26988) );
nor I_1252 (I26564,I26988,I26618);
not I_1253 (I27019,I26988);
and I_1254 (I27036,I26830,I27019);
nor I_1255 (I26570,I26635,I27036);
and I_1256 (I27067,I26988,I26957);
or I_1257 (I27084,I26635,I27067);
DFFARX1 I_1258  ( .D(I27084), .CLK(I5694_clk), .RSTB(I26584_rst), .Q(I26549) );
nand I_1259 (I26552,I26988,I26799);
not I_1260 (I27162_rst,I5701);
nand I_1261 (I27179,I2775,I4767);
and I_1262 (I27196,I27179,I1903);
DFFARX1 I_1263  ( .D(I27196), .CLK(I5694_clk), .RSTB(I27162_rst), .Q(I27213) );
nor I_1264 (I27230,I4647,I4767);
nor I_1265 (I27247,I27230,I27213);
not I_1266 (I27145,I27230);
DFFARX1 I_1267  ( .D(I2047), .CLK(I5694_clk), .RSTB(I27162_rst), .Q(I27278) );
not I_1268 (I27295,I27278);
nor I_1269 (I27312,I27230,I27295);
nand I_1270 (I27148,I27278,I27247);
DFFARX1 I_1271  ( .D(I27278), .CLK(I5694_clk), .RSTB(I27162_rst), .Q(I27130) );
nand I_1272 (I27357,I5151,I1751);
and I_1273 (I27374,I27357,I4815);
DFFARX1 I_1274  ( .D(I27374), .CLK(I5694_clk), .RSTB(I27162_rst), .Q(I27391) );
nor I_1275 (I27151,I27391,I27213);
nand I_1276 (I27142,I27391,I27312);
DFFARX1 I_1277  ( .D(I2895), .CLK(I5694_clk), .RSTB(I27162_rst), .Q(I27436) );
and I_1278 (I27453,I27436,I2695);
DFFARX1 I_1279  ( .D(I27453), .CLK(I5694_clk), .RSTB(I27162_rst), .Q(I27470) );
not I_1280 (I27133,I27470);
nand I_1281 (I27501,I27453,I27391);
and I_1282 (I27518,I27213,I27501);
DFFARX1 I_1283  ( .D(I27518), .CLK(I5694_clk), .RSTB(I27162_rst), .Q(I27124) );
DFFARX1 I_1284  ( .D(I1223), .CLK(I5694_clk), .RSTB(I27162_rst), .Q(I27549) );
nand I_1285 (I27566,I27549,I27213);
and I_1286 (I27583,I27391,I27566);
DFFARX1 I_1287  ( .D(I27583), .CLK(I5694_clk), .RSTB(I27162_rst), .Q(I27154) );
not I_1288 (I27614,I27549);
nor I_1289 (I27631,I27230,I27614);
and I_1290 (I27648,I27549,I27631);
or I_1291 (I27665,I27453,I27648);
DFFARX1 I_1292  ( .D(I27665), .CLK(I5694_clk), .RSTB(I27162_rst), .Q(I27139) );
nand I_1293 (I27136,I27549,I27295);
DFFARX1 I_1294  ( .D(I27549), .CLK(I5694_clk), .RSTB(I27162_rst), .Q(I27127) );
not I_1295 (I27757_rst,I5701);
nand I_1296 (I27774,I3527,I3127);
and I_1297 (I27791,I27774,I2191);
DFFARX1 I_1298  ( .D(I27791), .CLK(I5694_clk), .RSTB(I27757_rst), .Q(I27808) );
nor I_1299 (I27825,I2767,I3127);
nor I_1300 (I27842,I27825,I27808);
not I_1301 (I27740,I27825);
DFFARX1 I_1302  ( .D(I1767), .CLK(I5694_clk), .RSTB(I27757_rst), .Q(I27873) );
not I_1303 (I27890,I27873);
nor I_1304 (I27907,I27825,I27890);
nand I_1305 (I27743,I27873,I27842);
DFFARX1 I_1306  ( .D(I27873), .CLK(I5694_clk), .RSTB(I27757_rst), .Q(I27725) );
nand I_1307 (I27952,I5247,I4463);
and I_1308 (I27969,I27952,I3543);
DFFARX1 I_1309  ( .D(I27969), .CLK(I5694_clk), .RSTB(I27757_rst), .Q(I27986) );
nor I_1310 (I27746,I27986,I27808);
nand I_1311 (I27737,I27986,I27907);
DFFARX1 I_1312  ( .D(I4783), .CLK(I5694_clk), .RSTB(I27757_rst), .Q(I28031) );
and I_1313 (I28048,I28031,I2663);
DFFARX1 I_1314  ( .D(I28048), .CLK(I5694_clk), .RSTB(I27757_rst), .Q(I28065) );
not I_1315 (I27728,I28065);
nand I_1316 (I28096,I28048,I27986);
and I_1317 (I28113,I27808,I28096);
DFFARX1 I_1318  ( .D(I28113), .CLK(I5694_clk), .RSTB(I27757_rst), .Q(I27719) );
DFFARX1 I_1319  ( .D(I3655), .CLK(I5694_clk), .RSTB(I27757_rst), .Q(I28144) );
nand I_1320 (I28161,I28144,I27808);
and I_1321 (I28178,I27986,I28161);
DFFARX1 I_1322  ( .D(I28178), .CLK(I5694_clk), .RSTB(I27757_rst), .Q(I27749) );
not I_1323 (I28209,I28144);
nor I_1324 (I28226,I27825,I28209);
and I_1325 (I28243,I28144,I28226);
or I_1326 (I28260,I28048,I28243);
DFFARX1 I_1327  ( .D(I28260), .CLK(I5694_clk), .RSTB(I27757_rst), .Q(I27734) );
nand I_1328 (I27731,I28144,I27890);
DFFARX1 I_1329  ( .D(I28144), .CLK(I5694_clk), .RSTB(I27757_rst), .Q(I27722) );
not I_1330 (I28352_rst,I5701);
nand I_1331 (I28369,I3567,I4183);
and I_1332 (I28386,I28369,I2007);
DFFARX1 I_1333  ( .D(I28386), .CLK(I5694_clk), .RSTB(I28352_rst), .Q(I28403) );
nor I_1334 (I28420,I3311,I4183);
DFFARX1 I_1335  ( .D(I3647), .CLK(I5694_clk), .RSTB(I28352_rst), .Q(I28437) );
nand I_1336 (I28454,I28437,I28420);
DFFARX1 I_1337  ( .D(I28437), .CLK(I5694_clk), .RSTB(I28352_rst), .Q(I28323) );
nand I_1338 (I28485,I4399,I1519);
and I_1339 (I28502,I28485,I3359);
DFFARX1 I_1340  ( .D(I28502), .CLK(I5694_clk), .RSTB(I28352_rst), .Q(I28519) );
not I_1341 (I28536,I28519);
nor I_1342 (I28553,I28403,I28536);
and I_1343 (I28570,I28420,I28553);
and I_1344 (I28587,I28519,I28454);
DFFARX1 I_1345  ( .D(I28587), .CLK(I5694_clk), .RSTB(I28352_rst), .Q(I28320) );
DFFARX1 I_1346  ( .D(I28519), .CLK(I5694_clk), .RSTB(I28352_rst), .Q(I28314) );
DFFARX1 I_1347  ( .D(I4711), .CLK(I5694_clk), .RSTB(I28352_rst), .Q(I28632) );
and I_1348 (I28649,I28632,I1775);
nand I_1349 (I28666,I28649,I28519);
nor I_1350 (I28341,I28649,I28420);
not I_1351 (I28697,I28649);
nor I_1352 (I28714,I28403,I28697);
nand I_1353 (I28332,I28437,I28714);
nand I_1354 (I28326,I28519,I28697);
or I_1355 (I28759,I28649,I28570);
DFFARX1 I_1356  ( .D(I28759), .CLK(I5694_clk), .RSTB(I28352_rst), .Q(I28329) );
DFFARX1 I_1357  ( .D(I3935), .CLK(I5694_clk), .RSTB(I28352_rst), .Q(I28790) );
and I_1358 (I28807,I28790,I28666);
DFFARX1 I_1359  ( .D(I28807), .CLK(I5694_clk), .RSTB(I28352_rst), .Q(I28344) );
nor I_1360 (I28838,I28790,I28403);
nand I_1361 (I28338,I28649,I28838);
not I_1362 (I28335,I28790);
DFFARX1 I_1363  ( .D(I28790), .CLK(I5694_clk), .RSTB(I28352_rst), .Q(I28883) );
and I_1364 (I28317,I28790,I28883);
not I_1365 (I28947_rst,I5701);
nand I_1366 (I28964,I3503,I3559);
and I_1367 (I28981,I28964,I3303);
DFFARX1 I_1368  ( .D(I28981), .CLK(I5694_clk), .RSTB(I28947_rst), .Q(I28998) );
nor I_1369 (I29015,I3239,I3559);
DFFARX1 I_1370  ( .D(I2255), .CLK(I5694_clk), .RSTB(I28947_rst), .Q(I29032) );
nand I_1371 (I29049,I29032,I29015);
DFFARX1 I_1372  ( .D(I29032), .CLK(I5694_clk), .RSTB(I28947_rst), .Q(I28918) );
nand I_1373 (I29080,I3079,I4703);
and I_1374 (I29097,I29080,I4391);
DFFARX1 I_1375  ( .D(I29097), .CLK(I5694_clk), .RSTB(I28947_rst), .Q(I29114) );
not I_1376 (I29131,I29114);
nor I_1377 (I29148,I28998,I29131);
and I_1378 (I29165,I29015,I29148);
and I_1379 (I29182,I29114,I29049);
DFFARX1 I_1380  ( .D(I29182), .CLK(I5694_clk), .RSTB(I28947_rst), .Q(I28915) );
DFFARX1 I_1381  ( .D(I29114), .CLK(I5694_clk), .RSTB(I28947_rst), .Q(I28909) );
DFFARX1 I_1382  ( .D(I3631), .CLK(I5694_clk), .RSTB(I28947_rst), .Q(I29227) );
and I_1383 (I29244,I29227,I4535);
nand I_1384 (I29261,I29244,I29114);
nor I_1385 (I28936,I29244,I29015);
not I_1386 (I29292,I29244);
nor I_1387 (I29309,I28998,I29292);
nand I_1388 (I28927,I29032,I29309);
nand I_1389 (I28921,I29114,I29292);
or I_1390 (I29354,I29244,I29165);
DFFARX1 I_1391  ( .D(I29354), .CLK(I5694_clk), .RSTB(I28947_rst), .Q(I28924) );
DFFARX1 I_1392  ( .D(I1303), .CLK(I5694_clk), .RSTB(I28947_rst), .Q(I29385) );
and I_1393 (I29402,I29385,I29261);
DFFARX1 I_1394  ( .D(I29402), .CLK(I5694_clk), .RSTB(I28947_rst), .Q(I28939) );
nor I_1395 (I29433,I29385,I28998);
nand I_1396 (I28933,I29244,I29433);
not I_1397 (I28930,I29385);
DFFARX1 I_1398  ( .D(I29385), .CLK(I5694_clk), .RSTB(I28947_rst), .Q(I29478) );
and I_1399 (I28912,I29385,I29478);
not I_1400 (I29542_rst,I5701);
nand I_1401 (I29559,I4671,I4423);
and I_1402 (I29576,I29559,I1343);
DFFARX1 I_1403  ( .D(I29576), .CLK(I5694_clk), .RSTB(I29542_rst), .Q(I29593) );
nor I_1404 (I29610,I2959,I4423);
DFFARX1 I_1405  ( .D(I4799), .CLK(I5694_clk), .RSTB(I29542_rst), .Q(I29627) );
nand I_1406 (I29644,I29627,I29610);
DFFARX1 I_1407  ( .D(I29627), .CLK(I5694_clk), .RSTB(I29542_rst), .Q(I29513) );
nand I_1408 (I29675,I1367,I4823);
and I_1409 (I29692,I29675,I2247);
DFFARX1 I_1410  ( .D(I29692), .CLK(I5694_clk), .RSTB(I29542_rst), .Q(I29709) );
not I_1411 (I29726,I29709);
nor I_1412 (I29743,I29593,I29726);
and I_1413 (I29760,I29610,I29743);
and I_1414 (I29777,I29709,I29644);
DFFARX1 I_1415  ( .D(I29777), .CLK(I5694_clk), .RSTB(I29542_rst), .Q(I29510) );
DFFARX1 I_1416  ( .D(I29709), .CLK(I5694_clk), .RSTB(I29542_rst), .Q(I29504) );
DFFARX1 I_1417  ( .D(I2071), .CLK(I5694_clk), .RSTB(I29542_rst), .Q(I29822) );
and I_1418 (I29839,I29822,I3471);
nand I_1419 (I29856,I29839,I29709);
nor I_1420 (I29531,I29839,I29610);
not I_1421 (I29887,I29839);
nor I_1422 (I29904,I29593,I29887);
nand I_1423 (I29522,I29627,I29904);
nand I_1424 (I29516,I29709,I29887);
or I_1425 (I29949,I29839,I29760);
DFFARX1 I_1426  ( .D(I29949), .CLK(I5694_clk), .RSTB(I29542_rst), .Q(I29519) );
DFFARX1 I_1427  ( .D(I4047), .CLK(I5694_clk), .RSTB(I29542_rst), .Q(I29980) );
and I_1428 (I29997,I29980,I29856);
DFFARX1 I_1429  ( .D(I29997), .CLK(I5694_clk), .RSTB(I29542_rst), .Q(I29534) );
nor I_1430 (I30028,I29980,I29593);
nand I_1431 (I29528,I29839,I30028);
not I_1432 (I29525,I29980);
DFFARX1 I_1433  ( .D(I29980), .CLK(I5694_clk), .RSTB(I29542_rst), .Q(I30073) );
and I_1434 (I29507,I29980,I30073);
not I_1435 (I30137_rst,I5701);
nand I_1436 (I30154,I3047,I4143);
and I_1437 (I30171,I30154,I3767);
DFFARX1 I_1438  ( .D(I30171), .CLK(I5694_clk), .RSTB(I30137_rst), .Q(I30188) );
nor I_1439 (I30205,I3783,I4143);
DFFARX1 I_1440  ( .D(I4735), .CLK(I5694_clk), .RSTB(I30137_rst), .Q(I30222) );
nand I_1441 (I30239,I30222,I30205);
DFFARX1 I_1442  ( .D(I30222), .CLK(I5694_clk), .RSTB(I30137_rst), .Q(I30108) );
nand I_1443 (I30270,I3879,I4719);
and I_1444 (I30287,I30270,I3855);
DFFARX1 I_1445  ( .D(I30287), .CLK(I5694_clk), .RSTB(I30137_rst), .Q(I30304) );
not I_1446 (I30321,I30304);
nor I_1447 (I30338,I30188,I30321);
and I_1448 (I30355,I30205,I30338);
and I_1449 (I30372,I30304,I30239);
DFFARX1 I_1450  ( .D(I30372), .CLK(I5694_clk), .RSTB(I30137_rst), .Q(I30105) );
DFFARX1 I_1451  ( .D(I30304), .CLK(I5694_clk), .RSTB(I30137_rst), .Q(I30099) );
DFFARX1 I_1452  ( .D(I5223), .CLK(I5694_clk), .RSTB(I30137_rst), .Q(I30417) );
and I_1453 (I30434,I30417,I3671);
nand I_1454 (I30451,I30434,I30304);
nor I_1455 (I30126,I30434,I30205);
not I_1456 (I30482,I30434);
nor I_1457 (I30499,I30188,I30482);
nand I_1458 (I30117,I30222,I30499);
nand I_1459 (I30111,I30304,I30482);
or I_1460 (I30544,I30434,I30355);
DFFARX1 I_1461  ( .D(I30544), .CLK(I5694_clk), .RSTB(I30137_rst), .Q(I30114) );
DFFARX1 I_1462  ( .D(I3775), .CLK(I5694_clk), .RSTB(I30137_rst), .Q(I30575) );
and I_1463 (I30592,I30575,I30451);
DFFARX1 I_1464  ( .D(I30592), .CLK(I5694_clk), .RSTB(I30137_rst), .Q(I30129) );
nor I_1465 (I30623,I30575,I30188);
nand I_1466 (I30123,I30434,I30623);
not I_1467 (I30120,I30575);
DFFARX1 I_1468  ( .D(I30575), .CLK(I5694_clk), .RSTB(I30137_rst), .Q(I30668) );
and I_1469 (I30102,I30575,I30668);
not I_1470 (I30732_rst,I5701);
not I_1471 (I30749,I1663);
nor I_1472 (I30766,I1919,I2039);
nand I_1473 (I30783,I30766,I2183);
nor I_1474 (I30800,I30749,I1919);
nand I_1475 (I30817,I30800,I4959);
not I_1476 (I30834,I1919);
not I_1477 (I30851,I30834);
not I_1478 (I30868,I4431);
nor I_1479 (I30885,I30868,I1631);
and I_1480 (I30902,I30885,I1399);
or I_1481 (I30919,I30902,I2607);
DFFARX1 I_1482  ( .D(I30919), .CLK(I5694_clk), .RSTB(I30732_rst), .Q(I30936) );
nand I_1483 (I30953,I30749,I4431);
or I_1484 (I30721,I30953,I30936);
not I_1485 (I30984,I30953);
nor I_1486 (I31001,I30936,I30984);
and I_1487 (I31018,I30834,I31001);
nand I_1488 (I30694,I30953,I30851);
DFFARX1 I_1489  ( .D(I2719), .CLK(I5694_clk), .RSTB(I30732_rst), .Q(I31049) );
or I_1490 (I30715,I31049,I30936);
nor I_1491 (I31080,I31049,I30817);
nor I_1492 (I31097,I31049,I30851);
nand I_1493 (I30700,I30783,I31097);
or I_1494 (I31128,I31049,I31018);
DFFARX1 I_1495  ( .D(I31128), .CLK(I5694_clk), .RSTB(I30732_rst), .Q(I30697) );
not I_1496 (I30703,I31049);
DFFARX1 I_1497  ( .D(I5159), .CLK(I5694_clk), .RSTB(I30732_rst), .Q(I31173) );
not I_1498 (I31190,I31173);
nor I_1499 (I31207,I31190,I30783);
DFFARX1 I_1500  ( .D(I31207), .CLK(I5694_clk), .RSTB(I30732_rst), .Q(I30709) );
nor I_1501 (I30724,I31049,I31190);
nor I_1502 (I30712,I31190,I30953);
not I_1503 (I31266,I31190);
and I_1504 (I31283,I30817,I31266);
nor I_1505 (I30718,I30953,I31283);
nand I_1506 (I30706,I31190,I31080);
not I_1507 (I31361_rst,I5701);
not I_1508 (I31378,I3959);
nor I_1509 (I31395,I4207,I4327);
nand I_1510 (I31412,I31395,I1407);
nor I_1511 (I31429,I31378,I4207);
nand I_1512 (I31446,I31429,I1983);
not I_1513 (I31463,I4207);
not I_1514 (I31480,I31463);
not I_1515 (I31497,I1719);
nor I_1516 (I31514,I31497,I1319);
and I_1517 (I31531,I31514,I5239);
or I_1518 (I31548,I31531,I1351);
DFFARX1 I_1519  ( .D(I31548), .CLK(I5694_clk), .RSTB(I31361_rst), .Q(I31565) );
nand I_1520 (I31582,I31378,I1719);
or I_1521 (I31350,I31582,I31565);
not I_1522 (I31613,I31582);
nor I_1523 (I31630,I31565,I31613);
and I_1524 (I31647,I31463,I31630);
nand I_1525 (I31323,I31582,I31480);
DFFARX1 I_1526  ( .D(I2135), .CLK(I5694_clk), .RSTB(I31361_rst), .Q(I31678) );
or I_1527 (I31344,I31678,I31565);
nor I_1528 (I31709,I31678,I31446);
nor I_1529 (I31726,I31678,I31480);
nand I_1530 (I31329,I31412,I31726);
or I_1531 (I31757,I31678,I31647);
DFFARX1 I_1532  ( .D(I31757), .CLK(I5694_clk), .RSTB(I31361_rst), .Q(I31326) );
not I_1533 (I31332,I31678);
DFFARX1 I_1534  ( .D(I4063), .CLK(I5694_clk), .RSTB(I31361_rst), .Q(I31802) );
not I_1535 (I31819,I31802);
nor I_1536 (I31836,I31819,I31412);
DFFARX1 I_1537  ( .D(I31836), .CLK(I5694_clk), .RSTB(I31361_rst), .Q(I31338) );
nor I_1538 (I31353,I31678,I31819);
nor I_1539 (I31341,I31819,I31582);
not I_1540 (I31895,I31819);
and I_1541 (I31912,I31446,I31895);
nor I_1542 (I31347,I31582,I31912);
nand I_1543 (I31335,I31819,I31709);
not I_1544 (I31990_rst,I5701);
not I_1545 (I32007,I2751);
nor I_1546 (I32024,I2471,I2935);
nand I_1547 (I32041,I32024,I4239);
nor I_1548 (I32058,I32007,I2471);
nand I_1549 (I32075,I32058,I3551);
not I_1550 (I32092,I2471);
not I_1551 (I32109,I32092);
not I_1552 (I32126,I1543);
nor I_1553 (I32143,I32126,I2759);
and I_1554 (I32160,I32143,I2015);
or I_1555 (I32177,I32160,I3599);
DFFARX1 I_1556  ( .D(I32177), .CLK(I5694_clk), .RSTB(I31990_rst), .Q(I32194) );
nand I_1557 (I32211,I32007,I1543);
or I_1558 (I31979,I32211,I32194);
not I_1559 (I32242,I32211);
nor I_1560 (I32259,I32194,I32242);
and I_1561 (I32276,I32092,I32259);
nand I_1562 (I31952,I32211,I32109);
DFFARX1 I_1563  ( .D(I3087), .CLK(I5694_clk), .RSTB(I31990_rst), .Q(I32307) );
or I_1564 (I31973,I32307,I32194);
nor I_1565 (I32338,I32307,I32075);
nor I_1566 (I32355,I32307,I32109);
nand I_1567 (I31958,I32041,I32355);
or I_1568 (I32386,I32307,I32276);
DFFARX1 I_1569  ( .D(I32386), .CLK(I5694_clk), .RSTB(I31990_rst), .Q(I31955) );
not I_1570 (I31961,I32307);
DFFARX1 I_1571  ( .D(I5375), .CLK(I5694_clk), .RSTB(I31990_rst), .Q(I32431) );
not I_1572 (I32448,I32431);
nor I_1573 (I32465,I32448,I32041);
DFFARX1 I_1574  ( .D(I32465), .CLK(I5694_clk), .RSTB(I31990_rst), .Q(I31967) );
nor I_1575 (I31982,I32307,I32448);
nor I_1576 (I31970,I32448,I32211);
not I_1577 (I32524,I32448);
and I_1578 (I32541,I32075,I32524);
nor I_1579 (I31976,I32211,I32541);
nand I_1580 (I31964,I32448,I32338);
not I_1581 (I32619_rst,I5701);
not I_1582 (I32636,I3759);
nor I_1583 (I32653,I2287,I2863);
nand I_1584 (I32670,I32653,I4007);
nor I_1585 (I32687,I32636,I2287);
nand I_1586 (I32704,I32687,I4567);
not I_1587 (I32721,I2287);
not I_1588 (I32738,I32721);
not I_1589 (I32755,I5463);
nor I_1590 (I32772,I32755,I5063);
and I_1591 (I32789,I32772,I2703);
or I_1592 (I32806,I32789,I4855);
DFFARX1 I_1593  ( .D(I32806), .CLK(I5694_clk), .RSTB(I32619_rst), .Q(I32823) );
nand I_1594 (I32840,I32636,I5463);
or I_1595 (I32608,I32840,I32823);
not I_1596 (I32871,I32840);
nor I_1597 (I32888,I32823,I32871);
and I_1598 (I32905,I32721,I32888);
nand I_1599 (I32581,I32840,I32738);
DFFARX1 I_1600  ( .D(I4991), .CLK(I5694_clk), .RSTB(I32619_rst), .Q(I32936) );
or I_1601 (I32602,I32936,I32823);
nor I_1602 (I32967,I32936,I32704);
nor I_1603 (I32984,I32936,I32738);
nand I_1604 (I32587,I32670,I32984);
or I_1605 (I33015,I32936,I32905);
DFFARX1 I_1606  ( .D(I33015), .CLK(I5694_clk), .RSTB(I32619_rst), .Q(I32584) );
not I_1607 (I32590,I32936);
DFFARX1 I_1608  ( .D(I5191), .CLK(I5694_clk), .RSTB(I32619_rst), .Q(I33060) );
not I_1609 (I33077,I33060);
nor I_1610 (I33094,I33077,I32670);
DFFARX1 I_1611  ( .D(I33094), .CLK(I5694_clk), .RSTB(I32619_rst), .Q(I32596) );
nor I_1612 (I32611,I32936,I33077);
nor I_1613 (I32599,I33077,I32840);
not I_1614 (I33153,I33077);
and I_1615 (I33170,I32704,I33153);
nor I_1616 (I32605,I32840,I33170);
nand I_1617 (I32593,I33077,I32967);
not I_1618 (I33248_rst,I5701);
not I_1619 (I33265,I2335);
nor I_1620 (I33282,I3271,I3423);
nand I_1621 (I33299,I33282,I1815);
nor I_1622 (I33316,I33265,I3271);
nand I_1623 (I33333,I33316,I2551);
not I_1624 (I33350,I3271);
not I_1625 (I33367,I33350);
not I_1626 (I33384,I4359);
nor I_1627 (I33401,I33384,I1239);
and I_1628 (I33418,I33401,I4743);
or I_1629 (I33435,I33418,I4407);
DFFARX1 I_1630  ( .D(I33435), .CLK(I5694_clk), .RSTB(I33248_rst), .Q(I33452) );
nand I_1631 (I33469,I33265,I4359);
or I_1632 (I33237,I33469,I33452);
not I_1633 (I33500,I33469);
nor I_1634 (I33517,I33452,I33500);
and I_1635 (I33534,I33350,I33517);
nand I_1636 (I33210,I33469,I33367);
DFFARX1 I_1637  ( .D(I1487), .CLK(I5694_clk), .RSTB(I33248_rst), .Q(I33565) );
or I_1638 (I33231,I33565,I33452);
nor I_1639 (I33596,I33565,I33333);
nor I_1640 (I33613,I33565,I33367);
nand I_1641 (I33216,I33299,I33613);
or I_1642 (I33644,I33565,I33534);
DFFARX1 I_1643  ( .D(I33644), .CLK(I5694_clk), .RSTB(I33248_rst), .Q(I33213) );
not I_1644 (I33219,I33565);
DFFARX1 I_1645  ( .D(I2711), .CLK(I5694_clk), .RSTB(I33248_rst), .Q(I33689) );
not I_1646 (I33706,I33689);
nor I_1647 (I33723,I33706,I33299);
DFFARX1 I_1648  ( .D(I33723), .CLK(I5694_clk), .RSTB(I33248_rst), .Q(I33225) );
nor I_1649 (I33240,I33565,I33706);
nor I_1650 (I33228,I33706,I33469);
not I_1651 (I33782,I33706);
and I_1652 (I33799,I33333,I33782);
nor I_1653 (I33234,I33469,I33799);
nand I_1654 (I33222,I33706,I33596);
not I_1655 (I33877_rst,I5701);
nand I_1656 (I33894,I2975,I4839);
and I_1657 (I33911,I33894,I1383);
DFFARX1 I_1658  ( .D(I33911), .CLK(I5694_clk), .RSTB(I33877_rst), .Q(I33928) );
not I_1659 (I33866,I33928);
DFFARX1 I_1660  ( .D(I33928), .CLK(I5694_clk), .RSTB(I33877_rst), .Q(I33959) );
not I_1661 (I33854,I33959);
nor I_1662 (I33990,I5687,I4839);
not I_1663 (I34007,I33990);
nor I_1664 (I34024,I33928,I34007);
DFFARX1 I_1665  ( .D(I1991), .CLK(I5694_clk), .RSTB(I33877_rst), .Q(I34041) );
not I_1666 (I34058,I34041);
nand I_1667 (I33857,I34041,I34007);
DFFARX1 I_1668  ( .D(I34041), .CLK(I5694_clk), .RSTB(I33877_rst), .Q(I34089) );
and I_1669 (I33842,I33928,I34089);
nand I_1670 (I34120,I2383,I4023);
and I_1671 (I34137,I34120,I5679);
DFFARX1 I_1672  ( .D(I34137), .CLK(I5694_clk), .RSTB(I33877_rst), .Q(I34154) );
nor I_1673 (I34171,I34154,I34058);
and I_1674 (I34188,I33990,I34171);
nor I_1675 (I34205,I34154,I33928);
DFFARX1 I_1676  ( .D(I34154), .CLK(I5694_clk), .RSTB(I33877_rst), .Q(I33848) );
DFFARX1 I_1677  ( .D(I2599), .CLK(I5694_clk), .RSTB(I33877_rst), .Q(I34236) );
and I_1678 (I34253,I34236,I3015);
or I_1679 (I34270,I34253,I34188);
DFFARX1 I_1680  ( .D(I34270), .CLK(I5694_clk), .RSTB(I33877_rst), .Q(I33860) );
nand I_1681 (I33869,I34253,I34205);
DFFARX1 I_1682  ( .D(I34253), .CLK(I5694_clk), .RSTB(I33877_rst), .Q(I33839) );
DFFARX1 I_1683  ( .D(I5207), .CLK(I5694_clk), .RSTB(I33877_rst), .Q(I34329) );
nand I_1684 (I33863,I34329,I34024);
DFFARX1 I_1685  ( .D(I34329), .CLK(I5694_clk), .RSTB(I33877_rst), .Q(I33851) );
nand I_1686 (I34374,I34329,I33990);
and I_1687 (I34391,I34041,I34374);
DFFARX1 I_1688  ( .D(I34391), .CLK(I5694_clk), .RSTB(I33877_rst), .Q(I33845) );
not I_1689 (I34455_rst,I5701);
nand I_1690 (I34472,I4455,I1295);
and I_1691 (I34489,I34472,I2911);
DFFARX1 I_1692  ( .D(I34489), .CLK(I5694_clk), .RSTB(I34455_rst), .Q(I34506) );
not I_1693 (I34444,I34506);
DFFARX1 I_1694  ( .D(I34506), .CLK(I5694_clk), .RSTB(I34455_rst), .Q(I34537) );
not I_1695 (I34432,I34537);
nor I_1696 (I34568,I5303,I1295);
not I_1697 (I34585,I34568);
nor I_1698 (I34602,I34506,I34585);
DFFARX1 I_1699  ( .D(I4215), .CLK(I5694_clk), .RSTB(I34455_rst), .Q(I34619) );
not I_1700 (I34636,I34619);
nand I_1701 (I34435,I34619,I34585);
DFFARX1 I_1702  ( .D(I34619), .CLK(I5694_clk), .RSTB(I34455_rst), .Q(I34667) );
and I_1703 (I34420,I34506,I34667);
nand I_1704 (I34698,I5623,I3407);
and I_1705 (I34715,I34698,I4847);
DFFARX1 I_1706  ( .D(I34715), .CLK(I5694_clk), .RSTB(I34455_rst), .Q(I34732) );
nor I_1707 (I34749,I34732,I34636);
and I_1708 (I34766,I34568,I34749);
nor I_1709 (I34783,I34732,I34506);
DFFARX1 I_1710  ( .D(I34732), .CLK(I5694_clk), .RSTB(I34455_rst), .Q(I34426) );
DFFARX1 I_1711  ( .D(I3815), .CLK(I5694_clk), .RSTB(I34455_rst), .Q(I34814) );
and I_1712 (I34831,I34814,I4807);
or I_1713 (I34848,I34831,I34766);
DFFARX1 I_1714  ( .D(I34848), .CLK(I5694_clk), .RSTB(I34455_rst), .Q(I34438) );
nand I_1715 (I34447,I34831,I34783);
DFFARX1 I_1716  ( .D(I34831), .CLK(I5694_clk), .RSTB(I34455_rst), .Q(I34417) );
DFFARX1 I_1717  ( .D(I4551), .CLK(I5694_clk), .RSTB(I34455_rst), .Q(I34907) );
nand I_1718 (I34441,I34907,I34602);
DFFARX1 I_1719  ( .D(I34907), .CLK(I5694_clk), .RSTB(I34455_rst), .Q(I34429) );
nand I_1720 (I34952,I34907,I34568);
and I_1721 (I34969,I34619,I34952);
DFFARX1 I_1722  ( .D(I34969), .CLK(I5694_clk), .RSTB(I34455_rst), .Q(I34423) );
not I_1723 (I35033_rst,I5701);
nand I_1724 (I35050,I2727,I1567);
and I_1725 (I35067,I35050,I3167);
DFFARX1 I_1726  ( .D(I35067), .CLK(I5694_clk), .RSTB(I35033_rst), .Q(I35084) );
not I_1727 (I35022,I35084);
DFFARX1 I_1728  ( .D(I35084), .CLK(I5694_clk), .RSTB(I35033_rst), .Q(I35115) );
not I_1729 (I35010,I35115);
nor I_1730 (I35146,I5143,I1567);
not I_1731 (I35163,I35146);
nor I_1732 (I35180,I35084,I35163);
DFFARX1 I_1733  ( .D(I4879), .CLK(I5694_clk), .RSTB(I35033_rst), .Q(I35197) );
not I_1734 (I35214,I35197);
nand I_1735 (I35013,I35197,I35163);
DFFARX1 I_1736  ( .D(I35197), .CLK(I5694_clk), .RSTB(I35033_rst), .Q(I35245) );
and I_1737 (I34998,I35084,I35245);
nand I_1738 (I35276,I2359,I2999);
and I_1739 (I35293,I35276,I3903);
DFFARX1 I_1740  ( .D(I35293), .CLK(I5694_clk), .RSTB(I35033_rst), .Q(I35310) );
nor I_1741 (I35327,I35310,I35214);
and I_1742 (I35344,I35146,I35327);
nor I_1743 (I35361,I35310,I35084);
DFFARX1 I_1744  ( .D(I35310), .CLK(I5694_clk), .RSTB(I35033_rst), .Q(I35004) );
DFFARX1 I_1745  ( .D(I4575), .CLK(I5694_clk), .RSTB(I35033_rst), .Q(I35392) );
and I_1746 (I35409,I35392,I2847);
or I_1747 (I35426,I35409,I35344);
DFFARX1 I_1748  ( .D(I35426), .CLK(I5694_clk), .RSTB(I35033_rst), .Q(I35016) );
nand I_1749 (I35025,I35409,I35361);
DFFARX1 I_1750  ( .D(I35409), .CLK(I5694_clk), .RSTB(I35033_rst), .Q(I34995) );
DFFARX1 I_1751  ( .D(I5231), .CLK(I5694_clk), .RSTB(I35033_rst), .Q(I35485) );
nand I_1752 (I35019,I35485,I35180);
DFFARX1 I_1753  ( .D(I35485), .CLK(I5694_clk), .RSTB(I35033_rst), .Q(I35007) );
nand I_1754 (I35530,I35485,I35146);
and I_1755 (I35547,I35197,I35530);
DFFARX1 I_1756  ( .D(I35547), .CLK(I5694_clk), .RSTB(I35033_rst), .Q(I35001) );
not I_1757 (I35611_rst,I5701);
nand I_1758 (I35628,I4303,I3823);
and I_1759 (I35645,I35628,I2087);
DFFARX1 I_1760  ( .D(I35645), .CLK(I5694_clk), .RSTB(I35611_rst), .Q(I35662) );
not I_1761 (I35600,I35662);
DFFARX1 I_1762  ( .D(I35662), .CLK(I5694_clk), .RSTB(I35611_rst), .Q(I35693) );
not I_1763 (I35588,I35693);
nor I_1764 (I35724,I3967,I3823);
not I_1765 (I35741,I35724);
nor I_1766 (I35758,I35662,I35741);
DFFARX1 I_1767  ( .D(I5199), .CLK(I5694_clk), .RSTB(I35611_rst), .Q(I35775) );
not I_1768 (I35792,I35775);
nand I_1769 (I35591,I35775,I35741);
DFFARX1 I_1770  ( .D(I35775), .CLK(I5694_clk), .RSTB(I35611_rst), .Q(I35823) );
and I_1771 (I35576,I35662,I35823);
nand I_1772 (I35854,I2631,I2311);
and I_1773 (I35871,I35854,I3591);
DFFARX1 I_1774  ( .D(I35871), .CLK(I5694_clk), .RSTB(I35611_rst), .Q(I35888) );
nor I_1775 (I35905,I35888,I35792);
and I_1776 (I35922,I35724,I35905);
nor I_1777 (I35939,I35888,I35662);
DFFARX1 I_1778  ( .D(I35888), .CLK(I5694_clk), .RSTB(I35611_rst), .Q(I35582) );
DFFARX1 I_1779  ( .D(I2983), .CLK(I5694_clk), .RSTB(I35611_rst), .Q(I35970) );
and I_1780 (I35987,I35970,I5095);
or I_1781 (I36004,I35987,I35922);
DFFARX1 I_1782  ( .D(I36004), .CLK(I5694_clk), .RSTB(I35611_rst), .Q(I35594) );
nand I_1783 (I35603,I35987,I35939);
DFFARX1 I_1784  ( .D(I35987), .CLK(I5694_clk), .RSTB(I35611_rst), .Q(I35573) );
DFFARX1 I_1785  ( .D(I5255), .CLK(I5694_clk), .RSTB(I35611_rst), .Q(I36063) );
nand I_1786 (I35597,I36063,I35758);
DFFARX1 I_1787  ( .D(I36063), .CLK(I5694_clk), .RSTB(I35611_rst), .Q(I35585) );
nand I_1788 (I36108,I36063,I35724);
and I_1789 (I36125,I35775,I36108);
DFFARX1 I_1790  ( .D(I36125), .CLK(I5694_clk), .RSTB(I35611_rst), .Q(I35579) );
not I_1791 (I36189_rst,I5701);
nand I_1792 (I36206,I5407,I3199);
and I_1793 (I36223,I36206,I5071);
DFFARX1 I_1794  ( .D(I36223), .CLK(I5694_clk), .RSTB(I36189_rst), .Q(I36240) );
not I_1795 (I36178,I36240);
DFFARX1 I_1796  ( .D(I36240), .CLK(I5694_clk), .RSTB(I36189_rst), .Q(I36271) );
not I_1797 (I36166,I36271);
nor I_1798 (I36302,I2415,I3199);
not I_1799 (I36319,I36302);
nor I_1800 (I36336,I36240,I36319);
DFFARX1 I_1801  ( .D(I2143), .CLK(I5694_clk), .RSTB(I36189_rst), .Q(I36353) );
not I_1802 (I36370,I36353);
nand I_1803 (I36169,I36353,I36319);
DFFARX1 I_1804  ( .D(I36353), .CLK(I5694_clk), .RSTB(I36189_rst), .Q(I36401) );
and I_1805 (I36154,I36240,I36401);
nand I_1806 (I36432,I2463,I5487);
and I_1807 (I36449,I36432,I5495);
DFFARX1 I_1808  ( .D(I36449), .CLK(I5694_clk), .RSTB(I36189_rst), .Q(I36466) );
nor I_1809 (I36483,I36466,I36370);
and I_1810 (I36500,I36302,I36483);
nor I_1811 (I36517,I36466,I36240);
DFFARX1 I_1812  ( .D(I36466), .CLK(I5694_clk), .RSTB(I36189_rst), .Q(I36160) );
DFFARX1 I_1813  ( .D(I1807), .CLK(I5694_clk), .RSTB(I36189_rst), .Q(I36548) );
and I_1814 (I36565,I36548,I4015);
or I_1815 (I36582,I36565,I36500);
DFFARX1 I_1816  ( .D(I36582), .CLK(I5694_clk), .RSTB(I36189_rst), .Q(I36172) );
nand I_1817 (I36181,I36565,I36517);
DFFARX1 I_1818  ( .D(I36565), .CLK(I5694_clk), .RSTB(I36189_rst), .Q(I36151) );
DFFARX1 I_1819  ( .D(I5535), .CLK(I5694_clk), .RSTB(I36189_rst), .Q(I36641) );
nand I_1820 (I36175,I36641,I36336);
DFFARX1 I_1821  ( .D(I36641), .CLK(I5694_clk), .RSTB(I36189_rst), .Q(I36163) );
nand I_1822 (I36686,I36641,I36302);
and I_1823 (I36703,I36353,I36686);
DFFARX1 I_1824  ( .D(I36703), .CLK(I5694_clk), .RSTB(I36189_rst), .Q(I36157) );
not I_1825 (I36767_rst,I5701);
nand I_1826 (I36784,I1511,I1391);
and I_1827 (I36801,I36784,I2519);
DFFARX1 I_1828  ( .D(I36801), .CLK(I5694_clk), .RSTB(I36767_rst), .Q(I36818) );
not I_1829 (I36756,I36818);
DFFARX1 I_1830  ( .D(I36818), .CLK(I5694_clk), .RSTB(I36767_rst), .Q(I36849) );
not I_1831 (I36744,I36849);
nor I_1832 (I36880,I3623,I1391);
not I_1833 (I36897,I36880);
nor I_1834 (I36914,I36818,I36897);
DFFARX1 I_1835  ( .D(I1679), .CLK(I5694_clk), .RSTB(I36767_rst), .Q(I36931) );
not I_1836 (I36948,I36931);
nand I_1837 (I36747,I36931,I36897);
DFFARX1 I_1838  ( .D(I36931), .CLK(I5694_clk), .RSTB(I36767_rst), .Q(I36979) );
and I_1839 (I36732,I36818,I36979);
nand I_1840 (I37010,I2487,I2559);
and I_1841 (I37027,I37010,I4599);
DFFARX1 I_1842  ( .D(I37027), .CLK(I5694_clk), .RSTB(I36767_rst), .Q(I37044) );
nor I_1843 (I37061,I37044,I36948);
and I_1844 (I37078,I36880,I37061);
nor I_1845 (I37095,I37044,I36818);
DFFARX1 I_1846  ( .D(I37044), .CLK(I5694_clk), .RSTB(I36767_rst), .Q(I36738) );
DFFARX1 I_1847  ( .D(I2215), .CLK(I5694_clk), .RSTB(I36767_rst), .Q(I37126) );
and I_1848 (I37143,I37126,I4039);
or I_1849 (I37160,I37143,I37078);
DFFARX1 I_1850  ( .D(I37160), .CLK(I5694_clk), .RSTB(I36767_rst), .Q(I36750) );
nand I_1851 (I36759,I37143,I37095);
DFFARX1 I_1852  ( .D(I37143), .CLK(I5694_clk), .RSTB(I36767_rst), .Q(I36729) );
DFFARX1 I_1853  ( .D(I1583), .CLK(I5694_clk), .RSTB(I36767_rst), .Q(I37219) );
nand I_1854 (I36753,I37219,I36914);
DFFARX1 I_1855  ( .D(I37219), .CLK(I5694_clk), .RSTB(I36767_rst), .Q(I36741) );
nand I_1856 (I37264,I37219,I36880);
and I_1857 (I37281,I36931,I37264);
DFFARX1 I_1858  ( .D(I37281), .CLK(I5694_clk), .RSTB(I36767_rst), .Q(I36735) );
not I_1859 (I37345_rst,I5701);
nand I_1860 (I37362,I21195,I21189);
and I_1861 (I37379,I37362,I21201);
DFFARX1 I_1862  ( .D(I37379), .CLK(I5694_clk), .RSTB(I37345_rst), .Q(I37396) );
not I_1863 (I37413,I37396);
nor I_1864 (I37430,I21198,I21189);
or I_1865 (I37328,I37430,I37396);
not I_1866 (I37316,I37430);
DFFARX1 I_1867  ( .D(I21177), .CLK(I5694_clk), .RSTB(I37345_rst), .Q(I37475) );
nor I_1868 (I37492,I37475,I37430);
nand I_1869 (I37509,I21183,I21192);
and I_1870 (I37526,I37509,I21180);
DFFARX1 I_1871  ( .D(I37526), .CLK(I5694_clk), .RSTB(I37345_rst), .Q(I37543) );
nor I_1872 (I37325,I37543,I37396);
not I_1873 (I37574,I37543);
nor I_1874 (I37591,I37475,I37574);
DFFARX1 I_1875  ( .D(I21204), .CLK(I5694_clk), .RSTB(I37345_rst), .Q(I37608) );
and I_1876 (I37625,I37608,I21174);
or I_1877 (I37334,I37625,I37430);
nand I_1878 (I37313,I37625,I37591);
DFFARX1 I_1879  ( .D(I21186), .CLK(I5694_clk), .RSTB(I37345_rst), .Q(I37670) );
and I_1880 (I37687,I37670,I37413);
nor I_1881 (I37331,I37625,I37687);
nor I_1882 (I37718,I37670,I37475);
DFFARX1 I_1883  ( .D(I37718), .CLK(I5694_clk), .RSTB(I37345_rst), .Q(I37322) );
nor I_1884 (I37337,I37670,I37396);
not I_1885 (I37763,I37670);
nor I_1886 (I37780,I37543,I37763);
and I_1887 (I37797,I37430,I37780);
or I_1888 (I37814,I37625,I37797);
DFFARX1 I_1889  ( .D(I37814), .CLK(I5694_clk), .RSTB(I37345_rst), .Q(I37310) );
nand I_1890 (I37319,I37670,I37492);
nand I_1891 (I37307,I37670,I37574);
not I_1892 (I37906_rst,I5701);
nand I_1893 (I37923,I33210,I33213);
and I_1894 (I37940,I37923,I33219);
DFFARX1 I_1895  ( .D(I37940), .CLK(I5694_clk), .RSTB(I37906_rst), .Q(I37957) );
not I_1896 (I37974,I37957);
nor I_1897 (I37991,I33231,I33213);
or I_1898 (I37889,I37991,I37957);
not I_1899 (I37877,I37991);
DFFARX1 I_1900  ( .D(I33240), .CLK(I5694_clk), .RSTB(I37906_rst), .Q(I38036) );
nor I_1901 (I38053,I38036,I37991);
nand I_1902 (I38070,I33228,I33225);
and I_1903 (I38087,I38070,I33237);
DFFARX1 I_1904  ( .D(I38087), .CLK(I5694_clk), .RSTB(I37906_rst), .Q(I38104) );
nor I_1905 (I37886,I38104,I37957);
not I_1906 (I38135,I38104);
nor I_1907 (I38152,I38036,I38135);
DFFARX1 I_1908  ( .D(I33234), .CLK(I5694_clk), .RSTB(I37906_rst), .Q(I38169) );
and I_1909 (I38186,I38169,I33222);
or I_1910 (I37895,I38186,I37991);
nand I_1911 (I37874,I38186,I38152);
DFFARX1 I_1912  ( .D(I33216), .CLK(I5694_clk), .RSTB(I37906_rst), .Q(I38231) );
and I_1913 (I38248,I38231,I37974);
nor I_1914 (I37892,I38186,I38248);
nor I_1915 (I38279,I38231,I38036);
DFFARX1 I_1916  ( .D(I38279), .CLK(I5694_clk), .RSTB(I37906_rst), .Q(I37883) );
nor I_1917 (I37898,I38231,I37957);
not I_1918 (I38324,I38231);
nor I_1919 (I38341,I38104,I38324);
and I_1920 (I38358,I37991,I38341);
or I_1921 (I38375,I38186,I38358);
DFFARX1 I_1922  ( .D(I38375), .CLK(I5694_clk), .RSTB(I37906_rst), .Q(I37871) );
nand I_1923 (I37880,I38231,I38053);
nand I_1924 (I37868,I38231,I38135);
not I_1925 (I38467_rst,I5701);
nand I_1926 (I38484,I10796,I10793);
and I_1927 (I38501,I38484,I10790);
DFFARX1 I_1928  ( .D(I38501), .CLK(I5694_clk), .RSTB(I38467_rst), .Q(I38518) );
not I_1929 (I38535,I38518);
nor I_1930 (I38552,I10814,I10793);
or I_1931 (I38450,I38552,I38518);
not I_1932 (I38438,I38552);
DFFARX1 I_1933  ( .D(I10808), .CLK(I5694_clk), .RSTB(I38467_rst), .Q(I38597) );
nor I_1934 (I38614,I38597,I38552);
nand I_1935 (I38631,I10787,I10799);
and I_1936 (I38648,I38631,I10802);
DFFARX1 I_1937  ( .D(I38648), .CLK(I5694_clk), .RSTB(I38467_rst), .Q(I38665) );
nor I_1938 (I38447,I38665,I38518);
not I_1939 (I38696,I38665);
nor I_1940 (I38713,I38597,I38696);
DFFARX1 I_1941  ( .D(I10811), .CLK(I5694_clk), .RSTB(I38467_rst), .Q(I38730) );
and I_1942 (I38747,I38730,I10817);
or I_1943 (I38456,I38747,I38552);
nand I_1944 (I38435,I38747,I38713);
DFFARX1 I_1945  ( .D(I10805), .CLK(I5694_clk), .RSTB(I38467_rst), .Q(I38792) );
and I_1946 (I38809,I38792,I38535);
nor I_1947 (I38453,I38747,I38809);
nor I_1948 (I38840,I38792,I38597);
DFFARX1 I_1949  ( .D(I38840), .CLK(I5694_clk), .RSTB(I38467_rst), .Q(I38444) );
nor I_1950 (I38459,I38792,I38518);
not I_1951 (I38885,I38792);
nor I_1952 (I38902,I38665,I38885);
and I_1953 (I38919,I38552,I38902);
or I_1954 (I38936,I38747,I38919);
DFFARX1 I_1955  ( .D(I38936), .CLK(I5694_clk), .RSTB(I38467_rst), .Q(I38432) );
nand I_1956 (I38441,I38792,I38614);
nand I_1957 (I38429,I38792,I38696);
not I_1958 (I39028_rst,I5701);
nand I_1959 (I39045,I25352,I25334);
and I_1960 (I39062,I39045,I25343);
DFFARX1 I_1961  ( .D(I39062), .CLK(I5694_clk), .RSTB(I39028_rst), .Q(I39079) );
not I_1962 (I39096,I39079);
nor I_1963 (I39113,I25328,I25334);
or I_1964 (I39011,I39113,I39079);
not I_1965 (I38999,I39113);
DFFARX1 I_1966  ( .D(I25337), .CLK(I5694_clk), .RSTB(I39028_rst), .Q(I39158) );
nor I_1967 (I39175,I39158,I39113);
nand I_1968 (I39192,I25325,I25331);
and I_1969 (I39209,I39192,I25340);
DFFARX1 I_1970  ( .D(I39209), .CLK(I5694_clk), .RSTB(I39028_rst), .Q(I39226) );
nor I_1971 (I39008,I39226,I39079);
not I_1972 (I39257,I39226);
nor I_1973 (I39274,I39158,I39257);
DFFARX1 I_1974  ( .D(I25349), .CLK(I5694_clk), .RSTB(I39028_rst), .Q(I39291) );
and I_1975 (I39308,I39291,I25322);
or I_1976 (I39017,I39308,I39113);
nand I_1977 (I38996,I39308,I39274);
DFFARX1 I_1978  ( .D(I25346), .CLK(I5694_clk), .RSTB(I39028_rst), .Q(I39353) );
and I_1979 (I39370,I39353,I39096);
nor I_1980 (I39014,I39308,I39370);
nor I_1981 (I39401,I39353,I39158);
DFFARX1 I_1982  ( .D(I39401), .CLK(I5694_clk), .RSTB(I39028_rst), .Q(I39005) );
nor I_1983 (I39020,I39353,I39079);
not I_1984 (I39446,I39353);
nor I_1985 (I39463,I39226,I39446);
and I_1986 (I39480,I39113,I39463);
or I_1987 (I39497,I39308,I39480);
DFFARX1 I_1988  ( .D(I39497), .CLK(I5694_clk), .RSTB(I39028_rst), .Q(I38993) );
nand I_1989 (I39002,I39353,I39175);
nand I_1990 (I38990,I39353,I39257);
not I_1991 (I39589_rst,I5701);
not I_1992 (I39606,I23025);
nor I_1993 (I39623,I23013,I23019);
nand I_1994 (I39640,I39623,I23010);
DFFARX1 I_1995  ( .D(I39640), .CLK(I5694_clk), .RSTB(I39589_rst), .Q(I39563) );
nor I_1996 (I39671,I39606,I23013);
nand I_1997 (I39688,I39671,I23016);
not I_1998 (I39578,I39688);
DFFARX1 I_1999  ( .D(I39688), .CLK(I5694_clk), .RSTB(I39589_rst), .Q(I39560) );
not I_2000 (I39733,I23013);
not I_2001 (I39750,I39733);
not I_2002 (I39767,I23028);
nor I_2003 (I39784,I39767,I23040);
and I_2004 (I39801,I39784,I23022);
or I_2005 (I39818,I39801,I23037);
DFFARX1 I_2006  ( .D(I39818), .CLK(I5694_clk), .RSTB(I39589_rst), .Q(I39835) );
nor I_2007 (I39852,I39835,I39688);
nor I_2008 (I39869,I39835,I39750);
nand I_2009 (I39575,I39640,I39869);
nand I_2010 (I39900,I39606,I23028);
nand I_2011 (I39917,I39900,I39835);
and I_2012 (I39934,I39900,I39917);
DFFARX1 I_2013  ( .D(I39934), .CLK(I5694_clk), .RSTB(I39589_rst), .Q(I39557) );
DFFARX1 I_2014  ( .D(I39900), .CLK(I5694_clk), .RSTB(I39589_rst), .Q(I39965) );
and I_2015 (I39554,I39733,I39965);
DFFARX1 I_2016  ( .D(I23031), .CLK(I5694_clk), .RSTB(I39589_rst), .Q(I39996) );
not I_2017 (I40013,I39996);
nor I_2018 (I40030,I39688,I40013);
and I_2019 (I40047,I39996,I40030);
nand I_2020 (I39569,I39996,I39750);
DFFARX1 I_2021  ( .D(I39996), .CLK(I5694_clk), .RSTB(I39589_rst), .Q(I40078) );
not I_2022 (I39566,I40078);
DFFARX1 I_2023  ( .D(I23034), .CLK(I5694_clk), .RSTB(I39589_rst), .Q(I40109) );
not I_2024 (I40126,I40109);
or I_2025 (I40143,I40126,I40047);
DFFARX1 I_2026  ( .D(I40143), .CLK(I5694_clk), .RSTB(I39589_rst), .Q(I39572) );
nand I_2027 (I39581,I40126,I39852);
DFFARX1 I_2028  ( .D(I40126), .CLK(I5694_clk), .RSTB(I39589_rst), .Q(I39551) );
not I_2029 (I40235_rst,I5701);
not I_2030 (I40252,I12045);
nor I_2031 (I40269,I12075,I12054);
nand I_2032 (I40286,I40269,I12066);
DFFARX1 I_2033  ( .D(I40286), .CLK(I5694_clk), .RSTB(I40235_rst), .Q(I40209) );
nor I_2034 (I40317,I40252,I12075);
nand I_2035 (I40334,I40317,I12048);
not I_2036 (I40224,I40334);
DFFARX1 I_2037  ( .D(I40334), .CLK(I5694_clk), .RSTB(I40235_rst), .Q(I40206) );
not I_2038 (I40379,I12075);
not I_2039 (I40396,I40379);
not I_2040 (I40413,I12051);
nor I_2041 (I40430,I40413,I12069);
and I_2042 (I40447,I40430,I12060);
or I_2043 (I40464,I40447,I12057);
DFFARX1 I_2044  ( .D(I40464), .CLK(I5694_clk), .RSTB(I40235_rst), .Q(I40481) );
nor I_2045 (I40498,I40481,I40334);
nor I_2046 (I40515,I40481,I40396);
nand I_2047 (I40221,I40286,I40515);
nand I_2048 (I40546,I40252,I12051);
nand I_2049 (I40563,I40546,I40481);
and I_2050 (I40580,I40546,I40563);
DFFARX1 I_2051  ( .D(I40580), .CLK(I5694_clk), .RSTB(I40235_rst), .Q(I40203) );
DFFARX1 I_2052  ( .D(I40546), .CLK(I5694_clk), .RSTB(I40235_rst), .Q(I40611) );
and I_2053 (I40200,I40379,I40611);
DFFARX1 I_2054  ( .D(I12063), .CLK(I5694_clk), .RSTB(I40235_rst), .Q(I40642) );
not I_2055 (I40659,I40642);
nor I_2056 (I40676,I40334,I40659);
and I_2057 (I40693,I40642,I40676);
nand I_2058 (I40215,I40642,I40396);
DFFARX1 I_2059  ( .D(I40642), .CLK(I5694_clk), .RSTB(I40235_rst), .Q(I40724) );
not I_2060 (I40212,I40724);
DFFARX1 I_2061  ( .D(I12072), .CLK(I5694_clk), .RSTB(I40235_rst), .Q(I40755) );
not I_2062 (I40772,I40755);
or I_2063 (I40789,I40772,I40693);
DFFARX1 I_2064  ( .D(I40789), .CLK(I5694_clk), .RSTB(I40235_rst), .Q(I40218) );
nand I_2065 (I40227,I40772,I40498);
DFFARX1 I_2066  ( .D(I40772), .CLK(I5694_clk), .RSTB(I40235_rst), .Q(I40197) );
not I_2067 (I40881_rst,I5701);
not I_2068 (I40898,I30694);
nor I_2069 (I40915,I30709,I30724);
nand I_2070 (I40932,I40915,I30712);
DFFARX1 I_2071  ( .D(I40932), .CLK(I5694_clk), .RSTB(I40881_rst), .Q(I40855) );
nor I_2072 (I40963,I40898,I30709);
nand I_2073 (I40980,I40963,I30715);
not I_2074 (I40870,I40980);
DFFARX1 I_2075  ( .D(I40980), .CLK(I5694_clk), .RSTB(I40881_rst), .Q(I40852) );
not I_2076 (I41025,I30709);
not I_2077 (I41042,I41025);
not I_2078 (I41059,I30721);
nor I_2079 (I41076,I41059,I30718);
and I_2080 (I41093,I41076,I30697);
or I_2081 (I41110,I41093,I30706);
DFFARX1 I_2082  ( .D(I41110), .CLK(I5694_clk), .RSTB(I40881_rst), .Q(I41127) );
nor I_2083 (I41144,I41127,I40980);
nor I_2084 (I41161,I41127,I41042);
nand I_2085 (I40867,I40932,I41161);
nand I_2086 (I41192,I40898,I30721);
nand I_2087 (I41209,I41192,I41127);
and I_2088 (I41226,I41192,I41209);
DFFARX1 I_2089  ( .D(I41226), .CLK(I5694_clk), .RSTB(I40881_rst), .Q(I40849) );
DFFARX1 I_2090  ( .D(I41192), .CLK(I5694_clk), .RSTB(I40881_rst), .Q(I41257) );
and I_2091 (I40846,I41025,I41257);
DFFARX1 I_2092  ( .D(I30703), .CLK(I5694_clk), .RSTB(I40881_rst), .Q(I41288) );
not I_2093 (I41305,I41288);
nor I_2094 (I41322,I40980,I41305);
and I_2095 (I41339,I41288,I41322);
nand I_2096 (I40861,I41288,I41042);
DFFARX1 I_2097  ( .D(I41288), .CLK(I5694_clk), .RSTB(I40881_rst), .Q(I41370) );
not I_2098 (I40858,I41370);
DFFARX1 I_2099  ( .D(I30700), .CLK(I5694_clk), .RSTB(I40881_rst), .Q(I41401) );
not I_2100 (I41418,I41401);
or I_2101 (I41435,I41418,I41339);
DFFARX1 I_2102  ( .D(I41435), .CLK(I5694_clk), .RSTB(I40881_rst), .Q(I40864) );
nand I_2103 (I40873,I41418,I41144);
DFFARX1 I_2104  ( .D(I41418), .CLK(I5694_clk), .RSTB(I40881_rst), .Q(I40843) );
not I_2105 (I41527_rst,I5701);
not I_2106 (I41544,I31323);
nor I_2107 (I41561,I31338,I31353);
nand I_2108 (I41578,I41561,I31341);
DFFARX1 I_2109  ( .D(I41578), .CLK(I5694_clk), .RSTB(I41527_rst), .Q(I41501) );
nor I_2110 (I41609,I41544,I31338);
nand I_2111 (I41626,I41609,I31344);
not I_2112 (I41516,I41626);
DFFARX1 I_2113  ( .D(I41626), .CLK(I5694_clk), .RSTB(I41527_rst), .Q(I41498) );
not I_2114 (I41671,I31338);
not I_2115 (I41688,I41671);
not I_2116 (I41705,I31350);
nor I_2117 (I41722,I41705,I31347);
and I_2118 (I41739,I41722,I31326);
or I_2119 (I41756,I41739,I31335);
DFFARX1 I_2120  ( .D(I41756), .CLK(I5694_clk), .RSTB(I41527_rst), .Q(I41773) );
nor I_2121 (I41790,I41773,I41626);
nor I_2122 (I41807,I41773,I41688);
nand I_2123 (I41513,I41578,I41807);
nand I_2124 (I41838,I41544,I31350);
nand I_2125 (I41855,I41838,I41773);
and I_2126 (I41872,I41838,I41855);
DFFARX1 I_2127  ( .D(I41872), .CLK(I5694_clk), .RSTB(I41527_rst), .Q(I41495) );
DFFARX1 I_2128  ( .D(I41838), .CLK(I5694_clk), .RSTB(I41527_rst), .Q(I41903) );
and I_2129 (I41492,I41671,I41903);
DFFARX1 I_2130  ( .D(I31332), .CLK(I5694_clk), .RSTB(I41527_rst), .Q(I41934) );
not I_2131 (I41951,I41934);
nor I_2132 (I41968,I41626,I41951);
and I_2133 (I41985,I41934,I41968);
nand I_2134 (I41507,I41934,I41688);
DFFARX1 I_2135  ( .D(I41934), .CLK(I5694_clk), .RSTB(I41527_rst), .Q(I42016) );
not I_2136 (I41504,I42016);
DFFARX1 I_2137  ( .D(I31329), .CLK(I5694_clk), .RSTB(I41527_rst), .Q(I42047) );
not I_2138 (I42064,I42047);
or I_2139 (I42081,I42064,I41985);
DFFARX1 I_2140  ( .D(I42081), .CLK(I5694_clk), .RSTB(I41527_rst), .Q(I41510) );
nand I_2141 (I41519,I42064,I41790);
DFFARX1 I_2142  ( .D(I42064), .CLK(I5694_clk), .RSTB(I41527_rst), .Q(I41489) );
not I_2143 (I42173_rst,I5701);
not I_2144 (I42190,I15310);
nor I_2145 (I42207,I15307,I15295);
nand I_2146 (I42224,I42207,I15298);
DFFARX1 I_2147  ( .D(I42224), .CLK(I5694_clk), .RSTB(I42173_rst), .Q(I42147) );
nor I_2148 (I42255,I42190,I15307);
nand I_2149 (I42272,I42255,I15304);
not I_2150 (I42162,I42272);
DFFARX1 I_2151  ( .D(I42272), .CLK(I5694_clk), .RSTB(I42173_rst), .Q(I42144) );
not I_2152 (I42317,I15307);
not I_2153 (I42334,I42317);
not I_2154 (I42351,I15316);
nor I_2155 (I42368,I42351,I15292);
and I_2156 (I42385,I42368,I15313);
or I_2157 (I42402,I42385,I15301);
DFFARX1 I_2158  ( .D(I42402), .CLK(I5694_clk), .RSTB(I42173_rst), .Q(I42419) );
nor I_2159 (I42436,I42419,I42272);
nor I_2160 (I42453,I42419,I42334);
nand I_2161 (I42159,I42224,I42453);
nand I_2162 (I42484,I42190,I15316);
nand I_2163 (I42501,I42484,I42419);
and I_2164 (I42518,I42484,I42501);
DFFARX1 I_2165  ( .D(I42518), .CLK(I5694_clk), .RSTB(I42173_rst), .Q(I42141) );
DFFARX1 I_2166  ( .D(I42484), .CLK(I5694_clk), .RSTB(I42173_rst), .Q(I42549) );
and I_2167 (I42138,I42317,I42549);
DFFARX1 I_2168  ( .D(I15322), .CLK(I5694_clk), .RSTB(I42173_rst), .Q(I42580) );
not I_2169 (I42597,I42580);
nor I_2170 (I42614,I42272,I42597);
and I_2171 (I42631,I42580,I42614);
nand I_2172 (I42153,I42580,I42334);
DFFARX1 I_2173  ( .D(I42580), .CLK(I5694_clk), .RSTB(I42173_rst), .Q(I42662) );
not I_2174 (I42150,I42662);
DFFARX1 I_2175  ( .D(I15319), .CLK(I5694_clk), .RSTB(I42173_rst), .Q(I42693) );
not I_2176 (I42710,I42693);
or I_2177 (I42727,I42710,I42631);
DFFARX1 I_2178  ( .D(I42727), .CLK(I5694_clk), .RSTB(I42173_rst), .Q(I42156) );
nand I_2179 (I42165,I42710,I42436);
DFFARX1 I_2180  ( .D(I42710), .CLK(I5694_clk), .RSTB(I42173_rst), .Q(I42135) );
not I_2181 (I42819_rst,I5701);
not I_2182 (I42836,I16636);
nor I_2183 (I42853,I16633,I16621);
nand I_2184 (I42870,I42853,I16624);
DFFARX1 I_2185  ( .D(I42870), .CLK(I5694_clk), .RSTB(I42819_rst), .Q(I42793) );
nor I_2186 (I42901,I42836,I16633);
nand I_2187 (I42918,I42901,I16630);
not I_2188 (I42808,I42918);
DFFARX1 I_2189  ( .D(I42918), .CLK(I5694_clk), .RSTB(I42819_rst), .Q(I42790) );
not I_2190 (I42963,I16633);
not I_2191 (I42980,I42963);
not I_2192 (I42997,I16642);
nor I_2193 (I43014,I42997,I16618);
and I_2194 (I43031,I43014,I16639);
or I_2195 (I43048,I43031,I16627);
DFFARX1 I_2196  ( .D(I43048), .CLK(I5694_clk), .RSTB(I42819_rst), .Q(I43065) );
nor I_2197 (I43082,I43065,I42918);
nor I_2198 (I43099,I43065,I42980);
nand I_2199 (I42805,I42870,I43099);
nand I_2200 (I43130,I42836,I16642);
nand I_2201 (I43147,I43130,I43065);
and I_2202 (I43164,I43130,I43147);
DFFARX1 I_2203  ( .D(I43164), .CLK(I5694_clk), .RSTB(I42819_rst), .Q(I42787) );
DFFARX1 I_2204  ( .D(I43130), .CLK(I5694_clk), .RSTB(I42819_rst), .Q(I43195) );
and I_2205 (I42784,I42963,I43195);
DFFARX1 I_2206  ( .D(I16648), .CLK(I5694_clk), .RSTB(I42819_rst), .Q(I43226) );
not I_2207 (I43243,I43226);
nor I_2208 (I43260,I42918,I43243);
and I_2209 (I43277,I43226,I43260);
nand I_2210 (I42799,I43226,I42980);
DFFARX1 I_2211  ( .D(I43226), .CLK(I5694_clk), .RSTB(I42819_rst), .Q(I43308) );
not I_2212 (I42796,I43308);
DFFARX1 I_2213  ( .D(I16645), .CLK(I5694_clk), .RSTB(I42819_rst), .Q(I43339) );
not I_2214 (I43356,I43339);
or I_2215 (I43373,I43356,I43277);
DFFARX1 I_2216  ( .D(I43373), .CLK(I5694_clk), .RSTB(I42819_rst), .Q(I42802) );
nand I_2217 (I42811,I43356,I43082);
DFFARX1 I_2218  ( .D(I43356), .CLK(I5694_clk), .RSTB(I42819_rst), .Q(I42781) );
not I_2219 (I43465_rst,I5701);
not I_2220 (I43482,I5707);
nor I_2221 (I43499,I5719,I5704);
nand I_2222 (I43516,I43499,I5716);
DFFARX1 I_2223  ( .D(I43516), .CLK(I5694_clk), .RSTB(I43465_rst), .Q(I43439) );
nor I_2224 (I43547,I43482,I5719);
nand I_2225 (I43564,I43547,I5734);
not I_2226 (I43454,I43564);
DFFARX1 I_2227  ( .D(I43564), .CLK(I5694_clk), .RSTB(I43465_rst), .Q(I43436) );
not I_2228 (I43609,I5719);
not I_2229 (I43626,I43609);
not I_2230 (I43643,I5710);
nor I_2231 (I43660,I43643,I5722);
and I_2232 (I43677,I43660,I5713);
or I_2233 (I43694,I43677,I5728);
DFFARX1 I_2234  ( .D(I43694), .CLK(I5694_clk), .RSTB(I43465_rst), .Q(I43711) );
nor I_2235 (I43728,I43711,I43564);
nor I_2236 (I43745,I43711,I43626);
nand I_2237 (I43451,I43516,I43745);
nand I_2238 (I43776,I43482,I5710);
nand I_2239 (I43793,I43776,I43711);
and I_2240 (I43810,I43776,I43793);
DFFARX1 I_2241  ( .D(I43810), .CLK(I5694_clk), .RSTB(I43465_rst), .Q(I43433) );
DFFARX1 I_2242  ( .D(I43776), .CLK(I5694_clk), .RSTB(I43465_rst), .Q(I43841) );
and I_2243 (I43430,I43609,I43841);
DFFARX1 I_2244  ( .D(I5731), .CLK(I5694_clk), .RSTB(I43465_rst), .Q(I43872) );
not I_2245 (I43889,I43872);
nor I_2246 (I43906,I43564,I43889);
and I_2247 (I43923,I43872,I43906);
nand I_2248 (I43445,I43872,I43626);
DFFARX1 I_2249  ( .D(I43872), .CLK(I5694_clk), .RSTB(I43465_rst), .Q(I43954) );
not I_2250 (I43442,I43954);
DFFARX1 I_2251  ( .D(I5725), .CLK(I5694_clk), .RSTB(I43465_rst), .Q(I43985) );
not I_2252 (I44002,I43985);
or I_2253 (I44019,I44002,I43923);
DFFARX1 I_2254  ( .D(I44019), .CLK(I5694_clk), .RSTB(I43465_rst), .Q(I43448) );
nand I_2255 (I43457,I44002,I43728);
DFFARX1 I_2256  ( .D(I44002), .CLK(I5694_clk), .RSTB(I43465_rst), .Q(I43427) );
not I_2257 (I44111_rst,I5701);
not I_2258 (I44128,I12658);
nor I_2259 (I44145,I12655,I12643);
nand I_2260 (I44162,I44145,I12646);
DFFARX1 I_2261  ( .D(I44162), .CLK(I5694_clk), .RSTB(I44111_rst), .Q(I44085) );
nor I_2262 (I44193,I44128,I12655);
nand I_2263 (I44210,I44193,I12652);
not I_2264 (I44100,I44210);
DFFARX1 I_2265  ( .D(I44210), .CLK(I5694_clk), .RSTB(I44111_rst), .Q(I44082) );
not I_2266 (I44255,I12655);
not I_2267 (I44272,I44255);
not I_2268 (I44289,I12664);
nor I_2269 (I44306,I44289,I12640);
and I_2270 (I44323,I44306,I12661);
or I_2271 (I44340,I44323,I12649);
DFFARX1 I_2272  ( .D(I44340), .CLK(I5694_clk), .RSTB(I44111_rst), .Q(I44357) );
nor I_2273 (I44374,I44357,I44210);
nor I_2274 (I44391,I44357,I44272);
nand I_2275 (I44097,I44162,I44391);
nand I_2276 (I44422,I44128,I12664);
nand I_2277 (I44439,I44422,I44357);
and I_2278 (I44456,I44422,I44439);
DFFARX1 I_2279  ( .D(I44456), .CLK(I5694_clk), .RSTB(I44111_rst), .Q(I44079) );
DFFARX1 I_2280  ( .D(I44422), .CLK(I5694_clk), .RSTB(I44111_rst), .Q(I44487) );
and I_2281 (I44076,I44255,I44487);
DFFARX1 I_2282  ( .D(I12670), .CLK(I5694_clk), .RSTB(I44111_rst), .Q(I44518) );
not I_2283 (I44535,I44518);
nor I_2284 (I44552,I44210,I44535);
and I_2285 (I44569,I44518,I44552);
nand I_2286 (I44091,I44518,I44272);
DFFARX1 I_2287  ( .D(I44518), .CLK(I5694_clk), .RSTB(I44111_rst), .Q(I44600) );
not I_2288 (I44088,I44600);
DFFARX1 I_2289  ( .D(I12667), .CLK(I5694_clk), .RSTB(I44111_rst), .Q(I44631) );
not I_2290 (I44648,I44631);
or I_2291 (I44665,I44648,I44569);
DFFARX1 I_2292  ( .D(I44665), .CLK(I5694_clk), .RSTB(I44111_rst), .Q(I44094) );
nand I_2293 (I44103,I44648,I44374);
DFFARX1 I_2294  ( .D(I44648), .CLK(I5694_clk), .RSTB(I44111_rst), .Q(I44073) );
not I_2295 (I44757_rst,I5701);
not I_2296 (I44774,I17962);
nor I_2297 (I44791,I17971,I17944);
nand I_2298 (I44808,I44791,I17956);
DFFARX1 I_2299  ( .D(I44808), .CLK(I5694_clk), .RSTB(I44757_rst), .Q(I44728) );
nor I_2300 (I44839,I44774,I17971);
nand I_2301 (I44856,I44839,I17968);
nand I_2302 (I44873,I44856,I44808);
not I_2303 (I44890,I17971);
not I_2304 (I44907,I17947);
nor I_2305 (I44924,I44907,I17953);
and I_2306 (I44941,I44924,I17965);
or I_2307 (I44958,I44941,I17950);
DFFARX1 I_2308  ( .D(I44958), .CLK(I5694_clk), .RSTB(I44757_rst), .Q(I44975) );
nor I_2309 (I44992,I44975,I44856);
nand I_2310 (I44743,I44890,I44992);
not I_2311 (I44740,I44975);
and I_2312 (I45037,I44975,I44873);
DFFARX1 I_2313  ( .D(I45037), .CLK(I5694_clk), .RSTB(I44757_rst), .Q(I44725) );
DFFARX1 I_2314  ( .D(I44975), .CLK(I5694_clk), .RSTB(I44757_rst), .Q(I45068) );
and I_2315 (I44722,I44890,I45068);
nand I_2316 (I45099,I44774,I17947);
not I_2317 (I45116,I45099);
nor I_2318 (I45133,I44975,I45116);
DFFARX1 I_2319  ( .D(I17974), .CLK(I5694_clk), .RSTB(I44757_rst), .Q(I45150) );
nand I_2320 (I45167,I45150,I45099);
and I_2321 (I45184,I44890,I45167);
DFFARX1 I_2322  ( .D(I45184), .CLK(I5694_clk), .RSTB(I44757_rst), .Q(I44749) );
not I_2323 (I45215,I45150);
nand I_2324 (I44737,I45150,I45133);
nand I_2325 (I44731,I45150,I45116);
DFFARX1 I_2326  ( .D(I17959), .CLK(I5694_clk), .RSTB(I44757_rst), .Q(I45260) );
not I_2327 (I45277,I45260);
nor I_2328 (I44746,I45150,I45277);
nor I_2329 (I45308,I45277,I45215);
and I_2330 (I45325,I44856,I45308);
or I_2331 (I45342,I45099,I45325);
DFFARX1 I_2332  ( .D(I45342), .CLK(I5694_clk), .RSTB(I44757_rst), .Q(I44734) );
DFFARX1 I_2333  ( .D(I45277), .CLK(I5694_clk), .RSTB(I44757_rst), .Q(I44719) );
not I_2334 (I45420_rst,I5701);
not I_2335 (I45437,I42796);
nor I_2336 (I45454,I42784,I42808);
nand I_2337 (I45471,I45454,I42793);
DFFARX1 I_2338  ( .D(I45471), .CLK(I5694_clk), .RSTB(I45420_rst), .Q(I45391) );
nor I_2339 (I45502,I45437,I42784);
nand I_2340 (I45519,I45502,I42811);
nand I_2341 (I45536,I45519,I45471);
not I_2342 (I45553,I42784);
not I_2343 (I45570,I42781);
nor I_2344 (I45587,I45570,I42790);
and I_2345 (I45604,I45587,I42805);
or I_2346 (I45621,I45604,I42787);
DFFARX1 I_2347  ( .D(I45621), .CLK(I5694_clk), .RSTB(I45420_rst), .Q(I45638) );
nor I_2348 (I45655,I45638,I45519);
nand I_2349 (I45406,I45553,I45655);
not I_2350 (I45403,I45638);
and I_2351 (I45700,I45638,I45536);
DFFARX1 I_2352  ( .D(I45700), .CLK(I5694_clk), .RSTB(I45420_rst), .Q(I45388) );
DFFARX1 I_2353  ( .D(I45638), .CLK(I5694_clk), .RSTB(I45420_rst), .Q(I45731) );
and I_2354 (I45385,I45553,I45731);
nand I_2355 (I45762,I45437,I42781);
not I_2356 (I45779,I45762);
nor I_2357 (I45796,I45638,I45779);
DFFARX1 I_2358  ( .D(I42802), .CLK(I5694_clk), .RSTB(I45420_rst), .Q(I45813) );
nand I_2359 (I45830,I45813,I45762);
and I_2360 (I45847,I45553,I45830);
DFFARX1 I_2361  ( .D(I45847), .CLK(I5694_clk), .RSTB(I45420_rst), .Q(I45412) );
not I_2362 (I45878,I45813);
nand I_2363 (I45400,I45813,I45796);
nand I_2364 (I45394,I45813,I45779);
DFFARX1 I_2365  ( .D(I42799), .CLK(I5694_clk), .RSTB(I45420_rst), .Q(I45923) );
not I_2366 (I45940,I45923);
nor I_2367 (I45409,I45813,I45940);
nor I_2368 (I45971,I45940,I45878);
and I_2369 (I45988,I45519,I45971);
or I_2370 (I46005,I45762,I45988);
DFFARX1 I_2371  ( .D(I46005), .CLK(I5694_clk), .RSTB(I45420_rst), .Q(I45397) );
DFFARX1 I_2372  ( .D(I45940), .CLK(I5694_clk), .RSTB(I45420_rst), .Q(I45382) );
not I_2373 (I46083_rst,I5701);
not I_2374 (I46100,I29510);
nor I_2375 (I46117,I29525,I29507);
nand I_2376 (I46134,I46117,I29519);
DFFARX1 I_2377  ( .D(I46134), .CLK(I5694_clk), .RSTB(I46083_rst), .Q(I46054) );
nor I_2378 (I46165,I46100,I29525);
nand I_2379 (I46182,I46165,I29516);
nand I_2380 (I46199,I46182,I46134);
not I_2381 (I46216,I29525);
not I_2382 (I46233,I29534);
nor I_2383 (I46250,I46233,I29504);
and I_2384 (I46267,I46250,I29513);
or I_2385 (I46284,I46267,I29531);
DFFARX1 I_2386  ( .D(I46284), .CLK(I5694_clk), .RSTB(I46083_rst), .Q(I46301) );
nor I_2387 (I46318,I46301,I46182);
nand I_2388 (I46069,I46216,I46318);
not I_2389 (I46066,I46301);
and I_2390 (I46363,I46301,I46199);
DFFARX1 I_2391  ( .D(I46363), .CLK(I5694_clk), .RSTB(I46083_rst), .Q(I46051) );
DFFARX1 I_2392  ( .D(I46301), .CLK(I5694_clk), .RSTB(I46083_rst), .Q(I46394) );
and I_2393 (I46048,I46216,I46394);
nand I_2394 (I46425,I46100,I29534);
not I_2395 (I46442,I46425);
nor I_2396 (I46459,I46301,I46442);
DFFARX1 I_2397  ( .D(I29522), .CLK(I5694_clk), .RSTB(I46083_rst), .Q(I46476) );
nand I_2398 (I46493,I46476,I46425);
and I_2399 (I46510,I46216,I46493);
DFFARX1 I_2400  ( .D(I46510), .CLK(I5694_clk), .RSTB(I46083_rst), .Q(I46075) );
not I_2401 (I46541,I46476);
nand I_2402 (I46063,I46476,I46459);
nand I_2403 (I46057,I46476,I46442);
DFFARX1 I_2404  ( .D(I29528), .CLK(I5694_clk), .RSTB(I46083_rst), .Q(I46586) );
not I_2405 (I46603,I46586);
nor I_2406 (I46072,I46476,I46603);
nor I_2407 (I46634,I46603,I46541);
and I_2408 (I46651,I46182,I46634);
or I_2409 (I46668,I46425,I46651);
DFFARX1 I_2410  ( .D(I46668), .CLK(I5694_clk), .RSTB(I46083_rst), .Q(I46060) );
DFFARX1 I_2411  ( .D(I46603), .CLK(I5694_clk), .RSTB(I46083_rst), .Q(I46045) );
not I_2412 (I46746_rst,I5701);
or I_2413 (I46763,I37889,I37898);
or I_2414 (I46780,I37892,I37889);
DFFARX1 I_2415  ( .D(I46780), .CLK(I5694_clk), .RSTB(I46746_rst), .Q(I46720) );
nor I_2416 (I46811,I37868,I37871);
not I_2417 (I46828,I46811);
not I_2418 (I46845,I37868);
and I_2419 (I46862,I46845,I37880);
nor I_2420 (I46879,I46862,I37898);
nor I_2421 (I46896,I37886,I37877);
DFFARX1 I_2422  ( .D(I46896), .CLK(I5694_clk), .RSTB(I46746_rst), .Q(I46913) );
nand I_2423 (I46930,I46913,I46763);
and I_2424 (I46947,I46879,I46930);
DFFARX1 I_2425  ( .D(I46947), .CLK(I5694_clk), .RSTB(I46746_rst), .Q(I46714) );
nor I_2426 (I46978,I37886,I37892);
DFFARX1 I_2427  ( .D(I46978), .CLK(I5694_clk), .RSTB(I46746_rst), .Q(I46995) );
and I_2428 (I46711,I46811,I46995);
DFFARX1 I_2429  ( .D(I37883), .CLK(I5694_clk), .RSTB(I46746_rst), .Q(I47026) );
and I_2430 (I47043,I47026,I37874);
DFFARX1 I_2431  ( .D(I47043), .CLK(I5694_clk), .RSTB(I46746_rst), .Q(I47060) );
not I_2432 (I46723,I47060);
DFFARX1 I_2433  ( .D(I47043), .CLK(I5694_clk), .RSTB(I46746_rst), .Q(I46708) );
DFFARX1 I_2434  ( .D(I37895), .CLK(I5694_clk), .RSTB(I46746_rst), .Q(I47105) );
not I_2435 (I47122,I47105);
nor I_2436 (I47139,I46780,I47122);
and I_2437 (I47156,I47043,I47139);
or I_2438 (I47173,I46763,I47156);
DFFARX1 I_2439  ( .D(I47173), .CLK(I5694_clk), .RSTB(I46746_rst), .Q(I46729) );
nor I_2440 (I47204,I47105,I46913);
nand I_2441 (I46738,I46879,I47204);
nor I_2442 (I47235,I47105,I46828);
nand I_2443 (I46732,I46978,I47235);
not I_2444 (I46735,I47105);
nand I_2445 (I46726,I47105,I46828);
DFFARX1 I_2446  ( .D(I47105), .CLK(I5694_clk), .RSTB(I46746_rst), .Q(I46717) );
not I_2447 (I47341_rst,I5701);
or I_2448 (I47358,I32584,I32581);
or I_2449 (I47375,I32611,I32584);
DFFARX1 I_2450  ( .D(I47375), .CLK(I5694_clk), .RSTB(I47341_rst), .Q(I47315) );
nor I_2451 (I47406,I32590,I32596);
not I_2452 (I47423,I47406);
not I_2453 (I47440,I32590);
and I_2454 (I47457,I47440,I32587);
nor I_2455 (I47474,I47457,I32581);
nor I_2456 (I47491,I32599,I32608);
DFFARX1 I_2457  ( .D(I47491), .CLK(I5694_clk), .RSTB(I47341_rst), .Q(I47508) );
nand I_2458 (I47525,I47508,I47358);
and I_2459 (I47542,I47474,I47525);
DFFARX1 I_2460  ( .D(I47542), .CLK(I5694_clk), .RSTB(I47341_rst), .Q(I47309) );
nor I_2461 (I47573,I32599,I32611);
DFFARX1 I_2462  ( .D(I47573), .CLK(I5694_clk), .RSTB(I47341_rst), .Q(I47590) );
and I_2463 (I47306,I47406,I47590);
DFFARX1 I_2464  ( .D(I32602), .CLK(I5694_clk), .RSTB(I47341_rst), .Q(I47621) );
and I_2465 (I47638,I47621,I32593);
DFFARX1 I_2466  ( .D(I47638), .CLK(I5694_clk), .RSTB(I47341_rst), .Q(I47655) );
not I_2467 (I47318,I47655);
DFFARX1 I_2468  ( .D(I47638), .CLK(I5694_clk), .RSTB(I47341_rst), .Q(I47303) );
DFFARX1 I_2469  ( .D(I32605), .CLK(I5694_clk), .RSTB(I47341_rst), .Q(I47700) );
not I_2470 (I47717,I47700);
nor I_2471 (I47734,I47375,I47717);
and I_2472 (I47751,I47638,I47734);
or I_2473 (I47768,I47358,I47751);
DFFARX1 I_2474  ( .D(I47768), .CLK(I5694_clk), .RSTB(I47341_rst), .Q(I47324) );
nor I_2475 (I47799,I47700,I47508);
nand I_2476 (I47333,I47474,I47799);
nor I_2477 (I47830,I47700,I47423);
nand I_2478 (I47327,I47573,I47830);
not I_2479 (I47330,I47700);
nand I_2480 (I47321,I47700,I47423);
DFFARX1 I_2481  ( .D(I47700), .CLK(I5694_clk), .RSTB(I47341_rst), .Q(I47312) );
not I_2482 (I47936_rst,I5701);
or I_2483 (I47953,I24196,I24181);
or I_2484 (I47970,I24193,I24196);
DFFARX1 I_2485  ( .D(I47970), .CLK(I5694_clk), .RSTB(I47936_rst), .Q(I47910) );
nor I_2486 (I48001,I24175,I24166);
not I_2487 (I48018,I48001);
not I_2488 (I48035,I24175);
and I_2489 (I48052,I48035,I24190);
nor I_2490 (I48069,I48052,I24181);
nor I_2491 (I48086,I24169,I24187);
DFFARX1 I_2492  ( .D(I48086), .CLK(I5694_clk), .RSTB(I47936_rst), .Q(I48103) );
nand I_2493 (I48120,I48103,I47953);
and I_2494 (I48137,I48069,I48120);
DFFARX1 I_2495  ( .D(I48137), .CLK(I5694_clk), .RSTB(I47936_rst), .Q(I47904) );
nor I_2496 (I48168,I24169,I24193);
DFFARX1 I_2497  ( .D(I48168), .CLK(I5694_clk), .RSTB(I47936_rst), .Q(I48185) );
and I_2498 (I47901,I48001,I48185);
DFFARX1 I_2499  ( .D(I24178), .CLK(I5694_clk), .RSTB(I47936_rst), .Q(I48216) );
and I_2500 (I48233,I48216,I24172);
DFFARX1 I_2501  ( .D(I48233), .CLK(I5694_clk), .RSTB(I47936_rst), .Q(I48250) );
not I_2502 (I47913,I48250);
DFFARX1 I_2503  ( .D(I48233), .CLK(I5694_clk), .RSTB(I47936_rst), .Q(I47898) );
DFFARX1 I_2504  ( .D(I24184), .CLK(I5694_clk), .RSTB(I47936_rst), .Q(I48295) );
not I_2505 (I48312,I48295);
nor I_2506 (I48329,I47970,I48312);
and I_2507 (I48346,I48233,I48329);
or I_2508 (I48363,I47953,I48346);
DFFARX1 I_2509  ( .D(I48363), .CLK(I5694_clk), .RSTB(I47936_rst), .Q(I47919) );
nor I_2510 (I48394,I48295,I48103);
nand I_2511 (I47928,I48069,I48394);
nor I_2512 (I48425,I48295,I48018);
nand I_2513 (I47922,I48168,I48425);
not I_2514 (I47925,I48295);
nand I_2515 (I47916,I48295,I48018);
DFFARX1 I_2516  ( .D(I48295), .CLK(I5694_clk), .RSTB(I47936_rst), .Q(I47907) );
not I_2517 (I48531_rst,I5701);
or I_2518 (I48548,I44749,I44734);
or I_2519 (I48565,I44731,I44749);
DFFARX1 I_2520  ( .D(I48565), .CLK(I5694_clk), .RSTB(I48531_rst), .Q(I48505) );
nor I_2521 (I48596,I44719,I44728);
not I_2522 (I48613,I48596);
not I_2523 (I48630,I44719);
and I_2524 (I48647,I48630,I44743);
nor I_2525 (I48664,I48647,I44734);
nor I_2526 (I48681,I44722,I44737);
DFFARX1 I_2527  ( .D(I48681), .CLK(I5694_clk), .RSTB(I48531_rst), .Q(I48698) );
nand I_2528 (I48715,I48698,I48548);
and I_2529 (I48732,I48664,I48715);
DFFARX1 I_2530  ( .D(I48732), .CLK(I5694_clk), .RSTB(I48531_rst), .Q(I48499) );
nor I_2531 (I48763,I44722,I44731);
DFFARX1 I_2532  ( .D(I48763), .CLK(I5694_clk), .RSTB(I48531_rst), .Q(I48780) );
and I_2533 (I48496,I48596,I48780);
DFFARX1 I_2534  ( .D(I44725), .CLK(I5694_clk), .RSTB(I48531_rst), .Q(I48811) );
and I_2535 (I48828,I48811,I44746);
DFFARX1 I_2536  ( .D(I48828), .CLK(I5694_clk), .RSTB(I48531_rst), .Q(I48845) );
not I_2537 (I48508,I48845);
DFFARX1 I_2538  ( .D(I48828), .CLK(I5694_clk), .RSTB(I48531_rst), .Q(I48493) );
DFFARX1 I_2539  ( .D(I44740), .CLK(I5694_clk), .RSTB(I48531_rst), .Q(I48890) );
not I_2540 (I48907,I48890);
nor I_2541 (I48924,I48565,I48907);
and I_2542 (I48941,I48828,I48924);
or I_2543 (I48958,I48548,I48941);
DFFARX1 I_2544  ( .D(I48958), .CLK(I5694_clk), .RSTB(I48531_rst), .Q(I48514) );
nor I_2545 (I48989,I48890,I48698);
nand I_2546 (I48523,I48664,I48989);
nor I_2547 (I49020,I48890,I48613);
nand I_2548 (I48517,I48763,I49020);
not I_2549 (I48520,I48890);
nand I_2550 (I48511,I48890,I48613);
DFFARX1 I_2551  ( .D(I48890), .CLK(I5694_clk), .RSTB(I48531_rst), .Q(I48502) );
not I_2552 (I49126_rst,I5701);
or I_2553 (I49143,I35016,I34998);
not I_2554 (I49109,I49143);
DFFARX1 I_2555  ( .D(I49143), .CLK(I5694_clk), .RSTB(I49126_rst), .Q(I49088) );
or I_2556 (I49188,I35025,I35016);
nor I_2557 (I49205,I35007,I35022);
nor I_2558 (I49222,I49205,I49143);
not I_2559 (I49239,I35007);
and I_2560 (I49256,I49239,I35004);
nor I_2561 (I49273,I49256,I34998);
DFFARX1 I_2562  ( .D(I49273), .CLK(I5694_clk), .RSTB(I49126_rst), .Q(I49290) );
nor I_2563 (I49307,I35019,I34995);
DFFARX1 I_2564  ( .D(I49307), .CLK(I5694_clk), .RSTB(I49126_rst), .Q(I49324) );
nor I_2565 (I49115,I49324,I49273);
not I_2566 (I49355,I49324);
nor I_2567 (I49372,I35019,I35025);
nand I_2568 (I49389,I49273,I49372);
and I_2569 (I49406,I49188,I49389);
DFFARX1 I_2570  ( .D(I49406), .CLK(I5694_clk), .RSTB(I49126_rst), .Q(I49118) );
DFFARX1 I_2571  ( .D(I35013), .CLK(I5694_clk), .RSTB(I49126_rst), .Q(I49437) );
and I_2572 (I49454,I49437,I35001);
nor I_2573 (I49471,I49454,I49355);
and I_2574 (I49488,I49372,I49471);
or I_2575 (I49505,I49205,I49488);
DFFARX1 I_2576  ( .D(I49505), .CLK(I5694_clk), .RSTB(I49126_rst), .Q(I49103) );
not I_2577 (I49536,I49454);
nor I_2578 (I49553,I49143,I49536);
nand I_2579 (I49106,I49188,I49553);
nand I_2580 (I49100,I49324,I49536);
DFFARX1 I_2581  ( .D(I49454), .CLK(I5694_clk), .RSTB(I49126_rst), .Q(I49094) );
DFFARX1 I_2582  ( .D(I35010), .CLK(I5694_clk), .RSTB(I49126_rst), .Q(I49612) );
nand I_2583 (I49112,I49612,I49222);
DFFARX1 I_2584  ( .D(I49612), .CLK(I5694_clk), .RSTB(I49126_rst), .Q(I49643) );
not I_2585 (I49097,I49643);
and I_2586 (I49091,I49612,I49290);
not I_2587 (I49721_rst,I5701);
not I_2588 (I49738,I26549);
nor I_2589 (I49755,I26570,I26576);
nand I_2590 (I49772,I49755,I26564);
nor I_2591 (I49789,I49738,I26570);
nand I_2592 (I49806,I49789,I26546);
not I_2593 (I49823,I49806);
not I_2594 (I49840,I26570);
nor I_2595 (I49710,I49806,I49840);
not I_2596 (I49871,I49840);
nand I_2597 (I49695,I49806,I49871);
not I_2598 (I49902,I26552);
nor I_2599 (I49919,I49902,I26573);
and I_2600 (I49936,I49919,I26561);
or I_2601 (I49953,I49936,I26567);
DFFARX1 I_2602  ( .D(I49953), .CLK(I5694_clk), .RSTB(I49721_rst), .Q(I49970) );
nor I_2603 (I49987,I49970,I49823);
DFFARX1 I_2604  ( .D(I49970), .CLK(I5694_clk), .RSTB(I49721_rst), .Q(I50004) );
not I_2605 (I49692,I50004);
nand I_2606 (I50035,I49738,I26552);
and I_2607 (I50052,I50035,I49987);
DFFARX1 I_2608  ( .D(I50035), .CLK(I5694_clk), .RSTB(I49721_rst), .Q(I49689) );
DFFARX1 I_2609  ( .D(I26558), .CLK(I5694_clk), .RSTB(I49721_rst), .Q(I50083) );
nor I_2610 (I50100,I50083,I49806);
nand I_2611 (I49707,I49970,I50100);
nor I_2612 (I50131,I50083,I49871);
not I_2613 (I49704,I50083);
nand I_2614 (I50162,I50083,I49772);
and I_2615 (I50179,I49840,I50162);
DFFARX1 I_2616  ( .D(I50179), .CLK(I5694_clk), .RSTB(I49721_rst), .Q(I49683) );
DFFARX1 I_2617  ( .D(I50083), .CLK(I5694_clk), .RSTB(I49721_rst), .Q(I49686) );
DFFARX1 I_2618  ( .D(I26555), .CLK(I5694_clk), .RSTB(I49721_rst), .Q(I50224) );
not I_2619 (I50241,I50224);
nand I_2620 (I50258,I50241,I49806);
and I_2621 (I50275,I50035,I50258);
DFFARX1 I_2622  ( .D(I50275), .CLK(I5694_clk), .RSTB(I49721_rst), .Q(I49713) );
or I_2623 (I50306,I50241,I50052);
DFFARX1 I_2624  ( .D(I50306), .CLK(I5694_clk), .RSTB(I49721_rst), .Q(I49698) );
nand I_2625 (I49701,I50241,I50131);
not I_2626 (I50384_rst,I5701);
not I_2627 (I50401,I19894);
nor I_2628 (I50418,I19891,I19909);
nand I_2629 (I50435,I50418,I19912);
nor I_2630 (I50452,I50401,I19891);
nand I_2631 (I50469,I50452,I19897);
not I_2632 (I50486,I50469);
not I_2633 (I50503,I19891);
nor I_2634 (I50373,I50469,I50503);
not I_2635 (I50534,I50503);
nand I_2636 (I50358,I50469,I50534);
not I_2637 (I50565,I19906);
nor I_2638 (I50582,I50565,I19888);
and I_2639 (I50599,I50582,I19882);
or I_2640 (I50616,I50599,I19900);
DFFARX1 I_2641  ( .D(I50616), .CLK(I5694_clk), .RSTB(I50384_rst), .Q(I50633) );
nor I_2642 (I50650,I50633,I50486);
DFFARX1 I_2643  ( .D(I50633), .CLK(I5694_clk), .RSTB(I50384_rst), .Q(I50667) );
not I_2644 (I50355,I50667);
nand I_2645 (I50698,I50401,I19906);
and I_2646 (I50715,I50698,I50650);
DFFARX1 I_2647  ( .D(I50698), .CLK(I5694_clk), .RSTB(I50384_rst), .Q(I50352) );
DFFARX1 I_2648  ( .D(I19885), .CLK(I5694_clk), .RSTB(I50384_rst), .Q(I50746) );
nor I_2649 (I50763,I50746,I50469);
nand I_2650 (I50370,I50633,I50763);
nor I_2651 (I50794,I50746,I50534);
not I_2652 (I50367,I50746);
nand I_2653 (I50825,I50746,I50435);
and I_2654 (I50842,I50503,I50825);
DFFARX1 I_2655  ( .D(I50842), .CLK(I5694_clk), .RSTB(I50384_rst), .Q(I50346) );
DFFARX1 I_2656  ( .D(I50746), .CLK(I5694_clk), .RSTB(I50384_rst), .Q(I50349) );
DFFARX1 I_2657  ( .D(I19903), .CLK(I5694_clk), .RSTB(I50384_rst), .Q(I50887) );
not I_2658 (I50904,I50887);
nand I_2659 (I50921,I50904,I50469);
and I_2660 (I50938,I50698,I50921);
DFFARX1 I_2661  ( .D(I50938), .CLK(I5694_clk), .RSTB(I50384_rst), .Q(I50376) );
or I_2662 (I50969,I50904,I50715);
DFFARX1 I_2663  ( .D(I50969), .CLK(I5694_clk), .RSTB(I50384_rst), .Q(I50361) );
nand I_2664 (I50364,I50904,I50794);
not I_2665 (I51047_rst,I5701);
not I_2666 (I51064,I36741);
nor I_2667 (I51081,I36732,I36738);
nand I_2668 (I51098,I51081,I36750);
nor I_2669 (I51115,I51064,I36732);
nand I_2670 (I51132,I51115,I36735);
not I_2671 (I51149,I51132);
not I_2672 (I51166,I36732);
nor I_2673 (I51036,I51132,I51166);
not I_2674 (I51197,I51166);
nand I_2675 (I51021,I51132,I51197);
not I_2676 (I51228,I36759);
nor I_2677 (I51245,I51228,I36753);
and I_2678 (I51262,I51245,I36744);
or I_2679 (I51279,I51262,I36729);
DFFARX1 I_2680  ( .D(I51279), .CLK(I5694_clk), .RSTB(I51047_rst), .Q(I51296) );
nor I_2681 (I51313,I51296,I51149);
DFFARX1 I_2682  ( .D(I51296), .CLK(I5694_clk), .RSTB(I51047_rst), .Q(I51330) );
not I_2683 (I51018,I51330);
nand I_2684 (I51361,I51064,I36759);
and I_2685 (I51378,I51361,I51313);
DFFARX1 I_2686  ( .D(I51361), .CLK(I5694_clk), .RSTB(I51047_rst), .Q(I51015) );
DFFARX1 I_2687  ( .D(I36747), .CLK(I5694_clk), .RSTB(I51047_rst), .Q(I51409) );
nor I_2688 (I51426,I51409,I51132);
nand I_2689 (I51033,I51296,I51426);
nor I_2690 (I51457,I51409,I51197);
not I_2691 (I51030,I51409);
nand I_2692 (I51488,I51409,I51098);
and I_2693 (I51505,I51166,I51488);
DFFARX1 I_2694  ( .D(I51505), .CLK(I5694_clk), .RSTB(I51047_rst), .Q(I51009) );
DFFARX1 I_2695  ( .D(I51409), .CLK(I5694_clk), .RSTB(I51047_rst), .Q(I51012) );
DFFARX1 I_2696  ( .D(I36756), .CLK(I5694_clk), .RSTB(I51047_rst), .Q(I51550) );
not I_2697 (I51567,I51550);
nand I_2698 (I51584,I51567,I51132);
and I_2699 (I51601,I51361,I51584);
DFFARX1 I_2700  ( .D(I51601), .CLK(I5694_clk), .RSTB(I51047_rst), .Q(I51039) );
or I_2701 (I51632,I51567,I51378);
DFFARX1 I_2702  ( .D(I51632), .CLK(I5694_clk), .RSTB(I51047_rst), .Q(I51024) );
nand I_2703 (I51027,I51567,I51457);
not I_2704 (I51710_rst,I5701);
not I_2705 (I51727,I43433);
nor I_2706 (I51744,I43430,I43454);
nand I_2707 (I51761,I51744,I43451);
nor I_2708 (I51778,I51727,I43430);
nand I_2709 (I51795,I51778,I43457);
not I_2710 (I51812,I51795);
not I_2711 (I51829,I43430);
nor I_2712 (I51699,I51795,I51829);
not I_2713 (I51860,I51829);
nand I_2714 (I51684,I51795,I51860);
not I_2715 (I51891,I43448);
nor I_2716 (I51908,I51891,I43439);
and I_2717 (I51925,I51908,I43436);
or I_2718 (I51942,I51925,I43445);
DFFARX1 I_2719  ( .D(I51942), .CLK(I5694_clk), .RSTB(I51710_rst), .Q(I51959) );
nor I_2720 (I51976,I51959,I51812);
DFFARX1 I_2721  ( .D(I51959), .CLK(I5694_clk), .RSTB(I51710_rst), .Q(I51993) );
not I_2722 (I51681,I51993);
nand I_2723 (I52024,I51727,I43448);
and I_2724 (I52041,I52024,I51976);
DFFARX1 I_2725  ( .D(I52024), .CLK(I5694_clk), .RSTB(I51710_rst), .Q(I51678) );
DFFARX1 I_2726  ( .D(I43427), .CLK(I5694_clk), .RSTB(I51710_rst), .Q(I52072) );
nor I_2727 (I52089,I52072,I51795);
nand I_2728 (I51696,I51959,I52089);
nor I_2729 (I52120,I52072,I51860);
not I_2730 (I51693,I52072);
nand I_2731 (I52151,I52072,I51761);
and I_2732 (I52168,I51829,I52151);
DFFARX1 I_2733  ( .D(I52168), .CLK(I5694_clk), .RSTB(I51710_rst), .Q(I51672) );
DFFARX1 I_2734  ( .D(I52072), .CLK(I5694_clk), .RSTB(I51710_rst), .Q(I51675) );
DFFARX1 I_2735  ( .D(I43442), .CLK(I5694_clk), .RSTB(I51710_rst), .Q(I52213) );
not I_2736 (I52230,I52213);
nand I_2737 (I52247,I52230,I51795);
and I_2738 (I52264,I52024,I52247);
DFFARX1 I_2739  ( .D(I52264), .CLK(I5694_clk), .RSTB(I51710_rst), .Q(I51702) );
or I_2740 (I52295,I52230,I52041);
DFFARX1 I_2741  ( .D(I52295), .CLK(I5694_clk), .RSTB(I51710_rst), .Q(I51687) );
nand I_2742 (I51690,I52230,I52120);
not I_2743 (I52373_rst,I5701);
not I_2744 (I52390,I18602);
nor I_2745 (I52407,I18599,I18617);
nand I_2746 (I52424,I52407,I18620);
nor I_2747 (I52441,I52390,I18599);
nand I_2748 (I52458,I52441,I18605);
not I_2749 (I52475,I52458);
not I_2750 (I52492,I18599);
nor I_2751 (I52362,I52458,I52492);
not I_2752 (I52523,I52492);
nand I_2753 (I52347,I52458,I52523);
not I_2754 (I52554,I18614);
nor I_2755 (I52571,I52554,I18596);
and I_2756 (I52588,I52571,I18590);
or I_2757 (I52605,I52588,I18608);
DFFARX1 I_2758  ( .D(I52605), .CLK(I5694_clk), .RSTB(I52373_rst), .Q(I52622) );
nor I_2759 (I52639,I52622,I52475);
DFFARX1 I_2760  ( .D(I52622), .CLK(I5694_clk), .RSTB(I52373_rst), .Q(I52656) );
not I_2761 (I52344,I52656);
nand I_2762 (I52687,I52390,I18614);
and I_2763 (I52704,I52687,I52639);
DFFARX1 I_2764  ( .D(I52687), .CLK(I5694_clk), .RSTB(I52373_rst), .Q(I52341) );
DFFARX1 I_2765  ( .D(I18593), .CLK(I5694_clk), .RSTB(I52373_rst), .Q(I52735) );
nor I_2766 (I52752,I52735,I52458);
nand I_2767 (I52359,I52622,I52752);
nor I_2768 (I52783,I52735,I52523);
not I_2769 (I52356,I52735);
nand I_2770 (I52814,I52735,I52424);
and I_2771 (I52831,I52492,I52814);
DFFARX1 I_2772  ( .D(I52831), .CLK(I5694_clk), .RSTB(I52373_rst), .Q(I52335) );
DFFARX1 I_2773  ( .D(I52735), .CLK(I5694_clk), .RSTB(I52373_rst), .Q(I52338) );
DFFARX1 I_2774  ( .D(I18611), .CLK(I5694_clk), .RSTB(I52373_rst), .Q(I52876) );
not I_2775 (I52893,I52876);
nand I_2776 (I52910,I52893,I52458);
and I_2777 (I52927,I52687,I52910);
DFFARX1 I_2778  ( .D(I52927), .CLK(I5694_clk), .RSTB(I52373_rst), .Q(I52365) );
or I_2779 (I52958,I52893,I52704);
DFFARX1 I_2780  ( .D(I52958), .CLK(I5694_clk), .RSTB(I52373_rst), .Q(I52350) );
nand I_2781 (I52353,I52893,I52783);
not I_2782 (I53036_rst,I5701);
not I_2783 (I53053,I27737);
nor I_2784 (I53070,I27746,I27728);
nand I_2785 (I53087,I53070,I27749);
nor I_2786 (I53104,I53053,I27746);
nand I_2787 (I53121,I53104,I27740);
not I_2788 (I53138,I53121);
not I_2789 (I53155,I27746);
nor I_2790 (I53025,I53121,I53155);
not I_2791 (I53186,I53155);
nand I_2792 (I53010,I53121,I53186);
not I_2793 (I53217,I27734);
nor I_2794 (I53234,I53217,I27725);
and I_2795 (I53251,I53234,I27722);
or I_2796 (I53268,I53251,I27719);
DFFARX1 I_2797  ( .D(I53268), .CLK(I5694_clk), .RSTB(I53036_rst), .Q(I53285) );
nor I_2798 (I53302,I53285,I53138);
DFFARX1 I_2799  ( .D(I53285), .CLK(I5694_clk), .RSTB(I53036_rst), .Q(I53319) );
not I_2800 (I53007,I53319);
nand I_2801 (I53350,I53053,I27734);
and I_2802 (I53367,I53350,I53302);
DFFARX1 I_2803  ( .D(I53350), .CLK(I5694_clk), .RSTB(I53036_rst), .Q(I53004) );
DFFARX1 I_2804  ( .D(I27743), .CLK(I5694_clk), .RSTB(I53036_rst), .Q(I53398) );
nor I_2805 (I53415,I53398,I53121);
nand I_2806 (I53022,I53285,I53415);
nor I_2807 (I53446,I53398,I53186);
not I_2808 (I53019,I53398);
nand I_2809 (I53477,I53398,I53087);
and I_2810 (I53494,I53155,I53477);
DFFARX1 I_2811  ( .D(I53494), .CLK(I5694_clk), .RSTB(I53036_rst), .Q(I52998) );
DFFARX1 I_2812  ( .D(I53398), .CLK(I5694_clk), .RSTB(I53036_rst), .Q(I53001) );
DFFARX1 I_2813  ( .D(I27731), .CLK(I5694_clk), .RSTB(I53036_rst), .Q(I53539) );
not I_2814 (I53556,I53539);
nand I_2815 (I53573,I53556,I53121);
and I_2816 (I53590,I53350,I53573);
DFFARX1 I_2817  ( .D(I53590), .CLK(I5694_clk), .RSTB(I53036_rst), .Q(I53028) );
or I_2818 (I53621,I53556,I53367);
DFFARX1 I_2819  ( .D(I53621), .CLK(I5694_clk), .RSTB(I53036_rst), .Q(I53013) );
nand I_2820 (I53016,I53556,I53446);
not I_2821 (I53699_rst,I5701);
not I_2822 (I53716,I42141);
nor I_2823 (I53733,I42138,I42162);
nand I_2824 (I53750,I53733,I42159);
nor I_2825 (I53767,I53716,I42138);
nand I_2826 (I53784,I53767,I42165);
not I_2827 (I53801,I53784);
not I_2828 (I53818,I42138);
nor I_2829 (I53688,I53784,I53818);
not I_2830 (I53849,I53818);
nand I_2831 (I53673,I53784,I53849);
not I_2832 (I53880,I42156);
nor I_2833 (I53897,I53880,I42147);
and I_2834 (I53914,I53897,I42144);
or I_2835 (I53931,I53914,I42153);
DFFARX1 I_2836  ( .D(I53931), .CLK(I5694_clk), .RSTB(I53699_rst), .Q(I53948) );
nor I_2837 (I53965,I53948,I53801);
DFFARX1 I_2838  ( .D(I53948), .CLK(I5694_clk), .RSTB(I53699_rst), .Q(I53982) );
not I_2839 (I53670,I53982);
nand I_2840 (I54013,I53716,I42156);
and I_2841 (I54030,I54013,I53965);
DFFARX1 I_2842  ( .D(I54013), .CLK(I5694_clk), .RSTB(I53699_rst), .Q(I53667) );
DFFARX1 I_2843  ( .D(I42135), .CLK(I5694_clk), .RSTB(I53699_rst), .Q(I54061) );
nor I_2844 (I54078,I54061,I53784);
nand I_2845 (I53685,I53948,I54078);
nor I_2846 (I54109,I54061,I53849);
not I_2847 (I53682,I54061);
nand I_2848 (I54140,I54061,I53750);
and I_2849 (I54157,I53818,I54140);
DFFARX1 I_2850  ( .D(I54157), .CLK(I5694_clk), .RSTB(I53699_rst), .Q(I53661) );
DFFARX1 I_2851  ( .D(I54061), .CLK(I5694_clk), .RSTB(I53699_rst), .Q(I53664) );
DFFARX1 I_2852  ( .D(I42150), .CLK(I5694_clk), .RSTB(I53699_rst), .Q(I54202) );
not I_2853 (I54219,I54202);
nand I_2854 (I54236,I54219,I53784);
and I_2855 (I54253,I54013,I54236);
DFFARX1 I_2856  ( .D(I54253), .CLK(I5694_clk), .RSTB(I53699_rst), .Q(I53691) );
or I_2857 (I54284,I54219,I54030);
DFFARX1 I_2858  ( .D(I54284), .CLK(I5694_clk), .RSTB(I53699_rst), .Q(I53676) );
nand I_2859 (I53679,I54219,I54109);
not I_2860 (I54362_rst,I5701);
not I_2861 (I54379,I6283);
nor I_2862 (I54396,I6289,I6292);
nand I_2863 (I54413,I54396,I6268);
nor I_2864 (I54430,I54379,I6289);
nand I_2865 (I54447,I54430,I6277);
not I_2866 (I54464,I54447);
not I_2867 (I54481,I6289);
nor I_2868 (I54351,I54447,I54481);
not I_2869 (I54512,I54481);
nand I_2870 (I54336,I54447,I54512);
not I_2871 (I54543,I6271);
nor I_2872 (I54560,I54543,I6295);
and I_2873 (I54577,I54560,I6265);
or I_2874 (I54594,I54577,I6274);
DFFARX1 I_2875  ( .D(I54594), .CLK(I5694_clk), .RSTB(I54362_rst), .Q(I54611) );
nor I_2876 (I54628,I54611,I54464);
DFFARX1 I_2877  ( .D(I54611), .CLK(I5694_clk), .RSTB(I54362_rst), .Q(I54645) );
not I_2878 (I54333,I54645);
nand I_2879 (I54676,I54379,I6271);
and I_2880 (I54693,I54676,I54628);
DFFARX1 I_2881  ( .D(I54676), .CLK(I5694_clk), .RSTB(I54362_rst), .Q(I54330) );
DFFARX1 I_2882  ( .D(I6280), .CLK(I5694_clk), .RSTB(I54362_rst), .Q(I54724) );
nor I_2883 (I54741,I54724,I54447);
nand I_2884 (I54348,I54611,I54741);
nor I_2885 (I54772,I54724,I54512);
not I_2886 (I54345,I54724);
nand I_2887 (I54803,I54724,I54413);
and I_2888 (I54820,I54481,I54803);
DFFARX1 I_2889  ( .D(I54820), .CLK(I5694_clk), .RSTB(I54362_rst), .Q(I54324) );
DFFARX1 I_2890  ( .D(I54724), .CLK(I5694_clk), .RSTB(I54362_rst), .Q(I54327) );
DFFARX1 I_2891  ( .D(I6286), .CLK(I5694_clk), .RSTB(I54362_rst), .Q(I54865) );
not I_2892 (I54882,I54865);
nand I_2893 (I54899,I54882,I54447);
and I_2894 (I54916,I54676,I54899);
DFFARX1 I_2895  ( .D(I54916), .CLK(I5694_clk), .RSTB(I54362_rst), .Q(I54354) );
or I_2896 (I54947,I54882,I54693);
DFFARX1 I_2897  ( .D(I54947), .CLK(I5694_clk), .RSTB(I54362_rst), .Q(I54339) );
nand I_2898 (I54342,I54882,I54772);
not I_2899 (I55025_rst,I5701);
not I_2900 (I55042,I45385);
nor I_2901 (I55059,I45391,I45397);
nand I_2902 (I55076,I55059,I45400);
nor I_2903 (I55093,I55042,I45391);
nand I_2904 (I55110,I55093,I45382);
not I_2905 (I55127,I55110);
not I_2906 (I55144,I45391);
nor I_2907 (I55014,I55110,I55144);
not I_2908 (I55175,I55144);
nand I_2909 (I54999,I55110,I55175);
not I_2910 (I55206,I45394);
nor I_2911 (I55223,I55206,I45388);
and I_2912 (I55240,I55223,I45403);
or I_2913 (I55257,I55240,I45409);
DFFARX1 I_2914  ( .D(I55257), .CLK(I5694_clk), .RSTB(I55025_rst), .Q(I55274) );
nor I_2915 (I55291,I55274,I55127);
DFFARX1 I_2916  ( .D(I55274), .CLK(I5694_clk), .RSTB(I55025_rst), .Q(I55308) );
not I_2917 (I54996,I55308);
nand I_2918 (I55339,I55042,I45394);
and I_2919 (I55356,I55339,I55291);
DFFARX1 I_2920  ( .D(I55339), .CLK(I5694_clk), .RSTB(I55025_rst), .Q(I54993) );
DFFARX1 I_2921  ( .D(I45406), .CLK(I5694_clk), .RSTB(I55025_rst), .Q(I55387) );
nor I_2922 (I55404,I55387,I55110);
nand I_2923 (I55011,I55274,I55404);
nor I_2924 (I55435,I55387,I55175);
not I_2925 (I55008,I55387);
nand I_2926 (I55466,I55387,I55076);
and I_2927 (I55483,I55144,I55466);
DFFARX1 I_2928  ( .D(I55483), .CLK(I5694_clk), .RSTB(I55025_rst), .Q(I54987) );
DFFARX1 I_2929  ( .D(I55387), .CLK(I5694_clk), .RSTB(I55025_rst), .Q(I54990) );
DFFARX1 I_2930  ( .D(I45412), .CLK(I5694_clk), .RSTB(I55025_rst), .Q(I55528) );
not I_2931 (I55545,I55528);
nand I_2932 (I55562,I55545,I55110);
and I_2933 (I55579,I55339,I55562);
DFFARX1 I_2934  ( .D(I55579), .CLK(I5694_clk), .RSTB(I55025_rst), .Q(I55017) );
or I_2935 (I55610,I55545,I55356);
DFFARX1 I_2936  ( .D(I55610), .CLK(I5694_clk), .RSTB(I55025_rst), .Q(I55002) );
nand I_2937 (I55005,I55545,I55435);
not I_2938 (I55688_rst,I5701);
not I_2939 (I55705,I35585);
nor I_2940 (I55722,I35576,I35582);
nand I_2941 (I55739,I55722,I35594);
nor I_2942 (I55756,I55705,I35576);
nand I_2943 (I55773,I55756,I35579);
not I_2944 (I55790,I55773);
not I_2945 (I55807,I35576);
nor I_2946 (I55677,I55773,I55807);
not I_2947 (I55838,I55807);
nand I_2948 (I55662,I55773,I55838);
not I_2949 (I55869,I35603);
nor I_2950 (I55886,I55869,I35597);
and I_2951 (I55903,I55886,I35588);
or I_2952 (I55920,I55903,I35573);
DFFARX1 I_2953  ( .D(I55920), .CLK(I5694_clk), .RSTB(I55688_rst), .Q(I55937) );
nor I_2954 (I55954,I55937,I55790);
DFFARX1 I_2955  ( .D(I55937), .CLK(I5694_clk), .RSTB(I55688_rst), .Q(I55971) );
not I_2956 (I55659,I55971);
nand I_2957 (I56002,I55705,I35603);
and I_2958 (I56019,I56002,I55954);
DFFARX1 I_2959  ( .D(I56002), .CLK(I5694_clk), .RSTB(I55688_rst), .Q(I55656) );
DFFARX1 I_2960  ( .D(I35591), .CLK(I5694_clk), .RSTB(I55688_rst), .Q(I56050) );
nor I_2961 (I56067,I56050,I55773);
nand I_2962 (I55674,I55937,I56067);
nor I_2963 (I56098,I56050,I55838);
not I_2964 (I55671,I56050);
nand I_2965 (I56129,I56050,I55739);
and I_2966 (I56146,I55807,I56129);
DFFARX1 I_2967  ( .D(I56146), .CLK(I5694_clk), .RSTB(I55688_rst), .Q(I55650) );
DFFARX1 I_2968  ( .D(I56050), .CLK(I5694_clk), .RSTB(I55688_rst), .Q(I55653) );
DFFARX1 I_2969  ( .D(I35600), .CLK(I5694_clk), .RSTB(I55688_rst), .Q(I56191) );
not I_2970 (I56208,I56191);
nand I_2971 (I56225,I56208,I55773);
and I_2972 (I56242,I56002,I56225);
DFFARX1 I_2973  ( .D(I56242), .CLK(I5694_clk), .RSTB(I55688_rst), .Q(I55680) );
or I_2974 (I56273,I56208,I56019);
DFFARX1 I_2975  ( .D(I56273), .CLK(I5694_clk), .RSTB(I55688_rst), .Q(I55665) );
nand I_2976 (I55668,I56208,I56098);
not I_2977 (I56351_rst,I5701);
not I_2978 (I56368,I31973);
nor I_2979 (I56385,I31970,I31955);
nand I_2980 (I56402,I56385,I31964);
nor I_2981 (I56419,I56368,I31970);
nand I_2982 (I56436,I56419,I31979);
DFFARX1 I_2983  ( .D(I56436), .CLK(I5694_clk), .RSTB(I56351_rst), .Q(I56453) );
not I_2984 (I56322,I56453);
not I_2985 (I56484,I31970);
not I_2986 (I56501,I56484);
not I_2987 (I56518,I31952);
nor I_2988 (I56535,I56518,I31958);
and I_2989 (I56552,I56535,I31982);
or I_2990 (I56569,I56552,I31976);
DFFARX1 I_2991  ( .D(I56569), .CLK(I5694_clk), .RSTB(I56351_rst), .Q(I56586) );
DFFARX1 I_2992  ( .D(I56586), .CLK(I5694_clk), .RSTB(I56351_rst), .Q(I56319) );
DFFARX1 I_2993  ( .D(I56586), .CLK(I5694_clk), .RSTB(I56351_rst), .Q(I56617) );
DFFARX1 I_2994  ( .D(I56586), .CLK(I5694_clk), .RSTB(I56351_rst), .Q(I56313) );
nand I_2995 (I56648,I56368,I31952);
nand I_2996 (I56665,I56648,I56402);
and I_2997 (I56682,I56484,I56665);
DFFARX1 I_2998  ( .D(I56682), .CLK(I5694_clk), .RSTB(I56351_rst), .Q(I56343) );
and I_2999 (I56316,I56648,I56617);
DFFARX1 I_3000  ( .D(I31961), .CLK(I5694_clk), .RSTB(I56351_rst), .Q(I56727) );
nor I_3001 (I56340,I56727,I56648);
nor I_3002 (I56758,I56727,I56402);
nand I_3003 (I56337,I56436,I56758);
not I_3004 (I56334,I56727);
DFFARX1 I_3005  ( .D(I31967), .CLK(I5694_clk), .RSTB(I56351_rst), .Q(I56803) );
not I_3006 (I56820,I56803);
nor I_3007 (I56837,I56820,I56501);
and I_3008 (I56854,I56727,I56837);
or I_3009 (I56871,I56648,I56854);
DFFARX1 I_3010  ( .D(I56871), .CLK(I5694_clk), .RSTB(I56351_rst), .Q(I56328) );
not I_3011 (I56902,I56820);
nor I_3012 (I56919,I56727,I56902);
nand I_3013 (I56331,I56820,I56919);
nand I_3014 (I56325,I56484,I56902);
not I_3015 (I56997_rst,I5701);
not I_3016 (I57014,I8801);
nor I_3017 (I57031,I8822,I8804);
nand I_3018 (I57048,I57031,I8828);
nor I_3019 (I57065,I57014,I8822);
nand I_3020 (I57082,I57065,I8825);
DFFARX1 I_3021  ( .D(I57082), .CLK(I5694_clk), .RSTB(I56997_rst), .Q(I57099) );
not I_3022 (I56968,I57099);
not I_3023 (I57130,I8822);
not I_3024 (I57147,I57130);
not I_3025 (I57164,I8819);
nor I_3026 (I57181,I57164,I8798);
and I_3027 (I57198,I57181,I8810);
or I_3028 (I57215,I57198,I8807);
DFFARX1 I_3029  ( .D(I57215), .CLK(I5694_clk), .RSTB(I56997_rst), .Q(I57232) );
DFFARX1 I_3030  ( .D(I57232), .CLK(I5694_clk), .RSTB(I56997_rst), .Q(I56965) );
DFFARX1 I_3031  ( .D(I57232), .CLK(I5694_clk), .RSTB(I56997_rst), .Q(I57263) );
DFFARX1 I_3032  ( .D(I57232), .CLK(I5694_clk), .RSTB(I56997_rst), .Q(I56959) );
nand I_3033 (I57294,I57014,I8819);
nand I_3034 (I57311,I57294,I57048);
and I_3035 (I57328,I57130,I57311);
DFFARX1 I_3036  ( .D(I57328), .CLK(I5694_clk), .RSTB(I56997_rst), .Q(I56989) );
and I_3037 (I56962,I57294,I57263);
DFFARX1 I_3038  ( .D(I8813), .CLK(I5694_clk), .RSTB(I56997_rst), .Q(I57373) );
nor I_3039 (I56986,I57373,I57294);
nor I_3040 (I57404,I57373,I57048);
nand I_3041 (I56983,I57082,I57404);
not I_3042 (I56980,I57373);
DFFARX1 I_3043  ( .D(I8816), .CLK(I5694_clk), .RSTB(I56997_rst), .Q(I57449) );
not I_3044 (I57466,I57449);
nor I_3045 (I57483,I57466,I57147);
and I_3046 (I57500,I57373,I57483);
or I_3047 (I57517,I57294,I57500);
DFFARX1 I_3048  ( .D(I57517), .CLK(I5694_clk), .RSTB(I56997_rst), .Q(I56974) );
not I_3049 (I57548,I57466);
nor I_3050 (I57565,I57373,I57548);
nand I_3051 (I56977,I57466,I57565);
nand I_3052 (I56971,I57130,I57548);
not I_3053 (I57643_rst,I5701);
not I_3054 (I57660,I53022);
nor I_3055 (I57677,I53001,I53013);
nand I_3056 (I57694,I57677,I53016);
nor I_3057 (I57711,I57660,I53001);
nand I_3058 (I57728,I57711,I52998);
DFFARX1 I_3059  ( .D(I57728), .CLK(I5694_clk), .RSTB(I57643_rst), .Q(I57745) );
not I_3060 (I57614,I57745);
not I_3061 (I57776,I53001);
not I_3062 (I57793,I57776);
not I_3063 (I57810,I53019);
nor I_3064 (I57827,I57810,I53010);
and I_3065 (I57844,I57827,I53004);
or I_3066 (I57861,I57844,I53028);
DFFARX1 I_3067  ( .D(I57861), .CLK(I5694_clk), .RSTB(I57643_rst), .Q(I57878) );
DFFARX1 I_3068  ( .D(I57878), .CLK(I5694_clk), .RSTB(I57643_rst), .Q(I57611) );
DFFARX1 I_3069  ( .D(I57878), .CLK(I5694_clk), .RSTB(I57643_rst), .Q(I57909) );
DFFARX1 I_3070  ( .D(I57878), .CLK(I5694_clk), .RSTB(I57643_rst), .Q(I57605) );
nand I_3071 (I57940,I57660,I53019);
nand I_3072 (I57957,I57940,I57694);
and I_3073 (I57974,I57776,I57957);
DFFARX1 I_3074  ( .D(I57974), .CLK(I5694_clk), .RSTB(I57643_rst), .Q(I57635) );
and I_3075 (I57608,I57940,I57909);
DFFARX1 I_3076  ( .D(I53025), .CLK(I5694_clk), .RSTB(I57643_rst), .Q(I58019) );
nor I_3077 (I57632,I58019,I57940);
nor I_3078 (I58050,I58019,I57694);
nand I_3079 (I57629,I57728,I58050);
not I_3080 (I57626,I58019);
DFFARX1 I_3081  ( .D(I53007), .CLK(I5694_clk), .RSTB(I57643_rst), .Q(I58095) );
not I_3082 (I58112,I58095);
nor I_3083 (I58129,I58112,I57793);
and I_3084 (I58146,I58019,I58129);
or I_3085 (I58163,I57940,I58146);
DFFARX1 I_3086  ( .D(I58163), .CLK(I5694_clk), .RSTB(I57643_rst), .Q(I57620) );
not I_3087 (I58194,I58112);
nor I_3088 (I58211,I58019,I58194);
nand I_3089 (I57623,I58112,I58211);
nand I_3090 (I57617,I57776,I58194);
not I_3091 (I58289_rst,I5701);
not I_3092 (I58306,I11456);
nor I_3093 (I58323,I11462,I11459);
nand I_3094 (I58340,I58323,I11453);
nor I_3095 (I58357,I58306,I11462);
nand I_3096 (I58374,I58357,I11477);
DFFARX1 I_3097  ( .D(I58374), .CLK(I5694_clk), .RSTB(I58289_rst), .Q(I58391) );
not I_3098 (I58260,I58391);
not I_3099 (I58422,I11462);
not I_3100 (I58439,I58422);
not I_3101 (I58456,I11474);
nor I_3102 (I58473,I58456,I11465);
and I_3103 (I58490,I58473,I11450);
or I_3104 (I58507,I58490,I11471);
DFFARX1 I_3105  ( .D(I58507), .CLK(I5694_clk), .RSTB(I58289_rst), .Q(I58524) );
DFFARX1 I_3106  ( .D(I58524), .CLK(I5694_clk), .RSTB(I58289_rst), .Q(I58257) );
DFFARX1 I_3107  ( .D(I58524), .CLK(I5694_clk), .RSTB(I58289_rst), .Q(I58555) );
DFFARX1 I_3108  ( .D(I58524), .CLK(I5694_clk), .RSTB(I58289_rst), .Q(I58251) );
nand I_3109 (I58586,I58306,I11474);
nand I_3110 (I58603,I58586,I58340);
and I_3111 (I58620,I58422,I58603);
DFFARX1 I_3112  ( .D(I58620), .CLK(I5694_clk), .RSTB(I58289_rst), .Q(I58281) );
and I_3113 (I58254,I58586,I58555);
DFFARX1 I_3114  ( .D(I11468), .CLK(I5694_clk), .RSTB(I58289_rst), .Q(I58665) );
nor I_3115 (I58278,I58665,I58586);
nor I_3116 (I58696,I58665,I58340);
nand I_3117 (I58275,I58374,I58696);
not I_3118 (I58272,I58665);
DFFARX1 I_3119  ( .D(I11480), .CLK(I5694_clk), .RSTB(I58289_rst), .Q(I58741) );
not I_3120 (I58758,I58741);
nor I_3121 (I58775,I58758,I58439);
and I_3122 (I58792,I58665,I58775);
or I_3123 (I58809,I58586,I58792);
DFFARX1 I_3124  ( .D(I58809), .CLK(I5694_clk), .RSTB(I58289_rst), .Q(I58266) );
not I_3125 (I58840,I58758);
nor I_3126 (I58857,I58665,I58840);
nand I_3127 (I58269,I58758,I58857);
nand I_3128 (I58263,I58422,I58840);
not I_3129 (I58935_rst,I5701);
not I_3130 (I58952,I36169);
nor I_3131 (I58969,I36154,I36160);
nand I_3132 (I58986,I58969,I36157);
nor I_3133 (I59003,I58952,I36154);
nand I_3134 (I59020,I59003,I36166);
DFFARX1 I_3135  ( .D(I59020), .CLK(I5694_clk), .RSTB(I58935_rst), .Q(I59037) );
not I_3136 (I58906,I59037);
not I_3137 (I59068,I36154);
not I_3138 (I59085,I59068);
not I_3139 (I59102,I36181);
nor I_3140 (I59119,I59102,I36175);
and I_3141 (I59136,I59119,I36172);
or I_3142 (I59153,I59136,I36151);
DFFARX1 I_3143  ( .D(I59153), .CLK(I5694_clk), .RSTB(I58935_rst), .Q(I59170) );
DFFARX1 I_3144  ( .D(I59170), .CLK(I5694_clk), .RSTB(I58935_rst), .Q(I58903) );
DFFARX1 I_3145  ( .D(I59170), .CLK(I5694_clk), .RSTB(I58935_rst), .Q(I59201) );
DFFARX1 I_3146  ( .D(I59170), .CLK(I5694_clk), .RSTB(I58935_rst), .Q(I58897) );
nand I_3147 (I59232,I58952,I36181);
nand I_3148 (I59249,I59232,I58986);
and I_3149 (I59266,I59068,I59249);
DFFARX1 I_3150  ( .D(I59266), .CLK(I5694_clk), .RSTB(I58935_rst), .Q(I58927) );
and I_3151 (I58900,I59232,I59201);
DFFARX1 I_3152  ( .D(I36178), .CLK(I5694_clk), .RSTB(I58935_rst), .Q(I59311) );
nor I_3153 (I58924,I59311,I59232);
nor I_3154 (I59342,I59311,I58986);
nand I_3155 (I58921,I59020,I59342);
not I_3156 (I58918,I59311);
DFFARX1 I_3157  ( .D(I36163), .CLK(I5694_clk), .RSTB(I58935_rst), .Q(I59387) );
not I_3158 (I59404,I59387);
nor I_3159 (I59421,I59404,I59085);
and I_3160 (I59438,I59311,I59421);
or I_3161 (I59455,I59232,I59438);
DFFARX1 I_3162  ( .D(I59455), .CLK(I5694_clk), .RSTB(I58935_rst), .Q(I58912) );
not I_3163 (I59486,I59404);
nor I_3164 (I59503,I59311,I59486);
nand I_3165 (I58915,I59404,I59503);
nand I_3166 (I58909,I59068,I59486);
not I_3167 (I59581_rst,I5701);
not I_3168 (I59598,I13990);
nor I_3169 (I59615,I13969,I13981);
nand I_3170 (I59632,I59615,I13984);
nor I_3171 (I59649,I59598,I13969);
nand I_3172 (I59666,I59649,I13966);
DFFARX1 I_3173  ( .D(I59666), .CLK(I5694_clk), .RSTB(I59581_rst), .Q(I59683) );
not I_3174 (I59552,I59683);
not I_3175 (I59714,I13969);
not I_3176 (I59731,I59714);
not I_3177 (I59748,I13987);
nor I_3178 (I59765,I59748,I13978);
and I_3179 (I59782,I59765,I13972);
or I_3180 (I59799,I59782,I13996);
DFFARX1 I_3181  ( .D(I59799), .CLK(I5694_clk), .RSTB(I59581_rst), .Q(I59816) );
DFFARX1 I_3182  ( .D(I59816), .CLK(I5694_clk), .RSTB(I59581_rst), .Q(I59549) );
DFFARX1 I_3183  ( .D(I59816), .CLK(I5694_clk), .RSTB(I59581_rst), .Q(I59847) );
DFFARX1 I_3184  ( .D(I59816), .CLK(I5694_clk), .RSTB(I59581_rst), .Q(I59543) );
nand I_3185 (I59878,I59598,I13987);
nand I_3186 (I59895,I59878,I59632);
and I_3187 (I59912,I59714,I59895);
DFFARX1 I_3188  ( .D(I59912), .CLK(I5694_clk), .RSTB(I59581_rst), .Q(I59573) );
and I_3189 (I59546,I59878,I59847);
DFFARX1 I_3190  ( .D(I13993), .CLK(I5694_clk), .RSTB(I59581_rst), .Q(I59957) );
nor I_3191 (I59570,I59957,I59878);
nor I_3192 (I59988,I59957,I59632);
nand I_3193 (I59567,I59666,I59988);
not I_3194 (I59564,I59957);
DFFARX1 I_3195  ( .D(I13975), .CLK(I5694_clk), .RSTB(I59581_rst), .Q(I60033) );
not I_3196 (I60050,I60033);
nor I_3197 (I60067,I60050,I59731);
and I_3198 (I60084,I59957,I60067);
or I_3199 (I60101,I59878,I60084);
DFFARX1 I_3200  ( .D(I60101), .CLK(I5694_clk), .RSTB(I59581_rst), .Q(I59558) );
not I_3201 (I60132,I60050);
nor I_3202 (I60149,I59957,I60132);
nand I_3203 (I59561,I60050,I60149);
nand I_3204 (I59555,I59714,I60132);
not I_3205 (I60227_rst,I5701);
not I_3206 (I60244,I49103);
nor I_3207 (I60261,I49091,I49094);
nand I_3208 (I60278,I60261,I49118);
nor I_3209 (I60295,I60244,I49091);
nand I_3210 (I60312,I60295,I49100);
DFFARX1 I_3211  ( .D(I60312), .CLK(I5694_clk), .RSTB(I60227_rst), .Q(I60329) );
not I_3212 (I60198,I60329);
not I_3213 (I60360,I49091);
not I_3214 (I60377,I60360);
not I_3215 (I60394,I49097);
nor I_3216 (I60411,I60394,I49112);
and I_3217 (I60428,I60411,I49088);
or I_3218 (I60445,I60428,I49115);
DFFARX1 I_3219  ( .D(I60445), .CLK(I5694_clk), .RSTB(I60227_rst), .Q(I60462) );
DFFARX1 I_3220  ( .D(I60462), .CLK(I5694_clk), .RSTB(I60227_rst), .Q(I60195) );
DFFARX1 I_3221  ( .D(I60462), .CLK(I5694_clk), .RSTB(I60227_rst), .Q(I60493) );
DFFARX1 I_3222  ( .D(I60462), .CLK(I5694_clk), .RSTB(I60227_rst), .Q(I60189) );
nand I_3223 (I60524,I60244,I49097);
nand I_3224 (I60541,I60524,I60278);
and I_3225 (I60558,I60360,I60541);
DFFARX1 I_3226  ( .D(I60558), .CLK(I5694_clk), .RSTB(I60227_rst), .Q(I60219) );
and I_3227 (I60192,I60524,I60493);
DFFARX1 I_3228  ( .D(I49106), .CLK(I5694_clk), .RSTB(I60227_rst), .Q(I60603) );
nor I_3229 (I60216,I60603,I60524);
nor I_3230 (I60634,I60603,I60278);
nand I_3231 (I60213,I60312,I60634);
not I_3232 (I60210,I60603);
DFFARX1 I_3233  ( .D(I49109), .CLK(I5694_clk), .RSTB(I60227_rst), .Q(I60679) );
not I_3234 (I60696,I60679);
nor I_3235 (I60713,I60696,I60377);
and I_3236 (I60730,I60603,I60713);
or I_3237 (I60747,I60524,I60730);
DFFARX1 I_3238  ( .D(I60747), .CLK(I5694_clk), .RSTB(I60227_rst), .Q(I60204) );
not I_3239 (I60778,I60696);
nor I_3240 (I60795,I60603,I60778);
nand I_3241 (I60207,I60696,I60795);
nand I_3242 (I60201,I60360,I60778);
not I_3243 (I60873_rst,I5701);
not I_3244 (I60890,I41510);
nor I_3245 (I60907,I41501,I41492);
nand I_3246 (I60924,I60907,I41507);
nor I_3247 (I60941,I60890,I41501);
nand I_3248 (I60958,I60941,I41504);
DFFARX1 I_3249  ( .D(I60958), .CLK(I5694_clk), .RSTB(I60873_rst), .Q(I60975) );
not I_3250 (I60844,I60975);
not I_3251 (I61006,I41501);
not I_3252 (I61023,I61006);
not I_3253 (I61040,I41513);
nor I_3254 (I61057,I61040,I41498);
and I_3255 (I61074,I61057,I41516);
or I_3256 (I61091,I61074,I41489);
DFFARX1 I_3257  ( .D(I61091), .CLK(I5694_clk), .RSTB(I60873_rst), .Q(I61108) );
DFFARX1 I_3258  ( .D(I61108), .CLK(I5694_clk), .RSTB(I60873_rst), .Q(I60841) );
DFFARX1 I_3259  ( .D(I61108), .CLK(I5694_clk), .RSTB(I60873_rst), .Q(I61139) );
DFFARX1 I_3260  ( .D(I61108), .CLK(I5694_clk), .RSTB(I60873_rst), .Q(I60835) );
nand I_3261 (I61170,I60890,I41513);
nand I_3262 (I61187,I61170,I60924);
and I_3263 (I61204,I61006,I61187);
DFFARX1 I_3264  ( .D(I61204), .CLK(I5694_clk), .RSTB(I60873_rst), .Q(I60865) );
and I_3265 (I60838,I61170,I61139);
DFFARX1 I_3266  ( .D(I41519), .CLK(I5694_clk), .RSTB(I60873_rst), .Q(I61249) );
nor I_3267 (I60862,I61249,I61170);
nor I_3268 (I61280,I61249,I60924);
nand I_3269 (I60859,I60958,I61280);
not I_3270 (I60856,I61249);
DFFARX1 I_3271  ( .D(I41495), .CLK(I5694_clk), .RSTB(I60873_rst), .Q(I61325) );
not I_3272 (I61342,I61325);
nor I_3273 (I61359,I61342,I61023);
and I_3274 (I61376,I61249,I61359);
or I_3275 (I61393,I61170,I61376);
DFFARX1 I_3276  ( .D(I61393), .CLK(I5694_clk), .RSTB(I60873_rst), .Q(I60850) );
not I_3277 (I61424,I61342);
nor I_3278 (I61441,I61249,I61424);
nand I_3279 (I60853,I61342,I61441);
nand I_3280 (I60847,I61006,I61424);
not I_3281 (I61519_rst,I5701);
not I_3282 (I61536,I49707);
nor I_3283 (I61553,I49686,I49698);
nand I_3284 (I61570,I61553,I49701);
nor I_3285 (I61587,I61536,I49686);
nand I_3286 (I61604,I61587,I49683);
DFFARX1 I_3287  ( .D(I61604), .CLK(I5694_clk), .RSTB(I61519_rst), .Q(I61621) );
not I_3288 (I61490,I61621);
not I_3289 (I61652,I49686);
not I_3290 (I61669,I61652);
not I_3291 (I61686,I49704);
nor I_3292 (I61703,I61686,I49695);
and I_3293 (I61720,I61703,I49689);
or I_3294 (I61737,I61720,I49713);
DFFARX1 I_3295  ( .D(I61737), .CLK(I5694_clk), .RSTB(I61519_rst), .Q(I61754) );
DFFARX1 I_3296  ( .D(I61754), .CLK(I5694_clk), .RSTB(I61519_rst), .Q(I61487) );
DFFARX1 I_3297  ( .D(I61754), .CLK(I5694_clk), .RSTB(I61519_rst), .Q(I61785) );
DFFARX1 I_3298  ( .D(I61754), .CLK(I5694_clk), .RSTB(I61519_rst), .Q(I61481) );
nand I_3299 (I61816,I61536,I49704);
nand I_3300 (I61833,I61816,I61570);
and I_3301 (I61850,I61652,I61833);
DFFARX1 I_3302  ( .D(I61850), .CLK(I5694_clk), .RSTB(I61519_rst), .Q(I61511) );
and I_3303 (I61484,I61816,I61785);
DFFARX1 I_3304  ( .D(I49710), .CLK(I5694_clk), .RSTB(I61519_rst), .Q(I61895) );
nor I_3305 (I61508,I61895,I61816);
nor I_3306 (I61926,I61895,I61570);
nand I_3307 (I61505,I61604,I61926);
not I_3308 (I61502,I61895);
DFFARX1 I_3309  ( .D(I49692), .CLK(I5694_clk), .RSTB(I61519_rst), .Q(I61971) );
not I_3310 (I61988,I61971);
nor I_3311 (I62005,I61988,I61669);
and I_3312 (I62022,I61895,I62005);
or I_3313 (I62039,I61816,I62022);
DFFARX1 I_3314  ( .D(I62039), .CLK(I5694_clk), .RSTB(I61519_rst), .Q(I61496) );
not I_3315 (I62070,I61988);
nor I_3316 (I62087,I61895,I62070);
nand I_3317 (I61499,I61988,I62087);
nand I_3318 (I61493,I61652,I62070);
not I_3319 (I62165_rst,I5701);
not I_3320 (I62182,I10127);
nor I_3321 (I62199,I10148,I10130);
nand I_3322 (I62216,I62199,I10154);
nor I_3323 (I62233,I62182,I10148);
nand I_3324 (I62250,I62233,I10151);
DFFARX1 I_3325  ( .D(I62250), .CLK(I5694_clk), .RSTB(I62165_rst), .Q(I62267) );
not I_3326 (I62136,I62267);
not I_3327 (I62298,I10148);
not I_3328 (I62315,I62298);
not I_3329 (I62332,I10145);
nor I_3330 (I62349,I62332,I10124);
and I_3331 (I62366,I62349,I10136);
or I_3332 (I62383,I62366,I10133);
DFFARX1 I_3333  ( .D(I62383), .CLK(I5694_clk), .RSTB(I62165_rst), .Q(I62400) );
DFFARX1 I_3334  ( .D(I62400), .CLK(I5694_clk), .RSTB(I62165_rst), .Q(I62133) );
DFFARX1 I_3335  ( .D(I62400), .CLK(I5694_clk), .RSTB(I62165_rst), .Q(I62431) );
DFFARX1 I_3336  ( .D(I62400), .CLK(I5694_clk), .RSTB(I62165_rst), .Q(I62127) );
nand I_3337 (I62462,I62182,I10145);
nand I_3338 (I62479,I62462,I62216);
and I_3339 (I62496,I62298,I62479);
DFFARX1 I_3340  ( .D(I62496), .CLK(I5694_clk), .RSTB(I62165_rst), .Q(I62157) );
and I_3341 (I62130,I62462,I62431);
DFFARX1 I_3342  ( .D(I10139), .CLK(I5694_clk), .RSTB(I62165_rst), .Q(I62541) );
nor I_3343 (I62154,I62541,I62462);
nor I_3344 (I62572,I62541,I62216);
nand I_3345 (I62151,I62250,I62572);
not I_3346 (I62148,I62541);
DFFARX1 I_3347  ( .D(I10142), .CLK(I5694_clk), .RSTB(I62165_rst), .Q(I62617) );
not I_3348 (I62634,I62617);
nor I_3349 (I62651,I62634,I62315);
and I_3350 (I62668,I62541,I62651);
or I_3351 (I62685,I62462,I62668);
DFFARX1 I_3352  ( .D(I62685), .CLK(I5694_clk), .RSTB(I62165_rst), .Q(I62142) );
not I_3353 (I62716,I62634);
nor I_3354 (I62733,I62541,I62716);
nand I_3355 (I62145,I62634,I62733);
nand I_3356 (I62139,I62298,I62716);
not I_3357 (I62811_rst,I5701);
not I_3358 (I62828,I8138);
nor I_3359 (I62845,I8159,I8141);
nand I_3360 (I62862,I62845,I8165);
nor I_3361 (I62879,I62828,I8159);
nand I_3362 (I62896,I62879,I8162);
DFFARX1 I_3363  ( .D(I62896), .CLK(I5694_clk), .RSTB(I62811_rst), .Q(I62913) );
not I_3364 (I62782,I62913);
not I_3365 (I62944,I8159);
not I_3366 (I62961,I62944);
not I_3367 (I62978,I8156);
nor I_3368 (I62995,I62978,I8135);
and I_3369 (I63012,I62995,I8147);
or I_3370 (I63029,I63012,I8144);
DFFARX1 I_3371  ( .D(I63029), .CLK(I5694_clk), .RSTB(I62811_rst), .Q(I63046) );
DFFARX1 I_3372  ( .D(I63046), .CLK(I5694_clk), .RSTB(I62811_rst), .Q(I62779) );
DFFARX1 I_3373  ( .D(I63046), .CLK(I5694_clk), .RSTB(I62811_rst), .Q(I63077) );
DFFARX1 I_3374  ( .D(I63046), .CLK(I5694_clk), .RSTB(I62811_rst), .Q(I62773) );
nand I_3375 (I63108,I62828,I8156);
nand I_3376 (I63125,I63108,I62862);
and I_3377 (I63142,I62944,I63125);
DFFARX1 I_3378  ( .D(I63142), .CLK(I5694_clk), .RSTB(I62811_rst), .Q(I62803) );
and I_3379 (I62776,I63108,I63077);
DFFARX1 I_3380  ( .D(I8150), .CLK(I5694_clk), .RSTB(I62811_rst), .Q(I63187) );
nor I_3381 (I62800,I63187,I63108);
nor I_3382 (I63218,I63187,I62862);
nand I_3383 (I62797,I62896,I63218);
not I_3384 (I62794,I63187);
DFFARX1 I_3385  ( .D(I8153), .CLK(I5694_clk), .RSTB(I62811_rst), .Q(I63263) );
not I_3386 (I63280,I63263);
nor I_3387 (I63297,I63280,I62961);
and I_3388 (I63314,I63187,I63297);
or I_3389 (I63331,I63108,I63314);
DFFARX1 I_3390  ( .D(I63331), .CLK(I5694_clk), .RSTB(I62811_rst), .Q(I62788) );
not I_3391 (I63362,I63280);
nor I_3392 (I63379,I63187,I63362);
nand I_3393 (I62791,I63280,I63379);
nand I_3394 (I62785,I62944,I63362);
not I_3395 (I63457_rst,I5701);
not I_3396 (I63474,I23603);
nor I_3397 (I63491,I23606,I23588);
nand I_3398 (I63508,I63491,I23615);
nor I_3399 (I63525,I63474,I23606);
nand I_3400 (I63542,I63525,I23594);
DFFARX1 I_3401  ( .D(I63542), .CLK(I5694_clk), .RSTB(I63457_rst), .Q(I63559) );
not I_3402 (I63428,I63559);
not I_3403 (I63590,I23606);
not I_3404 (I63607,I63590);
not I_3405 (I63624,I23600);
nor I_3406 (I63641,I63624,I23612);
and I_3407 (I63658,I63641,I23618);
or I_3408 (I63675,I63658,I23597);
DFFARX1 I_3409  ( .D(I63675), .CLK(I5694_clk), .RSTB(I63457_rst), .Q(I63692) );
DFFARX1 I_3410  ( .D(I63692), .CLK(I5694_clk), .RSTB(I63457_rst), .Q(I63425) );
DFFARX1 I_3411  ( .D(I63692), .CLK(I5694_clk), .RSTB(I63457_rst), .Q(I63723) );
DFFARX1 I_3412  ( .D(I63692), .CLK(I5694_clk), .RSTB(I63457_rst), .Q(I63419) );
nand I_3413 (I63754,I63474,I23600);
nand I_3414 (I63771,I63754,I63508);
and I_3415 (I63788,I63590,I63771);
DFFARX1 I_3416  ( .D(I63788), .CLK(I5694_clk), .RSTB(I63457_rst), .Q(I63449) );
and I_3417 (I63422,I63754,I63723);
DFFARX1 I_3418  ( .D(I23609), .CLK(I5694_clk), .RSTB(I63457_rst), .Q(I63833) );
nor I_3419 (I63446,I63833,I63754);
nor I_3420 (I63864,I63833,I63508);
nand I_3421 (I63443,I63542,I63864);
not I_3422 (I63440,I63833);
DFFARX1 I_3423  ( .D(I23591), .CLK(I5694_clk), .RSTB(I63457_rst), .Q(I63909) );
not I_3424 (I63926,I63909);
nor I_3425 (I63943,I63926,I63607);
and I_3426 (I63960,I63833,I63943);
or I_3427 (I63977,I63754,I63960);
DFFARX1 I_3428  ( .D(I63977), .CLK(I5694_clk), .RSTB(I63457_rst), .Q(I63434) );
not I_3429 (I64008,I63926);
nor I_3430 (I64025,I63833,I64008);
nand I_3431 (I63437,I63926,I64025);
nand I_3432 (I63431,I63590,I64008);
not I_3433 (I64103_rst,I5701);
not I_3434 (I64120,I55674);
nor I_3435 (I64137,I55653,I55665);
nand I_3436 (I64154,I64137,I55668);
nor I_3437 (I64171,I64120,I55653);
nand I_3438 (I64188,I64171,I55650);
DFFARX1 I_3439  ( .D(I64188), .CLK(I5694_clk), .RSTB(I64103_rst), .Q(I64205) );
not I_3440 (I64074,I64205);
not I_3441 (I64236,I55653);
not I_3442 (I64253,I64236);
not I_3443 (I64270,I55671);
nor I_3444 (I64287,I64270,I55662);
and I_3445 (I64304,I64287,I55656);
or I_3446 (I64321,I64304,I55680);
DFFARX1 I_3447  ( .D(I64321), .CLK(I5694_clk), .RSTB(I64103_rst), .Q(I64338) );
DFFARX1 I_3448  ( .D(I64338), .CLK(I5694_clk), .RSTB(I64103_rst), .Q(I64071) );
DFFARX1 I_3449  ( .D(I64338), .CLK(I5694_clk), .RSTB(I64103_rst), .Q(I64369) );
DFFARX1 I_3450  ( .D(I64338), .CLK(I5694_clk), .RSTB(I64103_rst), .Q(I64065) );
nand I_3451 (I64400,I64120,I55671);
nand I_3452 (I64417,I64400,I64154);
and I_3453 (I64434,I64236,I64417);
DFFARX1 I_3454  ( .D(I64434), .CLK(I5694_clk), .RSTB(I64103_rst), .Q(I64095) );
and I_3455 (I64068,I64400,I64369);
DFFARX1 I_3456  ( .D(I55677), .CLK(I5694_clk), .RSTB(I64103_rst), .Q(I64479) );
nor I_3457 (I64092,I64479,I64400);
nor I_3458 (I64510,I64479,I64154);
nand I_3459 (I64089,I64188,I64510);
not I_3460 (I64086,I64479);
DFFARX1 I_3461  ( .D(I55659), .CLK(I5694_clk), .RSTB(I64103_rst), .Q(I64555) );
not I_3462 (I64572,I64555);
nor I_3463 (I64589,I64572,I64253);
and I_3464 (I64606,I64479,I64589);
or I_3465 (I64623,I64400,I64606);
DFFARX1 I_3466  ( .D(I64623), .CLK(I5694_clk), .RSTB(I64103_rst), .Q(I64080) );
not I_3467 (I64654,I64572);
nor I_3468 (I64671,I64479,I64654);
nand I_3469 (I64083,I64572,I64671);
nand I_3470 (I64077,I64236,I64654);
not I_3471 (I64749_rst,I5701);
not I_3472 (I64766,I14653);
nor I_3473 (I64783,I14632,I14644);
nand I_3474 (I64800,I64783,I14647);
nor I_3475 (I64817,I64766,I14632);
nand I_3476 (I64834,I64817,I14629);
DFFARX1 I_3477  ( .D(I64834), .CLK(I5694_clk), .RSTB(I64749_rst), .Q(I64851) );
not I_3478 (I64720,I64851);
not I_3479 (I64882,I14632);
not I_3480 (I64899,I64882);
not I_3481 (I64916,I14650);
nor I_3482 (I64933,I64916,I14641);
and I_3483 (I64950,I64933,I14635);
or I_3484 (I64967,I64950,I14659);
DFFARX1 I_3485  ( .D(I64967), .CLK(I5694_clk), .RSTB(I64749_rst), .Q(I64984) );
DFFARX1 I_3486  ( .D(I64984), .CLK(I5694_clk), .RSTB(I64749_rst), .Q(I64717) );
DFFARX1 I_3487  ( .D(I64984), .CLK(I5694_clk), .RSTB(I64749_rst), .Q(I65015) );
DFFARX1 I_3488  ( .D(I64984), .CLK(I5694_clk), .RSTB(I64749_rst), .Q(I64711) );
nand I_3489 (I65046,I64766,I14650);
nand I_3490 (I65063,I65046,I64800);
and I_3491 (I65080,I64882,I65063);
DFFARX1 I_3492  ( .D(I65080), .CLK(I5694_clk), .RSTB(I64749_rst), .Q(I64741) );
and I_3493 (I64714,I65046,I65015);
DFFARX1 I_3494  ( .D(I14656), .CLK(I5694_clk), .RSTB(I64749_rst), .Q(I65125) );
nor I_3495 (I64738,I65125,I65046);
nor I_3496 (I65156,I65125,I64800);
nand I_3497 (I64735,I64834,I65156);
not I_3498 (I64732,I65125);
DFFARX1 I_3499  ( .D(I14638), .CLK(I5694_clk), .RSTB(I64749_rst), .Q(I65201) );
not I_3500 (I65218,I65201);
nor I_3501 (I65235,I65218,I64899);
and I_3502 (I65252,I65125,I65235);
or I_3503 (I65269,I65046,I65252);
DFFARX1 I_3504  ( .D(I65269), .CLK(I5694_clk), .RSTB(I64749_rst), .Q(I64726) );
not I_3505 (I65300,I65218);
nor I_3506 (I65317,I65125,I65300);
nand I_3507 (I64729,I65218,I65317);
nand I_3508 (I64723,I64882,I65300);
not I_3509 (I65395_rst,I5701);
or I_3510 (I65412,I38456,I38441);
or I_3511 (I65429,I38429,I38456);
nor I_3512 (I65446,I38435,I38459);
DFFARX1 I_3513  ( .D(I65446), .CLK(I5694_clk), .RSTB(I65395_rst), .Q(I65463) );
DFFARX1 I_3514  ( .D(I65446), .CLK(I5694_clk), .RSTB(I65395_rst), .Q(I65357) );
not I_3515 (I65494,I38435);
and I_3516 (I65511,I65494,I38432);
nor I_3517 (I65528,I65511,I38441);
nor I_3518 (I65545,I38447,I38444);
DFFARX1 I_3519  ( .D(I65545), .CLK(I5694_clk), .RSTB(I65395_rst), .Q(I65562) );
not I_3520 (I65579,I65562);
DFFARX1 I_3521  ( .D(I65562), .CLK(I5694_clk), .RSTB(I65395_rst), .Q(I65366) );
nor I_3522 (I65610,I38447,I38429);
and I_3523 (I65360,I65610,I65463);
DFFARX1 I_3524  ( .D(I38438), .CLK(I5694_clk), .RSTB(I65395_rst), .Q(I65641) );
and I_3525 (I65658,I65641,I38453);
nand I_3526 (I65675,I65658,I65429);
and I_3527 (I65692,I65562,I65675);
DFFARX1 I_3528  ( .D(I65692), .CLK(I5694_clk), .RSTB(I65395_rst), .Q(I65387) );
nor I_3529 (I65384,I65658,I65528);
not I_3530 (I65737,I65658);
nor I_3531 (I65754,I65412,I65737);
nor I_3532 (I65771,I65658,I65610);
nand I_3533 (I65381,I65429,I65771);
nor I_3534 (I65802,I65658,I65579);
not I_3535 (I65378,I65658);
nand I_3536 (I65369,I65658,I65579);
DFFARX1 I_3537  ( .D(I38450), .CLK(I5694_clk), .RSTB(I65395_rst), .Q(I65847) );
and I_3538 (I65864,I65847,I65754);
or I_3539 (I65881,I65412,I65864);
DFFARX1 I_3540  ( .D(I65881), .CLK(I5694_clk), .RSTB(I65395_rst), .Q(I65372) );
nand I_3541 (I65375,I65847,I65802);
nand I_3542 (I65926,I65847,I65528);
and I_3543 (I65943,I65446,I65926);
DFFARX1 I_3544  ( .D(I65943), .CLK(I5694_clk), .RSTB(I65395_rst), .Q(I65363) );
not I_3545 (I66007_rst,I5701);
or I_3546 (I66024,I54336,I54324);
or I_3547 (I66041,I54333,I54336);
nor I_3548 (I66058,I54327,I54348);
DFFARX1 I_3549  ( .D(I66058), .CLK(I5694_clk), .RSTB(I66007_rst), .Q(I66075) );
DFFARX1 I_3550  ( .D(I66058), .CLK(I5694_clk), .RSTB(I66007_rst), .Q(I65969) );
not I_3551 (I66106,I54327);
and I_3552 (I66123,I66106,I54342);
nor I_3553 (I66140,I66123,I54324);
nor I_3554 (I66157,I54339,I54354);
DFFARX1 I_3555  ( .D(I66157), .CLK(I5694_clk), .RSTB(I66007_rst), .Q(I66174) );
not I_3556 (I66191,I66174);
DFFARX1 I_3557  ( .D(I66174), .CLK(I5694_clk), .RSTB(I66007_rst), .Q(I65978) );
nor I_3558 (I66222,I54339,I54333);
and I_3559 (I65972,I66222,I66075);
DFFARX1 I_3560  ( .D(I54351), .CLK(I5694_clk), .RSTB(I66007_rst), .Q(I66253) );
and I_3561 (I66270,I66253,I54330);
nand I_3562 (I66287,I66270,I66041);
and I_3563 (I66304,I66174,I66287);
DFFARX1 I_3564  ( .D(I66304), .CLK(I5694_clk), .RSTB(I66007_rst), .Q(I65999) );
nor I_3565 (I65996,I66270,I66140);
not I_3566 (I66349,I66270);
nor I_3567 (I66366,I66024,I66349);
nor I_3568 (I66383,I66270,I66222);
nand I_3569 (I65993,I66041,I66383);
nor I_3570 (I66414,I66270,I66191);
not I_3571 (I65990,I66270);
nand I_3572 (I65981,I66270,I66191);
DFFARX1 I_3573  ( .D(I54345), .CLK(I5694_clk), .RSTB(I66007_rst), .Q(I66459) );
and I_3574 (I66476,I66459,I66366);
or I_3575 (I66493,I66024,I66476);
DFFARX1 I_3576  ( .D(I66493), .CLK(I5694_clk), .RSTB(I66007_rst), .Q(I65984) );
nand I_3577 (I65987,I66459,I66414);
nand I_3578 (I66538,I66459,I66140);
and I_3579 (I66555,I66058,I66538);
DFFARX1 I_3580  ( .D(I66555), .CLK(I5694_clk), .RSTB(I66007_rst), .Q(I65975) );
not I_3581 (I66619_rst,I5701);
nand I_3582 (I66636,I62142,I62139);
and I_3583 (I66653,I66636,I62151);
DFFARX1 I_3584  ( .D(I66653), .CLK(I5694_clk), .RSTB(I66619_rst), .Q(I66670) );
not I_3585 (I66687,I66670);
DFFARX1 I_3586  ( .D(I66670), .CLK(I5694_clk), .RSTB(I66619_rst), .Q(I66587) );
nor I_3587 (I66718,I62148,I62139);
DFFARX1 I_3588  ( .D(I62154), .CLK(I5694_clk), .RSTB(I66619_rst), .Q(I66735) );
DFFARX1 I_3589  ( .D(I66735), .CLK(I5694_clk), .RSTB(I66619_rst), .Q(I66752) );
not I_3590 (I66590,I66752);
DFFARX1 I_3591  ( .D(I66735), .CLK(I5694_clk), .RSTB(I66619_rst), .Q(I66783) );
and I_3592 (I66584,I66670,I66783);
nand I_3593 (I66814,I62130,I62133);
and I_3594 (I66831,I66814,I62157);
DFFARX1 I_3595  ( .D(I66831), .CLK(I5694_clk), .RSTB(I66619_rst), .Q(I66848) );
nor I_3596 (I66865,I66848,I66687);
not I_3597 (I66882,I66848);
nand I_3598 (I66593,I66670,I66882);
DFFARX1 I_3599  ( .D(I62136), .CLK(I5694_clk), .RSTB(I66619_rst), .Q(I66913) );
and I_3600 (I66930,I66913,I62127);
nor I_3601 (I66947,I66930,I66848);
nor I_3602 (I66964,I66930,I66882);
nand I_3603 (I66599,I66718,I66964);
not I_3604 (I66602,I66930);
DFFARX1 I_3605  ( .D(I66930), .CLK(I5694_clk), .RSTB(I66619_rst), .Q(I66581) );
DFFARX1 I_3606  ( .D(I62145), .CLK(I5694_clk), .RSTB(I66619_rst), .Q(I67023) );
nand I_3607 (I67040,I67023,I66735);
and I_3608 (I67057,I66718,I67040);
DFFARX1 I_3609  ( .D(I67057), .CLK(I5694_clk), .RSTB(I66619_rst), .Q(I66611) );
nor I_3610 (I66608,I67023,I66930);
and I_3611 (I67102,I67023,I66865);
or I_3612 (I67119,I66718,I67102);
DFFARX1 I_3613  ( .D(I67119), .CLK(I5694_clk), .RSTB(I66619_rst), .Q(I66596) );
nand I_3614 (I66605,I67023,I66947);
not I_3615 (I67197_rst,I5701);
nand I_3616 (I67214,I7499,I7478);
and I_3617 (I67231,I67214,I7475);
DFFARX1 I_3618  ( .D(I67231), .CLK(I5694_clk), .RSTB(I67197_rst), .Q(I67248) );
not I_3619 (I67265,I67248);
DFFARX1 I_3620  ( .D(I67248), .CLK(I5694_clk), .RSTB(I67197_rst), .Q(I67165) );
nor I_3621 (I67296,I7484,I7478);
DFFARX1 I_3622  ( .D(I7472), .CLK(I5694_clk), .RSTB(I67197_rst), .Q(I67313) );
DFFARX1 I_3623  ( .D(I67313), .CLK(I5694_clk), .RSTB(I67197_rst), .Q(I67330) );
not I_3624 (I67168,I67330);
DFFARX1 I_3625  ( .D(I67313), .CLK(I5694_clk), .RSTB(I67197_rst), .Q(I67361) );
and I_3626 (I67162,I67248,I67361);
nand I_3627 (I67392,I7502,I7493);
and I_3628 (I67409,I67392,I7490);
DFFARX1 I_3629  ( .D(I67409), .CLK(I5694_clk), .RSTB(I67197_rst), .Q(I67426) );
nor I_3630 (I67443,I67426,I67265);
not I_3631 (I67460,I67426);
nand I_3632 (I67171,I67248,I67460);
DFFARX1 I_3633  ( .D(I7487), .CLK(I5694_clk), .RSTB(I67197_rst), .Q(I67491) );
and I_3634 (I67508,I67491,I7496);
nor I_3635 (I67525,I67508,I67426);
nor I_3636 (I67542,I67508,I67460);
nand I_3637 (I67177,I67296,I67542);
not I_3638 (I67180,I67508);
DFFARX1 I_3639  ( .D(I67508), .CLK(I5694_clk), .RSTB(I67197_rst), .Q(I67159) );
DFFARX1 I_3640  ( .D(I7481), .CLK(I5694_clk), .RSTB(I67197_rst), .Q(I67601) );
nand I_3641 (I67618,I67601,I67313);
and I_3642 (I67635,I67296,I67618);
DFFARX1 I_3643  ( .D(I67635), .CLK(I5694_clk), .RSTB(I67197_rst), .Q(I67189) );
nor I_3644 (I67186,I67601,I67508);
and I_3645 (I67680,I67601,I67443);
or I_3646 (I67697,I67296,I67680);
DFFARX1 I_3647  ( .D(I67697), .CLK(I5694_clk), .RSTB(I67197_rst), .Q(I67174) );
nand I_3648 (I67183,I67601,I67525);
not I_3649 (I67775_rst,I5701);
nand I_3650 (I67792,I60204,I60201);
and I_3651 (I67809,I67792,I60213);
DFFARX1 I_3652  ( .D(I67809), .CLK(I5694_clk), .RSTB(I67775_rst), .Q(I67826) );
not I_3653 (I67843,I67826);
DFFARX1 I_3654  ( .D(I67826), .CLK(I5694_clk), .RSTB(I67775_rst), .Q(I67743) );
nor I_3655 (I67874,I60210,I60201);
DFFARX1 I_3656  ( .D(I60216), .CLK(I5694_clk), .RSTB(I67775_rst), .Q(I67891) );
DFFARX1 I_3657  ( .D(I67891), .CLK(I5694_clk), .RSTB(I67775_rst), .Q(I67908) );
not I_3658 (I67746,I67908);
DFFARX1 I_3659  ( .D(I67891), .CLK(I5694_clk), .RSTB(I67775_rst), .Q(I67939) );
and I_3660 (I67740,I67826,I67939);
nand I_3661 (I67970,I60192,I60195);
and I_3662 (I67987,I67970,I60219);
DFFARX1 I_3663  ( .D(I67987), .CLK(I5694_clk), .RSTB(I67775_rst), .Q(I68004) );
nor I_3664 (I68021,I68004,I67843);
not I_3665 (I68038,I68004);
nand I_3666 (I67749,I67826,I68038);
DFFARX1 I_3667  ( .D(I60198), .CLK(I5694_clk), .RSTB(I67775_rst), .Q(I68069) );
and I_3668 (I68086,I68069,I60189);
nor I_3669 (I68103,I68086,I68004);
nor I_3670 (I68120,I68086,I68038);
nand I_3671 (I67755,I67874,I68120);
not I_3672 (I67758,I68086);
DFFARX1 I_3673  ( .D(I68086), .CLK(I5694_clk), .RSTB(I67775_rst), .Q(I67737) );
DFFARX1 I_3674  ( .D(I60207), .CLK(I5694_clk), .RSTB(I67775_rst), .Q(I68179) );
nand I_3675 (I68196,I68179,I67891);
and I_3676 (I68213,I67874,I68196);
DFFARX1 I_3677  ( .D(I68213), .CLK(I5694_clk), .RSTB(I67775_rst), .Q(I67767) );
nor I_3678 (I67764,I68179,I68086);
and I_3679 (I68258,I68179,I68021);
or I_3680 (I68275,I67874,I68258);
DFFARX1 I_3681  ( .D(I68275), .CLK(I5694_clk), .RSTB(I67775_rst), .Q(I67752) );
nand I_3682 (I67761,I68179,I68103);
not I_3683 (I68353_rst,I5701);
nand I_3684 (I68370,I34432,I34444);
and I_3685 (I68387,I68370,I34417);
DFFARX1 I_3686  ( .D(I68387), .CLK(I5694_clk), .RSTB(I68353_rst), .Q(I68404) );
not I_3687 (I68421,I68404);
DFFARX1 I_3688  ( .D(I68404), .CLK(I5694_clk), .RSTB(I68353_rst), .Q(I68321) );
nor I_3689 (I68452,I34435,I34444);
DFFARX1 I_3690  ( .D(I34426), .CLK(I5694_clk), .RSTB(I68353_rst), .Q(I68469) );
DFFARX1 I_3691  ( .D(I68469), .CLK(I5694_clk), .RSTB(I68353_rst), .Q(I68486) );
not I_3692 (I68324,I68486);
DFFARX1 I_3693  ( .D(I68469), .CLK(I5694_clk), .RSTB(I68353_rst), .Q(I68517) );
and I_3694 (I68318,I68404,I68517);
nand I_3695 (I68548,I34423,I34429);
and I_3696 (I68565,I68548,I34441);
DFFARX1 I_3697  ( .D(I68565), .CLK(I5694_clk), .RSTB(I68353_rst), .Q(I68582) );
nor I_3698 (I68599,I68582,I68421);
not I_3699 (I68616,I68582);
nand I_3700 (I68327,I68404,I68616);
DFFARX1 I_3701  ( .D(I34447), .CLK(I5694_clk), .RSTB(I68353_rst), .Q(I6864_rst7) );
and I_3702 (I68664,I6864_rst7,I34438);
nor I_3703 (I68681,I68664,I68582);
nor I_3704 (I68698,I68664,I68616);
nand I_3705 (I68333,I68452,I68698);
not I_3706 (I68336,I68664);
DFFARX1 I_3707  ( .D(I68664), .CLK(I5694_clk), .RSTB(I68353_rst), .Q(I68315) );
DFFARX1 I_3708  ( .D(I34420), .CLK(I5694_clk), .RSTB(I68353_rst), .Q(I68757) );
nand I_3709 (I68774,I68757,I68469);
and I_3710 (I68791,I68452,I68774);
DFFARX1 I_3711  ( .D(I68791), .CLK(I5694_clk), .RSTB(I68353_rst), .Q(I68345) );
nor I_3712 (I68342,I68757,I68664);
and I_3713 (I68836,I68757,I68599);
or I_3714 (I68853,I68452,I68836);
DFFARX1 I_3715  ( .D(I68853), .CLK(I5694_clk), .RSTB(I68353_rst), .Q(I68330) );
nand I_3716 (I68339,I68757,I68681);
not I_3717 (I68931_rst,I5701);
nand I_3718 (I68948,I19251,I19248);
and I_3719 (I68965,I68948,I19260);
DFFARX1 I_3720  ( .D(I68965), .CLK(I5694_clk), .RSTB(I68931_rst), .Q(I68982) );
not I_3721 (I68999,I68982);
DFFARX1 I_3722  ( .D(I68982), .CLK(I5694_clk), .RSTB(I68931_rst), .Q(I68899) );
nor I_3723 (I69030,I19257,I19248);
DFFARX1 I_3724  ( .D(I19263), .CLK(I5694_clk), .RSTB(I68931_rst), .Q(I69047) );
DFFARX1 I_3725  ( .D(I69047), .CLK(I5694_clk), .RSTB(I68931_rst), .Q(I69064) );
not I_3726 (I68902,I69064);
DFFARX1 I_3727  ( .D(I69047), .CLK(I5694_clk), .RSTB(I68931_rst), .Q(I69095) );
and I_3728 (I68896,I68982,I69095);
nand I_3729 (I69126,I19239,I19242);
and I_3730 (I69143,I69126,I19266);
DFFARX1 I_3731  ( .D(I69143), .CLK(I5694_clk), .RSTB(I68931_rst), .Q(I69160) );
nor I_3732 (I69177,I69160,I68999);
not I_3733 (I69194,I69160);
nand I_3734 (I68905,I68982,I69194);
DFFARX1 I_3735  ( .D(I19245), .CLK(I5694_clk), .RSTB(I68931_rst), .Q(I69225) );
and I_3736 (I69242,I69225,I19236);
nor I_3737 (I69259,I69242,I69160);
nor I_3738 (I69276,I69242,I69194);
nand I_3739 (I68911,I69030,I69276);
not I_3740 (I68914,I69242);
DFFARX1 I_3741  ( .D(I69242), .CLK(I5694_clk), .RSTB(I68931_rst), .Q(I68893) );
DFFARX1 I_3742  ( .D(I19254), .CLK(I5694_clk), .RSTB(I68931_rst), .Q(I69335) );
nand I_3743 (I69352,I69335,I69047);
and I_3744 (I69369,I69030,I69352);
DFFARX1 I_3745  ( .D(I69369), .CLK(I5694_clk), .RSTB(I68931_rst), .Q(I68923) );
nor I_3746 (I68920,I69335,I69242);
and I_3747 (I69414,I69335,I69177);
or I_3748 (I69431,I69030,I69414);
DFFARX1 I_3749  ( .D(I69431), .CLK(I5694_clk), .RSTB(I68931_rst), .Q(I68908) );
nand I_3750 (I68917,I69335,I69259);
not I_3751 (I69509_rst,I5701);
nand I_3752 (I69526,I37322,I37337);
and I_3753 (I69543,I69526,I37325);
DFFARX1 I_3754  ( .D(I69543), .CLK(I5694_clk), .RSTB(I69509_rst), .Q(I69560) );
not I_3755 (I69577,I69560);
DFFARX1 I_3756  ( .D(I69560), .CLK(I5694_clk), .RSTB(I69509_rst), .Q(I69477) );
nor I_3757 (I69608,I37334,I37337);
DFFARX1 I_3758  ( .D(I37319), .CLK(I5694_clk), .RSTB(I69509_rst), .Q(I69625) );
DFFARX1 I_3759  ( .D(I69625), .CLK(I5694_clk), .RSTB(I69509_rst), .Q(I69642) );
not I_3760 (I69480,I69642);
DFFARX1 I_3761  ( .D(I69625), .CLK(I5694_clk), .RSTB(I69509_rst), .Q(I69673) );
and I_3762 (I69474,I69560,I69673);
nand I_3763 (I69704,I37310,I37307);
and I_3764 (I69721,I69704,I37313);
DFFARX1 I_3765  ( .D(I69721), .CLK(I5694_clk), .RSTB(I69509_rst), .Q(I69738) );
nor I_3766 (I69755,I69738,I69577);
not I_3767 (I69772,I69738);
nand I_3768 (I69483,I69560,I69772);
DFFARX1 I_3769  ( .D(I37316), .CLK(I5694_clk), .RSTB(I69509_rst), .Q(I69803) );
and I_3770 (I69820,I69803,I37328);
nor I_3771 (I69837,I69820,I69738);
nor I_3772 (I69854,I69820,I69772);
nand I_3773 (I69489,I69608,I69854);
not I_3774 (I69492,I69820);
DFFARX1 I_3775  ( .D(I69820), .CLK(I5694_clk), .RSTB(I69509_rst), .Q(I69471) );
DFFARX1 I_3776  ( .D(I37331), .CLK(I5694_clk), .RSTB(I69509_rst), .Q(I69913) );
nand I_3777 (I69930,I69913,I69625);
and I_3778 (I69947,I69608,I69930);
DFFARX1 I_3779  ( .D(I69947), .CLK(I5694_clk), .RSTB(I69509_rst), .Q(I69501) );
nor I_3780 (I69498,I69913,I69820);
and I_3781 (I69992,I69913,I69755);
or I_3782 (I70009,I69608,I69992);
DFFARX1 I_3783  ( .D(I70009), .CLK(I5694_clk), .RSTB(I69509_rst), .Q(I69486) );
nand I_3784 (I69495,I69913,I69837);
not I_3785 (I70087_rst,I5701);
nand I_3786 (I70104,I44094,I44076);
and I_3787 (I70121,I70104,I44088);
DFFARX1 I_3788  ( .D(I70121), .CLK(I5694_clk), .RSTB(I70087_rst), .Q(I70138) );
not I_3789 (I70155,I70138);
DFFARX1 I_3790  ( .D(I70138), .CLK(I5694_clk), .RSTB(I70087_rst), .Q(I70055) );
nor I_3791 (I70186,I44091,I44076);
DFFARX1 I_3792  ( .D(I44100), .CLK(I5694_clk), .RSTB(I70087_rst), .Q(I70203) );
DFFARX1 I_3793  ( .D(I70203), .CLK(I5694_clk), .RSTB(I70087_rst), .Q(I70220) );
not I_3794 (I70058,I70220);
DFFARX1 I_3795  ( .D(I70203), .CLK(I5694_clk), .RSTB(I70087_rst), .Q(I70251) );
and I_3796 (I70052,I70138,I70251);
nand I_3797 (I70282,I44079,I44103);
and I_3798 (I70299,I70282,I44082);
DFFARX1 I_3799  ( .D(I70299), .CLK(I5694_clk), .RSTB(I70087_rst), .Q(I70316) );
nor I_3800 (I70333,I70316,I70155);
not I_3801 (I70350,I70316);
nand I_3802 (I70061,I70138,I70350);
DFFARX1 I_3803  ( .D(I44085), .CLK(I5694_clk), .RSTB(I70087_rst), .Q(I70381) );
and I_3804 (I70398,I70381,I44097);
nor I_3805 (I70415,I70398,I70316);
nor I_3806 (I70432,I70398,I70350);
nand I_3807 (I70067,I70186,I70432);
not I_3808 (I70070,I70398);
DFFARX1 I_3809  ( .D(I70398), .CLK(I5694_clk), .RSTB(I70087_rst), .Q(I70049) );
DFFARX1 I_3810  ( .D(I44073), .CLK(I5694_clk), .RSTB(I70087_rst), .Q(I70491) );
nand I_3811 (I70508,I70491,I70203);
and I_3812 (I70525,I70186,I70508);
DFFARX1 I_3813  ( .D(I70525), .CLK(I5694_clk), .RSTB(I70087_rst), .Q(I70079) );
nor I_3814 (I70076,I70491,I70398);
and I_3815 (I70570,I70491,I70333);
or I_3816 (I70587,I70186,I70570);
DFFARX1 I_3817  ( .D(I70587), .CLK(I5694_clk), .RSTB(I70087_rst), .Q(I70064) );
nand I_3818 (I70073,I70491,I70415);
not I_3819 (I70665_rst,I5701);
nand I_3820 (I70682,I58266,I58263);
and I_3821 (I70699,I70682,I58275);
DFFARX1 I_3822  ( .D(I70699), .CLK(I5694_clk), .RSTB(I70665_rst), .Q(I70716) );
not I_3823 (I70733,I70716);
DFFARX1 I_3824  ( .D(I70716), .CLK(I5694_clk), .RSTB(I70665_rst), .Q(I70633) );
nor I_3825 (I70764,I58272,I58263);
DFFARX1 I_3826  ( .D(I58278), .CLK(I5694_clk), .RSTB(I70665_rst), .Q(I70781) );
DFFARX1 I_3827  ( .D(I70781), .CLK(I5694_clk), .RSTB(I70665_rst), .Q(I70798) );
not I_3828 (I70636,I70798);
DFFARX1 I_3829  ( .D(I70781), .CLK(I5694_clk), .RSTB(I70665_rst), .Q(I70829) );
and I_3830 (I70630,I70716,I70829);
nand I_3831 (I70860,I58254,I58257);
and I_3832 (I70877,I70860,I58281);
DFFARX1 I_3833  ( .D(I70877), .CLK(I5694_clk), .RSTB(I70665_rst), .Q(I70894) );
nor I_3834 (I70911,I70894,I70733);
not I_3835 (I70928,I70894);
nand I_3836 (I70639,I70716,I70928);
DFFARX1 I_3837  ( .D(I58260), .CLK(I5694_clk), .RSTB(I70665_rst), .Q(I70959) );
and I_3838 (I70976,I70959,I58251);
nor I_3839 (I70993,I70976,I70894);
nor I_3840 (I71010,I70976,I70928);
nand I_3841 (I70645,I70764,I71010);
not I_3842 (I70648,I70976);
DFFARX1 I_3843  ( .D(I70976), .CLK(I5694_clk), .RSTB(I70665_rst), .Q(I70627) );
DFFARX1 I_3844  ( .D(I58269), .CLK(I5694_clk), .RSTB(I70665_rst), .Q(I71069) );
nand I_3845 (I71086,I71069,I70781);
and I_3846 (I71103,I70764,I71086);
DFFARX1 I_3847  ( .D(I71103), .CLK(I5694_clk), .RSTB(I70665_rst), .Q(I70657) );
nor I_3848 (I70654,I71069,I70976);
and I_3849 (I71148,I71069,I70911);
or I_3850 (I71165,I70764,I71148);
DFFARX1 I_3851  ( .D(I71165), .CLK(I5694_clk), .RSTB(I70665_rst), .Q(I70642) );
nand I_3852 (I70651,I71069,I70993);
not I_3853 (I71243_rst,I5701);
nand I_3854 (I71260,I25940,I25964);
and I_3855 (I71277,I71260,I25946);
DFFARX1 I_3856  ( .D(I71277), .CLK(I5694_clk), .RSTB(I71243_rst), .Q(I71294) );
not I_3857 (I71311,I71294);
DFFARX1 I_3858  ( .D(I71294), .CLK(I5694_clk), .RSTB(I71243_rst), .Q(I71211) );
nor I_3859 (I71342,I25934,I25964);
DFFARX1 I_3860  ( .D(I25949), .CLK(I5694_clk), .RSTB(I71243_rst), .Q(I71359) );
DFFARX1 I_3861  ( .D(I71359), .CLK(I5694_clk), .RSTB(I71243_rst), .Q(I71376) );
not I_3862 (I71214,I71376);
DFFARX1 I_3863  ( .D(I71359), .CLK(I5694_clk), .RSTB(I71243_rst), .Q(I71407) );
and I_3864 (I71208,I71294,I71407);
nand I_3865 (I71438,I25955,I25937);
and I_3866 (I71455,I71438,I25958);
DFFARX1 I_3867  ( .D(I71455), .CLK(I5694_clk), .RSTB(I71243_rst), .Q(I71472) );
nor I_3868 (I71489,I71472,I71311);
not I_3869 (I71506,I71472);
nand I_3870 (I71217,I71294,I71506);
DFFARX1 I_3871  ( .D(I25943), .CLK(I5694_clk), .RSTB(I71243_rst), .Q(I71537) );
and I_3872 (I71554,I71537,I25952);
nor I_3873 (I71571,I71554,I71472);
nor I_3874 (I71588,I71554,I71506);
nand I_3875 (I71223,I71342,I71588);
not I_3876 (I71226,I71554);
DFFARX1 I_3877  ( .D(I71554), .CLK(I5694_clk), .RSTB(I71243_rst), .Q(I71205) );
DFFARX1 I_3878  ( .D(I25961), .CLK(I5694_clk), .RSTB(I71243_rst), .Q(I71647) );
nand I_3879 (I71664,I71647,I71359);
and I_3880 (I71681,I71342,I71664);
DFFARX1 I_3881  ( .D(I71681), .CLK(I5694_clk), .RSTB(I71243_rst), .Q(I71235) );
nor I_3882 (I71232,I71647,I71554);
and I_3883 (I71726,I71647,I71489);
or I_3884 (I71743,I71342,I71726);
DFFARX1 I_3885  ( .D(I71743), .CLK(I5694_clk), .RSTB(I71243_rst), .Q(I71220) );
nand I_3886 (I71229,I71647,I71571);
not I_3887 (I71821_rst,I5701);
or I_3888 (I71838,I30114,I30099);
or I_3889 (I71855,I30126,I30114);
nor I_3890 (I71872,I30108,I30102);
not I_3891 (I71889,I71872);
DFFARX1 I_3892  ( .D(I71872), .CLK(I5694_clk), .RSTB(I71821_rst), .Q(I71789) );
nand I_3893 (I71920,I71872,I71838);
not I_3894 (I71937,I30108);
and I_3895 (I71954,I71937,I30105);
nor I_3896 (I71971,I71954,I30099);
nor I_3897 (I71988,I30120,I30129);
DFFARX1 I_3898  ( .D(I71988), .CLK(I5694_clk), .RSTB(I71821_rst), .Q(I72005) );
nor I_3899 (I72022,I72005,I71889);
not I_3900 (I72039,I72005);
nand I_3901 (I71795,I71872,I72039);
DFFARX1 I_3902  ( .D(I72005), .CLK(I5694_clk), .RSTB(I71821_rst), .Q(I71786) );
nor I_3903 (I72084,I30120,I30126);
nand I_3904 (I72101,I71855,I72084);
nor I_3905 (I71810,I71838,I72084);
and I_3906 (I72132,I72084,I72022);
or I_3907 (I72149,I71971,I72132);
DFFARX1 I_3908  ( .D(I72149), .CLK(I5694_clk), .RSTB(I71821_rst), .Q(I71798) );
DFFARX1 I_3909  ( .D(I30111), .CLK(I5694_clk), .RSTB(I71821_rst), .Q(I72180) );
and I_3910 (I72197,I72180,I30117);
not I_3911 (I71804,I72197);
DFFARX1 I_3912  ( .D(I72197), .CLK(I5694_clk), .RSTB(I71821_rst), .Q(I72228) );
not I_3913 (I71792,I72228);
and I_3914 (I72259,I72197,I71920);
DFFARX1 I_3915  ( .D(I72259), .CLK(I5694_clk), .RSTB(I71821_rst), .Q(I71783) );
DFFARX1 I_3916  ( .D(I30123), .CLK(I5694_clk), .RSTB(I71821_rst), .Q(I72290) );
and I_3917 (I72307,I72290,I72101);
DFFARX1 I_3918  ( .D(I72307), .CLK(I5694_clk), .RSTB(I71821_rst), .Q(I71813) );
nor I_3919 (I72338,I72290,I72197);
nand I_3920 (I71807,I71971,I72338);
nor I_3921 (I72369,I72290,I72039);
nand I_3922 (I71801,I71855,I72369);
not I_3923 (I72433_rst,I5701);
nand I_3924 (I72450,I21816,I21804);
and I_3925 (I72467,I72450,I21810);
DFFARX1 I_3926  ( .D(I72467), .CLK(I5694_clk), .RSTB(I72433_rst), .Q(I72484) );
nor I_3927 (I72501,I21801,I21804);
nor I_3928 (I72518,I72501,I72484);
not I_3929 (I72416,I72501);
DFFARX1 I_3930  ( .D(I21786), .CLK(I5694_clk), .RSTB(I72433_rst), .Q(I72549) );
not I_3931 (I72566,I72549);
nor I_3932 (I72583,I72501,I72566);
nand I_3933 (I72419,I72549,I72518);
DFFARX1 I_3934  ( .D(I72549), .CLK(I5694_clk), .RSTB(I72433_rst), .Q(I72401) );
nand I_3935 (I72628,I21795,I21813);
and I_3936 (I72645,I72628,I21807);
DFFARX1 I_3937  ( .D(I72645), .CLK(I5694_clk), .RSTB(I72433_rst), .Q(I72662) );
nor I_3938 (I72422,I72662,I72484);
nand I_3939 (I72413,I72662,I72583);
DFFARX1 I_3940  ( .D(I21798), .CLK(I5694_clk), .RSTB(I72433_rst), .Q(I72707) );
and I_3941 (I72724,I72707,I21792);
DFFARX1 I_3942  ( .D(I72724), .CLK(I5694_clk), .RSTB(I72433_rst), .Q(I72741) );
not I_3943 (I72404,I72741);
nand I_3944 (I72772,I72724,I72662);
and I_3945 (I72789,I72484,I72772);
DFFARX1 I_3946  ( .D(I72789), .CLK(I5694_clk), .RSTB(I72433_rst), .Q(I72395) );
DFFARX1 I_3947  ( .D(I21789), .CLK(I5694_clk), .RSTB(I72433_rst), .Q(I72820) );
nand I_3948 (I72837,I72820,I72484);
and I_3949 (I72854,I72662,I72837);
DFFARX1 I_3950  ( .D(I72854), .CLK(I5694_clk), .RSTB(I72433_rst), .Q(I72425) );
not I_3951 (I72885,I72820);
nor I_3952 (I72902,I72501,I72885);
and I_3953 (I72919,I72820,I72902);
or I_3954 (I72936,I72724,I72919);
DFFARX1 I_3955  ( .D(I72936), .CLK(I5694_clk), .RSTB(I72433_rst), .Q(I72410) );
nand I_3956 (I72407,I72820,I72566);
DFFARX1 I_3957  ( .D(I72820), .CLK(I5694_clk), .RSTB(I72433_rst), .Q(I72398) );
not I_3958 (I73028_rst,I5701);
nand I_3959 (I73045,I28924,I28915);
and I_3960 (I73062,I73045,I28933);
DFFARX1 I_3961  ( .D(I73062), .CLK(I5694_clk), .RSTB(I73028_rst), .Q(I73079) );
nor I_3962 (I73096,I28912,I28915);
nor I_3963 (I73113,I73096,I73079);
not I_3964 (I73011,I73096);
DFFARX1 I_3965  ( .D(I28921), .CLK(I5694_clk), .RSTB(I73028_rst), .Q(I73144) );
not I_3966 (I73161,I73144);
nor I_3967 (I73178,I73096,I73161);
nand I_3968 (I73014,I73144,I73113);
DFFARX1 I_3969  ( .D(I73144), .CLK(I5694_clk), .RSTB(I73028_rst), .Q(I72996) );
nand I_3970 (I73223,I28936,I28918);
and I_3971 (I73240,I73223,I28939);
DFFARX1 I_3972  ( .D(I73240), .CLK(I5694_clk), .RSTB(I73028_rst), .Q(I73257) );
nor I_3973 (I73017,I73257,I73079);
nand I_3974 (I73008,I73257,I73178);
DFFARX1 I_3975  ( .D(I28927), .CLK(I5694_clk), .RSTB(I73028_rst), .Q(I73302) );
and I_3976 (I73319,I73302,I28909);
DFFARX1 I_3977  ( .D(I73319), .CLK(I5694_clk), .RSTB(I73028_rst), .Q(I73336) );
not I_3978 (I72999,I73336);
nand I_3979 (I73367,I73319,I73257);
and I_3980 (I73384,I73079,I73367);
DFFARX1 I_3981  ( .D(I73384), .CLK(I5694_clk), .RSTB(I73028_rst), .Q(I72990) );
DFFARX1 I_3982  ( .D(I28930), .CLK(I5694_clk), .RSTB(I73028_rst), .Q(I73415) );
nand I_3983 (I73432,I73415,I73079);
and I_3984 (I73449,I73257,I73432);
DFFARX1 I_3985  ( .D(I73449), .CLK(I5694_clk), .RSTB(I73028_rst), .Q(I73020) );
not I_3986 (I73480,I73415);
nor I_3987 (I73497,I73096,I73480);
and I_3988 (I73514,I73415,I73497);
or I_3989 (I73531,I73319,I73514);
DFFARX1 I_3990  ( .D(I73531), .CLK(I5694_clk), .RSTB(I73028_rst), .Q(I73005) );
nand I_3991 (I73002,I73415,I73161);
DFFARX1 I_3992  ( .D(I73415), .CLK(I5694_clk), .RSTB(I73028_rst), .Q(I72993) );
not I_3993 (I73623_rst,I5701);
nand I_3994 (I73640,I28329,I28320);
and I_3995 (I73657,I73640,I28338);
DFFARX1 I_3996  ( .D(I73657), .CLK(I5694_clk), .RSTB(I73623_rst), .Q(I73674) );
nor I_3997 (I73691,I28317,I28320);
nor I_3998 (I73708,I73691,I73674);
not I_3999 (I73606,I73691);
DFFARX1 I_4000  ( .D(I28326), .CLK(I5694_clk), .RSTB(I73623_rst), .Q(I73739) );
not I_4001 (I73756,I73739);
nor I_4002 (I73773,I73691,I73756);
nand I_4003 (I73609,I73739,I73708);
DFFARX1 I_4004  ( .D(I73739), .CLK(I5694_clk), .RSTB(I73623_rst), .Q(I73591) );
nand I_4005 (I73818,I28341,I28323);
and I_4006 (I73835,I73818,I28344);
DFFARX1 I_4007  ( .D(I73835), .CLK(I5694_clk), .RSTB(I73623_rst), .Q(I73852) );
nor I_4008 (I73612,I73852,I73674);
nand I_4009 (I73603,I73852,I73773);
DFFARX1 I_4010  ( .D(I28332), .CLK(I5694_clk), .RSTB(I73623_rst), .Q(I73897) );
and I_4011 (I73914,I73897,I28314);
DFFARX1 I_4012  ( .D(I73914), .CLK(I5694_clk), .RSTB(I73623_rst), .Q(I73931) );
not I_4013 (I73594,I73931);
nand I_4014 (I73962,I73914,I73852);
and I_4015 (I73979,I73674,I73962);
DFFARX1 I_4016  ( .D(I73979), .CLK(I5694_clk), .RSTB(I73623_rst), .Q(I73585) );
DFFARX1 I_4017  ( .D(I28335), .CLK(I5694_clk), .RSTB(I73623_rst), .Q(I74010) );
nand I_4018 (I74027,I74010,I73674);
and I_4019 (I74044,I73852,I74027);
DFFARX1 I_4020  ( .D(I74044), .CLK(I5694_clk), .RSTB(I73623_rst), .Q(I73615) );
not I_4021 (I74075,I74010);
nor I_4022 (I74092,I73691,I74075);
and I_4023 (I74109,I74010,I74092);
or I_4024 (I74126,I73914,I74109);
DFFARX1 I_4025  ( .D(I74126), .CLK(I5694_clk), .RSTB(I73623_rst), .Q(I73600) );
nand I_4026 (I73597,I74010,I73756);
DFFARX1 I_4027  ( .D(I74010), .CLK(I5694_clk), .RSTB(I73623_rst), .Q(I73588) );
not I_4028 (I74218_rst,I5701);
nand I_4029 (I74235,I52353,I52359);
and I_4030 (I74252,I74235,I52341);
DFFARX1 I_4031  ( .D(I74252), .CLK(I5694_clk), .RSTB(I74218_rst), .Q(I74269) );
nor I_4032 (I74286,I52335,I52359);
nor I_4033 (I74303,I74286,I74269);
not I_4034 (I74201,I74286);
DFFARX1 I_4035  ( .D(I52365), .CLK(I5694_clk), .RSTB(I74218_rst), .Q(I74334) );
not I_4036 (I74351,I74334);
nor I_4037 (I74368,I74286,I74351);
nand I_4038 (I74204,I74334,I74303);
DFFARX1 I_4039  ( .D(I74334), .CLK(I5694_clk), .RSTB(I74218_rst), .Q(I74186) );
nand I_4040 (I74413,I52356,I52347);
and I_4041 (I74430,I74413,I52350);
DFFARX1 I_4042  ( .D(I74430), .CLK(I5694_clk), .RSTB(I74218_rst), .Q(I74447) );
nor I_4043 (I74207,I74447,I74269);
nand I_4044 (I74198,I74447,I74368);
DFFARX1 I_4045  ( .D(I52362), .CLK(I5694_clk), .RSTB(I74218_rst), .Q(I74492) );
and I_4046 (I74509,I74492,I52338);
DFFARX1 I_4047  ( .D(I74509), .CLK(I5694_clk), .RSTB(I74218_rst), .Q(I74526) );
not I_4048 (I74189,I74526);
nand I_4049 (I74557,I74509,I74447);
and I_4050 (I74574,I74269,I74557);
DFFARX1 I_4051  ( .D(I74574), .CLK(I5694_clk), .RSTB(I74218_rst), .Q(I74180) );
DFFARX1 I_4052  ( .D(I52344), .CLK(I5694_clk), .RSTB(I74218_rst), .Q(I74605) );
nand I_4053 (I74622,I74605,I74269);
and I_4054 (I74639,I74447,I74622);
DFFARX1 I_4055  ( .D(I74639), .CLK(I5694_clk), .RSTB(I74218_rst), .Q(I74210) );
not I_4056 (I74670,I74605);
nor I_4057 (I74687,I74286,I74670);
and I_4058 (I74704,I74605,I74687);
or I_4059 (I74721,I74509,I74704);
DFFARX1 I_4060  ( .D(I74721), .CLK(I5694_clk), .RSTB(I74218_rst), .Q(I74195) );
nand I_4061 (I74192,I74605,I74351);
DFFARX1 I_4062  ( .D(I74605), .CLK(I5694_clk), .RSTB(I74218_rst), .Q(I74183) );
not I_4063 (I74813_rst,I5701);
nand I_4064 (I74830,I61499,I61511);
and I_4065 (I74847,I74830,I61493);
DFFARX1 I_4066  ( .D(I74847), .CLK(I5694_clk), .RSTB(I74813_rst), .Q(I74864) );
nor I_4067 (I74881,I61505,I61511);
nor I_4068 (I74898,I74881,I74864);
not I_4069 (I74796,I74881);
DFFARX1 I_4070  ( .D(I61490), .CLK(I5694_clk), .RSTB(I74813_rst), .Q(I74929) );
not I_4071 (I74946,I74929);
nor I_4072 (I74963,I74881,I74946);
nand I_4073 (I74799,I74929,I74898);
DFFARX1 I_4074  ( .D(I74929), .CLK(I5694_clk), .RSTB(I74813_rst), .Q(I74781) );
nand I_4075 (I75008,I61481,I61496);
and I_4076 (I75025,I75008,I61487);
DFFARX1 I_4077  ( .D(I75025), .CLK(I5694_clk), .RSTB(I74813_rst), .Q(I75042) );
nor I_4078 (I74802,I75042,I74864);
nand I_4079 (I74793,I75042,I74963);
DFFARX1 I_4080  ( .D(I61508), .CLK(I5694_clk), .RSTB(I74813_rst), .Q(I75087) );
and I_4081 (I7510_rst4,I75087,I61502);
DFFARX1 I_4082  ( .D(I7510_rst4), .CLK(I5694_clk), .RSTB(I74813_rst), .Q(I75121) );
not I_4083 (I74784,I75121);
nand I_4084 (I75152,I7510_rst4,I75042);
and I_4085 (I75169,I74864,I75152);
DFFARX1 I_4086  ( .D(I75169), .CLK(I5694_clk), .RSTB(I74813_rst), .Q(I74775) );
DFFARX1 I_4087  ( .D(I61484), .CLK(I5694_clk), .RSTB(I74813_rst), .Q(I75200) );
nand I_4088 (I75217,I75200,I74864);
and I_4089 (I75234,I75042,I75217);
DFFARX1 I_4090  ( .D(I75234), .CLK(I5694_clk), .RSTB(I74813_rst), .Q(I74805) );
not I_4091 (I75265,I75200);
nor I_4092 (I75282,I74881,I75265);
and I_4093 (I75299,I75200,I75282);
or I_4094 (I75316,I7510_rst4,I75299);
DFFARX1 I_4095  ( .D(I75316), .CLK(I5694_clk), .RSTB(I74813_rst), .Q(I74790) );
nand I_4096 (I74787,I75200,I74946);
DFFARX1 I_4097  ( .D(I75200), .CLK(I5694_clk), .RSTB(I74813_rst), .Q(I74778) );
not I_4098 (I75408_rst,I5701);
nand I_4099 (I75425,I15973,I15979);
and I_4100 (I75442,I75425,I15961);
DFFARX1 I_4101  ( .D(I75442), .CLK(I5694_clk), .RSTB(I75408_rst), .Q(I75459) );
nor I_4102 (I75476,I15955,I15979);
nor I_4103 (I75493,I75476,I75459);
not I_4104 (I75391,I75476);
DFFARX1 I_4105  ( .D(I15985), .CLK(I5694_clk), .RSTB(I75408_rst), .Q(I75524) );
not I_4106 (I75541,I75524);
nor I_4107 (I75558,I75476,I75541);
nand I_4108 (I75394,I75524,I75493);
DFFARX1 I_4109  ( .D(I75524), .CLK(I5694_clk), .RSTB(I75408_rst), .Q(I75376) );
nand I_4110 (I75603,I15976,I15967);
and I_4111 (I75620,I75603,I15970);
DFFARX1 I_4112  ( .D(I75620), .CLK(I5694_clk), .RSTB(I75408_rst), .Q(I75637) );
nor I_4113 (I75397,I75637,I75459);
nand I_4114 (I75388,I75637,I75558);
DFFARX1 I_4115  ( .D(I15982), .CLK(I5694_clk), .RSTB(I75408_rst), .Q(I75682) );
and I_4116 (I75699,I75682,I15958);
DFFARX1 I_4117  ( .D(I75699), .CLK(I5694_clk), .RSTB(I75408_rst), .Q(I75716) );
not I_4118 (I75379,I75716);
nand I_4119 (I75747,I75699,I75637);
and I_4120 (I75764,I75459,I75747);
DFFARX1 I_4121  ( .D(I75764), .CLK(I5694_clk), .RSTB(I75408_rst), .Q(I75370) );
DFFARX1 I_4122  ( .D(I15964), .CLK(I5694_clk), .RSTB(I75408_rst), .Q(I75795) );
nand I_4123 (I75812,I75795,I75459);
and I_4124 (I75829,I75637,I75812);
DFFARX1 I_4125  ( .D(I75829), .CLK(I5694_clk), .RSTB(I75408_rst), .Q(I75400) );
not I_4126 (I75860,I75795);
nor I_4127 (I75877,I75476,I75860);
and I_4128 (I75894,I75795,I75877);
or I_4129 (I75911,I75699,I75894);
DFFARX1 I_4130  ( .D(I75911), .CLK(I5694_clk), .RSTB(I75408_rst), .Q(I75385) );
nand I_4131 (I75382,I75795,I75541);
DFFARX1 I_4132  ( .D(I75795), .CLK(I5694_clk), .RSTB(I75408_rst), .Q(I75373) );
not I_4133 (I76003_rst,I5701);
nand I_4134 (I76020,I65387,I65375);
and I_4135 (I76037,I76020,I65381);
DFFARX1 I_4136  ( .D(I76037), .CLK(I5694_clk), .RSTB(I76003_rst), .Q(I76054) );
nor I_4137 (I76071,I65372,I65375);
nor I_4138 (I76088,I76071,I76054);
not I_4139 (I75986,I76071);
DFFARX1 I_4140  ( .D(I65357), .CLK(I5694_clk), .RSTB(I76003_rst), .Q(I76119) );
not I_4141 (I76136,I76119);
nor I_4142 (I76153,I76071,I76136);
nand I_4143 (I75989,I76119,I76088);
DFFARX1 I_4144  ( .D(I76119), .CLK(I5694_clk), .RSTB(I76003_rst), .Q(I75971) );
nand I_4145 (I76198,I65366,I65384);
and I_4146 (I76215,I76198,I65378);
DFFARX1 I_4147  ( .D(I76215), .CLK(I5694_clk), .RSTB(I76003_rst), .Q(I76232) );
nor I_4148 (I75992,I76232,I76054);
nand I_4149 (I75983,I76232,I76153);
DFFARX1 I_4150  ( .D(I65369), .CLK(I5694_clk), .RSTB(I76003_rst), .Q(I76277) );
and I_4151 (I76294,I76277,I65363);
DFFARX1 I_4152  ( .D(I76294), .CLK(I5694_clk), .RSTB(I76003_rst), .Q(I76311) );
not I_4153 (I75974,I76311);
nand I_4154 (I76342,I76294,I76232);
and I_4155 (I76359,I76054,I76342);
DFFARX1 I_4156  ( .D(I76359), .CLK(I5694_clk), .RSTB(I76003_rst), .Q(I75965) );
DFFARX1 I_4157  ( .D(I65360), .CLK(I5694_clk), .RSTB(I76003_rst), .Q(I76390) );
nand I_4158 (I76407,I76390,I76054);
and I_4159 (I76424,I76232,I76407);
DFFARX1 I_4160  ( .D(I76424), .CLK(I5694_clk), .RSTB(I76003_rst), .Q(I75995) );
not I_4161 (I76455,I76390);
nor I_4162 (I76472,I76071,I76455);
and I_4163 (I76489,I76390,I76472);
or I_4164 (I76506,I76294,I76489);
DFFARX1 I_4165  ( .D(I76506), .CLK(I5694_clk), .RSTB(I76003_rst), .Q(I75980) );
nand I_4166 (I75977,I76390,I76136);
DFFARX1 I_4167  ( .D(I76390), .CLK(I5694_clk), .RSTB(I76003_rst), .Q(I75968) );
not I_4168 (I76598_rst,I5701);
nand I_4169 (I76615,I22428,I22416);
and I_4170 (I76632,I76615,I22422);
DFFARX1 I_4171  ( .D(I76632), .CLK(I5694_clk), .RSTB(I76598_rst), .Q(I76649) );
nor I_4172 (I76666,I22413,I22416);
nor I_4173 (I76683,I76666,I76649);
not I_4174 (I76581,I76666);
DFFARX1 I_4175  ( .D(I22398), .CLK(I5694_clk), .RSTB(I76598_rst), .Q(I76714) );
not I_4176 (I76731,I76714);
nor I_4177 (I76748,I76666,I76731);
nand I_4178 (I76584,I76714,I76683);
DFFARX1 I_4179  ( .D(I76714), .CLK(I5694_clk), .RSTB(I76598_rst), .Q(I76566) );
nand I_4180 (I76793,I22407,I22425);
and I_4181 (I76810,I76793,I22419);
DFFARX1 I_4182  ( .D(I76810), .CLK(I5694_clk), .RSTB(I76598_rst), .Q(I76827) );
nor I_4183 (I76587,I76827,I76649);
nand I_4184 (I76578,I76827,I76748);
DFFARX1 I_4185  ( .D(I22410), .CLK(I5694_clk), .RSTB(I76598_rst), .Q(I76872) );
and I_4186 (I76889,I76872,I22404);
DFFARX1 I_4187  ( .D(I76889), .CLK(I5694_clk), .RSTB(I76598_rst), .Q(I76906) );
not I_4188 (I76569,I76906);
nand I_4189 (I76937,I76889,I76827);
and I_4190 (I76954,I76649,I76937);
DFFARX1 I_4191  ( .D(I76954), .CLK(I5694_clk), .RSTB(I76598_rst), .Q(I76560) );
DFFARX1 I_4192  ( .D(I22401), .CLK(I5694_clk), .RSTB(I76598_rst), .Q(I76985) );
nand I_4193 (I77002,I76985,I76649);
and I_4194 (I77019,I76827,I77002);
DFFARX1 I_4195  ( .D(I77019), .CLK(I5694_clk), .RSTB(I76598_rst), .Q(I76590) );
not I_4196 (I77050,I76985);
nor I_4197 (I77067,I76666,I77050);
and I_4198 (I77084,I76985,I77067);
or I_4199 (I77101,I76889,I77084);
DFFARX1 I_4200  ( .D(I77101), .CLK(I5694_clk), .RSTB(I76598_rst), .Q(I76575) );
nand I_4201 (I76572,I76985,I76731);
DFFARX1 I_4202  ( .D(I76985), .CLK(I5694_clk), .RSTB(I76598_rst), .Q(I76563) );
not I_4203 (I77193_rst,I5701);
nand I_4204 (I77210,I33839,I33842);
and I_4205 (I77227,I77210,I33851);
DFFARX1 I_4206  ( .D(I77227), .CLK(I5694_clk), .RSTB(I77193_rst), .Q(I77244) );
nor I_4207 (I77261,I33845,I33842);
DFFARX1 I_4208  ( .D(I33866), .CLK(I5694_clk), .RSTB(I77193_rst), .Q(I77278) );
nand I_4209 (I77295,I77278,I77261);
DFFARX1 I_4210  ( .D(I77278), .CLK(I5694_clk), .RSTB(I77193_rst), .Q(I77164) );
nand I_4211 (I77326,I33863,I33869);
and I_4212 (I77343,I77326,I33854);
DFFARX1 I_4213  ( .D(I77343), .CLK(I5694_clk), .RSTB(I77193_rst), .Q(I77360) );
not I_4214 (I77377,I77360);
nor I_4215 (I77394,I77244,I77377);
and I_4216 (I77411,I77261,I77394);
and I_4217 (I77428,I77360,I77295);
DFFARX1 I_4218  ( .D(I77428), .CLK(I5694_clk), .RSTB(I77193_rst), .Q(I77161) );
DFFARX1 I_4219  ( .D(I77360), .CLK(I5694_clk), .RSTB(I77193_rst), .Q(I77155) );
DFFARX1 I_4220  ( .D(I33857), .CLK(I5694_clk), .RSTB(I77193_rst), .Q(I77473) );
and I_4221 (I77490,I77473,I33860);
nand I_4222 (I77507,I77490,I77360);
nor I_4223 (I77182,I77490,I77261);
not I_4224 (I77538,I77490);
nor I_4225 (I77555,I77244,I77538);
nand I_4226 (I77173,I77278,I77555);
nand I_4227 (I77167,I77360,I77538);
or I_4228 (I77600,I77490,I77411);
DFFARX1 I_4229  ( .D(I77600), .CLK(I5694_clk), .RSTB(I77193_rst), .Q(I77170) );
DFFARX1 I_4230  ( .D(I33848), .CLK(I5694_clk), .RSTB(I77193_rst), .Q(I77631) );
and I_4231 (I77648,I77631,I77507);
DFFARX1 I_4232  ( .D(I77648), .CLK(I5694_clk), .RSTB(I77193_rst), .Q(I77185) );
nor I_4233 (I77679,I77631,I77244);
nand I_4234 (I77179,I77490,I77679);
not I_4235 (I77176,I77631);
DFFARX1 I_4236  ( .D(I77631), .CLK(I5694_clk), .RSTB(I77193_rst), .Q(I77724) );
and I_4237 (I77158,I77631,I77724);
not I_4238 (I77788_rst,I5701);
nand I_4239 (I77805,I68327,I68342);
and I_4240 (I77822,I77805,I68339);
DFFARX1 I_4241  ( .D(I77822), .CLK(I5694_clk), .RSTB(I77788_rst), .Q(I77839) );
nor I_4242 (I77856,I68315,I68342);
DFFARX1 I_4243  ( .D(I68333), .CLK(I5694_clk), .RSTB(I77788_rst), .Q(I77873) );
nand I_4244 (I77890,I77873,I77856);
DFFARX1 I_4245  ( .D(I77873), .CLK(I5694_clk), .RSTB(I77788_rst), .Q(I77759) );
nand I_4246 (I77921,I68336,I68324);
and I_4247 (I77938,I77921,I68330);
DFFARX1 I_4248  ( .D(I77938), .CLK(I5694_clk), .RSTB(I77788_rst), .Q(I77955) );
not I_4249 (I77972,I77955);
nor I_4250 (I77989,I77839,I77972);
and I_4251 (I78006,I77856,I77989);
and I_4252 (I78023,I77955,I77890);
DFFARX1 I_4253  ( .D(I78023), .CLK(I5694_clk), .RSTB(I77788_rst), .Q(I77756) );
DFFARX1 I_4254  ( .D(I77955), .CLK(I5694_clk), .RSTB(I77788_rst), .Q(I77750) );
DFFARX1 I_4255  ( .D(I68321), .CLK(I5694_clk), .RSTB(I77788_rst), .Q(I78068) );
and I_4256 (I78085,I78068,I68345);
nand I_4257 (I78102,I78085,I77955);
nor I_4258 (I77777,I78085,I77856);
not I_4259 (I78133,I78085);
nor I_4260 (I78150,I77839,I78133);
nand I_4261 (I77768,I77873,I78150);
nand I_4262 (I77762,I77955,I78133);
or I_4263 (I78195,I78085,I78006);
DFFARX1 I_4264  ( .D(I78195), .CLK(I5694_clk), .RSTB(I77788_rst), .Q(I77765) );
DFFARX1 I_4265  ( .D(I68318), .CLK(I5694_clk), .RSTB(I77788_rst), .Q(I78226) );
and I_4266 (I78243,I78226,I78102);
DFFARX1 I_4267  ( .D(I78243), .CLK(I5694_clk), .RSTB(I77788_rst), .Q(I77780) );
nor I_4268 (I78274,I78226,I77839);
nand I_4269 (I77774,I78085,I78274);
not I_4270 (I77771,I78226);
DFFARX1 I_4271  ( .D(I78226), .CLK(I5694_clk), .RSTB(I77788_rst), .Q(I78319) );
and I_4272 (I77753,I78226,I78319);
not I_4273 (I78383_rst,I5701);
nand I_4274 (I78400,I24756,I24771);
and I_4275 (I78417,I78400,I24768);
DFFARX1 I_4276  ( .D(I78417), .CLK(I5694_clk), .RSTB(I78383_rst), .Q(I78434) );
nor I_4277 (I78451,I24744,I24771);
DFFARX1 I_4278  ( .D(I24762), .CLK(I5694_clk), .RSTB(I78383_rst), .Q(I78468) );
nand I_4279 (I78485,I78468,I78451);
DFFARX1 I_4280  ( .D(I78468), .CLK(I5694_clk), .RSTB(I78383_rst), .Q(I78354) );
nand I_4281 (I78516,I24765,I24753);
and I_4282 (I78533,I78516,I24759);
DFFARX1 I_4283  ( .D(I78533), .CLK(I5694_clk), .RSTB(I78383_rst), .Q(I78550) );
not I_4284 (I78567,I78550);
nor I_4285 (I78584,I78434,I78567);
and I_4286 (I78601,I78451,I78584);
and I_4287 (I78618,I78550,I78485);
DFFARX1 I_4288  ( .D(I78618), .CLK(I5694_clk), .RSTB(I78383_rst), .Q(I78351) );
DFFARX1 I_4289  ( .D(I78550), .CLK(I5694_clk), .RSTB(I78383_rst), .Q(I78345) );
DFFARX1 I_4290  ( .D(I24750), .CLK(I5694_clk), .RSTB(I78383_rst), .Q(I78663) );
and I_4291 (I78680,I78663,I24774);
nand I_4292 (I78697,I78680,I78550);
nor I_4293 (I78372,I78680,I78451);
not I_4294 (I78728,I78680);
nor I_4295 (I78745,I78434,I78728);
nand I_4296 (I78363,I78468,I78745);
nand I_4297 (I78357,I78550,I78728);
or I_4298 (I78790,I78680,I78601);
DFFARX1 I_4299  ( .D(I78790), .CLK(I5694_clk), .RSTB(I78383_rst), .Q(I78360) );
DFFARX1 I_4300  ( .D(I24747), .CLK(I5694_clk), .RSTB(I78383_rst), .Q(I78821) );
and I_4301 (I78838,I78821,I78697);
DFFARX1 I_4302  ( .D(I78838), .CLK(I5694_clk), .RSTB(I78383_rst), .Q(I78375) );
nor I_4303 (I78869,I78821,I78434);
nand I_4304 (I78369,I78680,I78869);
not I_4305 (I78366,I78821);
DFFARX1 I_4306  ( .D(I78821), .CLK(I5694_clk), .RSTB(I78383_rst), .Q(I78914) );
and I_4307 (I78348,I78821,I78914);
not I_4308 (I78978_rst,I5701);
nand I_4309 (I78995,I40224,I40200);
and I_4310 (I79012,I78995,I40209);
DFFARX1 I_4311  ( .D(I79012), .CLK(I5694_clk), .RSTB(I78978_rst), .Q(I79029) );
nor I_4312 (I79046,I40203,I40200);
DFFARX1 I_4313  ( .D(I40218), .CLK(I5694_clk), .RSTB(I78978_rst), .Q(I79063) );
nand I_4314 (I79080,I79063,I79046);
DFFARX1 I_4315  ( .D(I79063), .CLK(I5694_clk), .RSTB(I78978_rst), .Q(I78949) );
nand I_4316 (I79111,I40212,I40227);
and I_4317 (I79128,I79111,I40206);
DFFARX1 I_4318  ( .D(I79128), .CLK(I5694_clk), .RSTB(I78978_rst), .Q(I79145) );
not I_4319 (I79162,I79145);
nor I_4320 (I79179,I79029,I79162);
and I_4321 (I79196,I79046,I79179);
and I_4322 (I79213,I79145,I79080);
DFFARX1 I_4323  ( .D(I79213), .CLK(I5694_clk), .RSTB(I78978_rst), .Q(I78946) );
DFFARX1 I_4324  ( .D(I79145), .CLK(I5694_clk), .RSTB(I78978_rst), .Q(I78940) );
DFFARX1 I_4325  ( .D(I40197), .CLK(I5694_clk), .RSTB(I78978_rst), .Q(I79258) );
and I_4326 (I79275,I79258,I40215);
nand I_4327 (I79292,I79275,I79145);
nor I_4328 (I78967,I79275,I79046);
not I_4329 (I79323,I79275);
nor I_4330 (I79340,I79029,I79323);
nand I_4331 (I78958,I79063,I79340);
nand I_4332 (I78952,I79145,I79323);
or I_4333 (I79385,I79275,I79196);
DFFARX1 I_4334  ( .D(I79385), .CLK(I5694_clk), .RSTB(I78978_rst), .Q(I78955) );
DFFARX1 I_4335  ( .D(I40221), .CLK(I5694_clk), .RSTB(I78978_rst), .Q(I79416) );
and I_4336 (I79433,I79416,I79292);
DFFARX1 I_4337  ( .D(I79433), .CLK(I5694_clk), .RSTB(I78978_rst), .Q(I78970) );
nor I_4338 (I79464,I79416,I79029);
nand I_4339 (I78964,I79275,I79464);
not I_4340 (I78961,I79416);
DFFARX1 I_4341  ( .D(I79416), .CLK(I5694_clk), .RSTB(I78978_rst), .Q(I79509) );
and I_4342 (I78943,I79416,I79509);
not I_4343 (I79573_rst,I5701);
nand I_4344 (I79590,I27139,I27124);
and I_4345 (I79607,I79590,I27130);
DFFARX1 I_4346  ( .D(I79607), .CLK(I5694_clk), .RSTB(I79573_rst), .Q(I79624) );
nor I_4347 (I79641,I27133,I27124);
DFFARX1 I_4348  ( .D(I27145), .CLK(I5694_clk), .RSTB(I79573_rst), .Q(I79658) );
nand I_4349 (I79675,I79658,I79641);
DFFARX1 I_4350  ( .D(I79658), .CLK(I5694_clk), .RSTB(I79573_rst), .Q(I79544) );
nand I_4351 (I79706,I27136,I27127);
and I_4352 (I79723,I79706,I27154);
DFFARX1 I_4353  ( .D(I79723), .CLK(I5694_clk), .RSTB(I79573_rst), .Q(I79740) );
not I_4354 (I79757,I79740);
nor I_4355 (I79774,I79624,I79757);
and I_4356 (I79791,I79641,I79774);
and I_4357 (I79808,I79740,I79675);
DFFARX1 I_4358  ( .D(I79808), .CLK(I5694_clk), .RSTB(I79573_rst), .Q(I79541) );
DFFARX1 I_4359  ( .D(I79740), .CLK(I5694_clk), .RSTB(I79573_rst), .Q(I79535) );
DFFARX1 I_4360  ( .D(I27142), .CLK(I5694_clk), .RSTB(I79573_rst), .Q(I79853) );
and I_4361 (I79870,I79853,I27148);
nand I_4362 (I79887,I79870,I79740);
nor I_4363 (I79562,I79870,I79641);
not I_4364 (I79918,I79870);
nor I_4365 (I79935,I79624,I79918);
nand I_4366 (I79553,I79658,I79935);
nand I_4367 (I79547,I79740,I79918);
or I_4368 (I79980,I79870,I79791);
DFFARX1 I_4369  ( .D(I79980), .CLK(I5694_clk), .RSTB(I79573_rst), .Q(I79550) );
DFFARX1 I_4370  ( .D(I27151), .CLK(I5694_clk), .RSTB(I79573_rst), .Q(I80011) );
and I_4371 (I80028,I80011,I79887);
DFFARX1 I_4372  ( .D(I80028), .CLK(I5694_clk), .RSTB(I79573_rst), .Q(I79565) );
nor I_4373 (I80059,I80011,I79624);
nand I_4374 (I79559,I79870,I80059);
not I_4375 (I79556,I80011);
DFFARX1 I_4376  ( .D(I80011), .CLK(I5694_clk), .RSTB(I79573_rst), .Q(I80104) );
and I_4377 (I79538,I80011,I80104);
not I_4378 (I80168_rst,I5701);
nand I_4379 (I80185,I6853,I6829);
and I_4380 (I80202,I80185,I6838);
DFFARX1 I_4381  ( .D(I80202), .CLK(I5694_clk), .RSTB(I80168_rst), .Q(I80219) );
nor I_4382 (I80236,I6832,I6829);
DFFARX1 I_4383  ( .D(I6847), .CLK(I5694_clk), .RSTB(I80168_rst), .Q(I80253) );
nand I_4384 (I80270,I80253,I80236);
DFFARX1 I_4385  ( .D(I80253), .CLK(I5694_clk), .RSTB(I80168_rst), .Q(I80139) );
nand I_4386 (I80301,I6841,I6856);
and I_4387 (I80318,I80301,I6835);
DFFARX1 I_4388  ( .D(I80318), .CLK(I5694_clk), .RSTB(I80168_rst), .Q(I80335) );
not I_4389 (I80352,I80335);
nor I_4390 (I80369,I80219,I80352);
and I_4391 (I80386,I80236,I80369);
and I_4392 (I80403,I80335,I80270);
DFFARX1 I_4393  ( .D(I80403), .CLK(I5694_clk), .RSTB(I80168_rst), .Q(I80136) );
DFFARX1 I_4394  ( .D(I80335), .CLK(I5694_clk), .RSTB(I80168_rst), .Q(I80130) );
DFFARX1 I_4395  ( .D(I6826), .CLK(I5694_clk), .RSTB(I80168_rst), .Q(I80448) );
and I_4396 (I80465,I80448,I6844);
nand I_4397 (I80482,I80465,I80335);
nor I_4398 (I80157,I80465,I80236);
not I_4399 (I80513,I80465);
nor I_4400 (I80530,I80219,I80513);
nand I_4401 (I80148,I80253,I80530);
nand I_4402 (I80142,I80335,I80513);
or I_4403 (I80575,I80465,I80386);
DFFARX1 I_4404  ( .D(I80575), .CLK(I5694_clk), .RSTB(I80168_rst), .Q(I80145) );
DFFARX1 I_4405  ( .D(I6850), .CLK(I5694_clk), .RSTB(I80168_rst), .Q(I80606) );
and I_4406 (I80623,I80606,I80482);
DFFARX1 I_4407  ( .D(I80623), .CLK(I5694_clk), .RSTB(I80168_rst), .Q(I80160) );
nor I_4408 (I80654,I80606,I80219);
nand I_4409 (I80154,I80465,I80654);
not I_4410 (I80151,I80606);
DFFARX1 I_4411  ( .D(I80606), .CLK(I5694_clk), .RSTB(I80168_rst), .Q(I80699) );
and I_4412 (I80133,I80606,I80699);
not I_4413 (I80763_rst,I5701);
nand I_4414 (I80780,I20546,I20558);
and I_4415 (I80797,I80780,I20549);
DFFARX1 I_4416  ( .D(I80797), .CLK(I5694_clk), .RSTB(I80763_rst), .Q(I80814) );
nor I_4417 (I80831,I20543,I20558);
DFFARX1 I_4418  ( .D(I20534), .CLK(I5694_clk), .RSTB(I80763_rst), .Q(I80848) );
nand I_4419 (I80865,I80848,I80831);
DFFARX1 I_4420  ( .D(I80848), .CLK(I5694_clk), .RSTB(I80763_rst), .Q(I80734) );
nand I_4421 (I80896,I20540,I20531);
and I_4422 (I80913,I80896,I20537);
DFFARX1 I_4423  ( .D(I80913), .CLK(I5694_clk), .RSTB(I80763_rst), .Q(I80930) );
not I_4424 (I80947,I80930);
nor I_4425 (I80964,I80814,I80947);
and I_4426 (I80981,I80831,I80964);
and I_4427 (I80998,I80930,I80865);
DFFARX1 I_4428  ( .D(I80998), .CLK(I5694_clk), .RSTB(I80763_rst), .Q(I80731) );
DFFARX1 I_4429  ( .D(I80930), .CLK(I5694_clk), .RSTB(I80763_rst), .Q(I80725) );
DFFARX1 I_4430  ( .D(I20552), .CLK(I5694_clk), .RSTB(I80763_rst), .Q(I81043) );
and I_4431 (I81060,I81043,I20528);
nand I_4432 (I81077,I81060,I80930);
nor I_4433 (I80752,I81060,I80831);
not I_4434 (I81108,I81060);
nor I_4435 (I81125,I80814,I81108);
nand I_4436 (I80743,I80848,I81125);
nand I_4437 (I80737,I80930,I81108);
or I_4438 (I81170,I81060,I80981);
DFFARX1 I_4439  ( .D(I81170), .CLK(I5694_clk), .RSTB(I80763_rst), .Q(I80740) );
DFFARX1 I_4440  ( .D(I20555), .CLK(I5694_clk), .RSTB(I80763_rst), .Q(I81201) );
and I_4441 (I81218,I81201,I81077);
DFFARX1 I_4442  ( .D(I81218), .CLK(I5694_clk), .RSTB(I80763_rst), .Q(I80755) );
nor I_4443 (I81249,I81201,I80814);
nand I_4444 (I80749,I81060,I81249);
not I_4445 (I80746,I81201);
DFFARX1 I_4446  ( .D(I81201), .CLK(I5694_clk), .RSTB(I80763_rst), .Q(I81294) );
and I_4447 (I80728,I81201,I81294);
not I_4448 (I81358_rst,I5701);
nand I_4449 (I81375,I48523,I48508);
and I_4450 (I81392,I81375,I48520);
DFFARX1 I_4451  ( .D(I81392), .CLK(I5694_clk), .RSTB(I81358_rst), .Q(I81409) );
nor I_4452 (I81426,I48511,I48508);
DFFARX1 I_4453  ( .D(I48502), .CLK(I5694_clk), .RSTB(I81358_rst), .Q(I81443) );
nand I_4454 (I81460,I81443,I81426);
DFFARX1 I_4455  ( .D(I81443), .CLK(I5694_clk), .RSTB(I81358_rst), .Q(I81329) );
nand I_4456 (I81491,I48493,I48517);
and I_4457 (I81508,I81491,I48496);
DFFARX1 I_4458  ( .D(I81508), .CLK(I5694_clk), .RSTB(I81358_rst), .Q(I81525) );
not I_4459 (I81542,I81525);
nor I_4460 (I81559,I81409,I81542);
and I_4461 (I81576,I81426,I81559);
and I_4462 (I81593,I81525,I81460);
DFFARX1 I_4463  ( .D(I81593), .CLK(I5694_clk), .RSTB(I81358_rst), .Q(I81326) );
DFFARX1 I_4464  ( .D(I81525), .CLK(I5694_clk), .RSTB(I81358_rst), .Q(I81320) );
DFFARX1 I_4465  ( .D(I48514), .CLK(I5694_clk), .RSTB(I81358_rst), .Q(I81638) );
and I_4466 (I81655,I81638,I48499);
nand I_4467 (I81672,I81655,I81525);
nor I_4468 (I81347,I81655,I81426);
not I_4469 (I81703,I81655);
nor I_4470 (I81720,I81409,I81703);
nand I_4471 (I81338,I81443,I81720);
nand I_4472 (I81332,I81525,I81703);
or I_4473 (I81765,I81655,I81576);
DFFARX1 I_4474  ( .D(I81765), .CLK(I5694_clk), .RSTB(I81358_rst), .Q(I81335) );
DFFARX1 I_4475  ( .D(I48505), .CLK(I5694_clk), .RSTB(I81358_rst), .Q(I81796) );
and I_4476 (I81813,I81796,I81672);
DFFARX1 I_4477  ( .D(I81813), .CLK(I5694_clk), .RSTB(I81358_rst), .Q(I81350) );
nor I_4478 (I81844,I81796,I81409);
nand I_4479 (I81344,I81655,I81844);
not I_4480 (I81341,I81796);
DFFARX1 I_4481  ( .D(I81796), .CLK(I5694_clk), .RSTB(I81358_rst), .Q(I81889) );
and I_4482 (I81323,I81796,I81889);
not I_4483 (I81953_rst,I5701);
nand I_4484 (I81970,I9464,I9485);
and I_4485 (I81987,I81970,I9470);
DFFARX1 I_4486  ( .D(I81987), .CLK(I5694_clk), .RSTB(I81953_rst), .Q(I82004) );
nor I_4487 (I82021,I9488,I9485);
DFFARX1 I_4488  ( .D(I9491), .CLK(I5694_clk), .RSTB(I81953_rst), .Q(I82038) );
nand I_4489 (I82055,I82038,I82021);
DFFARX1 I_4490  ( .D(I82038), .CLK(I5694_clk), .RSTB(I81953_rst), .Q(I81924) );
nand I_4491 (I82086,I9461,I9473);
and I_4492 (I82103,I82086,I9482);
DFFARX1 I_4493  ( .D(I82103), .CLK(I5694_clk), .RSTB(I81953_rst), .Q(I82120) );
not I_4494 (I82137,I82120);
nor I_4495 (I82154,I82004,I82137);
and I_4496 (I82171,I82021,I82154);
and I_4497 (I82188,I82120,I82055);
DFFARX1 I_4498  ( .D(I82188), .CLK(I5694_clk), .RSTB(I81953_rst), .Q(I81921) );
DFFARX1 I_4499  ( .D(I82120), .CLK(I5694_clk), .RSTB(I81953_rst), .Q(I81915) );
DFFARX1 I_4500  ( .D(I9476), .CLK(I5694_clk), .RSTB(I81953_rst), .Q(I82233) );
and I_4501 (I82250,I82233,I9479);
nand I_4502 (I82267,I82250,I82120);
nor I_4503 (I81942,I82250,I82021);
not I_4504 (I82298,I82250);
nor I_4505 (I82315,I82004,I82298);
nand I_4506 (I81933,I82038,I82315);
nand I_4507 (I81927,I82120,I82298);
or I_4508 (I82360,I82250,I82171);
DFFARX1 I_4509  ( .D(I82360), .CLK(I5694_clk), .RSTB(I81953_rst), .Q(I81930) );
DFFARX1 I_4510  ( .D(I9467), .CLK(I5694_clk), .RSTB(I81953_rst), .Q(I82391) );
and I_4511 (I82408,I82391,I82267);
DFFARX1 I_4512  ( .D(I82408), .CLK(I5694_clk), .RSTB(I81953_rst), .Q(I81945) );
nor I_4513 (I82439,I82391,I82004);
nand I_4514 (I81939,I82250,I82439);
not I_4515 (I81936,I82391);
DFFARX1 I_4516  ( .D(I82391), .CLK(I5694_clk), .RSTB(I81953_rst), .Q(I82484) );
and I_4517 (I81918,I82391,I82484);
not I_4518 (I82548_rst,I5701);
not I_4519 (I82565,I77759);
nor I_4520 (I82582,I77762,I77771);
nand I_4521 (I82599,I82582,I77756);
nor I_4522 (I82616,I82565,I77762);
nand I_4523 (I82633,I82616,I77765);
not I_4524 (I82650,I77762);
not I_4525 (I82667,I82650);
not I_4526 (I82684,I77780);
nor I_4527 (I82701,I82684,I77768);
and I_4528 (I82718,I82701,I77753);
or I_4529 (I82735,I82718,I77750);
DFFARX1 I_4530  ( .D(I82735), .CLK(I5694_clk), .RSTB(I82548_rst), .Q(I82752) );
nand I_4531 (I82769,I82565,I77780);
or I_4532 (I82537,I82769,I82752);
not I_4533 (I82800,I82769);
nor I_4534 (I82817,I82752,I82800);
and I_4535 (I82834,I82650,I82817);
nand I_4536 (I82510,I82769,I82667);
DFFARX1 I_4537  ( .D(I77774), .CLK(I5694_clk), .RSTB(I82548_rst), .Q(I82865) );
or I_4538 (I82531,I82865,I82752);
nor I_4539 (I82896,I82865,I82633);
nor I_4540 (I82913,I82865,I82667);
nand I_4541 (I82516,I82599,I82913);
or I_4542 (I82944,I82865,I82834);
DFFARX1 I_4543  ( .D(I82944), .CLK(I5694_clk), .RSTB(I82548_rst), .Q(I82513) );
not I_4544 (I82519,I82865);
DFFARX1 I_4545  ( .D(I77777), .CLK(I5694_clk), .RSTB(I82548_rst), .Q(I82989) );
not I_4546 (I83006,I82989);
nor I_4547 (I83023,I83006,I82599);
DFFARX1 I_4548  ( .D(I83023), .CLK(I5694_clk), .RSTB(I82548_rst), .Q(I82525) );
nor I_4549 (I82540,I82865,I83006);
nor I_4550 (I82528,I83006,I82769);
not I_4551 (I83082,I83006);
and I_4552 (I83099,I82633,I83082);
nor I_4553 (I82534,I82769,I83099);
nand I_4554 (I82522,I83006,I82896);
not I_4555 (I83177_rst,I5701);
not I_4556 (I83194,I13321);
nor I_4557 (I83211,I13327,I13306);
nand I_4558 (I83228,I83211,I13312);
nor I_4559 (I83245,I83194,I13327);
nand I_4560 (I83262,I83245,I13318);
not I_4561 (I83279,I13327);
not I_4562 (I83296,I83279);
not I_4563 (I83313,I13315);
nor I_4564 (I83330,I83313,I13333);
and I_4565 (I83347,I83330,I13324);
or I_4566 (I83364,I83347,I13303);
DFFARX1 I_4567  ( .D(I83364), .CLK(I5694_clk), .RSTB(I83177_rst), .Q(I83381) );
nand I_4568 (I83398,I83194,I13315);
or I_4569 (I83166,I83398,I83381);
not I_4570 (I83429,I83398);
nor I_4571 (I83446,I83381,I83429);
and I_4572 (I83463,I83279,I83446);
nand I_4573 (I83139,I83398,I83296);
DFFARX1 I_4574  ( .D(I13330), .CLK(I5694_clk), .RSTB(I83177_rst), .Q(I83494) );
or I_4575 (I83160,I83494,I83381);
nor I_4576 (I83525,I83494,I83262);
nor I_4577 (I83542,I83494,I83296);
nand I_4578 (I83145,I83228,I83542);
or I_4579 (I83573,I83494,I83463);
DFFARX1 I_4580  ( .D(I83573), .CLK(I5694_clk), .RSTB(I83177_rst), .Q(I83142) );
not I_4581 (I83148,I83494);
DFFARX1 I_4582  ( .D(I13309), .CLK(I5694_clk), .RSTB(I83177_rst), .Q(I83618) );
not I_4583 (I83635,I83618);
nor I_4584 (I83652,I83635,I83228);
DFFARX1 I_4585  ( .D(I83652), .CLK(I5694_clk), .RSTB(I83177_rst), .Q(I83154) );
nor I_4586 (I83169,I83494,I83635);
nor I_4587 (I83157,I83635,I83398);
not I_4588 (I83711,I83635);
and I_4589 (I83728,I83262,I83711);
nor I_4590 (I83163,I83398,I83728);
nand I_4591 (I83151,I83635,I83525);
not I_4592 (I83806_rst,I5701);
not I_4593 (I83823,I72996);
nor I_4594 (I83840,I73014,I72993);
nand I_4595 (I83857,I83840,I73017);
nor I_4596 (I83874,I83823,I73014);
nand I_4597 (I83891,I83874,I73011);
not I_4598 (I83908,I73014);
not I_4599 (I83925,I83908);
not I_4600 (I83942,I73002);
nor I_4601 (I83959,I83942,I72990);
and I_4602 (I83976,I83959,I73008);
or I_4603 (I83993,I83976,I73020);
DFFARX1 I_4604  ( .D(I83993), .CLK(I5694_clk), .RSTB(I83806_rst), .Q(I84010) );
nand I_4605 (I84027,I83823,I73002);
or I_4606 (I83795,I84027,I84010);
not I_4607 (I84058,I84027);
nor I_4608 (I84075,I84010,I84058);
and I_4609 (I84092,I83908,I84075);
nand I_4610 (I83768,I84027,I83925);
DFFARX1 I_4611  ( .D(I72999), .CLK(I5694_clk), .RSTB(I83806_rst), .Q(I84123) );
or I_4612 (I83789,I84123,I84010);
nor I_4613 (I84154,I84123,I83891);
nor I_4614 (I84171,I84123,I83925);
nand I_4615 (I83774,I83857,I84171);
or I_4616 (I84202,I84123,I84092);
DFFARX1 I_4617  ( .D(I84202), .CLK(I5694_clk), .RSTB(I83806_rst), .Q(I83771) );
not I_4618 (I83777,I84123);
DFFARX1 I_4619  ( .D(I73005), .CLK(I5694_clk), .RSTB(I83806_rst), .Q(I84247) );
not I_4620 (I84264,I84247);
nor I_4621 (I84281,I84264,I83857);
DFFARX1 I_4622  ( .D(I84281), .CLK(I5694_clk), .RSTB(I83806_rst), .Q(I83783) );
nor I_4623 (I83798,I84123,I84264);
nor I_4624 (I83786,I84264,I84027);
not I_4625 (I84340,I84264);
and I_4626 (I84357,I83891,I84340);
nor I_4627 (I83792,I84027,I84357);
nand I_4628 (I83780,I84264,I84154);
not I_4629 (I84435_rst,I5701);
not I_4630 (I84452,I78949);
nor I_4631 (I84469,I78952,I78961);
nand I_4632 (I84486,I84469,I78946);
nor I_4633 (I84503,I84452,I78952);
nand I_4634 (I84520,I84503,I78955);
not I_4635 (I84537,I78952);
not I_4636 (I84554,I84537);
not I_4637 (I84571,I78970);
nor I_4638 (I84588,I84571,I78958);
and I_4639 (I84605,I84588,I78943);
or I_4640 (I84622,I84605,I78940);
DFFARX1 I_4641  ( .D(I84622), .CLK(I5694_clk), .RSTB(I84435_rst), .Q(I84639) );
nand I_4642 (I84656,I84452,I78970);
or I_4643 (I84424,I84656,I84639);
not I_4644 (I84687,I84656);
nor I_4645 (I84704,I84639,I84687);
and I_4646 (I84721,I84537,I84704);
nand I_4647 (I84397,I84656,I84554);
DFFARX1 I_4648  ( .D(I78964), .CLK(I5694_clk), .RSTB(I84435_rst), .Q(I84752) );
or I_4649 (I84418,I84752,I84639);
nor I_4650 (I84783,I84752,I84520);
nor I_4651 (I84800,I84752,I84554);
nand I_4652 (I84403,I84486,I84800);
or I_4653 (I84831,I84752,I84721);
DFFARX1 I_4654  ( .D(I84831), .CLK(I5694_clk), .RSTB(I84435_rst), .Q(I84400) );
not I_4655 (I84406,I84752);
DFFARX1 I_4656  ( .D(I78967), .CLK(I5694_clk), .RSTB(I84435_rst), .Q(I84876) );
not I_4657 (I84893,I84876);
nor I_4658 (I84910,I84893,I84486);
DFFARX1 I_4659  ( .D(I84910), .CLK(I5694_clk), .RSTB(I84435_rst), .Q(I84412) );
nor I_4660 (I84427,I84752,I84893);
nor I_4661 (I84415,I84893,I84656);
not I_4662 (I84969,I84893);
and I_4663 (I84986,I84520,I84969);
nor I_4664 (I84421,I84656,I84986);
nand I_4665 (I84409,I84893,I84783);
not I_4666 (I85064_rst,I5701);
not I_4667 (I85081,I63437);
nor I_4668 (I85098,I63446,I63449);
nand I_4669 (I85115,I85098,I63434);
nor I_4670 (I85132,I85081,I63446);
nand I_4671 (I85149,I85132,I63431);
not I_4672 (I85166,I63446);
not I_4673 (I85183,I85166);
not I_4674 (I85200,I63419);
nor I_4675 (I85217,I85200,I63425);
and I_4676 (I85234,I85217,I63422);
or I_4677 (I85251,I85234,I63443);
DFFARX1 I_4678  ( .D(I85251), .CLK(I5694_clk), .RSTB(I85064_rst), .Q(I85268) );
nand I_4679 (I85285,I85081,I63419);
or I_4680 (I85053,I85285,I85268);
not I_4681 (I85316,I85285);
nor I_4682 (I85333,I85268,I85316);
and I_4683 (I85350,I85166,I85333);
nand I_4684 (I85026,I85285,I85183);
DFFARX1 I_4685  ( .D(I63428), .CLK(I5694_clk), .RSTB(I85064_rst), .Q(I85381) );
or I_4686 (I85047,I85381,I85268);
nor I_4687 (I85412,I85381,I85149);
nor I_4688 (I85429,I85381,I85183);
nand I_4689 (I85032,I85115,I85429);
or I_4690 (I85460,I85381,I85350);
DFFARX1 I_4691  ( .D(I85460), .CLK(I5694_clk), .RSTB(I85064_rst), .Q(I85029) );
not I_4692 (I85035,I85381);
DFFARX1 I_4693  ( .D(I63440), .CLK(I5694_clk), .RSTB(I85064_rst), .Q(I85505) );
not I_4694 (I85522,I85505);
nor I_4695 (I85539,I85522,I85115);
DFFARX1 I_4696  ( .D(I85539), .CLK(I5694_clk), .RSTB(I85064_rst), .Q(I85041) );
nor I_4697 (I85056,I85381,I85522);
nor I_4698 (I85044,I85522,I85285);
not I_4699 (I85598,I85522);
and I_4700 (I85615,I85149,I85598);
nor I_4701 (I85050,I85285,I85615);
nand I_4702 (I85038,I85522,I85412);
not I_4703 (I85693_rst,I5701);
not I_4704 (I85710,I76566);
nor I_4705 (I85727,I76584,I76563);
nand I_4706 (I85744,I85727,I76587);
nor I_4707 (I85761,I85710,I76584);
nand I_4708 (I85778,I85761,I76581);
not I_4709 (I85795,I76584);
not I_4710 (I85812,I85795);
not I_4711 (I85829,I76572);
nor I_4712 (I85846,I85829,I76560);
and I_4713 (I85863,I85846,I76578);
or I_4714 (I85880,I85863,I76590);
DFFARX1 I_4715  ( .D(I85880), .CLK(I5694_clk), .RSTB(I85693_rst), .Q(I85897) );
nand I_4716 (I85914,I85710,I76572);
or I_4717 (I85682,I85914,I85897);
not I_4718 (I85945,I85914);
nor I_4719 (I85962,I85897,I85945);
and I_4720 (I85979,I85795,I85962);
nand I_4721 (I85655,I85914,I85812);
DFFARX1 I_4722  ( .D(I76569), .CLK(I5694_clk), .RSTB(I85693_rst), .Q(I86010) );
or I_4723 (I85676,I86010,I85897);
nor I_4724 (I86041,I86010,I85778);
nor I_4725 (I86058,I86010,I85812);
nand I_4726 (I85661,I85744,I86058);
or I_4727 (I86089,I86010,I85979);
DFFARX1 I_4728  ( .D(I86089), .CLK(I5694_clk), .RSTB(I85693_rst), .Q(I85658) );
not I_4729 (I85664,I86010);
DFFARX1 I_4730  ( .D(I76575), .CLK(I5694_clk), .RSTB(I85693_rst), .Q(I86134) );
not I_4731 (I86151,I86134);
nor I_4732 (I86168,I86151,I85744);
DFFARX1 I_4733  ( .D(I86168), .CLK(I5694_clk), .RSTB(I85693_rst), .Q(I85670) );
nor I_4734 (I85685,I86010,I86151);
nor I_4735 (I85673,I86151,I85914);
not I_4736 (I86227,I86151);
and I_4737 (I86244,I85778,I86227);
nor I_4738 (I85679,I85914,I86244);
nand I_4739 (I85667,I86151,I86041);
not I_4740 (I86322_rst,I5701);
not I_4741 (I86339,I67767);
nor I_4742 (I86356,I67740,I67758);
nand I_4743 (I86373,I86356,I67743);
nor I_4744 (I86390,I86339,I67740);
nand I_4745 (I86407,I86390,I67761);
not I_4746 (I86424,I67740);
not I_4747 (I86441,I86424);
not I_4748 (I86458,I67737);
nor I_4749 (I86475,I86458,I67764);
and I_4750 (I86492,I86475,I67755);
or I_4751 (I86509,I86492,I67746);
DFFARX1 I_4752  ( .D(I86509), .CLK(I5694_clk), .RSTB(I86322_rst), .Q(I86526) );
nand I_4753 (I86543,I86339,I67737);
or I_4754 (I86311,I86543,I86526);
not I_4755 (I86574,I86543);
nor I_4756 (I86591,I86526,I86574);
and I_4757 (I86608,I86424,I86591);
nand I_4758 (I86284,I86543,I86441);
DFFARX1 I_4759  ( .D(I67749), .CLK(I5694_clk), .RSTB(I86322_rst), .Q(I86639) );
or I_4760 (I86305,I86639,I86526);
nor I_4761 (I86670,I86639,I86407);
nor I_4762 (I86687,I86639,I86441);
nand I_4763 (I86290,I86373,I86687);
or I_4764 (I86718,I86639,I86608);
DFFARX1 I_4765  ( .D(I86718), .CLK(I5694_clk), .RSTB(I86322_rst), .Q(I86287) );
not I_4766 (I86293,I86639);
DFFARX1 I_4767  ( .D(I67752), .CLK(I5694_clk), .RSTB(I86322_rst), .Q(I86763) );
not I_4768 (I86780,I86763);
nor I_4769 (I86797,I86780,I86373);
DFFARX1 I_4770  ( .D(I86797), .CLK(I5694_clk), .RSTB(I86322_rst), .Q(I86299) );
nor I_4771 (I86314,I86639,I86780);
nor I_4772 (I86302,I86780,I86543);
not I_4773 (I86856,I86780);
and I_4774 (I86873,I86407,I86856);
nor I_4775 (I86308,I86543,I86873);
nand I_4776 (I86296,I86780,I86670);
not I_4777 (I86951_rst,I5701);
not I_4778 (I86968,I79544);
nor I_4779 (I86985,I79547,I79556);
nand I_4780 (I87002,I86985,I79541);
nor I_4781 (I87019,I86968,I79547);
nand I_4782 (I87036,I87019,I79550);
not I_4783 (I87053,I79547);
not I_4784 (I87070,I87053);
not I_4785 (I87087,I79565);
nor I_4786 (I87104,I87087,I79553);
and I_4787 (I87121,I87104,I79538);
or I_4788 (I87138,I87121,I79535);
DFFARX1 I_4789  ( .D(I87138), .CLK(I5694_clk), .RSTB(I86951_rst), .Q(I87155) );
nand I_4790 (I87172,I86968,I79565);
or I_4791 (I86940,I87172,I87155);
not I_4792 (I87203,I87172);
nor I_4793 (I87220,I87155,I87203);
and I_4794 (I87237,I87053,I87220);
nand I_4795 (I86913,I87172,I87070);
DFFARX1 I_4796  ( .D(I79559), .CLK(I5694_clk), .RSTB(I86951_rst), .Q(I87268) );
or I_4797 (I86934,I87268,I87155);
nor I_4798 (I87299,I87268,I87036);
nor I_4799 (I87316,I87268,I87070);
nand I_4800 (I86919,I87002,I87316);
or I_4801 (I87347,I87268,I87237);
DFFARX1 I_4802  ( .D(I87347), .CLK(I5694_clk), .RSTB(I86951_rst), .Q(I86916) );
not I_4803 (I86922,I87268);
DFFARX1 I_4804  ( .D(I79562), .CLK(I5694_clk), .RSTB(I86951_rst), .Q(I87392) );
not I_4805 (I87409,I87392);
nor I_4806 (I87426,I87409,I87002);
DFFARX1 I_4807  ( .D(I87426), .CLK(I5694_clk), .RSTB(I86951_rst), .Q(I86928) );
nor I_4808 (I86943,I87268,I87409);
nor I_4809 (I86931,I87409,I87172);
not I_4810 (I87485,I87409);
and I_4811 (I87502,I87036,I87485);
nor I_4812 (I86937,I87172,I87502);
nand I_4813 (I86925,I87409,I87299);
not I_4814 (I87580_rst,I5701);
not I_4815 (I87597,I70079);
nor I_4816 (I87614,I70052,I70070);
nand I_4817 (I87631,I87614,I70055);
nor I_4818 (I87648,I87597,I70052);
nand I_4819 (I87665,I87648,I70073);
not I_4820 (I87682,I70052);
not I_4821 (I87699,I87682);
not I_4822 (I87716,I70049);
nor I_4823 (I87733,I87716,I70076);
and I_4824 (I87750,I87733,I70067);
or I_4825 (I87767,I87750,I70058);
DFFARX1 I_4826  ( .D(I87767), .CLK(I5694_clk), .RSTB(I87580_rst), .Q(I87784) );
nand I_4827 (I87801,I87597,I70049);
or I_4828 (I87569,I87801,I87784);
not I_4829 (I87832,I87801);
nor I_4830 (I87849,I87784,I87832);
and I_4831 (I87866,I87682,I87849);
nand I_4832 (I87542,I87801,I87699);
DFFARX1 I_4833  ( .D(I70061), .CLK(I5694_clk), .RSTB(I87580_rst), .Q(I87897) );
or I_4834 (I87563,I87897,I87784);
nor I_4835 (I87928,I87897,I87665);
nor I_4836 (I87945,I87897,I87699);
nand I_4837 (I87548,I87631,I87945);
or I_4838 (I87976,I87897,I87866);
DFFARX1 I_4839  ( .D(I87976), .CLK(I5694_clk), .RSTB(I87580_rst), .Q(I87545) );
not I_4840 (I87551,I87897);
DFFARX1 I_4841  ( .D(I70064), .CLK(I5694_clk), .RSTB(I87580_rst), .Q(I88021) );
not I_4842 (I88038,I88021);
nor I_4843 (I88055,I88038,I87631);
DFFARX1 I_4844  ( .D(I88055), .CLK(I5694_clk), .RSTB(I87580_rst), .Q(I87557) );
nor I_4845 (I87572,I87897,I88038);
nor I_4846 (I87560,I88038,I87801);
not I_4847 (I88114,I88038);
and I_4848 (I88131,I87665,I88114);
nor I_4849 (I87566,I87801,I88131);
nand I_4850 (I87554,I88038,I87928);
not I_4851 (I88209_rst,I5701);
not I_4852 (I88226,I46057);
nor I_4853 (I88243,I46048,I46072);
nand I_4854 (I88260,I88243,I46075);
nor I_4855 (I88277,I88226,I46048);
nand I_4856 (I88294,I88277,I46066);
not I_4857 (I88311,I46048);
not I_4858 (I88328,I88311);
not I_4859 (I88345,I46060);
nor I_4860 (I8836_rst2,I88345,I46054);
and I_4861 (I88379,I8836_rst2,I46063);
or I_4862 (I88396,I88379,I46051);
DFFARX1 I_4863  ( .D(I88396), .CLK(I5694_clk), .RSTB(I88209_rst), .Q(I88413) );
nand I_4864 (I88430,I88226,I46060);
or I_4865 (I88198,I88430,I88413);
not I_4866 (I88461,I88430);
nor I_4867 (I88478,I88413,I88461);
and I_4868 (I88495,I88311,I88478);
nand I_4869 (I88171,I88430,I88328);
DFFARX1 I_4870  ( .D(I46045), .CLK(I5694_clk), .RSTB(I88209_rst), .Q(I88526) );
or I_4871 (I88192,I88526,I88413);
nor I_4872 (I88557,I88526,I88294);
nor I_4873 (I88574,I88526,I88328);
nand I_4874 (I88177,I88260,I88574);
or I_4875 (I88605,I88526,I88495);
DFFARX1 I_4876  ( .D(I88605), .CLK(I5694_clk), .RSTB(I88209_rst), .Q(I88174) );
not I_4877 (I88180,I88526);
DFFARX1 I_4878  ( .D(I46069), .CLK(I5694_clk), .RSTB(I88209_rst), .Q(I88650) );
not I_4879 (I88667,I88650);
nor I_4880 (I88684,I88667,I88260);
DFFARX1 I_4881  ( .D(I88684), .CLK(I5694_clk), .RSTB(I88209_rst), .Q(I88186) );
nor I_4882 (I88201,I88526,I88667);
nor I_4883 (I88189,I88667,I88430);
not I_4884 (I88743,I88667);
and I_4885 (I88760,I88294,I88743);
nor I_4886 (I88195,I88430,I88760);
nand I_4887 (I88183,I88667,I88557);
not I_4888 (I88838_rst,I5701);
not I_4889 (I88855,I39557);
nor I_4890 (I88872,I39575,I39554);
nand I_4891 (I88889,I88872,I39572);
nor I_4892 (I88906,I88855,I39575);
nand I_4893 (I88923,I88906,I39566);
not I_4894 (I88940,I39575);
not I_4895 (I88957,I88940);
not I_4896 (I88974,I39569);
nor I_4897 (I88991,I88974,I39563);
and I_4898 (I89008,I88991,I39560);
or I_4899 (I89025,I89008,I39551);
DFFARX1 I_4900  ( .D(I89025), .CLK(I5694_clk), .RSTB(I88838_rst), .Q(I89042) );
nand I_4901 (I89059,I88855,I39569);
or I_4902 (I88827,I89059,I89042);
not I_4903 (I89090,I89059);
nor I_4904 (I89107,I89042,I89090);
and I_4905 (I89124,I88940,I89107);
nand I_4906 (I88800,I89059,I88957);
DFFARX1 I_4907  ( .D(I39581), .CLK(I5694_clk), .RSTB(I88838_rst), .Q(I89155) );
or I_4908 (I88821,I89155,I89042);
nor I_4909 (I89186,I89155,I88923);
nor I_4910 (I89203,I89155,I88957);
nand I_4911 (I88806,I88889,I89203);
or I_4912 (I89234,I89155,I89124);
DFFARX1 I_4913  ( .D(I89234), .CLK(I5694_clk), .RSTB(I88838_rst), .Q(I88803) );
not I_4914 (I88809,I89155);
DFFARX1 I_4915  ( .D(I39578), .CLK(I5694_clk), .RSTB(I88838_rst), .Q(I89279) );
not I_4916 (I89296,I89279);
nor I_4917 (I89313,I89296,I88889);
DFFARX1 I_4918  ( .D(I89313), .CLK(I5694_clk), .RSTB(I88838_rst), .Q(I88815) );
nor I_4919 (I88830,I89155,I89296);
nor I_4920 (I88818,I89296,I89059);
not I_4921 (I89372,I89296);
and I_4922 (I89389,I88923,I89372);
nor I_4923 (I88824,I89059,I89389);
nand I_4924 (I88812,I89296,I89186);
not I_4925 (I89467_rst,I5701);
not I_4926 (I89484,I65975);
nor I_4927 (I89501,I65999,I65978);
nand I_4928 (I89518,I89501,I65984);
nor I_4929 (I89535,I89484,I65999);
nand I_4930 (I89552,I89535,I65996);
not I_4931 (I89569,I65999);
not I_4932 (I89586,I89569);
not I_4933 (I89603,I65993);
nor I_4934 (I89620,I89603,I65972);
and I_4935 (I89637,I89620,I65969);
or I_4936 (I89654,I89637,I65981);
DFFARX1 I_4937  ( .D(I89654), .CLK(I5694_clk), .RSTB(I89467_rst), .Q(I89671) );
nand I_4938 (I89688,I89484,I65993);
or I_4939 (I89456,I89688,I89671);
not I_4940 (I89719,I89688);
nor I_4941 (I89736,I89671,I89719);
and I_4942 (I89753,I89569,I89736);
nand I_4943 (I89429,I89688,I89586);
DFFARX1 I_4944  ( .D(I65987), .CLK(I5694_clk), .RSTB(I89467_rst), .Q(I89784) );
or I_4945 (I89450,I89784,I89671);
nor I_4946 (I89815,I89784,I89552);
nor I_4947 (I89832,I89784,I89586);
nand I_4948 (I89435,I89518,I89832);
or I_4949 (I89863,I89784,I89753);
DFFARX1 I_4950  ( .D(I89863), .CLK(I5694_clk), .RSTB(I89467_rst), .Q(I89432) );
not I_4951 (I89438,I89784);
DFFARX1 I_4952  ( .D(I65990), .CLK(I5694_clk), .RSTB(I89467_rst), .Q(I89908) );
not I_4953 (I89925,I89908);
nor I_4954 (I89942,I89925,I89518);
DFFARX1 I_4955  ( .D(I89942), .CLK(I5694_clk), .RSTB(I89467_rst), .Q(I89444) );
nor I_4956 (I89459,I89784,I89925);
nor I_4957 (I89447,I89925,I89688);
not I_4958 (I90001,I89925);
and I_4959 (I90018,I89552,I90001);
nor I_4960 (I89453,I89688,I90018);
nand I_4961 (I89441,I89925,I89815);
not I_4962 (I90096_rst,I5701);
not I_4963 (I90113,I51027);
nor I_4964 (I90130,I51033,I51012);
nand I_4965 (I90147,I90130,I51018);
nor I_4966 (I90164,I90113,I51033);
nand I_4967 (I90181,I90164,I51024);
not I_4968 (I90198,I51033);
not I_4969 (I90215,I90198);
not I_4970 (I90232,I51021);
nor I_4971 (I90249,I90232,I51039);
and I_4972 (I90266,I90249,I51030);
or I_4973 (I90283,I90266,I51009);
DFFARX1 I_4974  ( .D(I90283), .CLK(I5694_clk), .RSTB(I90096_rst), .Q(I90300) );
nand I_4975 (I90317,I90113,I51021);
or I_4976 (I90085,I90317,I90300);
not I_4977 (I90348,I90317);
nor I_4978 (I90365,I90300,I90348);
and I_4979 (I90382,I90198,I90365);
nand I_4980 (I90058,I90317,I90215);
DFFARX1 I_4981  ( .D(I51036), .CLK(I5694_clk), .RSTB(I90096_rst), .Q(I90413) );
or I_4982 (I90079,I90413,I90300);
nor I_4983 (I90444,I90413,I90181);
nor I_4984 (I90461,I90413,I90215);
nand I_4985 (I90064,I90147,I90461);
or I_4986 (I90492,I90413,I90382);
DFFARX1 I_4987  ( .D(I90492), .CLK(I5694_clk), .RSTB(I90096_rst), .Q(I90061) );
not I_4988 (I90067,I90413);
DFFARX1 I_4989  ( .D(I51015), .CLK(I5694_clk), .RSTB(I90096_rst), .Q(I90537) );
not I_4990 (I90554,I90537);
nor I_4991 (I90571,I90554,I90147);
DFFARX1 I_4992  ( .D(I90571), .CLK(I5694_clk), .RSTB(I90096_rst), .Q(I90073) );
nor I_4993 (I90088,I90413,I90554);
nor I_4994 (I90076,I90554,I90317);
not I_4995 (I90630,I90554);
and I_4996 (I90647,I90181,I90630);
nor I_4997 (I90082,I90317,I90647);
nand I_4998 (I90070,I90554,I90444);
not I_4999 (I90725_rst,I5701);
nand I_5000 (I90742,I74201,I74183);
and I_5001 (I90759,I90742,I74198);
DFFARX1 I_5002  ( .D(I90759), .CLK(I5694_clk), .RSTB(I90725_rst), .Q(I90776) );
not I_5003 (I90714,I90776);
DFFARX1 I_5004  ( .D(I90776), .CLK(I5694_clk), .RSTB(I90725_rst), .Q(I90807) );
not I_5005 (I90702,I90807);
nor I_5006 (I90838,I74189,I74183);
not I_5007 (I90855,I90838);
nor I_5008 (I90872,I90776,I90855);
DFFARX1 I_5009  ( .D(I74204), .CLK(I5694_clk), .RSTB(I90725_rst), .Q(I90889) );
not I_5010 (I90906,I90889);
nand I_5011 (I90705,I90889,I90855);
DFFARX1 I_5012  ( .D(I90889), .CLK(I5694_clk), .RSTB(I90725_rst), .Q(I90937) );
and I_5013 (I90690,I90776,I90937);
nand I_5014 (I90968,I74180,I74186);
and I_5015 (I90985,I90968,I74192);
DFFARX1 I_5016  ( .D(I90985), .CLK(I5694_clk), .RSTB(I90725_rst), .Q(I91002) );
nor I_5017 (I91019,I91002,I90906);
and I_5018 (I91036,I90838,I91019);
nor I_5019 (I91053,I91002,I90776);
DFFARX1 I_5020  ( .D(I91002), .CLK(I5694_clk), .RSTB(I90725_rst), .Q(I90696) );
DFFARX1 I_5021  ( .D(I74207), .CLK(I5694_clk), .RSTB(I90725_rst), .Q(I91084) );
and I_5022 (I91101,I91084,I74195);
or I_5023 (I91118,I91101,I91036);
DFFARX1 I_5024  ( .D(I91118), .CLK(I5694_clk), .RSTB(I90725_rst), .Q(I90708) );
nand I_5025 (I90717,I91101,I91053);
DFFARX1 I_5026  ( .D(I91101), .CLK(I5694_clk), .RSTB(I90725_rst), .Q(I90687) );
DFFARX1 I_5027  ( .D(I74210), .CLK(I5694_clk), .RSTB(I90725_rst), .Q(I91177) );
nand I_5028 (I90711,I91177,I90872);
DFFARX1 I_5029  ( .D(I91177), .CLK(I5694_clk), .RSTB(I90725_rst), .Q(I90699) );
nand I_5030 (I91222,I91177,I90838);
and I_5031 (I91239,I90889,I91222);
DFFARX1 I_5032  ( .D(I91239), .CLK(I5694_clk), .RSTB(I90725_rst), .Q(I90693) );
not I_5033 (I91303_rst,I5701);
nand I_5034 (I91320,I57623,I57626);
and I_5035 (I91337,I91320,I57605);
DFFARX1 I_5036  ( .D(I91337), .CLK(I5694_clk), .RSTB(I91303_rst), .Q(I91354) );
not I_5037 (I91292,I91354);
DFFARX1 I_5038  ( .D(I91354), .CLK(I5694_clk), .RSTB(I91303_rst), .Q(I91385) );
not I_5039 (I91280,I91385);
nor I_5040 (I91416,I57620,I57626);
not I_5041 (I91433,I91416);
nor I_5042 (I91450,I91354,I91433);
DFFARX1 I_5043  ( .D(I57629), .CLK(I5694_clk), .RSTB(I91303_rst), .Q(I91467) );
not I_5044 (I91484,I91467);
nand I_5045 (I91283,I91467,I91433);
DFFARX1 I_5046  ( .D(I91467), .CLK(I5694_clk), .RSTB(I91303_rst), .Q(I91515) );
and I_5047 (I91268,I91354,I91515);
nand I_5048 (I91546,I57617,I57635);
and I_5049 (I91563,I91546,I57611);
DFFARX1 I_5050  ( .D(I91563), .CLK(I5694_clk), .RSTB(I91303_rst), .Q(I91580) );
nor I_5051 (I91597,I91580,I91484);
and I_5052 (I91614,I91416,I91597);
nor I_5053 (I91631,I91580,I91354);
DFFARX1 I_5054  ( .D(I91580), .CLK(I5694_clk), .RSTB(I91303_rst), .Q(I91274) );
DFFARX1 I_5055  ( .D(I57608), .CLK(I5694_clk), .RSTB(I91303_rst), .Q(I91662) );
and I_5056 (I91679,I91662,I57614);
or I_5057 (I91696,I91679,I91614);
DFFARX1 I_5058  ( .D(I91696), .CLK(I5694_clk), .RSTB(I91303_rst), .Q(I91286) );
nand I_5059 (I91295,I91679,I91631);
DFFARX1 I_5060  ( .D(I91679), .CLK(I5694_clk), .RSTB(I91303_rst), .Q(I91265) );
DFFARX1 I_5061  ( .D(I57632), .CLK(I5694_clk), .RSTB(I91303_rst), .Q(I91755) );
nand I_5062 (I91289,I91755,I91450);
DFFARX1 I_5063  ( .D(I91755), .CLK(I5694_clk), .RSTB(I91303_rst), .Q(I91277) );
nand I_5064 (I91800,I91755,I91416);
and I_5065 (I91817,I91467,I91800);
DFFARX1 I_5066  ( .D(I91817), .CLK(I5694_clk), .RSTB(I91303_rst), .Q(I91271) );
not I_5067 (I91881_rst,I5701);
nand I_5068 (I91898,I40864,I40849);
and I_5069 (I91915,I91898,I40843);
DFFARX1 I_5070  ( .D(I91915), .CLK(I5694_clk), .RSTB(I91881_rst), .Q(I91932) );
not I_5071 (I91870,I91932);
DFFARX1 I_5072  ( .D(I91932), .CLK(I5694_clk), .RSTB(I91881_rst), .Q(I91963) );
not I_5073 (I91858,I91963);
nor I_5074 (I91994,I40870,I40849);
not I_5075 (I92011,I91994);
nor I_5076 (I92028,I91932,I92011);
DFFARX1 I_5077  ( .D(I40873), .CLK(I5694_clk), .RSTB(I91881_rst), .Q(I92045) );
not I_5078 (I92062,I92045);
nand I_5079 (I91861,I92045,I92011);
DFFARX1 I_5080  ( .D(I92045), .CLK(I5694_clk), .RSTB(I91881_rst), .Q(I92093) );
and I_5081 (I91846,I91932,I92093);
nand I_5082 (I92124,I40855,I40858);
and I_5083 (I92141,I92124,I40861);
DFFARX1 I_5084  ( .D(I92141), .CLK(I5694_clk), .RSTB(I91881_rst), .Q(I92158) );
nor I_5085 (I92175,I92158,I92062);
and I_5086 (I92192,I91994,I92175);
nor I_5087 (I92209,I92158,I91932);
DFFARX1 I_5088  ( .D(I92158), .CLK(I5694_clk), .RSTB(I91881_rst), .Q(I91852) );
DFFARX1 I_5089  ( .D(I40867), .CLK(I5694_clk), .RSTB(I91881_rst), .Q(I92240) );
and I_5090 (I92257,I92240,I40852);
or I_5091 (I92274,I92257,I92192);
DFFARX1 I_5092  ( .D(I92274), .CLK(I5694_clk), .RSTB(I91881_rst), .Q(I91864) );
nand I_5093 (I91873,I92257,I92209);
DFFARX1 I_5094  ( .D(I92257), .CLK(I5694_clk), .RSTB(I91881_rst), .Q(I91843) );
DFFARX1 I_5095  ( .D(I40846), .CLK(I5694_clk), .RSTB(I91881_rst), .Q(I92333) );
nand I_5096 (I91867,I92333,I92028);
DFFARX1 I_5097  ( .D(I92333), .CLK(I5694_clk), .RSTB(I91881_rst), .Q(I91855) );
nand I_5098 (I92378,I92333,I91994);
and I_5099 (I92395,I92045,I92378);
DFFARX1 I_5100  ( .D(I92395), .CLK(I5694_clk), .RSTB(I91881_rst), .Q(I91849) );
not I_5101 (I92459_rst,I5701);
nand I_5102 (I92476,I47907,I47904);
and I_5103 (I92493,I92476,I47916);
DFFARX1 I_5104  ( .D(I92493), .CLK(I5694_clk), .RSTB(I92459_rst), .Q(I92510) );
not I_5105 (I92448,I92510);
DFFARX1 I_5106  ( .D(I92510), .CLK(I5694_clk), .RSTB(I92459_rst), .Q(I92541) );
not I_5107 (I92436,I92541);
nor I_5108 (I92572,I47919,I47904);
not I_5109 (I92589,I92572);
nor I_5110 (I92606,I92510,I92589);
DFFARX1 I_5111  ( .D(I47925), .CLK(I5694_clk), .RSTB(I92459_rst), .Q(I92623) );
not I_5112 (I92640,I92623);
nand I_5113 (I92439,I92623,I92589);
DFFARX1 I_5114  ( .D(I92623), .CLK(I5694_clk), .RSTB(I92459_rst), .Q(I92671) );
and I_5115 (I92424,I92510,I92671);
nand I_5116 (I92702,I47898,I47901);
and I_5117 (I92719,I92702,I47910);
DFFARX1 I_5118  ( .D(I92719), .CLK(I5694_clk), .RSTB(I92459_rst), .Q(I92736) );
nor I_5119 (I92753,I92736,I92640);
and I_5120 (I92770,I92572,I92753);
nor I_5121 (I92787,I92736,I92510);
DFFARX1 I_5122  ( .D(I92736), .CLK(I5694_clk), .RSTB(I92459_rst), .Q(I92430) );
DFFARX1 I_5123  ( .D(I47928), .CLK(I5694_clk), .RSTB(I92459_rst), .Q(I92818) );
and I_5124 (I92835,I92818,I47922);
or I_5125 (I92852,I92835,I92770);
DFFARX1 I_5126  ( .D(I92852), .CLK(I5694_clk), .RSTB(I92459_rst), .Q(I92442) );
nand I_5127 (I92451,I92835,I92787);
DFFARX1 I_5128  ( .D(I92835), .CLK(I5694_clk), .RSTB(I92459_rst), .Q(I92421) );
DFFARX1 I_5129  ( .D(I47913), .CLK(I5694_clk), .RSTB(I92459_rst), .Q(I92911) );
nand I_5130 (I92445,I92911,I92606);
DFFARX1 I_5131  ( .D(I92911), .CLK(I5694_clk), .RSTB(I92459_rst), .Q(I92433) );
nand I_5132 (I92956,I92911,I92572);
and I_5133 (I92973,I92623,I92956);
DFFARX1 I_5134  ( .D(I92973), .CLK(I5694_clk), .RSTB(I92459_rst), .Q(I92427) );
not I_5135 (I93037_rst,I5701);
nand I_5136 (I93054,I39014,I38999);
and I_5137 (I93071,I93054,I39008);
DFFARX1 I_5138  ( .D(I93071), .CLK(I5694_clk), .RSTB(I93037_rst), .Q(I93088) );
not I_5139 (I93026,I93088);
DFFARX1 I_5140  ( .D(I93088), .CLK(I5694_clk), .RSTB(I93037_rst), .Q(I93119) );
not I_5141 (I93014,I93119);
nor I_5142 (I93150,I39020,I38999);
not I_5143 (I93167,I93150);
nor I_5144 (I93184,I93088,I93167);
DFFARX1 I_5145  ( .D(I39011), .CLK(I5694_clk), .RSTB(I93037_rst), .Q(I93201) );
not I_5146 (I93218,I93201);
nand I_5147 (I93017,I93201,I93167);
DFFARX1 I_5148  ( .D(I93201), .CLK(I5694_clk), .RSTB(I93037_rst), .Q(I93249) );
and I_5149 (I93002,I93088,I93249);
nand I_5150 (I93280,I38996,I38990);
and I_5151 (I93297,I93280,I39005);
DFFARX1 I_5152  ( .D(I93297), .CLK(I5694_clk), .RSTB(I93037_rst), .Q(I93314) );
nor I_5153 (I93331,I93314,I93218);
and I_5154 (I93348,I93150,I93331);
nor I_5155 (I93365,I93314,I93088);
DFFARX1 I_5156  ( .D(I93314), .CLK(I5694_clk), .RSTB(I93037_rst), .Q(I93008) );
DFFARX1 I_5157  ( .D(I38993), .CLK(I5694_clk), .RSTB(I93037_rst), .Q(I93396) );
and I_5158 (I93413,I93396,I39017);
or I_5159 (I93430,I93413,I93348);
DFFARX1 I_5160  ( .D(I93430), .CLK(I5694_clk), .RSTB(I93037_rst), .Q(I93020) );
nand I_5161 (I93029,I93413,I93365);
DFFARX1 I_5162  ( .D(I93413), .CLK(I5694_clk), .RSTB(I93037_rst), .Q(I92999) );
DFFARX1 I_5163  ( .D(I39002), .CLK(I5694_clk), .RSTB(I93037_rst), .Q(I93489) );
nand I_5164 (I93023,I93489,I93184);
DFFARX1 I_5165  ( .D(I93489), .CLK(I5694_clk), .RSTB(I93037_rst), .Q(I93011) );
nand I_5166 (I93534,I93489,I93150);
and I_5167 (I93551,I93201,I93534);
DFFARX1 I_5168  ( .D(I93551), .CLK(I5694_clk), .RSTB(I93037_rst), .Q(I93005) );
not I_5169 (I93615_rst,I5701);
nand I_5170 (I93632,I17290,I17287);
and I_5171 (I93649,I93632,I17311);
DFFARX1 I_5172  ( .D(I93649), .CLK(I5694_clk), .RSTB(I93615_rst), .Q(I93666) );
not I_5173 (I93604,I93666);
DFFARX1 I_5174  ( .D(I93666), .CLK(I5694_clk), .RSTB(I93615_rst), .Q(I93697) );
not I_5175 (I93592,I93697);
nor I_5176 (I93728,I17293,I17287);
not I_5177 (I93745,I93728);
nor I_5178 (I93762,I93666,I93745);
DFFARX1 I_5179  ( .D(I17308), .CLK(I5694_clk), .RSTB(I93615_rst), .Q(I93779) );
not I_5180 (I93796,I93779);
nand I_5181 (I93595,I93779,I93745);
DFFARX1 I_5182  ( .D(I93779), .CLK(I5694_clk), .RSTB(I93615_rst), .Q(I93827) );
and I_5183 (I93580,I93666,I93827);
nand I_5184 (I93858,I17296,I17281);
and I_5185 (I93875,I93858,I17299);
DFFARX1 I_5186  ( .D(I93875), .CLK(I5694_clk), .RSTB(I93615_rst), .Q(I93892) );
nor I_5187 (I93909,I93892,I93796);
and I_5188 (I93926,I93728,I93909);
nor I_5189 (I93943,I93892,I93666);
DFFARX1 I_5190  ( .D(I93892), .CLK(I5694_clk), .RSTB(I93615_rst), .Q(I93586) );
DFFARX1 I_5191  ( .D(I17302), .CLK(I5694_clk), .RSTB(I93615_rst), .Q(I93974) );
and I_5192 (I93991,I93974,I17305);
or I_5193 (I94008,I93991,I93926);
DFFARX1 I_5194  ( .D(I94008), .CLK(I5694_clk), .RSTB(I93615_rst), .Q(I93598) );
nand I_5195 (I93607,I93991,I93943);
DFFARX1 I_5196  ( .D(I93991), .CLK(I5694_clk), .RSTB(I93615_rst), .Q(I93577) );
DFFARX1 I_5197  ( .D(I17284), .CLK(I5694_clk), .RSTB(I93615_rst), .Q(I94067) );
nand I_5198 (I93601,I94067,I93762);
DFFARX1 I_5199  ( .D(I94067), .CLK(I5694_clk), .RSTB(I93615_rst), .Q(I93589) );
nand I_5200 (I94112,I94067,I93728);
and I_5201 (I94129,I93779,I94112);
DFFARX1 I_5202  ( .D(I94129), .CLK(I5694_clk), .RSTB(I93615_rst), .Q(I93583) );
not I_5203 (I94193_rst,I5701);
nand I_5204 (I94210,I78366,I78345);
and I_5205 (I94227,I94210,I78363);
DFFARX1 I_5206  ( .D(I94227), .CLK(I5694_clk), .RSTB(I94193_rst), .Q(I94244) );
not I_5207 (I94182,I94244);
DFFARX1 I_5208  ( .D(I94244), .CLK(I5694_clk), .RSTB(I94193_rst), .Q(I94275) );
not I_5209 (I94170,I94275);
nor I_5210 (I94306,I78375,I78345);
not I_5211 (I94323,I94306);
nor I_5212 (I94340,I94244,I94323);
DFFARX1 I_5213  ( .D(I78351), .CLK(I5694_clk), .RSTB(I94193_rst), .Q(I94357) );
not I_5214 (I94374,I94357);
nand I_5215 (I94173,I94357,I94323);
DFFARX1 I_5216  ( .D(I94357), .CLK(I5694_clk), .RSTB(I94193_rst), .Q(I94405) );
and I_5217 (I94158,I94244,I94405);
nand I_5218 (I94436,I78360,I78348);
and I_5219 (I94453,I94436,I78372);
DFFARX1 I_5220  ( .D(I94453), .CLK(I5694_clk), .RSTB(I94193_rst), .Q(I94470) );
nor I_5221 (I94487,I94470,I94374);
and I_5222 (I94504,I94306,I94487);
nor I_5223 (I94521,I94470,I94244);
DFFARX1 I_5224  ( .D(I94470), .CLK(I5694_clk), .RSTB(I94193_rst), .Q(I94164) );
DFFARX1 I_5225  ( .D(I78357), .CLK(I5694_clk), .RSTB(I94193_rst), .Q(I94552) );
and I_5226 (I94569,I94552,I78369);
or I_5227 (I94586,I94569,I94504);
DFFARX1 I_5228  ( .D(I94586), .CLK(I5694_clk), .RSTB(I94193_rst), .Q(I94176) );
nand I_5229 (I94185,I94569,I94521);
DFFARX1 I_5230  ( .D(I94569), .CLK(I5694_clk), .RSTB(I94193_rst), .Q(I94155) );
DFFARX1 I_5231  ( .D(I78354), .CLK(I5694_clk), .RSTB(I94193_rst), .Q(I94645) );
nand I_5232 (I94179,I94645,I94340);
DFFARX1 I_5233  ( .D(I94645), .CLK(I5694_clk), .RSTB(I94193_rst), .Q(I94167) );
nand I_5234 (I94690,I94645,I94306);
and I_5235 (I94707,I94357,I94690);
DFFARX1 I_5236  ( .D(I94707), .CLK(I5694_clk), .RSTB(I94193_rst), .Q(I94161) );
not I_5237 (I94771_rst,I5701);
nand I_5238 (I94788,I90058,I90061);
and I_5239 (I94805,I94788,I90067);
DFFARX1 I_5240  ( .D(I94805), .CLK(I5694_clk), .RSTB(I94771_rst), .Q(I94822) );
not I_5241 (I94839,I94822);
nor I_5242 (I94856,I90079,I90061);
or I_5243 (I94754,I94856,I94822);
not I_5244 (I94742,I94856);
DFFARX1 I_5245  ( .D(I90088), .CLK(I5694_clk), .RSTB(I94771_rst), .Q(I94901) );
nor I_5246 (I94918,I94901,I94856);
nand I_5247 (I94935,I90076,I90073);
and I_5248 (I94952,I94935,I90085);
DFFARX1 I_5249  ( .D(I94952), .CLK(I5694_clk), .RSTB(I94771_rst), .Q(I94969) );
nor I_5250 (I94751,I94969,I94822);
not I_5251 (I95000,I94969);
nor I_5252 (I95017,I94901,I95000);
DFFARX1 I_5253  ( .D(I90082), .CLK(I5694_clk), .RSTB(I94771_rst), .Q(I95034) );
and I_5254 (I95051,I95034,I90070);
or I_5255 (I94760,I95051,I94856);
nand I_5256 (I94739,I95051,I95017);
DFFARX1 I_5257  ( .D(I90064), .CLK(I5694_clk), .RSTB(I94771_rst), .Q(I95096) );
and I_5258 (I95113,I95096,I94839);
nor I_5259 (I94757,I95051,I95113);
nor I_5260 (I95144,I95096,I94901);
DFFARX1 I_5261  ( .D(I95144), .CLK(I5694_clk), .RSTB(I94771_rst), .Q(I94748) );
nor I_5262 (I94763,I95096,I94822);
not I_5263 (I95189,I95096);
nor I_5264 (I95206,I94969,I95189);
and I_5265 (I95223,I94856,I95206);
or I_5266 (I95240,I95051,I95223);
DFFARX1 I_5267  ( .D(I95240), .CLK(I5694_clk), .RSTB(I94771_rst), .Q(I94736) );
nand I_5268 (I94745,I95096,I94918);
nand I_5269 (I94733,I95096,I95000);
not I_5270 (I95332_rst,I5701);
nand I_5271 (I95349,I56989,I56980);
and I_5272 (I95366,I95349,I56983);
DFFARX1 I_5273  ( .D(I95366), .CLK(I5694_clk), .RSTB(I95332_rst), .Q(I95383) );
not I_5274 (I95400,I95383);
nor I_5275 (I95417,I56959,I56980);
or I_5276 (I95315,I95417,I95383);
not I_5277 (I95303,I95417);
DFFARX1 I_5278  ( .D(I56974), .CLK(I5694_clk), .RSTB(I95332_rst), .Q(I95462) );
nor I_5279 (I95479,I95462,I95417);
nand I_5280 (I95496,I56962,I56977);
and I_5281 (I95513,I95496,I56971);
DFFARX1 I_5282  ( .D(I95513), .CLK(I5694_clk), .RSTB(I95332_rst), .Q(I95530) );
nor I_5283 (I95312,I95530,I95383);
not I_5284 (I95561,I95530);
nor I_5285 (I95578,I95462,I95561);
DFFARX1 I_5286  ( .D(I56986), .CLK(I5694_clk), .RSTB(I95332_rst), .Q(I95595) );
and I_5287 (I95612,I95595,I56965);
or I_5288 (I95321,I95612,I95417);
nand I_5289 (I95300,I95612,I95578);
DFFARX1 I_5290  ( .D(I56968), .CLK(I5694_clk), .RSTB(I95332_rst), .Q(I95657) );
and I_5291 (I95674,I95657,I95400);
nor I_5292 (I95318,I95612,I95674);
nor I_5293 (I95705,I95657,I95462);
DFFARX1 I_5294  ( .D(I95705), .CLK(I5694_clk), .RSTB(I95332_rst), .Q(I95309) );
nor I_5295 (I95324,I95657,I95383);
not I_5296 (I95750,I95657);
nor I_5297 (I95767,I95530,I95750);
and I_5298 (I95784,I95417,I95767);
or I_5299 (I95801,I95612,I95784);
DFFARX1 I_5300  ( .D(I95801), .CLK(I5694_clk), .RSTB(I95332_rst), .Q(I95297) );
nand I_5301 (I95306,I95657,I95479);
nand I_5302 (I95294,I95657,I95561);
not I_5303 (I95893_rst,I5701);
nand I_5304 (I95910,I64095,I64086);
and I_5305 (I95927,I95910,I64089);
DFFARX1 I_5306  ( .D(I95927), .CLK(I5694_clk), .RSTB(I95893_rst), .Q(I95944) );
not I_5307 (I95961,I95944);
nor I_5308 (I95978,I64065,I64086);
or I_5309 (I95876,I95978,I95944);
not I_5310 (I95864,I95978);
DFFARX1 I_5311  ( .D(I64080), .CLK(I5694_clk), .RSTB(I95893_rst), .Q(I96023) );
nor I_5312 (I96040,I96023,I95978);
nand I_5313 (I96057,I64068,I64083);
and I_5314 (I96074,I96057,I64077);
DFFARX1 I_5315  ( .D(I96074), .CLK(I5694_clk), .RSTB(I95893_rst), .Q(I96091) );
nor I_5316 (I95873,I96091,I95944);
not I_5317 (I96122,I96091);
nor I_5318 (I96139,I96023,I96122);
DFFARX1 I_5319  ( .D(I64092), .CLK(I5694_clk), .RSTB(I95893_rst), .Q(I96156) );
and I_5320 (I96173,I96156,I64071);
or I_5321 (I95882,I96173,I95978);
nand I_5322 (I95861,I96173,I96139);
DFFARX1 I_5323  ( .D(I64074), .CLK(I5694_clk), .RSTB(I95893_rst), .Q(I96218) );
and I_5324 (I96235,I96218,I95961);
nor I_5325 (I95879,I96173,I96235);
nor I_5326 (I96266,I96218,I96023);
DFFARX1 I_5327  ( .D(I96266), .CLK(I5694_clk), .RSTB(I95893_rst), .Q(I95870) );
nor I_5328 (I95885,I96218,I95944);
not I_5329 (I96311,I96218);
nor I_5330 (I96328,I96091,I96311);
and I_5331 (I96345,I95978,I96328);
or I_5332 (I96362,I96173,I96345);
DFFARX1 I_5333  ( .D(I96362), .CLK(I5694_clk), .RSTB(I95893_rst), .Q(I95858) );
nand I_5334 (I95867,I96218,I96040);
nand I_5335 (I95855,I96218,I96122);
not I_5336 (I96454_rst,I5701);
nand I_5337 (I96471,I47327,I47330);
and I_5338 (I96488,I96471,I47324);
DFFARX1 I_5339  ( .D(I96488), .CLK(I5694_clk), .RSTB(I96454_rst), .Q(I96505) );
not I_5340 (I96522,I96505);
nor I_5341 (I96539,I47315,I47330);
or I_5342 (I96437,I96539,I96505);
not I_5343 (I96425,I96539);
DFFARX1 I_5344  ( .D(I47303), .CLK(I5694_clk), .RSTB(I96454_rst), .Q(I96584) );
nor I_5345 (I96601,I96584,I96539);
nand I_5346 (I96618,I47312,I47306);
and I_5347 (I96635,I96618,I47318);
DFFARX1 I_5348  ( .D(I96635), .CLK(I5694_clk), .RSTB(I96454_rst), .Q(I96652) );
nor I_5349 (I96434,I96652,I96505);
not I_5350 (I96683,I96652);
nor I_5351 (I96700,I96584,I96683);
DFFARX1 I_5352  ( .D(I47333), .CLK(I5694_clk), .RSTB(I96454_rst), .Q(I96717) );
and I_5353 (I96734,I96717,I47321);
or I_5354 (I96443,I96734,I96539);
nand I_5355 (I96422,I96734,I96700);
DFFARX1 I_5356  ( .D(I47309), .CLK(I5694_clk), .RSTB(I96454_rst), .Q(I96779) );
and I_5357 (I96796,I96779,I96522);
nor I_5358 (I96440,I96734,I96796);
nor I_5359 (I96827,I96779,I96584);
DFFARX1 I_5360  ( .D(I96827), .CLK(I5694_clk), .RSTB(I96454_rst), .Q(I96431) );
nor I_5361 (I96446,I96779,I96505);
not I_5362 (I96872,I96779);
nor I_5363 (I96889,I96652,I96872);
and I_5364 (I96906,I96539,I96889);
or I_5365 (I96923,I96734,I96906);
DFFARX1 I_5366  ( .D(I96923), .CLK(I5694_clk), .RSTB(I96454_rst), .Q(I96419) );
nand I_5367 (I96428,I96779,I96601);
nand I_5368 (I96416,I96779,I96683);
not I_5369 (I97015_rst,I5701);
nand I_5370 (I97032,I81341,I81329);
and I_5371 (I97049,I97032,I81326);
DFFARX1 I_5372  ( .D(I97049), .CLK(I5694_clk), .RSTB(I97015_rst), .Q(I97066) );
not I_5373 (I97083,I97066);
nor I_5374 (I97100,I81347,I81329);
or I_5375 (I96998,I97100,I97066);
not I_5376 (I96986,I97100);
DFFARX1 I_5377  ( .D(I81350), .CLK(I5694_clk), .RSTB(I97015_rst), .Q(I97145) );
nor I_5378 (I97162,I97145,I97100);
nand I_5379 (I97179,I81320,I81338);
and I_5380 (I97196,I97179,I81335);
DFFARX1 I_5381  ( .D(I97196), .CLK(I5694_clk), .RSTB(I97015_rst), .Q(I97213) );
nor I_5382 (I96995,I97213,I97066);
not I_5383 (I97244,I97213);
nor I_5384 (I97261,I97145,I97244);
DFFARX1 I_5385  ( .D(I81344), .CLK(I5694_clk), .RSTB(I97015_rst), .Q(I97278) );
and I_5386 (I97295,I97278,I81332);
or I_5387 (I97004,I97295,I97100);
nand I_5388 (I96983,I97295,I97261);
DFFARX1 I_5389  ( .D(I81323), .CLK(I5694_clk), .RSTB(I97015_rst), .Q(I97340) );
and I_5390 (I97357,I97340,I97083);
nor I_5391 (I97001,I97295,I97357);
nor I_5392 (I97388,I97340,I97145);
DFFARX1 I_5393  ( .D(I97388), .CLK(I5694_clk), .RSTB(I97015_rst), .Q(I96992) );
nor I_5394 (I97007,I97340,I97066);
not I_5395 (I97433,I97340);
nor I_5396 (I97450,I97213,I97433);
and I_5397 (I97467,I97100,I97450);
or I_5398 (I97484,I97295,I97467);
DFFARX1 I_5399  ( .D(I97484), .CLK(I5694_clk), .RSTB(I97015_rst), .Q(I96980) );
nand I_5400 (I96989,I97340,I97162);
nand I_5401 (I96977,I97340,I97244);
not I_5402 (I97576_rst,I5701);
nand I_5403 (I97593,I67171,I67168);
and I_5404 (I97610,I97593,I67162);
DFFARX1 I_5405  ( .D(I97610), .CLK(I5694_clk), .RSTB(I97576_rst), .Q(I97627) );
not I_5406 (I97644,I97627);
nor I_5407 (I97661,I67174,I67168);
or I_5408 (I97559,I97661,I97627);
not I_5409 (I97547,I97661);
DFFARX1 I_5410  ( .D(I67186), .CLK(I5694_clk), .RSTB(I97576_rst), .Q(I97706) );
nor I_5411 (I97723,I97706,I97661);
nand I_5412 (I97740,I67177,I67159);
and I_5413 (I97757,I97740,I67189);
DFFARX1 I_5414  ( .D(I97757), .CLK(I5694_clk), .RSTB(I97576_rst), .Q(I97774) );
nor I_5415 (I97556,I97774,I97627);
not I_5416 (I97805,I97774);
nor I_5417 (I97822,I97706,I97805);
DFFARX1 I_5418  ( .D(I67165), .CLK(I5694_clk), .RSTB(I97576_rst), .Q(I97839) );
and I_5419 (I97856,I97839,I67183);
or I_5420 (I97565,I97856,I97661);
nand I_5421 (I97544,I97856,I97822);
DFFARX1 I_5422  ( .D(I67180), .CLK(I5694_clk), .RSTB(I97576_rst), .Q(I97901) );
and I_5423 (I97918,I97901,I97644);
nor I_5424 (I97562,I97856,I97918);
nor I_5425 (I97949,I97901,I97706);
DFFARX1 I_5426  ( .D(I97949), .CLK(I5694_clk), .RSTB(I97576_rst), .Q(I97553) );
nor I_5427 (I97568,I97901,I97627);
not I_5428 (I97994,I97901);
nor I_5429 (I98011,I97774,I97994);
and I_5430 (I98028,I97661,I98011);
or I_5431 (I98045,I97856,I98028);
DFFARX1 I_5432  ( .D(I98045), .CLK(I5694_clk), .RSTB(I97576_rst), .Q(I97541) );
nand I_5433 (I97550,I97901,I97723);
nand I_5434 (I97538,I97901,I97805);
not I_5435 (I98137_rst,I5701);
nand I_5436 (I98154,I84397,I84400);
and I_5437 (I98171,I98154,I84406);
DFFARX1 I_5438  ( .D(I98171), .CLK(I5694_clk), .RSTB(I98137_rst), .Q(I98188) );
not I_5439 (I98205,I98188);
nor I_5440 (I98222,I84418,I84400);
or I_5441 (I98120,I98222,I98188);
not I_5442 (I98108,I98222);
DFFARX1 I_5443  ( .D(I84427), .CLK(I5694_clk), .RSTB(I98137_rst), .Q(I98267) );
nor I_5444 (I98284,I98267,I98222);
nand I_5445 (I98301,I84415,I84412);
and I_5446 (I98318,I98301,I84424);
DFFARX1 I_5447  ( .D(I98318), .CLK(I5694_clk), .RSTB(I98137_rst), .Q(I98335) );
nor I_5448 (I98117,I98335,I98188);
not I_5449 (I98366,I98335);
nor I_5450 (I98383,I98267,I98366);
DFFARX1 I_5451  ( .D(I84421), .CLK(I5694_clk), .RSTB(I98137_rst), .Q(I98400) );
and I_5452 (I98417,I98400,I84409);
or I_5453 (I98126,I98417,I98222);
nand I_5454 (I98105,I98417,I98383);
DFFARX1 I_5455  ( .D(I84403), .CLK(I5694_clk), .RSTB(I98137_rst), .Q(I98462) );
and I_5456 (I98479,I98462,I98205);
nor I_5457 (I98123,I98417,I98479);
nor I_5458 (I98510,I98462,I98267);
DFFARX1 I_5459  ( .D(I98510), .CLK(I5694_clk), .RSTB(I98137_rst), .Q(I98114) );
nor I_5460 (I98129,I98462,I98188);
not I_5461 (I98555,I98462);
nor I_5462 (I98572,I98335,I98555);
and I_5463 (I98589,I98222,I98572);
or I_5464 (I98606,I98417,I98589);
DFFARX1 I_5465  ( .D(I98606), .CLK(I5694_clk), .RSTB(I98137_rst), .Q(I98102) );
nand I_5466 (I98111,I98462,I98284);
nand I_5467 (I98099,I98462,I98366);
not I_5468 (I98698_rst,I5701);
not I_5469 (I98715,I85026);
nor I_5470 (I98732,I85041,I85056);
nand I_5471 (I98749,I98732,I85044);
DFFARX1 I_5472  ( .D(I98749), .CLK(I5694_clk), .RSTB(I98698_rst), .Q(I98672) );
nor I_5473 (I98780,I98715,I85041);
nand I_5474 (I98797,I98780,I85047);
not I_5475 (I98687,I98797);
DFFARX1 I_5476  ( .D(I98797), .CLK(I5694_clk), .RSTB(I98698_rst), .Q(I98669) );
not I_5477 (I98842,I85041);
not I_5478 (I98859,I98842);
not I_5479 (I98876,I85053);
nor I_5480 (I98893,I98876,I85050);
and I_5481 (I98910,I98893,I85029);
or I_5482 (I98927,I98910,I85038);
DFFARX1 I_5483  ( .D(I98927), .CLK(I5694_clk), .RSTB(I98698_rst), .Q(I98944) );
nor I_5484 (I98961,I98944,I98797);
nor I_5485 (I98978,I98944,I98859);
nand I_5486 (I98684,I98749,I98978);
nand I_5487 (I99009,I98715,I85053);
nand I_5488 (I99026,I99009,I98944);
and I_5489 (I99043,I99009,I99026);
DFFARX1 I_5490  ( .D(I99043), .CLK(I5694_clk), .RSTB(I98698_rst), .Q(I98666) );
DFFARX1 I_5491  ( .D(I99009), .CLK(I5694_clk), .RSTB(I98698_rst), .Q(I99074) );
and I_5492 (I98663,I98842,I99074);
DFFARX1 I_5493  ( .D(I85035), .CLK(I5694_clk), .RSTB(I98698_rst), .Q(I99105) );
not I_5494 (I99122,I99105);
nor I_5495 (I99139,I98797,I99122);
and I_5496 (I99156,I99105,I99139);
nand I_5497 (I98678,I99105,I98859);
DFFARX1 I_5498  ( .D(I99105), .CLK(I5694_clk), .RSTB(I98698_rst), .Q(I99187) );
not I_5499 (I98675,I99187);
DFFARX1 I_5500  ( .D(I85032), .CLK(I5694_clk), .RSTB(I98698_rst), .Q(I99218) );
not I_5501 (I99235,I99218);
or I_5502 (I99252,I99235,I99156);
DFFARX1 I_5503  ( .D(I99252), .CLK(I5694_clk), .RSTB(I98698_rst), .Q(I98681) );
nand I_5504 (I98690,I99235,I98961);
DFFARX1 I_5505  ( .D(I99235), .CLK(I5694_clk), .RSTB(I98698_rst), .Q(I98660) );
not I_5506 (I99344_rst,I5701);
not I_5507 (I99361,I71807);
nor I_5508 (I99378,I71789,I71798);
nand I_5509 (I99395,I99378,I71810);
DFFARX1 I_5510  ( .D(I99395), .CLK(I5694_clk), .RSTB(I99344_rst), .Q(I99318) );
nor I_5511 (I99426,I99361,I71789);
nand I_5512 (I99443,I99426,I71795);
not I_5513 (I99333,I99443);
DFFARX1 I_5514  ( .D(I99443), .CLK(I5694_clk), .RSTB(I99344_rst), .Q(I99315) );
not I_5515 (I99488,I71789);
not I_5516 (I99505,I99488);
not I_5517 (I99522,I71786);
nor I_5518 (I99539,I99522,I71804);
and I_5519 (I99556,I99539,I71792);
or I_5520 (I99573,I99556,I71813);
DFFARX1 I_5521  ( .D(I99573), .CLK(I5694_clk), .RSTB(I99344_rst), .Q(I99590) );
nor I_5522 (I99607,I99590,I99443);
nor I_5523 (I99624,I99590,I99505);
nand I_5524 (I99330,I99395,I99624);
nand I_5525 (I99655,I99361,I71786);
nand I_5526 (I99672,I99655,I99590);
and I_5527 (I99689,I99655,I99672);
DFFARX1 I_5528  ( .D(I99689), .CLK(I5694_clk), .RSTB(I99344_rst), .Q(I99312) );
DFFARX1 I_5529  ( .D(I99655), .CLK(I5694_clk), .RSTB(I99344_rst), .Q(I99720) );
and I_5530 (I99309,I99488,I99720);
DFFARX1 I_5531  ( .D(I71801), .CLK(I5694_clk), .RSTB(I99344_rst), .Q(I99751) );
not I_5532 (I99768,I99751);
nor I_5533 (I99785,I99443,I99768);
and I_5534 (I99802,I99751,I99785);
nand I_5535 (I99324,I99751,I99505);
DFFARX1 I_5536  ( .D(I99751), .CLK(I5694_clk), .RSTB(I99344_rst), .Q(I99833) );
not I_5537 (I99321,I99833);
DFFARX1 I_5538  ( .D(I71783), .CLK(I5694_clk), .RSTB(I99344_rst), .Q(I99864) );
not I_5539 (I99881,I99864);
or I_5540 (I99898,I99881,I99802);
DFFARX1 I_5541  ( .D(I99898), .CLK(I5694_clk), .RSTB(I99344_rst), .Q(I99327) );
nand I_5542 (I99336,I99881,I99607);
DFFARX1 I_5543  ( .D(I99881), .CLK(I5694_clk), .RSTB(I99344_rst), .Q(I99306) );
not I_5544 (I99990_rst,I5701);
not I_5545 (I100007,I66596);
nor I_5546 (I100024,I66584,I66590);
nand I_5547 (I100041,I100024,I66581);
DFFARX1 I_5548  ( .D(I100041), .CLK(I5694_clk), .RSTB(I99990_rst), .Q(I99964) );
nor I_5549 (I100072,I100007,I66584);
nand I_5550 (I100089,I100072,I66587);
not I_5551 (I99979,I100089);
DFFARX1 I_5552  ( .D(I100089), .CLK(I5694_clk), .RSTB(I99990_rst), .Q(I99961) );
not I_5553 (I100134,I66584);
not I_5554 (I100151,I100134);
not I_5555 (I100168,I66599);
nor I_5556 (I100185,I100168,I66611);
and I_5557 (I100202,I100185,I66593);
or I_5558 (I100219,I100202,I66608);
DFFARX1 I_5559  ( .D(I100219), .CLK(I5694_clk), .RSTB(I99990_rst), .Q(I100236) );
nor I_5560 (I100253,I100236,I100089);
nor I_5561 (I100270,I100236,I100151);
nand I_5562 (I99976,I100041,I100270);
nand I_5563 (I100301,I100007,I66599);
nand I_5564 (I100318,I100301,I100236);
and I_5565 (I100335,I100301,I100318);
DFFARX1 I_5566  ( .D(I100335), .CLK(I5694_clk), .RSTB(I99990_rst), .Q(I99958) );
DFFARX1 I_5567  ( .D(I100301), .CLK(I5694_clk), .RSTB(I99990_rst), .Q(I100366) );
and I_5568 (I99955,I100134,I100366);
DFFARX1 I_5569  ( .D(I66602), .CLK(I5694_clk), .RSTB(I99990_rst), .Q(I100397) );
not I_5570 (I100414,I100397);
nor I_5571 (I100431,I100089,I100414);
and I_5572 (I100448,I100397,I100431);
nand I_5573 (I99970,I100397,I100151);
DFFARX1 I_5574  ( .D(I100397), .CLK(I5694_clk), .RSTB(I99990_rst), .Q(I100479) );
not I_5575 (I99967,I100479);
DFFARX1 I_5576  ( .D(I66605), .CLK(I5694_clk), .RSTB(I99990_rst), .Q(I100510) );
not I_5577 (I100527,I100510);
or I_5578 (I100544,I100527,I100448);
DFFARX1 I_5579  ( .D(I100544), .CLK(I5694_clk), .RSTB(I99990_rst), .Q(I99973) );
nand I_5580 (I99982,I100527,I100253);
DFFARX1 I_5581  ( .D(I100527), .CLK(I5694_clk), .RSTB(I99990_rst), .Q(I99952) );
not I_5582 (I100636_rst,I5701);
not I_5583 (I100653,I46708);
nor I_5584 (I100670,I46738,I46717);
nand I_5585 (I100687,I100670,I46729);
DFFARX1 I_5586  ( .D(I100687), .CLK(I5694_clk), .RSTB(I100636_rst), .Q(I100610) );
nor I_5587 (I100718,I100653,I46738);
nand I_5588 (I100735,I100718,I46711);
not I_5589 (I100625,I100735);
DFFARX1 I_5590  ( .D(I100735), .CLK(I5694_clk), .RSTB(I100636_rst), .Q(I100607) );
not I_5591 (I100780,I46738);
not I_5592 (I100797,I100780);
not I_5593 (I100814,I46714);
nor I_5594 (I100831,I100814,I46732);
and I_5595 (I100848,I100831,I46723);
or I_5596 (I100865,I100848,I46720);
DFFARX1 I_5597  ( .D(I100865), .CLK(I5694_clk), .RSTB(I100636_rst), .Q(I100882) );
nor I_5598 (I100899,I100882,I100735);
nor I_5599 (I100916,I100882,I100797);
nand I_5600 (I100622,I100687,I100916);
nand I_5601 (I100947,I100653,I46714);
nand I_5602 (I100964,I100947,I100882);
and I_5603 (I100981,I100947,I100964);
DFFARX1 I_5604  ( .D(I100981), .CLK(I5694_clk), .RSTB(I100636_rst), .Q(I100604) );
DFFARX1 I_5605  ( .D(I100947), .CLK(I5694_clk), .RSTB(I100636_rst), .Q(I101012) );
and I_5606 (I100601,I100780,I101012);
DFFARX1 I_5607  ( .D(I46726), .CLK(I5694_clk), .RSTB(I100636_rst), .Q(I101043) );
not I_5608 (I101060,I101043);
nor I_5609 (I101077,I100735,I101060);
and I_5610 (I101094,I101043,I101077);
nand I_5611 (I100616,I101043,I100797);
DFFARX1 I_5612  ( .D(I101043), .CLK(I5694_clk), .RSTB(I100636_rst), .Q(I101125) );
not I_5613 (I100613,I101125);
DFFARX1 I_5614  ( .D(I46735), .CLK(I5694_clk), .RSTB(I100636_rst), .Q(I101156) );
not I_5615 (I101173,I101156);
or I_5616 (I101190,I101173,I101094);
DFFARX1 I_5617  ( .D(I101190), .CLK(I5694_clk), .RSTB(I100636_rst), .Q(I100619) );
nand I_5618 (I100628,I101173,I100899);
DFFARX1 I_5619  ( .D(I101173), .CLK(I5694_clk), .RSTB(I100636_rst), .Q(I100598) );
not I_5620 (I101282_rst,I5701);
not I_5621 (I101299,I74802);
nor I_5622 (I101316,I74778,I74784);
nand I_5623 (I101333,I101316,I74787);
DFFARX1 I_5624  ( .D(I101333), .CLK(I5694_clk), .RSTB(I101282_rst), .Q(I101256) );
nor I_5625 (I101364,I101299,I74778);
nand I_5626 (I101381,I101364,I74796);
not I_5627 (I101271,I101381);
DFFARX1 I_5628  ( .D(I101381), .CLK(I5694_clk), .RSTB(I101282_rst), .Q(I101253) );
not I_5629 (I101426,I74778);
not I_5630 (I101443,I101426);
not I_5631 (I101460,I74775);
nor I_5632 (I101477,I101460,I74790);
and I_5633 (I101494,I101477,I74781);
or I_5634 (I101511,I101494,I74793);
DFFARX1 I_5635  ( .D(I101511), .CLK(I5694_clk), .RSTB(I101282_rst), .Q(I101528) );
nor I_5636 (I101545,I101528,I101381);
nor I_5637 (I101562,I101528,I101443);
nand I_5638 (I101268,I101333,I101562);
nand I_5639 (I101593,I101299,I74775);
nand I_5640 (I101610,I101593,I101528);
and I_5641 (I10162_rst7,I101593,I101610);
DFFARX1 I_5642  ( .D(I10162_rst7), .CLK(I5694_clk), .RSTB(I101282_rst), .Q(I101250) );
DFFARX1 I_5643  ( .D(I101593), .CLK(I5694_clk), .RSTB(I101282_rst), .Q(I101658) );
and I_5644 (I101247,I101426,I101658);
DFFARX1 I_5645  ( .D(I74805), .CLK(I5694_clk), .RSTB(I101282_rst), .Q(I101689) );
not I_5646 (I101706,I101689);
nor I_5647 (I101723,I101381,I101706);
and I_5648 (I101740,I101689,I101723);
nand I_5649 (I101262,I101689,I101443);
DFFARX1 I_5650  ( .D(I101689), .CLK(I5694_clk), .RSTB(I101282_rst), .Q(I101771) );
not I_5651 (I101259,I101771);
DFFARX1 I_5652  ( .D(I74799), .CLK(I5694_clk), .RSTB(I101282_rst), .Q(I101802) );
not I_5653 (I101819,I101802);
or I_5654 (I101836,I101819,I101740);
DFFARX1 I_5655  ( .D(I101836), .CLK(I5694_clk), .RSTB(I101282_rst), .Q(I101265) );
nand I_5656 (I101274,I101819,I101545);
DFFARX1 I_5657  ( .D(I101819), .CLK(I5694_clk), .RSTB(I101282_rst), .Q(I101244) );
not I_5658 (I101928_rst,I5701);
not I_5659 (I101945,I80145);
nor I_5660 (I101962,I80130,I80157);
nand I_5661 (I101979,I101962,I80133);
DFFARX1 I_5662  ( .D(I101979), .CLK(I5694_clk), .RSTB(I101928_rst), .Q(I101902) );
nor I_5663 (I102010,I101945,I80130);
nand I_5664 (I102027,I102010,I80148);
not I_5665 (I101917,I102027);
DFFARX1 I_5666  ( .D(I102027), .CLK(I5694_clk), .RSTB(I101928_rst), .Q(I101899) );
not I_5667 (I102072,I80130);
not I_5668 (I102089,I102072);
not I_5669 (I102106,I80160);
nor I_5670 (I102123,I102106,I80142);
and I_5671 (I102140,I102123,I80151);
or I_5672 (I102157,I102140,I80136);
DFFARX1 I_5673  ( .D(I102157), .CLK(I5694_clk), .RSTB(I101928_rst), .Q(I102174) );
nor I_5674 (I102191,I102174,I102027);
nor I_5675 (I102208,I102174,I102089);
nand I_5676 (I101914,I101979,I102208);
nand I_5677 (I102239,I101945,I80160);
nand I_5678 (I102256,I102239,I102174);
and I_5679 (I102273,I102239,I102256);
DFFARX1 I_5680  ( .D(I102273), .CLK(I5694_clk), .RSTB(I101928_rst), .Q(I101896) );
DFFARX1 I_5681  ( .D(I102239), .CLK(I5694_clk), .RSTB(I101928_rst), .Q(I102304) );
and I_5682 (I101893,I102072,I102304);
DFFARX1 I_5683  ( .D(I80139), .CLK(I5694_clk), .RSTB(I101928_rst), .Q(I102335) );
not I_5684 (I102352,I102335);
nor I_5685 (I102369,I102027,I102352);
and I_5686 (I102386,I102335,I102369);
nand I_5687 (I101908,I102335,I102089);
DFFARX1 I_5688  ( .D(I102335), .CLK(I5694_clk), .RSTB(I101928_rst), .Q(I102417) );
not I_5689 (I101905,I102417);
DFFARX1 I_5690  ( .D(I80154), .CLK(I5694_clk), .RSTB(I101928_rst), .Q(I102448) );
not I_5691 (I102465,I102448);
or I_5692 (I102482,I102465,I102386);
DFFARX1 I_5693  ( .D(I102482), .CLK(I5694_clk), .RSTB(I101928_rst), .Q(I101911) );
nand I_5694 (I101920,I102465,I102191);
DFFARX1 I_5695  ( .D(I102465), .CLK(I5694_clk), .RSTB(I101928_rst), .Q(I101890) );
not I_5696 (I102574_rst,I5701);
not I_5697 (I102591,I94164);
nor I_5698 (I102608,I94161,I94158);
nand I_5699 (I102625,I102608,I94179);
DFFARX1 I_5700  ( .D(I102625), .CLK(I5694_clk), .RSTB(I102574_rst), .Q(I102548) );
nor I_5701 (I102656,I102591,I94161);
nand I_5702 (I102673,I102656,I94182);
not I_5703 (I102563,I102673);
DFFARX1 I_5704  ( .D(I102673), .CLK(I5694_clk), .RSTB(I102574_rst), .Q(I102545) );
not I_5705 (I102718,I94161);
not I_5706 (I102735,I102718);
not I_5707 (I102752,I94155);
nor I_5708 (I102769,I102752,I94167);
and I_5709 (I102786,I102769,I94176);
or I_5710 (I102803,I102786,I94170);
DFFARX1 I_5711  ( .D(I102803), .CLK(I5694_clk), .RSTB(I102574_rst), .Q(I102820) );
nor I_5712 (I102837,I102820,I102673);
nor I_5713 (I102854,I102820,I102735);
nand I_5714 (I102560,I102625,I102854);
nand I_5715 (I102885,I102591,I94155);
nand I_5716 (I102902,I102885,I102820);
and I_5717 (I102919,I102885,I102902);
DFFARX1 I_5718  ( .D(I102919), .CLK(I5694_clk), .RSTB(I102574_rst), .Q(I102542) );
DFFARX1 I_5719  ( .D(I102885), .CLK(I5694_clk), .RSTB(I102574_rst), .Q(I102950) );
and I_5720 (I102539,I102718,I102950);
DFFARX1 I_5721  ( .D(I94185), .CLK(I5694_clk), .RSTB(I102574_rst), .Q(I102981) );
not I_5722 (I102998,I102981);
nor I_5723 (I103015,I102673,I102998);
and I_5724 (I103032,I102981,I103015);
nand I_5725 (I102554,I102981,I102735);
DFFARX1 I_5726  ( .D(I102981), .CLK(I5694_clk), .RSTB(I102574_rst), .Q(I103063) );
not I_5727 (I102551,I103063);
DFFARX1 I_5728  ( .D(I94173), .CLK(I5694_clk), .RSTB(I102574_rst), .Q(I103094) );
not I_5729 (I103111,I103094);
or I_5730 (I103128,I103111,I103032);
DFFARX1 I_5731  ( .D(I103128), .CLK(I5694_clk), .RSTB(I102574_rst), .Q(I102557) );
nand I_5732 (I102566,I103111,I102837);
DFFARX1 I_5733  ( .D(I103111), .CLK(I5694_clk), .RSTB(I102574_rst), .Q(I102536) );
not I_5734 (I103220_rst,I5701);
not I_5735 (I103237,I96980);
nor I_5736 (I103254,I96992,I96977);
nand I_5737 (I103271,I103254,I96989);
DFFARX1 I_5738  ( .D(I103271), .CLK(I5694_clk), .RSTB(I103220_rst), .Q(I103194) );
nor I_5739 (I103302,I103237,I96992);
nand I_5740 (I103319,I103302,I97007);
not I_5741 (I103209,I103319);
DFFARX1 I_5742  ( .D(I103319), .CLK(I5694_clk), .RSTB(I103220_rst), .Q(I103191) );
not I_5743 (I103364,I96992);
not I_5744 (I103381,I103364);
not I_5745 (I103398,I96983);
nor I_5746 (I103415,I103398,I96995);
and I_5747 (I103432,I103415,I96986);
or I_5748 (I103449,I103432,I97001);
DFFARX1 I_5749  ( .D(I103449), .CLK(I5694_clk), .RSTB(I103220_rst), .Q(I103466) );
nor I_5750 (I103483,I103466,I103319);
nor I_5751 (I103500,I103466,I103381);
nand I_5752 (I103206,I103271,I103500);
nand I_5753 (I103531,I103237,I96983);
nand I_5754 (I103548,I103531,I103466);
and I_5755 (I103565,I103531,I103548);
DFFARX1 I_5756  ( .D(I103565), .CLK(I5694_clk), .RSTB(I103220_rst), .Q(I103188) );
DFFARX1 I_5757  ( .D(I103531), .CLK(I5694_clk), .RSTB(I103220_rst), .Q(I103596) );
and I_5758 (I103185,I103364,I103596);
DFFARX1 I_5759  ( .D(I97004), .CLK(I5694_clk), .RSTB(I103220_rst), .Q(I103627) );
not I_5760 (I103644,I103627);
nor I_5761 (I103661,I103319,I103644);
and I_5762 (I103678,I103627,I103661);
nand I_5763 (I103200,I103627,I103381);
DFFARX1 I_5764  ( .D(I103627), .CLK(I5694_clk), .RSTB(I103220_rst), .Q(I103709) );
not I_5765 (I103197,I103709);
DFFARX1 I_5766  ( .D(I96998), .CLK(I5694_clk), .RSTB(I103220_rst), .Q(I103740) );
not I_5767 (I103757,I103740);
or I_5768 (I103774,I103757,I103678);
DFFARX1 I_5769  ( .D(I103774), .CLK(I5694_clk), .RSTB(I103220_rst), .Q(I103203) );
nand I_5770 (I103212,I103757,I103483);
DFFARX1 I_5771  ( .D(I103757), .CLK(I5694_clk), .RSTB(I103220_rst), .Q(I103182) );
not I_5772 (I103866_rst,I5701);
not I_5773 (I103883,I55005);
nor I_5774 (I103900,I55002,I54990);
nand I_5775 (I103917,I103900,I54993);
DFFARX1 I_5776  ( .D(I103917), .CLK(I5694_clk), .RSTB(I103866_rst), .Q(I103840) );
nor I_5777 (I103948,I103883,I55002);
nand I_5778 (I103965,I103948,I54999);
not I_5779 (I103855,I103965);
DFFARX1 I_5780  ( .D(I103965), .CLK(I5694_clk), .RSTB(I103866_rst), .Q(I103837) );
not I_5781 (I104010,I55002);
not I_5782 (I104027,I104010);
not I_5783 (I104044,I55011);
nor I_5784 (I104061,I104044,I54987);
and I_5785 (I104078,I104061,I55008);
or I_5786 (I104095,I104078,I54996);
DFFARX1 I_5787  ( .D(I104095), .CLK(I5694_clk), .RSTB(I103866_rst), .Q(I104112) );
nor I_5788 (I104129,I104112,I103965);
nor I_5789 (I104146,I104112,I104027);
nand I_5790 (I103852,I103917,I104146);
nand I_5791 (I104177,I103883,I55011);
nand I_5792 (I104194,I104177,I104112);
and I_5793 (I104211,I104177,I104194);
DFFARX1 I_5794  ( .D(I104211), .CLK(I5694_clk), .RSTB(I103866_rst), .Q(I103834) );
DFFARX1 I_5795  ( .D(I104177), .CLK(I5694_clk), .RSTB(I103866_rst), .Q(I104242) );
and I_5796 (I103831,I104010,I104242);
DFFARX1 I_5797  ( .D(I55017), .CLK(I5694_clk), .RSTB(I103866_rst), .Q(I104273) );
not I_5798 (I104290,I104273);
nor I_5799 (I104307,I103965,I104290);
and I_5800 (I104324,I104273,I104307);
nand I_5801 (I103846,I104273,I104027);
DFFARX1 I_5802  ( .D(I104273), .CLK(I5694_clk), .RSTB(I103866_rst), .Q(I104355) );
not I_5803 (I103843,I104355);
DFFARX1 I_5804  ( .D(I55014), .CLK(I5694_clk), .RSTB(I103866_rst), .Q(I104386) );
not I_5805 (I104403,I104386);
or I_5806 (I104420,I104403,I104324);
DFFARX1 I_5807  ( .D(I104420), .CLK(I5694_clk), .RSTB(I103866_rst), .Q(I103849) );
nand I_5808 (I103858,I104403,I104129);
DFFARX1 I_5809  ( .D(I104403), .CLK(I5694_clk), .RSTB(I103866_rst), .Q(I103828) );
not I_5810 (I104512_rst,I5701);
not I_5811 (I104529,I87542);
nor I_5812 (I104546,I87557,I87572);
nand I_5813 (I104563,I104546,I87560);
DFFARX1 I_5814  ( .D(I104563), .CLK(I5694_clk), .RSTB(I104512_rst), .Q(I104486) );
nor I_5815 (I104594,I104529,I87557);
nand I_5816 (I104611,I104594,I87563);
not I_5817 (I104501,I104611);
DFFARX1 I_5818  ( .D(I104611), .CLK(I5694_clk), .RSTB(I104512_rst), .Q(I104483) );
not I_5819 (I104656,I87557);
not I_5820 (I104673,I104656);
not I_5821 (I104690,I87569);
nor I_5822 (I104707,I104690,I87566);
and I_5823 (I104724,I104707,I87545);
or I_5824 (I104741,I104724,I87554);
DFFARX1 I_5825  ( .D(I104741), .CLK(I5694_clk), .RSTB(I104512_rst), .Q(I104758) );
nor I_5826 (I104775,I104758,I104611);
nor I_5827 (I104792,I104758,I104673);
nand I_5828 (I104498,I104563,I104792);
nand I_5829 (I104823,I104529,I87569);
nand I_5830 (I104840,I104823,I104758);
and I_5831 (I104857,I104823,I104840);
DFFARX1 I_5832  ( .D(I104857), .CLK(I5694_clk), .RSTB(I104512_rst), .Q(I104480) );
DFFARX1 I_5833  ( .D(I104823), .CLK(I5694_clk), .RSTB(I104512_rst), .Q(I104888) );
and I_5834 (I104477,I104656,I104888);
DFFARX1 I_5835  ( .D(I87551), .CLK(I5694_clk), .RSTB(I104512_rst), .Q(I104919) );
not I_5836 (I104936,I104919);
nor I_5837 (I104953,I104611,I104936);
and I_5838 (I104970,I104919,I104953);
nand I_5839 (I104492,I104919,I104673);
DFFARX1 I_5840  ( .D(I104919), .CLK(I5694_clk), .RSTB(I104512_rst), .Q(I105001) );
not I_5841 (I104489,I105001);
DFFARX1 I_5842  ( .D(I87548), .CLK(I5694_clk), .RSTB(I104512_rst), .Q(I105032) );
not I_5843 (I105049,I105032);
or I_5844 (I105066,I105049,I104970);
DFFARX1 I_5845  ( .D(I105066), .CLK(I5694_clk), .RSTB(I104512_rst), .Q(I104495) );
nand I_5846 (I104504,I105049,I104775);
DFFARX1 I_5847  ( .D(I105049), .CLK(I5694_clk), .RSTB(I104512_rst), .Q(I104474) );
not I_5848 (I105158_rst,I5701);
not I_5849 (I105175,I71220);
nor I_5850 (I105192,I71208,I71214);
nand I_5851 (I105209,I105192,I71205);
DFFARX1 I_5852  ( .D(I105209), .CLK(I5694_clk), .RSTB(I105158_rst), .Q(I105132) );
nor I_5853 (I105240,I105175,I71208);
nand I_5854 (I105257,I105240,I71211);
not I_5855 (I105147,I105257);
DFFARX1 I_5856  ( .D(I105257), .CLK(I5694_clk), .RSTB(I105158_rst), .Q(I105129) );
not I_5857 (I105302,I71208);
not I_5858 (I105319,I105302);
not I_5859 (I105336,I71223);
nor I_5860 (I105353,I105336,I71235);
and I_5861 (I105370,I105353,I71217);
or I_5862 (I105387,I105370,I71232);
DFFARX1 I_5863  ( .D(I105387), .CLK(I5694_clk), .RSTB(I105158_rst), .Q(I105404) );
nor I_5864 (I105421,I105404,I105257);
nor I_5865 (I105438,I105404,I105319);
nand I_5866 (I105144,I105209,I105438);
nand I_5867 (I105469,I105175,I71223);
nand I_5868 (I105486,I105469,I105404);
and I_5869 (I105503,I105469,I105486);
DFFARX1 I_5870  ( .D(I105503), .CLK(I5694_clk), .RSTB(I105158_rst), .Q(I105126) );
DFFARX1 I_5871  ( .D(I105469), .CLK(I5694_clk), .RSTB(I105158_rst), .Q(I105534) );
and I_5872 (I105123,I105302,I105534);
DFFARX1 I_5873  ( .D(I71226), .CLK(I5694_clk), .RSTB(I105158_rst), .Q(I105565) );
not I_5874 (I105582,I105565);
nor I_5875 (I105599,I105257,I105582);
and I_5876 (I105616,I105565,I105599);
nand I_5877 (I105138,I105565,I105319);
DFFARX1 I_5878  ( .D(I105565), .CLK(I5694_clk), .RSTB(I105158_rst), .Q(I105647) );
not I_5879 (I105135,I105647);
DFFARX1 I_5880  ( .D(I71229), .CLK(I5694_clk), .RSTB(I105158_rst), .Q(I105678) );
not I_5881 (I105695,I105678);
or I_5882 (I105712,I105695,I105616);
DFFARX1 I_5883  ( .D(I105712), .CLK(I5694_clk), .RSTB(I105158_rst), .Q(I105141) );
nand I_5884 (I105150,I105695,I105421);
DFFARX1 I_5885  ( .D(I105695), .CLK(I5694_clk), .RSTB(I105158_rst), .Q(I105120) );
not I_5886 (I105804_rst,I5701);
not I_5887 (I105821,I93008);
nor I_5888 (I105838,I93005,I93002);
nand I_5889 (I105855,I105838,I93023);
DFFARX1 I_5890  ( .D(I105855), .CLK(I5694_clk), .RSTB(I105804_rst), .Q(I105778) );
nor I_5891 (I105886,I105821,I93005);
nand I_5892 (I105903,I105886,I93026);
not I_5893 (I105793,I105903);
DFFARX1 I_5894  ( .D(I105903), .CLK(I5694_clk), .RSTB(I105804_rst), .Q(I105775) );
not I_5895 (I105948,I93005);
not I_5896 (I105965,I105948);
not I_5897 (I105982,I92999);
nor I_5898 (I105999,I105982,I93011);
and I_5899 (I106016,I105999,I93020);
or I_5900 (I106033,I106016,I93014);
DFFARX1 I_5901  ( .D(I106033), .CLK(I5694_clk), .RSTB(I105804_rst), .Q(I106050) );
nor I_5902 (I106067,I106050,I105903);
nor I_5903 (I106084,I106050,I105965);
nand I_5904 (I105790,I105855,I106084);
nand I_5905 (I106115,I105821,I92999);
nand I_5906 (I106132,I106115,I106050);
and I_5907 (I106149,I106115,I106132);
DFFARX1 I_5908  ( .D(I106149), .CLK(I5694_clk), .RSTB(I105804_rst), .Q(I105772) );
DFFARX1 I_5909  ( .D(I106115), .CLK(I5694_clk), .RSTB(I105804_rst), .Q(I106180) );
and I_5910 (I105769,I105948,I106180);
DFFARX1 I_5911  ( .D(I93029), .CLK(I5694_clk), .RSTB(I105804_rst), .Q(I106211) );
not I_5912 (I106228,I106211);
nor I_5913 (I106245,I105903,I106228);
and I_5914 (I106262,I106211,I106245);
nand I_5915 (I105784,I106211,I105965);
DFFARX1 I_5916  ( .D(I106211), .CLK(I5694_clk), .RSTB(I105804_rst), .Q(I106293) );
not I_5917 (I105781,I106293);
DFFARX1 I_5918  ( .D(I93017), .CLK(I5694_clk), .RSTB(I105804_rst), .Q(I106324) );
not I_5919 (I106341,I106324);
or I_5920 (I106358,I106341,I106262);
DFFARX1 I_5921  ( .D(I106358), .CLK(I5694_clk), .RSTB(I105804_rst), .Q(I105787) );
nand I_5922 (I105796,I106341,I106067);
DFFARX1 I_5923  ( .D(I106341), .CLK(I5694_clk), .RSTB(I105804_rst), .Q(I105766) );
not I_5924 (I106450_rst,I5701);
not I_5925 (I106467,I95297);
nor I_5926 (I106484,I95309,I95294);
nand I_5927 (I106501,I106484,I95306);
DFFARX1 I_5928  ( .D(I106501), .CLK(I5694_clk), .RSTB(I106450_rst), .Q(I106424) );
nor I_5929 (I106532,I106467,I95309);
nand I_5930 (I106549,I106532,I95324);
not I_5931 (I106439,I106549);
DFFARX1 I_5932  ( .D(I106549), .CLK(I5694_clk), .RSTB(I106450_rst), .Q(I106421) );
not I_5933 (I106594,I95309);
not I_5934 (I106611,I106594);
not I_5935 (I106628,I95300);
nor I_5936 (I106645,I106628,I95312);
and I_5937 (I106662,I106645,I95303);
or I_5938 (I106679,I106662,I95318);
DFFARX1 I_5939  ( .D(I106679), .CLK(I5694_clk), .RSTB(I106450_rst), .Q(I106696) );
nor I_5940 (I106713,I106696,I106549);
nor I_5941 (I106730,I106696,I106611);
nand I_5942 (I106436,I106501,I106730);
nand I_5943 (I106761,I106467,I95300);
nand I_5944 (I106778,I106761,I106696);
and I_5945 (I106795,I106761,I106778);
DFFARX1 I_5946  ( .D(I106795), .CLK(I5694_clk), .RSTB(I106450_rst), .Q(I106418) );
DFFARX1 I_5947  ( .D(I106761), .CLK(I5694_clk), .RSTB(I106450_rst), .Q(I106826) );
and I_5948 (I106415,I106594,I106826);
DFFARX1 I_5949  ( .D(I95321), .CLK(I5694_clk), .RSTB(I106450_rst), .Q(I106857) );
not I_5950 (I106874,I106857);
nor I_5951 (I106891,I106549,I106874);
and I_5952 (I106908,I106857,I106891);
nand I_5953 (I106430,I106857,I106611);
DFFARX1 I_5954  ( .D(I106857), .CLK(I5694_clk), .RSTB(I106450_rst), .Q(I106939) );
not I_5955 (I106427,I106939);
DFFARX1 I_5956  ( .D(I95315), .CLK(I5694_clk), .RSTB(I106450_rst), .Q(I106970) );
not I_5957 (I106987,I106970);
or I_5958 (I107004,I106987,I106908);
DFFARX1 I_5959  ( .D(I107004), .CLK(I5694_clk), .RSTB(I106450_rst), .Q(I106433) );
nand I_5960 (I106442,I106987,I106713);
DFFARX1 I_5961  ( .D(I106987), .CLK(I5694_clk), .RSTB(I106450_rst), .Q(I106412) );
not I_5962 (I107096_rst,I5701);
not I_5963 (I107113,I86284);
nor I_5964 (I107130,I86299,I86314);
nand I_5965 (I107147,I107130,I86302);
DFFARX1 I_5966  ( .D(I107147), .CLK(I5694_clk), .RSTB(I107096_rst), .Q(I107070) );
nor I_5967 (I107178,I107113,I86299);
nand I_5968 (I107195,I107178,I86305);
not I_5969 (I107085,I107195);
DFFARX1 I_5970  ( .D(I107195), .CLK(I5694_clk), .RSTB(I107096_rst), .Q(I107067) );
not I_5971 (I107240,I86299);
not I_5972 (I107257,I107240);
not I_5973 (I107274,I86311);
nor I_5974 (I107291,I107274,I86308);
and I_5975 (I107308,I107291,I86287);
or I_5976 (I107325,I107308,I86296);
DFFARX1 I_5977  ( .D(I107325), .CLK(I5694_clk), .RSTB(I107096_rst), .Q(I107342) );
nor I_5978 (I107359,I107342,I107195);
nor I_5979 (I107376,I107342,I107257);
nand I_5980 (I107082,I107147,I107376);
nand I_5981 (I107407,I107113,I86311);
nand I_5982 (I107424,I107407,I107342);
and I_5983 (I107441,I107407,I107424);
DFFARX1 I_5984  ( .D(I107441), .CLK(I5694_clk), .RSTB(I107096_rst), .Q(I107064) );
DFFARX1 I_5985  ( .D(I107407), .CLK(I5694_clk), .RSTB(I107096_rst), .Q(I107472) );
and I_5986 (I107061,I107240,I107472);
DFFARX1 I_5987  ( .D(I86293), .CLK(I5694_clk), .RSTB(I107096_rst), .Q(I107503) );
not I_5988 (I107520,I107503);
nor I_5989 (I107537,I107195,I107520);
and I_5990 (I107554,I107503,I107537);
nand I_5991 (I107076,I107503,I107257);
DFFARX1 I_5992  ( .D(I107503), .CLK(I5694_clk), .RSTB(I107096_rst), .Q(I107585) );
not I_5993 (I107073,I107585);
DFFARX1 I_5994  ( .D(I86290), .CLK(I5694_clk), .RSTB(I107096_rst), .Q(I107616) );
not I_5995 (I107633,I107616);
or I_5996 (I107650,I107633,I107554);
DFFARX1 I_5997  ( .D(I107650), .CLK(I5694_clk), .RSTB(I107096_rst), .Q(I107079) );
nand I_5998 (I107088,I107633,I107359);
DFFARX1 I_5999  ( .D(I107633), .CLK(I5694_clk), .RSTB(I107096_rst), .Q(I107058) );
not I_6000 (I107742_rst,I5701);
not I_6001 (I107759,I92445);
nor I_6002 (I107776,I92424,I92436);
nand I_6003 (I107793,I107776,I92430);
DFFARX1 I_6004  ( .D(I107793), .CLK(I5694_clk), .RSTB(I107742_rst), .Q(I107713) );
nor I_6005 (I107824,I107759,I92424);
nand I_6006 (I107841,I107824,I92451);
nand I_6007 (I107858,I107841,I107793);
not I_6008 (I107875,I92424);
not I_6009 (I107892,I92427);
nor I_6010 (I107909,I107892,I92439);
and I_6011 (I107926,I107909,I92442);
or I_6012 (I107943,I107926,I92448);
DFFARX1 I_6013  ( .D(I107943), .CLK(I5694_clk), .RSTB(I107742_rst), .Q(I107960) );
nor I_6014 (I107977,I107960,I107841);
nand I_6015 (I107728,I107875,I107977);
not I_6016 (I107725,I107960);
and I_6017 (I108022,I107960,I107858);
DFFARX1 I_6018  ( .D(I108022), .CLK(I5694_clk), .RSTB(I107742_rst), .Q(I107710) );
DFFARX1 I_6019  ( .D(I107960), .CLK(I5694_clk), .RSTB(I107742_rst), .Q(I108053) );
and I_6020 (I107707,I107875,I108053);
nand I_6021 (I108084,I107759,I92427);
not I_6022 (I108101,I108084);
nor I_6023 (I108118,I107960,I108101);
DFFARX1 I_6024  ( .D(I92421), .CLK(I5694_clk), .RSTB(I107742_rst), .Q(I108135) );
nand I_6025 (I108152,I108135,I108084);
and I_6026 (I108169,I107875,I108152);
DFFARX1 I_6027  ( .D(I108169), .CLK(I5694_clk), .RSTB(I107742_rst), .Q(I107734) );
not I_6028 (I108200,I108135);
nand I_6029 (I107722,I108135,I108118);
nand I_6030 (I107716,I108135,I108101);
DFFARX1 I_6031  ( .D(I92433), .CLK(I5694_clk), .RSTB(I107742_rst), .Q(I108245) );
not I_6032 (I108262,I108245);
nor I_6033 (I107731,I108135,I108262);
nor I_6034 (I108293,I108262,I108200);
and I_6035 (I108310,I107841,I108293);
or I_6036 (I108327,I108084,I108310);
DFFARX1 I_6037  ( .D(I108327), .CLK(I5694_clk), .RSTB(I107742_rst), .Q(I107719) );
DFFARX1 I_6038  ( .D(I108262), .CLK(I5694_clk), .RSTB(I107742_rst), .Q(I107704) );
not I_6039 (I108405_rst,I5701);
not I_6040 (I108422,I60853);
nor I_6041 (I108439,I60862,I60835);
nand I_6042 (I108456,I108439,I60847);
DFFARX1 I_6043  ( .D(I108456), .CLK(I5694_clk), .RSTB(I108405_rst), .Q(I108376) );
nor I_6044 (I108487,I108422,I60862);
nand I_6045 (I108504,I108487,I60859);
nand I_6046 (I108521,I108504,I108456);
not I_6047 (I108538,I60862);
not I_6048 (I108555,I60838);
nor I_6049 (I108572,I108555,I60844);
and I_6050 (I108589,I108572,I60856);
or I_6051 (I108606,I108589,I60841);
DFFARX1 I_6052  ( .D(I108606), .CLK(I5694_clk), .RSTB(I108405_rst), .Q(I108623) );
nor I_6053 (I108640,I108623,I108504);
nand I_6054 (I108391,I108538,I108640);
not I_6055 (I108388,I108623);
and I_6056 (I108685,I108623,I108521);
DFFARX1 I_6057  ( .D(I108685), .CLK(I5694_clk), .RSTB(I108405_rst), .Q(I108373) );
DFFARX1 I_6058  ( .D(I108623), .CLK(I5694_clk), .RSTB(I108405_rst), .Q(I108716) );
and I_6059 (I108370,I108538,I108716);
nand I_6060 (I108747,I108422,I60838);
not I_6061 (I108764,I108747);
nor I_6062 (I108781,I108623,I108764);
DFFARX1 I_6063  ( .D(I60865), .CLK(I5694_clk), .RSTB(I108405_rst), .Q(I108798) );
nand I_6064 (I108815,I108798,I108747);
and I_6065 (I108832,I108538,I108815);
DFFARX1 I_6066  ( .D(I108832), .CLK(I5694_clk), .RSTB(I108405_rst), .Q(I108397) );
not I_6067 (I108863,I108798);
nand I_6068 (I108385,I108798,I108781);
nand I_6069 (I108379,I108798,I108764);
DFFARX1 I_6070  ( .D(I60850), .CLK(I5694_clk), .RSTB(I108405_rst), .Q(I108908) );
not I_6071 (I108925,I108908);
nor I_6072 (I108394,I108798,I108925);
nor I_6073 (I108956,I108925,I108863);
and I_6074 (I108973,I108504,I108956);
or I_6075 (I108990,I108747,I108973);
DFFARX1 I_6076  ( .D(I108990), .CLK(I5694_clk), .RSTB(I108405_rst), .Q(I108382) );
DFFARX1 I_6077  ( .D(I108925), .CLK(I5694_clk), .RSTB(I108405_rst), .Q(I108367) );
not I_6078 (I109068_rst,I5701);
not I_6079 (I109085,I102551);
nor I_6080 (I109102,I102539,I102563);
nand I_6081 (I109119,I109102,I102548);
DFFARX1 I_6082  ( .D(I109119), .CLK(I5694_clk), .RSTB(I109068_rst), .Q(I109039) );
nor I_6083 (I109150,I109085,I102539);
nand I_6084 (I109167,I109150,I102566);
nand I_6085 (I109184,I109167,I109119);
not I_6086 (I109201,I102539);
not I_6087 (I109218,I102536);
nor I_6088 (I109235,I109218,I102545);
and I_6089 (I109252,I109235,I102560);
or I_6090 (I109269,I109252,I102542);
DFFARX1 I_6091  ( .D(I109269), .CLK(I5694_clk), .RSTB(I109068_rst), .Q(I109286) );
nor I_6092 (I109303,I109286,I109167);
nand I_6093 (I109054,I109201,I109303);
not I_6094 (I109051,I109286);
and I_6095 (I109348,I109286,I109184);
DFFARX1 I_6096  ( .D(I109348), .CLK(I5694_clk), .RSTB(I109068_rst), .Q(I109036) );
DFFARX1 I_6097  ( .D(I109286), .CLK(I5694_clk), .RSTB(I109068_rst), .Q(I109379) );
and I_6098 (I109033,I109201,I109379);
nand I_6099 (I109410,I109085,I102536);
not I_6100 (I109427,I109410);
nor I_6101 (I109444,I109286,I109427);
DFFARX1 I_6102  ( .D(I102557), .CLK(I5694_clk), .RSTB(I109068_rst), .Q(I109461) );
nand I_6103 (I109478,I109461,I109410);
and I_6104 (I109495,I109201,I109478);
DFFARX1 I_6105  ( .D(I109495), .CLK(I5694_clk), .RSTB(I109068_rst), .Q(I109060) );
not I_6106 (I109526,I109461);
nand I_6107 (I109048,I109461,I109444);
nand I_6108 (I109042,I109461,I109427);
DFFARX1 I_6109  ( .D(I102554), .CLK(I5694_clk), .RSTB(I109068_rst), .Q(I109571) );
not I_6110 (I109588,I109571);
nor I_6111 (I109057,I109461,I109588);
nor I_6112 (I109619,I109588,I109526);
and I_6113 (I109636,I109167,I109619);
or I_6114 (I109653,I109410,I109636);
DFFARX1 I_6115  ( .D(I109653), .CLK(I5694_clk), .RSTB(I109068_rst), .Q(I109045) );
DFFARX1 I_6116  ( .D(I109588), .CLK(I5694_clk), .RSTB(I109068_rst), .Q(I109030) );
not I_6117 (I109731_rst,I5701);
not I_6118 (I109748,I53661);
nor I_6119 (I109765,I53670,I53682);
nand I_6120 (I109782,I109765,I53673);
DFFARX1 I_6121  ( .D(I109782), .CLK(I5694_clk), .RSTB(I109731_rst), .Q(I109702) );
nor I_6122 (I109813,I109748,I53670);
nand I_6123 (I109830,I109813,I53685);
nand I_6124 (I109847,I109830,I109782);
not I_6125 (I109864,I53670);
not I_6126 (I109881,I53691);
nor I_6127 (I109898,I109881,I53667);
and I_6128 (I109915,I109898,I53676);
or I_6129 (I109932,I109915,I53664);
DFFARX1 I_6130  ( .D(I109932), .CLK(I5694_clk), .RSTB(I109731_rst), .Q(I109949) );
nor I_6131 (I109966,I109949,I109830);
nand I_6132 (I109717,I109864,I109966);
not I_6133 (I109714,I109949);
and I_6134 (I110011,I109949,I109847);
DFFARX1 I_6135  ( .D(I110011), .CLK(I5694_clk), .RSTB(I109731_rst), .Q(I109699) );
DFFARX1 I_6136  ( .D(I109949), .CLK(I5694_clk), .RSTB(I109731_rst), .Q(I110042) );
and I_6137 (I109696,I109864,I110042);
nand I_6138 (I110073,I109748,I53691);
not I_6139 (I110090,I110073);
nor I_6140 (I110107,I109949,I110090);
DFFARX1 I_6141  ( .D(I53688), .CLK(I5694_clk), .RSTB(I109731_rst), .Q(I110124) );
nand I_6142 (I110141,I110124,I110073);
and I_6143 (I110158,I109864,I110141);
DFFARX1 I_6144  ( .D(I110158), .CLK(I5694_clk), .RSTB(I109731_rst), .Q(I109723) );
not I_6145 (I110189,I110124);
nand I_6146 (I109711,I110124,I110107);
nand I_6147 (I109705,I110124,I110090);
DFFARX1 I_6148  ( .D(I53679), .CLK(I5694_clk), .RSTB(I109731_rst), .Q(I110234) );
not I_6149 (I110251,I110234);
nor I_6150 (I109720,I110124,I110251);
nor I_6151 (I110282,I110251,I110189);
and I_6152 (I110299,I109830,I110282);
or I_6153 (I110316,I110073,I110299);
DFFARX1 I_6154  ( .D(I110316), .CLK(I5694_clk), .RSTB(I109731_rst), .Q(I109708) );
DFFARX1 I_6155  ( .D(I110251), .CLK(I5694_clk), .RSTB(I109731_rst), .Q(I109693) );
not I_6156 (I110394_rst,I5701);
not I_6157 (I110411,I69471);
nor I_6158 (I110428,I69477,I69474);
nand I_6159 (I110445,I110428,I69492);
DFFARX1 I_6160  ( .D(I110445), .CLK(I5694_clk), .RSTB(I110394_rst), .Q(I110365) );
nor I_6161 (I110476,I110411,I69477);
nand I_6162 (I110493,I110476,I69501);
nand I_6163 (I110510,I110493,I110445);
not I_6164 (I110527,I69477);
not I_6165 (I110544,I69495);
nor I_6166 (I110561,I110544,I69486);
and I_6167 (I110578,I110561,I69489);
or I_6168 (I110595,I110578,I69480);
DFFARX1 I_6169  ( .D(I110595), .CLK(I5694_clk), .RSTB(I110394_rst), .Q(I110612) );
nor I_6170 (I110629,I110612,I110493);
nand I_6171 (I110380,I110527,I110629);
not I_6172 (I110377,I110612);
and I_6173 (I110674,I110612,I110510);
DFFARX1 I_6174  ( .D(I110674), .CLK(I5694_clk), .RSTB(I110394_rst), .Q(I110362) );
DFFARX1 I_6175  ( .D(I110612), .CLK(I5694_clk), .RSTB(I110394_rst), .Q(I110705) );
and I_6176 (I110359,I110527,I110705);
nand I_6177 (I110736,I110411,I69495);
not I_6178 (I110753,I110736);
nor I_6179 (I110770,I110612,I110753);
DFFARX1 I_6180  ( .D(I69498), .CLK(I5694_clk), .RSTB(I110394_rst), .Q(I110787) );
nand I_6181 (I110804,I110787,I110736);
and I_6182 (I110821,I110527,I110804);
DFFARX1 I_6183  ( .D(I110821), .CLK(I5694_clk), .RSTB(I110394_rst), .Q(I110386) );
not I_6184 (I110852,I110787);
nand I_6185 (I110374,I110787,I110770);
nand I_6186 (I110368,I110787,I110753);
DFFARX1 I_6187  ( .D(I69483), .CLK(I5694_clk), .RSTB(I110394_rst), .Q(I110897) );
not I_6188 (I110914,I110897);
nor I_6189 (I110383,I110787,I110914);
nor I_6190 (I110945,I110914,I110852);
and I_6191 (I110962,I110493,I110945);
or I_6192 (I110979,I110736,I110962);
DFFARX1 I_6193  ( .D(I110979), .CLK(I5694_clk), .RSTB(I110394_rst), .Q(I110371) );
DFFARX1 I_6194  ( .D(I110914), .CLK(I5694_clk), .RSTB(I110394_rst), .Q(I110356) );
not I_6195 (I111057_rst,I5701);
not I_6196 (I111074,I51672);
nor I_6197 (I111091,I51681,I51693);
nand I_6198 (I111108,I111091,I51684);
DFFARX1 I_6199  ( .D(I111108), .CLK(I5694_clk), .RSTB(I111057_rst), .Q(I111028) );
nor I_6200 (I111139,I111074,I51681);
nand I_6201 (I111156,I111139,I51696);
nand I_6202 (I111173,I111156,I111108);
not I_6203 (I111190,I51681);
not I_6204 (I111207,I51702);
nor I_6205 (I111224,I111207,I51678);
and I_6206 (I111241,I111224,I51687);
or I_6207 (I111258,I111241,I51675);
DFFARX1 I_6208  ( .D(I111258), .CLK(I5694_clk), .RSTB(I111057_rst), .Q(I111275) );
nor I_6209 (I111292,I111275,I111156);
nand I_6210 (I111043,I111190,I111292);
not I_6211 (I111040,I111275);
and I_6212 (I111337,I111275,I111173);
DFFARX1 I_6213  ( .D(I111337), .CLK(I5694_clk), .RSTB(I111057_rst), .Q(I111025) );
DFFARX1 I_6214  ( .D(I111275), .CLK(I5694_clk), .RSTB(I111057_rst), .Q(I111368) );
and I_6215 (I111022,I111190,I111368);
nand I_6216 (I111399,I111074,I51702);
not I_6217 (I111416,I111399);
nor I_6218 (I111433,I111275,I111416);
DFFARX1 I_6219  ( .D(I51699), .CLK(I5694_clk), .RSTB(I111057_rst), .Q(I111450) );
nand I_6220 (I111467,I111450,I111399);
and I_6221 (I111484,I111190,I111467);
DFFARX1 I_6222  ( .D(I111484), .CLK(I5694_clk), .RSTB(I111057_rst), .Q(I111049) );
not I_6223 (I111515,I111450);
nand I_6224 (I111037,I111450,I111433);
nand I_6225 (I111031,I111450,I111416);
DFFARX1 I_6226  ( .D(I51690), .CLK(I5694_clk), .RSTB(I111057_rst), .Q(I111560) );
not I_6227 (I111577,I111560);
nor I_6228 (I111046,I111450,I111577);
nor I_6229 (I111608,I111577,I111515);
and I_6230 (I111625,I111156,I111608);
or I_6231 (I111642,I111399,I111625);
DFFARX1 I_6232  ( .D(I111642), .CLK(I5694_clk), .RSTB(I111057_rst), .Q(I111034) );
DFFARX1 I_6233  ( .D(I111577), .CLK(I5694_clk), .RSTB(I111057_rst), .Q(I111019) );
not I_6234 (I111720_rst,I5701);
not I_6235 (I111737,I86925);
nor I_6236 (I111754,I86931,I86943);
nand I_6237 (I111771,I111754,I86934);
DFFARX1 I_6238  ( .D(I111771), .CLK(I5694_clk), .RSTB(I111720_rst), .Q(I111691) );
nor I_6239 (I111802,I111737,I86931);
nand I_6240 (I111819,I111802,I86913);
nand I_6241 (I111836,I111819,I111771);
not I_6242 (I111853,I86931);
not I_6243 (I111870,I86928);
nor I_6244 (I111887,I111870,I86916);
and I_6245 (I111904,I111887,I86937);
or I_6246 (I111921,I111904,I86919);
DFFARX1 I_6247  ( .D(I111921), .CLK(I5694_clk), .RSTB(I111720_rst), .Q(I111938) );
nor I_6248 (I111955,I111938,I111819);
nand I_6249 (I111706,I111853,I111955);
not I_6250 (I111703,I111938);
and I_6251 (I112000,I111938,I111836);
DFFARX1 I_6252  ( .D(I112000), .CLK(I5694_clk), .RSTB(I111720_rst), .Q(I111688) );
DFFARX1 I_6253  ( .D(I111938), .CLK(I5694_clk), .RSTB(I111720_rst), .Q(I112031) );
and I_6254 (I111685,I111853,I112031);
nand I_6255 (I112062,I111737,I86928);
not I_6256 (I112079,I112062);
nor I_6257 (I112096,I111938,I112079);
DFFARX1 I_6258  ( .D(I86940), .CLK(I5694_clk), .RSTB(I111720_rst), .Q(I112113) );
nand I_6259 (I112130,I112113,I112062);
and I_6260 (I112147,I111853,I112130);
DFFARX1 I_6261  ( .D(I112147), .CLK(I5694_clk), .RSTB(I111720_rst), .Q(I111712) );
not I_6262 (I112178,I112113);
nand I_6263 (I111700,I112113,I112096);
nand I_6264 (I111694,I112113,I112079);
DFFARX1 I_6265  ( .D(I86922), .CLK(I5694_clk), .RSTB(I111720_rst), .Q(I112223) );
not I_6266 (I112240,I112223);
nor I_6267 (I111709,I112113,I112240);
nor I_6268 (I112271,I112240,I112178);
and I_6269 (I112288,I111819,I112271);
or I_6270 (I112305,I112062,I112288);
DFFARX1 I_6271  ( .D(I112305), .CLK(I5694_clk), .RSTB(I111720_rst), .Q(I111697) );
DFFARX1 I_6272  ( .D(I112240), .CLK(I5694_clk), .RSTB(I111720_rst), .Q(I111682) );
not I_6273 (I112383_rst,I5701);
not I_6274 (I112400,I50346);
nor I_6275 (I112417,I50355,I50367);
nand I_6276 (I112434,I112417,I50358);
DFFARX1 I_6277  ( .D(I112434), .CLK(I5694_clk), .RSTB(I112383_rst), .Q(I112354) );
nor I_6278 (I112465,I112400,I50355);
nand I_6279 (I112482,I112465,I50370);
nand I_6280 (I112499,I112482,I112434);
not I_6281 (I112516,I50355);
not I_6282 (I112533,I50376);
nor I_6283 (I112550,I112533,I50352);
and I_6284 (I112567,I112550,I50361);
or I_6285 (I112584,I112567,I50349);
DFFARX1 I_6286  ( .D(I112584), .CLK(I5694_clk), .RSTB(I112383_rst), .Q(I112601) );
nor I_6287 (I112618,I112601,I112482);
nand I_6288 (I112369,I112516,I112618);
not I_6289 (I112366,I112601);
and I_6290 (I112663,I112601,I112499);
DFFARX1 I_6291  ( .D(I112663), .CLK(I5694_clk), .RSTB(I112383_rst), .Q(I112351) );
DFFARX1 I_6292  ( .D(I112601), .CLK(I5694_clk), .RSTB(I112383_rst), .Q(I112694) );
and I_6293 (I112348,I112516,I112694);
nand I_6294 (I112725,I112400,I50376);
not I_6295 (I112742,I112725);
nor I_6296 (I112759,I112601,I112742);
DFFARX1 I_6297  ( .D(I50373), .CLK(I5694_clk), .RSTB(I112383_rst), .Q(I112776) );
nand I_6298 (I112793,I112776,I112725);
and I_6299 (I112810,I112516,I112793);
DFFARX1 I_6300  ( .D(I112810), .CLK(I5694_clk), .RSTB(I112383_rst), .Q(I112375) );
not I_6301 (I112841,I112776);
nand I_6302 (I112363,I112776,I112759);
nand I_6303 (I112357,I112776,I112742);
DFFARX1 I_6304  ( .D(I50364), .CLK(I5694_clk), .RSTB(I112383_rst), .Q(I112886) );
not I_6305 (I112903,I112886);
nor I_6306 (I112372,I112776,I112903);
nor I_6307 (I112934,I112903,I112841);
and I_6308 (I112951,I112482,I112934);
or I_6309 (I112968,I112725,I112951);
DFFARX1 I_6310  ( .D(I112968), .CLK(I5694_clk), .RSTB(I112383_rst), .Q(I112360) );
DFFARX1 I_6311  ( .D(I112903), .CLK(I5694_clk), .RSTB(I112383_rst), .Q(I112345) );
not I_6312 (I113046_rst,I5701);
not I_6313 (I113063,I90711);
nor I_6314 (I113080,I90690,I90702);
nand I_6315 (I113097,I113080,I90696);
DFFARX1 I_6316  ( .D(I113097), .CLK(I5694_clk), .RSTB(I113046_rst), .Q(I113017) );
nor I_6317 (I113128,I113063,I90690);
nand I_6318 (I113145,I113128,I90717);
nand I_6319 (I113162,I113145,I113097);
not I_6320 (I113179,I90690);
not I_6321 (I113196,I90693);
nor I_6322 (I113213,I113196,I90705);
and I_6323 (I113230,I113213,I90708);
or I_6324 (I113247,I113230,I90714);
DFFARX1 I_6325  ( .D(I113247), .CLK(I5694_clk), .RSTB(I113046_rst), .Q(I113264) );
nor I_6326 (I113281,I113264,I113145);
nand I_6327 (I113032,I113179,I113281);
not I_6328 (I113029,I113264);
and I_6329 (I113326,I113264,I113162);
DFFARX1 I_6330  ( .D(I113326), .CLK(I5694_clk), .RSTB(I113046_rst), .Q(I113014) );
DFFARX1 I_6331  ( .D(I113264), .CLK(I5694_clk), .RSTB(I113046_rst), .Q(I113357) );
and I_6332 (I113011,I113179,I113357);
nand I_6333 (I113388,I113063,I90693);
not I_6334 (I113405,I113388);
nor I_6335 (I113422,I113264,I113405);
DFFARX1 I_6336  ( .D(I90687), .CLK(I5694_clk), .RSTB(I113046_rst), .Q(I113439) );
nand I_6337 (I113456,I113439,I113388);
and I_6338 (I113473,I113179,I113456);
DFFARX1 I_6339  ( .D(I113473), .CLK(I5694_clk), .RSTB(I113046_rst), .Q(I113038) );
not I_6340 (I113504,I113439);
nand I_6341 (I113026,I113439,I113422);
nand I_6342 (I113020,I113439,I113405);
DFFARX1 I_6343  ( .D(I90699), .CLK(I5694_clk), .RSTB(I113046_rst), .Q(I113549) );
not I_6344 (I113566,I113549);
nor I_6345 (I113035,I113439,I113566);
nor I_6346 (I113597,I113566,I113504);
and I_6347 (I113614,I113145,I113597);
or I_6348 (I113631,I113388,I113614);
DFFARX1 I_6349  ( .D(I113631), .CLK(I5694_clk), .RSTB(I113046_rst), .Q(I113023) );
DFFARX1 I_6350  ( .D(I113566), .CLK(I5694_clk), .RSTB(I113046_rst), .Q(I113008) );
not I_6351 (I113709_rst,I5701);
or I_6352 (I113726,I59561,I59558);
or I_6353 (I113743,I59543,I59561);
DFFARX1 I_6354  ( .D(I113743), .CLK(I5694_clk), .RSTB(I113709_rst), .Q(I113683) );
nor I_6355 (I113774,I59552,I59555);
not I_6356 (I113791,I113774);
not I_6357 (I113808,I59552);
and I_6358 (I113825,I113808,I59567);
nor I_6359 (I113842,I113825,I59558);
nor I_6360 (I113859,I59573,I59549);
DFFARX1 I_6361  ( .D(I113859), .CLK(I5694_clk), .RSTB(I113709_rst), .Q(I113876) );
nand I_6362 (I113893,I113876,I113726);
and I_6363 (I113910,I113842,I113893);
DFFARX1 I_6364  ( .D(I113910), .CLK(I5694_clk), .RSTB(I113709_rst), .Q(I113677) );
nor I_6365 (I113941,I59573,I59543);
DFFARX1 I_6366  ( .D(I113941), .CLK(I5694_clk), .RSTB(I113709_rst), .Q(I113958) );
and I_6367 (I113674,I113774,I113958);
DFFARX1 I_6368  ( .D(I59564), .CLK(I5694_clk), .RSTB(I113709_rst), .Q(I113989) );
and I_6369 (I114006,I113989,I59570);
DFFARX1 I_6370  ( .D(I114006), .CLK(I5694_clk), .RSTB(I113709_rst), .Q(I114023) );
not I_6371 (I113686,I114023);
DFFARX1 I_6372  ( .D(I114006), .CLK(I5694_clk), .RSTB(I113709_rst), .Q(I113671) );
DFFARX1 I_6373  ( .D(I59546), .CLK(I5694_clk), .RSTB(I113709_rst), .Q(I114068) );
not I_6374 (I114085,I114068);
nor I_6375 (I114102,I113743,I114085);
and I_6376 (I114119,I114006,I114102);
or I_6377 (I114136,I113726,I114119);
DFFARX1 I_6378  ( .D(I114136), .CLK(I5694_clk), .RSTB(I113709_rst), .Q(I113692) );
nor I_6379 (I114167,I114068,I113876);
nand I_6380 (I113701,I113842,I114167);
nor I_6381 (I114198,I114068,I113791);
nand I_6382 (I113695,I113941,I114198);
not I_6383 (I113698,I114068);
nand I_6384 (I113689,I114068,I113791);
DFFARX1 I_6385  ( .D(I114068), .CLK(I5694_clk), .RSTB(I113709_rst), .Q(I113680) );
not I_6386 (I114304_rst,I5701);
or I_6387 (I114321,I89432,I89429);
or I_6388 (I114338,I89459,I89432);
DFFARX1 I_6389  ( .D(I114338), .CLK(I5694_clk), .RSTB(I114304_rst), .Q(I114278) );
nor I_6390 (I114369,I89438,I89444);
not I_6391 (I114386,I114369);
not I_6392 (I114403,I89438);
and I_6393 (I114420,I114403,I89435);
nor I_6394 (I114437,I114420,I89429);
nor I_6395 (I114454,I89447,I89456);
DFFARX1 I_6396  ( .D(I114454), .CLK(I5694_clk), .RSTB(I114304_rst), .Q(I114471) );
nand I_6397 (I114488,I114471,I114321);
and I_6398 (I114505,I114437,I114488);
DFFARX1 I_6399  ( .D(I114505), .CLK(I5694_clk), .RSTB(I114304_rst), .Q(I114272) );
nor I_6400 (I114536,I89447,I89459);
DFFARX1 I_6401  ( .D(I114536), .CLK(I5694_clk), .RSTB(I114304_rst), .Q(I114553) );
and I_6402 (I114269,I114369,I114553);
DFFARX1 I_6403  ( .D(I89450), .CLK(I5694_clk), .RSTB(I114304_rst), .Q(I114584) );
and I_6404 (I114601,I114584,I89441);
DFFARX1 I_6405  ( .D(I114601), .CLK(I5694_clk), .RSTB(I114304_rst), .Q(I114618) );
not I_6406 (I114281,I114618);
DFFARX1 I_6407  ( .D(I114601), .CLK(I5694_clk), .RSTB(I114304_rst), .Q(I114266) );
DFFARX1 I_6408  ( .D(I89453), .CLK(I5694_clk), .RSTB(I114304_rst), .Q(I114663) );
not I_6409 (I114680,I114663);
nor I_6410 (I114697,I114338,I114680);
and I_6411 (I114714,I114601,I114697);
or I_6412 (I114731,I114321,I114714);
DFFARX1 I_6413  ( .D(I114731), .CLK(I5694_clk), .RSTB(I114304_rst), .Q(I114287) );
nor I_6414 (I114762,I114663,I114471);
nand I_6415 (I114296,I114437,I114762);
nor I_6416 (I114793,I114663,I114386);
nand I_6417 (I114290,I114536,I114793);
not I_6418 (I114293,I114663);
nand I_6419 (I114284,I114663,I114386);
DFFARX1 I_6420  ( .D(I114663), .CLK(I5694_clk), .RSTB(I114304_rst), .Q(I114275) );
not I_6421 (I114899_rst,I5701);
or I_6422 (I114916,I95876,I95885);
or I_6423 (I114933,I95879,I95876);
DFFARX1 I_6424  ( .D(I114933), .CLK(I5694_clk), .RSTB(I114899_rst), .Q(I114873) );
nor I_6425 (I114964,I95855,I95858);
not I_6426 (I114981,I114964);
not I_6427 (I114998,I95855);
and I_6428 (I115015,I114998,I95867);
nor I_6429 (I115032,I115015,I95885);
nor I_6430 (I115049,I95873,I95864);
DFFARX1 I_6431  ( .D(I115049), .CLK(I5694_clk), .RSTB(I114899_rst), .Q(I115066) );
nand I_6432 (I115083,I115066,I114916);
and I_6433 (I115100,I115032,I115083);
DFFARX1 I_6434  ( .D(I115100), .CLK(I5694_clk), .RSTB(I114899_rst), .Q(I114867) );
nor I_6435 (I115131,I95873,I95879);
DFFARX1 I_6436  ( .D(I115131), .CLK(I5694_clk), .RSTB(I114899_rst), .Q(I115148) );
and I_6437 (I114864,I114964,I115148);
DFFARX1 I_6438  ( .D(I95870), .CLK(I5694_clk), .RSTB(I114899_rst), .Q(I115179) );
and I_6439 (I115196,I115179,I95861);
DFFARX1 I_6440  ( .D(I115196), .CLK(I5694_clk), .RSTB(I114899_rst), .Q(I115213) );
not I_6441 (I114876,I115213);
DFFARX1 I_6442  ( .D(I115196), .CLK(I5694_clk), .RSTB(I114899_rst), .Q(I114861) );
DFFARX1 I_6443  ( .D(I95882), .CLK(I5694_clk), .RSTB(I114899_rst), .Q(I115258) );
not I_6444 (I115275,I115258);
nor I_6445 (I115292,I114933,I115275);
and I_6446 (I115309,I115196,I115292);
or I_6447 (I115326,I114916,I115309);
DFFARX1 I_6448  ( .D(I115326), .CLK(I5694_clk), .RSTB(I114899_rst), .Q(I11488_rst2) );
nor I_6449 (I115357,I115258,I115066);
nand I_6450 (I114891,I115032,I115357);
nor I_6451 (I115388,I115258,I114981);
nand I_6452 (I11488_rst5,I115131,I115388);
not I_6453 (I11488_rst8,I115258);
nand I_6454 (I114879,I115258,I114981);
DFFARX1 I_6455  ( .D(I115258), .CLK(I5694_clk), .RSTB(I114899_rst), .Q(I114870) );
not I_6456 (I115494_rst,I5701);
or I_6457 (I115511,I98681,I98675);
or I_6458 (I115528,I98669,I98681);
DFFARX1 I_6459  ( .D(I115528), .CLK(I5694_clk), .RSTB(I115494_rst), .Q(I115468) );
nor I_6460 (I115559,I98687,I98678);
not I_6461 (I115576,I115559);
not I_6462 (I115593,I98687);
and I_6463 (I115610,I115593,I98684);
nor I_6464 (I115627,I115610,I98675);
nor I_6465 (I115644,I98660,I98666);
DFFARX1 I_6466  ( .D(I115644), .CLK(I5694_clk), .RSTB(I115494_rst), .Q(I115661) );
nand I_6467 (I115678,I115661,I115511);
and I_6468 (I115695,I115627,I115678);
DFFARX1 I_6469  ( .D(I115695), .CLK(I5694_clk), .RSTB(I115494_rst), .Q(I115462) );
nor I_6470 (I115726,I98660,I98669);
DFFARX1 I_6471  ( .D(I115726), .CLK(I5694_clk), .RSTB(I115494_rst), .Q(I115743) );
and I_6472 (I115459,I115559,I115743);
DFFARX1 I_6473  ( .D(I98672), .CLK(I5694_clk), .RSTB(I115494_rst), .Q(I115774) );
and I_6474 (I115791,I115774,I98690);
DFFARX1 I_6475  ( .D(I115791), .CLK(I5694_clk), .RSTB(I115494_rst), .Q(I115808) );
not I_6476 (I115471,I115808);
DFFARX1 I_6477  ( .D(I115791), .CLK(I5694_clk), .RSTB(I115494_rst), .Q(I115456) );
DFFARX1 I_6478  ( .D(I98663), .CLK(I5694_clk), .RSTB(I115494_rst), .Q(I115853) );
not I_6479 (I115870,I115853);
nor I_6480 (I115887,I115528,I115870);
and I_6481 (I115904,I115791,I115887);
or I_6482 (I115921,I115511,I115904);
DFFARX1 I_6483  ( .D(I115921), .CLK(I5694_clk), .RSTB(I115494_rst), .Q(I115477) );
nor I_6484 (I115952,I115853,I115661);
nand I_6485 (I115486,I115627,I115952);
nor I_6486 (I115983,I115853,I115576);
nand I_6487 (I115480,I115726,I115983);
not I_6488 (I115483,I115853);
nand I_6489 (I115474,I115853,I115576);
DFFARX1 I_6490  ( .D(I115853), .CLK(I5694_clk), .RSTB(I115494_rst), .Q(I115465) );
not I_6491 (I116089_rst,I5701);
or I_6492 (I116106,I56331,I56328);
or I_6493 (I116123,I56313,I56331);
DFFARX1 I_6494  ( .D(I116123), .CLK(I5694_clk), .RSTB(I116089_rst), .Q(I116063) );
nor I_6495 (I116154,I56322,I56325);
not I_6496 (I116171,I116154);
not I_6497 (I116188,I56322);
and I_6498 (I116205,I116188,I56337);
nor I_6499 (I116222,I116205,I56328);
nor I_6500 (I116239,I56343,I56319);
DFFARX1 I_6501  ( .D(I116239), .CLK(I5694_clk), .RSTB(I116089_rst), .Q(I116256) );
nand I_6502 (I116273,I116256,I116106);
and I_6503 (I116290,I116222,I116273);
DFFARX1 I_6504  ( .D(I116290), .CLK(I5694_clk), .RSTB(I116089_rst), .Q(I116057) );
nor I_6505 (I116321,I56343,I56313);
DFFARX1 I_6506  ( .D(I116321), .CLK(I5694_clk), .RSTB(I116089_rst), .Q(I116338) );
and I_6507 (I116054,I116154,I116338);
DFFARX1 I_6508  ( .D(I56334), .CLK(I5694_clk), .RSTB(I116089_rst), .Q(I116369) );
and I_6509 (I116386,I116369,I56340);
DFFARX1 I_6510  ( .D(I116386), .CLK(I5694_clk), .RSTB(I116089_rst), .Q(I116403) );
not I_6511 (I116066,I116403);
DFFARX1 I_6512  ( .D(I116386), .CLK(I5694_clk), .RSTB(I116089_rst), .Q(I116051) );
DFFARX1 I_6513  ( .D(I56316), .CLK(I5694_clk), .RSTB(I116089_rst), .Q(I116448) );
not I_6514 (I116465,I116448);
nor I_6515 (I116482,I116123,I116465);
and I_6516 (I116499,I116386,I116482);
or I_6517 (I116516,I116106,I116499);
DFFARX1 I_6518  ( .D(I116516), .CLK(I5694_clk), .RSTB(I116089_rst), .Q(I116072) );
nor I_6519 (I116547,I116448,I116256);
nand I_6520 (I116081,I116222,I116547);
nor I_6521 (I116578,I116448,I116171);
nand I_6522 (I116075,I116321,I116578);
not I_6523 (I116078,I116448);
nand I_6524 (I116069,I116448,I116171);
DFFARX1 I_6525  ( .D(I116448), .CLK(I5694_clk), .RSTB(I116089_rst), .Q(I116060) );
not I_6526 (I116684_rst,I5701);
or I_6527 (I116701,I72410,I72395);
or I_6528 (I116718,I72416,I72410);
DFFARX1 I_6529  ( .D(I116718), .CLK(I5694_clk), .RSTB(I116684_rst), .Q(I116658) );
nor I_6530 (I116749,I72422,I72404);
not I_6531 (I116766,I116749);
not I_6532 (I116783,I72422);
and I_6533 (I116800,I116783,I72401);
nor I_6534 (I116817,I116800,I72395);
nor I_6535 (I116834,I72398,I72407);
DFFARX1 I_6536  ( .D(I116834), .CLK(I5694_clk), .RSTB(I116684_rst), .Q(I116851) );
nand I_6537 (I116868,I116851,I116701);
and I_6538 (I116885,I116817,I116868);
DFFARX1 I_6539  ( .D(I116885), .CLK(I5694_clk), .RSTB(I116684_rst), .Q(I116652) );
nor I_6540 (I116916,I72398,I72416);
DFFARX1 I_6541  ( .D(I116916), .CLK(I5694_clk), .RSTB(I116684_rst), .Q(I116933) );
and I_6542 (I116649,I116749,I116933);
DFFARX1 I_6543  ( .D(I72425), .CLK(I5694_clk), .RSTB(I116684_rst), .Q(I116964) );
and I_6544 (I116981,I116964,I72413);
DFFARX1 I_6545  ( .D(I116981), .CLK(I5694_clk), .RSTB(I116684_rst), .Q(I116998) );
not I_6546 (I116661,I116998);
DFFARX1 I_6547  ( .D(I116981), .CLK(I5694_clk), .RSTB(I116684_rst), .Q(I116646) );
DFFARX1 I_6548  ( .D(I72419), .CLK(I5694_clk), .RSTB(I116684_rst), .Q(I117043) );
not I_6549 (I117060,I117043);
nor I_6550 (I117077,I116718,I117060);
and I_6551 (I117094,I116981,I117077);
or I_6552 (I117111,I116701,I117094);
DFFARX1 I_6553  ( .D(I117111), .CLK(I5694_clk), .RSTB(I116684_rst), .Q(I116667) );
nor I_6554 (I117142,I117043,I116851);
nand I_6555 (I116676,I116817,I117142);
nor I_6556 (I117173,I117043,I116766);
nand I_6557 (I116670,I116916,I117173);
not I_6558 (I116673,I117043);
nand I_6559 (I116664,I117043,I116766);
DFFARX1 I_6560  ( .D(I117043), .CLK(I5694_clk), .RSTB(I116684_rst), .Q(I116655) );
not I_6561 (I117279_rst,I5701);
or I_6562 (I117296,I80737,I80731);
or I_6563 (I117313,I80725,I80737);
DFFARX1 I_6564  ( .D(I117313), .CLK(I5694_clk), .RSTB(I117279_rst), .Q(I117253) );
nor I_6565 (I117344,I80728,I80734);
not I_6566 (I117361,I117344);
not I_6567 (I117378,I80728);
and I_6568 (I117395,I117378,I80752);
nor I_6569 (I117412,I117395,I80731);
nor I_6570 (I117429,I80755,I80746);
DFFARX1 I_6571  ( .D(I117429), .CLK(I5694_clk), .RSTB(I117279_rst), .Q(I117446) );
nand I_6572 (I117463,I117446,I117296);
and I_6573 (I117480,I117412,I117463);
DFFARX1 I_6574  ( .D(I117480), .CLK(I5694_clk), .RSTB(I117279_rst), .Q(I117247) );
nor I_6575 (I117511,I80755,I80725);
DFFARX1 I_6576  ( .D(I117511), .CLK(I5694_clk), .RSTB(I117279_rst), .Q(I117528) );
and I_6577 (I117244,I117344,I117528);
DFFARX1 I_6578  ( .D(I80743), .CLK(I5694_clk), .RSTB(I117279_rst), .Q(I117559) );
and I_6579 (I117576,I117559,I80740);
DFFARX1 I_6580  ( .D(I117576), .CLK(I5694_clk), .RSTB(I117279_rst), .Q(I117593) );
not I_6581 (I117256,I117593);
DFFARX1 I_6582  ( .D(I117576), .CLK(I5694_clk), .RSTB(I117279_rst), .Q(I117241) );
DFFARX1 I_6583  ( .D(I80749), .CLK(I5694_clk), .RSTB(I117279_rst), .Q(I117638) );
not I_6584 (I117655,I117638);
nor I_6585 (I117672,I117313,I117655);
and I_6586 (I117689,I117576,I117672);
or I_6587 (I117706,I117296,I117689);
DFFARX1 I_6588  ( .D(I117706), .CLK(I5694_clk), .RSTB(I117279_rst), .Q(I117262) );
nor I_6589 (I117737,I117638,I117446);
nand I_6590 (I117271,I117412,I117737);
nor I_6591 (I117768,I117638,I117361);
nand I_6592 (I117265,I117511,I117768);
not I_6593 (I117268,I117638);
nand I_6594 (I117259,I117638,I117361);
DFFARX1 I_6595  ( .D(I117638), .CLK(I5694_clk), .RSTB(I117279_rst), .Q(I117250) );
not I_6596 (I117874_rst,I5701);
or I_6597 (I117891,I91843,I91861);
or I_6598 (I117908,I91846,I91843);
DFFARX1 I_6599  ( .D(I117908), .CLK(I5694_clk), .RSTB(I117874_rst), .Q(I117848) );
nor I_6600 (I117939,I91855,I91858);
not I_6601 (I117956,I117939);
not I_6602 (I117973,I91855);
and I_6603 (I117990,I117973,I91864);
nor I_6604 (I118007,I117990,I91861);
nor I_6605 (I118024,I91870,I91849);
DFFARX1 I_6606  ( .D(I118024), .CLK(I5694_clk), .RSTB(I117874_rst), .Q(I118041) );
nand I_6607 (I118058,I118041,I117891);
and I_6608 (I118075,I118007,I118058);
DFFARX1 I_6609  ( .D(I118075), .CLK(I5694_clk), .RSTB(I117874_rst), .Q(I117842) );
nor I_6610 (I118106,I91870,I91846);
DFFARX1 I_6611  ( .D(I118106), .CLK(I5694_clk), .RSTB(I117874_rst), .Q(I118123) );
and I_6612 (I117839,I117939,I118123);
DFFARX1 I_6613  ( .D(I91873), .CLK(I5694_clk), .RSTB(I117874_rst), .Q(I118154) );
and I_6614 (I118171,I118154,I91867);
DFFARX1 I_6615  ( .D(I118171), .CLK(I5694_clk), .RSTB(I117874_rst), .Q(I118188) );
not I_6616 (I117851,I118188);
DFFARX1 I_6617  ( .D(I118171), .CLK(I5694_clk), .RSTB(I117874_rst), .Q(I117836) );
DFFARX1 I_6618  ( .D(I91852), .CLK(I5694_clk), .RSTB(I117874_rst), .Q(I118233) );
not I_6619 (I118250,I118233);
nor I_6620 (I118267,I117908,I118250);
and I_6621 (I118284,I118171,I118267);
or I_6622 (I118301,I117891,I118284);
DFFARX1 I_6623  ( .D(I118301), .CLK(I5694_clk), .RSTB(I117874_rst), .Q(I117857) );
nor I_6624 (I118332,I118233,I118041);
nand I_6625 (I117866,I118007,I118332);
nor I_6626 (I118363,I118233,I117956);
nand I_6627 (I117860,I118106,I118363);
not I_6628 (I117863,I118233);
nand I_6629 (I117854,I118233,I117956);
DFFARX1 I_6630  ( .D(I118233), .CLK(I5694_clk), .RSTB(I117874_rst), .Q(I117845) );
not I_6631 (I118469_rst,I5701);
or I_6632 (I118486,I91286,I91268);
not I_6633 (I118452,I118486);
DFFARX1 I_6634  ( .D(I118486), .CLK(I5694_clk), .RSTB(I118469_rst), .Q(I118431) );
or I_6635 (I118531,I91295,I91286);
nor I_6636 (I118548,I91277,I91292);
nor I_6637 (I118565,I118548,I118486);
not I_6638 (I118582,I91277);
and I_6639 (I118599,I118582,I91274);
nor I_6640 (I118616,I118599,I91268);
DFFARX1 I_6641  ( .D(I118616), .CLK(I5694_clk), .RSTB(I118469_rst), .Q(I118633) );
nor I_6642 (I118650,I91289,I91265);
DFFARX1 I_6643  ( .D(I118650), .CLK(I5694_clk), .RSTB(I118469_rst), .Q(I118667) );
nor I_6644 (I118458,I118667,I118616);
not I_6645 (I118698,I118667);
nor I_6646 (I118715,I91289,I91295);
nand I_6647 (I118732,I118616,I118715);
and I_6648 (I118749,I118531,I118732);
DFFARX1 I_6649  ( .D(I118749), .CLK(I5694_clk), .RSTB(I118469_rst), .Q(I118461) );
DFFARX1 I_6650  ( .D(I91283), .CLK(I5694_clk), .RSTB(I118469_rst), .Q(I118780) );
and I_6651 (I118797,I118780,I91271);
nor I_6652 (I118814,I118797,I118698);
and I_6653 (I118831,I118715,I118814);
or I_6654 (I118848,I118548,I118831);
DFFARX1 I_6655  ( .D(I118848), .CLK(I5694_clk), .RSTB(I118469_rst), .Q(I118446) );
not I_6656 (I118879,I118797);
nor I_6657 (I118896,I118486,I118879);
nand I_6658 (I118449,I118531,I118896);
nand I_6659 (I118443,I118667,I118879);
DFFARX1 I_6660  ( .D(I118797), .CLK(I5694_clk), .RSTB(I118469_rst), .Q(I118437) );
DFFARX1 I_6661  ( .D(I91280), .CLK(I5694_clk), .RSTB(I118469_rst), .Q(I118955) );
nand I_6662 (I118455,I118955,I118565);
DFFARX1 I_6663  ( .D(I118955), .CLK(I5694_clk), .RSTB(I118469_rst), .Q(I118986) );
not I_6664 (I118440,I118986);
and I_6665 (I118434,I118955,I118633);
not I_6666 (I119064_rst,I5701);
not I_6667 (I119081,I64723);
nor I_6668 (I119098,I64720,I64738);
nand I_6669 (I119115,I119098,I64741);
nor I_6670 (I119132,I119081,I64720);
nand I_6671 (I119149,I119132,I64726);
not I_6672 (I119166,I119149);
not I_6673 (I119183,I64720);
nor I_6674 (I119053,I119149,I119183);
not I_6675 (I119214,I119183);
nand I_6676 (I119038,I119149,I119214);
not I_6677 (I119245,I64735);
nor I_6678 (I119262,I119245,I64717);
and I_6679 (I119279,I119262,I64711);
or I_6680 (I119296,I119279,I64729);
DFFARX1 I_6681  ( .D(I119296), .CLK(I5694_clk), .RSTB(I119064_rst), .Q(I119313) );
nor I_6682 (I119330,I119313,I119166);
DFFARX1 I_6683  ( .D(I119313), .CLK(I5694_clk), .RSTB(I119064_rst), .Q(I119347) );
not I_6684 (I119035,I119347);
nand I_6685 (I119378,I119081,I64735);
and I_6686 (I119395,I119378,I119330);
DFFARX1 I_6687  ( .D(I119378), .CLK(I5694_clk), .RSTB(I119064_rst), .Q(I119032) );
DFFARX1 I_6688  ( .D(I64714), .CLK(I5694_clk), .RSTB(I119064_rst), .Q(I119426) );
nor I_6689 (I119443,I119426,I119149);
nand I_6690 (I119050,I119313,I119443);
nor I_6691 (I119474,I119426,I119214);
not I_6692 (I119047,I119426);
nand I_6693 (I119505,I119426,I119115);
and I_6694 (I119522,I119183,I119505);
DFFARX1 I_6695  ( .D(I119522), .CLK(I5694_clk), .RSTB(I119064_rst), .Q(I119026) );
DFFARX1 I_6696  ( .D(I119426), .CLK(I5694_clk), .RSTB(I119064_rst), .Q(I119029) );
DFFARX1 I_6697  ( .D(I64732), .CLK(I5694_clk), .RSTB(I119064_rst), .Q(I119567) );
not I_6698 (I119584,I119567);
nand I_6699 (I119601,I119584,I119149);
and I_6700 (I119618,I119378,I119601);
DFFARX1 I_6701  ( .D(I119618), .CLK(I5694_clk), .RSTB(I119064_rst), .Q(I119056) );
or I_6702 (I119649,I119584,I119395);
DFFARX1 I_6703  ( .D(I119649), .CLK(I5694_clk), .RSTB(I119064_rst), .Q(I119041) );
nand I_6704 (I119044,I119584,I119474);
not I_6705 (I119727_rst,I5701);
not I_6706 (I119744,I99312);
nor I_6707 (I119761,I99309,I99333);
nand I_6708 (I119778,I119761,I99330);
nor I_6709 (I119795,I119744,I99309);
nand I_6710 (I119812,I119795,I99336);
not I_6711 (I119829,I119812);
not I_6712 (I119846,I99309);
nor I_6713 (I119716,I119812,I119846);
not I_6714 (I119877,I119846);
nand I_6715 (I119701,I119812,I119877);
not I_6716 (I119908,I99327);
nor I_6717 (I119925,I119908,I99318);
and I_6718 (I119942,I119925,I99315);
or I_6719 (I119959,I119942,I99324);
DFFARX1 I_6720  ( .D(I119959), .CLK(I5694_clk), .RSTB(I119727_rst), .Q(I119976) );
nor I_6721 (I119993,I119976,I119829);
DFFARX1 I_6722  ( .D(I119976), .CLK(I5694_clk), .RSTB(I119727_rst), .Q(I120010) );
not I_6723 (I119698,I120010);
nand I_6724 (I120041,I119744,I99327);
and I_6725 (I120058,I120041,I119993);
DFFARX1 I_6726  ( .D(I120041), .CLK(I5694_clk), .RSTB(I119727_rst), .Q(I119695) );
DFFARX1 I_6727  ( .D(I99306), .CLK(I5694_clk), .RSTB(I119727_rst), .Q(I120089) );
nor I_6728 (I120106,I120089,I119812);
nand I_6729 (I119713,I119976,I120106);
nor I_6730 (I120137,I120089,I119877);
not I_6731 (I119710,I120089);
nand I_6732 (I120168,I120089,I119778);
and I_6733 (I120185,I119846,I120168);
DFFARX1 I_6734  ( .D(I120185), .CLK(I5694_clk), .RSTB(I119727_rst), .Q(I119689) );
DFFARX1 I_6735  ( .D(I120089), .CLK(I5694_clk), .RSTB(I119727_rst), .Q(I119692) );
DFFARX1 I_6736  ( .D(I99321), .CLK(I5694_clk), .RSTB(I119727_rst), .Q(I120230) );
not I_6737 (I120247,I120230);
nand I_6738 (I120264,I120247,I119812);
and I_6739 (I120281,I120041,I120264);
DFFARX1 I_6740  ( .D(I120281), .CLK(I5694_clk), .RSTB(I119727_rst), .Q(I119719) );
or I_6741 (I120312,I120247,I120058);
DFFARX1 I_6742  ( .D(I120312), .CLK(I5694_clk), .RSTB(I119727_rst), .Q(I119704) );
nand I_6743 (I119707,I120247,I120137);
not I_6744 (I120390_rst,I5701);
not I_6745 (I120407,I107064);
nor I_6746 (I120424,I107061,I107085);
nand I_6747 (I120441,I120424,I107082);
nor I_6748 (I120458,I120407,I107061);
nand I_6749 (I120475,I120458,I107088);
not I_6750 (I120492,I120475);
not I_6751 (I120509,I107061);
nor I_6752 (I120379,I120475,I120509);
not I_6753 (I120540,I120509);
nand I_6754 (I120364,I120475,I120540);
not I_6755 (I120571,I107079);
nor I_6756 (I120588,I120571,I107070);
and I_6757 (I120605,I120588,I107067);
or I_6758 (I120622,I120605,I107076);
DFFARX1 I_6759  ( .D(I120622), .CLK(I5694_clk), .RSTB(I120390_rst), .Q(I120639) );
nor I_6760 (I120656,I120639,I120492);
DFFARX1 I_6761  ( .D(I120639), .CLK(I5694_clk), .RSTB(I120390_rst), .Q(I120673) );
not I_6762 (I120361,I120673);
nand I_6763 (I120704,I120407,I107079);
and I_6764 (I120721,I120704,I120656);
DFFARX1 I_6765  ( .D(I120704), .CLK(I5694_clk), .RSTB(I120390_rst), .Q(I120358) );
DFFARX1 I_6766  ( .D(I107058), .CLK(I5694_clk), .RSTB(I120390_rst), .Q(I120752) );
nor I_6767 (I120769,I120752,I120475);
nand I_6768 (I120376,I120639,I120769);
nor I_6769 (I120800,I120752,I120540);
not I_6770 (I120373,I120752);
nand I_6771 (I12083_rst1,I120752,I120441);
and I_6772 (I120848,I120509,I12083_rst1);
DFFARX1 I_6773  ( .D(I120848), .CLK(I5694_clk), .RSTB(I120390_rst), .Q(I120352) );
DFFARX1 I_6774  ( .D(I120752), .CLK(I5694_clk), .RSTB(I120390_rst), .Q(I120355) );
DFFARX1 I_6775  ( .D(I107073), .CLK(I5694_clk), .RSTB(I120390_rst), .Q(I120893) );
not I_6776 (I120910,I120893);
nand I_6777 (I120927,I120910,I120475);
and I_6778 (I120944,I120704,I120927);
DFFARX1 I_6779  ( .D(I120944), .CLK(I5694_clk), .RSTB(I120390_rst), .Q(I120382) );
or I_6780 (I120975,I120910,I120721);
DFFARX1 I_6781  ( .D(I120975), .CLK(I5694_clk), .RSTB(I120390_rst), .Q(I120367) );
nand I_6782 (I120370,I120910,I120800);
not I_6783 (I121053_rst,I5701);
not I_6784 (I121070,I62785);
nor I_6785 (I121087,I62782,I62800);
nand I_6786 (I121104,I121087,I62803);
nor I_6787 (I121121,I121070,I62782);
nand I_6788 (I121138,I121121,I62788);
not I_6789 (I121155,I121138);
not I_6790 (I121172,I62782);
nor I_6791 (I121042,I121138,I121172);
not I_6792 (I121203,I121172);
nand I_6793 (I121027,I121138,I121203);
not I_6794 (I121234,I62797);
nor I_6795 (I121251,I121234,I62779);
and I_6796 (I121268,I121251,I62773);
or I_6797 (I121285,I121268,I62791);
DFFARX1 I_6798  ( .D(I121285), .CLK(I5694_clk), .RSTB(I121053_rst), .Q(I121302) );
nor I_6799 (I121319,I121302,I121155);
DFFARX1 I_6800  ( .D(I121302), .CLK(I5694_clk), .RSTB(I121053_rst), .Q(I121336) );
not I_6801 (I121024,I121336);
nand I_6802 (I121367,I121070,I62797);
and I_6803 (I121384,I121367,I121319);
DFFARX1 I_6804  ( .D(I121367), .CLK(I5694_clk), .RSTB(I121053_rst), .Q(I121021) );
DFFARX1 I_6805  ( .D(I62776), .CLK(I5694_clk), .RSTB(I121053_rst), .Q(I121415) );
nor I_6806 (I121432,I121415,I121138);
nand I_6807 (I121039,I121302,I121432);
nor I_6808 (I121463,I121415,I121203);
not I_6809 (I121036,I121415);
nand I_6810 (I121494,I121415,I121104);
and I_6811 (I121511,I121172,I121494);
DFFARX1 I_6812  ( .D(I121511), .CLK(I5694_clk), .RSTB(I121053_rst), .Q(I121015) );
DFFARX1 I_6813  ( .D(I121415), .CLK(I5694_clk), .RSTB(I121053_rst), .Q(I121018) );
DFFARX1 I_6814  ( .D(I62794), .CLK(I5694_clk), .RSTB(I121053_rst), .Q(I121556) );
not I_6815 (I121573,I121556);
nand I_6816 (I121590,I121573,I121138);
and I_6817 (I121607,I121367,I121590);
DFFARX1 I_6818  ( .D(I121607), .CLK(I5694_clk), .RSTB(I121053_rst), .Q(I121045) );
or I_6819 (I121638,I121573,I121384);
DFFARX1 I_6820  ( .D(I121638), .CLK(I5694_clk), .RSTB(I121053_rst), .Q(I121030) );
nand I_6821 (I121033,I121573,I121463);
not I_6822 (I121716_rst,I5701);
not I_6823 (I121733,I75388);
nor I_6824 (I121750,I75397,I75379);
nand I_6825 (I121767,I121750,I75400);
nor I_6826 (I121784,I121733,I75397);
nand I_6827 (I121801,I121784,I75391);
not I_6828 (I121818,I121801);
not I_6829 (I121835,I75397);
nor I_6830 (I121705,I121801,I121835);
not I_6831 (I121866,I121835);
nand I_6832 (I121690,I121801,I121866);
not I_6833 (I121897,I75385);
nor I_6834 (I121914,I121897,I75376);
and I_6835 (I121931,I121914,I75373);
or I_6836 (I121948,I121931,I75370);
DFFARX1 I_6837  ( .D(I121948), .CLK(I5694_clk), .RSTB(I121716_rst), .Q(I121965) );
nor I_6838 (I121982,I121965,I121818);
DFFARX1 I_6839  ( .D(I121965), .CLK(I5694_clk), .RSTB(I121716_rst), .Q(I121999) );
not I_6840 (I121687,I121999);
nand I_6841 (I122030,I121733,I75385);
and I_6842 (I122047,I122030,I121982);
DFFARX1 I_6843  ( .D(I122030), .CLK(I5694_clk), .RSTB(I121716_rst), .Q(I121684) );
DFFARX1 I_6844  ( .D(I75394), .CLK(I5694_clk), .RSTB(I121716_rst), .Q(I122078) );
nor I_6845 (I122095,I122078,I121801);
nand I_6846 (I121702,I121965,I122095);
nor I_6847 (I122126,I122078,I121866);
not I_6848 (I121699,I122078);
nand I_6849 (I122157,I122078,I121767);
and I_6850 (I122174,I121835,I122157);
DFFARX1 I_6851  ( .D(I122174), .CLK(I5694_clk), .RSTB(I121716_rst), .Q(I121678) );
DFFARX1 I_6852  ( .D(I122078), .CLK(I5694_clk), .RSTB(I121716_rst), .Q(I121681) );
DFFARX1 I_6853  ( .D(I75382), .CLK(I5694_clk), .RSTB(I121716_rst), .Q(I122219) );
not I_6854 (I122236,I122219);
nand I_6855 (I122253,I122236,I121801);
and I_6856 (I122270,I122030,I122253);
DFFARX1 I_6857  ( .D(I122270), .CLK(I5694_clk), .RSTB(I121716_rst), .Q(I121708) );
or I_6858 (I122301,I122236,I122047);
DFFARX1 I_6859  ( .D(I122301), .CLK(I5694_clk), .RSTB(I121716_rst), .Q(I121693) );
nand I_6860 (I121696,I122236,I122126);
not I_6861 (I122379_rst,I5701);
not I_6862 (I122396,I105126);
nor I_6863 (I122413,I105123,I105147);
nand I_6864 (I122430,I122413,I105144);
nor I_6865 (I122447,I122396,I105123);
nand I_6866 (I122464,I122447,I105150);
not I_6867 (I122481,I122464);
not I_6868 (I122498,I105123);
nor I_6869 (I122368,I122464,I122498);
not I_6870 (I122529,I122498);
nand I_6871 (I122353,I122464,I122529);
not I_6872 (I122560,I105141);
nor I_6873 (I122577,I122560,I105132);
and I_6874 (I122594,I122577,I105129);
or I_6875 (I122611,I122594,I105138);
DFFARX1 I_6876  ( .D(I122611), .CLK(I5694_clk), .RSTB(I122379_rst), .Q(I122628) );
nor I_6877 (I122645,I122628,I122481);
DFFARX1 I_6878  ( .D(I122628), .CLK(I5694_clk), .RSTB(I122379_rst), .Q(I122662) );
not I_6879 (I122350,I122662);
nand I_6880 (I122693,I122396,I105141);
and I_6881 (I122710,I122693,I122645);
DFFARX1 I_6882  ( .D(I122693), .CLK(I5694_clk), .RSTB(I122379_rst), .Q(I122347) );
DFFARX1 I_6883  ( .D(I105120), .CLK(I5694_clk), .RSTB(I122379_rst), .Q(I122741) );
nor I_6884 (I122758,I122741,I122464);
nand I_6885 (I122365,I122628,I122758);
nor I_6886 (I122789,I122741,I122529);
not I_6887 (I122362,I122741);
nand I_6888 (I122820,I122741,I122430);
and I_6889 (I122837,I122498,I122820);
DFFARX1 I_6890  ( .D(I122837), .CLK(I5694_clk), .RSTB(I122379_rst), .Q(I122341) );
DFFARX1 I_6891  ( .D(I122741), .CLK(I5694_clk), .RSTB(I122379_rst), .Q(I122344) );
DFFARX1 I_6892  ( .D(I105135), .CLK(I5694_clk), .RSTB(I122379_rst), .Q(I122882) );
not I_6893 (I122899,I122882);
nand I_6894 (I122916,I122899,I122464);
and I_6895 (I122933,I122693,I122916);
DFFARX1 I_6896  ( .D(I122933), .CLK(I5694_clk), .RSTB(I122379_rst), .Q(I122371) );
or I_6897 (I122964,I122899,I122710);
DFFARX1 I_6898  ( .D(I122964), .CLK(I5694_clk), .RSTB(I122379_rst), .Q(I122356) );
nand I_6899 (I122359,I122899,I122789);
not I_6900 (I123042_rst,I5701);
not I_6901 (I123059,I82516);
nor I_6902 (I123076,I82534,I82525);
nand I_6903 (I123093,I123076,I82531);
nor I_6904 (I123110,I123059,I82534);
nand I_6905 (I123127,I123110,I82537);
not I_6906 (I123144,I123127);
not I_6907 (I123161,I82534);
nor I_6908 (I123031,I123127,I123161);
not I_6909 (I123192,I123161);
nand I_6910 (I123016,I123127,I123192);
not I_6911 (I123223,I82513);
nor I_6912 (I123240,I123223,I82528);
and I_6913 (I123257,I123240,I82510);
or I_6914 (I123274,I123257,I82519);
DFFARX1 I_6915  ( .D(I123274), .CLK(I5694_clk), .RSTB(I123042_rst), .Q(I123291) );
nor I_6916 (I123308,I123291,I123144);
DFFARX1 I_6917  ( .D(I123291), .CLK(I5694_clk), .RSTB(I123042_rst), .Q(I123325) );
not I_6918 (I123013,I123325);
nand I_6919 (I123356,I123059,I82513);
and I_6920 (I123373,I123356,I123308);
DFFARX1 I_6921  ( .D(I123356), .CLK(I5694_clk), .RSTB(I123042_rst), .Q(I123010) );
DFFARX1 I_6922  ( .D(I82522), .CLK(I5694_clk), .RSTB(I123042_rst), .Q(I123404) );
nor I_6923 (I123421,I123404,I123127);
nand I_6924 (I123028,I123291,I123421);
nor I_6925 (I123452,I123404,I123192);
not I_6926 (I123025,I123404);
nand I_6927 (I123483,I123404,I123093);
and I_6928 (I123500,I123161,I123483);
DFFARX1 I_6929  ( .D(I123500), .CLK(I5694_clk), .RSTB(I123042_rst), .Q(I123004) );
DFFARX1 I_6930  ( .D(I123404), .CLK(I5694_clk), .RSTB(I123042_rst), .Q(I123007) );
DFFARX1 I_6931  ( .D(I82540), .CLK(I5694_clk), .RSTB(I123042_rst), .Q(I123545) );
not I_6932 (I123562,I123545);
nand I_6933 (I123579,I123562,I123127);
and I_6934 (I123596,I123356,I123579);
DFFARX1 I_6935  ( .D(I123596), .CLK(I5694_clk), .RSTB(I123042_rst), .Q(I123034) );
or I_6936 (I123627,I123562,I123373);
DFFARX1 I_6937  ( .D(I123627), .CLK(I5694_clk), .RSTB(I123042_rst), .Q(I123019) );
nand I_6938 (I123022,I123562,I123452);
not I_6939 (I123705_rst,I5701);
not I_6940 (I123722,I109033);
nor I_6941 (I123739,I109039,I109045);
nand I_6942 (I123756,I123739,I109048);
nor I_6943 (I123773,I123722,I109039);
nand I_6944 (I123790,I123773,I109030);
not I_6945 (I123807,I123790);
not I_6946 (I123824,I109039);
nor I_6947 (I123694,I123790,I123824);
not I_6948 (I123855,I123824);
nand I_6949 (I123679,I123790,I123855);
not I_6950 (I123886,I109042);
nor I_6951 (I123903,I123886,I109036);
and I_6952 (I123920,I123903,I109051);
or I_6953 (I123937,I123920,I109057);
DFFARX1 I_6954  ( .D(I123937), .CLK(I5694_clk), .RSTB(I123705_rst), .Q(I123954) );
nor I_6955 (I123971,I123954,I123807);
DFFARX1 I_6956  ( .D(I123954), .CLK(I5694_clk), .RSTB(I123705_rst), .Q(I123988) );
not I_6957 (I123676,I123988);
nand I_6958 (I124019,I123722,I109042);
and I_6959 (I124036,I124019,I123971);
DFFARX1 I_6960  ( .D(I124019), .CLK(I5694_clk), .RSTB(I123705_rst), .Q(I123673) );
DFFARX1 I_6961  ( .D(I109054), .CLK(I5694_clk), .RSTB(I123705_rst), .Q(I124067) );
nor I_6962 (I124084,I124067,I123790);
nand I_6963 (I123691,I123954,I124084);
nor I_6964 (I124115,I124067,I123855);
not I_6965 (I123688,I124067);
nand I_6966 (I124146,I124067,I123756);
and I_6967 (I124163,I123824,I124146);
DFFARX1 I_6968  ( .D(I124163), .CLK(I5694_clk), .RSTB(I123705_rst), .Q(I123667) );
DFFARX1 I_6969  ( .D(I124067), .CLK(I5694_clk), .RSTB(I123705_rst), .Q(I123670) );
DFFARX1 I_6970  ( .D(I109060), .CLK(I5694_clk), .RSTB(I123705_rst), .Q(I124208) );
not I_6971 (I124225,I124208);
nand I_6972 (I124242,I124225,I123790);
and I_6973 (I124259,I124019,I124242);
DFFARX1 I_6974  ( .D(I124259), .CLK(I5694_clk), .RSTB(I123705_rst), .Q(I123697) );
or I_6975 (I124290,I124225,I124036);
DFFARX1 I_6976  ( .D(I124290), .CLK(I5694_clk), .RSTB(I123705_rst), .Q(I123682) );
nand I_6977 (I123685,I124225,I124115);
not I_6978 (I124368_rst,I5701);
not I_6979 (I124385,I58909);
nor I_6980 (I124402,I58906,I58924);
nand I_6981 (I124419,I124402,I58927);
nor I_6982 (I124436,I124385,I58906);
nand I_6983 (I124453,I124436,I58912);
not I_6984 (I124470,I124453);
not I_6985 (I124487,I58906);
nor I_6986 (I124357,I124453,I124487);
not I_6987 (I124518,I124487);
nand I_6988 (I124342,I124453,I124518);
not I_6989 (I124549,I58921);
nor I_6990 (I124566,I124549,I58903);
and I_6991 (I124583,I124566,I58897);
or I_6992 (I124600,I124583,I58915);
DFFARX1 I_6993  ( .D(I124600), .CLK(I5694_clk), .RSTB(I124368_rst), .Q(I124617) );
nor I_6994 (I124634,I124617,I124470);
DFFARX1 I_6995  ( .D(I124617), .CLK(I5694_clk), .RSTB(I124368_rst), .Q(I124651) );
not I_6996 (I124339,I124651);
nand I_6997 (I124682,I124385,I58921);
and I_6998 (I124699,I124682,I124634);
DFFARX1 I_6999  ( .D(I124682), .CLK(I5694_clk), .RSTB(I124368_rst), .Q(I124336) );
DFFARX1 I_7000  ( .D(I58900), .CLK(I5694_clk), .RSTB(I124368_rst), .Q(I124730) );
nor I_7001 (I124747,I124730,I124453);
nand I_7002 (I124354,I124617,I124747);
nor I_7003 (I124778,I124730,I124518);
not I_7004 (I124351,I124730);
nand I_7005 (I124809,I124730,I124419);
and I_7006 (I124826,I124487,I124809);
DFFARX1 I_7007  ( .D(I124826), .CLK(I5694_clk), .RSTB(I124368_rst), .Q(I124330) );
DFFARX1 I_7008  ( .D(I124730), .CLK(I5694_clk), .RSTB(I124368_rst), .Q(I124333) );
DFFARX1 I_7009  ( .D(I58918), .CLK(I5694_clk), .RSTB(I124368_rst), .Q(I124871) );
not I_7010 (I124888,I124871);
nand I_7011 (I124905,I124888,I124453);
and I_7012 (I124922,I124682,I124905);
DFFARX1 I_7013  ( .D(I124922), .CLK(I5694_clk), .RSTB(I124368_rst), .Q(I124360) );
or I_7014 (I124953,I124888,I124699);
DFFARX1 I_7015  ( .D(I124953), .CLK(I5694_clk), .RSTB(I124368_rst), .Q(I124345) );
nand I_7016 (I124348,I124888,I124778);
not I_7017 (I125031_rst,I5701);
not I_7018 (I125048,I96434);
nor I_7019 (I125065,I96440,I96443);
nand I_7020 (I125082,I125065,I96419);
nor I_7021 (I125099,I125048,I96440);
nand I_7022 (I125116,I125099,I96428);
not I_7023 (I125133,I125116);
not I_7024 (I125150,I96440);
nor I_7025 (I125020,I125116,I125150);
not I_7026 (I125181,I125150);
nand I_7027 (I125005,I125116,I125181);
not I_7028 (I125212,I96422);
nor I_7029 (I125229,I125212,I96446);
and I_7030 (I125246,I125229,I96416);
or I_7031 (I125263,I125246,I96425);
DFFARX1 I_7032  ( .D(I125263), .CLK(I5694_clk), .RSTB(I125031_rst), .Q(I125280) );
nor I_7033 (I125297,I125280,I125133);
DFFARX1 I_7034  ( .D(I125280), .CLK(I5694_clk), .RSTB(I125031_rst), .Q(I125314) );
not I_7035 (I125002,I125314);
nand I_7036 (I125345,I125048,I96422);
and I_7037 (I125362,I125345,I125297);
DFFARX1 I_7038  ( .D(I125345), .CLK(I5694_clk), .RSTB(I125031_rst), .Q(I124999) );
DFFARX1 I_7039  ( .D(I96431), .CLK(I5694_clk), .RSTB(I125031_rst), .Q(I125393) );
nor I_7040 (I125410,I125393,I125116);
nand I_7041 (I125017,I125280,I125410);
nor I_7042 (I125441,I125393,I125181);
not I_7043 (I125014,I125393);
nand I_7044 (I125472,I125393,I125082);
and I_7045 (I125489,I125150,I125472);
DFFARX1 I_7046  ( .D(I125489), .CLK(I5694_clk), .RSTB(I125031_rst), .Q(I124993) );
DFFARX1 I_7047  ( .D(I125393), .CLK(I5694_clk), .RSTB(I125031_rst), .Q(I124996) );
DFFARX1 I_7048  ( .D(I96437), .CLK(I5694_clk), .RSTB(I125031_rst), .Q(I125534) );
not I_7049 (I125551,I125534);
nand I_7050 (I125568,I125551,I125116);
and I_7051 (I125585,I125345,I125568);
DFFARX1 I_7052  ( .D(I125585), .CLK(I5694_clk), .RSTB(I125031_rst), .Q(I125023) );
or I_7053 (I125616,I125551,I125362);
DFFARX1 I_7054  ( .D(I125616), .CLK(I5694_clk), .RSTB(I125031_rst), .Q(I125008) );
nand I_7055 (I125011,I125551,I125441);
not I_7056 (I125694_rst,I5701);
not I_7057 (I125711,I103188);
nor I_7058 (I125728,I103185,I103209);
nand I_7059 (I125745,I125728,I103206);
nor I_7060 (I125762,I125711,I103185);
nand I_7061 (I125779,I125762,I103212);
not I_7062 (I125796,I125779);
not I_7063 (I125813,I103185);
nor I_7064 (I125683,I125779,I125813);
not I_7065 (I125844,I125813);
nand I_7066 (I125668,I125779,I125844);
not I_7067 (I125875,I103203);
nor I_7068 (I125892,I125875,I103194);
and I_7069 (I125909,I125892,I103191);
or I_7070 (I125926,I125909,I103200);
DFFARX1 I_7071  ( .D(I125926), .CLK(I5694_clk), .RSTB(I125694_rst), .Q(I125943) );
nor I_7072 (I125960,I125943,I125796);
DFFARX1 I_7073  ( .D(I125943), .CLK(I5694_clk), .RSTB(I125694_rst), .Q(I125977) );
not I_7074 (I125665,I125977);
nand I_7075 (I126008,I125711,I103203);
and I_7076 (I126025,I126008,I125960);
DFFARX1 I_7077  ( .D(I126008), .CLK(I5694_clk), .RSTB(I125694_rst), .Q(I125662) );
DFFARX1 I_7078  ( .D(I103182), .CLK(I5694_clk), .RSTB(I125694_rst), .Q(I126056) );
nor I_7079 (I126073,I126056,I125779);
nand I_7080 (I125680,I125943,I126073);
nor I_7081 (I126104,I126056,I125844);
not I_7082 (I125677,I126056);
nand I_7083 (I126135,I126056,I125745);
and I_7084 (I126152,I125813,I126135);
DFFARX1 I_7085  ( .D(I126152), .CLK(I5694_clk), .RSTB(I125694_rst), .Q(I125656) );
DFFARX1 I_7086  ( .D(I126056), .CLK(I5694_clk), .RSTB(I125694_rst), .Q(I125659) );
DFFARX1 I_7087  ( .D(I103197), .CLK(I5694_clk), .RSTB(I125694_rst), .Q(I126197) );
not I_7088 (I126214,I126197);
nand I_7089 (I126231,I126214,I125779);
and I_7090 (I126248,I126008,I126231);
DFFARX1 I_7091  ( .D(I126248), .CLK(I5694_clk), .RSTB(I125694_rst), .Q(I125686) );
or I_7092 (I126279,I126214,I126025);
DFFARX1 I_7093  ( .D(I126279), .CLK(I5694_clk), .RSTB(I125694_rst), .Q(I125671) );
nand I_7094 (I125674,I126214,I126104);
not I_7095 (I126357_rst,I5701);
not I_7096 (I126374,I113689);
nor I_7097 (I126391,I113683,I113674);
nand I_7098 (I126408,I126391,I113686);
nor I_7099 (I126425,I126374,I113683);
nand I_7100 (I126442,I126425,I113701);
not I_7101 (I126459,I126442);
not I_7102 (I126476,I113683);
nor I_7103 (I126346,I126442,I126476);
not I_7104 (I126507,I126476);
nand I_7105 (I126331,I126442,I126507);
not I_7106 (I126538,I113677);
nor I_7107 (I126555,I126538,I113671);
and I_7108 (I126572,I126555,I113698);
or I_7109 (I126589,I126572,I113695);
DFFARX1 I_7110  ( .D(I126589), .CLK(I5694_clk), .RSTB(I126357_rst), .Q(I126606) );
nor I_7111 (I126623,I126606,I126459);
DFFARX1 I_7112  ( .D(I126606), .CLK(I5694_clk), .RSTB(I126357_rst), .Q(I126640) );
not I_7113 (I126328,I126640);
nand I_7114 (I126671,I126374,I113677);
and I_7115 (I126688,I126671,I126623);
DFFARX1 I_7116  ( .D(I126671), .CLK(I5694_clk), .RSTB(I126357_rst), .Q(I126325) );
DFFARX1 I_7117  ( .D(I113692), .CLK(I5694_clk), .RSTB(I126357_rst), .Q(I126719) );
nor I_7118 (I126736,I126719,I126442);
nand I_7119 (I126343,I126606,I126736);
nor I_7120 (I126767,I126719,I126507);
not I_7121 (I126340,I126719);
nand I_7122 (I126798,I126719,I126408);
and I_7123 (I126815,I126476,I126798);
DFFARX1 I_7124  ( .D(I126815), .CLK(I5694_clk), .RSTB(I126357_rst), .Q(I126319) );
DFFARX1 I_7125  ( .D(I126719), .CLK(I5694_clk), .RSTB(I126357_rst), .Q(I126322) );
DFFARX1 I_7126  ( .D(I113680), .CLK(I5694_clk), .RSTB(I126357_rst), .Q(I126860) );
not I_7127 (I126877,I126860);
nand I_7128 (I126894,I126877,I126442);
and I_7129 (I126911,I126671,I126894);
DFFARX1 I_7130  ( .D(I126911), .CLK(I5694_clk), .RSTB(I126357_rst), .Q(I126349) );
or I_7131 (I126942,I126877,I126688);
DFFARX1 I_7132  ( .D(I126942), .CLK(I5694_clk), .RSTB(I126357_rst), .Q(I126334) );
nand I_7133 (I126337,I126877,I126767);
not I_7134 (I127020_rst,I5701);
not I_7135 (I127037,I110359);
nor I_7136 (I127054,I110365,I110371);
nand I_7137 (I127071,I127054,I110374);
nor I_7138 (I127088,I127037,I110365);
nand I_7139 (I127105,I127088,I110356);
not I_7140 (I127122,I127105);
not I_7141 (I127139,I110365);
nor I_7142 (I127009,I127105,I127139);
not I_7143 (I127170,I127139);
nand I_7144 (I126994,I127105,I127170);
not I_7145 (I127201,I110368);
nor I_7146 (I127218,I127201,I110362);
and I_7147 (I127235,I127218,I110377);
or I_7148 (I127252,I127235,I110383);
DFFARX1 I_7149  ( .D(I127252), .CLK(I5694_clk), .RSTB(I127020_rst), .Q(I127269) );
nor I_7150 (I127286,I127269,I127122);
DFFARX1 I_7151  ( .D(I127269), .CLK(I5694_clk), .RSTB(I127020_rst), .Q(I127303) );
not I_7152 (I126991,I127303);
nand I_7153 (I127334,I127037,I110368);
and I_7154 (I127351,I127334,I127286);
DFFARX1 I_7155  ( .D(I127334), .CLK(I5694_clk), .RSTB(I127020_rst), .Q(I126988) );
DFFARX1 I_7156  ( .D(I110380), .CLK(I5694_clk), .RSTB(I127020_rst), .Q(I127382) );
nor I_7157 (I127399,I127382,I127105);
nand I_7158 (I127006,I127269,I127399);
nor I_7159 (I127430,I127382,I127170);
not I_7160 (I127003,I127382);
nand I_7161 (I127461,I127382,I127071);
and I_7162 (I127478,I127139,I127461);
DFFARX1 I_7163  ( .D(I127478), .CLK(I5694_clk), .RSTB(I127020_rst), .Q(I126982) );
DFFARX1 I_7164  ( .D(I127382), .CLK(I5694_clk), .RSTB(I127020_rst), .Q(I126985) );
DFFARX1 I_7165  ( .D(I110386), .CLK(I5694_clk), .RSTB(I127020_rst), .Q(I127523) );
not I_7166 (I127540,I127523);
nand I_7167 (I127557,I127540,I127105);
and I_7168 (I127574,I127334,I127557);
DFFARX1 I_7169  ( .D(I127574), .CLK(I5694_clk), .RSTB(I127020_rst), .Q(I127012) );
or I_7170 (I127605,I127540,I127351);
DFFARX1 I_7171  ( .D(I127605), .CLK(I5694_clk), .RSTB(I127020_rst), .Q(I126997) );
nand I_7172 (I127000,I127540,I127430);
not I_7173 (I127683_rst,I5701);
not I_7174 (I127700,I116652);
nor I_7175 (I127717,I116658,I116655);
nand I_7176 (I127734,I127717,I116649);
nor I_7177 (I127751,I127700,I116658);
nand I_7178 (I127768,I127751,I116673);
DFFARX1 I_7179  ( .D(I127768), .CLK(I5694_clk), .RSTB(I127683_rst), .Q(I127785) );
not I_7180 (I127654,I127785);
not I_7181 (I127816,I116658);
not I_7182 (I127833,I127816);
not I_7183 (I127850,I116670);
nor I_7184 (I127867,I127850,I116661);
and I_7185 (I127884,I127867,I116646);
or I_7186 (I127901,I127884,I116667);
DFFARX1 I_7187  ( .D(I127901), .CLK(I5694_clk), .RSTB(I127683_rst), .Q(I127918) );
DFFARX1 I_7188  ( .D(I127918), .CLK(I5694_clk), .RSTB(I127683_rst), .Q(I127651) );
DFFARX1 I_7189  ( .D(I127918), .CLK(I5694_clk), .RSTB(I127683_rst), .Q(I127949) );
DFFARX1 I_7190  ( .D(I127918), .CLK(I5694_clk), .RSTB(I127683_rst), .Q(I127645) );
nand I_7191 (I127980,I127700,I116670);
nand I_7192 (I127997,I127980,I127734);
and I_7193 (I128014,I127816,I127997);
DFFARX1 I_7194  ( .D(I128014), .CLK(I5694_clk), .RSTB(I127683_rst), .Q(I127675) );
and I_7195 (I127648,I127980,I127949);
DFFARX1 I_7196  ( .D(I116664), .CLK(I5694_clk), .RSTB(I127683_rst), .Q(I128059) );
nor I_7197 (I127672,I128059,I127980);
nor I_7198 (I128090,I128059,I127734);
nand I_7199 (I127669,I127768,I128090);
not I_7200 (I127666,I128059);
DFFARX1 I_7201  ( .D(I116676), .CLK(I5694_clk), .RSTB(I127683_rst), .Q(I128135) );
not I_7202 (I128152,I128135);
nor I_7203 (I128169,I128152,I127833);
and I_7204 (I128186,I128059,I128169);
or I_7205 (I128203,I127980,I128186);
DFFARX1 I_7206  ( .D(I128203), .CLK(I5694_clk), .RSTB(I127683_rst), .Q(I127660) );
not I_7207 (I128234,I128152);
nor I_7208 (I128251,I128059,I128234);
nand I_7209 (I127663,I128152,I128251);
nand I_7210 (I127657,I127816,I128234);
not I_7211 (I128329_rst,I5701);
not I_7212 (I128346,I98108);
nor I_7213 (I128363,I98123,I98117);
nand I_7214 (I128380,I128363,I98126);
nor I_7215 (I128397,I128346,I98123);
nand I_7216 (I128414,I128397,I98102);
DFFARX1 I_7217  ( .D(I128414), .CLK(I5694_clk), .RSTB(I128329_rst), .Q(I128431) );
not I_7218 (I128300,I128431);
not I_7219 (I128462,I98123);
not I_7220 (I128479,I128462);
not I_7221 (I128496,I98099);
nor I_7222 (I128513,I128496,I98114);
and I_7223 (I128530,I128513,I98120);
or I_7224 (I128547,I128530,I98129);
DFFARX1 I_7225  ( .D(I128547), .CLK(I5694_clk), .RSTB(I128329_rst), .Q(I128564) );
DFFARX1 I_7226  ( .D(I128564), .CLK(I5694_clk), .RSTB(I128329_rst), .Q(I128297) );
DFFARX1 I_7227  ( .D(I128564), .CLK(I5694_clk), .RSTB(I128329_rst), .Q(I128595) );
DFFARX1 I_7228  ( .D(I128564), .CLK(I5694_clk), .RSTB(I128329_rst), .Q(I128291) );
nand I_7229 (I128626,I128346,I98099);
nand I_7230 (I128643,I128626,I128380);
and I_7231 (I128660,I128462,I128643);
DFFARX1 I_7232  ( .D(I128660), .CLK(I5694_clk), .RSTB(I128329_rst), .Q(I128321) );
and I_7233 (I128294,I128626,I128595);
DFFARX1 I_7234  ( .D(I98111), .CLK(I5694_clk), .RSTB(I128329_rst), .Q(I128705) );
nor I_7235 (I128318,I128705,I128626);
nor I_7236 (I128736,I128705,I128380);
nand I_7237 (I128315,I128414,I128736);
not I_7238 (I128312,I128705);
DFFARX1 I_7239  ( .D(I98105), .CLK(I5694_clk), .RSTB(I128329_rst), .Q(I128781) );
not I_7240 (I128798,I128781);
nor I_7241 (I128815,I128798,I128479);
and I_7242 (I128832,I128705,I128815);
or I_7243 (I128849,I128626,I128832);
DFFARX1 I_7244  ( .D(I128849), .CLK(I5694_clk), .RSTB(I128329_rst), .Q(I128306) );
not I_7245 (I128880,I128798);
nor I_7246 (I128897,I128705,I128880);
nand I_7247 (I128309,I128798,I128897);
nand I_7248 (I128303,I128462,I128880);
not I_7249 (I128975_rst,I5701);
not I_7250 (I128992,I81933);
nor I_7251 (I129009,I81921,I81930);
nand I_7252 (I129026,I129009,I81945);
nor I_7253 (I129043,I128992,I81921);
nand I_7254 (I129060,I129043,I81927);
DFFARX1 I_7255  ( .D(I129060), .CLK(I5694_clk), .RSTB(I128975_rst), .Q(I129077) );
not I_7256 (I128946,I129077);
not I_7257 (I129108,I81921);
not I_7258 (I129125,I129108);
not I_7259 (I129142,I81915);
nor I_7260 (I129159,I129142,I81936);
and I_7261 (I129176,I129159,I81918);
or I_7262 (I129193,I129176,I81924);
DFFARX1 I_7263  ( .D(I129193), .CLK(I5694_clk), .RSTB(I128975_rst), .Q(I129210) );
DFFARX1 I_7264  ( .D(I129210), .CLK(I5694_clk), .RSTB(I128975_rst), .Q(I128943) );
DFFARX1 I_7265  ( .D(I129210), .CLK(I5694_clk), .RSTB(I128975_rst), .Q(I129241) );
DFFARX1 I_7266  ( .D(I129210), .CLK(I5694_clk), .RSTB(I128975_rst), .Q(I128937) );
nand I_7267 (I129272,I128992,I81915);
nand I_7268 (I129289,I129272,I129026);
and I_7269 (I129306,I129108,I129289);
DFFARX1 I_7270  ( .D(I129306), .CLK(I5694_clk), .RSTB(I128975_rst), .Q(I128967) );
and I_7271 (I128940,I129272,I129241);
DFFARX1 I_7272  ( .D(I81942), .CLK(I5694_clk), .RSTB(I128975_rst), .Q(I129351) );
nor I_7273 (I128964,I129351,I129272);
nor I_7274 (I129382,I129351,I129026);
nand I_7275 (I128961,I129060,I129382);
not I_7276 (I128958,I129351);
DFFARX1 I_7277  ( .D(I81939), .CLK(I5694_clk), .RSTB(I128975_rst), .Q(I129427) );
not I_7278 (I129444,I129427);
nor I_7279 (I129461,I129444,I129125);
and I_7280 (I129478,I129351,I129461);
or I_7281 (I129495,I129272,I129478);
DFFARX1 I_7282  ( .D(I129495), .CLK(I5694_clk), .RSTB(I128975_rst), .Q(I128952) );
not I_7283 (I129526,I129444);
nor I_7284 (I129543,I129351,I129526);
nand I_7285 (I128955,I129444,I129543);
nand I_7286 (I128949,I129108,I129526);
not I_7287 (I129621_rst,I5701);
not I_7288 (I129638,I70642);
nor I_7289 (I129655,I70645,I70627);
nand I_7290 (I129672,I129655,I70654);
nor I_7291 (I129689,I129638,I70645);
nand I_7292 (I129706,I129689,I70633);
DFFARX1 I_7293  ( .D(I129706), .CLK(I5694_clk), .RSTB(I129621_rst), .Q(I129723) );
not I_7294 (I129592,I129723);
not I_7295 (I129754,I70645);
not I_7296 (I129771,I129754);
not I_7297 (I129788,I70639);
nor I_7298 (I129805,I129788,I70651);
and I_7299 (I129822,I129805,I70657);
or I_7300 (I129839,I129822,I70636);
DFFARX1 I_7301  ( .D(I129839), .CLK(I5694_clk), .RSTB(I129621_rst), .Q(I129856) );
DFFARX1 I_7302  ( .D(I129856), .CLK(I5694_clk), .RSTB(I129621_rst), .Q(I129589) );
DFFARX1 I_7303  ( .D(I129856), .CLK(I5694_clk), .RSTB(I129621_rst), .Q(I129887) );
DFFARX1 I_7304  ( .D(I129856), .CLK(I5694_clk), .RSTB(I129621_rst), .Q(I129583) );
nand I_7305 (I129918,I129638,I70639);
nand I_7306 (I129935,I129918,I129672);
and I_7307 (I129952,I129754,I129935);
DFFARX1 I_7308  ( .D(I129952), .CLK(I5694_clk), .RSTB(I129621_rst), .Q(I129613) );
and I_7309 (I129586,I129918,I129887);
DFFARX1 I_7310  ( .D(I70648), .CLK(I5694_clk), .RSTB(I129621_rst), .Q(I129997) );
nor I_7311 (I129610,I129997,I129918);
nor I_7312 (I130028,I129997,I129672);
nand I_7313 (I129607,I129706,I130028);
not I_7314 (I129604,I129997);
DFFARX1 I_7315  ( .D(I70630), .CLK(I5694_clk), .RSTB(I129621_rst), .Q(I130073) );
not I_7316 (I130090,I130073);
nor I_7317 (I130107,I130090,I129771);
and I_7318 (I130124,I129997,I130107);
or I_7319 (I130141,I129918,I130124);
DFFARX1 I_7320  ( .D(I130141), .CLK(I5694_clk), .RSTB(I129621_rst), .Q(I129598) );
not I_7321 (I130172,I130090);
nor I_7322 (I130189,I129997,I130172);
nand I_7323 (I129601,I130090,I130189);
nand I_7324 (I129595,I129754,I130172);
not I_7325 (I130267_rst,I5701);
not I_7326 (I130284,I83789);
nor I_7327 (I130301,I83786,I83771);
nand I_7328 (I130318,I130301,I83780);
nor I_7329 (I130335,I130284,I83786);
nand I_7330 (I130352,I130335,I83795);
DFFARX1 I_7331  ( .D(I130352), .CLK(I5694_clk), .RSTB(I130267_rst), .Q(I130369) );
not I_7332 (I130238,I130369);
not I_7333 (I130400,I83786);
not I_7334 (I130417,I130400);
not I_7335 (I130434,I83768);
nor I_7336 (I130451,I130434,I83774);
and I_7337 (I130468,I130451,I83798);
or I_7338 (I130485,I130468,I83792);
DFFARX1 I_7339  ( .D(I130485), .CLK(I5694_clk), .RSTB(I130267_rst), .Q(I130502) );
DFFARX1 I_7340  ( .D(I130502), .CLK(I5694_clk), .RSTB(I130267_rst), .Q(I130235) );
DFFARX1 I_7341  ( .D(I130502), .CLK(I5694_clk), .RSTB(I130267_rst), .Q(I130533) );
DFFARX1 I_7342  ( .D(I130502), .CLK(I5694_clk), .RSTB(I130267_rst), .Q(I130229) );
nand I_7343 (I130564,I130284,I83768);
nand I_7344 (I130581,I130564,I130318);
and I_7345 (I130598,I130400,I130581);
DFFARX1 I_7346  ( .D(I130598), .CLK(I5694_clk), .RSTB(I130267_rst), .Q(I130259) );
and I_7347 (I130232,I130564,I130533);
DFFARX1 I_7348  ( .D(I83777), .CLK(I5694_clk), .RSTB(I130267_rst), .Q(I130643) );
nor I_7349 (I130256,I130643,I130564);
nor I_7350 (I130674,I130643,I130318);
nand I_7351 (I130253,I130352,I130674);
not I_7352 (I130250,I130643);
DFFARX1 I_7353  ( .D(I83783), .CLK(I5694_clk), .RSTB(I130267_rst), .Q(I130719) );
not I_7354 (I130736,I130719);
nor I_7355 (I130753,I130736,I130417);
and I_7356 (I130770,I130643,I130753);
or I_7357 (I130787,I130564,I130770);
DFFARX1 I_7358  ( .D(I130787), .CLK(I5694_clk), .RSTB(I130267_rst), .Q(I130244) );
not I_7359 (I130818,I130736);
nor I_7360 (I130835,I130643,I130818);
nand I_7361 (I130247,I130736,I130835);
nand I_7362 (I130241,I130400,I130818);
not I_7363 (I130913_rst,I5701);
not I_7364 (I130930,I68908);
nor I_7365 (I130947,I68911,I68893);
nand I_7366 (I130964,I130947,I68920);
nor I_7367 (I130981,I130930,I68911);
nand I_7368 (I130998,I130981,I68899);
DFFARX1 I_7369  ( .D(I130998), .CLK(I5694_clk), .RSTB(I130913_rst), .Q(I131015) );
not I_7370 (I130884,I131015);
not I_7371 (I131046,I68911);
not I_7372 (I131063,I131046);
not I_7373 (I131080,I68905);
nor I_7374 (I131097,I131080,I68917);
and I_7375 (I131114,I131097,I68923);
or I_7376 (I131131,I131114,I68902);
DFFARX1 I_7377  ( .D(I131131), .CLK(I5694_clk), .RSTB(I130913_rst), .Q(I131148) );
DFFARX1 I_7378  ( .D(I131148), .CLK(I5694_clk), .RSTB(I130913_rst), .Q(I130881) );
DFFARX1 I_7379  ( .D(I131148), .CLK(I5694_clk), .RSTB(I130913_rst), .Q(I131179) );
DFFARX1 I_7380  ( .D(I131148), .CLK(I5694_clk), .RSTB(I130913_rst), .Q(I130875) );
nand I_7381 (I131210,I130930,I68905);
nand I_7382 (I131227,I131210,I130964);
and I_7383 (I131244,I131046,I131227);
DFFARX1 I_7384  ( .D(I131244), .CLK(I5694_clk), .RSTB(I130913_rst), .Q(I130905) );
and I_7385 (I130878,I131210,I131179);
DFFARX1 I_7386  ( .D(I68914), .CLK(I5694_clk), .RSTB(I130913_rst), .Q(I131289) );
nor I_7387 (I130902,I131289,I131210);
nor I_7388 (I131320,I131289,I130964);
nand I_7389 (I130899,I130998,I131320);
not I_7390 (I130896,I131289);
DFFARX1 I_7391  ( .D(I68896), .CLK(I5694_clk), .RSTB(I130913_rst), .Q(I131365) );
not I_7392 (I131382,I131365);
nor I_7393 (I131399,I131382,I131063);
and I_7394 (I131416,I131289,I131399);
or I_7395 (I131433,I131210,I131416);
DFFARX1 I_7396  ( .D(I131433), .CLK(I5694_clk), .RSTB(I130913_rst), .Q(I130890) );
not I_7397 (I131464,I131382);
nor I_7398 (I131481,I131289,I131464);
nand I_7399 (I130893,I131382,I131481);
nand I_7400 (I130887,I131046,I131464);
not I_7401 (I131559_rst,I5701);
not I_7402 (I131576,I108370);
nor I_7403 (I131593,I108391,I108373);
nand I_7404 (I131610,I131593,I108397);
nor I_7405 (I131627,I131576,I108391);
nand I_7406 (I131644,I131627,I108394);
DFFARX1 I_7407  ( .D(I131644), .CLK(I5694_clk), .RSTB(I131559_rst), .Q(I131661) );
not I_7408 (I131530,I131661);
not I_7409 (I131692,I108391);
not I_7410 (I131709,I131692);
not I_7411 (I131726,I108388);
nor I_7412 (I131743,I131726,I108367);
and I_7413 (I131760,I131743,I108379);
or I_7414 (I131777,I131760,I108376);
DFFARX1 I_7415  ( .D(I131777), .CLK(I5694_clk), .RSTB(I131559_rst), .Q(I131794) );
DFFARX1 I_7416  ( .D(I131794), .CLK(I5694_clk), .RSTB(I131559_rst), .Q(I131527) );
DFFARX1 I_7417  ( .D(I131794), .CLK(I5694_clk), .RSTB(I131559_rst), .Q(I131825) );
DFFARX1 I_7418  ( .D(I131794), .CLK(I5694_clk), .RSTB(I131559_rst), .Q(I131521) );
nand I_7419 (I131856,I131576,I108388);
nand I_7420 (I131873,I131856,I131610);
and I_7421 (I131890,I131692,I131873);
DFFARX1 I_7422  ( .D(I131890), .CLK(I5694_clk), .RSTB(I131559_rst), .Q(I131551) );
and I_7423 (I131524,I131856,I131825);
DFFARX1 I_7424  ( .D(I108382), .CLK(I5694_clk), .RSTB(I131559_rst), .Q(I131935) );
nor I_7425 (I131548,I131935,I131856);
nor I_7426 (I131966,I131935,I131610);
nand I_7427 (I131545,I131644,I131966);
not I_7428 (I131542,I131935);
DFFARX1 I_7429  ( .D(I108385), .CLK(I5694_clk), .RSTB(I131559_rst), .Q(I132011) );
not I_7430 (I132028,I132011);
nor I_7431 (I132045,I132028,I131709);
and I_7432 (I132062,I131935,I132045);
or I_7433 (I132079,I131856,I132062);
DFFARX1 I_7434  ( .D(I132079), .CLK(I5694_clk), .RSTB(I131559_rst), .Q(I131536) );
not I_7435 (I132110,I132028);
nor I_7436 (I132127,I131935,I132110);
nand I_7437 (I131539,I132028,I132127);
nand I_7438 (I131533,I131692,I132110);
not I_7439 (I132205_rst,I5701);
not I_7440 (I132222,I126343);
nor I_7441 (I132239,I126322,I126334);
nand I_7442 (I132256,I132239,I126337);
nor I_7443 (I132273,I132222,I126322);
nand I_7444 (I132290,I132273,I126319);
DFFARX1 I_7445  ( .D(I132290), .CLK(I5694_clk), .RSTB(I132205_rst), .Q(I132307) );
not I_7446 (I132176,I132307);
not I_7447 (I132338,I126322);
not I_7448 (I132355,I132338);
not I_7449 (I132372,I126340);
nor I_7450 (I132389,I132372,I126331);
and I_7451 (I132406,I132389,I126325);
or I_7452 (I132423,I132406,I126349);
DFFARX1 I_7453  ( .D(I132423), .CLK(I5694_clk), .RSTB(I132205_rst), .Q(I132440) );
DFFARX1 I_7454  ( .D(I132440), .CLK(I5694_clk), .RSTB(I132205_rst), .Q(I132173) );
DFFARX1 I_7455  ( .D(I132440), .CLK(I5694_clk), .RSTB(I132205_rst), .Q(I132471) );
DFFARX1 I_7456  ( .D(I132440), .CLK(I5694_clk), .RSTB(I132205_rst), .Q(I132167) );
nand I_7457 (I132502,I132222,I126340);
nand I_7458 (I132519,I132502,I132256);
and I_7459 (I132536,I132338,I132519);
DFFARX1 I_7460  ( .D(I132536), .CLK(I5694_clk), .RSTB(I132205_rst), .Q(I132197) );
and I_7461 (I132170,I132502,I132471);
DFFARX1 I_7462  ( .D(I126346), .CLK(I5694_clk), .RSTB(I132205_rst), .Q(I132581) );
nor I_7463 (I132194,I132581,I132502);
nor I_7464 (I132612,I132581,I132256);
nand I_7465 (I132191,I132290,I132612);
not I_7466 (I132188,I132581);
DFFARX1 I_7467  ( .D(I126328), .CLK(I5694_clk), .RSTB(I132205_rst), .Q(I132657) );
not I_7468 (I132674,I132657);
nor I_7469 (I132691,I132674,I132355);
and I_7470 (I132708,I132581,I132691);
or I_7471 (I132725,I132502,I132708);
DFFARX1 I_7472  ( .D(I132725), .CLK(I5694_clk), .RSTB(I132205_rst), .Q(I132182) );
not I_7473 (I132756,I132674);
nor I_7474 (I132773,I132581,I132756);
nand I_7475 (I132185,I132674,I132773);
nand I_7476 (I132179,I132338,I132756);
not I_7477 (I132851_rst,I5701);
not I_7478 (I132868,I107707);
nor I_7479 (I132885,I107728,I107710);
nand I_7480 (I132902,I132885,I107734);
nor I_7481 (I132919,I132868,I107728);
nand I_7482 (I132936,I132919,I107731);
DFFARX1 I_7483  ( .D(I132936), .CLK(I5694_clk), .RSTB(I132851_rst), .Q(I132953) );
not I_7484 (I132822,I132953);
not I_7485 (I132984,I107728);
not I_7486 (I133001,I132984);
not I_7487 (I133018,I107725);
nor I_7488 (I133035,I133018,I107704);
and I_7489 (I133052,I133035,I107716);
or I_7490 (I133069,I133052,I107713);
DFFARX1 I_7491  ( .D(I133069), .CLK(I5694_clk), .RSTB(I132851_rst), .Q(I133086) );
DFFARX1 I_7492  ( .D(I133086), .CLK(I5694_clk), .RSTB(I132851_rst), .Q(I132819) );
DFFARX1 I_7493  ( .D(I133086), .CLK(I5694_clk), .RSTB(I132851_rst), .Q(I133117) );
DFFARX1 I_7494  ( .D(I133086), .CLK(I5694_clk), .RSTB(I132851_rst), .Q(I132813) );
nand I_7495 (I133148,I132868,I107725);
nand I_7496 (I133165,I133148,I132902);
and I_7497 (I133182,I132984,I133165);
DFFARX1 I_7498  ( .D(I133182), .CLK(I5694_clk), .RSTB(I132851_rst), .Q(I132843) );
and I_7499 (I132816,I133148,I133117);
DFFARX1 I_7500  ( .D(I107719), .CLK(I5694_clk), .RSTB(I132851_rst), .Q(I133227) );
nor I_7501 (I132840,I133227,I133148);
nor I_7502 (I133258,I133227,I132902);
nand I_7503 (I132837,I132936,I133258);
not I_7504 (I132834,I133227);
DFFARX1 I_7505  ( .D(I107722), .CLK(I5694_clk), .RSTB(I132851_rst), .Q(I133303) );
not I_7506 (I133320,I133303);
nor I_7507 (I133337,I133320,I133001);
and I_7508 (I133354,I133227,I133337);
or I_7509 (I133371,I133148,I133354);
DFFARX1 I_7510  ( .D(I133371), .CLK(I5694_clk), .RSTB(I132851_rst), .Q(I132828) );
not I_7511 (I133402,I133320);
nor I_7512 (I13341_rst9,I133227,I133402);
nand I_7513 (I132831,I133320,I13341_rst9);
nand I_7514 (I132825,I132984,I133402);
not I_7515 (I133497_rst,I5701);
not I_7516 (I133514,I120376);
nor I_7517 (I133531,I120355,I120367);
nand I_7518 (I133548,I133531,I120370);
nor I_7519 (I133565,I133514,I120355);
nand I_7520 (I133582,I133565,I120352);
DFFARX1 I_7521  ( .D(I133582), .CLK(I5694_clk), .RSTB(I133497_rst), .Q(I133599) );
not I_7522 (I133468,I133599);
not I_7523 (I133630,I120355);
not I_7524 (I133647,I133630);
not I_7525 (I133664,I120373);
nor I_7526 (I133681,I133664,I120364);
and I_7527 (I133698,I133681,I120358);
or I_7528 (I133715,I133698,I120382);
DFFARX1 I_7529  ( .D(I133715), .CLK(I5694_clk), .RSTB(I133497_rst), .Q(I133732) );
DFFARX1 I_7530  ( .D(I133732), .CLK(I5694_clk), .RSTB(I133497_rst), .Q(I133465) );
DFFARX1 I_7531  ( .D(I133732), .CLK(I5694_clk), .RSTB(I133497_rst), .Q(I133763) );
DFFARX1 I_7532  ( .D(I133732), .CLK(I5694_clk), .RSTB(I133497_rst), .Q(I133459) );
nand I_7533 (I133794,I133514,I120373);
nand I_7534 (I133811,I133794,I133548);
and I_7535 (I133828,I133630,I133811);
DFFARX1 I_7536  ( .D(I133828), .CLK(I5694_clk), .RSTB(I133497_rst), .Q(I133489) );
and I_7537 (I133462,I133794,I133763);
DFFARX1 I_7538  ( .D(I120379), .CLK(I5694_clk), .RSTB(I133497_rst), .Q(I133873) );
nor I_7539 (I133486,I133873,I133794);
nor I_7540 (I133904,I133873,I133548);
nand I_7541 (I133483,I133582,I133904);
not I_7542 (I133480,I133873);
DFFARX1 I_7543  ( .D(I120361), .CLK(I5694_clk), .RSTB(I133497_rst), .Q(I133949) );
not I_7544 (I133966,I133949);
nor I_7545 (I133983,I133966,I133647);
and I_7546 (I134000,I133873,I133983);
or I_7547 (I134017,I133794,I134000);
DFFARX1 I_7548  ( .D(I134017), .CLK(I5694_clk), .RSTB(I133497_rst), .Q(I133474) );
not I_7549 (I134048,I133966);
nor I_7550 (I134065,I133873,I134048);
nand I_7551 (I133477,I133966,I134065);
nand I_7552 (I133471,I133630,I134048);
not I_7553 (I134143_rst,I5701);
not I_7554 (I134160,I101911);
nor I_7555 (I134177,I101902,I101893);
nand I_7556 (I134194,I134177,I101908);
nor I_7557 (I134211,I134160,I101902);
nand I_7558 (I134228,I134211,I101905);
DFFARX1 I_7559  ( .D(I134228), .CLK(I5694_clk), .RSTB(I134143_rst), .Q(I134245) );
not I_7560 (I134114,I134245);
not I_7561 (I134276,I101902);
not I_7562 (I134293,I134276);
not I_7563 (I134310,I101914);
nor I_7564 (I134327,I134310,I101899);
and I_7565 (I134344,I134327,I101917);
or I_7566 (I134361,I134344,I101890);
DFFARX1 I_7567  ( .D(I134361), .CLK(I5694_clk), .RSTB(I134143_rst), .Q(I134378) );
DFFARX1 I_7568  ( .D(I134378), .CLK(I5694_clk), .RSTB(I134143_rst), .Q(I134111) );
DFFARX1 I_7569  ( .D(I134378), .CLK(I5694_clk), .RSTB(I134143_rst), .Q(I134409) );
DFFARX1 I_7570  ( .D(I134378), .CLK(I5694_clk), .RSTB(I134143_rst), .Q(I134105) );
nand I_7571 (I134440,I134160,I101914);
nand I_7572 (I134457,I134440,I134194);
and I_7573 (I134474,I134276,I134457);
DFFARX1 I_7574  ( .D(I134474), .CLK(I5694_clk), .RSTB(I134143_rst), .Q(I134135) );
and I_7575 (I134108,I134440,I134409);
DFFARX1 I_7576  ( .D(I101920), .CLK(I5694_clk), .RSTB(I134143_rst), .Q(I134519) );
nor I_7577 (I134132,I134519,I134440);
nor I_7578 (I134550,I134519,I134194);
nand I_7579 (I134129,I134228,I134550);
not I_7580 (I134126,I134519);
DFFARX1 I_7581  ( .D(I101896), .CLK(I5694_clk), .RSTB(I134143_rst), .Q(I134595) );
not I_7582 (I134612,I134595);
nor I_7583 (I134629,I134612,I134293);
and I_7584 (I134646,I134519,I134629);
or I_7585 (I134663,I134440,I134646);
DFFARX1 I_7586  ( .D(I134663), .CLK(I5694_clk), .RSTB(I134143_rst), .Q(I134120) );
not I_7587 (I134694,I134612);
nor I_7588 (I134711,I134519,I134694);
nand I_7589 (I134123,I134612,I134711);
nand I_7590 (I134117,I134276,I134694);
not I_7591 (I134789_rst,I5701);
not I_7592 (I134806,I97547);
nor I_7593 (I134823,I97562,I97556);
nand I_7594 (I134840,I134823,I97565);
nor I_7595 (I134857,I134806,I97562);
nand I_7596 (I134874,I134857,I97541);
DFFARX1 I_7597  ( .D(I134874), .CLK(I5694_clk), .RSTB(I134789_rst), .Q(I134891) );
not I_7598 (I134760,I134891);
not I_7599 (I134922,I97562);
not I_7600 (I134939,I134922);
not I_7601 (I134956,I97538);
nor I_7602 (I134973,I134956,I97553);
and I_7603 (I134990,I134973,I97559);
or I_7604 (I135007,I134990,I97568);
DFFARX1 I_7605  ( .D(I135007), .CLK(I5694_clk), .RSTB(I134789_rst), .Q(I135024) );
DFFARX1 I_7606  ( .D(I135024), .CLK(I5694_clk), .RSTB(I134789_rst), .Q(I134757) );
DFFARX1 I_7607  ( .D(I135024), .CLK(I5694_clk), .RSTB(I134789_rst), .Q(I135055) );
DFFARX1 I_7608  ( .D(I135024), .CLK(I5694_clk), .RSTB(I134789_rst), .Q(I134751) );
nand I_7609 (I135086,I134806,I97538);
nand I_7610 (I135103,I135086,I134840);
and I_7611 (I135120,I134922,I135103);
DFFARX1 I_7612  ( .D(I135120), .CLK(I5694_clk), .RSTB(I134789_rst), .Q(I134781) );
and I_7613 (I134754,I135086,I135055);
DFFARX1 I_7614  ( .D(I97550), .CLK(I5694_clk), .RSTB(I134789_rst), .Q(I135165) );
nor I_7615 (I134778,I135165,I135086);
nor I_7616 (I135196,I135165,I134840);
nand I_7617 (I134775,I134874,I135196);
not I_7618 (I134772,I135165);
DFFARX1 I_7619  ( .D(I97544), .CLK(I5694_clk), .RSTB(I134789_rst), .Q(I135241) );
not I_7620 (I135258,I135241);
nor I_7621 (I135275,I135258,I134939);
and I_7622 (I135292,I135165,I135275);
or I_7623 (I135309,I135086,I135292);
DFFARX1 I_7624  ( .D(I135309), .CLK(I5694_clk), .RSTB(I134789_rst), .Q(I134766) );
not I_7625 (I135340,I135258);
nor I_7626 (I135357,I135165,I135340);
nand I_7627 (I134769,I135258,I135357);
nand I_7628 (I134763,I134922,I135340);
not I_7629 (I135435_rst,I5701);
not I_7630 (I135452,I111022);
nor I_7631 (I135469,I111043,I111025);
nand I_7632 (I135486,I135469,I111049);
nor I_7633 (I135503,I135452,I111043);
nand I_7634 (I135520,I135503,I111046);
DFFARX1 I_7635  ( .D(I135520), .CLK(I5694_clk), .RSTB(I135435_rst), .Q(I135537) );
not I_7636 (I135406,I135537);
not I_7637 (I135568,I111043);
not I_7638 (I135585,I135568);
not I_7639 (I135602,I111040);
nor I_7640 (I135619,I135602,I111019);
and I_7641 (I135636,I135619,I111031);
or I_7642 (I135653,I135636,I111028);
DFFARX1 I_7643  ( .D(I135653), .CLK(I5694_clk), .RSTB(I135435_rst), .Q(I135670) );
DFFARX1 I_7644  ( .D(I135670), .CLK(I5694_clk), .RSTB(I135435_rst), .Q(I135403) );
DFFARX1 I_7645  ( .D(I135670), .CLK(I5694_clk), .RSTB(I135435_rst), .Q(I135701) );
DFFARX1 I_7646  ( .D(I135670), .CLK(I5694_clk), .RSTB(I135435_rst), .Q(I135397) );
nand I_7647 (I135732,I135452,I111040);
nand I_7648 (I135749,I135732,I135486);
and I_7649 (I135766,I135568,I135749);
DFFARX1 I_7650  ( .D(I135766), .CLK(I5694_clk), .RSTB(I135435_rst), .Q(I135427) );
and I_7651 (I135400,I135732,I135701);
DFFARX1 I_7652  ( .D(I111034), .CLK(I5694_clk), .RSTB(I135435_rst), .Q(I135811) );
nor I_7653 (I135424,I135811,I135732);
nor I_7654 (I135842,I135811,I135486);
nand I_7655 (I135421,I135520,I135842);
not I_7656 (I135418,I135811);
DFFARX1 I_7657  ( .D(I111037), .CLK(I5694_clk), .RSTB(I135435_rst), .Q(I135887) );
not I_7658 (I135904,I135887);
nor I_7659 (I135921,I135904,I135585);
and I_7660 (I135938,I135811,I135921);
or I_7661 (I135955,I135732,I135938);
DFFARX1 I_7662  ( .D(I135955), .CLK(I5694_clk), .RSTB(I135435_rst), .Q(I135412) );
not I_7663 (I135986,I135904);
nor I_7664 (I136003,I135811,I135986);
nand I_7665 (I135415,I135904,I136003);
nand I_7666 (I135409,I135568,I135986);
not I_7667 (I136081_rst,I5701);
not I_7668 (I136098,I123028);
nor I_7669 (I136115,I123007,I123019);
nand I_7670 (I136132,I136115,I123022);
nor I_7671 (I136149,I136098,I123007);
nand I_7672 (I136166,I136149,I123004);
DFFARX1 I_7673  ( .D(I136166), .CLK(I5694_clk), .RSTB(I136081_rst), .Q(I136183) );
not I_7674 (I136052,I136183);
not I_7675 (I136214,I123007);
not I_7676 (I136231,I136214);
not I_7677 (I136248,I123025);
nor I_7678 (I136265,I136248,I123016);
and I_7679 (I136282,I136265,I123010);
or I_7680 (I136299,I136282,I123034);
DFFARX1 I_7681  ( .D(I136299), .CLK(I5694_clk), .RSTB(I136081_rst), .Q(I136316) );
DFFARX1 I_7682  ( .D(I136316), .CLK(I5694_clk), .RSTB(I136081_rst), .Q(I136049) );
DFFARX1 I_7683  ( .D(I136316), .CLK(I5694_clk), .RSTB(I136081_rst), .Q(I136347) );
DFFARX1 I_7684  ( .D(I136316), .CLK(I5694_clk), .RSTB(I136081_rst), .Q(I136043) );
nand I_7685 (I136378,I136098,I123025);
nand I_7686 (I136395,I136378,I136132);
and I_7687 (I136412,I136214,I136395);
DFFARX1 I_7688  ( .D(I136412), .CLK(I5694_clk), .RSTB(I136081_rst), .Q(I136073) );
and I_7689 (I136046,I136378,I136347);
DFFARX1 I_7690  ( .D(I123031), .CLK(I5694_clk), .RSTB(I136081_rst), .Q(I136457) );
nor I_7691 (I136070,I136457,I136378);
nor I_7692 (I136488,I136457,I136132);
nand I_7693 (I136067,I136166,I136488);
not I_7694 (I136064,I136457);
DFFARX1 I_7695  ( .D(I123013), .CLK(I5694_clk), .RSTB(I136081_rst), .Q(I136533) );
not I_7696 (I136550,I136533);
nor I_7697 (I136567,I136550,I136231);
and I_7698 (I136584,I136457,I136567);
or I_7699 (I136601,I136378,I136584);
DFFARX1 I_7700  ( .D(I136601), .CLK(I5694_clk), .RSTB(I136081_rst), .Q(I136058) );
not I_7701 (I136632,I136550);
nor I_7702 (I136649,I136457,I136632);
nand I_7703 (I136061,I136550,I136649);
nand I_7704 (I136055,I136214,I136632);
not I_7705 (I136727_rst,I5701);
or I_7706 (I136744,I75974,I75986);
or I_7707 (I136761,I75989,I75974);
nor I_7708 (I136778,I75971,I75965);
DFFARX1 I_7709  ( .D(I136778), .CLK(I5694_clk), .RSTB(I136727_rst), .Q(I136795) );
DFFARX1 I_7710  ( .D(I136778), .CLK(I5694_clk), .RSTB(I136727_rst), .Q(I136689) );
not I_7711 (I136826,I75971);
and I_7712 (I136843,I136826,I75977);
nor I_7713 (I136860,I136843,I75986);
nor I_7714 (I136877,I75980,I75983);
DFFARX1 I_7715  ( .D(I136877), .CLK(I5694_clk), .RSTB(I136727_rst), .Q(I136894) );
not I_7716 (I136911,I136894);
DFFARX1 I_7717  ( .D(I136894), .CLK(I5694_clk), .RSTB(I136727_rst), .Q(I136698) );
nor I_7718 (I136942,I75980,I75989);
and I_7719 (I136692,I136942,I136795);
DFFARX1 I_7720  ( .D(I75995), .CLK(I5694_clk), .RSTB(I136727_rst), .Q(I136973) );
and I_7721 (I136990,I136973,I75968);
nand I_7722 (I137007,I136990,I136761);
and I_7723 (I137024,I136894,I137007);
DFFARX1 I_7724  ( .D(I137024), .CLK(I5694_clk), .RSTB(I136727_rst), .Q(I136719) );
nor I_7725 (I136716,I136990,I136860);
not I_7726 (I137069,I136990);
nor I_7727 (I137086,I136744,I137069);
nor I_7728 (I137103,I136990,I136942);
nand I_7729 (I136713,I136761,I137103);
nor I_7730 (I137134,I136990,I136911);
not I_7731 (I136710,I136990);
nand I_7732 (I136701,I136990,I136911);
DFFARX1 I_7733  ( .D(I75992), .CLK(I5694_clk), .RSTB(I136727_rst), .Q(I137179) );
and I_7734 (I137196,I137179,I137086);
or I_7735 (I137213,I136744,I137196);
DFFARX1 I_7736  ( .D(I137213), .CLK(I5694_clk), .RSTB(I136727_rst), .Q(I136704) );
nand I_7737 (I136707,I137179,I137134);
nand I_7738 (I137258,I137179,I136860);
and I_7739 (I137275,I136778,I137258);
DFFARX1 I_7740  ( .D(I137275), .CLK(I5694_clk), .RSTB(I136727_rst), .Q(I136695) );
not I_7741 (I137339_rst,I5701);
or I_7742 (I137356,I105766,I105793);
or I_7743 (I137373,I105781,I105766);
nor I_7744 (I137390,I105790,I105769);
DFFARX1 I_7745  ( .D(I137390), .CLK(I5694_clk), .RSTB(I137339_rst), .Q(I137407) );
DFFARX1 I_7746  ( .D(I137390), .CLK(I5694_clk), .RSTB(I137339_rst), .Q(I137301) );
not I_7747 (I137438,I105790);
and I_7748 (I137455,I137438,I105787);
nor I_7749 (I137472,I137455,I105793);
nor I_7750 (I137489,I105784,I105772);
DFFARX1 I_7751  ( .D(I137489), .CLK(I5694_clk), .RSTB(I137339_rst), .Q(I137506) );
not I_7752 (I137523,I137506);
DFFARX1 I_7753  ( .D(I137506), .CLK(I5694_clk), .RSTB(I137339_rst), .Q(I137310) );
nor I_7754 (I137554,I105784,I105781);
and I_7755 (I137304,I137554,I137407);
DFFARX1 I_7756  ( .D(I105796), .CLK(I5694_clk), .RSTB(I137339_rst), .Q(I137585) );
and I_7757 (I137602,I137585,I105778);
nand I_7758 (I137619,I137602,I137373);
and I_7759 (I137636,I137506,I137619);
DFFARX1 I_7760  ( .D(I137636), .CLK(I5694_clk), .RSTB(I137339_rst), .Q(I137331) );
nor I_7761 (I137328,I137602,I137472);
not I_7762 (I137681,I137602);
nor I_7763 (I137698,I137356,I137681);
nor I_7764 (I137715,I137602,I137554);
nand I_7765 (I137325,I137373,I137715);
nor I_7766 (I137746,I137602,I137523);
not I_7767 (I137322,I137602);
nand I_7768 (I137313,I137602,I137523);
DFFARX1 I_7769  ( .D(I105775), .CLK(I5694_clk), .RSTB(I137339_rst), .Q(I137791) );
and I_7770 (I137808,I137791,I137698);
or I_7771 (I137825,I137356,I137808);
DFFARX1 I_7772  ( .D(I137825), .CLK(I5694_clk), .RSTB(I137339_rst), .Q(I137316) );
nand I_7773 (I137319,I137791,I137746);
nand I_7774 (I137870,I137791,I137472);
and I_7775 (I137887,I137390,I137870);
DFFARX1 I_7776  ( .D(I137887), .CLK(I5694_clk), .RSTB(I137339_rst), .Q(I137307) );
not I_7777 (I137951_rst,I5701);
nand I_7778 (I137968,I118431,I118434);
and I_7779 (I137985,I137968,I118440);
DFFARX1 I_7780  ( .D(I137985), .CLK(I5694_clk), .RSTB(I137951_rst), .Q(I138002) );
not I_7781 (I138019,I138002);
DFFARX1 I_7782  ( .D(I138002), .CLK(I5694_clk), .RSTB(I137951_rst), .Q(I137919) );
nor I_7783 (I138050,I118452,I118434);
DFFARX1 I_7784  ( .D(I118443), .CLK(I5694_clk), .RSTB(I137951_rst), .Q(I138067) );
DFFARX1 I_7785  ( .D(I138067), .CLK(I5694_clk), .RSTB(I137951_rst), .Q(I138084) );
not I_7786 (I137922,I138084);
DFFARX1 I_7787  ( .D(I138067), .CLK(I5694_clk), .RSTB(I137951_rst), .Q(I138115) );
and I_7788 (I137916,I138002,I138115);
nand I_7789 (I138146,I118449,I118446);
and I_7790 (I138163,I138146,I118458);
DFFARX1 I_7791  ( .D(I138163), .CLK(I5694_clk), .RSTB(I137951_rst), .Q(I138180) );
nor I_7792 (I138197,I138180,I138019);
not I_7793 (I138214,I138180);
nand I_7794 (I137925,I138002,I138214);
DFFARX1 I_7795  ( .D(I118455), .CLK(I5694_clk), .RSTB(I137951_rst), .Q(I138245) );
and I_7796 (I138262,I138245,I118461);
nor I_7797 (I138279,I138262,I138180);
nor I_7798 (I138296,I138262,I138214);
nand I_7799 (I137931,I138050,I138296);
not I_7800 (I137934,I138262);
DFFARX1 I_7801  ( .D(I138262), .CLK(I5694_clk), .RSTB(I137951_rst), .Q(I137913) );
DFFARX1 I_7802  ( .D(I118437), .CLK(I5694_clk), .RSTB(I137951_rst), .Q(I138355) );
nand I_7803 (I138372,I138355,I138067);
and I_7804 (I138389,I138050,I138372);
DFFARX1 I_7805  ( .D(I138389), .CLK(I5694_clk), .RSTB(I137951_rst), .Q(I137943) );
nor I_7806 (I137940,I138355,I138262);
and I_7807 (I138434,I138355,I138197);
or I_7808 (I138451,I138050,I138434);
DFFARX1 I_7809  ( .D(I138451), .CLK(I5694_clk), .RSTB(I137951_rst), .Q(I137928) );
nand I_7810 (I137937,I138355,I138279);
not I_7811 (I138529_rst,I5701);
nand I_7812 (I138546,I88189,I88192);
and I_7813 (I138563,I138546,I88198);
DFFARX1 I_7814  ( .D(I138563), .CLK(I5694_clk), .RSTB(I138529_rst), .Q(I138580) );
not I_7815 (I138597,I138580);
DFFARX1 I_7816  ( .D(I138580), .CLK(I5694_clk), .RSTB(I138529_rst), .Q(I138497) );
nor I_7817 (I138628,I88195,I88192);
DFFARX1 I_7818  ( .D(I88174), .CLK(I5694_clk), .RSTB(I138529_rst), .Q(I138645) );
DFFARX1 I_7819  ( .D(I138645), .CLK(I5694_clk), .RSTB(I138529_rst), .Q(I138662) );
not I_7820 (I138500,I138662);
DFFARX1 I_7821  ( .D(I138645), .CLK(I5694_clk), .RSTB(I138529_rst), .Q(I138693) );
and I_7822 (I138494,I138580,I138693);
nand I_7823 (I138724,I88171,I88186);
and I_7824 (I138741,I138724,I88183);
DFFARX1 I_7825  ( .D(I138741), .CLK(I5694_clk), .RSTB(I138529_rst), .Q(I138758) );
nor I_7826 (I138775,I138758,I138597);
not I_7827 (I138792,I138758);
nand I_7828 (I138503,I138580,I138792);
DFFARX1 I_7829  ( .D(I88201), .CLK(I5694_clk), .RSTB(I138529_rst), .Q(I138823) );
and I_7830 (I138840,I138823,I88180);
nor I_7831 (I138857,I138840,I138758);
nor I_7832 (I138874,I138840,I138792);
nand I_7833 (I138509,I138628,I138874);
not I_7834 (I138512,I138840);
DFFARX1 I_7835  ( .D(I138840), .CLK(I5694_clk), .RSTB(I138529_rst), .Q(I138491) );
DFFARX1 I_7836  ( .D(I88177), .CLK(I5694_clk), .RSTB(I138529_rst), .Q(I138933) );
nand I_7837 (I138950,I138933,I138645);
and I_7838 (I138967,I138628,I138950);
DFFARX1 I_7839  ( .D(I138967), .CLK(I5694_clk), .RSTB(I138529_rst), .Q(I138521) );
nor I_7840 (I138518,I138933,I138840);
and I_7841 (I139012,I138933,I138775);
or I_7842 (I139029,I138628,I139012);
DFFARX1 I_7843  ( .D(I139029), .CLK(I5694_clk), .RSTB(I138529_rst), .Q(I138506) );
nand I_7844 (I138515,I138933,I138857);
not I_7845 (I139107_rst,I5701);
nand I_7846 (I139124,I137301,I137331);
and I_7847 (I139141,I139124,I137328);
DFFARX1 I_7848  ( .D(I139141), .CLK(I5694_clk), .RSTB(I139107_rst), .Q(I139158) );
not I_7849 (I139175,I139158);
DFFARX1 I_7850  ( .D(I139158), .CLK(I5694_clk), .RSTB(I139107_rst), .Q(I139075) );
nor I_7851 (I139206,I137319,I137331);
DFFARX1 I_7852  ( .D(I137307), .CLK(I5694_clk), .RSTB(I139107_rst), .Q(I139223) );
DFFARX1 I_7853  ( .D(I139223), .CLK(I5694_clk), .RSTB(I139107_rst), .Q(I139240) );
not I_7854 (I139078,I139240);
DFFARX1 I_7855  ( .D(I139223), .CLK(I5694_clk), .RSTB(I139107_rst), .Q(I139271) );
and I_7856 (I139072,I139158,I139271);
nand I_7857 (I139302,I137310,I137316);
and I_7858 (I139319,I139302,I137322);
DFFARX1 I_7859  ( .D(I139319), .CLK(I5694_clk), .RSTB(I139107_rst), .Q(I139336) );
nor I_7860 (I139353,I139336,I139175);
not I_7861 (I139370,I139336);
nand I_7862 (I139081,I139158,I139370);
DFFARX1 I_7863  ( .D(I137313), .CLK(I5694_clk), .RSTB(I139107_rst), .Q(I139401) );
and I_7864 (I139418,I139401,I137304);
nor I_7865 (I139435,I139418,I139336);
nor I_7866 (I139452,I139418,I139370);
nand I_7867 (I139087,I139206,I139452);
not I_7868 (I139090,I139418);
DFFARX1 I_7869  ( .D(I139418), .CLK(I5694_clk), .RSTB(I139107_rst), .Q(I139069) );
DFFARX1 I_7870  ( .D(I137325), .CLK(I5694_clk), .RSTB(I139107_rst), .Q(I139511) );
nand I_7871 (I139528,I139511,I139223);
and I_7872 (I139545,I139206,I139528);
DFFARX1 I_7873  ( .D(I139545), .CLK(I5694_clk), .RSTB(I139107_rst), .Q(I139099) );
nor I_7874 (I139096,I139511,I139418);
and I_7875 (I139590,I139511,I139353);
or I_7876 (I139607,I139206,I139590);
DFFARX1 I_7877  ( .D(I139607), .CLK(I5694_clk), .RSTB(I139107_rst), .Q(I139084) );
nand I_7878 (I139093,I139511,I139435);
not I_7879 (I139685_rst,I5701);
nand I_7880 (I139702,I85673,I85676);
and I_7881 (I139719,I139702,I85682);
DFFARX1 I_7882  ( .D(I139719), .CLK(I5694_clk), .RSTB(I139685_rst), .Q(I139736) );
not I_7883 (I139753,I139736);
DFFARX1 I_7884  ( .D(I139736), .CLK(I5694_clk), .RSTB(I139685_rst), .Q(I139653) );
nor I_7885 (I139784,I85679,I85676);
DFFARX1 I_7886  ( .D(I85658), .CLK(I5694_clk), .RSTB(I139685_rst), .Q(I139801) );
DFFARX1 I_7887  ( .D(I139801), .CLK(I5694_clk), .RSTB(I139685_rst), .Q(I139818) );
not I_7888 (I139656,I139818);
DFFARX1 I_7889  ( .D(I139801), .CLK(I5694_clk), .RSTB(I139685_rst), .Q(I139849) );
and I_7890 (I139650,I139736,I139849);
nand I_7891 (I139880,I85655,I85670);
and I_7892 (I139897,I139880,I85667);
DFFARX1 I_7893  ( .D(I139897), .CLK(I5694_clk), .RSTB(I139685_rst), .Q(I139914) );
nor I_7894 (I139931,I139914,I139753);
not I_7895 (I139948,I139914);
nand I_7896 (I139659,I139736,I139948);
DFFARX1 I_7897  ( .D(I85685), .CLK(I5694_clk), .RSTB(I139685_rst), .Q(I139979) );
and I_7898 (I139996,I139979,I85664);
nor I_7899 (I140013,I139996,I139914);
nor I_7900 (I140030,I139996,I139948);
nand I_7901 (I139665,I139784,I140030);
not I_7902 (I139668,I139996);
DFFARX1 I_7903  ( .D(I139996), .CLK(I5694_clk), .RSTB(I139685_rst), .Q(I139647) );
DFFARX1 I_7904  ( .D(I85661), .CLK(I5694_clk), .RSTB(I139685_rst), .Q(I140089) );
nand I_7905 (I140106,I140089,I139801);
and I_7906 (I140123,I139784,I140106);
DFFARX1 I_7907  ( .D(I140123), .CLK(I5694_clk), .RSTB(I139685_rst), .Q(I139677) );
nor I_7908 (I139674,I140089,I139996);
and I_7909 (I140168,I140089,I139931);
or I_7910 (I140185,I139784,I140168);
DFFARX1 I_7911  ( .D(I140185), .CLK(I5694_clk), .RSTB(I139685_rst), .Q(I139662) );
nand I_7912 (I139671,I140089,I140013);
not I_7913 (I140263_rst,I5701);
or I_7914 (I140280,I88827,I88821);
or I_7915 (I140297,I88830,I88827);
nor I_7916 (I140314,I88824,I88806);
not I_7917 (I140331,I140314);
DFFARX1 I_7918  ( .D(I140314), .CLK(I5694_clk), .RSTB(I140263_rst), .Q(I140231) );
nand I_7919 (I140362,I140314,I140280);
not I_7920 (I140379,I88824);
and I_7921 (I140396,I140379,I88803);
nor I_7922 (I140413,I140396,I88821);
nor I_7923 (I140430,I88818,I88800);
DFFARX1 I_7924  ( .D(I140430), .CLK(I5694_clk), .RSTB(I140263_rst), .Q(I140447) );
nor I_7925 (I140464,I140447,I140331);
not I_7926 (I140481,I140447);
nand I_7927 (I140237,I140314,I140481);
DFFARX1 I_7928  ( .D(I140447), .CLK(I5694_clk), .RSTB(I140263_rst), .Q(I140228) );
nor I_7929 (I140526,I88818,I88830);
nand I_7930 (I140543,I140297,I140526);
nor I_7931 (I140252,I140280,I140526);
and I_7932 (I140574,I140526,I140464);
or I_7933 (I140591,I140413,I140574);
DFFARX1 I_7934  ( .D(I140591), .CLK(I5694_clk), .RSTB(I140263_rst), .Q(I140240) );
DFFARX1 I_7935  ( .D(I88812), .CLK(I5694_clk), .RSTB(I140263_rst), .Q(I140622) );
and I_7936 (I140639,I140622,I88815);
not I_7937 (I140246,I140639);
DFFARX1 I_7938  ( .D(I140639), .CLK(I5694_clk), .RSTB(I140263_rst), .Q(I140670) );
not I_7939 (I140234,I140670);
and I_7940 (I140701,I140639,I140362);
DFFARX1 I_7941  ( .D(I140701), .CLK(I5694_clk), .RSTB(I140263_rst), .Q(I140225) );
DFFARX1 I_7942  ( .D(I88809), .CLK(I5694_clk), .RSTB(I140263_rst), .Q(I140732) );
and I_7943 (I140749,I140732,I140543);
DFFARX1 I_7944  ( .D(I140749), .CLK(I5694_clk), .RSTB(I140263_rst), .Q(I140255) );
nor I_7945 (I140780,I140732,I140639);
nand I_7946 (I140249,I140413,I140780);
nor I_7947 (I140811,I140732,I140481);
nand I_7948 (I140243,I140297,I140811);
not I_7949 (I140875_rst,I5701);
or I_7950 (I140892,I113017,I113008);
or I_7951 (I140909,I113020,I113017);
nor I_7952 (I140926,I113035,I113011);
not I_7953 (I140943,I140926);
DFFARX1 I_7954  ( .D(I140926), .CLK(I5694_clk), .RSTB(I140875_rst), .Q(I140843) );
nand I_7955 (I140974,I140926,I140892);
not I_7956 (I140991,I113035);
and I_7957 (I141008,I140991,I113032);
nor I_7958 (I141025,I141008,I113008);
nor I_7959 (I141042,I113029,I113014);
DFFARX1 I_7960  ( .D(I141042), .CLK(I5694_clk), .RSTB(I140875_rst), .Q(I141059) );
nor I_7961 (I141076,I141059,I140943);
not I_7962 (I141093,I141059);
nand I_7963 (I140849,I140926,I141093);
DFFARX1 I_7964  ( .D(I141059), .CLK(I5694_clk), .RSTB(I140875_rst), .Q(I140840) );
nor I_7965 (I141138,I113029,I113020);
nand I_7966 (I141155,I140909,I141138);
nor I_7967 (I140864,I140892,I141138);
and I_7968 (I141186,I141138,I141076);
or I_7969 (I141203,I141025,I141186);
DFFARX1 I_7970  ( .D(I141203), .CLK(I5694_clk), .RSTB(I140875_rst), .Q(I140852) );
DFFARX1 I_7971  ( .D(I113038), .CLK(I5694_clk), .RSTB(I140875_rst), .Q(I141234) );
and I_7972 (I141251,I141234,I113023);
not I_7973 (I140858,I141251);
DFFARX1 I_7974  ( .D(I141251), .CLK(I5694_clk), .RSTB(I140875_rst), .Q(I141282) );
not I_7975 (I140846,I141282);
and I_7976 (I141313,I141251,I140974);
DFFARX1 I_7977  ( .D(I141313), .CLK(I5694_clk), .RSTB(I140875_rst), .Q(I140837) );
DFFARX1 I_7978  ( .D(I113026), .CLK(I5694_clk), .RSTB(I140875_rst), .Q(I141344) );
and I_7979 (I141361,I141344,I141155);
DFFARX1 I_7980  ( .D(I141361), .CLK(I5694_clk), .RSTB(I140875_rst), .Q(I140867) );
nor I_7981 (I141392,I141344,I141251);
nand I_7982 (I140861,I141025,I141392);
nor I_7983 (I141423,I141344,I141093);
nand I_7984 (I140855,I140909,I141423);
not I_7985 (I141487_rst,I5701);
or I_7986 (I141504,I104498,I104489);
or I_7987 (I141521,I104486,I104498);
nor I_7988 (I141538,I104483,I104501);
not I_7989 (I141555,I141538);
DFFARX1 I_7990  ( .D(I141538), .CLK(I5694_clk), .RSTB(I141487_rst), .Q(I141455) );
nand I_7991 (I141586,I141538,I141504);
not I_7992 (I141603,I104483);
and I_7993 (I141620,I141603,I104474);
nor I_7994 (I141637,I141620,I104489);
nor I_7995 (I141654,I104477,I104480);
DFFARX1 I_7996  ( .D(I141654), .CLK(I5694_clk), .RSTB(I141487_rst), .Q(I141671) );
nor I_7997 (I141688,I141671,I141555);
not I_7998 (I141705,I141671);
nand I_7999 (I141461,I141538,I141705);
DFFARX1 I_8000  ( .D(I141671), .CLK(I5694_clk), .RSTB(I141487_rst), .Q(I141452) );
nor I_8001 (I141750,I104477,I104486);
nand I_8002 (I141767,I141521,I141750);
nor I_8003 (I141476,I141504,I141750);
and I_8004 (I141798,I141750,I141688);
or I_8005 (I141815,I141637,I141798);
DFFARX1 I_8006  ( .D(I141815), .CLK(I5694_clk), .RSTB(I141487_rst), .Q(I141464) );
DFFARX1 I_8007  ( .D(I104492), .CLK(I5694_clk), .RSTB(I141487_rst), .Q(I141846) );
and I_8008 (I141863,I141846,I104504);
not I_8009 (I141470,I141863);
DFFARX1 I_8010  ( .D(I141863), .CLK(I5694_clk), .RSTB(I141487_rst), .Q(I141894) );
not I_8011 (I141458,I141894);
and I_8012 (I141925,I141863,I141586);
DFFARX1 I_8013  ( .D(I141925), .CLK(I5694_clk), .RSTB(I141487_rst), .Q(I141449) );
DFFARX1 I_8014  ( .D(I104495), .CLK(I5694_clk), .RSTB(I141487_rst), .Q(I141956) );
and I_8015 (I141973,I141956,I141767);
DFFARX1 I_8016  ( .D(I141973), .CLK(I5694_clk), .RSTB(I141487_rst), .Q(I141479) );
nor I_8017 (I142004,I141956,I141863);
nand I_8018 (I141473,I141637,I142004);
nor I_8019 (I142035,I141956,I141705);
nand I_8020 (I141467,I141521,I142035);
not I_8021 (I142099_rst,I5701);
or I_8022 (I142116,I73606,I73600);
or I_8023 (I142133,I73594,I73606);
nor I_8024 (I142150,I73615,I73603);
or I_8025 (I142088,I142150,I142116);
not I_8026 (I142181,I73615);
and I_8027 (I142198,I142181,I73588);
nor I_8028 (I142215,I142198,I73600);
not I_8029 (I142232,I142215);
nor I_8030 (I142249,I73591,I73585);
DFFARX1 I_8031  ( .D(I142249), .CLK(I5694_clk), .RSTB(I142099_rst), .Q(I142266) );
nor I_8032 (I142283,I142266,I142215);
nand I_8033 (I142073,I142116,I142283);
nor I_8034 (I142314,I142266,I142232);
not I_8035 (I142070,I142266);
nor I_8036 (I142345,I73591,I73594);
or I_8037 (I142082,I142116,I142345);
DFFARX1 I_8038  ( .D(I73612), .CLK(I5694_clk), .RSTB(I142099_rst), .Q(I142376) );
and I_8039 (I142393,I142376,I73609);
nor I_8040 (I142410,I142393,I142266);
DFFARX1 I_8041  ( .D(I142410), .CLK(I5694_clk), .RSTB(I142099_rst), .Q(I142076) );
nor I_8042 (I142091,I142393,I142345);
not I_8043 (I142455,I142393);
nor I_8044 (I142472,I142133,I142455);
nand I_8045 (I142061,I142393,I142232);
DFFARX1 I_8046  ( .D(I73597), .CLK(I5694_clk), .RSTB(I142099_rst), .Q(I142503) );
nor I_8047 (I142079,I142503,I142133);
not I_8048 (I142534,I142503);
and I_8049 (I142551,I142345,I142534);
nor I_8050 (I142085,I142150,I142551);
and I_8051 (I142582,I142503,I142472);
or I_8052 (I142599,I142150,I142582);
DFFARX1 I_8053  ( .D(I142599), .CLK(I5694_clk), .RSTB(I142099_rst), .Q(I142064) );
nand I_8054 (I142067,I142503,I142314);
not I_8055 (I142677_rst,I5701);
or I_8056 (I142694,I116051,I116057);
or I_8057 (I142711,I116060,I116051);
nor I_8058 (I142728,I116075,I116063);
or I_8059 (I142666,I142728,I142694);
not I_8060 (I142759,I116075);
and I_8061 (I142776,I142759,I116054);
nor I_8062 (I142793,I142776,I116057);
not I_8063 (I142810,I142793);
nor I_8064 (I142827,I116069,I116078);
DFFARX1 I_8065  ( .D(I142827), .CLK(I5694_clk), .RSTB(I142677_rst), .Q(I142844) );
nor I_8066 (I142861,I142844,I142793);
nand I_8067 (I142651,I142694,I142861);
nor I_8068 (I142892,I142844,I142810);
not I_8069 (I142648,I142844);
nor I_8070 (I142923,I116069,I116060);
or I_8071 (I142660,I142694,I142923);
DFFARX1 I_8072  ( .D(I116066), .CLK(I5694_clk), .RSTB(I142677_rst), .Q(I142954) );
and I_8073 (I142971,I142954,I116081);
nor I_8074 (I142988,I142971,I142844);
DFFARX1 I_8075  ( .D(I142988), .CLK(I5694_clk), .RSTB(I142677_rst), .Q(I142654) );
nor I_8076 (I142669,I142971,I142923);
not I_8077 (I143033,I142971);
nor I_8078 (I143050,I142711,I143033);
nand I_8079 (I142639,I142971,I142810);
DFFARX1 I_8080  ( .D(I116072), .CLK(I5694_clk), .RSTB(I142677_rst), .Q(I143081) );
nor I_8081 (I142657,I143081,I142711);
not I_8082 (I143112,I143081);
and I_8083 (I143129,I142923,I143112);
nor I_8084 (I142663,I142728,I143129);
and I_8085 (I143160,I143081,I143050);
or I_8086 (I143177,I142728,I143160);
DFFARX1 I_8087  ( .D(I143177), .CLK(I5694_clk), .RSTB(I142677_rst), .Q(I142642) );
nand I_8088 (I142645,I143081,I142892);
not I_8089 (I143255_rst,I5701);
nand I_8090 (I143272,I132185,I132197);
and I_8091 (I143289,I143272,I132179);
DFFARX1 I_8092  ( .D(I143289), .CLK(I5694_clk), .RSTB(I143255_rst), .Q(I143306) );
nor I_8093 (I143323,I132191,I132197);
nor I_8094 (I143340,I143323,I143306);
not I_8095 (I143238,I143323);
DFFARX1 I_8096  ( .D(I132176), .CLK(I5694_clk), .RSTB(I143255_rst), .Q(I143371) );
not I_8097 (I143388,I143371);
nor I_8098 (I143405,I143323,I143388);
nand I_8099 (I143241,I143371,I143340);
DFFARX1 I_8100  ( .D(I143371), .CLK(I5694_clk), .RSTB(I143255_rst), .Q(I143223) );
nand I_8101 (I143450,I132167,I132182);
and I_8102 (I143467,I143450,I132173);
DFFARX1 I_8103  ( .D(I143467), .CLK(I5694_clk), .RSTB(I143255_rst), .Q(I143484) );
nor I_8104 (I143244,I143484,I143306);
nand I_8105 (I143235,I143484,I143405);
DFFARX1 I_8106  ( .D(I132194), .CLK(I5694_clk), .RSTB(I143255_rst), .Q(I143529) );
and I_8107 (I143546,I143529,I132188);
DFFARX1 I_8108  ( .D(I143546), .CLK(I5694_clk), .RSTB(I143255_rst), .Q(I143563) );
not I_8109 (I143226,I143563);
nand I_8110 (I143594,I143546,I143484);
and I_8111 (I143611,I143306,I143594);
DFFARX1 I_8112  ( .D(I143611), .CLK(I5694_clk), .RSTB(I143255_rst), .Q(I143217) );
DFFARX1 I_8113  ( .D(I132170), .CLK(I5694_clk), .RSTB(I143255_rst), .Q(I143642) );
nand I_8114 (I143659,I143642,I143306);
and I_8115 (I143676,I143484,I143659);
DFFARX1 I_8116  ( .D(I143676), .CLK(I5694_clk), .RSTB(I143255_rst), .Q(I143247) );
not I_8117 (I143707,I143642);
nor I_8118 (I143724,I143323,I143707);
and I_8119 (I143741,I143642,I143724);
or I_8120 (I143758,I143546,I143741);
DFFARX1 I_8121  ( .D(I143758), .CLK(I5694_clk), .RSTB(I143255_rst), .Q(I143232) );
nand I_8122 (I143229,I143642,I143388);
DFFARX1 I_8123  ( .D(I143642), .CLK(I5694_clk), .RSTB(I143255_rst), .Q(I143220) );
not I_8124 (I143850_rst,I5701);
nand I_8125 (I143867,I83157,I83148);
and I_8126 (I143884,I143867,I83166);
DFFARX1 I_8127  ( .D(I143884), .CLK(I5694_clk), .RSTB(I143850_rst), .Q(I143901) );
nor I_8128 (I143918,I83163,I83148);
nor I_8129 (I143935,I143918,I143901);
not I_8130 (I143833,I143918);
DFFARX1 I_8131  ( .D(I83145), .CLK(I5694_clk), .RSTB(I143850_rst), .Q(I143966) );
not I_8132 (I143983,I143966);
nor I_8133 (I144000,I143918,I143983);
nand I_8134 (I143836,I143966,I143935);
DFFARX1 I_8135  ( .D(I143966), .CLK(I5694_clk), .RSTB(I143850_rst), .Q(I143818) );
nand I_8136 (I144045,I83154,I83169);
and I_8137 (I144062,I144045,I83160);
DFFARX1 I_8138  ( .D(I144062), .CLK(I5694_clk), .RSTB(I143850_rst), .Q(I144079) );
nor I_8139 (I143839,I144079,I143901);
nand I_8140 (I143830,I144079,I144000);
DFFARX1 I_8141  ( .D(I83142), .CLK(I5694_clk), .RSTB(I143850_rst), .Q(I144124) );
and I_8142 (I144141,I144124,I83151);
DFFARX1 I_8143  ( .D(I144141), .CLK(I5694_clk), .RSTB(I143850_rst), .Q(I144158) );
not I_8144 (I143821,I144158);
nand I_8145 (I144189,I144141,I144079);
and I_8146 (I144206,I143901,I144189);
DFFARX1 I_8147  ( .D(I144206), .CLK(I5694_clk), .RSTB(I143850_rst), .Q(I143812) );
DFFARX1 I_8148  ( .D(I83139), .CLK(I5694_clk), .RSTB(I143850_rst), .Q(I144237) );
nand I_8149 (I144254,I144237,I143901);
and I_8150 (I144271,I144079,I144254);
DFFARX1 I_8151  ( .D(I144271), .CLK(I5694_clk), .RSTB(I143850_rst), .Q(I143842) );
not I_8152 (I144302,I144237);
nor I_8153 (I144319,I143918,I144302);
and I_8154 (I144336,I144237,I144319);
or I_8155 (I144353,I144141,I144336);
DFFARX1 I_8156  ( .D(I144353), .CLK(I5694_clk), .RSTB(I143850_rst), .Q(I143827) );
nand I_8157 (I143824,I144237,I143983);
DFFARX1 I_8158  ( .D(I144237), .CLK(I5694_clk), .RSTB(I143850_rst), .Q(I143815) );
not I_8159 (I144445_rst,I5701);
nand I_8160 (I144462,I117256,I117253);
and I_8161 (I144479,I144462,I117250);
DFFARX1 I_8162  ( .D(I144479), .CLK(I5694_clk), .RSTB(I144445_rst), .Q(I144496) );
nor I_8163 (I144513,I117241,I117253);
nor I_8164 (I144530,I144513,I144496);
not I_8165 (I144428,I144513);
DFFARX1 I_8166  ( .D(I117259), .CLK(I5694_clk), .RSTB(I144445_rst), .Q(I144561) );
not I_8167 (I144578,I144561);
nor I_8168 (I144595,I144513,I144578);
nand I_8169 (I144431,I144561,I144530);
DFFARX1 I_8170  ( .D(I144561), .CLK(I5694_clk), .RSTB(I144445_rst), .Q(I144413) );
nand I_8171 (I144640,I117244,I117268);
and I_8172 (I144657,I144640,I117247);
DFFARX1 I_8173  ( .D(I144657), .CLK(I5694_clk), .RSTB(I144445_rst), .Q(I144674) );
nor I_8174 (I144434,I144674,I144496);
nand I_8175 (I144425,I144674,I144595);
DFFARX1 I_8176  ( .D(I117265), .CLK(I5694_clk), .RSTB(I144445_rst), .Q(I144719) );
and I_8177 (I144736,I144719,I117262);
DFFARX1 I_8178  ( .D(I144736), .CLK(I5694_clk), .RSTB(I144445_rst), .Q(I144753) );
not I_8179 (I144416,I144753);
nand I_8180 (I144784,I144736,I144674);
and I_8181 (I144801,I144496,I144784);
DFFARX1 I_8182  ( .D(I144801), .CLK(I5694_clk), .RSTB(I144445_rst), .Q(I144407) );
DFFARX1 I_8183  ( .D(I117271), .CLK(I5694_clk), .RSTB(I144445_rst), .Q(I144832) );
nand I_8184 (I144849,I144832,I144496);
and I_8185 (I144866,I144674,I144849);
DFFARX1 I_8186  ( .D(I144866), .CLK(I5694_clk), .RSTB(I144445_rst), .Q(I144437) );
not I_8187 (I144897,I144832);
nor I_8188 (I144914,I144513,I144897);
and I_8189 (I144931,I144832,I144914);
or I_8190 (I144948,I144736,I144931);
DFFARX1 I_8191  ( .D(I144948), .CLK(I5694_clk), .RSTB(I144445_rst), .Q(I144422) );
nand I_8192 (I144419,I144832,I144578);
DFFARX1 I_8193  ( .D(I144832), .CLK(I5694_clk), .RSTB(I144445_rst), .Q(I144410) );
not I_8194 (I145040_rst,I5701);
nand I_8195 (I145057,I127000,I127006);
and I_8196 (I145074,I145057,I126988);
DFFARX1 I_8197  ( .D(I145074), .CLK(I5694_clk), .RSTB(I145040_rst), .Q(I145091) );
nor I_8198 (I145108,I126982,I127006);
nor I_8199 (I145125,I145108,I145091);
not I_8200 (I145023,I145108);
DFFARX1 I_8201  ( .D(I127012), .CLK(I5694_clk), .RSTB(I145040_rst), .Q(I145156) );
not I_8202 (I145173,I145156);
nor I_8203 (I145190,I145108,I145173);
nand I_8204 (I145026,I145156,I145125);
DFFARX1 I_8205  ( .D(I145156), .CLK(I5694_clk), .RSTB(I145040_rst), .Q(I145008) );
nand I_8206 (I145235,I127003,I126994);
and I_8207 (I145252,I145235,I126997);
DFFARX1 I_8208  ( .D(I145252), .CLK(I5694_clk), .RSTB(I145040_rst), .Q(I145269) );
nor I_8209 (I145029,I145269,I145091);
nand I_8210 (I145020,I145269,I145190);
DFFARX1 I_8211  ( .D(I127009), .CLK(I5694_clk), .RSTB(I145040_rst), .Q(I145314) );
and I_8212 (I145331,I145314,I126985);
DFFARX1 I_8213  ( .D(I145331), .CLK(I5694_clk), .RSTB(I145040_rst), .Q(I145348) );
not I_8214 (I145011,I145348);
nand I_8215 (I145379,I145331,I145269);
and I_8216 (I145396,I145091,I145379);
DFFARX1 I_8217  ( .D(I145396), .CLK(I5694_clk), .RSTB(I145040_rst), .Q(I145002) );
DFFARX1 I_8218  ( .D(I126991), .CLK(I5694_clk), .RSTB(I145040_rst), .Q(I145427) );
nand I_8219 (I145444,I145427,I145091);
and I_8220 (I145461,I145269,I145444);
DFFARX1 I_8221  ( .D(I145461), .CLK(I5694_clk), .RSTB(I145040_rst), .Q(I145032) );
not I_8222 (I145492,I145427);
nor I_8223 (I145509,I145108,I145492);
and I_8224 (I145526,I145427,I145509);
or I_8225 (I145543,I145331,I145526);
DFFARX1 I_8226  ( .D(I145543), .CLK(I5694_clk), .RSTB(I145040_rst), .Q(I145017) );
nand I_8227 (I145014,I145427,I145173);
DFFARX1 I_8228  ( .D(I145427), .CLK(I5694_clk), .RSTB(I145040_rst), .Q(I145005) );
not I_8229 (I145635_rst,I5701);
nand I_8230 (I145652,I77170,I77161);
and I_8231 (I145669,I145652,I77179);
DFFARX1 I_8232  ( .D(I145669), .CLK(I5694_clk), .RSTB(I145635_rst), .Q(I145686) );
nor I_8233 (I145703,I77158,I77161);
nor I_8234 (I145720,I145703,I145686);
not I_8235 (I145618,I145703);
DFFARX1 I_8236  ( .D(I77167), .CLK(I5694_clk), .RSTB(I145635_rst), .Q(I145751) );
not I_8237 (I145768,I145751);
nor I_8238 (I145785,I145703,I145768);
nand I_8239 (I145621,I145751,I145720);
DFFARX1 I_8240  ( .D(I145751), .CLK(I5694_clk), .RSTB(I145635_rst), .Q(I145603) );
nand I_8241 (I145830,I77182,I77164);
and I_8242 (I145847,I145830,I77185);
DFFARX1 I_8243  ( .D(I145847), .CLK(I5694_clk), .RSTB(I145635_rst), .Q(I145864) );
nor I_8244 (I145624,I145864,I145686);
nand I_8245 (I145615,I145864,I145785);
DFFARX1 I_8246  ( .D(I77173), .CLK(I5694_clk), .RSTB(I145635_rst), .Q(I145909) );
and I_8247 (I145926,I145909,I77155);
DFFARX1 I_8248  ( .D(I145926), .CLK(I5694_clk), .RSTB(I145635_rst), .Q(I145943) );
not I_8249 (I145606,I145943);
nand I_8250 (I145974,I145926,I145864);
and I_8251 (I145991,I145686,I145974);
DFFARX1 I_8252  ( .D(I145991), .CLK(I5694_clk), .RSTB(I145635_rst), .Q(I145597) );
DFFARX1 I_8253  ( .D(I77176), .CLK(I5694_clk), .RSTB(I145635_rst), .Q(I146022) );
nand I_8254 (I146039,I146022,I145686);
and I_8255 (I146056,I145864,I146039);
DFFARX1 I_8256  ( .D(I146056), .CLK(I5694_clk), .RSTB(I145635_rst), .Q(I145627) );
not I_8257 (I146087,I146022);
nor I_8258 (I146104,I145703,I146087);
and I_8259 (I146121,I146022,I146104);
or I_8260 (I146138,I145926,I146121);
DFFARX1 I_8261  ( .D(I146138), .CLK(I5694_clk), .RSTB(I145635_rst), .Q(I145612) );
nand I_8262 (I145609,I146022,I145768);
DFFARX1 I_8263  ( .D(I146022), .CLK(I5694_clk), .RSTB(I145635_rst), .Q(I145600) );
not I_8264 (I146230_rst,I5701);
nand I_8265 (I146247,I119707,I119713);
and I_8266 (I146264,I146247,I119695);
DFFARX1 I_8267  ( .D(I146264), .CLK(I5694_clk), .RSTB(I146230_rst), .Q(I146281) );
nor I_8268 (I146298,I119689,I119713);
nor I_8269 (I146315,I146298,I146281);
not I_8270 (I146213,I146298);
DFFARX1 I_8271  ( .D(I119719), .CLK(I5694_clk), .RSTB(I146230_rst), .Q(I146346) );
not I_8272 (I146363,I146346);
nor I_8273 (I146380,I146298,I146363);
nand I_8274 (I146216,I146346,I146315);
DFFARX1 I_8275  ( .D(I146346), .CLK(I5694_clk), .RSTB(I146230_rst), .Q(I146198) );
nand I_8276 (I146425,I119710,I119701);
and I_8277 (I146442,I146425,I119704);
DFFARX1 I_8278  ( .D(I146442), .CLK(I5694_clk), .RSTB(I146230_rst), .Q(I146459) );
nor I_8279 (I146219,I146459,I146281);
nand I_8280 (I146210,I146459,I146380);
DFFARX1 I_8281  ( .D(I119716), .CLK(I5694_clk), .RSTB(I146230_rst), .Q(I146504) );
and I_8282 (I146521,I146504,I119692);
DFFARX1 I_8283  ( .D(I146521), .CLK(I5694_clk), .RSTB(I146230_rst), .Q(I146538) );
not I_8284 (I146201,I146538);
nand I_8285 (I146569,I146521,I146459);
and I_8286 (I146586,I146281,I146569);
DFFARX1 I_8287  ( .D(I146586), .CLK(I5694_clk), .RSTB(I146230_rst), .Q(I146192) );
DFFARX1 I_8288  ( .D(I119698), .CLK(I5694_clk), .RSTB(I146230_rst), .Q(I146617) );
nand I_8289 (I146634,I146617,I146281);
and I_8290 (I146651,I146459,I146634);
DFFARX1 I_8291  ( .D(I146651), .CLK(I5694_clk), .RSTB(I146230_rst), .Q(I146222) );
not I_8292 (I146682,I146617);
nor I_8293 (I146699,I146298,I146682);
and I_8294 (I146716,I146617,I146699);
or I_8295 (I146733,I146521,I146716);
DFFARX1 I_8296  ( .D(I146733), .CLK(I5694_clk), .RSTB(I146230_rst), .Q(I146207) );
nand I_8297 (I146204,I146617,I146363);
DFFARX1 I_8298  ( .D(I146617), .CLK(I5694_clk), .RSTB(I146230_rst), .Q(I146195) );
not I_8299 (I146825_rst,I5701);
nand I_8300 (I146842,I93589,I93595);
and I_8301 (I146859,I146842,I93586);
DFFARX1 I_8302  ( .D(I146859), .CLK(I5694_clk), .RSTB(I146825_rst), .Q(I146876) );
nor I_8303 (I146893,I93598,I93595);
nor I_8304 (I146910,I146893,I146876);
not I_8305 (I146808,I146893);
DFFARX1 I_8306  ( .D(I93577), .CLK(I5694_clk), .RSTB(I146825_rst), .Q(I146941) );
not I_8307 (I146958,I146941);
nor I_8308 (I146975,I146893,I146958);
nand I_8309 (I146811,I146941,I146910);
DFFARX1 I_8310  ( .D(I146941), .CLK(I5694_clk), .RSTB(I146825_rst), .Q(I146793) );
nand I_8311 (I147020,I93601,I93583);
and I_8312 (I147037,I147020,I93592);
DFFARX1 I_8313  ( .D(I147037), .CLK(I5694_clk), .RSTB(I146825_rst), .Q(I147054) );
nor I_8314 (I146814,I147054,I146876);
nand I_8315 (I146805,I147054,I146975);
DFFARX1 I_8316  ( .D(I93607), .CLK(I5694_clk), .RSTB(I146825_rst), .Q(I147099) );
and I_8317 (I147116,I147099,I93580);
DFFARX1 I_8318  ( .D(I147116), .CLK(I5694_clk), .RSTB(I146825_rst), .Q(I147133) );
not I_8319 (I146796,I147133);
nand I_8320 (I147164,I147116,I147054);
and I_8321 (I147181,I146876,I147164);
DFFARX1 I_8322  ( .D(I147181), .CLK(I5694_clk), .RSTB(I146825_rst), .Q(I146787) );
DFFARX1 I_8323  ( .D(I93604), .CLK(I5694_clk), .RSTB(I146825_rst), .Q(I147212) );
nand I_8324 (I147229,I147212,I146876);
and I_8325 (I147246,I147054,I147229);
DFFARX1 I_8326  ( .D(I147246), .CLK(I5694_clk), .RSTB(I146825_rst), .Q(I146817) );
not I_8327 (I147277,I147212);
nor I_8328 (I147294,I146893,I147277);
and I_8329 (I147311,I147212,I147294);
or I_8330 (I147328,I147116,I147311);
DFFARX1 I_8331  ( .D(I147328), .CLK(I5694_clk), .RSTB(I146825_rst), .Q(I146802) );
nand I_8332 (I146799,I147212,I146958);
DFFARX1 I_8333  ( .D(I147212), .CLK(I5694_clk), .RSTB(I146825_rst), .Q(I146790) );
not I_8334 (I147420_rst,I5701);
nand I_8335 (I147437,I134123,I134135);
and I_8336 (I147454,I147437,I134117);
DFFARX1 I_8337  ( .D(I147454), .CLK(I5694_clk), .RSTB(I147420_rst), .Q(I147471) );
nor I_8338 (I147488,I134129,I134135);
nor I_8339 (I147505,I147488,I147471);
not I_8340 (I147403,I147488);
DFFARX1 I_8341  ( .D(I134114), .CLK(I5694_clk), .RSTB(I147420_rst), .Q(I147536) );
not I_8342 (I147553,I147536);
nor I_8343 (I147570,I147488,I147553);
nand I_8344 (I147406,I147536,I147505);
DFFARX1 I_8345  ( .D(I147536), .CLK(I5694_clk), .RSTB(I147420_rst), .Q(I147388) );
nand I_8346 (I147615,I134105,I134120);
and I_8347 (I147632,I147615,I134111);
DFFARX1 I_8348  ( .D(I147632), .CLK(I5694_clk), .RSTB(I147420_rst), .Q(I147649) );
nor I_8349 (I147409,I147649,I147471);
nand I_8350 (I147400,I147649,I147570);
DFFARX1 I_8351  ( .D(I134132), .CLK(I5694_clk), .RSTB(I147420_rst), .Q(I147694) );
and I_8352 (I147711,I147694,I134126);
DFFARX1 I_8353  ( .D(I147711), .CLK(I5694_clk), .RSTB(I147420_rst), .Q(I147728) );
not I_8354 (I147391,I147728);
nand I_8355 (I147759,I147711,I147649);
and I_8356 (I147776,I147471,I147759);
DFFARX1 I_8357  ( .D(I147776), .CLK(I5694_clk), .RSTB(I147420_rst), .Q(I147382) );
DFFARX1 I_8358  ( .D(I134108), .CLK(I5694_clk), .RSTB(I147420_rst), .Q(I147807) );
nand I_8359 (I147824,I147807,I147471);
and I_8360 (I147841,I147649,I147824);
DFFARX1 I_8361  ( .D(I147841), .CLK(I5694_clk), .RSTB(I147420_rst), .Q(I147412) );
not I_8362 (I147872,I147807);
nor I_8363 (I147889,I147488,I147872);
and I_8364 (I147906,I147807,I147889);
or I_8365 (I147923,I147711,I147906);
DFFARX1 I_8366  ( .D(I147923), .CLK(I5694_clk), .RSTB(I147420_rst), .Q(I147397) );
nand I_8367 (I147394,I147807,I147553);
DFFARX1 I_8368  ( .D(I147807), .CLK(I5694_clk), .RSTB(I147420_rst), .Q(I147385) );
not I_8369 (I148015_rst,I5701);
nand I_8370 (I148032,I124348,I124354);
and I_8371 (I148049,I148032,I124336);
DFFARX1 I_8372  ( .D(I148049), .CLK(I5694_clk), .RSTB(I148015_rst), .Q(I148066) );
nor I_8373 (I148083,I124330,I124354);
nor I_8374 (I148100,I148083,I148066);
not I_8375 (I147998,I148083);
DFFARX1 I_8376  ( .D(I124360), .CLK(I5694_clk), .RSTB(I148015_rst), .Q(I148131) );
not I_8377 (I148148,I148131);
nor I_8378 (I148165,I148083,I148148);
nand I_8379 (I148001,I148131,I148100);
DFFARX1 I_8380  ( .D(I148131), .CLK(I5694_clk), .RSTB(I148015_rst), .Q(I147983) );
nand I_8381 (I148210,I124351,I124342);
and I_8382 (I148227,I148210,I124345);
DFFARX1 I_8383  ( .D(I148227), .CLK(I5694_clk), .RSTB(I148015_rst), .Q(I148244) );
nor I_8384 (I148004,I148244,I148066);
nand I_8385 (I147995,I148244,I148165);
DFFARX1 I_8386  ( .D(I124357), .CLK(I5694_clk), .RSTB(I148015_rst), .Q(I148289) );
and I_8387 (I148306,I148289,I124333);
DFFARX1 I_8388  ( .D(I148306), .CLK(I5694_clk), .RSTB(I148015_rst), .Q(I148323) );
not I_8389 (I147986,I148323);
nand I_8390 (I148354,I148306,I148244);
and I_8391 (I148371,I148066,I148354);
DFFARX1 I_8392  ( .D(I148371), .CLK(I5694_clk), .RSTB(I148015_rst), .Q(I147977) );
DFFARX1 I_8393  ( .D(I124339), .CLK(I5694_clk), .RSTB(I148015_rst), .Q(I148402) );
nand I_8394 (I148419,I148402,I148066);
and I_8395 (I148436,I148244,I148419);
DFFARX1 I_8396  ( .D(I148436), .CLK(I5694_clk), .RSTB(I148015_rst), .Q(I148007) );
not I_8397 (I148467,I148402);
nor I_8398 (I148484,I148083,I148467);
and I_8399 (I148501,I148402,I148484);
or I_8400 (I148518,I148306,I148501);
DFFARX1 I_8401  ( .D(I148518), .CLK(I5694_clk), .RSTB(I148015_rst), .Q(I147992) );
nand I_8402 (I147989,I148402,I148148);
DFFARX1 I_8403  ( .D(I148402), .CLK(I5694_clk), .RSTB(I148015_rst), .Q(I147980) );
not I_8404 (I148610_rst,I5701);
nand I_8405 (I148627,I133477,I133489);
and I_8406 (I148644,I148627,I133471);
DFFARX1 I_8407  ( .D(I148644), .CLK(I5694_clk), .RSTB(I148610_rst), .Q(I148661) );
nor I_8408 (I148678,I133483,I133489);
nor I_8409 (I148695,I148678,I148661);
not I_8410 (I148593,I148678);
DFFARX1 I_8411  ( .D(I133468), .CLK(I5694_clk), .RSTB(I148610_rst), .Q(I148726) );
not I_8412 (I148743,I148726);
nor I_8413 (I148760,I148678,I148743);
nand I_8414 (I148596,I148726,I148695);
DFFARX1 I_8415  ( .D(I148726), .CLK(I5694_clk), .RSTB(I148610_rst), .Q(I148578) );
nand I_8416 (I148805,I133459,I133474);
and I_8417 (I148822,I148805,I133465);
DFFARX1 I_8418  ( .D(I148822), .CLK(I5694_clk), .RSTB(I148610_rst), .Q(I148839) );
nor I_8419 (I148599,I148839,I148661);
nand I_8420 (I148590,I148839,I148760);
DFFARX1 I_8421  ( .D(I133486), .CLK(I5694_clk), .RSTB(I148610_rst), .Q(I148884) );
and I_8422 (I148901,I148884,I133480);
DFFARX1 I_8423  ( .D(I148901), .CLK(I5694_clk), .RSTB(I148610_rst), .Q(I148918) );
not I_8424 (I148581,I148918);
nand I_8425 (I148949,I148901,I148839);
and I_8426 (I148966,I148661,I148949);
DFFARX1 I_8427  ( .D(I148966), .CLK(I5694_clk), .RSTB(I148610_rst), .Q(I148572) );
DFFARX1 I_8428  ( .D(I133462), .CLK(I5694_clk), .RSTB(I148610_rst), .Q(I148997) );
nand I_8429 (I149014,I148997,I148661);
and I_8430 (I149031,I148839,I149014);
DFFARX1 I_8431  ( .D(I149031), .CLK(I5694_clk), .RSTB(I148610_rst), .Q(I148602) );
not I_8432 (I149062,I148997);
nor I_8433 (I149079,I148678,I149062);
and I_8434 (I149096,I148997,I149079);
or I_8435 (I149113,I148901,I149096);
DFFARX1 I_8436  ( .D(I149113), .CLK(I5694_clk), .RSTB(I148610_rst), .Q(I148587) );
nand I_8437 (I148584,I148997,I148743);
DFFARX1 I_8438  ( .D(I148997), .CLK(I5694_clk), .RSTB(I148610_rst), .Q(I148575) );
not I_8439 (I149205_rst,I5701);
nand I_8440 (I149222,I109696,I109717);
and I_8441 (I149239,I149222,I109702);
DFFARX1 I_8442  ( .D(I149239), .CLK(I5694_clk), .RSTB(I149205_rst), .Q(I149256) );
nor I_8443 (I149273,I109720,I109717);
DFFARX1 I_8444  ( .D(I109723), .CLK(I5694_clk), .RSTB(I149205_rst), .Q(I149290) );
nand I_8445 (I149307,I149290,I149273);
DFFARX1 I_8446  ( .D(I149290), .CLK(I5694_clk), .RSTB(I149205_rst), .Q(I149176) );
nand I_8447 (I149338,I109693,I109705);
and I_8448 (I149355,I149338,I109714);
DFFARX1 I_8449  ( .D(I149355), .CLK(I5694_clk), .RSTB(I149205_rst), .Q(I149372) );
not I_8450 (I149389,I149372);
nor I_8451 (I149406,I149256,I149389);
and I_8452 (I149423,I149273,I149406);
and I_8453 (I149440,I149372,I149307);
DFFARX1 I_8454  ( .D(I149440), .CLK(I5694_clk), .RSTB(I149205_rst), .Q(I149173) );
DFFARX1 I_8455  ( .D(I149372), .CLK(I5694_clk), .RSTB(I149205_rst), .Q(I149167) );
DFFARX1 I_8456  ( .D(I109708), .CLK(I5694_clk), .RSTB(I149205_rst), .Q(I149485) );
and I_8457 (I149502,I149485,I109711);
nand I_8458 (I149519,I149502,I149372);
nor I_8459 (I149194,I149502,I149273);
not I_8460 (I149550,I149502);
nor I_8461 (I149567,I149256,I149550);
nand I_8462 (I149185,I149290,I149567);
nand I_8463 (I149179,I149372,I149550);
or I_8464 (I149612,I149502,I149423);
DFFARX1 I_8465  ( .D(I149612), .CLK(I5694_clk), .RSTB(I149205_rst), .Q(I149182) );
DFFARX1 I_8466  ( .D(I109699), .CLK(I5694_clk), .RSTB(I149205_rst), .Q(I149643) );
and I_8467 (I149660,I149643,I149519);
DFFARX1 I_8468  ( .D(I149660), .CLK(I5694_clk), .RSTB(I149205_rst), .Q(I149197) );
nor I_8469 (I149691,I149643,I149256);
nand I_8470 (I149191,I149502,I149691);
not I_8471 (I149188,I149643);
DFFARX1 I_8472  ( .D(I149643), .CLK(I5694_clk), .RSTB(I149205_rst), .Q(I149736) );
and I_8473 (I149170,I149643,I149736);
not I_8474 (I149800_rst,I5701);
nand I_8475 (I149817,I127663,I127675);
and I_8476 (I149834,I149817,I127666);
DFFARX1 I_8477  ( .D(I149834), .CLK(I5694_clk), .RSTB(I149800_rst), .Q(I149851) );
nor I_8478 (I149868,I127660,I127675);
DFFARX1 I_8479  ( .D(I127651), .CLK(I5694_clk), .RSTB(I149800_rst), .Q(I149885) );
nand I_8480 (I149902,I149885,I149868);
DFFARX1 I_8481  ( .D(I149885), .CLK(I5694_clk), .RSTB(I149800_rst), .Q(I149771) );
nand I_8482 (I149933,I127657,I127648);
and I_8483 (I149950,I149933,I127654);
DFFARX1 I_8484  ( .D(I149950), .CLK(I5694_clk), .RSTB(I149800_rst), .Q(I149967) );
not I_8485 (I149984,I149967);
nor I_8486 (I150001,I149851,I149984);
and I_8487 (I150018,I149868,I150001);
and I_8488 (I150035,I149967,I149902);
DFFARX1 I_8489  ( .D(I150035), .CLK(I5694_clk), .RSTB(I149800_rst), .Q(I149768) );
DFFARX1 I_8490  ( .D(I149967), .CLK(I5694_clk), .RSTB(I149800_rst), .Q(I149762) );
DFFARX1 I_8491  ( .D(I127669), .CLK(I5694_clk), .RSTB(I149800_rst), .Q(I150080) );
and I_8492 (I150097,I150080,I127645);
nand I_8493 (I150114,I150097,I149967);
nor I_8494 (I149789,I150097,I149868);
not I_8495 (I150145,I150097);
nor I_8496 (I150162,I149851,I150145);
nand I_8497 (I149780,I149885,I150162);
nand I_8498 (I149774,I149967,I150145);
or I_8499 (I150207,I150097,I150018);
DFFARX1 I_8500  ( .D(I150207), .CLK(I5694_clk), .RSTB(I149800_rst), .Q(I149777) );
DFFARX1 I_8501  ( .D(I127672), .CLK(I5694_clk), .RSTB(I149800_rst), .Q(I150238) );
and I_8502 (I150255,I150238,I150114);
DFFARX1 I_8503  ( .D(I150255), .CLK(I5694_clk), .RSTB(I149800_rst), .Q(I149792) );
nor I_8504 (I150286,I150238,I149851);
nand I_8505 (I149786,I150097,I150286);
not I_8506 (I149783,I150238);
DFFARX1 I_8507  ( .D(I150238), .CLK(I5694_clk), .RSTB(I149800_rst), .Q(I150331) );
and I_8508 (I149765,I150238,I150331);
not I_8509 (I150395_rst,I5701);
nand I_8510 (I150412,I147397,I147382);
and I_8511 (I150429,I150412,I147388);
DFFARX1 I_8512  ( .D(I150429), .CLK(I5694_clk), .RSTB(I150395_rst), .Q(I150446) );
nor I_8513 (I150463,I147391,I147382);
DFFARX1 I_8514  ( .D(I147403), .CLK(I5694_clk), .RSTB(I150395_rst), .Q(I150480) );
nand I_8515 (I150497,I150480,I150463);
DFFARX1 I_8516  ( .D(I150480), .CLK(I5694_clk), .RSTB(I150395_rst), .Q(I150366) );
nand I_8517 (I150528,I147394,I147385);
and I_8518 (I150545,I150528,I147412);
DFFARX1 I_8519  ( .D(I150545), .CLK(I5694_clk), .RSTB(I150395_rst), .Q(I150562) );
not I_8520 (I150579,I150562);
nor I_8521 (I150596,I150446,I150579);
and I_8522 (I150613,I150463,I150596);
and I_8523 (I150630,I150562,I150497);
DFFARX1 I_8524  ( .D(I150630), .CLK(I5694_clk), .RSTB(I150395_rst), .Q(I150363) );
DFFARX1 I_8525  ( .D(I150562), .CLK(I5694_clk), .RSTB(I150395_rst), .Q(I150357) );
DFFARX1 I_8526  ( .D(I147400), .CLK(I5694_clk), .RSTB(I150395_rst), .Q(I150675) );
and I_8527 (I150692,I150675,I147406);
nand I_8528 (I150709,I150692,I150562);
nor I_8529 (I150384,I150692,I150463);
not I_8530 (I150740,I150692);
nor I_8531 (I150757,I150446,I150740);
nand I_8532 (I150375,I150480,I150757);
nand I_8533 (I150369,I150562,I150740);
or I_8534 (I150802,I150692,I150613);
DFFARX1 I_8535  ( .D(I150802), .CLK(I5694_clk), .RSTB(I150395_rst), .Q(I150372) );
DFFARX1 I_8536  ( .D(I147409), .CLK(I5694_clk), .RSTB(I150395_rst), .Q(I150833) );
and I_8537 (I150850,I150833,I150709);
DFFARX1 I_8538  ( .D(I150850), .CLK(I5694_clk), .RSTB(I150395_rst), .Q(I150387) );
nor I_8539 (I150881,I150833,I150446);
nand I_8540 (I150381,I150692,I150881);
not I_8541 (I150378,I150833);
DFFARX1 I_8542  ( .D(I150833), .CLK(I5694_clk), .RSTB(I150395_rst), .Q(I150926) );
and I_8543 (I150360,I150833,I150926);
not I_8544 (I150990_rst,I5701);
nand I_8545 (I151007,I142669,I142657);
and I_8546 (I151024,I151007,I142645);
DFFARX1 I_8547  ( .D(I151024), .CLK(I5694_clk), .RSTB(I150990_rst), .Q(I151041) );
nor I_8548 (I151058,I142642,I142657);
DFFARX1 I_8549  ( .D(I142654), .CLK(I5694_clk), .RSTB(I150990_rst), .Q(I151075) );
nand I_8550 (I151092,I151075,I151058);
DFFARX1 I_8551  ( .D(I151075), .CLK(I5694_clk), .RSTB(I150990_rst), .Q(I150961) );
nand I_8552 (I151123,I142651,I142648);
and I_8553 (I151140,I151123,I142666);
DFFARX1 I_8554  ( .D(I151140), .CLK(I5694_clk), .RSTB(I150990_rst), .Q(I151157) );
not I_8555 (I151174,I151157);
nor I_8556 (I151191,I151041,I151174);
and I_8557 (I151208,I151058,I151191);
and I_8558 (I151225,I151157,I151092);
DFFARX1 I_8559  ( .D(I151225), .CLK(I5694_clk), .RSTB(I150990_rst), .Q(I150958) );
DFFARX1 I_8560  ( .D(I151157), .CLK(I5694_clk), .RSTB(I150990_rst), .Q(I150952) );
DFFARX1 I_8561  ( .D(I142663), .CLK(I5694_clk), .RSTB(I150990_rst), .Q(I151270) );
and I_8562 (I151287,I151270,I142639);
nand I_8563 (I151304,I151287,I151157);
nor I_8564 (I150979,I151287,I151058);
not I_8565 (I151335,I151287);
nor I_8566 (I151352,I151041,I151335);
nand I_8567 (I150970,I151075,I151352);
nand I_8568 (I150964,I151157,I151335);
or I_8569 (I151397,I151287,I151208);
DFFARX1 I_8570  ( .D(I151397), .CLK(I5694_clk), .RSTB(I150990_rst), .Q(I150967) );
DFFARX1 I_8571  ( .D(I142660), .CLK(I5694_clk), .RSTB(I150990_rst), .Q(I151428) );
and I_8572 (I151445,I151428,I151304);
DFFARX1 I_8573  ( .D(I151445), .CLK(I5694_clk), .RSTB(I150990_rst), .Q(I150982) );
nor I_8574 (I151476,I151428,I151041);
nand I_8575 (I150976,I151287,I151476);
not I_8576 (I150973,I151428);
DFFARX1 I_8577  ( .D(I151428), .CLK(I5694_clk), .RSTB(I150990_rst), .Q(I151521) );
and I_8578 (I150955,I151428,I151521);
not I_8579 (I151585_rst,I5701);
nand I_8580 (I151602,I114891,I114876);
and I_8581 (I151619,I151602,I11488_rst8);
DFFARX1 I_8582  ( .D(I151619), .CLK(I5694_clk), .RSTB(I151585_rst), .Q(I151636) );
nor I_8583 (I151653,I114879,I114876);
DFFARX1 I_8584  ( .D(I114870), .CLK(I5694_clk), .RSTB(I151585_rst), .Q(I151670) );
nand I_8585 (I151687,I151670,I151653);
DFFARX1 I_8586  ( .D(I151670), .CLK(I5694_clk), .RSTB(I151585_rst), .Q(I151556) );
nand I_8587 (I151718,I114861,I11488_rst5);
and I_8588 (I151735,I151718,I114864);
DFFARX1 I_8589  ( .D(I151735), .CLK(I5694_clk), .RSTB(I151585_rst), .Q(I151752) );
not I_8590 (I151769,I151752);
nor I_8591 (I151786,I151636,I151769);
and I_8592 (I151803,I151653,I151786);
and I_8593 (I151820,I151752,I151687);
DFFARX1 I_8594  ( .D(I151820), .CLK(I5694_clk), .RSTB(I151585_rst), .Q(I151553) );
DFFARX1 I_8595  ( .D(I151752), .CLK(I5694_clk), .RSTB(I151585_rst), .Q(I151547) );
DFFARX1 I_8596  ( .D(I11488_rst2), .CLK(I5694_clk), .RSTB(I151585_rst), .Q(I151865) );
and I_8597 (I151882,I151865,I114867);
nand I_8598 (I151899,I151882,I151752);
nor I_8599 (I151574,I151882,I151653);
not I_8600 (I151930,I151882);
nor I_8601 (I151947,I151636,I151930);
nand I_8602 (I151565,I151670,I151947);
nand I_8603 (I151559,I151752,I151930);
or I_8604 (I151992,I151882,I151803);
DFFARX1 I_8605  ( .D(I151992), .CLK(I5694_clk), .RSTB(I151585_rst), .Q(I151562) );
DFFARX1 I_8606  ( .D(I114873), .CLK(I5694_clk), .RSTB(I151585_rst), .Q(I152023) );
and I_8607 (I152040,I152023,I151899);
DFFARX1 I_8608  ( .D(I152040), .CLK(I5694_clk), .RSTB(I151585_rst), .Q(I151577) );
nor I_8609 (I152071,I152023,I151636);
nand I_8610 (I151571,I151882,I152071);
not I_8611 (I151568,I152023);
DFFARX1 I_8612  ( .D(I152023), .CLK(I5694_clk), .RSTB(I151585_rst), .Q(I152116) );
and I_8613 (I151550,I152023,I152116);
not I_8614 (I152180_rst,I5701);
nand I_8615 (I152197,I106439,I106415);
and I_8616 (I152214,I152197,I106424);
DFFARX1 I_8617  ( .D(I152214), .CLK(I5694_clk), .RSTB(I152180_rst), .Q(I152231) );
nor I_8618 (I152248,I106418,I106415);
DFFARX1 I_8619  ( .D(I106433), .CLK(I5694_clk), .RSTB(I152180_rst), .Q(I152265) );
nand I_8620 (I152282,I152265,I152248);
DFFARX1 I_8621  ( .D(I152265), .CLK(I5694_clk), .RSTB(I152180_rst), .Q(I152151) );
nand I_8622 (I152313,I106427,I106442);
and I_8623 (I152330,I152313,I106421);
DFFARX1 I_8624  ( .D(I152330), .CLK(I5694_clk), .RSTB(I152180_rst), .Q(I152347) );
not I_8625 (I152364,I152347);
nor I_8626 (I152381,I152231,I152364);
and I_8627 (I152398,I152248,I152381);
and I_8628 (I152415,I152347,I152282);
DFFARX1 I_8629  ( .D(I152415), .CLK(I5694_clk), .RSTB(I152180_rst), .Q(I152148) );
DFFARX1 I_8630  ( .D(I152347), .CLK(I5694_clk), .RSTB(I152180_rst), .Q(I152142) );
DFFARX1 I_8631  ( .D(I106412), .CLK(I5694_clk), .RSTB(I152180_rst), .Q(I152460) );
and I_8632 (I152477,I152460,I106430);
nand I_8633 (I152494,I152477,I152347);
nor I_8634 (I152169,I152477,I152248);
not I_8635 (I152525,I152477);
nor I_8636 (I152542,I152231,I152525);
nand I_8637 (I152160,I152265,I152542);
nand I_8638 (I152154,I152347,I152525);
or I_8639 (I152587,I152477,I152398);
DFFARX1 I_8640  ( .D(I152587), .CLK(I5694_clk), .RSTB(I152180_rst), .Q(I152157) );
DFFARX1 I_8641  ( .D(I106436), .CLK(I5694_clk), .RSTB(I152180_rst), .Q(I152618) );
and I_8642 (I152635,I152618,I152494);
DFFARX1 I_8643  ( .D(I152635), .CLK(I5694_clk), .RSTB(I152180_rst), .Q(I152172) );
nor I_8644 (I152666,I152618,I152231);
nand I_8645 (I152166,I152477,I152666);
not I_8646 (I152163,I152618);
DFFARX1 I_8647  ( .D(I152618), .CLK(I5694_clk), .RSTB(I152180_rst), .Q(I152711) );
and I_8648 (I152145,I152618,I152711);
not I_8649 (I152775_rst,I5701);
nand I_8650 (I152792,I134769,I134781);
and I_8651 (I152809,I152792,I134772);
DFFARX1 I_8652  ( .D(I152809), .CLK(I5694_clk), .RSTB(I152775_rst), .Q(I152826) );
nor I_8653 (I152843,I134766,I134781);
DFFARX1 I_8654  ( .D(I134757), .CLK(I5694_clk), .RSTB(I152775_rst), .Q(I152860) );
nand I_8655 (I152877,I152860,I152843);
DFFARX1 I_8656  ( .D(I152860), .CLK(I5694_clk), .RSTB(I152775_rst), .Q(I152746) );
nand I_8657 (I152908,I134763,I134754);
and I_8658 (I152925,I152908,I134760);
DFFARX1 I_8659  ( .D(I152925), .CLK(I5694_clk), .RSTB(I152775_rst), .Q(I152942) );
not I_8660 (I152959,I152942);
nor I_8661 (I152976,I152826,I152959);
and I_8662 (I152993,I152843,I152976);
and I_8663 (I153010,I152942,I152877);
DFFARX1 I_8664  ( .D(I153010), .CLK(I5694_clk), .RSTB(I152775_rst), .Q(I152743) );
DFFARX1 I_8665  ( .D(I152942), .CLK(I5694_clk), .RSTB(I152775_rst), .Q(I152737) );
DFFARX1 I_8666  ( .D(I134775), .CLK(I5694_clk), .RSTB(I152775_rst), .Q(I153055) );
and I_8667 (I153072,I153055,I134751);
nand I_8668 (I153089,I153072,I152942);
nor I_8669 (I152764,I153072,I152843);
not I_8670 (I153120,I153072);
nor I_8671 (I153137,I152826,I153120);
nand I_8672 (I152755,I152860,I153137);
nand I_8673 (I152749,I152942,I153120);
or I_8674 (I153182,I153072,I152993);
DFFARX1 I_8675  ( .D(I153182), .CLK(I5694_clk), .RSTB(I152775_rst), .Q(I152752) );
DFFARX1 I_8676  ( .D(I134778), .CLK(I5694_clk), .RSTB(I152775_rst), .Q(I153213) );
and I_8677 (I153230,I153213,I153089);
DFFARX1 I_8678  ( .D(I153230), .CLK(I5694_clk), .RSTB(I152775_rst), .Q(I152767) );
nor I_8679 (I153261,I153213,I152826);
nand I_8680 (I152761,I153072,I153261);
not I_8681 (I152758,I153213);
DFFARX1 I_8682  ( .D(I153213), .CLK(I5694_clk), .RSTB(I152775_rst), .Q(I15330_rst6) );
and I_8683 (I152740,I153213,I15330_rst6);
not I_8684 (I153370_rst,I5701);
not I_8685 (I153387,I103834);
nor I_8686 (I153404,I103852,I103831);
nand I_8687 (I153421,I153404,I103849);
nor I_8688 (I153438,I153387,I103852);
nand I_8689 (I153455,I153438,I103843);
not I_8690 (I153472,I103852);
not I_8691 (I153489,I153472);
not I_8692 (I153506,I103846);
nor I_8693 (I153523,I153506,I103840);
and I_8694 (I153540,I153523,I103837);
or I_8695 (I153557,I153540,I103828);
DFFARX1 I_8696  ( .D(I153557), .CLK(I5694_clk), .RSTB(I153370_rst), .Q(I153574) );
nand I_8697 (I153591,I153387,I103846);
or I_8698 (I153359,I153591,I153574);
not I_8699 (I153622,I153591);
nor I_8700 (I153639,I153574,I153622);
and I_8701 (I153656,I153472,I153639);
nand I_8702 (I153332,I153591,I153489);
DFFARX1 I_8703  ( .D(I103858), .CLK(I5694_clk), .RSTB(I153370_rst), .Q(I153687) );
or I_8704 (I153353,I153687,I153574);
nor I_8705 (I153718,I153687,I153455);
nor I_8706 (I153735,I153687,I153489);
nand I_8707 (I153338,I153421,I153735);
or I_8708 (I153766,I153687,I153656);
DFFARX1 I_8709  ( .D(I153766), .CLK(I5694_clk), .RSTB(I153370_rst), .Q(I153335) );
not I_8710 (I153341,I153687);
DFFARX1 I_8711  ( .D(I103855), .CLK(I5694_clk), .RSTB(I153370_rst), .Q(I153811) );
not I_8712 (I153828,I153811);
nor I_8713 (I153845,I153828,I153421);
DFFARX1 I_8714  ( .D(I153845), .CLK(I5694_clk), .RSTB(I153370_rst), .Q(I153347) );
nor I_8715 (I153362,I153687,I153828);
nor I_8716 (I153350,I153828,I153591);
not I_8717 (I153904,I153828);
and I_8718 (I153921,I153455,I153904);
nor I_8719 (I153356,I153591,I153921);
nand I_8720 (I153344,I153828,I153718);
not I_8721 (I153999_rst,I5701);
not I_8722 (I154016,I125674);
nor I_8723 (I154033,I125680,I125659);
nand I_8724 (I154050,I154033,I125665);
nor I_8725 (I154067,I154016,I125680);
nand I_8726 (I154084,I154067,I125671);
not I_8727 (I154101,I125680);
not I_8728 (I154118,I154101);
not I_8729 (I154135,I125668);
nor I_8730 (I154152,I154135,I125686);
and I_8731 (I154169,I154152,I125677);
or I_8732 (I154186,I154169,I125656);
DFFARX1 I_8733  ( .D(I154186), .CLK(I5694_clk), .RSTB(I153999_rst), .Q(I154203) );
nand I_8734 (I154220,I154016,I125668);
or I_8735 (I153988,I154220,I154203);
not I_8736 (I154251,I154220);
nor I_8737 (I154268,I154203,I154251);
and I_8738 (I154285,I154101,I154268);
nand I_8739 (I153961,I154220,I154118);
DFFARX1 I_8740  ( .D(I125683), .CLK(I5694_clk), .RSTB(I153999_rst), .Q(I154316) );
or I_8741 (I153982,I154316,I154203);
nor I_8742 (I154347,I154316,I154084);
nor I_8743 (I154364,I154316,I154118);
nand I_8744 (I153967,I154050,I154364);
or I_8745 (I154395,I154316,I154285);
DFFARX1 I_8746  ( .D(I154395), .CLK(I5694_clk), .RSTB(I153999_rst), .Q(I153964) );
not I_8747 (I153970,I154316);
DFFARX1 I_8748  ( .D(I125662), .CLK(I5694_clk), .RSTB(I153999_rst), .Q(I154440) );
not I_8749 (I154457,I154440);
nor I_8750 (I154474,I154457,I154050);
DFFARX1 I_8751  ( .D(I154474), .CLK(I5694_clk), .RSTB(I153999_rst), .Q(I153976) );
nor I_8752 (I153991,I154316,I154457);
nor I_8753 (I153979,I154457,I154220);
not I_8754 (I154533,I154457);
and I_8755 (I154550,I154084,I154533);
nor I_8756 (I153985,I154220,I154550);
nand I_8757 (I153973,I154457,I154347);
not I_8758 (I154628_rst,I5701);
not I_8759 (I154645,I135415);
nor I_8760 (I154662,I135424,I135427);
nand I_8761 (I154679,I154662,I135412);
nor I_8762 (I154696,I154645,I135424);
nand I_8763 (I154713,I154696,I135409);
not I_8764 (I154730,I135424);
not I_8765 (I154747,I154730);
not I_8766 (I154764,I135397);
nor I_8767 (I154781,I154764,I135403);
and I_8768 (I154798,I154781,I135400);
or I_8769 (I154815,I154798,I135421);
DFFARX1 I_8770  ( .D(I154815), .CLK(I5694_clk), .RSTB(I154628_rst), .Q(I154832) );
nand I_8771 (I154849,I154645,I135397);
or I_8772 (I154617,I154849,I154832);
not I_8773 (I154880,I154849);
nor I_8774 (I154897,I154832,I154880);
and I_8775 (I154914,I154730,I154897);
nand I_8776 (I154590,I154849,I154747);
DFFARX1 I_8777  ( .D(I135406), .CLK(I5694_clk), .RSTB(I154628_rst), .Q(I154945) );
or I_8778 (I154611,I154945,I154832);
nor I_8779 (I154976,I154945,I154713);
nor I_8780 (I154993,I154945,I154747);
nand I_8781 (I154596,I154679,I154993);
or I_8782 (I155024,I154945,I154914);
DFFARX1 I_8783  ( .D(I155024), .CLK(I5694_clk), .RSTB(I154628_rst), .Q(I154593) );
not I_8784 (I154599,I154945);
DFFARX1 I_8785  ( .D(I135418), .CLK(I5694_clk), .RSTB(I154628_rst), .Q(I155069) );
not I_8786 (I155086,I155069);
nor I_8787 (I155103,I155086,I154679);
DFFARX1 I_8788  ( .D(I155103), .CLK(I5694_clk), .RSTB(I154628_rst), .Q(I154605) );
nor I_8789 (I154620,I154945,I155086);
nor I_8790 (I154608,I155086,I154849);
not I_8791 (I155162,I155086);
and I_8792 (I155179,I154713,I155162);
nor I_8793 (I154614,I154849,I155179);
nand I_8794 (I154602,I155086,I154976);
not I_8795 (I155257_rst,I5701);
not I_8796 (I155274,I138521);
nor I_8797 (I155291,I138494,I138512);
nand I_8798 (I155308,I155291,I138497);
nor I_8799 (I155325,I155274,I138494);
nand I_8800 (I155342,I155325,I138515);
not I_8801 (I155359,I138494);
not I_8802 (I155376,I155359);
not I_8803 (I155393,I138491);
nor I_8804 (I155410,I155393,I138518);
and I_8805 (I155427,I155410,I138509);
or I_8806 (I155444,I155427,I138500);
DFFARX1 I_8807  ( .D(I155444), .CLK(I5694_clk), .RSTB(I155257_rst), .Q(I155461) );
nand I_8808 (I155478,I155274,I138491);
or I_8809 (I155246,I155478,I155461);
not I_8810 (I155509,I155478);
nor I_8811 (I155526,I155461,I155509);
and I_8812 (I155543,I155359,I155526);
nand I_8813 (I155219,I155478,I155376);
DFFARX1 I_8814  ( .D(I138503), .CLK(I5694_clk), .RSTB(I155257_rst), .Q(I155574) );
or I_8815 (I155240,I155574,I155461);
nor I_8816 (I155605,I155574,I155342);
nor I_8817 (I155622,I155574,I155376);
nand I_8818 (I155225,I155308,I155622);
or I_8819 (I155653,I155574,I155543);
DFFARX1 I_8820  ( .D(I155653), .CLK(I5694_clk), .RSTB(I155257_rst), .Q(I155222) );
not I_8821 (I155228,I155574);
DFFARX1 I_8822  ( .D(I138506), .CLK(I5694_clk), .RSTB(I155257_rst), .Q(I155698) );
not I_8823 (I155715,I155698);
nor I_8824 (I155732,I155715,I155308);
DFFARX1 I_8825  ( .D(I155732), .CLK(I5694_clk), .RSTB(I155257_rst), .Q(I155234) );
nor I_8826 (I155249,I155574,I155715);
nor I_8827 (I155237,I155715,I155478);
not I_8828 (I155791,I155715);
and I_8829 (I155808,I155342,I155791);
nor I_8830 (I155243,I155478,I155808);
nand I_8831 (I155231,I155715,I155605);
not I_8832 (I155886_rst,I5701);
not I_8833 (I155903,I101250);
nor I_8834 (I155920,I101268,I101247);
nand I_8835 (I155937,I155920,I101265);
nor I_8836 (I155954,I155903,I101268);
nand I_8837 (I155971,I155954,I101259);
not I_8838 (I155988,I101268);
not I_8839 (I156005,I155988);
not I_8840 (I156022,I101262);
nor I_8841 (I156039,I156022,I101256);
and I_8842 (I156056,I156039,I101253);
or I_8843 (I156073,I156056,I101244);
DFFARX1 I_8844  ( .D(I156073), .CLK(I5694_clk), .RSTB(I155886_rst), .Q(I156090) );
nand I_8845 (I156107,I155903,I101262);
or I_8846 (I155875,I156107,I156090);
not I_8847 (I156138,I156107);
nor I_8848 (I156155,I156090,I156138);
and I_8849 (I156172,I155988,I156155);
nand I_8850 (I155848,I156107,I156005);
DFFARX1 I_8851  ( .D(I101274), .CLK(I5694_clk), .RSTB(I155886_rst), .Q(I156203) );
or I_8852 (I155869,I156203,I156090);
nor I_8853 (I156234,I156203,I155971);
nor I_8854 (I156251,I156203,I156005);
nand I_8855 (I155854,I155937,I156251);
or I_8856 (I156282,I156203,I156172);
DFFARX1 I_8857  ( .D(I156282), .CLK(I5694_clk), .RSTB(I155886_rst), .Q(I155851) );
not I_8858 (I155857,I156203);
DFFARX1 I_8859  ( .D(I101271), .CLK(I5694_clk), .RSTB(I155886_rst), .Q(I156327) );
not I_8860 (I156344,I156327);
nor I_8861 (I156361,I156344,I155937);
DFFARX1 I_8862  ( .D(I156361), .CLK(I5694_clk), .RSTB(I155886_rst), .Q(I155863) );
nor I_8863 (I155878,I156203,I156344);
nor I_8864 (I155866,I156344,I156107);
not I_8865 (I156420,I156344);
and I_8866 (I156437,I155971,I156420);
nor I_8867 (I155872,I156107,I156437);
nand I_8868 (I155860,I156344,I156234);
not I_8869 (I156515_rst,I5701);
not I_8870 (I156532,I142079);
nor I_8871 (I156549,I142064,I142085);
nand I_8872 (I156566,I156549,I142073);
nor I_8873 (I156583,I156532,I142064);
nand I_8874 (I156600,I156583,I142061);
not I_8875 (I156617,I142064);
not I_8876 (I156634,I156617);
not I_8877 (I156651,I142088);
nor I_8878 (I156668,I156651,I142076);
and I_8879 (I156685,I156668,I142070);
or I_8880 (I156702,I156685,I142067);
DFFARX1 I_8881  ( .D(I156702), .CLK(I5694_clk), .RSTB(I156515_rst), .Q(I156719) );
nand I_8882 (I156736,I156532,I142088);
or I_8883 (I156504,I156736,I156719);
not I_8884 (I156767,I156736);
nor I_8885 (I156784,I156719,I156767);
and I_8886 (I156801,I156617,I156784);
nand I_8887 (I156477,I156736,I156634);
DFFARX1 I_8888  ( .D(I142091), .CLK(I5694_clk), .RSTB(I156515_rst), .Q(I156832) );
or I_8889 (I156498,I156832,I156719);
nor I_8890 (I156863,I156832,I156600);
nor I_8891 (I156880,I156832,I156634);
nand I_8892 (I156483,I156566,I156880);
or I_8893 (I156911,I156832,I156801);
DFFARX1 I_8894  ( .D(I156911), .CLK(I5694_clk), .RSTB(I156515_rst), .Q(I156480) );
not I_8895 (I156486,I156832);
DFFARX1 I_8896  ( .D(I142082), .CLK(I5694_clk), .RSTB(I156515_rst), .Q(I156956) );
not I_8897 (I156973,I156956);
nor I_8898 (I156990,I156973,I156566);
DFFARX1 I_8899  ( .D(I156990), .CLK(I5694_clk), .RSTB(I156515_rst), .Q(I156492) );
nor I_8900 (I156507,I156832,I156973);
nor I_8901 (I156495,I156973,I156736);
not I_8902 (I157049,I156973);
and I_8903 (I157066,I156600,I157049);
nor I_8904 (I156501,I156736,I157066);
nand I_8905 (I156489,I156973,I156863);
not I_8906 (I157144_rst,I5701);
not I_8907 (I157161,I100604);
nor I_8908 (I157178,I100622,I100601);
nand I_8909 (I157195,I157178,I100619);
nor I_8910 (I157212,I157161,I100622);
nand I_8911 (I157229,I157212,I100613);
not I_8912 (I157246,I100622);
not I_8913 (I157263,I157246);
not I_8914 (I157280,I100616);
nor I_8915 (I157297,I157280,I100610);
and I_8916 (I157314,I157297,I100607);
or I_8917 (I157331,I157314,I100598);
DFFARX1 I_8918  ( .D(I157331), .CLK(I5694_clk), .RSTB(I157144_rst), .Q(I157348) );
nand I_8919 (I157365,I157161,I100616);
or I_8920 (I157133,I157365,I157348);
not I_8921 (I157396,I157365);
nor I_8922 (I157413,I157348,I157396);
and I_8923 (I157430,I157246,I157413);
nand I_8924 (I157106,I157365,I157263);
DFFARX1 I_8925  ( .D(I100628), .CLK(I5694_clk), .RSTB(I157144_rst), .Q(I157461) );
or I_8926 (I157127,I157461,I157348);
nor I_8927 (I157492,I157461,I157229);
nor I_8928 (I157509,I157461,I157263);
nand I_8929 (I157112,I157195,I157509);
or I_8930 (I157540,I157461,I157430);
DFFARX1 I_8931  ( .D(I157540), .CLK(I5694_clk), .RSTB(I157144_rst), .Q(I157109) );
not I_8932 (I157115,I157461);
DFFARX1 I_8933  ( .D(I100625), .CLK(I5694_clk), .RSTB(I157144_rst), .Q(I157585) );
not I_8934 (I157602,I157585);
nor I_8935 (I157619,I157602,I157195);
DFFARX1 I_8936  ( .D(I157619), .CLK(I5694_clk), .RSTB(I157144_rst), .Q(I157121) );
nor I_8937 (I157136,I157461,I157602);
nor I_8938 (I157124,I157602,I157365);
not I_8939 (I157678,I157602);
and I_8940 (I157695,I157229,I157678);
nor I_8941 (I157130,I157365,I157695);
nand I_8942 (I157118,I157602,I157492);
not I_8943 (I157773_rst,I5701);
not I_8944 (I157790,I139677);
nor I_8945 (I157807,I139650,I139668);
nand I_8946 (I157824,I157807,I139653);
nor I_8947 (I157841,I157790,I139650);
nand I_8948 (I157858,I157841,I139671);
not I_8949 (I157875,I139650);
not I_8950 (I157892,I157875);
not I_8951 (I157909,I139647);
nor I_8952 (I157926,I157909,I139674);
and I_8953 (I157943,I157926,I139665);
or I_8954 (I157960,I157943,I139656);
DFFARX1 I_8955  ( .D(I157960), .CLK(I5694_clk), .RSTB(I157773_rst), .Q(I157977) );
nand I_8956 (I157994,I157790,I139647);
or I_8957 (I157762,I157994,I157977);
not I_8958 (I158025,I157994);
nor I_8959 (I158042,I157977,I158025);
and I_8960 (I158059,I157875,I158042);
nand I_8961 (I157735,I157994,I157892);
DFFARX1 I_8962  ( .D(I139659), .CLK(I5694_clk), .RSTB(I157773_rst), .Q(I158090) );
or I_8963 (I157756,I158090,I157977);
nor I_8964 (I158121,I158090,I157858);
nor I_8965 (I158138,I158090,I157892);
nand I_8966 (I157741,I157824,I158138);
or I_8967 (I158169,I158090,I158059);
DFFARX1 I_8968  ( .D(I158169), .CLK(I5694_clk), .RSTB(I157773_rst), .Q(I157738) );
not I_8969 (I157744,I158090);
DFFARX1 I_8970  ( .D(I139662), .CLK(I5694_clk), .RSTB(I157773_rst), .Q(I158214) );
not I_8971 (I158231,I158214);
nor I_8972 (I158248,I158231,I157824);
DFFARX1 I_8973  ( .D(I158248), .CLK(I5694_clk), .RSTB(I157773_rst), .Q(I157750) );
nor I_8974 (I157765,I158090,I158231);
nor I_8975 (I157753,I158231,I157994);
not I_8976 (I158307,I158231);
and I_8977 (I158324,I157858,I158307);
nor I_8978 (I157759,I157994,I158324);
nand I_8979 (I157747,I158231,I158121);
not I_8980 (I158402_rst,I5701);
not I_8981 (I158419,I131539);
nor I_8982 (I158436,I131548,I131551);
nand I_8983 (I158453,I158436,I131536);
nor I_8984 (I158470,I158419,I131548);
nand I_8985 (I158487,I158470,I131533);
not I_8986 (I158504,I131548);
not I_8987 (I158521,I158504);
not I_8988 (I158538,I131521);
nor I_8989 (I158555,I158538,I131527);
and I_8990 (I158572,I158555,I131524);
or I_8991 (I158589,I158572,I131545);
DFFARX1 I_8992  ( .D(I158589), .CLK(I5694_clk), .RSTB(I158402_rst), .Q(I158606) );
nand I_8993 (I158623,I158419,I131521);
or I_8994 (I158391,I158623,I158606);
not I_8995 (I158654,I158623);
nor I_8996 (I158671,I158606,I158654);
and I_8997 (I158688,I158504,I158671);
nand I_8998 (I158364,I158623,I158521);
DFFARX1 I_8999  ( .D(I131530), .CLK(I5694_clk), .RSTB(I158402_rst), .Q(I158719) );
or I_9000 (I158385,I158719,I158606);
nor I_9001 (I158750,I158719,I158487);
nor I_9002 (I158767,I158719,I158521);
nand I_9003 (I158370,I158453,I158767);
or I_9004 (I158798,I158719,I158688);
DFFARX1 I_9005  ( .D(I158798), .CLK(I5694_clk), .RSTB(I158402_rst), .Q(I158367) );
not I_9006 (I158373,I158719);
DFFARX1 I_9007  ( .D(I131542), .CLK(I5694_clk), .RSTB(I158402_rst), .Q(I158843) );
not I_9008 (I158860,I158843);
nor I_9009 (I158877,I158860,I158453);
DFFARX1 I_9010  ( .D(I158877), .CLK(I5694_clk), .RSTB(I158402_rst), .Q(I158379) );
nor I_9011 (I158394,I158719,I158860);
nor I_9012 (I158382,I158860,I158623);
not I_9013 (I158936,I158860);
and I_9014 (I158953,I158487,I158936);
nor I_9015 (I158388,I158623,I158953);
nand I_9016 (I158376,I158860,I158750);
not I_9017 (I159031_rst,I5701);
nand I_9018 (I159048,I114275,I114272);
and I_9019 (I159065,I159048,I114284);
DFFARX1 I_9020  ( .D(I159065), .CLK(I5694_clk), .RSTB(I159031_rst), .Q(I159082) );
not I_9021 (I159020,I159082);
DFFARX1 I_9022  ( .D(I159082), .CLK(I5694_clk), .RSTB(I159031_rst), .Q(I159113) );
not I_9023 (I159008,I159113);
nor I_9024 (I159144,I114287,I114272);
not I_9025 (I159161,I159144);
nor I_9026 (I159178,I159082,I159161);
DFFARX1 I_9027  ( .D(I114293), .CLK(I5694_clk), .RSTB(I159031_rst), .Q(I159195) );
not I_9028 (I159212,I159195);
nand I_9029 (I159011,I159195,I159161);
DFFARX1 I_9030  ( .D(I159195), .CLK(I5694_clk), .RSTB(I159031_rst), .Q(I159243) );
and I_9031 (I158996,I159082,I159243);
nand I_9032 (I159274,I114266,I114269);
and I_9033 (I159291,I159274,I114278);
DFFARX1 I_9034  ( .D(I159291), .CLK(I5694_clk), .RSTB(I159031_rst), .Q(I159308) );
nor I_9035 (I159325,I159308,I159212);
and I_9036 (I159342,I159144,I159325);
nor I_9037 (I159359,I159308,I159082);
DFFARX1 I_9038  ( .D(I159308), .CLK(I5694_clk), .RSTB(I159031_rst), .Q(I159002) );
DFFARX1 I_9039  ( .D(I114296), .CLK(I5694_clk), .RSTB(I159031_rst), .Q(I159390) );
and I_9040 (I159407,I159390,I114290);
or I_9041 (I159424,I159407,I159342);
DFFARX1 I_9042  ( .D(I159424), .CLK(I5694_clk), .RSTB(I159031_rst), .Q(I159014) );
nand I_9043 (I159023,I159407,I159359);
DFFARX1 I_9044  ( .D(I159407), .CLK(I5694_clk), .RSTB(I159031_rst), .Q(I158993) );
DFFARX1 I_9045  ( .D(I114281), .CLK(I5694_clk), .RSTB(I159031_rst), .Q(I159483) );
nand I_9046 (I159017,I159483,I159178);
DFFARX1 I_9047  ( .D(I159483), .CLK(I5694_clk), .RSTB(I159031_rst), .Q(I159005) );
nand I_9048 (I159528,I159483,I159144);
and I_9049 (I159545,I159195,I159528);
DFFARX1 I_9050  ( .D(I159545), .CLK(I5694_clk), .RSTB(I159031_rst), .Q(I158999) );
not I_9051 (I159609_rst,I5701);
nand I_9052 (I159626,I94757,I94742);
and I_9053 (I159643,I159626,I94751);
DFFARX1 I_9054  ( .D(I159643), .CLK(I5694_clk), .RSTB(I159609_rst), .Q(I159660) );
not I_9055 (I159598,I159660);
DFFARX1 I_9056  ( .D(I159660), .CLK(I5694_clk), .RSTB(I159609_rst), .Q(I159691) );
not I_9057 (I159586,I159691);
nor I_9058 (I159722,I94763,I94742);
not I_9059 (I159739,I159722);
nor I_9060 (I159756,I159660,I159739);
DFFARX1 I_9061  ( .D(I94754), .CLK(I5694_clk), .RSTB(I159609_rst), .Q(I159773) );
not I_9062 (I159790,I159773);
nand I_9063 (I159589,I159773,I159739);
DFFARX1 I_9064  ( .D(I159773), .CLK(I5694_clk), .RSTB(I159609_rst), .Q(I159821) );
and I_9065 (I159574,I159660,I159821);
nand I_9066 (I159852,I94739,I94733);
and I_9067 (I159869,I159852,I94748);
DFFARX1 I_9068  ( .D(I159869), .CLK(I5694_clk), .RSTB(I159609_rst), .Q(I159886) );
nor I_9069 (I159903,I159886,I159790);
and I_9070 (I159920,I159722,I159903);
nor I_9071 (I15993_rst7,I159886,I159660);
DFFARX1 I_9072  ( .D(I159886), .CLK(I5694_clk), .RSTB(I159609_rst), .Q(I159580) );
DFFARX1 I_9073  ( .D(I94736), .CLK(I5694_clk), .RSTB(I159609_rst), .Q(I159968) );
and I_9074 (I159985,I159968,I94760);
or I_9075 (I160002,I159985,I159920);
DFFARX1 I_9076  ( .D(I160002), .CLK(I5694_clk), .RSTB(I159609_rst), .Q(I159592) );
nand I_9077 (I159601,I159985,I15993_rst7);
DFFARX1 I_9078  ( .D(I159985), .CLK(I5694_clk), .RSTB(I159609_rst), .Q(I159571) );
DFFARX1 I_9079  ( .D(I94745), .CLK(I5694_clk), .RSTB(I159609_rst), .Q(I160061) );
nand I_9080 (I159595,I160061,I159756);
DFFARX1 I_9081  ( .D(I160061), .CLK(I5694_clk), .RSTB(I159609_rst), .Q(I159583) );
nand I_9082 (I160106,I160061,I159722);
and I_9083 (I160123,I159773,I160106);
DFFARX1 I_9084  ( .D(I160123), .CLK(I5694_clk), .RSTB(I159609_rst), .Q(I159577) );
not I_9085 (I160187_rst,I5701);
nand I_9086 (I160204,I112345,I112375);
and I_9087 (I160221,I160204,I112357);
DFFARX1 I_9088  ( .D(I160221), .CLK(I5694_clk), .RSTB(I160187_rst), .Q(I160238) );
not I_9089 (I160176,I160238);
DFFARX1 I_9090  ( .D(I160238), .CLK(I5694_clk), .RSTB(I160187_rst), .Q(I160269) );
not I_9091 (I160164,I160269);
nor I_9092 (I160300,I112354,I112375);
not I_9093 (I160317,I160300);
nor I_9094 (I160334,I160238,I160317);
DFFARX1 I_9095  ( .D(I112348), .CLK(I5694_clk), .RSTB(I160187_rst), .Q(I160351) );
not I_9096 (I160368,I160351);
nand I_9097 (I160167,I160351,I160317);
DFFARX1 I_9098  ( .D(I160351), .CLK(I5694_clk), .RSTB(I160187_rst), .Q(I160399) );
and I_9099 (I160152,I160238,I160399);
nand I_9100 (I160430,I112351,I112366);
and I_9101 (I160447,I160430,I112363);
DFFARX1 I_9102  ( .D(I160447), .CLK(I5694_clk), .RSTB(I160187_rst), .Q(I160464) );
nor I_9103 (I160481,I160464,I160368);
and I_9104 (I160498,I160300,I160481);
nor I_9105 (I160515,I160464,I160238);
DFFARX1 I_9106  ( .D(I160464), .CLK(I5694_clk), .RSTB(I160187_rst), .Q(I160158) );
DFFARX1 I_9107  ( .D(I112360), .CLK(I5694_clk), .RSTB(I160187_rst), .Q(I160546) );
and I_9108 (I160563,I160546,I112372);
or I_9109 (I160580,I160563,I160498);
DFFARX1 I_9110  ( .D(I160580), .CLK(I5694_clk), .RSTB(I160187_rst), .Q(I160170) );
nand I_9111 (I160179,I160563,I160515);
DFFARX1 I_9112  ( .D(I160563), .CLK(I5694_clk), .RSTB(I160187_rst), .Q(I160149) );
DFFARX1 I_9113  ( .D(I112369), .CLK(I5694_clk), .RSTB(I160187_rst), .Q(I160639) );
nand I_9114 (I160173,I160639,I160334);
DFFARX1 I_9115  ( .D(I160639), .CLK(I5694_clk), .RSTB(I160187_rst), .Q(I160161) );
nand I_9116 (I160684,I160639,I160300);
and I_9117 (I160701,I160351,I160684);
DFFARX1 I_9118  ( .D(I160701), .CLK(I5694_clk), .RSTB(I160187_rst), .Q(I160155) );
not I_9119 (I160765_rst,I5701);
nand I_9120 (I160782,I99973,I99958);
and I_9121 (I160799,I160782,I99952);
DFFARX1 I_9122  ( .D(I160799), .CLK(I5694_clk), .RSTB(I160765_rst), .Q(I160816) );
not I_9123 (I160754,I160816);
DFFARX1 I_9124  ( .D(I160816), .CLK(I5694_clk), .RSTB(I160765_rst), .Q(I160847) );
not I_9125 (I160742,I160847);
nor I_9126 (I160878,I99979,I99958);
not I_9127 (I160895,I160878);
nor I_9128 (I160912,I160816,I160895);
DFFARX1 I_9129  ( .D(I99982), .CLK(I5694_clk), .RSTB(I160765_rst), .Q(I160929) );
not I_9130 (I160946,I160929);
nand I_9131 (I160745,I160929,I160895);
DFFARX1 I_9132  ( .D(I160929), .CLK(I5694_clk), .RSTB(I160765_rst), .Q(I160977) );
and I_9133 (I160730,I160816,I160977);
nand I_9134 (I161008,I99964,I99967);
and I_9135 (I161025,I161008,I99970);
DFFARX1 I_9136  ( .D(I161025), .CLK(I5694_clk), .RSTB(I160765_rst), .Q(I161042) );
nor I_9137 (I161059,I161042,I160946);
and I_9138 (I161076,I160878,I161059);
nor I_9139 (I161093,I161042,I160816);
DFFARX1 I_9140  ( .D(I161042), .CLK(I5694_clk), .RSTB(I160765_rst), .Q(I160736) );
DFFARX1 I_9141  ( .D(I99976), .CLK(I5694_clk), .RSTB(I160765_rst), .Q(I161124) );
and I_9142 (I161141,I161124,I99961);
or I_9143 (I161158,I161141,I161076);
DFFARX1 I_9144  ( .D(I161158), .CLK(I5694_clk), .RSTB(I160765_rst), .Q(I160748) );
nand I_9145 (I160757,I161141,I161093);
DFFARX1 I_9146  ( .D(I161141), .CLK(I5694_clk), .RSTB(I160765_rst), .Q(I160727) );
DFFARX1 I_9147  ( .D(I99955), .CLK(I5694_clk), .RSTB(I160765_rst), .Q(I161217) );
nand I_9148 (I160751,I161217,I160912);
DFFARX1 I_9149  ( .D(I161217), .CLK(I5694_clk), .RSTB(I160765_rst), .Q(I160739) );
nand I_9150 (I161262,I161217,I160878);
and I_9151 (I161279,I160929,I161262);
DFFARX1 I_9152  ( .D(I161279), .CLK(I5694_clk), .RSTB(I160765_rst), .Q(I160733) );
not I_9153 (I161343_rst,I5701);
nand I_9154 (I161360,I128967,I128958);
and I_9155 (I161377,I161360,I128961);
DFFARX1 I_9156  ( .D(I161377), .CLK(I5694_clk), .RSTB(I161343_rst), .Q(I161394) );
not I_9157 (I161411,I161394);
nor I_9158 (I161428,I128937,I128958);
or I_9159 (I161326,I161428,I161394);
not I_9160 (I161314,I161428);
DFFARX1 I_9161  ( .D(I128952), .CLK(I5694_clk), .RSTB(I161343_rst), .Q(I161473) );
nor I_9162 (I161490,I161473,I161428);
nand I_9163 (I161507,I128940,I128955);
and I_9164 (I161524,I161507,I128949);
DFFARX1 I_9165  ( .D(I161524), .CLK(I5694_clk), .RSTB(I161343_rst), .Q(I161541) );
nor I_9166 (I161323,I161541,I161394);
not I_9167 (I161572,I161541);
nor I_9168 (I161589,I161473,I161572);
DFFARX1 I_9169  ( .D(I128964), .CLK(I5694_clk), .RSTB(I161343_rst), .Q(I161606) );
and I_9170 (I161623,I161606,I128943);
or I_9171 (I161332,I161623,I161428);
nand I_9172 (I161311,I161623,I161589);
DFFARX1 I_9173  ( .D(I128946), .CLK(I5694_clk), .RSTB(I161343_rst), .Q(I161668) );
and I_9174 (I161685,I161668,I161411);
nor I_9175 (I161329,I161623,I161685);
nor I_9176 (I161716,I161668,I161473);
DFFARX1 I_9177  ( .D(I161716), .CLK(I5694_clk), .RSTB(I161343_rst), .Q(I161320) );
nor I_9178 (I161335,I161668,I161394);
not I_9179 (I161761,I161668);
nor I_9180 (I161778,I161541,I161761);
and I_9181 (I161795,I161428,I161778);
or I_9182 (I161812,I161623,I161795);
DFFARX1 I_9183  ( .D(I161812), .CLK(I5694_clk), .RSTB(I161343_rst), .Q(I161308) );
nand I_9184 (I161317,I161668,I161490);
nand I_9185 (I161305,I161668,I161572);
not I_9186 (I161904_rst,I5701);
nand I_9187 (I161921,I159002,I159023);
and I_9188 (I161938,I161921,I159011);
DFFARX1 I_9189  ( .D(I161938), .CLK(I5694_clk), .RSTB(I161904_rst), .Q(I161955) );
not I_9190 (I161972,I161955);
nor I_9191 (I161989,I159017,I159023);
or I_9192 (I161887,I161989,I161955);
not I_9193 (I161875,I161989);
DFFARX1 I_9194  ( .D(I159005), .CLK(I5694_clk), .RSTB(I161904_rst), .Q(I162034) );
nor I_9195 (I162051,I162034,I161989);
nand I_9196 (I162068,I158996,I159014);
and I_9197 (I162085,I162068,I159008);
DFFARX1 I_9198  ( .D(I162085), .CLK(I5694_clk), .RSTB(I161904_rst), .Q(I162102) );
nor I_9199 (I161884,I162102,I161955);
not I_9200 (I162133,I162102);
nor I_9201 (I162150,I162034,I162133);
DFFARX1 I_9202  ( .D(I159020), .CLK(I5694_clk), .RSTB(I161904_rst), .Q(I162167) );
and I_9203 (I162184,I162167,I158993);
or I_9204 (I161893,I162184,I161989);
nand I_9205 (I161872,I162184,I162150);
DFFARX1 I_9206  ( .D(I158999), .CLK(I5694_clk), .RSTB(I161904_rst), .Q(I162229) );
and I_9207 (I162246,I162229,I161972);
nor I_9208 (I161890,I162184,I162246);
nor I_9209 (I162277,I162229,I162034);
DFFARX1 I_9210  ( .D(I162277), .CLK(I5694_clk), .RSTB(I161904_rst), .Q(I161881) );
nor I_9211 (I161896,I162229,I161955);
not I_9212 (I162322,I162229);
nor I_9213 (I162339,I162102,I162322);
and I_9214 (I162356,I161989,I162339);
or I_9215 (I162373,I162184,I162356);
DFFARX1 I_9216  ( .D(I162373), .CLK(I5694_clk), .RSTB(I161904_rst), .Q(I161869) );
nand I_9217 (I161878,I162229,I162051);
nand I_9218 (I161866,I162229,I162133);
not I_9219 (I162465_rst,I5701);
nand I_9220 (I162482,I141479,I141461);
and I_9221 (I162499,I162482,I141470);
DFFARX1 I_9222  ( .D(I162499), .CLK(I5694_clk), .RSTB(I162465_rst), .Q(I162516) );
not I_9223 (I162533,I162516);
nor I_9224 (I162550,I141455,I141461);
or I_9225 (I162448,I162550,I162516);
not I_9226 (I162436,I162550);
DFFARX1 I_9227  ( .D(I141464), .CLK(I5694_clk), .RSTB(I162465_rst), .Q(I162595) );
nor I_9228 (I162612,I162595,I162550);
nand I_9229 (I162629,I141452,I141458);
and I_9230 (I162646,I162629,I141467);
DFFARX1 I_9231  ( .D(I162646), .CLK(I5694_clk), .RSTB(I162465_rst), .Q(I162663) );
nor I_9232 (I162445,I162663,I162516);
not I_9233 (I162694,I162663);
nor I_9234 (I162711,I162595,I162694);
DFFARX1 I_9235  ( .D(I141476), .CLK(I5694_clk), .RSTB(I162465_rst), .Q(I162728) );
and I_9236 (I162745,I162728,I141449);
or I_9237 (I162454,I162745,I162550);
nand I_9238 (I162433,I162745,I162711);
DFFARX1 I_9239  ( .D(I141473), .CLK(I5694_clk), .RSTB(I162465_rst), .Q(I162790) );
and I_9240 (I162807,I162790,I162533);
nor I_9241 (I162451,I162745,I162807);
nor I_9242 (I162838,I162790,I162595);
DFFARX1 I_9243  ( .D(I162838), .CLK(I5694_clk), .RSTB(I162465_rst), .Q(I162442) );
nor I_9244 (I162457,I162790,I162516);
not I_9245 (I162883,I162790);
nor I_9246 (I162900,I162663,I162883);
and I_9247 (I162917,I162550,I162900);
or I_9248 (I162934,I162745,I162917);
DFFARX1 I_9249  ( .D(I162934), .CLK(I5694_clk), .RSTB(I162465_rst), .Q(I162430) );
nand I_9250 (I162439,I162790,I162612);
nand I_9251 (I162427,I162790,I162694);
not I_9252 (I163026_rst,I5701);
nand I_9253 (I163043,I132843,I132834);
and I_9254 (I163060,I163043,I132837);
DFFARX1 I_9255  ( .D(I163060), .CLK(I5694_clk), .RSTB(I163026_rst), .Q(I163077) );
not I_9256 (I163094,I163077);
nor I_9257 (I163111,I132813,I132834);
or I_9258 (I163009,I163111,I163077);
not I_9259 (I162997,I163111);
DFFARX1 I_9260  ( .D(I132828), .CLK(I5694_clk), .RSTB(I163026_rst), .Q(I163156) );
nor I_9261 (I163173,I163156,I163111);
nand I_9262 (I163190,I132816,I132831);
and I_9263 (I163207,I163190,I132825);
DFFARX1 I_9264  ( .D(I163207), .CLK(I5694_clk), .RSTB(I163026_rst), .Q(I163224) );
nor I_9265 (I163006,I163224,I163077);
not I_9266 (I163255,I163224);
nor I_9267 (I163272,I163156,I163255);
DFFARX1 I_9268  ( .D(I132840), .CLK(I5694_clk), .RSTB(I163026_rst), .Q(I163289) );
and I_9269 (I163306,I163289,I132819);
or I_9270 (I163015,I163306,I163111);
nand I_9271 (I162994,I163306,I163272);
DFFARX1 I_9272  ( .D(I132822), .CLK(I5694_clk), .RSTB(I163026_rst), .Q(I163351) );
and I_9273 (I163368,I163351,I163094);
nor I_9274 (I163012,I163306,I163368);
nor I_9275 (I163399,I163351,I163156);
DFFARX1 I_9276  ( .D(I163399), .CLK(I5694_clk), .RSTB(I163026_rst), .Q(I163003) );
nor I_9277 (I163018,I163351,I163077);
not I_9278 (I163444,I163351);
nor I_9279 (I163461,I163224,I163444);
and I_9280 (I163478,I163111,I163461);
or I_9281 (I163495,I163306,I163478);
DFFARX1 I_9282  ( .D(I163495), .CLK(I5694_clk), .RSTB(I163026_rst), .Q(I162991) );
nand I_9283 (I163000,I163351,I163173);
nand I_9284 (I162988,I163351,I163255);
not I_9285 (I163587_rst,I5701);
nand I_9286 (I163604,I155848,I155851);
and I_9287 (I163621,I163604,I155857);
DFFARX1 I_9288  ( .D(I163621), .CLK(I5694_clk), .RSTB(I163587_rst), .Q(I163638) );
not I_9289 (I163655,I163638);
nor I_9290 (I163672,I155869,I155851);
or I_9291 (I163570,I163672,I163638);
not I_9292 (I163558,I163672);
DFFARX1 I_9293  ( .D(I155878), .CLK(I5694_clk), .RSTB(I163587_rst), .Q(I163717) );
nor I_9294 (I163734,I163717,I163672);
nand I_9295 (I163751,I155866,I155863);
and I_9296 (I163768,I163751,I155875);
DFFARX1 I_9297  ( .D(I163768), .CLK(I5694_clk), .RSTB(I163587_rst), .Q(I163785) );
nor I_9298 (I163567,I163785,I163638);
not I_9299 (I163816,I163785);
nor I_9300 (I163833,I163717,I163816);
DFFARX1 I_9301  ( .D(I155872), .CLK(I5694_clk), .RSTB(I163587_rst), .Q(I163850) );
and I_9302 (I163867,I163850,I155860);
or I_9303 (I163576,I163867,I163672);
nand I_9304 (I163555,I163867,I163833);
DFFARX1 I_9305  ( .D(I155854), .CLK(I5694_clk), .RSTB(I163587_rst), .Q(I163912) );
and I_9306 (I163929,I163912,I163655);
nor I_9307 (I163573,I163867,I163929);
nor I_9308 (I163960,I163912,I163717);
DFFARX1 I_9309  ( .D(I163960), .CLK(I5694_clk), .RSTB(I163587_rst), .Q(I163564) );
nor I_9310 (I163579,I163912,I163638);
not I_9311 (I164005,I163912);
nor I_9312 (I164022,I163785,I164005);
and I_9313 (I164039,I163672,I164022);
or I_9314 (I164056,I163867,I164039);
DFFARX1 I_9315  ( .D(I164056), .CLK(I5694_clk), .RSTB(I163587_rst), .Q(I163552) );
nand I_9316 (I163561,I163912,I163734);
nand I_9317 (I163549,I163912,I163816);
not I_9318 (I164148_rst,I5701);
nand I_9319 (I164165,I140867,I140849);
and I_9320 (I164182,I164165,I140858);
DFFARX1 I_9321  ( .D(I164182), .CLK(I5694_clk), .RSTB(I164148_rst), .Q(I164199) );
not I_9322 (I164216,I164199);
nor I_9323 (I164233,I140843,I140849);
or I_9324 (I164131,I164233,I164199);
not I_9325 (I164119,I164233);
DFFARX1 I_9326  ( .D(I140852), .CLK(I5694_clk), .RSTB(I164148_rst), .Q(I164278) );
nor I_9327 (I164295,I164278,I164233);
nand I_9328 (I164312,I140840,I140846);
and I_9329 (I164329,I164312,I140855);
DFFARX1 I_9330  ( .D(I164329), .CLK(I5694_clk), .RSTB(I164148_rst), .Q(I164346) );
nor I_9331 (I164128,I164346,I164199);
not I_9332 (I164377,I164346);
nor I_9333 (I164394,I164278,I164377);
DFFARX1 I_9334  ( .D(I140864), .CLK(I5694_clk), .RSTB(I164148_rst), .Q(I164411) );
and I_9335 (I164428,I164411,I140837);
or I_9336 (I164137,I164428,I164233);
nand I_9337 (I164116,I164428,I164394);
DFFARX1 I_9338  ( .D(I140861), .CLK(I5694_clk), .RSTB(I164148_rst), .Q(I164473) );
and I_9339 (I164490,I164473,I164216);
nor I_9340 (I164134,I164428,I164490);
nor I_9341 (I164521,I164473,I164278);
DFFARX1 I_9342  ( .D(I164521), .CLK(I5694_clk), .RSTB(I164148_rst), .Q(I164125) );
nor I_9343 (I164140,I164473,I164199);
not I_9344 (I164566,I164473);
nor I_9345 (I164583,I164346,I164566);
and I_9346 (I164600,I164233,I164583);
or I_9347 (I164617,I164428,I164600);
DFFARX1 I_9348  ( .D(I164617), .CLK(I5694_clk), .RSTB(I164148_rst), .Q(I164113) );
nand I_9349 (I164122,I164473,I164295);
nand I_9350 (I164110,I164473,I164377);
not I_9351 (I164709_rst,I5701);
not I_9352 (I164726,I164113);
nor I_9353 (I164743,I164125,I164110);
nand I_9354 (I164760,I164743,I164122);
DFFARX1 I_9355  ( .D(I164760), .CLK(I5694_clk), .RSTB(I164709_rst), .Q(I164683) );
nor I_9356 (I164791,I164726,I164125);
nand I_9357 (I164808,I164791,I164140);
not I_9358 (I164698,I164808);
DFFARX1 I_9359  ( .D(I164808), .CLK(I5694_clk), .RSTB(I164709_rst), .Q(I164680) );
not I_9360 (I164853,I164125);
not I_9361 (I164870,I164853);
not I_9362 (I164887,I164116);
nor I_9363 (I164904,I164887,I164128);
and I_9364 (I164921,I164904,I164119);
or I_9365 (I164938,I164921,I164134);
DFFARX1 I_9366  ( .D(I164938), .CLK(I5694_clk), .RSTB(I164709_rst), .Q(I164955) );
nor I_9367 (I164972,I164955,I164808);
nor I_9368 (I164989,I164955,I164870);
nand I_9369 (I164695,I164760,I164989);
nand I_9370 (I165020,I164726,I164116);
nand I_9371 (I165037,I165020,I164955);
and I_9372 (I165054,I165020,I165037);
DFFARX1 I_9373  ( .D(I165054), .CLK(I5694_clk), .RSTB(I164709_rst), .Q(I164677) );
DFFARX1 I_9374  ( .D(I165020), .CLK(I5694_clk), .RSTB(I164709_rst), .Q(I165085) );
and I_9375 (I164674,I164853,I165085);
DFFARX1 I_9376  ( .D(I164137), .CLK(I5694_clk), .RSTB(I164709_rst), .Q(I165116) );
not I_9377 (I165133,I165116);
nor I_9378 (I165150,I164808,I165133);
and I_9379 (I165167,I165116,I165150);
nand I_9380 (I164689,I165116,I164870);
DFFARX1 I_9381  ( .D(I165116), .CLK(I5694_clk), .RSTB(I164709_rst), .Q(I165198) );
not I_9382 (I164686,I165198);
DFFARX1 I_9383  ( .D(I164131), .CLK(I5694_clk), .RSTB(I164709_rst), .Q(I165229) );
not I_9384 (I165246,I165229);
or I_9385 (I165263,I165246,I165167);
DFFARX1 I_9386  ( .D(I165263), .CLK(I5694_clk), .RSTB(I164709_rst), .Q(I164692) );
nand I_9387 (I164701,I165246,I164972);
DFFARX1 I_9388  ( .D(I165246), .CLK(I5694_clk), .RSTB(I164709_rst), .Q(I164671) );
not I_9389 (I165355_rst,I5701);
not I_9390 (I165372,I111700);
nor I_9391 (I165389,I111688,I111694);
nand I_9392 (I165406,I165389,I111703);
DFFARX1 I_9393  ( .D(I165406), .CLK(I5694_clk), .RSTB(I165355_rst), .Q(I165329) );
nor I_9394 (I165437,I165372,I111688);
nand I_9395 (I165454,I165437,I111691);
not I_9396 (I165344,I165454);
DFFARX1 I_9397  ( .D(I165454), .CLK(I5694_clk), .RSTB(I165355_rst), .Q(I165326) );
not I_9398 (I165499,I111688);
not I_9399 (I165516,I165499);
not I_9400 (I165533,I111712);
nor I_9401 (I165550,I165533,I111685);
and I_9402 (I165567,I165550,I111706);
or I_9403 (I165584,I165567,I111697);
DFFARX1 I_9404  ( .D(I165584), .CLK(I5694_clk), .RSTB(I165355_rst), .Q(I165601) );
nor I_9405 (I165618,I165601,I165454);
nor I_9406 (I165635,I165601,I165516);
nand I_9407 (I165341,I165406,I165635);
nand I_9408 (I165666,I165372,I111712);
nand I_9409 (I165683,I165666,I165601);
and I_9410 (I165700,I165666,I165683);
DFFARX1 I_9411  ( .D(I165700), .CLK(I5694_clk), .RSTB(I165355_rst), .Q(I165323) );
DFFARX1 I_9412  ( .D(I165666), .CLK(I5694_clk), .RSTB(I165355_rst), .Q(I165731) );
and I_9413 (I165320,I165499,I165731);
DFFARX1 I_9414  ( .D(I111682), .CLK(I5694_clk), .RSTB(I165355_rst), .Q(I165762) );
not I_9415 (I165779,I165762);
nor I_9416 (I165796,I165454,I165779);
and I_9417 (I165813,I165762,I165796);
nand I_9418 (I165335,I165762,I165516);
DFFARX1 I_9419  ( .D(I165762), .CLK(I5694_clk), .RSTB(I165355_rst), .Q(I165844) );
not I_9420 (I165332,I165844);
DFFARX1 I_9421  ( .D(I111709), .CLK(I5694_clk), .RSTB(I165355_rst), .Q(I165875) );
not I_9422 (I165892,I165875);
or I_9423 (I165909,I165892,I165813);
DFFARX1 I_9424  ( .D(I165909), .CLK(I5694_clk), .RSTB(I165355_rst), .Q(I165338) );
nand I_9425 (I165347,I165892,I165618);
DFFARX1 I_9426  ( .D(I165892), .CLK(I5694_clk), .RSTB(I165355_rst), .Q(I165317) );
not I_9427 (I166001_rst,I5701);
not I_9428 (I166018,I130893);
nor I_9429 (I166035,I130905,I130887);
nand I_9430 (I166052,I166035,I130902);
DFFARX1 I_9431  ( .D(I166052), .CLK(I5694_clk), .RSTB(I166001_rst), .Q(I165975) );
nor I_9432 (I166083,I166018,I130905);
nand I_9433 (I166100,I166083,I130890);
not I_9434 (I165990,I166100);
DFFARX1 I_9435  ( .D(I166100), .CLK(I5694_clk), .RSTB(I166001_rst), .Q(I165972) );
not I_9436 (I166145,I130905);
not I_9437 (I166162,I166145);
not I_9438 (I166179,I130899);
nor I_9439 (I166196,I166179,I130878);
and I_9440 (I166213,I166196,I130881);
or I_9441 (I166230,I166213,I130884);
DFFARX1 I_9442  ( .D(I166230), .CLK(I5694_clk), .RSTB(I166001_rst), .Q(I166247) );
nor I_9443 (I166264,I166247,I166100);
nor I_9444 (I166281,I166247,I166162);
nand I_9445 (I165987,I166052,I166281);
nand I_9446 (I166312,I166018,I130899);
nand I_9447 (I166329,I166312,I166247);
and I_9448 (I166346,I166312,I166329);
DFFARX1 I_9449  ( .D(I166346), .CLK(I5694_clk), .RSTB(I166001_rst), .Q(I165969) );
DFFARX1 I_9450  ( .D(I166312), .CLK(I5694_clk), .RSTB(I166001_rst), .Q(I166377) );
and I_9451 (I165966,I166145,I166377);
DFFARX1 I_9452  ( .D(I130875), .CLK(I5694_clk), .RSTB(I166001_rst), .Q(I166408) );
not I_9453 (I166425,I166408);
nor I_9454 (I166442,I166100,I166425);
and I_9455 (I166459,I166408,I166442);
nand I_9456 (I165981,I166408,I166162);
DFFARX1 I_9457  ( .D(I166408), .CLK(I5694_clk), .RSTB(I166001_rst), .Q(I166490) );
not I_9458 (I165978,I166490);
DFFARX1 I_9459  ( .D(I130896), .CLK(I5694_clk), .RSTB(I166001_rst), .Q(I166521) );
not I_9460 (I166538,I166521);
or I_9461 (I166555,I166538,I166459);
DFFARX1 I_9462  ( .D(I166555), .CLK(I5694_clk), .RSTB(I166001_rst), .Q(I165984) );
nand I_9463 (I165993,I166538,I166264);
DFFARX1 I_9464  ( .D(I166538), .CLK(I5694_clk), .RSTB(I166001_rst), .Q(I165963) );
not I_9465 (I166647_rst,I5701);
not I_9466 (I166664,I145624);
nor I_9467 (I166681,I145600,I145606);
nand I_9468 (I166698,I166681,I145609);
DFFARX1 I_9469  ( .D(I166698), .CLK(I5694_clk), .RSTB(I166647_rst), .Q(I166621) );
nor I_9470 (I166729,I166664,I145600);
nand I_9471 (I166746,I166729,I145618);
not I_9472 (I166636,I166746);
DFFARX1 I_9473  ( .D(I166746), .CLK(I5694_clk), .RSTB(I166647_rst), .Q(I166618) );
not I_9474 (I166791,I145600);
not I_9475 (I166808,I166791);
not I_9476 (I166825,I145597);
nor I_9477 (I166842,I166825,I145612);
and I_9478 (I166859,I166842,I145603);
or I_9479 (I166876,I166859,I145615);
DFFARX1 I_9480  ( .D(I166876), .CLK(I5694_clk), .RSTB(I166647_rst), .Q(I166893) );
nor I_9481 (I166910,I166893,I166746);
nor I_9482 (I166927,I166893,I166808);
nand I_9483 (I166633,I166698,I166927);
nand I_9484 (I166958,I166664,I145597);
nand I_9485 (I166975,I166958,I166893);
and I_9486 (I166992,I166958,I166975);
DFFARX1 I_9487  ( .D(I166992), .CLK(I5694_clk), .RSTB(I166647_rst), .Q(I166615) );
DFFARX1 I_9488  ( .D(I166958), .CLK(I5694_clk), .RSTB(I166647_rst), .Q(I167023) );
and I_9489 (I166612,I166791,I167023);
DFFARX1 I_9490  ( .D(I145627), .CLK(I5694_clk), .RSTB(I166647_rst), .Q(I167054) );
not I_9491 (I167071,I167054);
nor I_9492 (I167088,I166746,I167071);
and I_9493 (I167105,I167054,I167088);
nand I_9494 (I166627,I167054,I166808);
DFFARX1 I_9495  ( .D(I167054), .CLK(I5694_clk), .RSTB(I166647_rst), .Q(I167136) );
not I_9496 (I166624,I167136);
DFFARX1 I_9497  ( .D(I145621), .CLK(I5694_clk), .RSTB(I166647_rst), .Q(I167167) );
not I_9498 (I167184,I167167);
or I_9499 (I167201,I167184,I167105);
DFFARX1 I_9500  ( .D(I167201), .CLK(I5694_clk), .RSTB(I166647_rst), .Q(I166630) );
nand I_9501 (I166639,I167184,I166910);
DFFARX1 I_9502  ( .D(I167184), .CLK(I5694_clk), .RSTB(I166647_rst), .Q(I166609) );
not I_9503 (I167293_rst,I5701);
not I_9504 (I167310,I125011);
nor I_9505 (I167327,I125008,I124996);
nand I_9506 (I167344,I167327,I124999);
DFFARX1 I_9507  ( .D(I167344), .CLK(I5694_clk), .RSTB(I167293_rst), .Q(I167267) );
nor I_9508 (I167375,I167310,I125008);
nand I_9509 (I167392,I167375,I125005);
not I_9510 (I167282,I167392);
DFFARX1 I_9511  ( .D(I167392), .CLK(I5694_clk), .RSTB(I167293_rst), .Q(I167264) );
not I_9512 (I167437,I125008);
not I_9513 (I167454,I167437);
not I_9514 (I167471,I125017);
nor I_9515 (I167488,I167471,I124993);
and I_9516 (I167505,I167488,I125014);
or I_9517 (I167522,I167505,I125002);
DFFARX1 I_9518  ( .D(I167522), .CLK(I5694_clk), .RSTB(I167293_rst), .Q(I167539) );
nor I_9519 (I167556,I167539,I167392);
nor I_9520 (I167573,I167539,I167454);
nand I_9521 (I167279,I167344,I167573);
nand I_9522 (I167604,I167310,I125017);
nand I_9523 (I167621,I167604,I167539);
and I_9524 (I167638,I167604,I167621);
DFFARX1 I_9525  ( .D(I167638), .CLK(I5694_clk), .RSTB(I167293_rst), .Q(I167261) );
DFFARX1 I_9526  ( .D(I167604), .CLK(I5694_clk), .RSTB(I167293_rst), .Q(I167669) );
and I_9527 (I167258,I167437,I167669);
DFFARX1 I_9528  ( .D(I125023), .CLK(I5694_clk), .RSTB(I167293_rst), .Q(I167700) );
not I_9529 (I167717,I167700);
nor I_9530 (I167734,I167392,I167717);
and I_9531 (I167751,I167700,I167734);
nand I_9532 (I167273,I167700,I167454);
DFFARX1 I_9533  ( .D(I167700), .CLK(I5694_clk), .RSTB(I167293_rst), .Q(I167782) );
not I_9534 (I167270,I167782);
DFFARX1 I_9535  ( .D(I125020), .CLK(I5694_clk), .RSTB(I167293_rst), .Q(I167813) );
not I_9536 (I167830,I167813);
or I_9537 (I167847,I167830,I167751);
DFFARX1 I_9538  ( .D(I167847), .CLK(I5694_clk), .RSTB(I167293_rst), .Q(I167276) );
nand I_9539 (I167285,I167830,I167556);
DFFARX1 I_9540  ( .D(I167830), .CLK(I5694_clk), .RSTB(I167293_rst), .Q(I167255) );
not I_9541 (I167939_rst,I5701);
not I_9542 (I167956,I154590);
nor I_9543 (I167973,I154605,I154620);
nand I_9544 (I167990,I167973,I154608);
DFFARX1 I_9545  ( .D(I167990), .CLK(I5694_clk), .RSTB(I167939_rst), .Q(I167913) );
nor I_9546 (I168021,I167956,I154605);
nand I_9547 (I168038,I168021,I154611);
not I_9548 (I167928,I168038);
DFFARX1 I_9549  ( .D(I168038), .CLK(I5694_clk), .RSTB(I167939_rst), .Q(I167910) );
not I_9550 (I168083,I154605);
not I_9551 (I168100,I168083);
not I_9552 (I168117,I154617);
nor I_9553 (I168134,I168117,I154614);
and I_9554 (I168151,I168134,I154593);
or I_9555 (I168168,I168151,I154602);
DFFARX1 I_9556  ( .D(I168168), .CLK(I5694_clk), .RSTB(I167939_rst), .Q(I168185) );
nor I_9557 (I168202,I168185,I168038);
nor I_9558 (I168219,I168185,I168100);
nand I_9559 (I167925,I167990,I168219);
nand I_9560 (I168250,I167956,I154617);
nand I_9561 (I168267,I168250,I168185);
and I_9562 (I168284,I168250,I168267);
DFFARX1 I_9563  ( .D(I168284), .CLK(I5694_clk), .RSTB(I167939_rst), .Q(I167907) );
DFFARX1 I_9564  ( .D(I168250), .CLK(I5694_clk), .RSTB(I167939_rst), .Q(I168315) );
and I_9565 (I167904,I168083,I168315);
DFFARX1 I_9566  ( .D(I154599), .CLK(I5694_clk), .RSTB(I167939_rst), .Q(I168346) );
not I_9567 (I168363,I168346);
nor I_9568 (I168380,I168038,I168363);
and I_9569 (I168397,I168346,I168380);
nand I_9570 (I167919,I168346,I168100);
DFFARX1 I_9571  ( .D(I168346), .CLK(I5694_clk), .RSTB(I167939_rst), .Q(I168428) );
not I_9572 (I167916,I168428);
DFFARX1 I_9573  ( .D(I154596), .CLK(I5694_clk), .RSTB(I167939_rst), .Q(I168459) );
not I_9574 (I168476,I168459);
or I_9575 (I168493,I168476,I168397);
DFFARX1 I_9576  ( .D(I168493), .CLK(I5694_clk), .RSTB(I167939_rst), .Q(I167922) );
nand I_9577 (I167931,I168476,I168202);
DFFARX1 I_9578  ( .D(I168476), .CLK(I5694_clk), .RSTB(I167939_rst), .Q(I167901) );
not I_9579 (I168585_rst,I5701);
not I_9580 (I168602,I115456);
nor I_9581 (I168619,I115486,I115465);
nand I_9582 (I168636,I168619,I115477);
DFFARX1 I_9583  ( .D(I168636), .CLK(I5694_clk), .RSTB(I168585_rst), .Q(I168559) );
nor I_9584 (I168667,I168602,I115486);
nand I_9585 (I168684,I168667,I115459);
not I_9586 (I168574,I168684);
DFFARX1 I_9587  ( .D(I168684), .CLK(I5694_clk), .RSTB(I168585_rst), .Q(I168556) );
not I_9588 (I168729,I115486);
not I_9589 (I168746,I168729);
not I_9590 (I168763,I115462);
nor I_9591 (I168780,I168763,I115480);
and I_9592 (I168797,I168780,I115471);
or I_9593 (I168814,I168797,I115468);
DFFARX1 I_9594  ( .D(I168814), .CLK(I5694_clk), .RSTB(I168585_rst), .Q(I168831) );
nor I_9595 (I168848,I168831,I168684);
nor I_9596 (I168865,I168831,I168746);
nand I_9597 (I168571,I168636,I168865);
nand I_9598 (I168896,I168602,I115462);
nand I_9599 (I168913,I168896,I168831);
and I_9600 (I168930,I168896,I168913);
DFFARX1 I_9601  ( .D(I168930), .CLK(I5694_clk), .RSTB(I168585_rst), .Q(I168553) );
DFFARX1 I_9602  ( .D(I168896), .CLK(I5694_clk), .RSTB(I168585_rst), .Q(I168961) );
and I_9603 (I168550,I168729,I168961);
DFFARX1 I_9604  ( .D(I115474), .CLK(I5694_clk), .RSTB(I168585_rst), .Q(I168992) );
not I_9605 (I169009,I168992);
nor I_9606 (I169026,I168684,I169009);
and I_9607 (I169043,I168992,I169026);
nand I_9608 (I168565,I168992,I168746);
DFFARX1 I_9609  ( .D(I168992), .CLK(I5694_clk), .RSTB(I168585_rst), .Q(I169074) );
not I_9610 (I168562,I169074);
DFFARX1 I_9611  ( .D(I115483), .CLK(I5694_clk), .RSTB(I168585_rst), .Q(I169105) );
not I_9612 (I169122,I169105);
or I_9613 (I169139,I169122,I169043);
DFFARX1 I_9614  ( .D(I169139), .CLK(I5694_clk), .RSTB(I168585_rst), .Q(I168568) );
nand I_9615 (I168577,I169122,I168848);
DFFARX1 I_9616  ( .D(I169122), .CLK(I5694_clk), .RSTB(I168585_rst), .Q(I168547) );
not I_9617 (I169231_rst,I5701);
not I_9618 (I169248,I123685);
nor I_9619 (I169265,I123682,I123670);
nand I_9620 (I169282,I169265,I123673);
DFFARX1 I_9621  ( .D(I169282), .CLK(I5694_clk), .RSTB(I169231_rst), .Q(I169205) );
nor I_9622 (I169313,I169248,I123682);
nand I_9623 (I169330,I169313,I123679);
not I_9624 (I169220,I169330);
DFFARX1 I_9625  ( .D(I169330), .CLK(I5694_clk), .RSTB(I169231_rst), .Q(I169202) );
not I_9626 (I169375,I123682);
not I_9627 (I169392,I169375);
not I_9628 (I169409,I123691);
nor I_9629 (I169426,I169409,I123667);
and I_9630 (I169443,I169426,I123688);
or I_9631 (I169460,I169443,I123676);
DFFARX1 I_9632  ( .D(I169460), .CLK(I5694_clk), .RSTB(I169231_rst), .Q(I169477) );
nor I_9633 (I169494,I169477,I169330);
nor I_9634 (I169511,I169477,I169392);
nand I_9635 (I169217,I169282,I169511);
nand I_9636 (I169542,I169248,I123691);
nand I_9637 (I169559,I169542,I169477);
and I_9638 (I169576,I169542,I169559);
DFFARX1 I_9639  ( .D(I169576), .CLK(I5694_clk), .RSTB(I169231_rst), .Q(I169199) );
DFFARX1 I_9640  ( .D(I169542), .CLK(I5694_clk), .RSTB(I169231_rst), .Q(I169607) );
and I_9641 (I169196,I169375,I169607);
DFFARX1 I_9642  ( .D(I123697), .CLK(I5694_clk), .RSTB(I169231_rst), .Q(I169638) );
not I_9643 (I169655,I169638);
nor I_9644 (I169672,I169330,I169655);
and I_9645 (I169689,I169638,I169672);
nand I_9646 (I169211,I169638,I169392);
DFFARX1 I_9647  ( .D(I169638), .CLK(I5694_clk), .RSTB(I169231_rst), .Q(I169720) );
not I_9648 (I169208,I169720);
DFFARX1 I_9649  ( .D(I123694), .CLK(I5694_clk), .RSTB(I169231_rst), .Q(I169751) );
not I_9650 (I169768,I169751);
or I_9651 (I169785,I169768,I169689);
DFFARX1 I_9652  ( .D(I169785), .CLK(I5694_clk), .RSTB(I169231_rst), .Q(I169214) );
nand I_9653 (I169223,I169768,I169494);
DFFARX1 I_9654  ( .D(I169768), .CLK(I5694_clk), .RSTB(I169231_rst), .Q(I169193) );
not I_9655 (I169877_rst,I5701);
not I_9656 (I169894,I117836);
nor I_9657 (I169911,I117866,I117845);
nand I_9658 (I169928,I169911,I117857);
DFFARX1 I_9659  ( .D(I169928), .CLK(I5694_clk), .RSTB(I169877_rst), .Q(I169851) );
nor I_9660 (I169959,I169894,I117866);
nand I_9661 (I169976,I169959,I117839);
not I_9662 (I169866,I169976);
DFFARX1 I_9663  ( .D(I169976), .CLK(I5694_clk), .RSTB(I169877_rst), .Q(I169848) );
not I_9664 (I170021,I117866);
not I_9665 (I170038,I170021);
not I_9666 (I170055,I117842);
nor I_9667 (I170072,I170055,I117860);
and I_9668 (I170089,I170072,I117851);
or I_9669 (I170106,I170089,I117848);
DFFARX1 I_9670  ( .D(I170106), .CLK(I5694_clk), .RSTB(I169877_rst), .Q(I170123) );
nor I_9671 (I170140,I170123,I169976);
nor I_9672 (I170157,I170123,I170038);
nand I_9673 (I169863,I169928,I170157);
nand I_9674 (I170188,I169894,I117842);
nand I_9675 (I170205,I170188,I170123);
and I_9676 (I170222,I170188,I170205);
DFFARX1 I_9677  ( .D(I170222), .CLK(I5694_clk), .RSTB(I169877_rst), .Q(I169845) );
DFFARX1 I_9678  ( .D(I170188), .CLK(I5694_clk), .RSTB(I169877_rst), .Q(I170253) );
and I_9679 (I169842,I170021,I170253);
DFFARX1 I_9680  ( .D(I117854), .CLK(I5694_clk), .RSTB(I169877_rst), .Q(I170284) );
not I_9681 (I170301,I170284);
nor I_9682 (I170318,I169976,I170301);
and I_9683 (I170335,I170284,I170318);
nand I_9684 (I169857,I170284,I170038);
DFFARX1 I_9685  ( .D(I170284), .CLK(I5694_clk), .RSTB(I169877_rst), .Q(I170366) );
not I_9686 (I169854,I170366);
DFFARX1 I_9687  ( .D(I117863), .CLK(I5694_clk), .RSTB(I169877_rst), .Q(I170397) );
not I_9688 (I170414,I170397);
or I_9689 (I170431,I170414,I170335);
DFFARX1 I_9690  ( .D(I170431), .CLK(I5694_clk), .RSTB(I169877_rst), .Q(I169860) );
nand I_9691 (I169869,I170414,I170140);
DFFARX1 I_9692  ( .D(I170414), .CLK(I5694_clk), .RSTB(I169877_rst), .Q(I169839) );
not I_9693 (I170523_rst,I5701);
not I_9694 (I170540,I157106);
nor I_9695 (I170557,I157121,I157136);
nand I_9696 (I170574,I170557,I157124);
DFFARX1 I_9697  ( .D(I170574), .CLK(I5694_clk), .RSTB(I170523_rst), .Q(I170497) );
nor I_9698 (I170605,I170540,I157121);
nand I_9699 (I170622,I170605,I157127);
not I_9700 (I170512,I170622);
DFFARX1 I_9701  ( .D(I170622), .CLK(I5694_clk), .RSTB(I170523_rst), .Q(I170494) );
not I_9702 (I170667,I157121);
not I_9703 (I170684,I170667);
not I_9704 (I170701,I157133);
nor I_9705 (I170718,I170701,I157130);
and I_9706 (I170735,I170718,I157109);
or I_9707 (I170752,I170735,I157118);
DFFARX1 I_9708  ( .D(I170752), .CLK(I5694_clk), .RSTB(I170523_rst), .Q(I170769) );
nor I_9709 (I170786,I170769,I170622);
nor I_9710 (I170803,I170769,I170684);
nand I_9711 (I170509,I170574,I170803);
nand I_9712 (I170834,I170540,I157133);
nand I_9713 (I170851,I170834,I170769);
and I_9714 (I170868,I170834,I170851);
DFFARX1 I_9715  ( .D(I170868), .CLK(I5694_clk), .RSTB(I170523_rst), .Q(I170491) );
DFFARX1 I_9716  ( .D(I170834), .CLK(I5694_clk), .RSTB(I170523_rst), .Q(I170899) );
and I_9717 (I170488,I170667,I170899);
DFFARX1 I_9718  ( .D(I157115), .CLK(I5694_clk), .RSTB(I170523_rst), .Q(I170930) );
not I_9719 (I170947,I170930);
nor I_9720 (I170964,I170622,I170947);
and I_9721 (I170981,I170930,I170964);
nand I_9722 (I170503,I170930,I170684);
DFFARX1 I_9723  ( .D(I170930), .CLK(I5694_clk), .RSTB(I170523_rst), .Q(I171012) );
not I_9724 (I170500,I171012);
DFFARX1 I_9725  ( .D(I157112), .CLK(I5694_clk), .RSTB(I170523_rst), .Q(I171043) );
not I_9726 (I171060,I171043);
or I_9727 (I171077,I171060,I170981);
DFFARX1 I_9728  ( .D(I171077), .CLK(I5694_clk), .RSTB(I170523_rst), .Q(I170506) );
nand I_9729 (I170515,I171060,I170786);
DFFARX1 I_9730  ( .D(I171060), .CLK(I5694_clk), .RSTB(I170523_rst), .Q(I170485) );
not I_9731 (I171169_rst,I5701);
not I_9732 (I171186,I143244);
nor I_9733 (I171203,I143220,I143226);
nand I_9734 (I171220,I171203,I143229);
DFFARX1 I_9735  ( .D(I171220), .CLK(I5694_clk), .RSTB(I171169_rst), .Q(I171143) );
nor I_9736 (I171251,I171186,I143220);
nand I_9737 (I171268,I171251,I143238);
not I_9738 (I171158,I171268);
DFFARX1 I_9739  ( .D(I171268), .CLK(I5694_clk), .RSTB(I171169_rst), .Q(I171140) );
not I_9740 (I171313,I143220);
not I_9741 (I171330,I171313);
not I_9742 (I171347,I143217);
nor I_9743 (I171364,I171347,I143232);
and I_9744 (I171381,I171364,I143223);
or I_9745 (I171398,I171381,I143235);
DFFARX1 I_9746  ( .D(I171398), .CLK(I5694_clk), .RSTB(I171169_rst), .Q(I171415) );
nor I_9747 (I171432,I171415,I171268);
nor I_9748 (I171449,I171415,I171330);
nand I_9749 (I171155,I171220,I171449);
nand I_9750 (I171480,I171186,I143217);
nand I_9751 (I171497,I171480,I171415);
and I_9752 (I171514,I171480,I171497);
DFFARX1 I_9753  ( .D(I171514), .CLK(I5694_clk), .RSTB(I171169_rst), .Q(I171137) );
DFFARX1 I_9754  ( .D(I171480), .CLK(I5694_clk), .RSTB(I171169_rst), .Q(I171545) );
and I_9755 (I171134,I171313,I171545);
DFFARX1 I_9756  ( .D(I143247), .CLK(I5694_clk), .RSTB(I171169_rst), .Q(I171576) );
not I_9757 (I171593,I171576);
nor I_9758 (I171610,I171268,I171593);
and I_9759 (I171627,I171576,I171610);
nand I_9760 (I171149,I171576,I171330);
DFFARX1 I_9761  ( .D(I171576), .CLK(I5694_clk), .RSTB(I171169_rst), .Q(I171658) );
not I_9762 (I171146,I171658);
DFFARX1 I_9763  ( .D(I143241), .CLK(I5694_clk), .RSTB(I171169_rst), .Q(I171689) );
not I_9764 (I171706,I171689);
or I_9765 (I171723,I171706,I171627);
DFFARX1 I_9766  ( .D(I171723), .CLK(I5694_clk), .RSTB(I171169_rst), .Q(I171152) );
nand I_9767 (I171161,I171706,I171432);
DFFARX1 I_9768  ( .D(I171706), .CLK(I5694_clk), .RSTB(I171169_rst), .Q(I171131) );
not I_9769 (I171815_rst,I5701);
not I_9770 (I171832,I122359);
nor I_9771 (I171849,I122356,I122344);
nand I_9772 (I171866,I171849,I122347);
DFFARX1 I_9773  ( .D(I171866), .CLK(I5694_clk), .RSTB(I171815_rst), .Q(I171789) );
nor I_9774 (I171897,I171832,I122356);
nand I_9775 (I171914,I171897,I122353);
not I_9776 (I171804,I171914);
DFFARX1 I_9777  ( .D(I171914), .CLK(I5694_clk), .RSTB(I171815_rst), .Q(I171786) );
not I_9778 (I171959,I122356);
not I_9779 (I171976,I171959);
not I_9780 (I171993,I122365);
nor I_9781 (I172010,I171993,I122341);
and I_9782 (I172027,I172010,I122362);
or I_9783 (I172044,I172027,I122350);
DFFARX1 I_9784  ( .D(I172044), .CLK(I5694_clk), .RSTB(I171815_rst), .Q(I172061) );
nor I_9785 (I172078,I172061,I171914);
nor I_9786 (I172095,I172061,I171976);
nand I_9787 (I171801,I171866,I172095);
nand I_9788 (I172126,I171832,I122365);
nand I_9789 (I172143,I172126,I172061);
and I_9790 (I172160,I172126,I172143);
DFFARX1 I_9791  ( .D(I172160), .CLK(I5694_clk), .RSTB(I171815_rst), .Q(I171783) );
DFFARX1 I_9792  ( .D(I172126), .CLK(I5694_clk), .RSTB(I171815_rst), .Q(I172191) );
and I_9793 (I171780,I171959,I172191);
DFFARX1 I_9794  ( .D(I122371), .CLK(I5694_clk), .RSTB(I171815_rst), .Q(I172222) );
not I_9795 (I172239,I172222);
nor I_9796 (I172256,I171914,I172239);
and I_9797 (I172273,I172222,I172256);
nand I_9798 (I171795,I172222,I171976);
DFFARX1 I_9799  ( .D(I172222), .CLK(I5694_clk), .RSTB(I171815_rst), .Q(I172304) );
not I_9800 (I171792,I172304);
DFFARX1 I_9801  ( .D(I122368), .CLK(I5694_clk), .RSTB(I171815_rst), .Q(I172335) );
not I_9802 (I172352,I172335);
or I_9803 (I172369,I172352,I172273);
DFFARX1 I_9804  ( .D(I172369), .CLK(I5694_clk), .RSTB(I171815_rst), .Q(I171798) );
nand I_9805 (I171807,I172352,I172078);
DFFARX1 I_9806  ( .D(I172352), .CLK(I5694_clk), .RSTB(I171815_rst), .Q(I171777) );
not I_9807 (I172461_rst,I5701);
not I_9808 (I172478,I153332);
nor I_9809 (I172495,I153347,I153362);
nand I_9810 (I172512,I172495,I153350);
DFFARX1 I_9811  ( .D(I172512), .CLK(I5694_clk), .RSTB(I172461_rst), .Q(I172435) );
nor I_9812 (I172543,I172478,I153347);
nand I_9813 (I172560,I172543,I153353);
not I_9814 (I172450,I172560);
DFFARX1 I_9815  ( .D(I172560), .CLK(I5694_clk), .RSTB(I172461_rst), .Q(I172432) );
not I_9816 (I172605,I153347);
not I_9817 (I172622,I172605);
not I_9818 (I172639,I153359);
nor I_9819 (I172656,I172639,I153356);
and I_9820 (I172673,I172656,I153335);
or I_9821 (I172690,I172673,I153344);
DFFARX1 I_9822  ( .D(I172690), .CLK(I5694_clk), .RSTB(I172461_rst), .Q(I172707) );
nor I_9823 (I172724,I172707,I172560);
nor I_9824 (I172741,I172707,I172622);
nand I_9825 (I172447,I172512,I172741);
nand I_9826 (I172772,I172478,I153359);
nand I_9827 (I172789,I172772,I172707);
and I_9828 (I172806,I172772,I172789);
DFFARX1 I_9829  ( .D(I172806), .CLK(I5694_clk), .RSTB(I172461_rst), .Q(I172429) );
DFFARX1 I_9830  ( .D(I172772), .CLK(I5694_clk), .RSTB(I172461_rst), .Q(I172837) );
and I_9831 (I172426,I172605,I172837);
DFFARX1 I_9832  ( .D(I153341), .CLK(I5694_clk), .RSTB(I172461_rst), .Q(I172868) );
not I_9833 (I172885,I172868);
nor I_9834 (I172902,I172560,I172885);
and I_9835 (I172919,I172868,I172902);
nand I_9836 (I172441,I172868,I172622);
DFFARX1 I_9837  ( .D(I172868), .CLK(I5694_clk), .RSTB(I172461_rst), .Q(I172950) );
not I_9838 (I172438,I172950);
DFFARX1 I_9839  ( .D(I153338), .CLK(I5694_clk), .RSTB(I172461_rst), .Q(I172981) );
not I_9840 (I172998,I172981);
or I_9841 (I173015,I172998,I172919);
DFFARX1 I_9842  ( .D(I173015), .CLK(I5694_clk), .RSTB(I172461_rst), .Q(I172444) );
nand I_9843 (I172453,I172998,I172724);
DFFARX1 I_9844  ( .D(I172998), .CLK(I5694_clk), .RSTB(I172461_rst), .Q(I172423) );
not I_9845 (I173107_rst,I5701);
not I_9846 (I173124,I121033);
nor I_9847 (I173141,I121030,I121018);
nand I_9848 (I173158,I173141,I121021);
DFFARX1 I_9849  ( .D(I173158), .CLK(I5694_clk), .RSTB(I173107_rst), .Q(I173081) );
nor I_9850 (I173189,I173124,I121030);
nand I_9851 (I173206,I173189,I121027);
not I_9852 (I173096,I173206);
DFFARX1 I_9853  ( .D(I173206), .CLK(I5694_clk), .RSTB(I173107_rst), .Q(I173078) );
not I_9854 (I173251,I121030);
not I_9855 (I173268,I173251);
not I_9856 (I173285,I121039);
nor I_9857 (I173302,I173285,I121015);
and I_9858 (I173319,I173302,I121036);
or I_9859 (I173336,I173319,I121024);
DFFARX1 I_9860  ( .D(I173336), .CLK(I5694_clk), .RSTB(I173107_rst), .Q(I173353) );
nor I_9861 (I173370,I173353,I173206);
nor I_9862 (I173387,I173353,I173268);
nand I_9863 (I173093,I173158,I173387);
nand I_9864 (I173418,I173124,I121039);
nand I_9865 (I173435,I173418,I173353);
and I_9866 (I173452,I173418,I173435);
DFFARX1 I_9867  ( .D(I173452), .CLK(I5694_clk), .RSTB(I173107_rst), .Q(I173075) );
DFFARX1 I_9868  ( .D(I173418), .CLK(I5694_clk), .RSTB(I173107_rst), .Q(I173483) );
and I_9869 (I173072,I173251,I173483);
DFFARX1 I_9870  ( .D(I121045), .CLK(I5694_clk), .RSTB(I173107_rst), .Q(I173514) );
not I_9871 (I173531,I173514);
nor I_9872 (I173548,I173206,I173531);
and I_9873 (I173565,I173514,I173548);
nand I_9874 (I173087,I173514,I173268);
DFFARX1 I_9875  ( .D(I173514), .CLK(I5694_clk), .RSTB(I173107_rst), .Q(I173596) );
not I_9876 (I173084,I173596);
DFFARX1 I_9877  ( .D(I121042), .CLK(I5694_clk), .RSTB(I173107_rst), .Q(I173627) );
not I_9878 (I173644,I173627);
or I_9879 (I173661,I173644,I173565);
DFFARX1 I_9880  ( .D(I173661), .CLK(I5694_clk), .RSTB(I173107_rst), .Q(I173090) );
nand I_9881 (I173099,I173644,I173370);
DFFARX1 I_9882  ( .D(I173644), .CLK(I5694_clk), .RSTB(I173107_rst), .Q(I173069) );
not I_9883 (I173753_rst,I5701);
not I_9884 (I173770,I153973);
nor I_9885 (I173787,I153979,I153991);
nand I_9886 (I173804,I173787,I153982);
DFFARX1 I_9887  ( .D(I173804), .CLK(I5694_clk), .RSTB(I173753_rst), .Q(I173724) );
nor I_9888 (I173835,I173770,I153979);
nand I_9889 (I173852,I173835,I153961);
nand I_9890 (I173869,I173852,I173804);
not I_9891 (I173886,I153979);
not I_9892 (I173903,I153976);
nor I_9893 (I173920,I173903,I153964);
and I_9894 (I173937,I173920,I153985);
or I_9895 (I173954,I173937,I153967);
DFFARX1 I_9896  ( .D(I173954), .CLK(I5694_clk), .RSTB(I173753_rst), .Q(I173971) );
nor I_9897 (I173988,I173971,I173852);
nand I_9898 (I173739,I173886,I173988);
not I_9899 (I173736,I173971);
and I_9900 (I174033,I173971,I173869);
DFFARX1 I_9901  ( .D(I174033), .CLK(I5694_clk), .RSTB(I173753_rst), .Q(I173721) );
DFFARX1 I_9902  ( .D(I173971), .CLK(I5694_clk), .RSTB(I173753_rst), .Q(I174064) );
and I_9903 (I173718,I173886,I174064);
nand I_9904 (I174095,I173770,I153976);
not I_9905 (I174112,I174095);
nor I_9906 (I174129,I173971,I174112);
DFFARX1 I_9907  ( .D(I153988), .CLK(I5694_clk), .RSTB(I173753_rst), .Q(I174146) );
nand I_9908 (I174163,I174146,I174095);
and I_9909 (I174180,I173886,I174163);
DFFARX1 I_9910  ( .D(I174180), .CLK(I5694_clk), .RSTB(I173753_rst), .Q(I173745) );
not I_9911 (I174211,I174146);
nand I_9912 (I173733,I174146,I174129);
nand I_9913 (I173727,I174146,I174112);
DFFARX1 I_9914  ( .D(I153970), .CLK(I5694_clk), .RSTB(I173753_rst), .Q(I174256) );
not I_9915 (I174273,I174256);
nor I_9916 (I173742,I174146,I174273);
nor I_9917 (I174304,I174273,I174211);
and I_9918 (I174321,I173852,I174304);
or I_9919 (I174338,I174095,I174321);
DFFARX1 I_9920  ( .D(I174338), .CLK(I5694_clk), .RSTB(I173753_rst), .Q(I173730) );
DFFARX1 I_9921  ( .D(I174273), .CLK(I5694_clk), .RSTB(I173753_rst), .Q(I173715) );
not I_9922 (I174416_rst,I5701);
not I_9923 (I174433,I173084);
nor I_9924 (I174450,I173072,I173096);
nand I_9925 (I174467,I174450,I173081);
DFFARX1 I_9926  ( .D(I174467), .CLK(I5694_clk), .RSTB(I174416_rst), .Q(I174387) );
nor I_9927 (I174498,I174433,I173072);
nand I_9928 (I174515,I174498,I173099);
nand I_9929 (I174532,I174515,I174467);
not I_9930 (I174549,I173072);
not I_9931 (I174566,I173069);
nor I_9932 (I174583,I174566,I173078);
and I_9933 (I174600,I174583,I173093);
or I_9934 (I174617,I174600,I173075);
DFFARX1 I_9935  ( .D(I174617), .CLK(I5694_clk), .RSTB(I174416_rst), .Q(I174634) );
nor I_9936 (I174651,I174634,I174515);
nand I_9937 (I174402,I174549,I174651);
not I_9938 (I174399,I174634);
and I_9939 (I174696,I174634,I174532);
DFFARX1 I_9940  ( .D(I174696), .CLK(I5694_clk), .RSTB(I174416_rst), .Q(I174384) );
DFFARX1 I_9941  ( .D(I174634), .CLK(I5694_clk), .RSTB(I174416_rst), .Q(I174727) );
and I_9942 (I174381,I174549,I174727);
nand I_9943 (I174758,I174433,I173069);
not I_9944 (I174775,I174758);
nor I_9945 (I174792,I174634,I174775);
DFFARX1 I_9946  ( .D(I173090), .CLK(I5694_clk), .RSTB(I174416_rst), .Q(I174809) );
nand I_9947 (I174826,I174809,I174758);
and I_9948 (I174843,I174549,I174826);
DFFARX1 I_9949  ( .D(I174843), .CLK(I5694_clk), .RSTB(I174416_rst), .Q(I174408) );
not I_9950 (I174874,I174809);
nand I_9951 (I174396,I174809,I174792);
nand I_9952 (I174390,I174809,I174775);
DFFARX1 I_9953  ( .D(I173087), .CLK(I5694_clk), .RSTB(I174416_rst), .Q(I174919) );
not I_9954 (I174936,I174919);
nor I_9955 (I174405,I174809,I174936);
nor I_9956 (I174967,I174936,I174874);
and I_9957 (I174984,I174515,I174967);
or I_9958 (I175001,I174758,I174984);
DFFARX1 I_9959  ( .D(I175001), .CLK(I5694_clk), .RSTB(I174416_rst), .Q(I174393) );
DFFARX1 I_9960  ( .D(I174936), .CLK(I5694_clk), .RSTB(I174416_rst), .Q(I174378) );
not I_9961 (I175079_rst,I5701);
not I_9962 (I175096,I121678);
nor I_9963 (I175113,I121687,I121699);
nand I_9964 (I175130,I175113,I121690);
DFFARX1 I_9965  ( .D(I175130), .CLK(I5694_clk), .RSTB(I175079_rst), .Q(I175050) );
nor I_9966 (I175161,I175096,I121687);
nand I_9967 (I175178,I175161,I121702);
nand I_9968 (I175195,I175178,I175130);
not I_9969 (I175212,I121687);
not I_9970 (I175229,I121708);
nor I_9971 (I175246,I175229,I121684);
and I_9972 (I175263,I175246,I121693);
or I_9973 (I175280,I175263,I121681);
DFFARX1 I_9974  ( .D(I175280), .CLK(I5694_clk), .RSTB(I175079_rst), .Q(I175297) );
nor I_9975 (I175314,I175297,I175178);
nand I_9976 (I175065,I175212,I175314);
not I_9977 (I175062,I175297);
and I_9978 (I175359,I175297,I175195);
DFFARX1 I_9979  ( .D(I175359), .CLK(I5694_clk), .RSTB(I175079_rst), .Q(I175047) );
DFFARX1 I_9980  ( .D(I175297), .CLK(I5694_clk), .RSTB(I175079_rst), .Q(I175390) );
and I_9981 (I175044,I175212,I175390);
nand I_9982 (I175421,I175096,I121708);
not I_9983 (I175438,I175421);
nor I_9984 (I175455,I175297,I175438);
DFFARX1 I_9985  ( .D(I121705), .CLK(I5694_clk), .RSTB(I175079_rst), .Q(I175472) );
nand I_9986 (I175489,I175472,I175421);
and I_9987 (I175506,I175212,I175489);
DFFARX1 I_9988  ( .D(I175506), .CLK(I5694_clk), .RSTB(I175079_rst), .Q(I175071) );
not I_9989 (I175537,I175472);
nand I_9990 (I175059,I175472,I175455);
nand I_9991 (I175053,I175472,I175438);
DFFARX1 I_9992  ( .D(I121696), .CLK(I5694_clk), .RSTB(I175079_rst), .Q(I175582) );
not I_9993 (I175599,I175582);
nor I_9994 (I175068,I175472,I175599);
nor I_9995 (I175630,I175599,I175537);
and I_9996 (I175647,I175178,I175630);
or I_9997 (I175664,I175421,I175647);
DFFARX1 I_9998  ( .D(I175664), .CLK(I5694_clk), .RSTB(I175079_rst), .Q(I175056) );
DFFARX1 I_9999  ( .D(I175599), .CLK(I5694_clk), .RSTB(I175079_rst), .Q(I175041) );
not I_10000 (I175742_rst,I5701);
not I_10001 (I175759,I130247);
nor I_10002 (I175776,I130256,I130229);
nand I_10003 (I175793,I175776,I130241);
DFFARX1 I_10004  ( .D(I175793), .CLK(I5694_clk), .RSTB(I175742_rst), .Q(I175713) );
nor I_10005 (I175824,I175759,I130256);
nand I_10006 (I175841,I175824,I130253);
nand I_10007 (I175858,I175841,I175793);
not I_10008 (I175875,I130256);
not I_10009 (I175892,I130232);
nor I_10010 (I175909,I175892,I130238);
and I_10011 (I175926,I175909,I130250);
or I_10012 (I175943,I175926,I130235);
DFFARX1 I_10013  ( .D(I175943), .CLK(I5694_clk), .RSTB(I175742_rst), .Q(I175960) );
nor I_10014 (I175977,I175960,I175841);
nand I_10015 (I175728,I175875,I175977);
not I_10016 (I175725,I175960);
and I_10017 (I176022,I175960,I175858);
DFFARX1 I_10018  ( .D(I176022), .CLK(I5694_clk), .RSTB(I175742_rst), .Q(I175710) );
DFFARX1 I_10019  ( .D(I175960), .CLK(I5694_clk), .RSTB(I175742_rst), .Q(I176053) );
and I_10020 (I175707,I175875,I176053);
nand I_10021 (I176084,I175759,I130232);
not I_10022 (I176101,I176084);
nor I_10023 (I176118,I175960,I176101);
DFFARX1 I_10024  ( .D(I130259), .CLK(I5694_clk), .RSTB(I175742_rst), .Q(I176135) );
nand I_10025 (I176152,I176135,I176084);
and I_10026 (I176169,I175875,I176152);
DFFARX1 I_10027  ( .D(I176169), .CLK(I5694_clk), .RSTB(I175742_rst), .Q(I175734) );
not I_10028 (I176200,I176135);
nand I_10029 (I175722,I176135,I176118);
nand I_10030 (I175716,I176135,I176101);
DFFARX1 I_10031  ( .D(I130244), .CLK(I5694_clk), .RSTB(I175742_rst), .Q(I176245) );
not I_10032 (I176262,I176245);
nor I_10033 (I175731,I176135,I176262);
nor I_10034 (I176293,I176262,I176200);
and I_10035 (I176310,I175841,I176293);
or I_10036 (I176327,I176084,I176310);
DFFARX1 I_10037  ( .D(I176327), .CLK(I5694_clk), .RSTB(I175742_rst), .Q(I175719) );
DFFARX1 I_10038  ( .D(I176262), .CLK(I5694_clk), .RSTB(I175742_rst), .Q(I175704) );
not I_10039 (I176405_rst,I5701);
not I_10040 (I176422,I163003);
nor I_10041 (I176439,I162991,I162994);
nand I_10042 (I176456,I176439,I163009);
DFFARX1 I_10043  ( .D(I176456), .CLK(I5694_clk), .RSTB(I176405_rst), .Q(I176376) );
nor I_10044 (I176487,I176422,I162991);
nand I_10045 (I176504,I176487,I163000);
nand I_10046 (I176521,I176504,I176456);
not I_10047 (I176538,I162991);
not I_10048 (I176555,I163012);
nor I_10049 (I176572,I176555,I162988);
and I_10050 (I176589,I176572,I162997);
or I_10051 (I176606,I176589,I163006);
DFFARX1 I_10052  ( .D(I176606), .CLK(I5694_clk), .RSTB(I176405_rst), .Q(I176623) );
nor I_10053 (I176640,I176623,I176504);
nand I_10054 (I176391,I176538,I176640);
not I_10055 (I176388,I176623);
and I_10056 (I176685,I176623,I176521);
DFFARX1 I_10057  ( .D(I176685), .CLK(I5694_clk), .RSTB(I176405_rst), .Q(I176373) );
DFFARX1 I_10058  ( .D(I176623), .CLK(I5694_clk), .RSTB(I176405_rst), .Q(I176716) );
and I_10059 (I176370,I176538,I176716);
nand I_10060 (I176747,I176422,I163012);
not I_10061 (I176764,I176747);
nor I_10062 (I176781,I176623,I176764);
DFFARX1 I_10063  ( .D(I163018), .CLK(I5694_clk), .RSTB(I176405_rst), .Q(I176798) );
nand I_10064 (I176815,I176798,I176747);
and I_10065 (I176832,I176538,I176815);
DFFARX1 I_10066  ( .D(I176832), .CLK(I5694_clk), .RSTB(I176405_rst), .Q(I176397) );
not I_10067 (I176863,I176798);
nand I_10068 (I176385,I176798,I176781);
nand I_10069 (I176379,I176798,I176764);
DFFARX1 I_10070  ( .D(I163015), .CLK(I5694_clk), .RSTB(I176405_rst), .Q(I176908) );
not I_10071 (I176925,I176908);
nor I_10072 (I176394,I176798,I176925);
nor I_10073 (I176956,I176925,I176863);
and I_10074 (I176973,I176504,I176956);
or I_10075 (I176990,I176747,I176973);
DFFARX1 I_10076  ( .D(I176990), .CLK(I5694_clk), .RSTB(I176405_rst), .Q(I176382) );
DFFARX1 I_10077  ( .D(I176925), .CLK(I5694_clk), .RSTB(I176405_rst), .Q(I176367) );
not I_10078 (I177068_rst,I5701);
not I_10079 (I177085,I136061);
nor I_10080 (I177102,I136070,I136043);
nand I_10081 (I177119,I177102,I136055);
DFFARX1 I_10082  ( .D(I177119), .CLK(I5694_clk), .RSTB(I177068_rst), .Q(I177039) );
nor I_10083 (I177150,I177085,I136070);
nand I_10084 (I177167,I177150,I136067);
nand I_10085 (I177184,I177167,I177119);
not I_10086 (I177201,I136070);
not I_10087 (I177218,I136046);
nor I_10088 (I177235,I177218,I136052);
and I_10089 (I177252,I177235,I136064);
or I_10090 (I177269,I177252,I136049);
DFFARX1 I_10091  ( .D(I177269), .CLK(I5694_clk), .RSTB(I177068_rst), .Q(I177286) );
nor I_10092 (I177303,I177286,I177167);
nand I_10093 (I177054,I177201,I177303);
not I_10094 (I177051,I177286);
and I_10095 (I177348,I177286,I177184);
DFFARX1 I_10096  ( .D(I177348), .CLK(I5694_clk), .RSTB(I177068_rst), .Q(I177036) );
DFFARX1 I_10097  ( .D(I177286), .CLK(I5694_clk), .RSTB(I177068_rst), .Q(I177379) );
and I_10098 (I177033,I177201,I177379);
nand I_10099 (I177410,I177085,I136046);
not I_10100 (I177427,I177410);
nor I_10101 (I177444,I177286,I177427);
DFFARX1 I_10102  ( .D(I136073), .CLK(I5694_clk), .RSTB(I177068_rst), .Q(I177461) );
nand I_10103 (I177478,I177461,I177410);
and I_10104 (I177495,I177201,I177478);
DFFARX1 I_10105  ( .D(I177495), .CLK(I5694_clk), .RSTB(I177068_rst), .Q(I177060) );
not I_10106 (I177526,I177461);
nand I_10107 (I177048,I177461,I177444);
nand I_10108 (I177042,I177461,I177427);
DFFARX1 I_10109  ( .D(I136058), .CLK(I5694_clk), .RSTB(I177068_rst), .Q(I177571) );
not I_10110 (I177588,I177571);
nor I_10111 (I177057,I177461,I177588);
nor I_10112 (I177619,I177588,I177526);
and I_10113 (I177636,I177167,I177619);
or I_10114 (I177653,I177410,I177636);
DFFARX1 I_10115  ( .D(I177653), .CLK(I5694_clk), .RSTB(I177068_rst), .Q(I177045) );
DFFARX1 I_10116  ( .D(I177588), .CLK(I5694_clk), .RSTB(I177068_rst), .Q(I177030) );
not I_10117 (I177731_rst,I5701);
not I_10118 (I177748,I150958);
nor I_10119 (I177765,I150973,I150955);
nand I_10120 (I177782,I177765,I150967);
DFFARX1 I_10121  ( .D(I177782), .CLK(I5694_clk), .RSTB(I177731_rst), .Q(I177702) );
nor I_10122 (I177813,I177748,I150973);
nand I_10123 (I177830,I177813,I150964);
nand I_10124 (I177847,I177830,I177782);
not I_10125 (I177864,I150973);
not I_10126 (I177881,I150982);
nor I_10127 (I177898,I177881,I150952);
and I_10128 (I177915,I177898,I150961);
or I_10129 (I177932,I177915,I150979);
DFFARX1 I_10130  ( .D(I177932), .CLK(I5694_clk), .RSTB(I177731_rst), .Q(I177949) );
nor I_10131 (I177966,I177949,I177830);
nand I_10132 (I177717,I177864,I177966);
not I_10133 (I177714,I177949);
and I_10134 (I178011,I177949,I177847);
DFFARX1 I_10135  ( .D(I178011), .CLK(I5694_clk), .RSTB(I177731_rst), .Q(I177699) );
DFFARX1 I_10136  ( .D(I177949), .CLK(I5694_clk), .RSTB(I177731_rst), .Q(I178042) );
and I_10137 (I177696,I177864,I178042);
nand I_10138 (I178073,I177748,I150982);
not I_10139 (I178090,I178073);
nor I_10140 (I178107,I177949,I178090);
DFFARX1 I_10141  ( .D(I150970), .CLK(I5694_clk), .RSTB(I177731_rst), .Q(I178124) );
nand I_10142 (I178141,I178124,I178073);
and I_10143 (I178158,I177864,I178141);
DFFARX1 I_10144  ( .D(I178158), .CLK(I5694_clk), .RSTB(I177731_rst), .Q(I177723) );
not I_10145 (I178189,I178124);
nand I_10146 (I177711,I178124,I178107);
nand I_10147 (I177705,I178124,I178090);
DFFARX1 I_10148  ( .D(I150976), .CLK(I5694_clk), .RSTB(I177731_rst), .Q(I178234) );
not I_10149 (I178251,I178234);
nor I_10150 (I177720,I178124,I178251);
nor I_10151 (I178282,I178251,I178189);
and I_10152 (I178299,I177830,I178282);
or I_10153 (I178316,I178073,I178299);
DFFARX1 I_10154  ( .D(I178316), .CLK(I5694_clk), .RSTB(I177731_rst), .Q(I177708) );
DFFARX1 I_10155  ( .D(I178251), .CLK(I5694_clk), .RSTB(I177731_rst), .Q(I177693) );
not I_10156 (I178394_rst,I5701);
not I_10157 (I178411,I146802);
nor I_10158 (I178428,I146814,I146817);
nand I_10159 (I178445,I178428,I146805);
DFFARX1 I_10160  ( .D(I178445), .CLK(I5694_clk), .RSTB(I178394_rst), .Q(I178365) );
nor I_10161 (I178476,I178411,I146814);
nand I_10162 (I178493,I178476,I146790);
nand I_10163 (I178510,I178493,I178445);
not I_10164 (I178527,I146814);
not I_10165 (I178544,I146793);
nor I_10166 (I178561,I178544,I146796);
and I_10167 (I178578,I178561,I146799);
or I_10168 (I178595,I178578,I146808);
DFFARX1 I_10169  ( .D(I178595), .CLK(I5694_clk), .RSTB(I178394_rst), .Q(I178612) );
nor I_10170 (I178629,I178612,I178493);
nand I_10171 (I178380,I178527,I178629);
not I_10172 (I178377,I178612);
and I_10173 (I178674,I178612,I178510);
DFFARX1 I_10174  ( .D(I178674), .CLK(I5694_clk), .RSTB(I178394_rst), .Q(I178362) );
DFFARX1 I_10175  ( .D(I178612), .CLK(I5694_clk), .RSTB(I178394_rst), .Q(I178705) );
and I_10176 (I178359,I178527,I178705);
nand I_10177 (I178736,I178411,I146793);
not I_10178 (I178753,I178736);
nor I_10179 (I178770,I178612,I178753);
DFFARX1 I_10180  ( .D(I146811), .CLK(I5694_clk), .RSTB(I178394_rst), .Q(I178787) );
nand I_10181 (I178804,I178787,I178736);
and I_10182 (I178821,I178527,I178804);
DFFARX1 I_10183  ( .D(I178821), .CLK(I5694_clk), .RSTB(I178394_rst), .Q(I178386) );
not I_10184 (I178852,I178787);
nand I_10185 (I178374,I178787,I178770);
nand I_10186 (I178368,I178787,I178753);
DFFARX1 I_10187  ( .D(I146787), .CLK(I5694_clk), .RSTB(I178394_rst), .Q(I178897) );
not I_10188 (I178914,I178897);
nor I_10189 (I178383,I178787,I178914);
nor I_10190 (I178945,I178914,I178852);
and I_10191 (I178962,I178493,I178945);
or I_10192 (I178979,I178736,I178962);
DFFARX1 I_10193  ( .D(I178979), .CLK(I5694_clk), .RSTB(I178394_rst), .Q(I178371) );
DFFARX1 I_10194  ( .D(I178914), .CLK(I5694_clk), .RSTB(I178394_rst), .Q(I178356) );
not I_10195 (I179057_rst,I5701);
not I_10196 (I179074,I152148);
nor I_10197 (I179091,I152163,I152145);
nand I_10198 (I179108,I179091,I152157);
DFFARX1 I_10199  ( .D(I179108), .CLK(I5694_clk), .RSTB(I179057_rst), .Q(I179028) );
nor I_10200 (I179139,I179074,I152163);
nand I_10201 (I179156,I179139,I152154);
nand I_10202 (I179173,I179156,I179108);
not I_10203 (I179190,I152163);
not I_10204 (I179207,I152172);
nor I_10205 (I179224,I179207,I152142);
and I_10206 (I179241,I179224,I152151);
or I_10207 (I179258,I179241,I152169);
DFFARX1 I_10208  ( .D(I179258), .CLK(I5694_clk), .RSTB(I179057_rst), .Q(I179275) );
nor I_10209 (I179292,I179275,I179156);
nand I_10210 (I179043,I179190,I179292);
not I_10211 (I179040,I179275);
and I_10212 (I179337,I179275,I179173);
DFFARX1 I_10213  ( .D(I179337), .CLK(I5694_clk), .RSTB(I179057_rst), .Q(I179025) );
DFFARX1 I_10214  ( .D(I179275), .CLK(I5694_clk), .RSTB(I179057_rst), .Q(I179368) );
and I_10215 (I179022,I179190,I179368);
nand I_10216 (I179399,I179074,I152172);
not I_10217 (I179416,I179399);
nor I_10218 (I179433,I179275,I179416);
DFFARX1 I_10219  ( .D(I152160), .CLK(I5694_clk), .RSTB(I179057_rst), .Q(I179450) );
nand I_10220 (I179467,I179450,I179399);
and I_10221 (I179484,I179190,I179467);
DFFARX1 I_10222  ( .D(I179484), .CLK(I5694_clk), .RSTB(I179057_rst), .Q(I179049) );
not I_10223 (I179515,I179450);
nand I_10224 (I179037,I179450,I179433);
nand I_10225 (I179031,I179450,I179416);
DFFARX1 I_10226  ( .D(I152166), .CLK(I5694_clk), .RSTB(I179057_rst), .Q(I179560) );
not I_10227 (I179577,I179560);
nor I_10228 (I179046,I179450,I179577);
nor I_10229 (I179608,I179577,I179515);
and I_10230 (I179625,I179156,I179608);
or I_10231 (I179642,I179399,I179625);
DFFARX1 I_10232  ( .D(I179642), .CLK(I5694_clk), .RSTB(I179057_rst), .Q(I179034) );
DFFARX1 I_10233  ( .D(I179577), .CLK(I5694_clk), .RSTB(I179057_rst), .Q(I179019) );
not I_10234 (I179720_rst,I5701);
or I_10235 (I179737,I159571,I159589);
or I_10236 (I179754,I159574,I159571);
DFFARX1 I_10237  ( .D(I179754), .CLK(I5694_clk), .RSTB(I179720_rst), .Q(I179694) );
nor I_10238 (I179785,I159583,I159586);
not I_10239 (I179802,I179785);
not I_10240 (I179819,I159583);
and I_10241 (I179836,I179819,I159592);
nor I_10242 (I179853,I179836,I159589);
nor I_10243 (I179870,I159598,I159577);
DFFARX1 I_10244  ( .D(I179870), .CLK(I5694_clk), .RSTB(I179720_rst), .Q(I179887) );
nand I_10245 (I179904,I179887,I179737);
and I_10246 (I179921,I179853,I179904);
DFFARX1 I_10247  ( .D(I179921), .CLK(I5694_clk), .RSTB(I179720_rst), .Q(I179688) );
nor I_10248 (I179952,I159598,I159574);
DFFARX1 I_10249  ( .D(I179952), .CLK(I5694_clk), .RSTB(I179720_rst), .Q(I179969) );
and I_10250 (I179685,I179785,I179969);
DFFARX1 I_10251  ( .D(I159601), .CLK(I5694_clk), .RSTB(I179720_rst), .Q(I180000) );
and I_10252 (I180017,I180000,I159595);
DFFARX1 I_10253  ( .D(I180017), .CLK(I5694_clk), .RSTB(I179720_rst), .Q(I180034) );
not I_10254 (I179697,I180034);
DFFARX1 I_10255  ( .D(I180017), .CLK(I5694_clk), .RSTB(I179720_rst), .Q(I179682) );
DFFARX1 I_10256  ( .D(I159580), .CLK(I5694_clk), .RSTB(I179720_rst), .Q(I180079) );
not I_10257 (I180096,I180079);
nor I_10258 (I180113,I179754,I180096);
and I_10259 (I180130,I180017,I180113);
or I_10260 (I180147,I179737,I180130);
DFFARX1 I_10261  ( .D(I180147), .CLK(I5694_clk), .RSTB(I179720_rst), .Q(I179703) );
nor I_10262 (I180178,I180079,I179887);
nand I_10263 (I179712,I179853,I180178);
nor I_10264 (I180209,I180079,I179802);
nand I_10265 (I179706,I179952,I180209);
not I_10266 (I179709,I180079);
nand I_10267 (I179700,I180079,I179802);
DFFARX1 I_10268  ( .D(I180079), .CLK(I5694_clk), .RSTB(I179720_rst), .Q(I179691) );
not I_10269 (I180315_rst,I5701);
or I_10270 (I180332,I165984,I165978);
or I_10271 (I180349,I165972,I165984);
DFFARX1 I_10272  ( .D(I180349), .CLK(I5694_clk), .RSTB(I180315_rst), .Q(I180289) );
nor I_10273 (I180380,I165990,I165981);
not I_10274 (I180397,I180380);
not I_10275 (I180414,I165990);
and I_10276 (I180431,I180414,I165987);
nor I_10277 (I180448,I180431,I165978);
nor I_10278 (I180465,I165963,I165969);
DFFARX1 I_10279  ( .D(I180465), .CLK(I5694_clk), .RSTB(I180315_rst), .Q(I180482) );
nand I_10280 (I180499,I180482,I180332);
and I_10281 (I180516,I180448,I180499);
DFFARX1 I_10282  ( .D(I180516), .CLK(I5694_clk), .RSTB(I180315_rst), .Q(I180283) );
nor I_10283 (I180547,I165963,I165972);
DFFARX1 I_10284  ( .D(I180547), .CLK(I5694_clk), .RSTB(I180315_rst), .Q(I180564) );
and I_10285 (I180280,I180380,I180564);
DFFARX1 I_10286  ( .D(I165975), .CLK(I5694_clk), .RSTB(I180315_rst), .Q(I180595) );
and I_10287 (I180612,I180595,I165993);
DFFARX1 I_10288  ( .D(I180612), .CLK(I5694_clk), .RSTB(I180315_rst), .Q(I180629) );
not I_10289 (I180292,I180629);
DFFARX1 I_10290  ( .D(I180612), .CLK(I5694_clk), .RSTB(I180315_rst), .Q(I180277) );
DFFARX1 I_10291  ( .D(I165966), .CLK(I5694_clk), .RSTB(I180315_rst), .Q(I180674) );
not I_10292 (I180691,I180674);
nor I_10293 (I180708,I180349,I180691);
and I_10294 (I180725,I180612,I180708);
or I_10295 (I180742,I180332,I180725);
DFFARX1 I_10296  ( .D(I180742), .CLK(I5694_clk), .RSTB(I180315_rst), .Q(I180298) );
nor I_10297 (I180773,I180674,I180482);
nand I_10298 (I180307,I180448,I180773);
nor I_10299 (I180804,I180674,I180397);
nand I_10300 (I180301,I180547,I180804);
not I_10301 (I180304,I180674);
nand I_10302 (I180295,I180674,I180397);
DFFARX1 I_10303  ( .D(I180674), .CLK(I5694_clk), .RSTB(I180315_rst), .Q(I180286) );
not I_10304 (I180910_rst,I5701);
or I_10305 (I180927,I147992,I147977);
or I_10306 (I180944,I147998,I147992);
DFFARX1 I_10307  ( .D(I180944), .CLK(I5694_clk), .RSTB(I180910_rst), .Q(I180884) );
nor I_10308 (I180975,I148004,I147986);
not I_10309 (I180992,I180975);
not I_10310 (I181009,I148004);
and I_10311 (I181026,I181009,I147983);
nor I_10312 (I181043,I181026,I147977);
nor I_10313 (I181060,I147980,I147989);
DFFARX1 I_10314  ( .D(I181060), .CLK(I5694_clk), .RSTB(I180910_rst), .Q(I181077) );
nand I_10315 (I181094,I181077,I180927);
and I_10316 (I181111,I181043,I181094);
DFFARX1 I_10317  ( .D(I181111), .CLK(I5694_clk), .RSTB(I180910_rst), .Q(I180878) );
nor I_10318 (I181142,I147980,I147998);
DFFARX1 I_10319  ( .D(I181142), .CLK(I5694_clk), .RSTB(I180910_rst), .Q(I181159) );
and I_10320 (I180875,I180975,I181159);
DFFARX1 I_10321  ( .D(I148007), .CLK(I5694_clk), .RSTB(I180910_rst), .Q(I181190) );
and I_10322 (I181207,I181190,I147995);
DFFARX1 I_10323  ( .D(I181207), .CLK(I5694_clk), .RSTB(I180910_rst), .Q(I181224) );
not I_10324 (I180887,I181224);
DFFARX1 I_10325  ( .D(I181207), .CLK(I5694_clk), .RSTB(I180910_rst), .Q(I180872) );
DFFARX1 I_10326  ( .D(I148001), .CLK(I5694_clk), .RSTB(I180910_rst), .Q(I181269) );
not I_10327 (I181286,I181269);
nor I_10328 (I181303,I180944,I181286);
and I_10329 (I181320,I181207,I181303);
or I_10330 (I181337,I180927,I181320);
DFFARX1 I_10331  ( .D(I181337), .CLK(I5694_clk), .RSTB(I180910_rst), .Q(I180893) );
nor I_10332 (I181368,I181269,I181077);
nand I_10333 (I180902,I181043,I181368);
nor I_10334 (I181399,I181269,I180992);
nand I_10335 (I180896,I181142,I181399);
not I_10336 (I180899,I181269);
nand I_10337 (I180890,I181269,I180992);
DFFARX1 I_10338  ( .D(I181269), .CLK(I5694_clk), .RSTB(I180910_rst), .Q(I180881) );
not I_10339 (I181505_rst,I5701);
or I_10340 (I181522,I119026,I119041);
or I_10341 (I181539,I119029,I119026);
DFFARX1 I_10342  ( .D(I181539), .CLK(I5694_clk), .RSTB(I181505_rst), .Q(I181479) );
nor I_10343 (I181570,I119032,I119047);
not I_10344 (I181587,I181570);
not I_10345 (I181604,I119032);
and I_10346 (I181621,I181604,I119035);
nor I_10347 (I181638,I181621,I119041);
nor I_10348 (I181655,I119038,I119056);
DFFARX1 I_10349  ( .D(I181655), .CLK(I5694_clk), .RSTB(I181505_rst), .Q(I181672) );
nand I_10350 (I181689,I181672,I181522);
and I_10351 (I181706,I181638,I181689);
DFFARX1 I_10352  ( .D(I181706), .CLK(I5694_clk), .RSTB(I181505_rst), .Q(I181473) );
nor I_10353 (I181737,I119038,I119029);
DFFARX1 I_10354  ( .D(I181737), .CLK(I5694_clk), .RSTB(I181505_rst), .Q(I181754) );
and I_10355 (I181470,I181570,I181754);
DFFARX1 I_10356  ( .D(I119053), .CLK(I5694_clk), .RSTB(I181505_rst), .Q(I181785) );
and I_10357 (I181802,I181785,I119044);
DFFARX1 I_10358  ( .D(I181802), .CLK(I5694_clk), .RSTB(I181505_rst), .Q(I181819) );
not I_10359 (I181482,I181819);
DFFARX1 I_10360  ( .D(I181802), .CLK(I5694_clk), .RSTB(I181505_rst), .Q(I181467) );
DFFARX1 I_10361  ( .D(I119050), .CLK(I5694_clk), .RSTB(I181505_rst), .Q(I181864) );
not I_10362 (I181881,I181864);
nor I_10363 (I181898,I181539,I181881);
and I_10364 (I181915,I181802,I181898);
or I_10365 (I181932,I181522,I181915);
DFFARX1 I_10366  ( .D(I181932), .CLK(I5694_clk), .RSTB(I181505_rst), .Q(I181488) );
nor I_10367 (I181963,I181864,I181672);
nand I_10368 (I181497,I181638,I181963);
nor I_10369 (I181994,I181864,I181587);
nand I_10370 (I181491,I181737,I181994);
not I_10371 (I181494,I181864);
nand I_10372 (I181485,I181864,I181587);
DFFARX1 I_10373  ( .D(I181864), .CLK(I5694_clk), .RSTB(I181505_rst), .Q(I181476) );
not I_10374 (I182100_rst,I5701);
or I_10375 (I182117,I164689,I164686);
not I_10376 (I182083,I182117);
DFFARX1 I_10377  ( .D(I182117), .CLK(I5694_clk), .RSTB(I182100_rst), .Q(I182062) );
or I_10378 (I182162,I164680,I164689);
nor I_10379 (I182179,I164698,I164671);
nor I_10380 (I182196,I182179,I182117);
not I_10381 (I182213,I164698);
and I_10382 (I182230,I182213,I164692);
nor I_10383 (I182247,I182230,I164686);
DFFARX1 I_10384  ( .D(I182247), .CLK(I5694_clk), .RSTB(I182100_rst), .Q(I182264) );
nor I_10385 (I182281,I164674,I164701);
DFFARX1 I_10386  ( .D(I182281), .CLK(I5694_clk), .RSTB(I182100_rst), .Q(I182298) );
nor I_10387 (I182089,I182298,I182247);
not I_10388 (I182329,I182298);
nor I_10389 (I182346,I164674,I164680);
nand I_10390 (I182363,I182247,I182346);
and I_10391 (I182380,I182162,I182363);
DFFARX1 I_10392  ( .D(I182380), .CLK(I5694_clk), .RSTB(I182100_rst), .Q(I182092) );
DFFARX1 I_10393  ( .D(I164677), .CLK(I5694_clk), .RSTB(I182100_rst), .Q(I182411) );
and I_10394 (I182428,I182411,I164683);
nor I_10395 (I182445,I182428,I182329);
and I_10396 (I182462,I182346,I182445);
or I_10397 (I182479,I182179,I182462);
DFFARX1 I_10398  ( .D(I182479), .CLK(I5694_clk), .RSTB(I182100_rst), .Q(I182077) );
not I_10399 (I182510,I182428);
nor I_10400 (I182527,I182117,I182510);
nand I_10401 (I182080,I182162,I182527);
nand I_10402 (I182074,I182298,I182510);
DFFARX1 I_10403  ( .D(I182428), .CLK(I5694_clk), .RSTB(I182100_rst), .Q(I182068) );
DFFARX1 I_10404  ( .D(I164695), .CLK(I5694_clk), .RSTB(I182100_rst), .Q(I182586) );
nand I_10405 (I182086,I182586,I182196);
DFFARX1 I_10406  ( .D(I182586), .CLK(I5694_clk), .RSTB(I182100_rst), .Q(I182617) );
not I_10407 (I182071,I182617);
and I_10408 (I182065,I182586,I182264);
not I_10409 (I182695_rst,I5701);
or I_10410 (I182712,I167273,I167270);
not I_10411 (I182678,I182712);
DFFARX1 I_10412  ( .D(I182712), .CLK(I5694_clk), .RSTB(I182695_rst), .Q(I182657) );
or I_10413 (I182757,I167264,I167273);
nor I_10414 (I182774,I167282,I167255);
nor I_10415 (I182791,I182774,I182712);
not I_10416 (I182808,I167282);
and I_10417 (I182825,I182808,I167276);
nor I_10418 (I182842,I182825,I167270);
DFFARX1 I_10419  ( .D(I182842), .CLK(I5694_clk), .RSTB(I182695_rst), .Q(I182859) );
nor I_10420 (I182876,I167258,I167285);
DFFARX1 I_10421  ( .D(I182876), .CLK(I5694_clk), .RSTB(I182695_rst), .Q(I182893) );
nor I_10422 (I182684,I182893,I182842);
not I_10423 (I182924,I182893);
nor I_10424 (I182941,I167258,I167264);
nand I_10425 (I182958,I182842,I182941);
and I_10426 (I182975,I182757,I182958);
DFFARX1 I_10427  ( .D(I182975), .CLK(I5694_clk), .RSTB(I182695_rst), .Q(I182687) );
DFFARX1 I_10428  ( .D(I167261), .CLK(I5694_clk), .RSTB(I182695_rst), .Q(I183006) );
and I_10429 (I183023,I183006,I167267);
nor I_10430 (I183040,I183023,I182924);
and I_10431 (I183057,I182941,I183040);
or I_10432 (I183074,I182774,I183057);
DFFARX1 I_10433  ( .D(I183074), .CLK(I5694_clk), .RSTB(I182695_rst), .Q(I182672) );
not I_10434 (I183105,I183023);
nor I_10435 (I183122,I182712,I183105);
nand I_10436 (I182675,I182757,I183122);
nand I_10437 (I182669,I182893,I183105);
DFFARX1 I_10438  ( .D(I183023), .CLK(I5694_clk), .RSTB(I182695_rst), .Q(I182663) );
DFFARX1 I_10439  ( .D(I167279), .CLK(I5694_clk), .RSTB(I182695_rst), .Q(I183181) );
nand I_10440 (I182681,I183181,I182791);
DFFARX1 I_10441  ( .D(I183181), .CLK(I5694_clk), .RSTB(I182695_rst), .Q(I183212) );
not I_10442 (I182666,I183212);
and I_10443 (I182660,I183181,I182859);
not I_10444 (I183290_rst,I5701);
not I_10445 (I183307,I177696);
nor I_10446 (I183324,I177702,I177708);
nand I_10447 (I183341,I183324,I177711);
nor I_10448 (I183358,I183307,I177702);
nand I_10449 (I183375,I183358,I177693);
not I_10450 (I183392,I183375);
not I_10451 (I183409,I177702);
nor I_10452 (I183279,I183375,I183409);
not I_10453 (I183440,I183409);
nand I_10454 (I183264,I183375,I183440);
not I_10455 (I183471,I177705);
nor I_10456 (I183488,I183471,I177699);
and I_10457 (I183505,I183488,I177714);
or I_10458 (I183522,I183505,I177720);
DFFARX1 I_10459  ( .D(I183522), .CLK(I5694_clk), .RSTB(I183290_rst), .Q(I183539) );
nor I_10460 (I183556,I183539,I183392);
DFFARX1 I_10461  ( .D(I183539), .CLK(I5694_clk), .RSTB(I183290_rst), .Q(I183573) );
not I_10462 (I183261,I183573);
nand I_10463 (I183604,I183307,I177705);
and I_10464 (I183621,I183604,I183556);
DFFARX1 I_10465  ( .D(I183604), .CLK(I5694_clk), .RSTB(I183290_rst), .Q(I183258) );
DFFARX1 I_10466  ( .D(I177717), .CLK(I5694_clk), .RSTB(I183290_rst), .Q(I183652) );
nor I_10467 (I183669,I183652,I183375);
nand I_10468 (I183276,I183539,I183669);
nor I_10469 (I183700,I183652,I183440);
not I_10470 (I183273,I183652);
nand I_10471 (I183731,I183652,I183341);
and I_10472 (I183748,I183409,I183731);
DFFARX1 I_10473  ( .D(I183748), .CLK(I5694_clk), .RSTB(I183290_rst), .Q(I183252) );
DFFARX1 I_10474  ( .D(I183652), .CLK(I5694_clk), .RSTB(I183290_rst), .Q(I183255) );
DFFARX1 I_10475  ( .D(I177723), .CLK(I5694_clk), .RSTB(I183290_rst), .Q(I183793) );
not I_10476 (I183810,I183793);
nand I_10477 (I183827,I183810,I183375);
and I_10478 (I183844,I183604,I183827);
DFFARX1 I_10479  ( .D(I183844), .CLK(I5694_clk), .RSTB(I183290_rst), .Q(I183282) );
or I_10480 (I183875,I183810,I183621);
DFFARX1 I_10481  ( .D(I183875), .CLK(I5694_clk), .RSTB(I183290_rst), .Q(I183267) );
nand I_10482 (I183270,I183810,I183700);
not I_10483 (I183953_rst,I5701);
not I_10484 (I183970,I149185);
nor I_10485 (I183987,I149182,I149173);
nand I_10486 (I184004,I183987,I149176);
nor I_10487 (I184021,I183970,I149182);
nand I_10488 (I184038,I184021,I149170);
not I_10489 (I184055,I184038);
not I_10490 (I184072,I149182);
nor I_10491 (I183942,I184038,I184072);
not I_10492 (I184103,I184072);
nand I_10493 (I183927,I184038,I184103);
not I_10494 (I184134,I149191);
nor I_10495 (I184151,I184134,I149194);
and I_10496 (I184168,I184151,I149179);
or I_10497 (I184185,I184168,I149167);
DFFARX1 I_10498  ( .D(I184185), .CLK(I5694_clk), .RSTB(I183953_rst), .Q(I184202) );
nor I_10499 (I184219,I184202,I184055);
DFFARX1 I_10500  ( .D(I184202), .CLK(I5694_clk), .RSTB(I183953_rst), .Q(I184236) );
not I_10501 (I183924,I184236);
nand I_10502 (I184267,I183970,I149191);
and I_10503 (I184284,I184267,I184219);
DFFARX1 I_10504  ( .D(I184267), .CLK(I5694_clk), .RSTB(I183953_rst), .Q(I183921) );
DFFARX1 I_10505  ( .D(I149188), .CLK(I5694_clk), .RSTB(I183953_rst), .Q(I184315) );
nor I_10506 (I184332,I184315,I184038);
nand I_10507 (I183939,I184202,I184332);
nor I_10508 (I184363,I184315,I184103);
not I_10509 (I183936,I184315);
nand I_10510 (I184394,I184315,I184004);
and I_10511 (I184411,I184072,I184394);
DFFARX1 I_10512  ( .D(I184411), .CLK(I5694_clk), .RSTB(I183953_rst), .Q(I183915) );
DFFARX1 I_10513  ( .D(I184315), .CLK(I5694_clk), .RSTB(I183953_rst), .Q(I183918) );
DFFARX1 I_10514  ( .D(I149197), .CLK(I5694_clk), .RSTB(I183953_rst), .Q(I184456) );
not I_10515 (I184473,I184456);
nand I_10516 (I184490,I184473,I184038);
and I_10517 (I184507,I184267,I184490);
DFFARX1 I_10518  ( .D(I184507), .CLK(I5694_clk), .RSTB(I183953_rst), .Q(I183945) );
or I_10519 (I184538,I184473,I184284);
DFFARX1 I_10520  ( .D(I184538), .CLK(I5694_clk), .RSTB(I183953_rst), .Q(I183930) );
nand I_10521 (I183933,I184473,I184363);
not I_10522 (I184616_rst,I5701);
not I_10523 (I184633,I169199);
nor I_10524 (I184650,I169196,I169220);
nand I_10525 (I184667,I184650,I169217);
nor I_10526 (I184684,I184633,I169196);
nand I_10527 (I184701,I184684,I169223);
not I_10528 (I184718,I184701);
not I_10529 (I184735,I169196);
nor I_10530 (I184605,I184701,I184735);
not I_10531 (I184766,I184735);
nand I_10532 (I184590,I184701,I184766);
not I_10533 (I184797,I169214);
nor I_10534 (I184814,I184797,I169205);
and I_10535 (I184831,I184814,I169202);
or I_10536 (I184848,I184831,I169211);
DFFARX1 I_10537  ( .D(I184848), .CLK(I5694_clk), .RSTB(I184616_rst), .Q(I184865) );
nor I_10538 (I184882,I184865,I184718);
DFFARX1 I_10539  ( .D(I184865), .CLK(I5694_clk), .RSTB(I184616_rst), .Q(I184899) );
not I_10540 (I184587,I184899);
nand I_10541 (I184930,I184633,I169214);
and I_10542 (I184947,I184930,I184882);
DFFARX1 I_10543  ( .D(I184930), .CLK(I5694_clk), .RSTB(I184616_rst), .Q(I184584) );
DFFARX1 I_10544  ( .D(I169193), .CLK(I5694_clk), .RSTB(I184616_rst), .Q(I184978) );
nor I_10545 (I184995,I184978,I184701);
nand I_10546 (I184602,I184865,I184995);
nor I_10547 (I185026,I184978,I184766);
not I_10548 (I184599,I184978);
nand I_10549 (I185057,I184978,I184667);
and I_10550 (I185074,I184735,I185057);
DFFARX1 I_10551  ( .D(I185074), .CLK(I5694_clk), .RSTB(I184616_rst), .Q(I184578) );
DFFARX1 I_10552  ( .D(I184978), .CLK(I5694_clk), .RSTB(I184616_rst), .Q(I184581) );
DFFARX1 I_10553  ( .D(I169208), .CLK(I5694_clk), .RSTB(I184616_rst), .Q(I185119) );
not I_10554 (I185136,I185119);
nand I_10555 (I185153,I185136,I184701);
and I_10556 (I185170,I184930,I185153);
DFFARX1 I_10557  ( .D(I185170), .CLK(I5694_clk), .RSTB(I184616_rst), .Q(I184608) );
or I_10558 (I185201,I185136,I184947);
DFFARX1 I_10559  ( .D(I185201), .CLK(I5694_clk), .RSTB(I184616_rst), .Q(I184593) );
nand I_10560 (I184596,I185136,I185026);
not I_10561 (I185279_rst,I5701);
not I_10562 (I185296,I171783);
nor I_10563 (I185313,I171780,I171804);
nand I_10564 (I185330,I185313,I171801);
nor I_10565 (I185347,I185296,I171780);
nand I_10566 (I185364,I185347,I171807);
not I_10567 (I185381,I185364);
not I_10568 (I185398,I171780);
nor I_10569 (I185268,I185364,I185398);
not I_10570 (I185429,I185398);
nand I_10571 (I185253,I185364,I185429);
not I_10572 (I185460,I171798);
nor I_10573 (I185477,I185460,I171789);
and I_10574 (I185494,I185477,I171786);
or I_10575 (I185511,I185494,I171795);
DFFARX1 I_10576  ( .D(I185511), .CLK(I5694_clk), .RSTB(I185279_rst), .Q(I185528) );
nor I_10577 (I185545,I185528,I185381);
DFFARX1 I_10578  ( .D(I185528), .CLK(I5694_clk), .RSTB(I185279_rst), .Q(I185562) );
not I_10579 (I185250,I185562);
nand I_10580 (I185593,I185296,I171798);
and I_10581 (I185610,I185593,I185545);
DFFARX1 I_10582  ( .D(I185593), .CLK(I5694_clk), .RSTB(I185279_rst), .Q(I185247) );
DFFARX1 I_10583  ( .D(I171777), .CLK(I5694_clk), .RSTB(I185279_rst), .Q(I185641) );
nor I_10584 (I185658,I185641,I185364);
nand I_10585 (I185265,I185528,I185658);
nor I_10586 (I185689,I185641,I185429);
not I_10587 (I185262,I185641);
nand I_10588 (I185720,I185641,I185330);
and I_10589 (I185737,I185398,I185720);
DFFARX1 I_10590  ( .D(I185737), .CLK(I5694_clk), .RSTB(I185279_rst), .Q(I185241) );
DFFARX1 I_10591  ( .D(I185641), .CLK(I5694_clk), .RSTB(I185279_rst), .Q(I185244) );
DFFARX1 I_10592  ( .D(I171792), .CLK(I5694_clk), .RSTB(I185279_rst), .Q(I185782) );
not I_10593 (I185799,I185782);
nand I_10594 (I185816,I185799,I185364);
and I_10595 (I185833,I185593,I185816);
DFFARX1 I_10596  ( .D(I185833), .CLK(I5694_clk), .RSTB(I185279_rst), .Q(I185271) );
or I_10597 (I185864,I185799,I185610);
DFFARX1 I_10598  ( .D(I185864), .CLK(I5694_clk), .RSTB(I185279_rst), .Q(I185256) );
nand I_10599 (I185259,I185799,I185689);
not I_10600 (I185942_rst,I5701);
not I_10601 (I185959,I182684);
nor I_10602 (I185976,I182657,I182660);
nand I_10603 (I185993,I185976,I182672);
nor I_10604 (I186010,I185959,I182657);
nand I_10605 (I186027,I186010,I182678);
not I_10606 (I186044,I186027);
not I_10607 (I186061,I182657);
nor I_10608 (I185931,I186027,I186061);
not I_10609 (I186092,I186061);
nand I_10610 (I185916,I186027,I186092);
not I_10611 (I186123,I182681);
nor I_10612 (I186140,I186123,I182663);
and I_10613 (I186157,I186140,I182666);
or I_10614 (I186174,I186157,I182687);
DFFARX1 I_10615  ( .D(I186174), .CLK(I5694_clk), .RSTB(I185942_rst), .Q(I186191) );
nor I_10616 (I186208,I186191,I186044);
DFFARX1 I_10617  ( .D(I186191), .CLK(I5694_clk), .RSTB(I185942_rst), .Q(I186225) );
not I_10618 (I185913,I186225);
nand I_10619 (I186256,I185959,I182681);
and I_10620 (I186273,I186256,I186208);
DFFARX1 I_10621  ( .D(I186256), .CLK(I5694_clk), .RSTB(I185942_rst), .Q(I185910) );
DFFARX1 I_10622  ( .D(I182669), .CLK(I5694_clk), .RSTB(I185942_rst), .Q(I186304) );
nor I_10623 (I186321,I186304,I186027);
nand I_10624 (I185928,I186191,I186321);
nor I_10625 (I186352,I186304,I186092);
not I_10626 (I185925,I186304);
nand I_10627 (I186383,I186304,I185993);
and I_10628 (I186400,I186061,I186383);
DFFARX1 I_10629  ( .D(I186400), .CLK(I5694_clk), .RSTB(I185942_rst), .Q(I185904) );
DFFARX1 I_10630  ( .D(I186304), .CLK(I5694_clk), .RSTB(I185942_rst), .Q(I185907) );
DFFARX1 I_10631  ( .D(I182675), .CLK(I5694_clk), .RSTB(I185942_rst), .Q(I186445) );
not I_10632 (I186462,I186445);
nand I_10633 (I186479,I186462,I186027);
and I_10634 (I186496,I186256,I186479);
DFFARX1 I_10635  ( .D(I186496), .CLK(I5694_clk), .RSTB(I185942_rst), .Q(I185934) );
or I_10636 (I186527,I186462,I186273);
DFFARX1 I_10637  ( .D(I186527), .CLK(I5694_clk), .RSTB(I185942_rst), .Q(I185919) );
nand I_10638 (I185922,I186462,I186352);
not I_10639 (I186605_rst,I5701);
not I_10640 (I186622,I129595);
nor I_10641 (I186639,I129592,I129610);
nand I_10642 (I186656,I186639,I129613);
nor I_10643 (I186673,I186622,I129592);
nand I_10644 (I186690,I186673,I129598);
not I_10645 (I186707,I186690);
not I_10646 (I186724,I129592);
nor I_10647 (I186594,I186690,I186724);
not I_10648 (I186755,I186724);
nand I_10649 (I186579,I186690,I186755);
not I_10650 (I186786,I129607);
nor I_10651 (I186803,I186786,I129589);
and I_10652 (I186820,I186803,I129583);
or I_10653 (I186837,I186820,I129601);
DFFARX1 I_10654  ( .D(I186837), .CLK(I5694_clk), .RSTB(I186605_rst), .Q(I186854) );
nor I_10655 (I186871,I186854,I186707);
DFFARX1 I_10656  ( .D(I186854), .CLK(I5694_clk), .RSTB(I186605_rst), .Q(I186888) );
not I_10657 (I186576,I186888);
nand I_10658 (I186919,I186622,I129607);
and I_10659 (I186936,I186919,I186871);
DFFARX1 I_10660  ( .D(I186919), .CLK(I5694_clk), .RSTB(I186605_rst), .Q(I186573) );
DFFARX1 I_10661  ( .D(I129586), .CLK(I5694_clk), .RSTB(I186605_rst), .Q(I186967) );
nor I_10662 (I186984,I186967,I186690);
nand I_10663 (I186591,I186854,I186984);
nor I_10664 (I187015,I186967,I186755);
not I_10665 (I186588,I186967);
nand I_10666 (I187046,I186967,I186656);
and I_10667 (I187063,I186724,I187046);
DFFARX1 I_10668  ( .D(I187063), .CLK(I5694_clk), .RSTB(I186605_rst), .Q(I186567) );
DFFARX1 I_10669  ( .D(I186967), .CLK(I5694_clk), .RSTB(I186605_rst), .Q(I186570) );
DFFARX1 I_10670  ( .D(I129604), .CLK(I5694_clk), .RSTB(I186605_rst), .Q(I187108) );
not I_10671 (I187125,I187108);
nand I_10672 (I187142,I187125,I186690);
and I_10673 (I187159,I186919,I187142);
DFFARX1 I_10674  ( .D(I187159), .CLK(I5694_clk), .RSTB(I186605_rst), .Q(I186597) );
or I_10675 (I187190,I187125,I186936);
DFFARX1 I_10676  ( .D(I187190), .CLK(I5694_clk), .RSTB(I186605_rst), .Q(I186582) );
nand I_10677 (I186585,I187125,I187015);
not I_10678 (I187268_rst,I5701);
not I_10679 (I187285,I160161);
nor I_10680 (I187302,I160152,I160158);
nand I_10681 (I187319,I187302,I160170);
nor I_10682 (I187336,I187285,I160152);
nand I_10683 (I187353,I187336,I160155);
not I_10684 (I187370,I187353);
not I_10685 (I187387,I160152);
nor I_10686 (I187257,I187353,I187387);
not I_10687 (I187418,I187387);
nand I_10688 (I187242,I187353,I187418);
not I_10689 (I187449,I160179);
nor I_10690 (I187466,I187449,I160173);
and I_10691 (I187483,I187466,I160164);
or I_10692 (I187500,I187483,I160149);
DFFARX1 I_10693  ( .D(I187500), .CLK(I5694_clk), .RSTB(I187268_rst), .Q(I187517) );
nor I_10694 (I187534,I187517,I187370);
DFFARX1 I_10695  ( .D(I187517), .CLK(I5694_clk), .RSTB(I187268_rst), .Q(I187551) );
not I_10696 (I187239,I187551);
nand I_10697 (I187582,I187285,I160179);
and I_10698 (I187599,I187582,I187534);
DFFARX1 I_10699  ( .D(I187582), .CLK(I5694_clk), .RSTB(I187268_rst), .Q(I187236) );
DFFARX1 I_10700  ( .D(I160167), .CLK(I5694_clk), .RSTB(I187268_rst), .Q(I187630) );
nor I_10701 (I187647,I187630,I187353);
nand I_10702 (I187254,I187517,I187647);
nor I_10703 (I187678,I187630,I187418);
not I_10704 (I187251,I187630);
nand I_10705 (I187709,I187630,I187319);
and I_10706 (I187726,I187387,I187709);
DFFARX1 I_10707  ( .D(I187726), .CLK(I5694_clk), .RSTB(I187268_rst), .Q(I187230) );
DFFARX1 I_10708  ( .D(I187630), .CLK(I5694_clk), .RSTB(I187268_rst), .Q(I187233) );
DFFARX1 I_10709  ( .D(I160176), .CLK(I5694_clk), .RSTB(I187268_rst), .Q(I187771) );
not I_10710 (I187788,I187771);
nand I_10711 (I187805,I187788,I187353);
and I_10712 (I187822,I187582,I187805);
DFFARX1 I_10713  ( .D(I187822), .CLK(I5694_clk), .RSTB(I187268_rst), .Q(I187260) );
or I_10714 (I187853,I187788,I187599);
DFFARX1 I_10715  ( .D(I187853), .CLK(I5694_clk), .RSTB(I187268_rst), .Q(I187245) );
nand I_10716 (I187248,I187788,I187678);
not I_10717 (I187931_rst,I5701);
not I_10718 (I187948,I155225);
nor I_10719 (I187965,I155243,I155234);
nand I_10720 (I187982,I187965,I155240);
nor I_10721 (I187999,I187948,I155243);
nand I_10722 (I188016,I187999,I155246);
not I_10723 (I188033,I188016);
not I_10724 (I188050,I155243);
nor I_10725 (I187920,I188016,I188050);
not I_10726 (I188081,I188050);
nand I_10727 (I187905,I188016,I188081);
not I_10728 (I188112,I155222);
nor I_10729 (I188129,I188112,I155237);
and I_10730 (I188146,I188129,I155219);
or I_10731 (I188163,I188146,I155228);
DFFARX1 I_10732  ( .D(I188163), .CLK(I5694_clk), .RSTB(I187931_rst), .Q(I188180) );
nor I_10733 (I188197,I188180,I188033);
DFFARX1 I_10734  ( .D(I188180), .CLK(I5694_clk), .RSTB(I187931_rst), .Q(I188214) );
not I_10735 (I187902,I188214);
nand I_10736 (I188245,I187948,I155222);
and I_10737 (I188262,I188245,I188197);
DFFARX1 I_10738  ( .D(I188245), .CLK(I5694_clk), .RSTB(I187931_rst), .Q(I187899) );
DFFARX1 I_10739  ( .D(I155231), .CLK(I5694_clk), .RSTB(I187931_rst), .Q(I188293) );
nor I_10740 (I188310,I188293,I188016);
nand I_10741 (I187917,I188180,I188310);
nor I_10742 (I188341,I188293,I188081);
not I_10743 (I187914,I188293);
nand I_10744 (I188372,I188293,I187982);
and I_10745 (I188389,I188050,I188372);
DFFARX1 I_10746  ( .D(I188389), .CLK(I5694_clk), .RSTB(I187931_rst), .Q(I187893) );
DFFARX1 I_10747  ( .D(I188293), .CLK(I5694_clk), .RSTB(I187931_rst), .Q(I187896) );
DFFARX1 I_10748  ( .D(I155249), .CLK(I5694_clk), .RSTB(I187931_rst), .Q(I188434) );
not I_10749 (I188451,I188434);
nand I_10750 (I188468,I188451,I188016);
and I_10751 (I188485,I188245,I188468);
DFFARX1 I_10752  ( .D(I188485), .CLK(I5694_clk), .RSTB(I187931_rst), .Q(I187923) );
or I_10753 (I188516,I188451,I188262);
DFFARX1 I_10754  ( .D(I188516), .CLK(I5694_clk), .RSTB(I187931_rst), .Q(I187908) );
nand I_10755 (I187911,I188451,I188341);
not I_10756 (I188594_rst,I5701);
not I_10757 (I188611,I161884);
nor I_10758 (I188628,I161890,I161893);
nand I_10759 (I188645,I188628,I161869);
nor I_10760 (I188662,I188611,I161890);
nand I_10761 (I188679,I188662,I161878);
not I_10762 (I188696,I188679);
not I_10763 (I188713,I161890);
nor I_10764 (I188583,I188679,I188713);
not I_10765 (I188744,I188713);
nand I_10766 (I188568,I188679,I188744);
not I_10767 (I188775,I161872);
nor I_10768 (I188792,I188775,I161896);
and I_10769 (I188809,I188792,I161866);
or I_10770 (I188826,I188809,I161875);
DFFARX1 I_10771  ( .D(I188826), .CLK(I5694_clk), .RSTB(I188594_rst), .Q(I188843) );
nor I_10772 (I188860,I188843,I188696);
DFFARX1 I_10773  ( .D(I188843), .CLK(I5694_clk), .RSTB(I188594_rst), .Q(I188877) );
not I_10774 (I188565,I188877);
nand I_10775 (I188908,I188611,I161872);
and I_10776 (I188925,I188908,I188860);
DFFARX1 I_10777  ( .D(I188908), .CLK(I5694_clk), .RSTB(I188594_rst), .Q(I188562) );
DFFARX1 I_10778  ( .D(I161881), .CLK(I5694_clk), .RSTB(I188594_rst), .Q(I188956) );
nor I_10779 (I188973,I188956,I188679);
nand I_10780 (I188580,I188843,I188973);
nor I_10781 (I189004,I188956,I188744);
not I_10782 (I188577,I188956);
nand I_10783 (I189035,I188956,I188645);
and I_10784 (I189052,I188713,I189035);
DFFARX1 I_10785  ( .D(I189052), .CLK(I5694_clk), .RSTB(I188594_rst), .Q(I188556) );
DFFARX1 I_10786  ( .D(I188956), .CLK(I5694_clk), .RSTB(I188594_rst), .Q(I188559) );
DFFARX1 I_10787  ( .D(I161887), .CLK(I5694_clk), .RSTB(I188594_rst), .Q(I189097) );
not I_10788 (I189114,I189097);
nand I_10789 (I189131,I189114,I188679);
and I_10790 (I189148,I188908,I189131);
DFFARX1 I_10791  ( .D(I189148), .CLK(I5694_clk), .RSTB(I188594_rst), .Q(I188586) );
or I_10792 (I189179,I189114,I188925);
DFFARX1 I_10793  ( .D(I189179), .CLK(I5694_clk), .RSTB(I188594_rst), .Q(I188571) );
nand I_10794 (I188574,I189114,I189004);
not I_10795 (I189257_rst,I5701);
not I_10796 (I189274,I150375);
nor I_10797 (I189291,I150372,I150363);
nand I_10798 (I189308,I189291,I150366);
nor I_10799 (I189325,I189274,I150372);
nand I_10800 (I189342,I189325,I150360);
not I_10801 (I189359,I189342);
not I_10802 (I189376,I150372);
nor I_10803 (I189246,I189342,I189376);
not I_10804 (I189407,I189376);
nand I_10805 (I189231,I189342,I189407);
not I_10806 (I189438,I150381);
nor I_10807 (I189455,I189438,I150384);
and I_10808 (I189472,I189455,I150369);
or I_10809 (I189489,I189472,I150357);
DFFARX1 I_10810  ( .D(I189489), .CLK(I5694_clk), .RSTB(I189257_rst), .Q(I189506) );
nor I_10811 (I189523,I189506,I189359);
DFFARX1 I_10812  ( .D(I189506), .CLK(I5694_clk), .RSTB(I189257_rst), .Q(I189540) );
not I_10813 (I189228,I189540);
nand I_10814 (I189571,I189274,I150381);
and I_10815 (I189588,I189571,I189523);
DFFARX1 I_10816  ( .D(I189571), .CLK(I5694_clk), .RSTB(I189257_rst), .Q(I189225) );
DFFARX1 I_10817  ( .D(I150378), .CLK(I5694_clk), .RSTB(I189257_rst), .Q(I189619) );
nor I_10818 (I189636,I189619,I189342);
nand I_10819 (I189243,I189506,I189636);
nor I_10820 (I189667,I189619,I189407);
not I_10821 (I189240,I189619);
nand I_10822 (I189698,I189619,I189308);
and I_10823 (I189715,I189376,I189698);
DFFARX1 I_10824  ( .D(I189715), .CLK(I5694_clk), .RSTB(I189257_rst), .Q(I189219) );
DFFARX1 I_10825  ( .D(I189619), .CLK(I5694_clk), .RSTB(I189257_rst), .Q(I189222) );
DFFARX1 I_10826  ( .D(I150387), .CLK(I5694_clk), .RSTB(I189257_rst), .Q(I189760) );
not I_10827 (I189777,I189760);
nand I_10828 (I189794,I189777,I189342);
and I_10829 (I189811,I189571,I189794);
DFFARX1 I_10830  ( .D(I189811), .CLK(I5694_clk), .RSTB(I189257_rst), .Q(I189249) );
or I_10831 (I189842,I189777,I189588);
DFFARX1 I_10832  ( .D(I189842), .CLK(I5694_clk), .RSTB(I189257_rst), .Q(I189234) );
nand I_10833 (I189237,I189777,I189667);
not I_10834 (I189920_rst,I5701);
not I_10835 (I189937,I136695);
nor I_10836 (I189954,I136698,I136704);
nand I_10837 (I189971,I189954,I136710);
nor I_10838 (I189988,I189937,I136698);
nand I_10839 (I190005,I189988,I136689);
not I_10840 (I190022,I190005);
not I_10841 (I190039,I136698);
nor I_10842 (I189909,I190005,I190039);
not I_10843 (I190070,I190039);
nand I_10844 (I189894,I190005,I190070);
not I_10845 (I190101,I136701);
nor I_10846 (I190118,I190101,I136716);
and I_10847 (I190135,I190118,I136719);
or I_10848 (I190152,I190135,I136692);
DFFARX1 I_10849  ( .D(I190152), .CLK(I5694_clk), .RSTB(I189920_rst), .Q(I190169) );
nor I_10850 (I190186,I190169,I190022);
DFFARX1 I_10851  ( .D(I190169), .CLK(I5694_clk), .RSTB(I189920_rst), .Q(I190203) );
not I_10852 (I189891,I190203);
nand I_10853 (I190234,I189937,I136701);
and I_10854 (I190251,I190234,I190186);
DFFARX1 I_10855  ( .D(I190234), .CLK(I5694_clk), .RSTB(I189920_rst), .Q(I189888) );
DFFARX1 I_10856  ( .D(I136713), .CLK(I5694_clk), .RSTB(I189920_rst), .Q(I190282) );
nor I_10857 (I190299,I190282,I190005);
nand I_10858 (I189906,I190169,I190299);
nor I_10859 (I190330,I190282,I190070);
not I_10860 (I189903,I190282);
nand I_10861 (I190361,I190282,I189971);
and I_10862 (I190378,I190039,I190361);
DFFARX1 I_10863  ( .D(I190378), .CLK(I5694_clk), .RSTB(I189920_rst), .Q(I189882) );
DFFARX1 I_10864  ( .D(I190282), .CLK(I5694_clk), .RSTB(I189920_rst), .Q(I189885) );
DFFARX1 I_10865  ( .D(I136707), .CLK(I5694_clk), .RSTB(I189920_rst), .Q(I190423) );
not I_10866 (I190440,I190423);
nand I_10867 (I190457,I190440,I190005);
and I_10868 (I190474,I190234,I190457);
DFFARX1 I_10869  ( .D(I190474), .CLK(I5694_clk), .RSTB(I189920_rst), .Q(I189912) );
or I_10870 (I190505,I190440,I190251);
DFFARX1 I_10871  ( .D(I190505), .CLK(I5694_clk), .RSTB(I189920_rst), .Q(I189897) );
nand I_10872 (I189900,I190440,I190330);
not I_10873 (I190583_rst,I5701);
not I_10874 (I190600,I139084);
nor I_10875 (I190617,I139096,I139078);
nand I_10876 (I190634,I190617,I139099);
nor I_10877 (I190651,I190600,I139096);
nand I_10878 (I190668,I190651,I139090);
not I_10879 (I190685,I190668);
not I_10880 (I190702,I139096);
nor I_10881 (I190572,I190668,I190702);
not I_10882 (I190733,I190702);
nand I_10883 (I190557,I190668,I190733);
not I_10884 (I190764,I139081);
nor I_10885 (I190781,I190764,I139075);
and I_10886 (I190798,I190781,I139087);
or I_10887 (I190815,I190798,I139072);
DFFARX1 I_10888  ( .D(I190815), .CLK(I5694_clk), .RSTB(I190583_rst), .Q(I190832) );
nor I_10889 (I190849,I190832,I190685);
DFFARX1 I_10890  ( .D(I190832), .CLK(I5694_clk), .RSTB(I190583_rst), .Q(I190866) );
not I_10891 (I190554,I190866);
nand I_10892 (I190897,I190600,I139081);
and I_10893 (I190914,I190897,I190849);
DFFARX1 I_10894  ( .D(I190897), .CLK(I5694_clk), .RSTB(I190583_rst), .Q(I190551) );
DFFARX1 I_10895  ( .D(I139069), .CLK(I5694_clk), .RSTB(I190583_rst), .Q(I190945) );
nor I_10896 (I190962,I190945,I190668);
nand I_10897 (I190569,I190832,I190962);
nor I_10898 (I190993,I190945,I190733);
not I_10899 (I190566,I190945);
nand I_10900 (I191024,I190945,I190634);
and I_10901 (I191041,I190702,I191024);
DFFARX1 I_10902  ( .D(I191041), .CLK(I5694_clk), .RSTB(I190583_rst), .Q(I190545) );
DFFARX1 I_10903  ( .D(I190945), .CLK(I5694_clk), .RSTB(I190583_rst), .Q(I190548) );
DFFARX1 I_10904  ( .D(I139093), .CLK(I5694_clk), .RSTB(I190583_rst), .Q(I191086) );
not I_10905 (I191103,I191086);
nand I_10906 (I191120,I191103,I190668);
and I_10907 (I191137,I190897,I191120);
DFFARX1 I_10908  ( .D(I191137), .CLK(I5694_clk), .RSTB(I190583_rst), .Q(I190575) );
or I_10909 (I191168,I191103,I190914);
DFFARX1 I_10910  ( .D(I191168), .CLK(I5694_clk), .RSTB(I190583_rst), .Q(I190560) );
nand I_10911 (I190563,I191103,I190993);
not I_10912 (I191246_rst,I5701);
not I_10913 (I191263,I163567);
nor I_10914 (I191280,I163573,I163576);
nand I_10915 (I191297,I191280,I163552);
nor I_10916 (I191314,I191263,I163573);
nand I_10917 (I191331,I191314,I163561);
not I_10918 (I191348,I191331);
not I_10919 (I191365,I163573);
nor I_10920 (I191235,I191331,I191365);
not I_10921 (I191396,I191365);
nand I_10922 (I191220,I191331,I191396);
not I_10923 (I191427,I163555);
nor I_10924 (I191444,I191427,I163579);
and I_10925 (I191461,I191444,I163549);
or I_10926 (I191478,I191461,I163558);
DFFARX1 I_10927  ( .D(I191478), .CLK(I5694_clk), .RSTB(I191246_rst), .Q(I191495) );
nor I_10928 (I191512,I191495,I191348);
DFFARX1 I_10929  ( .D(I191495), .CLK(I5694_clk), .RSTB(I191246_rst), .Q(I191529) );
not I_10930 (I191217,I191529);
nand I_10931 (I191560,I191263,I163555);
and I_10932 (I191577,I191560,I191512);
DFFARX1 I_10933  ( .D(I191560), .CLK(I5694_clk), .RSTB(I191246_rst), .Q(I191214) );
DFFARX1 I_10934  ( .D(I163564), .CLK(I5694_clk), .RSTB(I191246_rst), .Q(I191608) );
nor I_10935 (I191625,I191608,I191331);
nand I_10936 (I191232,I191495,I191625);
nor I_10937 (I191656,I191608,I191396);
not I_10938 (I191229,I191608);
nand I_10939 (I191687,I191608,I191297);
and I_10940 (I191704,I191365,I191687);
DFFARX1 I_10941  ( .D(I191704), .CLK(I5694_clk), .RSTB(I191246_rst), .Q(I191208) );
DFFARX1 I_10942  ( .D(I191608), .CLK(I5694_clk), .RSTB(I191246_rst), .Q(I191211) );
DFFARX1 I_10943  ( .D(I163570), .CLK(I5694_clk), .RSTB(I191246_rst), .Q(I191749) );
not I_10944 (I191766,I191749);
nand I_10945 (I191783,I191766,I191331);
and I_10946 (I191800,I191560,I191783);
DFFARX1 I_10947  ( .D(I191800), .CLK(I5694_clk), .RSTB(I191246_rst), .Q(I191238) );
or I_10948 (I191831,I191766,I191577);
DFFARX1 I_10949  ( .D(I191831), .CLK(I5694_clk), .RSTB(I191246_rst), .Q(I191223) );
nand I_10950 (I191226,I191766,I191656);
not I_10951 (I191909_rst,I5701);
not I_10952 (I191926,I165323);
nor I_10953 (I191943,I165320,I165344);
nand I_10954 (I191960,I191943,I165341);
nor I_10955 (I191977,I191926,I165320);
nand I_10956 (I191994,I191977,I165347);
not I_10957 (I192011,I191994);
not I_10958 (I192028,I165320);
nor I_10959 (I191898,I191994,I192028);
not I_10960 (I192059,I192028);
nand I_10961 (I191883,I191994,I192059);
not I_10962 (I192090,I165338);
nor I_10963 (I192107,I192090,I165329);
and I_10964 (I192124,I192107,I165326);
or I_10965 (I192141,I192124,I165335);
DFFARX1 I_10966  ( .D(I192141), .CLK(I5694_clk), .RSTB(I191909_rst), .Q(I192158) );
nor I_10967 (I192175,I192158,I192011);
DFFARX1 I_10968  ( .D(I192158), .CLK(I5694_clk), .RSTB(I191909_rst), .Q(I192192) );
not I_10969 (I191880,I192192);
nand I_10970 (I192223,I191926,I165338);
and I_10971 (I192240,I192223,I192175);
DFFARX1 I_10972  ( .D(I192223), .CLK(I5694_clk), .RSTB(I191909_rst), .Q(I191877) );
DFFARX1 I_10973  ( .D(I165317), .CLK(I5694_clk), .RSTB(I191909_rst), .Q(I192271) );
nor I_10974 (I192288,I192271,I191994);
nand I_10975 (I191895,I192158,I192288);
nor I_10976 (I192319,I192271,I192059);
not I_10977 (I191892,I192271);
nand I_10978 (I192350,I192271,I191960);
and I_10979 (I192367,I192028,I192350);
DFFARX1 I_10980  ( .D(I192367), .CLK(I5694_clk), .RSTB(I191909_rst), .Q(I191871) );
DFFARX1 I_10981  ( .D(I192271), .CLK(I5694_clk), .RSTB(I191909_rst), .Q(I191874) );
DFFARX1 I_10982  ( .D(I165332), .CLK(I5694_clk), .RSTB(I191909_rst), .Q(I192412) );
not I_10983 (I192429,I192412);
nand I_10984 (I192446,I192429,I191994);
and I_10985 (I192463,I192223,I192446);
DFFARX1 I_10986  ( .D(I192463), .CLK(I5694_clk), .RSTB(I191909_rst), .Q(I191901) );
or I_10987 (I192494,I192429,I192240);
DFFARX1 I_10988  ( .D(I192494), .CLK(I5694_clk), .RSTB(I191909_rst), .Q(I191886) );
nand I_10989 (I191889,I192429,I192319);
not I_10990 (I192572_rst,I5701);
not I_10991 (I192589,I128303);
nor I_10992 (I192606,I128300,I128318);
nand I_10993 (I192623,I192606,I128321);
nor I_10994 (I192640,I192589,I128300);
nand I_10995 (I192657,I192640,I128306);
not I_10996 (I192674,I192657);
not I_10997 (I192691,I128300);
nor I_10998 (I192561,I192657,I192691);
not I_10999 (I192722,I192691);
nand I_11000 (I192546,I192657,I192722);
not I_11001 (I192753,I128315);
nor I_11002 (I192770,I192753,I128297);
and I_11003 (I192787,I192770,I128291);
or I_11004 (I192804,I192787,I128309);
DFFARX1 I_11005  ( .D(I192804), .CLK(I5694_clk), .RSTB(I192572_rst), .Q(I192821) );
nor I_11006 (I192838,I192821,I192674);
DFFARX1 I_11007  ( .D(I192821), .CLK(I5694_clk), .RSTB(I192572_rst), .Q(I192855) );
not I_11008 (I192543,I192855);
nand I_11009 (I192886,I192589,I128315);
and I_11010 (I192903,I192886,I192838);
DFFARX1 I_11011  ( .D(I192886), .CLK(I5694_clk), .RSTB(I192572_rst), .Q(I192540) );
DFFARX1 I_11012  ( .D(I128294), .CLK(I5694_clk), .RSTB(I192572_rst), .Q(I192934) );
nor I_11013 (I192951,I192934,I192657);
nand I_11014 (I192558,I192821,I192951);
nor I_11015 (I192982,I192934,I192722);
not I_11016 (I192555,I192934);
nand I_11017 (I193013,I192934,I192623);
and I_11018 (I193030,I192691,I193013);
DFFARX1 I_11019  ( .D(I193030), .CLK(I5694_clk), .RSTB(I192572_rst), .Q(I192534) );
DFFARX1 I_11020  ( .D(I192934), .CLK(I5694_clk), .RSTB(I192572_rst), .Q(I192537) );
DFFARX1 I_11021  ( .D(I128312), .CLK(I5694_clk), .RSTB(I192572_rst), .Q(I193075) );
not I_11022 (I193092,I193075);
nand I_11023 (I193109,I193092,I192657);
and I_11024 (I193126,I192886,I193109);
DFFARX1 I_11025  ( .D(I193126), .CLK(I5694_clk), .RSTB(I192572_rst), .Q(I192564) );
or I_11026 (I193157,I193092,I192903);
DFFARX1 I_11027  ( .D(I193157), .CLK(I5694_clk), .RSTB(I192572_rst), .Q(I192549) );
nand I_11028 (I192552,I193092,I192982);
not I_11029 (I193235_rst,I5701);
not I_11030 (I193252,I140255);
nor I_11031 (I193269,I140243,I140234);
nand I_11032 (I193286,I193269,I140246);
nor I_11033 (I193303,I193252,I140243);
nand I_11034 (I193320,I193303,I140252);
DFFARX1 I_11035  ( .D(I193320), .CLK(I5694_clk), .RSTB(I193235_rst), .Q(I193337) );
not I_11036 (I193206,I193337);
not I_11037 (I193368,I140243);
not I_11038 (I193385,I193368);
not I_11039 (I193402,I140228);
nor I_11040 (I193419,I193402,I140249);
and I_11041 (I193436,I193419,I140240);
or I_11042 (I193453,I193436,I140237);
DFFARX1 I_11043  ( .D(I193453), .CLK(I5694_clk), .RSTB(I193235_rst), .Q(I193470) );
DFFARX1 I_11044  ( .D(I193470), .CLK(I5694_clk), .RSTB(I193235_rst), .Q(I193203) );
DFFARX1 I_11045  ( .D(I193470), .CLK(I5694_clk), .RSTB(I193235_rst), .Q(I193501) );
DFFARX1 I_11046  ( .D(I193470), .CLK(I5694_clk), .RSTB(I193235_rst), .Q(I193197) );
nand I_11047 (I193532,I193252,I140228);
nand I_11048 (I193549,I193532,I193286);
and I_11049 (I193566,I193368,I193549);
DFFARX1 I_11050  ( .D(I193566), .CLK(I5694_clk), .RSTB(I193235_rst), .Q(I193227) );
and I_11051 (I193200,I193532,I193501);
DFFARX1 I_11052  ( .D(I140225), .CLK(I5694_clk), .RSTB(I193235_rst), .Q(I193611) );
nor I_11053 (I193224,I193611,I193532);
nor I_11054 (I193642,I193611,I193286);
nand I_11055 (I193221,I193320,I193642);
not I_11056 (I193218,I193611);
DFFARX1 I_11057  ( .D(I140231), .CLK(I5694_clk), .RSTB(I193235_rst), .Q(I193687) );
not I_11058 (I193704,I193687);
nor I_11059 (I193721,I193704,I193385);
and I_11060 (I193738,I193611,I193721);
or I_11061 (I193755,I193532,I193738);
DFFARX1 I_11062  ( .D(I193755), .CLK(I5694_clk), .RSTB(I193235_rst), .Q(I193212) );
not I_11063 (I193786,I193704);
nor I_11064 (I193803,I193611,I193786);
nand I_11065 (I193215,I193704,I193803);
nand I_11066 (I193209,I193368,I193786);
not I_11067 (I193881_rst,I5701);
not I_11068 (I193898,I171152);
nor I_11069 (I193915,I171143,I171134);
nand I_11070 (I193932,I193915,I171149);
nor I_11071 (I193949,I193898,I171143);
nand I_11072 (I193966,I193949,I171146);
DFFARX1 I_11073  ( .D(I193966), .CLK(I5694_clk), .RSTB(I193881_rst), .Q(I193983) );
not I_11074 (I193852,I193983);
not I_11075 (I194014,I171143);
not I_11076 (I194031,I194014);
not I_11077 (I194048,I171155);
nor I_11078 (I194065,I194048,I171140);
and I_11079 (I194082,I194065,I171158);
or I_11080 (I194099,I194082,I171131);
DFFARX1 I_11081  ( .D(I194099), .CLK(I5694_clk), .RSTB(I193881_rst), .Q(I194116) );
DFFARX1 I_11082  ( .D(I194116), .CLK(I5694_clk), .RSTB(I193881_rst), .Q(I193849) );
DFFARX1 I_11083  ( .D(I194116), .CLK(I5694_clk), .RSTB(I193881_rst), .Q(I194147) );
DFFARX1 I_11084  ( .D(I194116), .CLK(I5694_clk), .RSTB(I193881_rst), .Q(I193843) );
nand I_11085 (I194178,I193898,I171155);
nand I_11086 (I194195,I194178,I193932);
and I_11087 (I194212,I194014,I194195);
DFFARX1 I_11088  ( .D(I194212), .CLK(I5694_clk), .RSTB(I193881_rst), .Q(I193873) );
and I_11089 (I193846,I194178,I194147);
DFFARX1 I_11090  ( .D(I171161), .CLK(I5694_clk), .RSTB(I193881_rst), .Q(I194257) );
nor I_11091 (I193870,I194257,I194178);
nor I_11092 (I194288,I194257,I193932);
nand I_11093 (I193867,I193966,I194288);
not I_11094 (I193864,I194257);
DFFARX1 I_11095  ( .D(I171137), .CLK(I5694_clk), .RSTB(I193881_rst), .Q(I194333) );
not I_11096 (I194350,I194333);
nor I_11097 (I194367,I194350,I194031);
and I_11098 (I194384,I194257,I194367);
or I_11099 (I194401,I194178,I194384);
DFFARX1 I_11100  ( .D(I194401), .CLK(I5694_clk), .RSTB(I193881_rst), .Q(I193858) );
not I_11101 (I194432,I194350);
nor I_11102 (I194449,I194257,I194432);
nand I_11103 (I193861,I194350,I194449);
nand I_11104 (I193855,I194014,I194432);
not I_11105 (I194527_rst,I5701);
not I_11106 (I194544,I175707);
nor I_11107 (I194561,I175728,I175710);
nand I_11108 (I194578,I194561,I175734);
nor I_11109 (I194595,I194544,I175728);
nand I_11110 (I194612,I194595,I175731);
DFFARX1 I_11111  ( .D(I194612), .CLK(I5694_clk), .RSTB(I194527_rst), .Q(I194629) );
not I_11112 (I194498,I194629);
not I_11113 (I194660,I175728);
not I_11114 (I194677,I194660);
not I_11115 (I194694,I175725);
nor I_11116 (I194711,I194694,I175704);
and I_11117 (I194728,I194711,I175716);
or I_11118 (I194745,I194728,I175713);
DFFARX1 I_11119  ( .D(I194745), .CLK(I5694_clk), .RSTB(I194527_rst), .Q(I194762) );
DFFARX1 I_11120  ( .D(I194762), .CLK(I5694_clk), .RSTB(I194527_rst), .Q(I194495) );
DFFARX1 I_11121  ( .D(I194762), .CLK(I5694_clk), .RSTB(I194527_rst), .Q(I194793) );
DFFARX1 I_11122  ( .D(I194762), .CLK(I5694_clk), .RSTB(I194527_rst), .Q(I194489) );
nand I_11123 (I194824,I194544,I175725);
nand I_11124 (I194841,I194824,I194578);
and I_11125 (I194858,I194660,I194841);
DFFARX1 I_11126  ( .D(I194858), .CLK(I5694_clk), .RSTB(I194527_rst), .Q(I194519) );
and I_11127 (I194492,I194824,I194793);
DFFARX1 I_11128  ( .D(I175719), .CLK(I5694_clk), .RSTB(I194527_rst), .Q(I194903) );
nor I_11129 (I194516,I194903,I194824);
nor I_11130 (I194934,I194903,I194578);
nand I_11131 (I194513,I194612,I194934);
not I_11132 (I194510,I194903);
DFFARX1 I_11133  ( .D(I175722), .CLK(I5694_clk), .RSTB(I194527_rst), .Q(I194979) );
not I_11134 (I194996,I194979);
nor I_11135 (I195013,I194996,I194677);
and I_11136 (I195030,I194903,I195013);
or I_11137 (I195047,I194824,I195030);
DFFARX1 I_11138  ( .D(I195047), .CLK(I5694_clk), .RSTB(I194527_rst), .Q(I194504) );
not I_11139 (I195078,I194996);
nor I_11140 (I195095,I194903,I195078);
nand I_11141 (I194507,I194996,I195095);
nand I_11142 (I194501,I194660,I195078);
not I_11143 (I195173_rst,I5701);
not I_11144 (I195190,I175044);
nor I_11145 (I195207,I175065,I175047);
nand I_11146 (I195224,I195207,I175071);
nor I_11147 (I195241,I195190,I175065);
nand I_11148 (I195258,I195241,I175068);
DFFARX1 I_11149  ( .D(I195258), .CLK(I5694_clk), .RSTB(I195173_rst), .Q(I195275) );
not I_11150 (I195144,I195275);
not I_11151 (I195306,I175065);
not I_11152 (I195323,I195306);
not I_11153 (I195340,I175062);
nor I_11154 (I195357,I195340,I175041);
and I_11155 (I195374,I195357,I175053);
or I_11156 (I195391,I195374,I175050);
DFFARX1 I_11157  ( .D(I195391), .CLK(I5694_clk), .RSTB(I195173_rst), .Q(I195408) );
DFFARX1 I_11158  ( .D(I195408), .CLK(I5694_clk), .RSTB(I195173_rst), .Q(I195141) );
DFFARX1 I_11159  ( .D(I195408), .CLK(I5694_clk), .RSTB(I195173_rst), .Q(I195439) );
DFFARX1 I_11160  ( .D(I195408), .CLK(I5694_clk), .RSTB(I195173_rst), .Q(I195135) );
nand I_11161 (I195470,I195190,I175062);
nand I_11162 (I195487,I195470,I195224);
and I_11163 (I195504,I195306,I195487);
DFFARX1 I_11164  ( .D(I195504), .CLK(I5694_clk), .RSTB(I195173_rst), .Q(I195165) );
and I_11165 (I195138,I195470,I195439);
DFFARX1 I_11166  ( .D(I175056), .CLK(I5694_clk), .RSTB(I195173_rst), .Q(I195549) );
nor I_11167 (I195162,I195549,I195470);
nor I_11168 (I195580,I195549,I195224);
nand I_11169 (I195159,I195258,I195580);
not I_11170 (I195156,I195549);
DFFARX1 I_11171  ( .D(I175059), .CLK(I5694_clk), .RSTB(I195173_rst), .Q(I195625) );
not I_11172 (I195642,I195625);
nor I_11173 (I195659,I195642,I195323);
and I_11174 (I195676,I195549,I195659);
or I_11175 (I195693,I195470,I195676);
DFFARX1 I_11176  ( .D(I195693), .CLK(I5694_clk), .RSTB(I195173_rst), .Q(I195150) );
not I_11177 (I195724,I195642);
nor I_11178 (I195741,I195549,I195724);
nand I_11179 (I195153,I195642,I195741);
nand I_11180 (I195147,I195306,I195724);
not I_11181 (I195819_rst,I5701);
not I_11182 (I195836,I160745);
nor I_11183 (I195853,I160730,I160736);
nand I_11184 (I195870,I195853,I160733);
nor I_11185 (I195887,I195836,I160730);
nand I_11186 (I195904,I195887,I160742);
DFFARX1 I_11187  ( .D(I195904), .CLK(I5694_clk), .RSTB(I195819_rst), .Q(I195921) );
not I_11188 (I195790,I195921);
not I_11189 (I195952,I160730);
not I_11190 (I195969,I195952);
not I_11191 (I195986,I160757);
nor I_11192 (I196003,I195986,I160751);
and I_11193 (I196020,I196003,I160748);
or I_11194 (I196037,I196020,I160727);
DFFARX1 I_11195  ( .D(I196037), .CLK(I5694_clk), .RSTB(I195819_rst), .Q(I196054) );
DFFARX1 I_11196  ( .D(I196054), .CLK(I5694_clk), .RSTB(I195819_rst), .Q(I195787) );
DFFARX1 I_11197  ( .D(I196054), .CLK(I5694_clk), .RSTB(I195819_rst), .Q(I196085) );
DFFARX1 I_11198  ( .D(I196054), .CLK(I5694_clk), .RSTB(I195819_rst), .Q(I195781) );
nand I_11199 (I196116,I195836,I160757);
nand I_11200 (I196133,I196116,I195870);
and I_11201 (I196150,I195952,I196133);
DFFARX1 I_11202  ( .D(I196150), .CLK(I5694_clk), .RSTB(I195819_rst), .Q(I195811) );
and I_11203 (I195784,I196116,I196085);
DFFARX1 I_11204  ( .D(I160754), .CLK(I5694_clk), .RSTB(I195819_rst), .Q(I196195) );
nor I_11205 (I195808,I196195,I196116);
nor I_11206 (I196226,I196195,I195870);
nand I_11207 (I195805,I195904,I196226);
not I_11208 (I195802,I196195);
DFFARX1 I_11209  ( .D(I160739), .CLK(I5694_clk), .RSTB(I195819_rst), .Q(I196271) );
not I_11210 (I196288,I196271);
nor I_11211 (I196305,I196288,I195969);
and I_11212 (I196322,I196195,I196305);
or I_11213 (I196339,I196116,I196322);
DFFARX1 I_11214  ( .D(I196339), .CLK(I5694_clk), .RSTB(I195819_rst), .Q(I195796) );
not I_11215 (I196370,I196288);
nor I_11216 (I196387,I196195,I196370);
nand I_11217 (I195799,I196288,I196387);
nand I_11218 (I195793,I195952,I196370);
not I_11219 (I196465_rst,I5701);
not I_11220 (I196482,I161314);
nor I_11221 (I196499,I161329,I161323);
nand I_11222 (I196516,I196499,I161332);
nor I_11223 (I196533,I196482,I161329);
nand I_11224 (I196550,I196533,I161308);
DFFARX1 I_11225  ( .D(I196550), .CLK(I5694_clk), .RSTB(I196465_rst), .Q(I196567) );
not I_11226 (I196436,I196567);
not I_11227 (I196598,I161329);
not I_11228 (I196615,I196598);
not I_11229 (I196632,I161305);
nor I_11230 (I196649,I196632,I161320);
and I_11231 (I196666,I196649,I161326);
or I_11232 (I196683,I196666,I161335);
DFFARX1 I_11233  ( .D(I196683), .CLK(I5694_clk), .RSTB(I196465_rst), .Q(I196700) );
DFFARX1 I_11234  ( .D(I196700), .CLK(I5694_clk), .RSTB(I196465_rst), .Q(I196433) );
DFFARX1 I_11235  ( .D(I196700), .CLK(I5694_clk), .RSTB(I196465_rst), .Q(I196731) );
DFFARX1 I_11236  ( .D(I196700), .CLK(I5694_clk), .RSTB(I196465_rst), .Q(I196427) );
nand I_11237 (I196762,I196482,I161305);
nand I_11238 (I196779,I196762,I196516);
and I_11239 (I196796,I196598,I196779);
DFFARX1 I_11240  ( .D(I196796), .CLK(I5694_clk), .RSTB(I196465_rst), .Q(I196457) );
and I_11241 (I196430,I196762,I196731);
DFFARX1 I_11242  ( .D(I161317), .CLK(I5694_clk), .RSTB(I196465_rst), .Q(I196841) );
nor I_11243 (I196454,I196841,I196762);
nor I_11244 (I196872,I196841,I196516);
nand I_11245 (I196451,I196550,I196872);
not I_11246 (I196448,I196841);
DFFARX1 I_11247  ( .D(I161311), .CLK(I5694_clk), .RSTB(I196465_rst), .Q(I196917) );
not I_11248 (I196934,I196917);
nor I_11249 (I196951,I196934,I196615);
and I_11250 (I196968,I196841,I196951);
or I_11251 (I196985,I196762,I196968);
DFFARX1 I_11252  ( .D(I196985), .CLK(I5694_clk), .RSTB(I196465_rst), .Q(I196442) );
not I_11253 (I197016,I196934);
nor I_11254 (I197033,I196841,I197016);
nand I_11255 (I196445,I196934,I197033);
nand I_11256 (I196439,I196598,I197016);
not I_11257 (I197111_rst,I5701);
not I_11258 (I197128,I156498);
nor I_11259 (I197145,I156495,I156480);
nand I_11260 (I197162,I197145,I156489);
nor I_11261 (I197179,I197128,I156495);
nand I_11262 (I197196,I197179,I156504);
DFFARX1 I_11263  ( .D(I197196), .CLK(I5694_clk), .RSTB(I197111_rst), .Q(I197213) );
not I_11264 (I197082,I197213);
not I_11265 (I197244,I156495);
not I_11266 (I197261,I197244);
not I_11267 (I197278,I156477);
nor I_11268 (I197295,I197278,I156483);
and I_11269 (I197312,I197295,I156507);
or I_11270 (I197329,I197312,I156501);
DFFARX1 I_11271  ( .D(I197329), .CLK(I5694_clk), .RSTB(I197111_rst), .Q(I197346) );
DFFARX1 I_11272  ( .D(I197346), .CLK(I5694_clk), .RSTB(I197111_rst), .Q(I197079) );
DFFARX1 I_11273  ( .D(I197346), .CLK(I5694_clk), .RSTB(I197111_rst), .Q(I197377) );
DFFARX1 I_11274  ( .D(I197346), .CLK(I5694_clk), .RSTB(I197111_rst), .Q(I197073) );
nand I_11275 (I197408,I197128,I156477);
nand I_11276 (I197425,I197408,I197162);
and I_11277 (I197442,I197244,I197425);
DFFARX1 I_11278  ( .D(I197442), .CLK(I5694_clk), .RSTB(I197111_rst), .Q(I197103) );
and I_11279 (I197076,I197408,I197377);
DFFARX1 I_11280  ( .D(I156486), .CLK(I5694_clk), .RSTB(I197111_rst), .Q(I197487) );
nor I_11281 (I197100,I197487,I197408);
nor I_11282 (I197518,I197487,I197162);
nand I_11283 (I197097,I197196,I197518);
not I_11284 (I197094,I197487);
DFFARX1 I_11285  ( .D(I156492), .CLK(I5694_clk), .RSTB(I197111_rst), .Q(I197563) );
not I_11286 (I197580,I197563);
nor I_11287 (I197597,I197580,I197261);
and I_11288 (I197614,I197487,I197597);
or I_11289 (I197631,I197408,I197614);
DFFARX1 I_11290  ( .D(I197631), .CLK(I5694_clk), .RSTB(I197111_rst), .Q(I197088) );
not I_11291 (I197662,I197580);
nor I_11292 (I197679,I197487,I197662);
nand I_11293 (I197091,I197580,I197679);
nand I_11294 (I197085,I197244,I197662);
not I_11295 (I197757_rst,I5701);
or I_11296 (I197774,I177036,I177057);
or I_11297 (I197791,I177054,I177036);
nor I_11298 (I197808,I177045,I177042);
DFFARX1 I_11299  ( .D(I197808), .CLK(I5694_clk), .RSTB(I197757_rst), .Q(I197825) );
DFFARX1 I_11300  ( .D(I197808), .CLK(I5694_clk), .RSTB(I197757_rst), .Q(I197719) );
not I_11301 (I197856,I177045);
and I_11302 (I197873,I197856,I177051);
nor I_11303 (I197890,I197873,I177057);
nor I_11304 (I197907,I177039,I177030);
DFFARX1 I_11305  ( .D(I197907), .CLK(I5694_clk), .RSTB(I197757_rst), .Q(I197924) );
not I_11306 (I197941,I197924);
DFFARX1 I_11307  ( .D(I197924), .CLK(I5694_clk), .RSTB(I197757_rst), .Q(I197728) );
nor I_11308 (I197972,I177039,I177054);
and I_11309 (I197722,I197972,I197825);
DFFARX1 I_11310  ( .D(I177033), .CLK(I5694_clk), .RSTB(I197757_rst), .Q(I198003) );
and I_11311 (I198020,I198003,I177048);
nand I_11312 (I198037,I198020,I197791);
and I_11313 (I198054,I197924,I198037);
DFFARX1 I_11314  ( .D(I198054), .CLK(I5694_clk), .RSTB(I197757_rst), .Q(I197749) );
nor I_11315 (I197746,I198020,I197890);
not I_11316 (I198099,I198020);
nor I_11317 (I198116,I197774,I198099);
nor I_11318 (I198133,I198020,I197972);
nand I_11319 (I197743,I197791,I198133);
nor I_11320 (I198164,I198020,I197941);
not I_11321 (I197740,I198020);
nand I_11322 (I197731,I198020,I197941);
DFFARX1 I_11323  ( .D(I177060), .CLK(I5694_clk), .RSTB(I197757_rst), .Q(I198209) );
and I_11324 (I198226,I198209,I198116);
or I_11325 (I198243,I197774,I198226);
DFFARX1 I_11326  ( .D(I198243), .CLK(I5694_clk), .RSTB(I197757_rst), .Q(I197734) );
nand I_11327 (I197737,I198209,I198164);
nand I_11328 (I198288,I198209,I197890);
and I_11329 (I198305,I197808,I198288);
DFFARX1 I_11330  ( .D(I198305), .CLK(I5694_clk), .RSTB(I197757_rst), .Q(I197725) );
not I_11331 (I198369_rst,I5701);
or I_11332 (I198386,I137913,I137928);
or I_11333 (I198403,I137943,I137913);
nor I_11334 (I198420,I137925,I137916);
DFFARX1 I_11335  ( .D(I198420), .CLK(I5694_clk), .RSTB(I198369_rst), .Q(I198437) );
DFFARX1 I_11336  ( .D(I198420), .CLK(I5694_clk), .RSTB(I198369_rst), .Q(I198331) );
not I_11337 (I198468,I137925);
and I_11338 (I198485,I198468,I137934);
nor I_11339 (I198502,I198485,I137928);
nor I_11340 (I198519,I137940,I137931);
DFFARX1 I_11341  ( .D(I198519), .CLK(I5694_clk), .RSTB(I198369_rst), .Q(I198536) );
not I_11342 (I198553,I198536);
DFFARX1 I_11343  ( .D(I198536), .CLK(I5694_clk), .RSTB(I198369_rst), .Q(I198340) );
nor I_11344 (I198584,I137940,I137943);
and I_11345 (I198334,I198584,I198437);
DFFARX1 I_11346  ( .D(I137919), .CLK(I5694_clk), .RSTB(I198369_rst), .Q(I198615) );
and I_11347 (I198632,I198615,I137922);
nand I_11348 (I198649,I198632,I198403);
and I_11349 (I198666,I198536,I198649);
DFFARX1 I_11350  ( .D(I198666), .CLK(I5694_clk), .RSTB(I198369_rst), .Q(I198361) );
nor I_11351 (I198358,I198632,I198502);
not I_11352 (I198711,I198632);
nor I_11353 (I198728,I198386,I198711);
nor I_11354 (I198745,I198632,I198584);
nand I_11355 (I198355,I198403,I198745);
nor I_11356 (I198776,I198632,I198553);
not I_11357 (I198352,I198632);
nand I_11358 (I198343,I198632,I198553);
DFFARX1 I_11359  ( .D(I137937), .CLK(I5694_clk), .RSTB(I198369_rst), .Q(I198821) );
and I_11360 (I198838,I198821,I198728);
or I_11361 (I198855,I198386,I198838);
DFFARX1 I_11362  ( .D(I198855), .CLK(I5694_clk), .RSTB(I198369_rst), .Q(I198346) );
nand I_11363 (I198349,I198821,I198776);
nand I_11364 (I198900,I198821,I198502);
and I_11365 (I198917,I198420,I198900);
DFFARX1 I_11366  ( .D(I198917), .CLK(I5694_clk), .RSTB(I198369_rst), .Q(I198337) );
not I_11367 (I198981_rst,I5701);
or I_11368 (I198998,I166609,I166636);
or I_11369 (I199015,I166624,I166609);
nor I_11370 (I199032,I166633,I166612);
DFFARX1 I_11371  ( .D(I199032), .CLK(I5694_clk), .RSTB(I198981_rst), .Q(I199049) );
DFFARX1 I_11372  ( .D(I199032), .CLK(I5694_clk), .RSTB(I198981_rst), .Q(I198943) );
not I_11373 (I199080,I166633);
and I_11374 (I199097,I199080,I166630);
nor I_11375 (I199114,I199097,I166636);
nor I_11376 (I199131,I166627,I166615);
DFFARX1 I_11377  ( .D(I199131), .CLK(I5694_clk), .RSTB(I198981_rst), .Q(I199148) );
not I_11378 (I199165,I199148);
DFFARX1 I_11379  ( .D(I199148), .CLK(I5694_clk), .RSTB(I198981_rst), .Q(I198952) );
nor I_11380 (I199196,I166627,I166624);
and I_11381 (I198946,I199196,I199049);
DFFARX1 I_11382  ( .D(I166639), .CLK(I5694_clk), .RSTB(I198981_rst), .Q(I199227) );
and I_11383 (I199244,I199227,I166621);
nand I_11384 (I199261,I199244,I199015);
and I_11385 (I199278,I199148,I199261);
DFFARX1 I_11386  ( .D(I199278), .CLK(I5694_clk), .RSTB(I198981_rst), .Q(I198973) );
nor I_11387 (I198970,I199244,I199114);
not I_11388 (I199323,I199244);
nor I_11389 (I199340,I198998,I199323);
nor I_11390 (I199357,I199244,I199196);
nand I_11391 (I198967,I199015,I199357);
nor I_11392 (I199388,I199244,I199165);
not I_11393 (I198964,I199244);
nand I_11394 (I198955,I199244,I199165);
DFFARX1 I_11395  ( .D(I166618), .CLK(I5694_clk), .RSTB(I198981_rst), .Q(I199433) );
and I_11396 (I199450,I199433,I199340);
or I_11397 (I199467,I198998,I199450);
DFFARX1 I_11398  ( .D(I199467), .CLK(I5694_clk), .RSTB(I198981_rst), .Q(I198958) );
nand I_11399 (I198961,I199433,I199388);
nand I_11400 (I199512,I199433,I199114);
and I_11401 (I199529,I199032,I199512);
DFFARX1 I_11402  ( .D(I199529), .CLK(I5694_clk), .RSTB(I198981_rst), .Q(I198949) );
not I_11403 (I199593_rst,I5701);
or I_11404 (I199610,I151553,I151574);
or I_11405 (I199627,I151559,I151553);
nor I_11406 (I199644,I151562,I151550);
DFFARX1 I_11407  ( .D(I199644), .CLK(I5694_clk), .RSTB(I199593_rst), .Q(I199661) );
DFFARX1 I_11408  ( .D(I199644), .CLK(I5694_clk), .RSTB(I199593_rst), .Q(I199555) );
not I_11409 (I199692,I151562);
and I_11410 (I199709,I199692,I151568);
nor I_11411 (I199726,I199709,I151574);
nor I_11412 (I199743,I151556,I151571);
DFFARX1 I_11413  ( .D(I199743), .CLK(I5694_clk), .RSTB(I199593_rst), .Q(I199760) );
not I_11414 (I199777,I199760);
DFFARX1 I_11415  ( .D(I199760), .CLK(I5694_clk), .RSTB(I199593_rst), .Q(I199564) );
nor I_11416 (I199808,I151556,I151559);
and I_11417 (I199558,I199808,I199661);
DFFARX1 I_11418  ( .D(I151547), .CLK(I5694_clk), .RSTB(I199593_rst), .Q(I199839) );
and I_11419 (I199856,I199839,I151577);
nand I_11420 (I199873,I199856,I199627);
and I_11421 (I199890,I199760,I199873);
DFFARX1 I_11422  ( .D(I199890), .CLK(I5694_clk), .RSTB(I199593_rst), .Q(I199585) );
nor I_11423 (I199582,I199856,I199726);
not I_11424 (I199935,I199856);
nor I_11425 (I199952,I199610,I199935);
nor I_11426 (I199969,I199856,I199808);
nand I_11427 (I199579,I199627,I199969);
nor I_11428 (I200000,I199856,I199777);
not I_11429 (I199576,I199856);
nand I_11430 (I199567,I199856,I199777);
DFFARX1 I_11431  ( .D(I151565), .CLK(I5694_clk), .RSTB(I199593_rst), .Q(I200045) );
and I_11432 (I200062,I200045,I199952);
or I_11433 (I200079,I199610,I200062);
DFFARX1 I_11434  ( .D(I200079), .CLK(I5694_clk), .RSTB(I199593_rst), .Q(I199570) );
nand I_11435 (I199573,I200045,I200000);
nand I_11436 (I200124,I200045,I199726);
and I_11437 (I200141,I199644,I200124);
DFFARX1 I_11438  ( .D(I200141), .CLK(I5694_clk), .RSTB(I199593_rst), .Q(I199561) );
not I_11439 (I200205_rst,I5701);
nand I_11440 (I200222,I148599,I148587);
and I_11441 (I200239,I200222,I148581);
DFFARX1 I_11442  ( .D(I200239), .CLK(I5694_clk), .RSTB(I200205_rst), .Q(I200256) );
not I_11443 (I200273,I200256);
DFFARX1 I_11444  ( .D(I200256), .CLK(I5694_clk), .RSTB(I200205_rst), .Q(I200173) );
nor I_11445 (I200304,I148578,I148587);
DFFARX1 I_11446  ( .D(I148572), .CLK(I5694_clk), .RSTB(I200205_rst), .Q(I200321) );
DFFARX1 I_11447  ( .D(I200321), .CLK(I5694_clk), .RSTB(I200205_rst), .Q(I200338) );
not I_11448 (I200176,I200338);
DFFARX1 I_11449  ( .D(I200321), .CLK(I5694_clk), .RSTB(I200205_rst), .Q(I200369) );
and I_11450 (I200170,I200256,I200369);
nand I_11451 (I200400,I148575,I148590);
and I_11452 (I200417,I200400,I148602);
DFFARX1 I_11453  ( .D(I200417), .CLK(I5694_clk), .RSTB(I200205_rst), .Q(I200434) );
nor I_11454 (I200451,I200434,I200273);
not I_11455 (I200468,I200434);
nand I_11456 (I200179,I200256,I200468);
DFFARX1 I_11457  ( .D(I148593), .CLK(I5694_clk), .RSTB(I200205_rst), .Q(I200499) );
and I_11458 (I200516,I200499,I148584);
nor I_11459 (I200533,I200516,I200434);
nor I_11460 (I200550,I200516,I200468);
nand I_11461 (I200185,I200304,I200550);
not I_11462 (I200188,I200516);
DFFARX1 I_11463  ( .D(I200516), .CLK(I5694_clk), .RSTB(I200205_rst), .Q(I200167) );
DFFARX1 I_11464  ( .D(I148596), .CLK(I5694_clk), .RSTB(I200205_rst), .Q(I200609) );
nand I_11465 (I200626,I200609,I200321);
and I_11466 (I200643,I200304,I200626);
DFFARX1 I_11467  ( .D(I200643), .CLK(I5694_clk), .RSTB(I200205_rst), .Q(I200197) );
nor I_11468 (I200194,I200609,I200516);
and I_11469 (I200688,I200609,I200451);
or I_11470 (I200705,I200304,I200688);
DFFARX1 I_11471  ( .D(I200705), .CLK(I5694_clk), .RSTB(I200205_rst), .Q(I200182) );
nand I_11472 (I200191,I200609,I200533);
not I_11473 (I200783_rst,I5701);
nand I_11474 (I200800,I143839,I143827);
and I_11475 (I200817,I200800,I143821);
DFFARX1 I_11476  ( .D(I200817), .CLK(I5694_clk), .RSTB(I200783_rst), .Q(I200834) );
not I_11477 (I200851,I200834);
DFFARX1 I_11478  ( .D(I200834), .CLK(I5694_clk), .RSTB(I200783_rst), .Q(I200751) );
nor I_11479 (I200882,I143818,I143827);
DFFARX1 I_11480  ( .D(I143812), .CLK(I5694_clk), .RSTB(I200783_rst), .Q(I200899) );
DFFARX1 I_11481  ( .D(I200899), .CLK(I5694_clk), .RSTB(I200783_rst), .Q(I200916) );
not I_11482 (I200754,I200916);
DFFARX1 I_11483  ( .D(I200899), .CLK(I5694_clk), .RSTB(I200783_rst), .Q(I200947) );
and I_11484 (I200748,I200834,I200947);
nand I_11485 (I200978,I143815,I143830);
and I_11486 (I200995,I200978,I143842);
DFFARX1 I_11487  ( .D(I200995), .CLK(I5694_clk), .RSTB(I200783_rst), .Q(I201012) );
nor I_11488 (I201029,I201012,I200851);
not I_11489 (I201046,I201012);
nand I_11490 (I200757,I200834,I201046);
DFFARX1 I_11491  ( .D(I143833), .CLK(I5694_clk), .RSTB(I200783_rst), .Q(I201077) );
and I_11492 (I201094,I201077,I143824);
nor I_11493 (I201111,I201094,I201012);
nor I_11494 (I201128,I201094,I201046);
nand I_11495 (I200763,I200882,I201128);
not I_11496 (I200766,I201094);
DFFARX1 I_11497  ( .D(I201094), .CLK(I5694_clk), .RSTB(I200783_rst), .Q(I200745) );
DFFARX1 I_11498  ( .D(I143836), .CLK(I5694_clk), .RSTB(I200783_rst), .Q(I201187) );
nand I_11499 (I201204,I201187,I200899);
and I_11500 (I201221,I200882,I201204);
DFFARX1 I_11501  ( .D(I201221), .CLK(I5694_clk), .RSTB(I200783_rst), .Q(I200775) );
nor I_11502 (I200772,I201187,I201094);
and I_11503 (I201266,I201187,I201029);
or I_11504 (I201283,I200882,I201266);
DFFARX1 I_11505  ( .D(I201283), .CLK(I5694_clk), .RSTB(I200783_rst), .Q(I200760) );
nand I_11506 (I200769,I201187,I201111);
not I_11507 (I201361_rst,I5701);
nand I_11508 (I201378,I149771,I149768);
and I_11509 (I201395,I201378,I149762);
DFFARX1 I_11510  ( .D(I201395), .CLK(I5694_clk), .RSTB(I201361_rst), .Q(I201412) );
not I_11511 (I201429,I201412);
DFFARX1 I_11512  ( .D(I201412), .CLK(I5694_clk), .RSTB(I201361_rst), .Q(I201329) );
nor I_11513 (I201460,I149783,I149768);
DFFARX1 I_11514  ( .D(I149786), .CLK(I5694_clk), .RSTB(I201361_rst), .Q(I201477) );
DFFARX1 I_11515  ( .D(I201477), .CLK(I5694_clk), .RSTB(I201361_rst), .Q(I201494) );
not I_11516 (I201332,I201494);
DFFARX1 I_11517  ( .D(I201477), .CLK(I5694_clk), .RSTB(I201361_rst), .Q(I201525) );
and I_11518 (I201326,I201412,I201525);
nand I_11519 (I201556,I149789,I149780);
and I_11520 (I201573,I201556,I149792);
DFFARX1 I_11521  ( .D(I201573), .CLK(I5694_clk), .RSTB(I201361_rst), .Q(I201590) );
nor I_11522 (I201607,I201590,I201429);
not I_11523 (I201624,I201590);
nand I_11524 (I201335,I201412,I201624);
DFFARX1 I_11525  ( .D(I149765), .CLK(I5694_clk), .RSTB(I201361_rst), .Q(I201655) );
and I_11526 (I201672,I201655,I149774);
nor I_11527 (I201689,I201672,I201590);
nor I_11528 (I201706,I201672,I201624);
nand I_11529 (I201341,I201460,I201706);
not I_11530 (I201344,I201672);
DFFARX1 I_11531  ( .D(I201672), .CLK(I5694_clk), .RSTB(I201361_rst), .Q(I201323) );
DFFARX1 I_11532  ( .D(I149777), .CLK(I5694_clk), .RSTB(I201361_rst), .Q(I201765) );
nand I_11533 (I201782,I201765,I201477);
and I_11534 (I201799,I201460,I201782);
DFFARX1 I_11535  ( .D(I201799), .CLK(I5694_clk), .RSTB(I201361_rst), .Q(I201353) );
nor I_11536 (I201350,I201765,I201672);
and I_11537 (I201844,I201765,I201607);
or I_11538 (I201861,I201460,I201844);
DFFARX1 I_11539  ( .D(I201861), .CLK(I5694_clk), .RSTB(I201361_rst), .Q(I201338) );
nand I_11540 (I201347,I201765,I201689);
not I_11541 (I201939_rst,I5701);
nand I_11542 (I201956,I197088,I197085);
and I_11543 (I201973,I201956,I197097);
DFFARX1 I_11544  ( .D(I201973), .CLK(I5694_clk), .RSTB(I201939_rst), .Q(I201990) );
not I_11545 (I202007,I201990);
DFFARX1 I_11546  ( .D(I201990), .CLK(I5694_clk), .RSTB(I201939_rst), .Q(I201907) );
nor I_11547 (I202038,I197094,I197085);
DFFARX1 I_11548  ( .D(I197100), .CLK(I5694_clk), .RSTB(I201939_rst), .Q(I202055) );
DFFARX1 I_11549  ( .D(I202055), .CLK(I5694_clk), .RSTB(I201939_rst), .Q(I202072) );
not I_11550 (I201910,I202072);
DFFARX1 I_11551  ( .D(I202055), .CLK(I5694_clk), .RSTB(I201939_rst), .Q(I202103) );
and I_11552 (I201904,I201990,I202103);
nand I_11553 (I202134,I197076,I197079);
and I_11554 (I202151,I202134,I197103);
DFFARX1 I_11555  ( .D(I202151), .CLK(I5694_clk), .RSTB(I201939_rst), .Q(I202168) );
nor I_11556 (I202185,I202168,I202007);
not I_11557 (I202202,I202168);
nand I_11558 (I201913,I201990,I202202);
DFFARX1 I_11559  ( .D(I197082), .CLK(I5694_clk), .RSTB(I201939_rst), .Q(I202233) );
and I_11560 (I202250,I202233,I197073);
nor I_11561 (I202267,I202250,I202168);
nor I_11562 (I202284,I202250,I202202);
nand I_11563 (I201919,I202038,I202284);
not I_11564 (I201922,I202250);
DFFARX1 I_11565  ( .D(I202250), .CLK(I5694_clk), .RSTB(I201939_rst), .Q(I201901) );
DFFARX1 I_11566  ( .D(I197091), .CLK(I5694_clk), .RSTB(I201939_rst), .Q(I202343) );
nand I_11567 (I202360,I202343,I202055);
and I_11568 (I202377,I202038,I202360);
DFFARX1 I_11569  ( .D(I202377), .CLK(I5694_clk), .RSTB(I201939_rst), .Q(I201931) );
nor I_11570 (I201928,I202343,I202250);
and I_11571 (I202422,I202343,I202185);
or I_11572 (I202439,I202038,I202422);
DFFARX1 I_11573  ( .D(I202439), .CLK(I5694_clk), .RSTB(I201939_rst), .Q(I201916) );
nand I_11574 (I201925,I202343,I202267);
not I_11575 (I202517_rst,I5701);
nand I_11576 (I202534,I182062,I182065);
and I_11577 (I202551,I202534,I182071);
DFFARX1 I_11578  ( .D(I202551), .CLK(I5694_clk), .RSTB(I202517_rst), .Q(I202568) );
not I_11579 (I202585,I202568);
DFFARX1 I_11580  ( .D(I202568), .CLK(I5694_clk), .RSTB(I202517_rst), .Q(I202485) );
nor I_11581 (I202616,I182083,I182065);
DFFARX1 I_11582  ( .D(I182074), .CLK(I5694_clk), .RSTB(I202517_rst), .Q(I202633) );
DFFARX1 I_11583  ( .D(I202633), .CLK(I5694_clk), .RSTB(I202517_rst), .Q(I202650) );
not I_11584 (I202488,I202650);
DFFARX1 I_11585  ( .D(I202633), .CLK(I5694_clk), .RSTB(I202517_rst), .Q(I202681) );
and I_11586 (I202482,I202568,I202681);
nand I_11587 (I202712,I182080,I182077);
and I_11588 (I202729,I202712,I182089);
DFFARX1 I_11589  ( .D(I202729), .CLK(I5694_clk), .RSTB(I202517_rst), .Q(I202746) );
nor I_11590 (I202763,I202746,I202585);
not I_11591 (I202780,I202746);
nand I_11592 (I202491,I202568,I202780);
DFFARX1 I_11593  ( .D(I182086), .CLK(I5694_clk), .RSTB(I202517_rst), .Q(I202811) );
and I_11594 (I202828,I202811,I182092);
nor I_11595 (I202845,I202828,I202746);
nor I_11596 (I202862,I202828,I202780);
nand I_11597 (I202497,I202616,I202862);
not I_11598 (I202500,I202828);
DFFARX1 I_11599  ( .D(I202828), .CLK(I5694_clk), .RSTB(I202517_rst), .Q(I202479) );
DFFARX1 I_11600  ( .D(I182068), .CLK(I5694_clk), .RSTB(I202517_rst), .Q(I202921) );
nand I_11601 (I202938,I202921,I202633);
and I_11602 (I202955,I202616,I202938);
DFFARX1 I_11603  ( .D(I202955), .CLK(I5694_clk), .RSTB(I202517_rst), .Q(I202509) );
nor I_11604 (I202506,I202921,I202828);
and I_11605 (I203000,I202921,I202763);
or I_11606 (I203017,I202616,I203000);
DFFARX1 I_11607  ( .D(I203017), .CLK(I5694_clk), .RSTB(I202517_rst), .Q(I202494) );
nand I_11608 (I202503,I202921,I202845);
not I_11609 (I203095_rst,I5701);
nand I_11610 (I203112,I180301,I180286);
and I_11611 (I203129,I203112,I180295);
DFFARX1 I_11612  ( .D(I203129), .CLK(I5694_clk), .RSTB(I203095_rst), .Q(I203146) );
not I_11613 (I203163,I203146);
DFFARX1 I_11614  ( .D(I203146), .CLK(I5694_clk), .RSTB(I203095_rst), .Q(I203063) );
nor I_11615 (I203194,I180304,I180286);
DFFARX1 I_11616  ( .D(I180283), .CLK(I5694_clk), .RSTB(I203095_rst), .Q(I203211) );
DFFARX1 I_11617  ( .D(I203211), .CLK(I5694_clk), .RSTB(I203095_rst), .Q(I203228) );
not I_11618 (I203066,I203228);
DFFARX1 I_11619  ( .D(I203211), .CLK(I5694_clk), .RSTB(I203095_rst), .Q(I203259) );
and I_11620 (I203060,I203146,I203259);
nand I_11621 (I203290,I180307,I180280);
and I_11622 (I203307,I203290,I180298);
DFFARX1 I_11623  ( .D(I203307), .CLK(I5694_clk), .RSTB(I203095_rst), .Q(I203324) );
nor I_11624 (I203341,I203324,I203163);
not I_11625 (I203358,I203324);
nand I_11626 (I203069,I203146,I203358);
DFFARX1 I_11627  ( .D(I180292), .CLK(I5694_clk), .RSTB(I203095_rst), .Q(I203389) );
and I_11628 (I203406,I203389,I180277);
nor I_11629 (I203423,I203406,I203324);
nor I_11630 (I203440,I203406,I203358);
nand I_11631 (I203075,I203194,I203440);
not I_11632 (I203078,I203406);
DFFARX1 I_11633  ( .D(I203406), .CLK(I5694_clk), .RSTB(I203095_rst), .Q(I203057) );
DFFARX1 I_11634  ( .D(I180289), .CLK(I5694_clk), .RSTB(I203095_rst), .Q(I203499) );
nand I_11635 (I203516,I203499,I203211);
and I_11636 (I203533,I203194,I203516);
DFFARX1 I_11637  ( .D(I203533), .CLK(I5694_clk), .RSTB(I203095_rst), .Q(I203087) );
nor I_11638 (I203084,I203499,I203406);
and I_11639 (I203578,I203499,I203341);
or I_11640 (I203595,I203194,I203578);
DFFARX1 I_11641  ( .D(I203595), .CLK(I5694_clk), .RSTB(I203095_rst), .Q(I203072) );
nand I_11642 (I203081,I203499,I203423);
not I_11643 (I203673_rst,I5701);
nand I_11644 (I203690,I144434,I144422);
and I_11645 (I203707,I203690,I144416);
DFFARX1 I_11646  ( .D(I203707), .CLK(I5694_clk), .RSTB(I203673_rst), .Q(I203724) );
not I_11647 (I203741,I203724);
DFFARX1 I_11648  ( .D(I203724), .CLK(I5694_clk), .RSTB(I203673_rst), .Q(I203641) );
nor I_11649 (I203772,I144413,I144422);
DFFARX1 I_11650  ( .D(I144407), .CLK(I5694_clk), .RSTB(I203673_rst), .Q(I203789) );
DFFARX1 I_11651  ( .D(I203789), .CLK(I5694_clk), .RSTB(I203673_rst), .Q(I203806) );
not I_11652 (I203644,I203806);
DFFARX1 I_11653  ( .D(I203789), .CLK(I5694_clk), .RSTB(I203673_rst), .Q(I203837) );
and I_11654 (I203638,I203724,I203837);
nand I_11655 (I203868,I144410,I144425);
and I_11656 (I203885,I203868,I144437);
DFFARX1 I_11657  ( .D(I203885), .CLK(I5694_clk), .RSTB(I203673_rst), .Q(I203902) );
nor I_11658 (I203919,I203902,I203741);
not I_11659 (I203936,I203902);
nand I_11660 (I203647,I203724,I203936);
DFFARX1 I_11661  ( .D(I144428), .CLK(I5694_clk), .RSTB(I203673_rst), .Q(I203967) );
and I_11662 (I203984,I203967,I144419);
nor I_11663 (I204001,I203984,I203902);
nor I_11664 (I204018,I203984,I203936);
nand I_11665 (I203653,I203772,I204018);
not I_11666 (I203656,I203984);
DFFARX1 I_11667  ( .D(I203984), .CLK(I5694_clk), .RSTB(I203673_rst), .Q(I203635) );
DFFARX1 I_11668  ( .D(I144431), .CLK(I5694_clk), .RSTB(I203673_rst), .Q(I204077) );
nand I_11669 (I204094,I204077,I203789);
and I_11670 (I204111,I203772,I204094);
DFFARX1 I_11671  ( .D(I204111), .CLK(I5694_clk), .RSTB(I203673_rst), .Q(I203665) );
nor I_11672 (I203662,I204077,I203984);
and I_11673 (I204156,I204077,I203919);
or I_11674 (I204173,I203772,I204156);
DFFARX1 I_11675  ( .D(I204173), .CLK(I5694_clk), .RSTB(I203673_rst), .Q(I203650) );
nand I_11676 (I203659,I204077,I204001);
not I_11677 (I204251_rst,I5701);
nand I_11678 (I204268,I179706,I179691);
and I_11679 (I204285,I204268,I179700);
DFFARX1 I_11680  ( .D(I204285), .CLK(I5694_clk), .RSTB(I204251_rst), .Q(I204302) );
not I_11681 (I204319,I204302);
DFFARX1 I_11682  ( .D(I204302), .CLK(I5694_clk), .RSTB(I204251_rst), .Q(I204219) );
nor I_11683 (I204350,I179709,I179691);
DFFARX1 I_11684  ( .D(I179688), .CLK(I5694_clk), .RSTB(I204251_rst), .Q(I204367) );
DFFARX1 I_11685  ( .D(I204367), .CLK(I5694_clk), .RSTB(I204251_rst), .Q(I204384) );
not I_11686 (I204222,I204384);
DFFARX1 I_11687  ( .D(I204367), .CLK(I5694_clk), .RSTB(I204251_rst), .Q(I204415) );
and I_11688 (I204216,I204302,I204415);
nand I_11689 (I204446,I179712,I179685);
and I_11690 (I204463,I204446,I179703);
DFFARX1 I_11691  ( .D(I204463), .CLK(I5694_clk), .RSTB(I204251_rst), .Q(I204480) );
nor I_11692 (I204497,I204480,I204319);
not I_11693 (I204514,I204480);
nand I_11694 (I204225,I204302,I204514);
DFFARX1 I_11695  ( .D(I179697), .CLK(I5694_clk), .RSTB(I204251_rst), .Q(I204545) );
and I_11696 (I204562,I204545,I179682);
nor I_11697 (I204579,I204562,I204480);
nor I_11698 (I204596,I204562,I204514);
nand I_11699 (I204231,I204350,I204596);
not I_11700 (I204234,I204562);
DFFARX1 I_11701  ( .D(I204562), .CLK(I5694_clk), .RSTB(I204251_rst), .Q(I204213) );
DFFARX1 I_11702  ( .D(I179694), .CLK(I5694_clk), .RSTB(I204251_rst), .Q(I204655) );
nand I_11703 (I204672,I204655,I204367);
and I_11704 (I204689,I204350,I204672);
DFFARX1 I_11705  ( .D(I204689), .CLK(I5694_clk), .RSTB(I204251_rst), .Q(I204243) );
nor I_11706 (I204240,I204655,I204562);
and I_11707 (I204734,I204655,I204497);
or I_11708 (I204751,I204350,I204734);
DFFARX1 I_11709  ( .D(I204751), .CLK(I5694_clk), .RSTB(I204251_rst), .Q(I204228) );
nand I_11710 (I204237,I204655,I204579);
not I_11711 (I204829_rst,I5701);
nand I_11712 (I204846,I162442,I162457);
and I_11713 (I204863,I204846,I162445);
DFFARX1 I_11714  ( .D(I204863), .CLK(I5694_clk), .RSTB(I204829_rst), .Q(I204880) );
not I_11715 (I204897,I204880);
DFFARX1 I_11716  ( .D(I204880), .CLK(I5694_clk), .RSTB(I204829_rst), .Q(I204797) );
nor I_11717 (I204928,I162454,I162457);
DFFARX1 I_11718  ( .D(I162439), .CLK(I5694_clk), .RSTB(I204829_rst), .Q(I204945) );
DFFARX1 I_11719  ( .D(I204945), .CLK(I5694_clk), .RSTB(I204829_rst), .Q(I204962) );
not I_11720 (I204800,I204962);
DFFARX1 I_11721  ( .D(I204945), .CLK(I5694_clk), .RSTB(I204829_rst), .Q(I204993) );
and I_11722 (I204794,I204880,I204993);
nand I_11723 (I205024,I162430,I162427);
and I_11724 (I205041,I205024,I162433);
DFFARX1 I_11725  ( .D(I205041), .CLK(I5694_clk), .RSTB(I204829_rst), .Q(I205058) );
nor I_11726 (I205075,I205058,I204897);
not I_11727 (I205092,I205058);
nand I_11728 (I204803,I204880,I205092);
DFFARX1 I_11729  ( .D(I162436), .CLK(I5694_clk), .RSTB(I204829_rst), .Q(I205123) );
and I_11730 (I205140,I205123,I162448);
nor I_11731 (I205157,I205140,I205058);
nor I_11732 (I205174,I205140,I205092);
nand I_11733 (I204809,I204928,I205174);
not I_11734 (I204812,I205140);
DFFARX1 I_11735  ( .D(I205140), .CLK(I5694_clk), .RSTB(I204829_rst), .Q(I204791) );
DFFARX1 I_11736  ( .D(I162451), .CLK(I5694_clk), .RSTB(I204829_rst), .Q(I205233) );
nand I_11737 (I205250,I205233,I204945);
and I_11738 (I205267,I204928,I205250);
DFFARX1 I_11739  ( .D(I205267), .CLK(I5694_clk), .RSTB(I204829_rst), .Q(I204821) );
nor I_11740 (I204818,I205233,I205140);
and I_11741 (I205312,I205233,I205075);
or I_11742 (I205329,I204928,I205312);
DFFARX1 I_11743  ( .D(I205329), .CLK(I5694_clk), .RSTB(I204829_rst), .Q(I204806) );
nand I_11744 (I204815,I205233,I205157);
not I_11745 (I205407_rst,I5701);
nand I_11746 (I205424,I152746,I152743);
and I_11747 (I205441,I205424,I152737);
DFFARX1 I_11748  ( .D(I205441), .CLK(I5694_clk), .RSTB(I205407_rst), .Q(I205458) );
not I_11749 (I205475,I205458);
DFFARX1 I_11750  ( .D(I205458), .CLK(I5694_clk), .RSTB(I205407_rst), .Q(I205375) );
nor I_11751 (I205506,I152758,I152743);
DFFARX1 I_11752  ( .D(I152761), .CLK(I5694_clk), .RSTB(I205407_rst), .Q(I205523) );
DFFARX1 I_11753  ( .D(I205523), .CLK(I5694_clk), .RSTB(I205407_rst), .Q(I205540) );
not I_11754 (I205378,I205540);
DFFARX1 I_11755  ( .D(I205523), .CLK(I5694_clk), .RSTB(I205407_rst), .Q(I205571) );
and I_11756 (I205372,I205458,I205571);
nand I_11757 (I205602,I152764,I152755);
and I_11758 (I205619,I205602,I152767);
DFFARX1 I_11759  ( .D(I205619), .CLK(I5694_clk), .RSTB(I205407_rst), .Q(I205636) );
nor I_11760 (I205653,I205636,I205475);
not I_11761 (I205670,I205636);
nand I_11762 (I205381,I205458,I205670);
DFFARX1 I_11763  ( .D(I152740), .CLK(I5694_clk), .RSTB(I205407_rst), .Q(I205701) );
and I_11764 (I205718,I205701,I152749);
nor I_11765 (I205735,I205718,I205636);
nor I_11766 (I205752,I205718,I205670);
nand I_11767 (I205387,I205506,I205752);
not I_11768 (I205390,I205718);
DFFARX1 I_11769  ( .D(I205718), .CLK(I5694_clk), .RSTB(I205407_rst), .Q(I205369) );
DFFARX1 I_11770  ( .D(I152752), .CLK(I5694_clk), .RSTB(I205407_rst), .Q(I205811) );
nand I_11771 (I205828,I205811,I205523);
and I_11772 (I205845,I205506,I205828);
DFFARX1 I_11773  ( .D(I205845), .CLK(I5694_clk), .RSTB(I205407_rst), .Q(I205399) );
nor I_11774 (I205396,I205811,I205718);
and I_11775 (I205890,I205811,I205653);
or I_11776 (I205907,I205506,I205890);
DFFARX1 I_11777  ( .D(I205907), .CLK(I5694_clk), .RSTB(I205407_rst), .Q(I205384) );
nand I_11778 (I205393,I205811,I205735);
not I_11779 (I205985_rst,I5701);
nand I_11780 (I206002,I185907,I185934);
and I_11781 (I206019,I206002,I185922);
DFFARX1 I_11782  ( .D(I206019), .CLK(I5694_clk), .RSTB(I205985_rst), .Q(I206036) );
not I_11783 (I206053,I206036);
DFFARX1 I_11784  ( .D(I206036), .CLK(I5694_clk), .RSTB(I205985_rst), .Q(I205953) );
nor I_11785 (I206084,I185910,I185934);
DFFARX1 I_11786  ( .D(I185925), .CLK(I5694_clk), .RSTB(I205985_rst), .Q(I206101) );
DFFARX1 I_11787  ( .D(I206101), .CLK(I5694_clk), .RSTB(I205985_rst), .Q(I206118) );
not I_11788 (I205956,I206118);
DFFARX1 I_11789  ( .D(I206101), .CLK(I5694_clk), .RSTB(I205985_rst), .Q(I206149) );
and I_11790 (I205950,I206036,I206149);
nand I_11791 (I206180,I185919,I185916);
and I_11792 (I206197,I206180,I185913);
DFFARX1 I_11793  ( .D(I206197), .CLK(I5694_clk), .RSTB(I205985_rst), .Q(I206214) );
nor I_11794 (I206231,I206214,I206053);
not I_11795 (I206248,I206214);
nand I_11796 (I205959,I206036,I206248);
DFFARX1 I_11797  ( .D(I185928), .CLK(I5694_clk), .RSTB(I205985_rst), .Q(I206279) );
and I_11798 (I206296,I206279,I185904);
nor I_11799 (I206313,I206296,I206214);
nor I_11800 (I206330,I206296,I206248);
nand I_11801 (I205965,I206084,I206330);
not I_11802 (I205968,I206296);
DFFARX1 I_11803  ( .D(I206296), .CLK(I5694_clk), .RSTB(I205985_rst), .Q(I205947) );
DFFARX1 I_11804  ( .D(I185931), .CLK(I5694_clk), .RSTB(I205985_rst), .Q(I206389) );
nand I_11805 (I206406,I206389,I206101);
and I_11806 (I206423,I206084,I206406);
DFFARX1 I_11807  ( .D(I206423), .CLK(I5694_clk), .RSTB(I205985_rst), .Q(I205977) );
nor I_11808 (I205974,I206389,I206296);
and I_11809 (I206468,I206389,I206231);
or I_11810 (I206485,I206084,I206468);
DFFARX1 I_11811  ( .D(I206485), .CLK(I5694_clk), .RSTB(I205985_rst), .Q(I205962) );
nand I_11812 (I205971,I206389,I206313);
not I_11813 (I206563_rst,I5701);
nand I_11814 (I206580,I195796,I195793);
and I_11815 (I206597,I206580,I195805);
DFFARX1 I_11816  ( .D(I206597), .CLK(I5694_clk), .RSTB(I206563_rst), .Q(I206614) );
not I_11817 (I206631,I206614);
DFFARX1 I_11818  ( .D(I206614), .CLK(I5694_clk), .RSTB(I206563_rst), .Q(I206531) );
nor I_11819 (I206662,I195802,I195793);
DFFARX1 I_11820  ( .D(I195808), .CLK(I5694_clk), .RSTB(I206563_rst), .Q(I206679) );
DFFARX1 I_11821  ( .D(I206679), .CLK(I5694_clk), .RSTB(I206563_rst), .Q(I206696) );
not I_11822 (I206534,I206696);
DFFARX1 I_11823  ( .D(I206679), .CLK(I5694_clk), .RSTB(I206563_rst), .Q(I206727) );
and I_11824 (I206528,I206614,I206727);
nand I_11825 (I206758,I195784,I195787);
and I_11826 (I206775,I206758,I195811);
DFFARX1 I_11827  ( .D(I206775), .CLK(I5694_clk), .RSTB(I206563_rst), .Q(I206792) );
nor I_11828 (I206809,I206792,I206631);
not I_11829 (I206826,I206792);
nand I_11830 (I206537,I206614,I206826);
DFFARX1 I_11831  ( .D(I195790), .CLK(I5694_clk), .RSTB(I206563_rst), .Q(I206857) );
and I_11832 (I206874,I206857,I195781);
nor I_11833 (I206891,I206874,I206792);
nor I_11834 (I206908,I206874,I206826);
nand I_11835 (I206543,I206662,I206908);
not I_11836 (I206546,I206874);
DFFARX1 I_11837  ( .D(I206874), .CLK(I5694_clk), .RSTB(I206563_rst), .Q(I206525) );
DFFARX1 I_11838  ( .D(I195799), .CLK(I5694_clk), .RSTB(I206563_rst), .Q(I206967) );
nand I_11839 (I206984,I206967,I206679);
and I_11840 (I207001,I206662,I206984);
DFFARX1 I_11841  ( .D(I207001), .CLK(I5694_clk), .RSTB(I206563_rst), .Q(I206555) );
nor I_11842 (I206552,I206967,I206874);
and I_11843 (I207046,I206967,I206809);
or I_11844 (I207063,I206662,I207046);
DFFARX1 I_11845  ( .D(I207063), .CLK(I5694_clk), .RSTB(I206563_rst), .Q(I206540) );
nand I_11846 (I206549,I206967,I206891);
not I_11847 (I207141_rst,I5701);
or I_11848 (I207158,I189222,I189219);
or I_11849 (I207175,I189234,I189222);
nor I_11850 (I207192,I189249,I189225);
not I_11851 (I207209,I207192);
DFFARX1 I_11852  ( .D(I207192), .CLK(I5694_clk), .RSTB(I207141_rst), .Q(I207109) );
nand I_11853 (I207240,I207192,I207158);
not I_11854 (I207257,I189249);
and I_11855 (I207274,I207257,I189243);
nor I_11856 (I207291,I207274,I189219);
nor I_11857 (I207308,I189237,I189246);
DFFARX1 I_11858  ( .D(I207308), .CLK(I5694_clk), .RSTB(I207141_rst), .Q(I207325) );
nor I_11859 (I207342,I207325,I207209);
not I_11860 (I207359,I207325);
nand I_11861 (I207115,I207192,I207359);
DFFARX1 I_11862  ( .D(I207325), .CLK(I5694_clk), .RSTB(I207141_rst), .Q(I207106) );
nor I_11863 (I207404,I189237,I189234);
nand I_11864 (I207421,I207175,I207404);
nor I_11865 (I207130,I207158,I207404);
and I_11866 (I207452,I207404,I207342);
or I_11867 (I207469,I207291,I207452);
DFFARX1 I_11868  ( .D(I207469), .CLK(I5694_clk), .RSTB(I207141_rst), .Q(I207118) );
DFFARX1 I_11869  ( .D(I189231), .CLK(I5694_clk), .RSTB(I207141_rst), .Q(I207500) );
and I_11870 (I207517,I207500,I189228);
not I_11871 (I207124,I207517);
DFFARX1 I_11872  ( .D(I207517), .CLK(I5694_clk), .RSTB(I207141_rst), .Q(I207548) );
not I_11873 (I207112,I207548);
and I_11874 (I207579,I207517,I207240);
DFFARX1 I_11875  ( .D(I207579), .CLK(I5694_clk), .RSTB(I207141_rst), .Q(I207103) );
DFFARX1 I_11876  ( .D(I189240), .CLK(I5694_clk), .RSTB(I207141_rst), .Q(I207610) );
and I_11877 (I207627,I207610,I207421);
DFFARX1 I_11878  ( .D(I207627), .CLK(I5694_clk), .RSTB(I207141_rst), .Q(I207133) );
nor I_11879 (I207658,I207610,I207517);
nand I_11880 (I207127,I207291,I207658);
nor I_11881 (I207689,I207610,I207359);
nand I_11882 (I207121,I207175,I207689);
not I_11883 (I207753_rst,I5701);
or I_11884 (I207770,I157762,I157756);
or I_11885 (I207787,I157765,I157762);
nor I_11886 (I207804,I157759,I157741);
not I_11887 (I207821,I207804);
DFFARX1 I_11888  ( .D(I207804), .CLK(I5694_clk), .RSTB(I207753_rst), .Q(I207721) );
nand I_11889 (I207852,I207804,I207770);
not I_11890 (I207869,I157759);
and I_11891 (I207886,I207869,I157738);
nor I_11892 (I207903,I207886,I157756);
nor I_11893 (I207920,I157753,I157735);
DFFARX1 I_11894  ( .D(I207920), .CLK(I5694_clk), .RSTB(I207753_rst), .Q(I207937) );
nor I_11895 (I207954,I207937,I207821);
not I_11896 (I207971,I207937);
nand I_11897 (I207727,I207804,I207971);
DFFARX1 I_11898  ( .D(I207937), .CLK(I5694_clk), .RSTB(I207753_rst), .Q(I207718) );
nor I_11899 (I208016,I157753,I157765);
nand I_11900 (I208033,I207787,I208016);
nor I_11901 (I207742,I207770,I208016);
and I_11902 (I208064,I208016,I207954);
or I_11903 (I208081,I207903,I208064);
DFFARX1 I_11904  ( .D(I208081), .CLK(I5694_clk), .RSTB(I207753_rst), .Q(I207730) );
DFFARX1 I_11905  ( .D(I157747), .CLK(I5694_clk), .RSTB(I207753_rst), .Q(I208112) );
and I_11906 (I208129,I208112,I157750);
not I_11907 (I207736,I208129);
DFFARX1 I_11908  ( .D(I208129), .CLK(I5694_clk), .RSTB(I207753_rst), .Q(I208160) );
not I_11909 (I207724,I208160);
and I_11910 (I208191,I208129,I207852);
DFFARX1 I_11911  ( .D(I208191), .CLK(I5694_clk), .RSTB(I207753_rst), .Q(I207715) );
DFFARX1 I_11912  ( .D(I157744), .CLK(I5694_clk), .RSTB(I207753_rst), .Q(I208222) );
and I_11913 (I208239,I208222,I208033);
DFFARX1 I_11914  ( .D(I208239), .CLK(I5694_clk), .RSTB(I207753_rst), .Q(I207745) );
nor I_11915 (I208270,I208222,I208129);
nand I_11916 (I207739,I207903,I208270);
nor I_11917 (I208301,I208222,I207971);
nand I_11918 (I207733,I207787,I208301);
not I_11919 (I208365_rst,I5701);
or I_11920 (I208382,I145026,I145032);
or I_11921 (I208399,I145029,I145026);
nor I_11922 (I208416,I145002,I145020);
not I_11923 (I208433,I208416);
DFFARX1 I_11924  ( .D(I208416), .CLK(I5694_clk), .RSTB(I208365_rst), .Q(I208333) );
nand I_11925 (I208464,I208416,I208382);
not I_11926 (I208481,I145002);
and I_11927 (I208498,I208481,I145014);
nor I_11928 (I208515,I208498,I145032);
nor I_11929 (I208532,I145017,I145005);
DFFARX1 I_11930  ( .D(I208532), .CLK(I5694_clk), .RSTB(I208365_rst), .Q(I208549) );
nor I_11931 (I208566,I208549,I208433);
not I_11932 (I208583,I208549);
nand I_11933 (I208339,I208416,I208583);
DFFARX1 I_11934  ( .D(I208549), .CLK(I5694_clk), .RSTB(I208365_rst), .Q(I208330) );
nor I_11935 (I208628,I145017,I145029);
nand I_11936 (I208645,I208399,I208628);
nor I_11937 (I208354,I208382,I208628);
and I_11938 (I208676,I208628,I208566);
or I_11939 (I208693,I208515,I208676);
DFFARX1 I_11940  ( .D(I208693), .CLK(I5694_clk), .RSTB(I208365_rst), .Q(I208342) );
DFFARX1 I_11941  ( .D(I145008), .CLK(I5694_clk), .RSTB(I208365_rst), .Q(I208724) );
and I_11942 (I208741,I208724,I145023);
not I_11943 (I208348,I208741);
DFFARX1 I_11944  ( .D(I208741), .CLK(I5694_clk), .RSTB(I208365_rst), .Q(I208772) );
not I_11945 (I208336,I208772);
and I_11946 (I208803,I208741,I208464);
DFFARX1 I_11947  ( .D(I208803), .CLK(I5694_clk), .RSTB(I208365_rst), .Q(I208327) );
DFFARX1 I_11948  ( .D(I145011), .CLK(I5694_clk), .RSTB(I208365_rst), .Q(I208834) );
and I_11949 (I208851,I208834,I208645);
DFFARX1 I_11950  ( .D(I208851), .CLK(I5694_clk), .RSTB(I208365_rst), .Q(I208357) );
nor I_11951 (I208882,I208834,I208741);
nand I_11952 (I208351,I208515,I208882);
nor I_11953 (I208913,I208834,I208583);
nand I_11954 (I208345,I208399,I208913);
not I_11955 (I208977_rst,I5701);
or I_11956 (I208994,I146213,I146207);
or I_11957 (I209011,I146201,I146213);
nor I_11958 (I209028,I146222,I146210);
or I_11959 (I208966,I209028,I208994);
not I_11960 (I209059,I146222);
and I_11961 (I209076,I209059,I146195);
nor I_11962 (I209093,I209076,I146207);
not I_11963 (I209110,I209093);
nor I_11964 (I209127,I146198,I146192);
DFFARX1 I_11965  ( .D(I209127), .CLK(I5694_clk), .RSTB(I208977_rst), .Q(I209144) );
nor I_11966 (I209161,I209144,I209093);
nand I_11967 (I208951,I208994,I209161);
nor I_11968 (I209192,I209144,I209110);
not I_11969 (I208948,I209144);
nor I_11970 (I209223,I146198,I146201);
or I_11971 (I208960,I208994,I209223);
DFFARX1 I_11972  ( .D(I146219), .CLK(I5694_clk), .RSTB(I208977_rst), .Q(I209254) );
and I_11973 (I209271,I209254,I146216);
nor I_11974 (I209288,I209271,I209144);
DFFARX1 I_11975  ( .D(I209288), .CLK(I5694_clk), .RSTB(I208977_rst), .Q(I208954) );
nor I_11976 (I208969,I209271,I209223);
not I_11977 (I209333,I209271);
nor I_11978 (I209350,I209011,I209333);
nand I_11979 (I208939,I209271,I209110);
DFFARX1 I_11980  ( .D(I146204), .CLK(I5694_clk), .RSTB(I208977_rst), .Q(I209381) );
nor I_11981 (I208957,I209381,I209011);
not I_11982 (I209412,I209381);
and I_11983 (I209429,I209223,I209412);
nor I_11984 (I208963,I209028,I209429);
and I_11985 (I209460,I209381,I209350);
or I_11986 (I209477,I209028,I209460);
DFFARX1 I_11987  ( .D(I209477), .CLK(I5694_clk), .RSTB(I208977_rst), .Q(I208942) );
nand I_11988 (I208945,I209381,I209192);
not I_11989 (I209555_rst,I5701);
nand I_11990 (I209572,I190563,I190569);
and I_11991 (I209589,I209572,I190551);
DFFARX1 I_11992  ( .D(I209589), .CLK(I5694_clk), .RSTB(I209555_rst), .Q(I209606) );
nor I_11993 (I209623,I190545,I190569);
nor I_11994 (I209640,I209623,I209606);
not I_11995 (I209538,I209623);
DFFARX1 I_11996  ( .D(I190575), .CLK(I5694_clk), .RSTB(I209555_rst), .Q(I209671) );
not I_11997 (I209688,I209671);
nor I_11998 (I209705,I209623,I209688);
nand I_11999 (I209541,I209671,I209640);
DFFARX1 I_12000  ( .D(I209671), .CLK(I5694_clk), .RSTB(I209555_rst), .Q(I209523) );
nand I_12001 (I209750,I190566,I190557);
and I_12002 (I209767,I209750,I190560);
DFFARX1 I_12003  ( .D(I209767), .CLK(I5694_clk), .RSTB(I209555_rst), .Q(I209784) );
nor I_12004 (I209544,I209784,I209606);
nand I_12005 (I209535,I209784,I209705);
DFFARX1 I_12006  ( .D(I190572), .CLK(I5694_clk), .RSTB(I209555_rst), .Q(I209829) );
and I_12007 (I209846,I209829,I190548);
DFFARX1 I_12008  ( .D(I209846), .CLK(I5694_clk), .RSTB(I209555_rst), .Q(I209863) );
not I_12009 (I209526,I209863);
nand I_12010 (I209894,I209846,I209784);
and I_12011 (I209911,I209606,I209894);
DFFARX1 I_12012  ( .D(I209911), .CLK(I5694_clk), .RSTB(I209555_rst), .Q(I209517) );
DFFARX1 I_12013  ( .D(I190554), .CLK(I5694_clk), .RSTB(I209555_rst), .Q(I209942) );
nand I_12014 (I209959,I209942,I209606);
and I_12015 (I209976,I209784,I209959);
DFFARX1 I_12016  ( .D(I209976), .CLK(I5694_clk), .RSTB(I209555_rst), .Q(I209547) );
not I_12017 (I210007,I209942);
nor I_12018 (I210024,I209623,I210007);
and I_12019 (I210041,I209942,I210024);
or I_12020 (I210058,I209846,I210041);
DFFARX1 I_12021  ( .D(I210058), .CLK(I5694_clk), .RSTB(I209555_rst), .Q(I209532) );
nand I_12022 (I209529,I209942,I209688);
DFFARX1 I_12023  ( .D(I209942), .CLK(I5694_clk), .RSTB(I209555_rst), .Q(I209520) );
not I_12024 (I210150_rst,I5701);
nand I_12025 (I210167,I187248,I187254);
and I_12026 (I210184,I210167,I187236);
DFFARX1 I_12027  ( .D(I210184), .CLK(I5694_clk), .RSTB(I210150_rst), .Q(I210201) );
nor I_12028 (I210218,I187230,I187254);
nor I_12029 (I210235,I210218,I210201);
not I_12030 (I210133,I210218);
DFFARX1 I_12031  ( .D(I187260), .CLK(I5694_clk), .RSTB(I210150_rst), .Q(I210266) );
not I_12032 (I210283,I210266);
nor I_12033 (I210300,I210218,I210283);
nand I_12034 (I210136,I210266,I210235);
DFFARX1 I_12035  ( .D(I210266), .CLK(I5694_clk), .RSTB(I210150_rst), .Q(I210118) );
nand I_12036 (I210345,I187251,I187242);
and I_12037 (I210362,I210345,I187245);
DFFARX1 I_12038  ( .D(I210362), .CLK(I5694_clk), .RSTB(I210150_rst), .Q(I210379) );
nor I_12039 (I210139,I210379,I210201);
nand I_12040 (I210130,I210379,I210300);
DFFARX1 I_12041  ( .D(I187257), .CLK(I5694_clk), .RSTB(I210150_rst), .Q(I210424) );
and I_12042 (I210441,I210424,I187233);
DFFARX1 I_12043  ( .D(I210441), .CLK(I5694_clk), .RSTB(I210150_rst), .Q(I210458) );
not I_12044 (I210121,I210458);
nand I_12045 (I210489,I210441,I210379);
and I_12046 (I210506,I210201,I210489);
DFFARX1 I_12047  ( .D(I210506), .CLK(I5694_clk), .RSTB(I210150_rst), .Q(I210112) );
DFFARX1 I_12048  ( .D(I187239), .CLK(I5694_clk), .RSTB(I210150_rst), .Q(I210537) );
nand I_12049 (I210554,I210537,I210201);
and I_12050 (I210571,I210379,I210554);
DFFARX1 I_12051  ( .D(I210571), .CLK(I5694_clk), .RSTB(I210150_rst), .Q(I210142) );
not I_12052 (I210602,I210537);
nor I_12053 (I210619,I210218,I210602);
and I_12054 (I210636,I210537,I210619);
or I_12055 (I210653,I210441,I210636);
DFFARX1 I_12056  ( .D(I210653), .CLK(I5694_clk), .RSTB(I210150_rst), .Q(I210127) );
nand I_12057 (I210124,I210537,I210283);
DFFARX1 I_12058  ( .D(I210537), .CLK(I5694_clk), .RSTB(I210150_rst), .Q(I210115) );
not I_12059 (I210745_rst,I5701);
nand I_12060 (I210762,I195153,I195165);
and I_12061 (I210779,I210762,I195147);
DFFARX1 I_12062  ( .D(I210779), .CLK(I5694_clk), .RSTB(I210745_rst), .Q(I210796) );
nor I_12063 (I210813,I195159,I195165);
nor I_12064 (I210830,I210813,I210796);
not I_12065 (I210728,I210813);
DFFARX1 I_12066  ( .D(I195144), .CLK(I5694_clk), .RSTB(I210745_rst), .Q(I210861) );
not I_12067 (I210878,I210861);
nor I_12068 (I210895,I210813,I210878);
nand I_12069 (I210731,I210861,I210830);
DFFARX1 I_12070  ( .D(I210861), .CLK(I5694_clk), .RSTB(I210745_rst), .Q(I210713) );
nand I_12071 (I210940,I195135,I195150);
and I_12072 (I210957,I210940,I195141);
DFFARX1 I_12073  ( .D(I210957), .CLK(I5694_clk), .RSTB(I210745_rst), .Q(I210974) );
nor I_12074 (I210734,I210974,I210796);
nand I_12075 (I210725,I210974,I210895);
DFFARX1 I_12076  ( .D(I195162), .CLK(I5694_clk), .RSTB(I210745_rst), .Q(I211019) );
and I_12077 (I211036,I211019,I195156);
DFFARX1 I_12078  ( .D(I211036), .CLK(I5694_clk), .RSTB(I210745_rst), .Q(I211053) );
not I_12079 (I210716,I211053);
nand I_12080 (I211084,I211036,I210974);
and I_12081 (I211101,I210796,I211084);
DFFARX1 I_12082  ( .D(I211101), .CLK(I5694_clk), .RSTB(I210745_rst), .Q(I210707) );
DFFARX1 I_12083  ( .D(I195138), .CLK(I5694_clk), .RSTB(I210745_rst), .Q(I211132) );
nand I_12084 (I211149,I211132,I210796);
and I_12085 (I211166,I210974,I211149);
DFFARX1 I_12086  ( .D(I211166), .CLK(I5694_clk), .RSTB(I210745_rst), .Q(I210737) );
not I_12087 (I211197,I211132);
nor I_12088 (I211214,I210813,I211197);
and I_12089 (I211231,I211132,I211214);
or I_12090 (I211248,I211036,I211231);
DFFARX1 I_12091  ( .D(I211248), .CLK(I5694_clk), .RSTB(I210745_rst), .Q(I210722) );
nand I_12092 (I210719,I211132,I210878);
DFFARX1 I_12093  ( .D(I211132), .CLK(I5694_clk), .RSTB(I210745_rst), .Q(I210710) );
not I_12094 (I211340_rst,I5701);
nand I_12095 (I211357,I173733,I173745);
and I_12096 (I211374,I211357,I173724);
DFFARX1 I_12097  ( .D(I211374), .CLK(I5694_clk), .RSTB(I211340_rst), .Q(I211391) );
nor I_12098 (I211408,I173715,I173745);
nor I_12099 (I211425,I211408,I211391);
not I_12100 (I211323,I211408);
DFFARX1 I_12101  ( .D(I173727), .CLK(I5694_clk), .RSTB(I211340_rst), .Q(I211456) );
not I_12102 (I211473,I211456);
nor I_12103 (I211490,I211408,I211473);
nand I_12104 (I211326,I211456,I211425);
DFFARX1 I_12105  ( .D(I211456), .CLK(I5694_clk), .RSTB(I211340_rst), .Q(I211308) );
nand I_12106 (I211535,I173742,I173730);
and I_12107 (I211552,I211535,I173718);
DFFARX1 I_12108  ( .D(I211552), .CLK(I5694_clk), .RSTB(I211340_rst), .Q(I211569) );
nor I_12109 (I211329,I211569,I211391);
nand I_12110 (I211320,I211569,I211490);
DFFARX1 I_12111  ( .D(I173736), .CLK(I5694_clk), .RSTB(I211340_rst), .Q(I211614) );
and I_12112 (I211631,I211614,I173721);
DFFARX1 I_12113  ( .D(I211631), .CLK(I5694_clk), .RSTB(I211340_rst), .Q(I211648) );
not I_12114 (I211311,I211648);
nand I_12115 (I211679,I211631,I211569);
and I_12116 (I211696,I211391,I211679);
DFFARX1 I_12117  ( .D(I211696), .CLK(I5694_clk), .RSTB(I211340_rst), .Q(I211302) );
DFFARX1 I_12118  ( .D(I173739), .CLK(I5694_clk), .RSTB(I211340_rst), .Q(I211727) );
nand I_12119 (I211744,I211727,I211391);
and I_12120 (I211761,I211569,I211744);
DFFARX1 I_12121  ( .D(I211761), .CLK(I5694_clk), .RSTB(I211340_rst), .Q(I211332) );
not I_12122 (I211792,I211727);
nor I_12123 (I211809,I211408,I211792);
and I_12124 (I211826,I211727,I211809);
or I_12125 (I211843,I211631,I211826);
DFFARX1 I_12126  ( .D(I211843), .CLK(I5694_clk), .RSTB(I211340_rst), .Q(I211317) );
nand I_12127 (I211314,I211727,I211473);
DFFARX1 I_12128  ( .D(I211727), .CLK(I5694_clk), .RSTB(I211340_rst), .Q(I211305) );
not I_12129 (I211935_rst,I5701);
nand I_12130 (I211952,I167910,I167922);
and I_12131 (I211969,I211952,I167931);
DFFARX1 I_12132  ( .D(I211969), .CLK(I5694_clk), .RSTB(I211935_rst), .Q(I211986) );
nor I_12133 (I212003,I167925,I167922);
nor I_12134 (I212020,I212003,I211986);
not I_12135 (I211918,I212003);
DFFARX1 I_12136  ( .D(I167919), .CLK(I5694_clk), .RSTB(I211935_rst), .Q(I212051) );
not I_12137 (I212068,I212051);
nor I_12138 (I212085,I212003,I212068);
nand I_12139 (I211921,I212051,I212020);
DFFARX1 I_12140  ( .D(I212051), .CLK(I5694_clk), .RSTB(I211935_rst), .Q(I211903) );
nand I_12141 (I212130,I167916,I167913);
and I_12142 (I212147,I212130,I167904);
DFFARX1 I_12143  ( .D(I212147), .CLK(I5694_clk), .RSTB(I211935_rst), .Q(I212164) );
nor I_12144 (I211924,I212164,I211986);
nand I_12145 (I211915,I212164,I212085);
DFFARX1 I_12146  ( .D(I167928), .CLK(I5694_clk), .RSTB(I211935_rst), .Q(I212209) );
and I_12147 (I212226,I212209,I167907);
DFFARX1 I_12148  ( .D(I212226), .CLK(I5694_clk), .RSTB(I211935_rst), .Q(I212243) );
not I_12149 (I211906,I212243);
nand I_12150 (I212274,I212226,I212164);
and I_12151 (I212291,I211986,I212274);
DFFARX1 I_12152  ( .D(I212291), .CLK(I5694_clk), .RSTB(I211935_rst), .Q(I211897) );
DFFARX1 I_12153  ( .D(I167901), .CLK(I5694_clk), .RSTB(I211935_rst), .Q(I212322) );
nand I_12154 (I212339,I212322,I211986);
and I_12155 (I212356,I212164,I212339);
DFFARX1 I_12156  ( .D(I212356), .CLK(I5694_clk), .RSTB(I211935_rst), .Q(I211927) );
not I_12157 (I212387,I212322);
nor I_12158 (I212404,I212003,I212387);
and I_12159 (I212421,I212322,I212404);
or I_12160 (I212438,I212226,I212421);
DFFARX1 I_12161  ( .D(I212438), .CLK(I5694_clk), .RSTB(I211935_rst), .Q(I211912) );
nand I_12162 (I211909,I212322,I212068);
DFFARX1 I_12163  ( .D(I212322), .CLK(I5694_clk), .RSTB(I211935_rst), .Q(I211900) );
not I_12164 (I212530_rst,I5701);
nand I_12165 (I212547,I158382,I158373);
and I_12166 (I212564,I212547,I158391);
DFFARX1 I_12167  ( .D(I212564), .CLK(I5694_clk), .RSTB(I212530_rst), .Q(I212581) );
nor I_12168 (I212598,I158388,I158373);
nor I_12169 (I212615,I212598,I212581);
not I_12170 (I212513,I212598);
DFFARX1 I_12171  ( .D(I158370), .CLK(I5694_clk), .RSTB(I212530_rst), .Q(I212646) );
not I_12172 (I212663,I212646);
nor I_12173 (I212680,I212598,I212663);
nand I_12174 (I212516,I212646,I212615);
DFFARX1 I_12175  ( .D(I212646), .CLK(I5694_clk), .RSTB(I212530_rst), .Q(I212498) );
nand I_12176 (I212725,I158379,I158394);
and I_12177 (I212742,I212725,I158385);
DFFARX1 I_12178  ( .D(I212742), .CLK(I5694_clk), .RSTB(I212530_rst), .Q(I212759) );
nor I_12179 (I212519,I212759,I212581);
nand I_12180 (I212510,I212759,I212680);
DFFARX1 I_12181  ( .D(I158367), .CLK(I5694_clk), .RSTB(I212530_rst), .Q(I212804) );
and I_12182 (I212821,I212804,I158376);
DFFARX1 I_12183  ( .D(I212821), .CLK(I5694_clk), .RSTB(I212530_rst), .Q(I212838) );
not I_12184 (I212501,I212838);
nand I_12185 (I212869,I212821,I212759);
and I_12186 (I212886,I212581,I212869);
DFFARX1 I_12187  ( .D(I212886), .CLK(I5694_clk), .RSTB(I212530_rst), .Q(I212492) );
DFFARX1 I_12188  ( .D(I158364), .CLK(I5694_clk), .RSTB(I212530_rst), .Q(I212917) );
nand I_12189 (I212934,I212917,I212581);
and I_12190 (I212951,I212759,I212934);
DFFARX1 I_12191  ( .D(I212951), .CLK(I5694_clk), .RSTB(I212530_rst), .Q(I212522) );
not I_12192 (I212982,I212917);
nor I_12193 (I212999,I212598,I212982);
and I_12194 (I213016,I212917,I212999);
or I_12195 (I213033,I212821,I213016);
DFFARX1 I_12196  ( .D(I213033), .CLK(I5694_clk), .RSTB(I212530_rst), .Q(I212507) );
nand I_12197 (I212504,I212917,I212663);
DFFARX1 I_12198  ( .D(I212917), .CLK(I5694_clk), .RSTB(I212530_rst), .Q(I212495) );
not I_12199 (I213125_rst,I5701);
nand I_12200 (I213142,I203084,I203087);
and I_12201 (I213159,I213142,I203081);
DFFARX1 I_12202  ( .D(I213159), .CLK(I5694_clk), .RSTB(I213125_rst), .Q(I213176) );
nor I_12203 (I213193,I203078,I203087);
nor I_12204 (I213210,I213193,I213176);
not I_12205 (I213108,I213193);
DFFARX1 I_12206  ( .D(I203060), .CLK(I5694_clk), .RSTB(I213125_rst), .Q(I213241) );
not I_12207 (I213258,I213241);
nor I_12208 (I213275,I213193,I213258);
nand I_12209 (I213111,I213241,I213210);
DFFARX1 I_12210  ( .D(I213241), .CLK(I5694_clk), .RSTB(I213125_rst), .Q(I213093) );
nand I_12211 (I213320,I203069,I203066);
and I_12212 (I213337,I213320,I203075);
DFFARX1 I_12213  ( .D(I213337), .CLK(I5694_clk), .RSTB(I213125_rst), .Q(I213354) );
nor I_12214 (I213114,I213354,I213176);
nand I_12215 (I213105,I213354,I213275);
DFFARX1 I_12216  ( .D(I203057), .CLK(I5694_clk), .RSTB(I213125_rst), .Q(I213399) );
and I_12217 (I213416,I213399,I203072);
DFFARX1 I_12218  ( .D(I213416), .CLK(I5694_clk), .RSTB(I213125_rst), .Q(I213433) );
not I_12219 (I213096,I213433);
nand I_12220 (I213464,I213416,I213354);
and I_12221 (I213481,I213176,I213464);
DFFARX1 I_12222  ( .D(I213481), .CLK(I5694_clk), .RSTB(I213125_rst), .Q(I213087) );
DFFARX1 I_12223  ( .D(I203063), .CLK(I5694_clk), .RSTB(I213125_rst), .Q(I213512) );
nand I_12224 (I213529,I213512,I213176);
and I_12225 (I213546,I213354,I213529);
DFFARX1 I_12226  ( .D(I213546), .CLK(I5694_clk), .RSTB(I213125_rst), .Q(I213117) );
not I_12227 (I213577,I213512);
nor I_12228 (I213594,I213193,I213577);
and I_12229 (I213611,I213512,I213594);
or I_12230 (I213628,I213416,I213611);
DFFARX1 I_12231  ( .D(I213628), .CLK(I5694_clk), .RSTB(I213125_rst), .Q(I213102) );
nand I_12232 (I213099,I213512,I213258);
DFFARX1 I_12233  ( .D(I213512), .CLK(I5694_clk), .RSTB(I213125_rst), .Q(I213090) );
not I_12234 (I213720_rst,I5701);
nand I_12235 (I213737,I170494,I170506);
and I_12236 (I213754,I213737,I170515);
DFFARX1 I_12237  ( .D(I213754), .CLK(I5694_clk), .RSTB(I213720_rst), .Q(I213771) );
nor I_12238 (I213788,I170509,I170506);
nor I_12239 (I213805,I213788,I213771);
not I_12240 (I213703,I213788);
DFFARX1 I_12241  ( .D(I170503), .CLK(I5694_clk), .RSTB(I213720_rst), .Q(I213836) );
not I_12242 (I213853,I213836);
nor I_12243 (I213870,I213788,I213853);
nand I_12244 (I213706,I213836,I213805);
DFFARX1 I_12245  ( .D(I213836), .CLK(I5694_clk), .RSTB(I213720_rst), .Q(I213688) );
nand I_12246 (I213915,I170500,I170497);
and I_12247 (I213932,I213915,I170488);
DFFARX1 I_12248  ( .D(I213932), .CLK(I5694_clk), .RSTB(I213720_rst), .Q(I213949) );
nor I_12249 (I213709,I213949,I213771);
nand I_12250 (I213700,I213949,I213870);
DFFARX1 I_12251  ( .D(I170512), .CLK(I5694_clk), .RSTB(I213720_rst), .Q(I213994) );
and I_12252 (I214011,I213994,I170491);
DFFARX1 I_12253  ( .D(I214011), .CLK(I5694_clk), .RSTB(I213720_rst), .Q(I214028) );
not I_12254 (I213691,I214028);
nand I_12255 (I214059,I214011,I213949);
and I_12256 (I214076,I213771,I214059);
DFFARX1 I_12257  ( .D(I214076), .CLK(I5694_clk), .RSTB(I213720_rst), .Q(I213682) );
DFFARX1 I_12258  ( .D(I170485), .CLK(I5694_clk), .RSTB(I213720_rst), .Q(I214107) );
nand I_12259 (I214124,I214107,I213771);
and I_12260 (I214141,I213949,I214124);
DFFARX1 I_12261  ( .D(I214141), .CLK(I5694_clk), .RSTB(I213720_rst), .Q(I213712) );
not I_12262 (I214172,I214107);
nor I_12263 (I214189,I213788,I214172);
and I_12264 (I214206,I214107,I214189);
or I_12265 (I214223,I214011,I214206);
DFFARX1 I_12266  ( .D(I214223), .CLK(I5694_clk), .RSTB(I213720_rst), .Q(I213697) );
nand I_12267 (I213694,I214107,I213853);
DFFARX1 I_12268  ( .D(I214107), .CLK(I5694_clk), .RSTB(I213720_rst), .Q(I213685) );
not I_12269 (I214315_rst,I5701);
nand I_12270 (I214332,I174381,I174402);
and I_12271 (I214349,I214332,I174387);
DFFARX1 I_12272  ( .D(I214349), .CLK(I5694_clk), .RSTB(I214315_rst), .Q(I214366) );
nor I_12273 (I214383,I174405,I174402);
DFFARX1 I_12274  ( .D(I174408), .CLK(I5694_clk), .RSTB(I214315_rst), .Q(I214400) );
nand I_12275 (I214417,I214400,I214383);
DFFARX1 I_12276  ( .D(I214400), .CLK(I5694_clk), .RSTB(I214315_rst), .Q(I214286) );
nand I_12277 (I214448,I174378,I174390);
and I_12278 (I214465,I214448,I174399);
DFFARX1 I_12279  ( .D(I214465), .CLK(I5694_clk), .RSTB(I214315_rst), .Q(I214482) );
not I_12280 (I214499,I214482);
nor I_12281 (I214516,I214366,I214499);
and I_12282 (I214533,I214383,I214516);
and I_12283 (I214550,I214482,I214417);
DFFARX1 I_12284  ( .D(I214550), .CLK(I5694_clk), .RSTB(I214315_rst), .Q(I214283) );
DFFARX1 I_12285  ( .D(I214482), .CLK(I5694_clk), .RSTB(I214315_rst), .Q(I214277) );
DFFARX1 I_12286  ( .D(I174393), .CLK(I5694_clk), .RSTB(I214315_rst), .Q(I214595) );
and I_12287 (I214612,I214595,I174396);
nand I_12288 (I214629,I214612,I214482);
nor I_12289 (I214304,I214612,I214383);
not I_12290 (I214660,I214612);
nor I_12291 (I214677,I214366,I214660);
nand I_12292 (I214295,I214400,I214677);
nand I_12293 (I214289,I214482,I214660);
or I_12294 (I214722,I214612,I214533);
DFFARX1 I_12295  ( .D(I214722), .CLK(I5694_clk), .RSTB(I214315_rst), .Q(I214292) );
DFFARX1 I_12296  ( .D(I174384), .CLK(I5694_clk), .RSTB(I214315_rst), .Q(I214753) );
and I_12297 (I214770,I214753,I214629);
DFFARX1 I_12298  ( .D(I214770), .CLK(I5694_clk), .RSTB(I214315_rst), .Q(I214307) );
nor I_12299 (I214801,I214753,I214366);
nand I_12300 (I214301,I214612,I214801);
not I_12301 (I214298,I214753);
DFFARX1 I_12302  ( .D(I214753), .CLK(I5694_clk), .RSTB(I214315_rst), .Q(I214846) );
and I_12303 (I214280,I214753,I214846);
not I_12304 (I214910_rst,I5701);
nand I_12305 (I214927,I169866,I169842);
and I_12306 (I214944,I214927,I169851);
DFFARX1 I_12307  ( .D(I214944), .CLK(I5694_clk), .RSTB(I214910_rst), .Q(I214961) );
nor I_12308 (I214978,I169845,I169842);
DFFARX1 I_12309  ( .D(I169860), .CLK(I5694_clk), .RSTB(I214910_rst), .Q(I214995) );
nand I_12310 (I215012,I214995,I214978);
DFFARX1 I_12311  ( .D(I214995), .CLK(I5694_clk), .RSTB(I214910_rst), .Q(I214881) );
nand I_12312 (I215043,I169854,I169869);
and I_12313 (I215060,I215043,I169848);
DFFARX1 I_12314  ( .D(I215060), .CLK(I5694_clk), .RSTB(I214910_rst), .Q(I215077) );
not I_12315 (I215094,I215077);
nor I_12316 (I215111,I214961,I215094);
and I_12317 (I215128,I214978,I215111);
and I_12318 (I215145,I215077,I215012);
DFFARX1 I_12319  ( .D(I215145), .CLK(I5694_clk), .RSTB(I214910_rst), .Q(I214878) );
DFFARX1 I_12320  ( .D(I215077), .CLK(I5694_clk), .RSTB(I214910_rst), .Q(I214872) );
DFFARX1 I_12321  ( .D(I169839), .CLK(I5694_clk), .RSTB(I214910_rst), .Q(I215190) );
and I_12322 (I215207,I215190,I169857);
nand I_12323 (I215224,I215207,I215077);
nor I_12324 (I214899,I215207,I214978);
not I_12325 (I215255,I215207);
nor I_12326 (I215272,I214961,I215255);
nand I_12327 (I214890,I214995,I215272);
nand I_12328 (I214884,I215077,I215255);
or I_12329 (I215317,I215207,I215128);
DFFARX1 I_12330  ( .D(I215317), .CLK(I5694_clk), .RSTB(I214910_rst), .Q(I214887) );
DFFARX1 I_12331  ( .D(I169863), .CLK(I5694_clk), .RSTB(I214910_rst), .Q(I215348) );
and I_12332 (I215365,I215348,I215224);
DFFARX1 I_12333  ( .D(I215365), .CLK(I5694_clk), .RSTB(I214910_rst), .Q(I214902) );
nor I_12334 (I215396,I215348,I214961);
nand I_12335 (I214896,I215207,I215396);
not I_12336 (I214893,I215348);
DFFARX1 I_12337  ( .D(I215348), .CLK(I5694_clk), .RSTB(I214910_rst), .Q(I215441) );
and I_12338 (I214875,I215348,I215441);
not I_12339 (I215505_rst,I5701);
nand I_12340 (I215522,I203647,I203662);
and I_12341 (I215539,I215522,I203659);
DFFARX1 I_12342  ( .D(I215539), .CLK(I5694_clk), .RSTB(I215505_rst), .Q(I215556) );
nor I_12343 (I215573,I203635,I203662);
DFFARX1 I_12344  ( .D(I203653), .CLK(I5694_clk), .RSTB(I215505_rst), .Q(I215590) );
nand I_12345 (I215607,I215590,I215573);
DFFARX1 I_12346  ( .D(I215590), .CLK(I5694_clk), .RSTB(I215505_rst), .Q(I215476) );
nand I_12347 (I215638,I203656,I203644);
and I_12348 (I215655,I215638,I203650);
DFFARX1 I_12349  ( .D(I215655), .CLK(I5694_clk), .RSTB(I215505_rst), .Q(I215672) );
not I_12350 (I215689,I215672);
nor I_12351 (I215706,I215556,I215689);
and I_12352 (I215723,I215573,I215706);
and I_12353 (I215740,I215672,I215607);
DFFARX1 I_12354  ( .D(I215740), .CLK(I5694_clk), .RSTB(I215505_rst), .Q(I215473) );
DFFARX1 I_12355  ( .D(I215672), .CLK(I5694_clk), .RSTB(I215505_rst), .Q(I215467) );
DFFARX1 I_12356  ( .D(I203641), .CLK(I5694_clk), .RSTB(I215505_rst), .Q(I215785) );
and I_12357 (I215802,I215785,I203665);
nand I_12358 (I215819,I215802,I215672);
nor I_12359 (I215494,I215802,I215573);
not I_12360 (I215850,I215802);
nor I_12361 (I215867,I215556,I215850);
nand I_12362 (I215485,I215590,I215867);
nand I_12363 (I215479,I215672,I215850);
or I_12364 (I215912,I215802,I215723);
DFFARX1 I_12365  ( .D(I215912), .CLK(I5694_clk), .RSTB(I215505_rst), .Q(I215482) );
DFFARX1 I_12366  ( .D(I203638), .CLK(I5694_clk), .RSTB(I215505_rst), .Q(I215943) );
and I_12367 (I215960,I215943,I215819);
DFFARX1 I_12368  ( .D(I215960), .CLK(I5694_clk), .RSTB(I215505_rst), .Q(I215497) );
nor I_12369 (I215991,I215943,I215556);
nand I_12370 (I215491,I215802,I215991);
not I_12371 (I215488,I215943);
DFFARX1 I_12372  ( .D(I215943), .CLK(I5694_clk), .RSTB(I215505_rst), .Q(I216036) );
and I_12373 (I215470,I215943,I216036);
not I_12374 (I216100_rst,I5701);
nand I_12375 (I216117,I191901,I191871);
and I_12376 (I216134,I216117,I191889);
DFFARX1 I_12377  ( .D(I216134), .CLK(I5694_clk), .RSTB(I216100_rst), .Q(I216151) );
nor I_12378 (I216168,I191883,I191871);
DFFARX1 I_12379  ( .D(I191880), .CLK(I5694_clk), .RSTB(I216100_rst), .Q(I216185) );
nand I_12380 (I216202,I216185,I216168);
DFFARX1 I_12381  ( .D(I216185), .CLK(I5694_clk), .RSTB(I216100_rst), .Q(I216071) );
nand I_12382 (I216233,I191874,I191877);
and I_12383 (I216250,I216233,I191895);
DFFARX1 I_12384  ( .D(I216250), .CLK(I5694_clk), .RSTB(I216100_rst), .Q(I216267) );
not I_12385 (I216284,I216267);
nor I_12386 (I216301,I216151,I216284);
and I_12387 (I216318,I216168,I216301);
and I_12388 (I216335,I216267,I216202);
DFFARX1 I_12389  ( .D(I216335), .CLK(I5694_clk), .RSTB(I216100_rst), .Q(I216068) );
DFFARX1 I_12390  ( .D(I216267), .CLK(I5694_clk), .RSTB(I216100_rst), .Q(I216062) );
DFFARX1 I_12391  ( .D(I191898), .CLK(I5694_clk), .RSTB(I216100_rst), .Q(I216380) );
and I_12392 (I216397,I216380,I191892);
nand I_12393 (I216414,I216397,I216267);
nor I_12394 (I216089,I216397,I216168);
not I_12395 (I216445,I216397);
nor I_12396 (I216462,I216151,I216445);
nand I_12397 (I216080,I216185,I216462);
nand I_12398 (I216074,I216267,I216445);
or I_12399 (I216507,I216397,I216318);
DFFARX1 I_12400  ( .D(I216507), .CLK(I5694_clk), .RSTB(I216100_rst), .Q(I216077) );
DFFARX1 I_12401  ( .D(I191886), .CLK(I5694_clk), .RSTB(I216100_rst), .Q(I216538) );
and I_12402 (I216555,I216538,I216414);
DFFARX1 I_12403  ( .D(I216555), .CLK(I5694_clk), .RSTB(I216100_rst), .Q(I216092) );
nor I_12404 (I216586,I216538,I216151);
nand I_12405 (I216086,I216397,I216586);
not I_12406 (I216083,I216538);
DFFARX1 I_12407  ( .D(I216538), .CLK(I5694_clk), .RSTB(I216100_rst), .Q(I216631) );
and I_12408 (I216065,I216538,I216631);
not I_12409 (I216695_rst,I5701);
nand I_12410 (I216712,I188586,I188556);
and I_12411 (I216729,I216712,I188574);
DFFARX1 I_12412  ( .D(I216729), .CLK(I5694_clk), .RSTB(I216695_rst), .Q(I216746) );
nor I_12413 (I216763,I188568,I188556);
DFFARX1 I_12414  ( .D(I188565), .CLK(I5694_clk), .RSTB(I216695_rst), .Q(I216780) );
nand I_12415 (I216797,I216780,I216763);
DFFARX1 I_12416  ( .D(I216780), .CLK(I5694_clk), .RSTB(I216695_rst), .Q(I216666) );
nand I_12417 (I216828,I188559,I188562);
and I_12418 (I216845,I216828,I188580);
DFFARX1 I_12419  ( .D(I216845), .CLK(I5694_clk), .RSTB(I216695_rst), .Q(I216862) );
not I_12420 (I216879,I216862);
nor I_12421 (I216896,I216746,I216879);
and I_12422 (I216913,I216763,I216896);
and I_12423 (I216930,I216862,I216797);
DFFARX1 I_12424  ( .D(I216930), .CLK(I5694_clk), .RSTB(I216695_rst), .Q(I216663) );
DFFARX1 I_12425  ( .D(I216862), .CLK(I5694_clk), .RSTB(I216695_rst), .Q(I216657) );
DFFARX1 I_12426  ( .D(I188583), .CLK(I5694_clk), .RSTB(I216695_rst), .Q(I216975) );
and I_12427 (I216992,I216975,I188577);
nand I_12428 (I217009,I216992,I216862);
nor I_12429 (I216684,I216992,I216763);
not I_12430 (I217040,I216992);
nor I_12431 (I217057,I216746,I217040);
nand I_12432 (I216675,I216780,I217057);
nand I_12433 (I216669,I216862,I217040);
or I_12434 (I217102,I216992,I216913);
DFFARX1 I_12435  ( .D(I217102), .CLK(I5694_clk), .RSTB(I216695_rst), .Q(I216672) );
DFFARX1 I_12436  ( .D(I188571), .CLK(I5694_clk), .RSTB(I216695_rst), .Q(I217133) );
and I_12437 (I217150,I217133,I217009);
DFFARX1 I_12438  ( .D(I217150), .CLK(I5694_clk), .RSTB(I216695_rst), .Q(I216687) );
nor I_12439 (I217181,I217133,I216746);
nand I_12440 (I216681,I216992,I217181);
not I_12441 (I216678,I217133);
DFFARX1 I_12442  ( .D(I217133), .CLK(I5694_clk), .RSTB(I216695_rst), .Q(I217226) );
and I_12443 (I216660,I217133,I217226);
not I_12444 (I217290_rst,I5701);
nand I_12445 (I217307,I185271,I185241);
and I_12446 (I217324,I217307,I185259);
DFFARX1 I_12447  ( .D(I217324), .CLK(I5694_clk), .RSTB(I217290_rst), .Q(I217341) );
nor I_12448 (I217358,I185253,I185241);
DFFARX1 I_12449  ( .D(I185250), .CLK(I5694_clk), .RSTB(I217290_rst), .Q(I217375) );
nand I_12450 (I217392,I217375,I217358);
DFFARX1 I_12451  ( .D(I217375), .CLK(I5694_clk), .RSTB(I217290_rst), .Q(I217261) );
nand I_12452 (I217423,I185244,I185247);
and I_12453 (I217440,I217423,I185265);
DFFARX1 I_12454  ( .D(I217440), .CLK(I5694_clk), .RSTB(I217290_rst), .Q(I217457) );
not I_12455 (I217474,I217457);
nor I_12456 (I217491,I217341,I217474);
and I_12457 (I217508,I217358,I217491);
and I_12458 (I217525,I217457,I217392);
DFFARX1 I_12459  ( .D(I217525), .CLK(I5694_clk), .RSTB(I217290_rst), .Q(I217258) );
DFFARX1 I_12460  ( .D(I217457), .CLK(I5694_clk), .RSTB(I217290_rst), .Q(I217252) );
DFFARX1 I_12461  ( .D(I185268), .CLK(I5694_clk), .RSTB(I217290_rst), .Q(I217570) );
and I_12462 (I217587,I217570,I185262);
nand I_12463 (I217604,I217587,I217457);
nor I_12464 (I217279,I217587,I217358);
not I_12465 (I217635,I217587);
nor I_12466 (I217652,I217341,I217635);
nand I_12467 (I217270,I217375,I217652);
nand I_12468 (I217264,I217457,I217635);
or I_12469 (I217697,I217587,I217508);
DFFARX1 I_12470  ( .D(I217697), .CLK(I5694_clk), .RSTB(I217290_rst), .Q(I217267) );
DFFARX1 I_12471  ( .D(I185256), .CLK(I5694_clk), .RSTB(I217290_rst), .Q(I217728) );
and I_12472 (I217745,I217728,I217604);
DFFARX1 I_12473  ( .D(I217745), .CLK(I5694_clk), .RSTB(I217290_rst), .Q(I217282) );
nor I_12474 (I217776,I217728,I217341);
nand I_12475 (I217276,I217587,I217776);
not I_12476 (I217273,I217728);
DFFARX1 I_12477  ( .D(I217728), .CLK(I5694_clk), .RSTB(I217290_rst), .Q(I217821) );
and I_12478 (I217255,I217728,I217821);
not I_12479 (I217885_rst,I5701);
not I_12480 (I217902,I176379);
nor I_12481 (I217919,I176370,I176394);
nand I_12482 (I217936,I217919,I176397);
nor I_12483 (I217953,I217902,I176370);
nand I_12484 (I217970,I217953,I176388);
not I_12485 (I217987,I176370);
not I_12486 (I218004,I217987);
not I_12487 (I218021,I176382);
nor I_12488 (I218038,I218021,I176376);
and I_12489 (I218055,I218038,I176385);
or I_12490 (I218072,I218055,I176373);
DFFARX1 I_12491  ( .D(I218072), .CLK(I5694_clk), .RSTB(I217885_rst), .Q(I218089) );
nand I_12492 (I218106,I217902,I176382);
or I_12493 (I217874,I218106,I218089);
not I_12494 (I218137,I218106);
nor I_12495 (I218154,I218089,I218137);
and I_12496 (I218171,I217987,I218154);
nand I_12497 (I217847,I218106,I218004);
DFFARX1 I_12498  ( .D(I176367), .CLK(I5694_clk), .RSTB(I217885_rst), .Q(I218202) );
or I_12499 (I217868,I218202,I218089);
nor I_12500 (I218233,I218202,I217970);
nor I_12501 (I218250,I218202,I218004);
nand I_12502 (I217853,I217936,I218250);
or I_12503 (I218281,I218202,I218171);
DFFARX1 I_12504  ( .D(I218281), .CLK(I5694_clk), .RSTB(I217885_rst), .Q(I217850) );
not I_12505 (I217856,I218202);
DFFARX1 I_12506  ( .D(I176391), .CLK(I5694_clk), .RSTB(I217885_rst), .Q(I218326) );
not I_12507 (I218343,I218326);
nor I_12508 (I218360,I218343,I217936);
DFFARX1 I_12509  ( .D(I218360), .CLK(I5694_clk), .RSTB(I217885_rst), .Q(I217862) );
nor I_12510 (I217877,I218202,I218343);
nor I_12511 (I217865,I218343,I218106);
not I_12512 (I218419,I218343);
and I_12513 (I218436,I217970,I218419);
nor I_12514 (I217871,I218106,I218436);
nand I_12515 (I217859,I218343,I218233);
not I_12516 (I218514_rst,I5701);
not I_12517 (I218531,I214881);
nor I_12518 (I218548,I214884,I214893);
nand I_12519 (I218565,I218548,I214878);
nor I_12520 (I218582,I218531,I214884);
nand I_12521 (I218599,I218582,I214887);
not I_12522 (I218616,I214884);
not I_12523 (I218633,I218616);
not I_12524 (I218650,I214902);
nor I_12525 (I218667,I218650,I214890);
and I_12526 (I218684,I218667,I214875);
or I_12527 (I218701,I218684,I214872);
DFFARX1 I_12528  ( .D(I218701), .CLK(I5694_clk), .RSTB(I218514_rst), .Q(I218718) );
nand I_12529 (I218735,I218531,I214902);
or I_12530 (I218503,I218735,I218718);
not I_12531 (I218766,I218735);
nor I_12532 (I218783,I218718,I218766);
and I_12533 (I218800,I218616,I218783);
nand I_12534 (I218476,I218735,I218633);
DFFARX1 I_12535  ( .D(I214896), .CLK(I5694_clk), .RSTB(I218514_rst), .Q(I218831) );
or I_12536 (I218497,I218831,I218718);
nor I_12537 (I218862,I218831,I218599);
nor I_12538 (I218879,I218831,I218633);
nand I_12539 (I218482,I218565,I218879);
or I_12540 (I218910,I218831,I218800);
DFFARX1 I_12541  ( .D(I218910), .CLK(I5694_clk), .RSTB(I218514_rst), .Q(I218479) );
not I_12542 (I218485,I218831);
DFFARX1 I_12543  ( .D(I214899), .CLK(I5694_clk), .RSTB(I218514_rst), .Q(I218955) );
not I_12544 (I218972,I218955);
nor I_12545 (I218989,I218972,I218565);
DFFARX1 I_12546  ( .D(I218989), .CLK(I5694_clk), .RSTB(I218514_rst), .Q(I218491) );
nor I_12547 (I218506,I218831,I218972);
nor I_12548 (I218494,I218972,I218735);
not I_12549 (I219048,I218972);
and I_12550 (I219065,I218599,I219048);
nor I_12551 (I218500,I218735,I219065);
nand I_12552 (I218488,I218972,I218862);
not I_12553 (I219143_rst,I5701);
not I_12554 (I219160,I200197);
nor I_12555 (I219177,I200170,I200188);
nand I_12556 (I219194,I219177,I200173);
nor I_12557 (I219211,I219160,I200170);
nand I_12558 (I219228,I219211,I200191);
not I_12559 (I219245,I200170);
not I_12560 (I219262,I219245);
not I_12561 (I219279,I200167);
nor I_12562 (I219296,I219279,I200194);
and I_12563 (I219313,I219296,I200185);
or I_12564 (I219330,I219313,I200176);
DFFARX1 I_12565  ( .D(I219330), .CLK(I5694_clk), .RSTB(I219143_rst), .Q(I219347) );
nand I_12566 (I219364,I219160,I200167);
or I_12567 (I219132,I219364,I219347);
not I_12568 (I219395,I219364);
nor I_12569 (I219412,I219347,I219395);
and I_12570 (I219429,I219245,I219412);
nand I_12571 (I219105,I219364,I219262);
DFFARX1 I_12572  ( .D(I200179), .CLK(I5694_clk), .RSTB(I219143_rst), .Q(I219460) );
or I_12573 (I219126,I219460,I219347);
nor I_12574 (I219491,I219460,I219228);
nor I_12575 (I219508,I219460,I219262);
nand I_12576 (I219111,I219194,I219508);
or I_12577 (I219539,I219460,I219429);
DFFARX1 I_12578  ( .D(I219539), .CLK(I5694_clk), .RSTB(I219143_rst), .Q(I219108) );
not I_12579 (I219114,I219460);
DFFARX1 I_12580  ( .D(I200182), .CLK(I5694_clk), .RSTB(I219143_rst), .Q(I219584) );
not I_12581 (I219601,I219584);
nor I_12582 (I219618,I219601,I219194);
DFFARX1 I_12583  ( .D(I219618), .CLK(I5694_clk), .RSTB(I219143_rst), .Q(I219120) );
nor I_12584 (I219135,I219460,I219601);
nor I_12585 (I219123,I219601,I219364);
not I_12586 (I219677,I219601);
and I_12587 (I219694,I219228,I219677);
nor I_12588 (I219129,I219364,I219694);
nand I_12589 (I219117,I219601,I219491);
not I_12590 (I219772_rst,I5701);
not I_12591 (I219789,I186585);
nor I_12592 (I219806,I186591,I186570);
nand I_12593 (I219823,I219806,I186576);
nor I_12594 (I219840,I219789,I186591);
nand I_12595 (I219857,I219840,I186582);
not I_12596 (I219874,I186591);
not I_12597 (I219891,I219874);
not I_12598 (I219908,I186579);
nor I_12599 (I219925,I219908,I186597);
and I_12600 (I219942,I219925,I186588);
or I_12601 (I219959,I219942,I186567);
DFFARX1 I_12602  ( .D(I219959), .CLK(I5694_clk), .RSTB(I219772_rst), .Q(I219976) );
nand I_12603 (I219993,I219789,I186579);
or I_12604 (I219761,I219993,I219976);
not I_12605 (I220024,I219993);
nor I_12606 (I220041,I219976,I220024);
and I_12607 (I220058,I219874,I220041);
nand I_12608 (I219734,I219993,I219891);
DFFARX1 I_12609  ( .D(I186594), .CLK(I5694_clk), .RSTB(I219772_rst), .Q(I220089) );
or I_12610 (I219755,I220089,I219976);
nor I_12611 (I220120,I220089,I219857);
nor I_12612 (I220137,I220089,I219891);
nand I_12613 (I219740,I219823,I220137);
or I_12614 (I220168,I220089,I220058);
DFFARX1 I_12615  ( .D(I220168), .CLK(I5694_clk), .RSTB(I219772_rst), .Q(I219737) );
not I_12616 (I219743,I220089);
DFFARX1 I_12617  ( .D(I186573), .CLK(I5694_clk), .RSTB(I219772_rst), .Q(I220213) );
not I_12618 (I220230,I220213);
nor I_12619 (I220247,I220230,I219823);
DFFARX1 I_12620  ( .D(I220247), .CLK(I5694_clk), .RSTB(I219772_rst), .Q(I219749) );
nor I_12621 (I219764,I220089,I220230);
nor I_12622 (I219752,I220230,I219993);
not I_12623 (I220306,I220230);
and I_12624 (I220323,I219857,I220306);
nor I_12625 (I219758,I219993,I220323);
nand I_12626 (I219746,I220230,I220120);
not I_12627 (I220401_rst,I5701);
not I_12628 (I220418,I204821);
nor I_12629 (I220435,I204794,I204812);
nand I_12630 (I220452,I220435,I204797);
nor I_12631 (I220469,I220418,I204794);
nand I_12632 (I220486,I220469,I204815);
not I_12633 (I220503,I204794);
not I_12634 (I220520,I220503);
not I_12635 (I220537,I204791);
nor I_12636 (I220554,I220537,I204818);
and I_12637 (I220571,I220554,I204809);
or I_12638 (I220588,I220571,I204800);
DFFARX1 I_12639  ( .D(I220588), .CLK(I5694_clk), .RSTB(I220401_rst), .Q(I220605) );
nand I_12640 (I220622,I220418,I204791);
or I_12641 (I220390,I220622,I220605);
not I_12642 (I220653,I220622);
nor I_12643 (I220670,I220605,I220653);
and I_12644 (I220687,I220503,I220670);
nand I_12645 (I220363,I220622,I220520);
DFFARX1 I_12646  ( .D(I204803), .CLK(I5694_clk), .RSTB(I220401_rst), .Q(I220718) );
or I_12647 (I220384,I220718,I220605);
nor I_12648 (I220749,I220718,I220486);
nor I_12649 (I220766,I220718,I220520);
nand I_12650 (I220369,I220452,I220766);
or I_12651 (I220797,I220718,I220687);
DFFARX1 I_12652  ( .D(I220797), .CLK(I5694_clk), .RSTB(I220401_rst), .Q(I220366) );
not I_12653 (I220372,I220718);
DFFARX1 I_12654  ( .D(I204806), .CLK(I5694_clk), .RSTB(I220401_rst), .Q(I220842) );
not I_12655 (I220859,I220842);
nor I_12656 (I220876,I220859,I220452);
DFFARX1 I_12657  ( .D(I220876), .CLK(I5694_clk), .RSTB(I220401_rst), .Q(I220378) );
nor I_12658 (I220393,I220718,I220859);
nor I_12659 (I220381,I220859,I220622);
not I_12660 (I220935,I220859);
and I_12661 (I220952,I220486,I220935);
nor I_12662 (I220387,I220622,I220952);
nand I_12663 (I220375,I220859,I220749);
not I_12664 (I221030_rst,I5701);
not I_12665 (I221047,I209523);
nor I_12666 (I221064,I209541,I209520);
nand I_12667 (I221081,I221064,I209544);
nor I_12668 (I221098,I221047,I209541);
nand I_12669 (I221115,I221098,I209538);
not I_12670 (I221132,I209541);
not I_12671 (I221149,I221132);
not I_12672 (I221166,I209529);
nor I_12673 (I221183,I221166,I209517);
and I_12674 (I221200,I221183,I209535);
or I_12675 (I221217,I221200,I209547);
DFFARX1 I_12676  ( .D(I221217), .CLK(I5694_clk), .RSTB(I221030_rst), .Q(I221234) );
nand I_12677 (I221251,I221047,I209529);
or I_12678 (I221019,I221251,I221234);
not I_12679 (I221282,I221251);
nor I_12680 (I221299,I221234,I221282);
and I_12681 (I221316,I221132,I221299);
nand I_12682 (I220992,I221251,I221149);
DFFARX1 I_12683  ( .D(I209526), .CLK(I5694_clk), .RSTB(I221030_rst), .Q(I221347) );
or I_12684 (I221013,I221347,I221234);
nor I_12685 (I221378,I221347,I221115);
nor I_12686 (I221395,I221347,I221149);
nand I_12687 (I220998,I221081,I221395);
or I_12688 (I221426,I221347,I221316);
DFFARX1 I_12689  ( .D(I221426), .CLK(I5694_clk), .RSTB(I221030_rst), .Q(I220995) );
not I_12690 (I221001,I221347);
DFFARX1 I_12691  ( .D(I209532), .CLK(I5694_clk), .RSTB(I221030_rst), .Q(I221471) );
not I_12692 (I221488,I221471);
nor I_12693 (I221505,I221488,I221081);
DFFARX1 I_12694  ( .D(I221505), .CLK(I5694_clk), .RSTB(I221030_rst), .Q(I221007) );
nor I_12695 (I221022,I221347,I221488);
nor I_12696 (I221010,I221488,I221251);
not I_12697 (I221564,I221488);
and I_12698 (I221581,I221115,I221564);
nor I_12699 (I221016,I221251,I221581);
nand I_12700 (I221004,I221488,I221378);
not I_12701 (I221659_rst,I5701);
nand I_12702 (I221676,I208339,I208357);
and I_12703 (I221693,I221676,I208333);
DFFARX1 I_12704  ( .D(I221693), .CLK(I5694_clk), .RSTB(I221659_rst), .Q(I221710) );
not I_12705 (I221648,I221710);
DFFARX1 I_12706  ( .D(I221710), .CLK(I5694_clk), .RSTB(I221659_rst), .Q(I221741) );
not I_12707 (I221636,I221741);
nor I_12708 (I221772,I208345,I208357);
not I_12709 (I221789,I221772);
nor I_12710 (I221806,I221710,I221789);
DFFARX1 I_12711  ( .D(I208336), .CLK(I5694_clk), .RSTB(I221659_rst), .Q(I221823) );
not I_12712 (I221840,I221823);
nand I_12713 (I221639,I221823,I221789);
DFFARX1 I_12714  ( .D(I221823), .CLK(I5694_clk), .RSTB(I221659_rst), .Q(I221871) );
and I_12715 (I221624,I221710,I221871);
nand I_12716 (I221902,I208351,I208330);
and I_12717 (I221919,I221902,I208348);
DFFARX1 I_12718  ( .D(I221919), .CLK(I5694_clk), .RSTB(I221659_rst), .Q(I221936) );
nor I_12719 (I221953,I221936,I221840);
and I_12720 (I221970,I221772,I221953);
nor I_12721 (I221987,I221936,I221710);
DFFARX1 I_12722  ( .D(I221936), .CLK(I5694_clk), .RSTB(I221659_rst), .Q(I221630) );
DFFARX1 I_12723  ( .D(I208354), .CLK(I5694_clk), .RSTB(I221659_rst), .Q(I222018) );
and I_12724 (I222035,I222018,I208342);
or I_12725 (I222052,I222035,I221970);
DFFARX1 I_12726  ( .D(I222052), .CLK(I5694_clk), .RSTB(I221659_rst), .Q(I221642) );
nand I_12727 (I221651,I222035,I221987);
DFFARX1 I_12728  ( .D(I222035), .CLK(I5694_clk), .RSTB(I221659_rst), .Q(I221621) );
DFFARX1 I_12729  ( .D(I208327), .CLK(I5694_clk), .RSTB(I221659_rst), .Q(I222111) );
nand I_12730 (I221645,I222111,I221806);
DFFARX1 I_12731  ( .D(I222111), .CLK(I5694_clk), .RSTB(I221659_rst), .Q(I221633) );
nand I_12732 (I222156,I222111,I221772);
and I_12733 (I222173,I221823,I222156);
DFFARX1 I_12734  ( .D(I222173), .CLK(I5694_clk), .RSTB(I221659_rst), .Q(I221627) );
not I_12735 (I222237_rst,I5701);
nand I_12736 (I222254,I193215,I193218);
and I_12737 (I222271,I222254,I193197);
DFFARX1 I_12738  ( .D(I222271), .CLK(I5694_clk), .RSTB(I222237_rst), .Q(I222288) );
not I_12739 (I222226,I222288);
DFFARX1 I_12740  ( .D(I222288), .CLK(I5694_clk), .RSTB(I222237_rst), .Q(I222319) );
not I_12741 (I222214,I222319);
nor I_12742 (I222350,I193212,I193218);
not I_12743 (I222367,I222350);
nor I_12744 (I222384,I222288,I222367);
DFFARX1 I_12745  ( .D(I193221), .CLK(I5694_clk), .RSTB(I222237_rst), .Q(I222401) );
not I_12746 (I222418,I222401);
nand I_12747 (I222217,I222401,I222367);
DFFARX1 I_12748  ( .D(I222401), .CLK(I5694_clk), .RSTB(I222237_rst), .Q(I222449) );
and I_12749 (I222202,I222288,I222449);
nand I_12750 (I222480,I193209,I193227);
and I_12751 (I222497,I222480,I193203);
DFFARX1 I_12752  ( .D(I222497), .CLK(I5694_clk), .RSTB(I222237_rst), .Q(I222514) );
nor I_12753 (I222531,I222514,I222418);
and I_12754 (I222548,I222350,I222531);
nor I_12755 (I222565,I222514,I222288);
DFFARX1 I_12756  ( .D(I222514), .CLK(I5694_clk), .RSTB(I222237_rst), .Q(I222208) );
DFFARX1 I_12757  ( .D(I193200), .CLK(I5694_clk), .RSTB(I222237_rst), .Q(I222596) );
and I_12758 (I222613,I222596,I193206);
or I_12759 (I222630,I222613,I222548);
DFFARX1 I_12760  ( .D(I222630), .CLK(I5694_clk), .RSTB(I222237_rst), .Q(I222220) );
nand I_12761 (I222229,I222613,I222565);
DFFARX1 I_12762  ( .D(I222613), .CLK(I5694_clk), .RSTB(I222237_rst), .Q(I222199) );
DFFARX1 I_12763  ( .D(I193224), .CLK(I5694_clk), .RSTB(I222237_rst), .Q(I222689) );
nand I_12764 (I222223,I222689,I222384);
DFFARX1 I_12765  ( .D(I222689), .CLK(I5694_clk), .RSTB(I222237_rst), .Q(I222211) );
nand I_12766 (I222734,I222689,I222350);
and I_12767 (I222751,I222401,I222734);
DFFARX1 I_12768  ( .D(I222751), .CLK(I5694_clk), .RSTB(I222237_rst), .Q(I222205) );
not I_12769 (I222815_rst,I5701);
nand I_12770 (I222832,I201904,I201922);
and I_12771 (I222849,I222832,I201913);
DFFARX1 I_12772  ( .D(I222849), .CLK(I5694_clk), .RSTB(I222815_rst), .Q(I222866) );
not I_12773 (I222804,I222866);
DFFARX1 I_12774  ( .D(I222866), .CLK(I5694_clk), .RSTB(I222815_rst), .Q(I222897) );
not I_12775 (I222792,I222897);
nor I_12776 (I222928,I201910,I201922);
not I_12777 (I222945,I222928);
nor I_12778 (I222962,I222866,I222945);
DFFARX1 I_12779  ( .D(I201901), .CLK(I5694_clk), .RSTB(I222815_rst), .Q(I222979) );
not I_12780 (I222996,I222979);
nand I_12781 (I222795,I222979,I222945);
DFFARX1 I_12782  ( .D(I222979), .CLK(I5694_clk), .RSTB(I222815_rst), .Q(I223027) );
and I_12783 (I222780,I222866,I223027);
nand I_12784 (I223058,I201919,I201931);
and I_12785 (I223075,I223058,I201925);
DFFARX1 I_12786  ( .D(I223075), .CLK(I5694_clk), .RSTB(I222815_rst), .Q(I223092) );
nor I_12787 (I223109,I223092,I222996);
and I_12788 (I223126,I222928,I223109);
nor I_12789 (I223143,I223092,I222866);
DFFARX1 I_12790  ( .D(I223092), .CLK(I5694_clk), .RSTB(I222815_rst), .Q(I222786) );
DFFARX1 I_12791  ( .D(I201907), .CLK(I5694_clk), .RSTB(I222815_rst), .Q(I223174) );
and I_12792 (I223191,I223174,I201916);
or I_12793 (I223208,I223191,I223126);
DFFARX1 I_12794  ( .D(I223208), .CLK(I5694_clk), .RSTB(I222815_rst), .Q(I222798) );
nand I_12795 (I222807,I223191,I223143);
DFFARX1 I_12796  ( .D(I223191), .CLK(I5694_clk), .RSTB(I222815_rst), .Q(I222777) );
DFFARX1 I_12797  ( .D(I201928), .CLK(I5694_clk), .RSTB(I222815_rst), .Q(I223267) );
nand I_12798 (I222801,I223267,I222962);
DFFARX1 I_12799  ( .D(I223267), .CLK(I5694_clk), .RSTB(I222815_rst), .Q(I222789) );
nand I_12800 (I223312,I223267,I222928);
and I_12801 (I223329,I222979,I223312);
DFFARX1 I_12802  ( .D(I223329), .CLK(I5694_clk), .RSTB(I222815_rst), .Q(I222783) );
not I_12803 (I223393_rst,I5701);
nand I_12804 (I223410,I178356,I178386);
and I_12805 (I223427,I223410,I178368);
DFFARX1 I_12806  ( .D(I223427), .CLK(I5694_clk), .RSTB(I223393_rst), .Q(I223444) );
not I_12807 (I223382,I223444);
DFFARX1 I_12808  ( .D(I223444), .CLK(I5694_clk), .RSTB(I223393_rst), .Q(I223475) );
not I_12809 (I223370,I223475);
nor I_12810 (I223506,I178365,I178386);
not I_12811 (I223523,I223506);
nor I_12812 (I223540,I223444,I223523);
DFFARX1 I_12813  ( .D(I178359), .CLK(I5694_clk), .RSTB(I223393_rst), .Q(I223557) );
not I_12814 (I223574,I223557);
nand I_12815 (I223373,I223557,I223523);
DFFARX1 I_12816  ( .D(I223557), .CLK(I5694_clk), .RSTB(I223393_rst), .Q(I223605) );
and I_12817 (I223358,I223444,I223605);
nand I_12818 (I223636,I178362,I178377);
and I_12819 (I223653,I223636,I178374);
DFFARX1 I_12820  ( .D(I223653), .CLK(I5694_clk), .RSTB(I223393_rst), .Q(I223670) );
nor I_12821 (I223687,I223670,I223574);
and I_12822 (I223704,I223506,I223687);
nor I_12823 (I223721,I223670,I223444);
DFFARX1 I_12824  ( .D(I223670), .CLK(I5694_clk), .RSTB(I223393_rst), .Q(I223364) );
DFFARX1 I_12825  ( .D(I178371), .CLK(I5694_clk), .RSTB(I223393_rst), .Q(I223752) );
and I_12826 (I223769,I223752,I178383);
or I_12827 (I223786,I223769,I223704);
DFFARX1 I_12828  ( .D(I223786), .CLK(I5694_clk), .RSTB(I223393_rst), .Q(I223376) );
nand I_12829 (I223385,I223769,I223721);
DFFARX1 I_12830  ( .D(I223769), .CLK(I5694_clk), .RSTB(I223393_rst), .Q(I223355) );
DFFARX1 I_12831  ( .D(I178380), .CLK(I5694_clk), .RSTB(I223393_rst), .Q(I223845) );
nand I_12832 (I223379,I223845,I223540);
DFFARX1 I_12833  ( .D(I223845), .CLK(I5694_clk), .RSTB(I223393_rst), .Q(I223367) );
nand I_12834 (I223890,I223845,I223506);
and I_12835 (I223907,I223557,I223890);
DFFARX1 I_12836  ( .D(I223907), .CLK(I5694_clk), .RSTB(I223393_rst), .Q(I223361) );
not I_12837 (I223971_rst,I5701);
nand I_12838 (I223988,I183924,I183921);
and I_12839 (I224005,I223988,I183945);
DFFARX1 I_12840  ( .D(I224005), .CLK(I5694_clk), .RSTB(I223971_rst), .Q(I224022) );
not I_12841 (I223960,I224022);
DFFARX1 I_12842  ( .D(I224022), .CLK(I5694_clk), .RSTB(I223971_rst), .Q(I224053) );
not I_12843 (I223948,I224053);
nor I_12844 (I224084,I183927,I183921);
not I_12845 (I224101,I224084);
nor I_12846 (I224118,I224022,I224101);
DFFARX1 I_12847  ( .D(I183942), .CLK(I5694_clk), .RSTB(I223971_rst), .Q(I224135) );
not I_12848 (I224152,I224135);
nand I_12849 (I223951,I224135,I224101);
DFFARX1 I_12850  ( .D(I224135), .CLK(I5694_clk), .RSTB(I223971_rst), .Q(I224183) );
and I_12851 (I223936,I224022,I224183);
nand I_12852 (I224214,I183930,I183915);
and I_12853 (I224231,I224214,I183933);
DFFARX1 I_12854  ( .D(I224231), .CLK(I5694_clk), .RSTB(I223971_rst), .Q(I224248) );
nor I_12855 (I224265,I224248,I224152);
and I_12856 (I224282,I224084,I224265);
nor I_12857 (I224299,I224248,I224022);
DFFARX1 I_12858  ( .D(I224248), .CLK(I5694_clk), .RSTB(I223971_rst), .Q(I223942) );
DFFARX1 I_12859  ( .D(I183936), .CLK(I5694_clk), .RSTB(I223971_rst), .Q(I224330) );
and I_12860 (I224347,I224330,I183939);
or I_12861 (I22436_rst4,I224347,I224282);
DFFARX1 I_12862  ( .D(I22436_rst4), .CLK(I5694_clk), .RSTB(I223971_rst), .Q(I223954) );
nand I_12863 (I223963,I224347,I224299);
DFFARX1 I_12864  ( .D(I224347), .CLK(I5694_clk), .RSTB(I223971_rst), .Q(I223933) );
DFFARX1 I_12865  ( .D(I183918), .CLK(I5694_clk), .RSTB(I223971_rst), .Q(I224423) );
nand I_12866 (I223957,I224423,I224118);
DFFARX1 I_12867  ( .D(I224423), .CLK(I5694_clk), .RSTB(I223971_rst), .Q(I223945) );
nand I_12868 (I224468,I224423,I224084);
and I_12869 (I224485,I224135,I224468);
DFFARX1 I_12870  ( .D(I224485), .CLK(I5694_clk), .RSTB(I223971_rst), .Q(I223939) );
not I_12871 (I224549_rst,I5701);
nand I_12872 (I224566,I168568,I168553);
and I_12873 (I224583,I224566,I168547);
DFFARX1 I_12874  ( .D(I224583), .CLK(I5694_clk), .RSTB(I224549_rst), .Q(I224600) );
not I_12875 (I224538,I224600);
DFFARX1 I_12876  ( .D(I224600), .CLK(I5694_clk), .RSTB(I224549_rst), .Q(I224631) );
not I_12877 (I224526,I224631);
nor I_12878 (I224662,I168574,I168553);
not I_12879 (I224679,I224662);
nor I_12880 (I224696,I224600,I224679);
DFFARX1 I_12881  ( .D(I168577), .CLK(I5694_clk), .RSTB(I224549_rst), .Q(I224713) );
not I_12882 (I224730,I224713);
nand I_12883 (I224529,I224713,I224679);
DFFARX1 I_12884  ( .D(I224713), .CLK(I5694_clk), .RSTB(I224549_rst), .Q(I224761) );
and I_12885 (I224514,I224600,I224761);
nand I_12886 (I224792,I168559,I168562);
and I_12887 (I224809,I224792,I168565);
DFFARX1 I_12888  ( .D(I224809), .CLK(I5694_clk), .RSTB(I224549_rst), .Q(I224826) );
nor I_12889 (I224843,I224826,I224730);
and I_12890 (I224860,I224662,I224843);
nor I_12891 (I224877,I224826,I224600);
DFFARX1 I_12892  ( .D(I224826), .CLK(I5694_clk), .RSTB(I224549_rst), .Q(I224520) );
DFFARX1 I_12893  ( .D(I168571), .CLK(I5694_clk), .RSTB(I224549_rst), .Q(I224908) );
and I_12894 (I224925,I224908,I168556);
or I_12895 (I224942,I224925,I224860);
DFFARX1 I_12896  ( .D(I224942), .CLK(I5694_clk), .RSTB(I224549_rst), .Q(I224532) );
nand I_12897 (I224541,I224925,I224877);
DFFARX1 I_12898  ( .D(I224925), .CLK(I5694_clk), .RSTB(I224549_rst), .Q(I224511) );
DFFARX1 I_12899  ( .D(I168550), .CLK(I5694_clk), .RSTB(I224549_rst), .Q(I225001) );
nand I_12900 (I224535,I225001,I224696);
DFFARX1 I_12901  ( .D(I225001), .CLK(I5694_clk), .RSTB(I224549_rst), .Q(I224523) );
nand I_12902 (I225046,I225001,I224662);
and I_12903 (I225063,I224713,I225046);
DFFARX1 I_12904  ( .D(I225063), .CLK(I5694_clk), .RSTB(I224549_rst), .Q(I224517) );
not I_12905 (I225127_rst,I5701);
nand I_12906 (I225144,I213108,I213090);
and I_12907 (I225161,I225144,I213105);
DFFARX1 I_12908  ( .D(I225161), .CLK(I5694_clk), .RSTB(I225127_rst), .Q(I225178) );
not I_12909 (I225116,I225178);
DFFARX1 I_12910  ( .D(I225178), .CLK(I5694_clk), .RSTB(I225127_rst), .Q(I225209) );
not I_12911 (I225104,I225209);
nor I_12912 (I225240,I213096,I213090);
not I_12913 (I225257,I225240);
nor I_12914 (I225274,I225178,I225257);
DFFARX1 I_12915  ( .D(I213111), .CLK(I5694_clk), .RSTB(I225127_rst), .Q(I225291) );
not I_12916 (I225308,I225291);
nand I_12917 (I225107,I225291,I225257);
DFFARX1 I_12918  ( .D(I225291), .CLK(I5694_clk), .RSTB(I225127_rst), .Q(I225339) );
and I_12919 (I225092,I225178,I225339);
nand I_12920 (I225370,I213087,I213093);
and I_12921 (I225387,I225370,I213099);
DFFARX1 I_12922  ( .D(I225387), .CLK(I5694_clk), .RSTB(I225127_rst), .Q(I225404) );
nor I_12923 (I225421,I225404,I225308);
and I_12924 (I225438,I225240,I225421);
nor I_12925 (I225455,I225404,I225178);
DFFARX1 I_12926  ( .D(I225404), .CLK(I5694_clk), .RSTB(I225127_rst), .Q(I225098) );
DFFARX1 I_12927  ( .D(I213114), .CLK(I5694_clk), .RSTB(I225127_rst), .Q(I225486) );
and I_12928 (I225503,I225486,I213102);
or I_12929 (I225520,I225503,I225438);
DFFARX1 I_12930  ( .D(I225520), .CLK(I5694_clk), .RSTB(I225127_rst), .Q(I225110) );
nand I_12931 (I225119,I225503,I225455);
DFFARX1 I_12932  ( .D(I225503), .CLK(I5694_clk), .RSTB(I225127_rst), .Q(I225089) );
DFFARX1 I_12933  ( .D(I213117), .CLK(I5694_clk), .RSTB(I225127_rst), .Q(I225579) );
nand I_12934 (I225113,I225579,I225274);
DFFARX1 I_12935  ( .D(I225579), .CLK(I5694_clk), .RSTB(I225127_rst), .Q(I225101) );
nand I_12936 (I225624,I225579,I225240);
and I_12937 (I225641,I225291,I225624);
DFFARX1 I_12938  ( .D(I225641), .CLK(I5694_clk), .RSTB(I225127_rst), .Q(I225095) );
not I_12939 (I225705_rst,I5701);
nand I_12940 (I225722,I206528,I206546);
and I_12941 (I225739,I225722,I206537);
DFFARX1 I_12942  ( .D(I225739), .CLK(I5694_clk), .RSTB(I225705_rst), .Q(I225756) );
not I_12943 (I225694,I225756);
DFFARX1 I_12944  ( .D(I225756), .CLK(I5694_clk), .RSTB(I225705_rst), .Q(I225787) );
not I_12945 (I225682,I225787);
nor I_12946 (I225818,I206534,I206546);
not I_12947 (I225835,I225818);
nor I_12948 (I225852,I225756,I225835);
DFFARX1 I_12949  ( .D(I206525), .CLK(I5694_clk), .RSTB(I225705_rst), .Q(I225869) );
not I_12950 (I225886,I225869);
nand I_12951 (I225685,I225869,I225835);
DFFARX1 I_12952  ( .D(I225869), .CLK(I5694_clk), .RSTB(I225705_rst), .Q(I225917) );
and I_12953 (I225670,I225756,I225917);
nand I_12954 (I225948,I206543,I206555);
and I_12955 (I225965,I225948,I206549);
DFFARX1 I_12956  ( .D(I225965), .CLK(I5694_clk), .RSTB(I225705_rst), .Q(I225982) );
nor I_12957 (I225999,I225982,I225886);
and I_12958 (I226016,I225818,I225999);
nor I_12959 (I226033,I225982,I225756);
DFFARX1 I_12960  ( .D(I225982), .CLK(I5694_clk), .RSTB(I225705_rst), .Q(I225676) );
DFFARX1 I_12961  ( .D(I206531), .CLK(I5694_clk), .RSTB(I225705_rst), .Q(I226064) );
and I_12962 (I226081,I226064,I206540);
or I_12963 (I226098,I226081,I226016);
DFFARX1 I_12964  ( .D(I226098), .CLK(I5694_clk), .RSTB(I225705_rst), .Q(I225688) );
nand I_12965 (I225697,I226081,I226033);
DFFARX1 I_12966  ( .D(I226081), .CLK(I5694_clk), .RSTB(I225705_rst), .Q(I225667) );
DFFARX1 I_12967  ( .D(I206552), .CLK(I5694_clk), .RSTB(I225705_rst), .Q(I226157) );
nand I_12968 (I225691,I226157,I225852);
DFFARX1 I_12969  ( .D(I226157), .CLK(I5694_clk), .RSTB(I225705_rst), .Q(I225679) );
nand I_12970 (I226202,I226157,I225818);
and I_12971 (I226219,I225869,I226202);
DFFARX1 I_12972  ( .D(I226219), .CLK(I5694_clk), .RSTB(I225705_rst), .Q(I225673) );
not I_12973 (I226283_rst,I5701);
nand I_12974 (I226300,I205959,I205956);
and I_12975 (I226317,I226300,I205950);
DFFARX1 I_12976  ( .D(I226317), .CLK(I5694_clk), .RSTB(I226283_rst), .Q(I226334) );
not I_12977 (I226351,I226334);
nor I_12978 (I226368,I205962,I205956);
or I_12979 (I226266,I226368,I226334);
not I_12980 (I226254,I226368);
DFFARX1 I_12981  ( .D(I205974), .CLK(I5694_clk), .RSTB(I226283_rst), .Q(I226413) );
nor I_12982 (I226430,I226413,I226368);
nand I_12983 (I226447,I205965,I205947);
and I_12984 (I226464,I226447,I205977);
DFFARX1 I_12985  ( .D(I226464), .CLK(I5694_clk), .RSTB(I226283_rst), .Q(I226481) );
nor I_12986 (I226263,I226481,I226334);
not I_12987 (I226512,I226481);
nor I_12988 (I226529,I226413,I226512);
DFFARX1 I_12989  ( .D(I205953), .CLK(I5694_clk), .RSTB(I226283_rst), .Q(I226546) );
and I_12990 (I226563,I226546,I205971);
or I_12991 (I226272,I226563,I226368);
nand I_12992 (I226251,I226563,I226529);
DFFARX1 I_12993  ( .D(I205968), .CLK(I5694_clk), .RSTB(I226283_rst), .Q(I226608) );
and I_12994 (I226625,I226608,I226351);
nor I_12995 (I226269,I226563,I226625);
nor I_12996 (I226656,I226608,I226413);
DFFARX1 I_12997  ( .D(I226656), .CLK(I5694_clk), .RSTB(I226283_rst), .Q(I226260) );
nor I_12998 (I226275,I226608,I226334);
not I_12999 (I226701,I226608);
nor I_13000 (I226718,I226481,I226701);
and I_13001 (I226735,I226368,I226718);
or I_13002 (I226752,I226563,I226735);
DFFARX1 I_13003  ( .D(I226752), .CLK(I5694_clk), .RSTB(I226283_rst), .Q(I226248) );
nand I_13004 (I226257,I226608,I226430);
nand I_13005 (I226245,I226608,I226512);
not I_13006 (I226844_rst,I5701);
nand I_13007 (I226861,I210115,I210118);
and I_13008 (I226878,I226861,I210130);
DFFARX1 I_13009  ( .D(I226878), .CLK(I5694_clk), .RSTB(I226844_rst), .Q(I226895) );
not I_13010 (I226912,I226895);
nor I_13011 (I226929,I210124,I210118);
or I_13012 (I226827,I226929,I226895);
not I_13013 (I226815,I226929);
DFFARX1 I_13014  ( .D(I210127), .CLK(I5694_clk), .RSTB(I226844_rst), .Q(I226974) );
nor I_13015 (I226991,I226974,I226929);
nand I_13016 (I227008,I210121,I210139);
and I_13017 (I227025,I227008,I210142);
DFFARX1 I_13018  ( .D(I227025), .CLK(I5694_clk), .RSTB(I226844_rst), .Q(I227042) );
nor I_13019 (I226824,I227042,I226895);
not I_13020 (I227073,I227042);
nor I_13021 (I227090,I226974,I227073);
DFFARX1 I_13022  ( .D(I210112), .CLK(I5694_clk), .RSTB(I226844_rst), .Q(I227107) );
and I_13023 (I227124,I227107,I210133);
or I_13024 (I226833,I227124,I226929);
nand I_13025 (I226812,I227124,I227090);
DFFARX1 I_13026  ( .D(I210136), .CLK(I5694_clk), .RSTB(I226844_rst), .Q(I227169) );
and I_13027 (I227186,I227169,I226912);
nor I_13028 (I226830,I227124,I227186);
nor I_13029 (I227217,I227169,I226974);
DFFARX1 I_13030  ( .D(I227217), .CLK(I5694_clk), .RSTB(I226844_rst), .Q(I226821) );
nor I_13031 (I226836,I227169,I226895);
not I_13032 (I227262,I227169);
nor I_13033 (I227279,I227042,I227262);
and I_13034 (I227296,I226929,I227279);
or I_13035 (I227313,I227124,I227296);
DFFARX1 I_13036  ( .D(I227313), .CLK(I5694_clk), .RSTB(I226844_rst), .Q(I226809) );
nand I_13037 (I226818,I227169,I226991);
nand I_13038 (I226806,I227169,I227073);
not I_13039 (I227405_rst,I5701);
nand I_13040 (I227422,I179028,I179025);
and I_13041 (I227439,I227422,I179022);
DFFARX1 I_13042  ( .D(I227439), .CLK(I5694_clk), .RSTB(I227405_rst), .Q(I227456) );
not I_13043 (I227473,I227456);
nor I_13044 (I227490,I179046,I179025);
or I_13045 (I227388,I227490,I227456);
not I_13046 (I227376,I227490);
DFFARX1 I_13047  ( .D(I179040), .CLK(I5694_clk), .RSTB(I227405_rst), .Q(I227535) );
nor I_13048 (I227552,I227535,I227490);
nand I_13049 (I227569,I179019,I179031);
and I_13050 (I227586,I227569,I179034);
DFFARX1 I_13051  ( .D(I227586), .CLK(I5694_clk), .RSTB(I227405_rst), .Q(I227603) );
nor I_13052 (I227385,I227603,I227456);
not I_13053 (I227634,I227603);
nor I_13054 (I227651,I227535,I227634);
DFFARX1 I_13055  ( .D(I179043), .CLK(I5694_clk), .RSTB(I227405_rst), .Q(I227668) );
and I_13056 (I227685,I227668,I179049);
or I_13057 (I227394,I227685,I227490);
nand I_13058 (I227373,I227685,I227651);
DFFARX1 I_13059  ( .D(I179037), .CLK(I5694_clk), .RSTB(I227405_rst), .Q(I227730) );
and I_13060 (I227747,I227730,I227473);
nor I_13061 (I227391,I227685,I227747);
nor I_13062 (I227778,I227730,I227535);
DFFARX1 I_13063  ( .D(I227778), .CLK(I5694_clk), .RSTB(I227405_rst), .Q(I227382) );
nor I_13064 (I227397,I227730,I227456);
not I_13065 (I227823,I227730);
nor I_13066 (I227840,I227603,I227823);
and I_13067 (I227857,I227490,I227840);
or I_13068 (I227874,I227685,I227857);
DFFARX1 I_13069  ( .D(I227874), .CLK(I5694_clk), .RSTB(I227405_rst), .Q(I227370) );
nand I_13070 (I227379,I227730,I227552);
nand I_13071 (I227367,I227730,I227634);
not I_13072 (I227966_rst,I5701);
nand I_13073 (I227983,I172444,I172447);
and I_13074 (I228000,I227983,I172429);
DFFARX1 I_13075  ( .D(I228000), .CLK(I5694_clk), .RSTB(I227966_rst), .Q(I228017) );
not I_13076 (I228034,I228017);
nor I_13077 (I228051,I172426,I172447);
or I_13078 (I227949,I228051,I228017);
not I_13079 (I227937,I228051);
DFFARX1 I_13080  ( .D(I172450), .CLK(I5694_clk), .RSTB(I227966_rst), .Q(I228096) );
nor I_13081 (I228113,I228096,I228051);
nand I_13082 (I228130,I172435,I172441);
and I_13083 (I228147,I228130,I172453);
DFFARX1 I_13084  ( .D(I228147), .CLK(I5694_clk), .RSTB(I227966_rst), .Q(I228164) );
nor I_13085 (I227946,I228164,I228017);
not I_13086 (I228195,I228164);
nor I_13087 (I228212,I228096,I228195);
DFFARX1 I_13088  ( .D(I172432), .CLK(I5694_clk), .RSTB(I227966_rst), .Q(I228229) );
and I_13089 (I228246,I228229,I172423);
or I_13090 (I227955,I228246,I228051);
nand I_13091 (I227934,I228246,I228212);
DFFARX1 I_13092  ( .D(I172438), .CLK(I5694_clk), .RSTB(I227966_rst), .Q(I228291) );
and I_13093 (I228308,I228291,I228034);
nor I_13094 (I227952,I228246,I228308);
nor I_13095 (I228339,I228291,I228096);
DFFARX1 I_13096  ( .D(I228339), .CLK(I5694_clk), .RSTB(I227966_rst), .Q(I227943) );
nor I_13097 (I227958,I228291,I228017);
not I_13098 (I228384,I228291);
nor I_13099 (I228401,I228164,I228384);
and I_13100 (I228418,I228051,I228401);
or I_13101 (I228435,I228246,I228418);
DFFARX1 I_13102  ( .D(I228435), .CLK(I5694_clk), .RSTB(I227966_rst), .Q(I227931) );
nand I_13103 (I227940,I228291,I228113);
nand I_13104 (I227928,I228291,I228195);
not I_13105 (I228527_rst,I5701);
not I_13106 (I228544,I191226);
nor I_13107 (I228561,I191223,I191211);
nand I_13108 (I228578,I228561,I191214);
DFFARX1 I_13109  ( .D(I228578), .CLK(I5694_clk), .RSTB(I228527_rst), .Q(I228501) );
nor I_13110 (I228609,I228544,I191223);
nand I_13111 (I228626,I228609,I191220);
not I_13112 (I228516,I228626);
DFFARX1 I_13113  ( .D(I228626), .CLK(I5694_clk), .RSTB(I228527_rst), .Q(I228498) );
not I_13114 (I228671,I191223);
not I_13115 (I228688,I228671);
not I_13116 (I228705,I191232);
nor I_13117 (I228722,I228705,I191208);
and I_13118 (I228739,I228722,I191229);
or I_13119 (I228756,I228739,I191217);
DFFARX1 I_13120  ( .D(I228756), .CLK(I5694_clk), .RSTB(I228527_rst), .Q(I228773) );
nor I_13121 (I228790,I228773,I228626);
nor I_13122 (I228807,I228773,I228688);
nand I_13123 (I228513,I228578,I228807);
nand I_13124 (I228838,I228544,I191232);
nand I_13125 (I228855,I228838,I228773);
and I_13126 (I228872,I228838,I228855);
DFFARX1 I_13127  ( .D(I228872), .CLK(I5694_clk), .RSTB(I228527_rst), .Q(I228495) );
DFFARX1 I_13128  ( .D(I228838), .CLK(I5694_clk), .RSTB(I228527_rst), .Q(I228903) );
and I_13129 (I228492,I228671,I228903);
DFFARX1 I_13130  ( .D(I191238), .CLK(I5694_clk), .RSTB(I228527_rst), .Q(I228934) );
not I_13131 (I228951,I228934);
nor I_13132 (I228968,I228626,I228951);
and I_13133 (I228985,I228934,I228968);
nand I_13134 (I228507,I228934,I228688);
DFFARX1 I_13135  ( .D(I228934), .CLK(I5694_clk), .RSTB(I228527_rst), .Q(I229016) );
not I_13136 (I228504,I229016);
DFFARX1 I_13137  ( .D(I191235), .CLK(I5694_clk), .RSTB(I228527_rst), .Q(I229047) );
not I_13138 (I229064,I229047);
or I_13139 (I229081,I229064,I228985);
DFFARX1 I_13140  ( .D(I229081), .CLK(I5694_clk), .RSTB(I228527_rst), .Q(I228510) );
nand I_13141 (I228519,I229064,I228790);
DFFARX1 I_13142  ( .D(I229064), .CLK(I5694_clk), .RSTB(I228527_rst), .Q(I228489) );
not I_13143 (I229173_rst,I5701);
not I_13144 (I229190,I198349);
nor I_13145 (I229207,I198331,I198346);
nand I_13146 (I229224,I229207,I198355);
DFFARX1 I_13147  ( .D(I229224), .CLK(I5694_clk), .RSTB(I229173_rst), .Q(I229147) );
nor I_13148 (I229255,I229190,I198331);
nand I_13149 (I229272,I229255,I198358);
not I_13150 (I229162,I229272);
DFFARX1 I_13151  ( .D(I229272), .CLK(I5694_clk), .RSTB(I229173_rst), .Q(I229144) );
not I_13152 (I229317,I198331);
not I_13153 (I229334,I229317);
not I_13154 (I229351,I198361);
nor I_13155 (I229368,I229351,I198337);
and I_13156 (I229385,I229368,I198340);
or I_13157 (I229402,I229385,I198334);
DFFARX1 I_13158  ( .D(I229402), .CLK(I5694_clk), .RSTB(I229173_rst), .Q(I229419) );
nor I_13159 (I229436,I229419,I229272);
nor I_13160 (I229453,I229419,I229334);
nand I_13161 (I229159,I229224,I229453);
nand I_13162 (I229484,I229190,I198361);
nand I_13163 (I229501,I229484,I229419);
and I_13164 (I229518,I229484,I229501);
DFFARX1 I_13165  ( .D(I229518), .CLK(I5694_clk), .RSTB(I229173_rst), .Q(I229141) );
DFFARX1 I_13166  ( .D(I229484), .CLK(I5694_clk), .RSTB(I229173_rst), .Q(I229549) );
and I_13167 (I229138,I229317,I229549);
DFFARX1 I_13168  ( .D(I198343), .CLK(I5694_clk), .RSTB(I229173_rst), .Q(I229580) );
not I_13169 (I229597,I229580);
nor I_13170 (I229614,I229272,I229597);
and I_13171 (I229631,I229580,I229614);
nand I_13172 (I229153,I229580,I229334);
DFFARX1 I_13173  ( .D(I229580), .CLK(I5694_clk), .RSTB(I229173_rst), .Q(I229662) );
not I_13174 (I229150,I229662);
DFFARX1 I_13175  ( .D(I198352), .CLK(I5694_clk), .RSTB(I229173_rst), .Q(I229693) );
not I_13176 (I229710,I229693);
or I_13177 (I229727,I229710,I229631);
DFFARX1 I_13178  ( .D(I229727), .CLK(I5694_clk), .RSTB(I229173_rst), .Q(I229156) );
nand I_13179 (I229165,I229710,I229436);
DFFARX1 I_13180  ( .D(I229710), .CLK(I5694_clk), .RSTB(I229173_rst), .Q(I229135) );
not I_13181 (I229819_rst,I5701);
not I_13182 (I229836,I187911);
nor I_13183 (I229853,I187908,I187896);
nand I_13184 (I229870,I229853,I187899);
DFFARX1 I_13185  ( .D(I229870), .CLK(I5694_clk), .RSTB(I229819_rst), .Q(I229793) );
nor I_13186 (I229901,I229836,I187908);
nand I_13187 (I229918,I229901,I187905);
not I_13188 (I229808,I229918);
DFFARX1 I_13189  ( .D(I229918), .CLK(I5694_clk), .RSTB(I229819_rst), .Q(I229790) );
not I_13190 (I229963,I187908);
not I_13191 (I229980,I229963);
not I_13192 (I229997,I187917);
nor I_13193 (I230014,I229997,I187893);
and I_13194 (I230031,I230014,I187914);
or I_13195 (I230048,I230031,I187902);
DFFARX1 I_13196  ( .D(I230048), .CLK(I5694_clk), .RSTB(I229819_rst), .Q(I230065) );
nor I_13197 (I230082,I230065,I229918);
nor I_13198 (I230099,I230065,I229980);
nand I_13199 (I229805,I229870,I230099);
nand I_13200 (I230130,I229836,I187917);
nand I_13201 (I230147,I230130,I230065);
and I_13202 (I230164,I230130,I230147);
DFFARX1 I_13203  ( .D(I230164), .CLK(I5694_clk), .RSTB(I229819_rst), .Q(I229787) );
DFFARX1 I_13204  ( .D(I230130), .CLK(I5694_clk), .RSTB(I229819_rst), .Q(I230195) );
and I_13205 (I229784,I229963,I230195);
DFFARX1 I_13206  ( .D(I187923), .CLK(I5694_clk), .RSTB(I229819_rst), .Q(I230226) );
not I_13207 (I230243,I230226);
nor I_13208 (I230260,I229918,I230243);
and I_13209 (I230277,I230226,I230260);
nand I_13210 (I229799,I230226,I229980);
DFFARX1 I_13211  ( .D(I230226), .CLK(I5694_clk), .RSTB(I229819_rst), .Q(I230308) );
not I_13212 (I229796,I230308);
DFFARX1 I_13213  ( .D(I187920), .CLK(I5694_clk), .RSTB(I229819_rst), .Q(I230339) );
not I_13214 (I230356,I230339);
or I_13215 (I230373,I230356,I230277);
DFFARX1 I_13216  ( .D(I230373), .CLK(I5694_clk), .RSTB(I229819_rst), .Q(I229802) );
nand I_13217 (I229811,I230356,I230082);
DFFARX1 I_13218  ( .D(I230356), .CLK(I5694_clk), .RSTB(I229819_rst), .Q(I229781) );
not I_13219 (I230465_rst,I5701);
not I_13220 (I23048_rst2,I189900);
nor I_13221 (I230499,I189897,I189885);
nand I_13222 (I230516,I230499,I189888);
DFFARX1 I_13223  ( .D(I230516), .CLK(I5694_clk), .RSTB(I230465_rst), .Q(I230439) );
nor I_13224 (I230547,I23048_rst2,I189897);
nand I_13225 (I230564,I230547,I189894);
not I_13226 (I230454,I230564);
DFFARX1 I_13227  ( .D(I230564), .CLK(I5694_clk), .RSTB(I230465_rst), .Q(I230436) );
not I_13228 (I230609,I189897);
not I_13229 (I230626,I230609);
not I_13230 (I230643,I189906);
nor I_13231 (I230660,I230643,I189882);
and I_13232 (I230677,I230660,I189903);
or I_13233 (I230694,I230677,I189891);
DFFARX1 I_13234  ( .D(I230694), .CLK(I5694_clk), .RSTB(I230465_rst), .Q(I230711) );
nor I_13235 (I230728,I230711,I230564);
nor I_13236 (I230745,I230711,I230626);
nand I_13237 (I230451,I230516,I230745);
nand I_13238 (I230776,I23048_rst2,I189906);
nand I_13239 (I230793,I230776,I230711);
and I_13240 (I230810,I230776,I230793);
DFFARX1 I_13241  ( .D(I230810), .CLK(I5694_clk), .RSTB(I230465_rst), .Q(I230433) );
DFFARX1 I_13242  ( .D(I230776), .CLK(I5694_clk), .RSTB(I230465_rst), .Q(I230841) );
and I_13243 (I230430,I230609,I230841);
DFFARX1 I_13244  ( .D(I189912), .CLK(I5694_clk), .RSTB(I230465_rst), .Q(I230872) );
not I_13245 (I230889,I230872);
nor I_13246 (I230906,I230564,I230889);
and I_13247 (I230923,I230872,I230906);
nand I_13248 (I230445,I230872,I230626);
DFFARX1 I_13249  ( .D(I230872), .CLK(I5694_clk), .RSTB(I230465_rst), .Q(I230954) );
not I_13250 (I230442,I230954);
DFFARX1 I_13251  ( .D(I189909), .CLK(I5694_clk), .RSTB(I230465_rst), .Q(I230985) );
not I_13252 (I231002,I230985);
or I_13253 (I231019,I231002,I230923);
DFFARX1 I_13254  ( .D(I231019), .CLK(I5694_clk), .RSTB(I230465_rst), .Q(I230448) );
nand I_13255 (I230457,I231002,I230728);
DFFARX1 I_13256  ( .D(I231002), .CLK(I5694_clk), .RSTB(I230465_rst), .Q(I230427) );
not I_13257 (I231111_rst,I5701);
not I_13258 (I231128,I212519);
nor I_13259 (I231145,I212495,I212501);
nand I_13260 (I231162,I231145,I212504);
DFFARX1 I_13261  ( .D(I231162), .CLK(I5694_clk), .RSTB(I231111_rst), .Q(I231085) );
nor I_13262 (I231193,I231128,I212495);
nand I_13263 (I231210,I231193,I212513);
not I_13264 (I231100,I231210);
DFFARX1 I_13265  ( .D(I231210), .CLK(I5694_clk), .RSTB(I231111_rst), .Q(I231082) );
not I_13266 (I231255,I212495);
not I_13267 (I231272,I231255);
not I_13268 (I231289,I212492);
nor I_13269 (I231306,I231289,I212507);
and I_13270 (I231323,I231306,I212498);
or I_13271 (I231340,I231323,I212510);
DFFARX1 I_13272  ( .D(I231340), .CLK(I5694_clk), .RSTB(I231111_rst), .Q(I231357) );
nor I_13273 (I231374,I231357,I231210);
nor I_13274 (I231391,I231357,I231272);
nand I_13275 (I231097,I231162,I231391);
nand I_13276 (I231422,I231128,I212492);
nand I_13277 (I231439,I231422,I231357);
and I_13278 (I231456,I231422,I231439);
DFFARX1 I_13279  ( .D(I231456), .CLK(I5694_clk), .RSTB(I231111_rst), .Q(I231079) );
DFFARX1 I_13280  ( .D(I231422), .CLK(I5694_clk), .RSTB(I231111_rst), .Q(I231487) );
and I_13281 (I231076,I231255,I231487);
DFFARX1 I_13282  ( .D(I212522), .CLK(I5694_clk), .RSTB(I231111_rst), .Q(I231518) );
not I_13283 (I231535,I231518);
nor I_13284 (I231552,I231210,I231535);
and I_13285 (I231569,I231518,I231552);
nand I_13286 (I231091,I231518,I231272);
DFFARX1 I_13287  ( .D(I231518), .CLK(I5694_clk), .RSTB(I231111_rst), .Q(I231600) );
not I_13288 (I231088,I231600);
DFFARX1 I_13289  ( .D(I212516), .CLK(I5694_clk), .RSTB(I231111_rst), .Q(I231631) );
not I_13290 (I231648,I231631);
or I_13291 (I231665,I231648,I231569);
DFFARX1 I_13292  ( .D(I231665), .CLK(I5694_clk), .RSTB(I231111_rst), .Q(I231094) );
nand I_13293 (I231103,I231648,I231374);
DFFARX1 I_13294  ( .D(I231648), .CLK(I5694_clk), .RSTB(I231111_rst), .Q(I231073) );
not I_13295 (I231757_rst,I5701);
not I_13296 (I231774,I225676);
nor I_13297 (I231791,I225673,I225670);
nand I_13298 (I231808,I231791,I225691);
DFFARX1 I_13299  ( .D(I231808), .CLK(I5694_clk), .RSTB(I231757_rst), .Q(I231731) );
nor I_13300 (I231839,I231774,I225673);
nand I_13301 (I231856,I231839,I225694);
not I_13302 (I231746,I231856);
DFFARX1 I_13303  ( .D(I231856), .CLK(I5694_clk), .RSTB(I231757_rst), .Q(I231728) );
not I_13304 (I231901,I225673);
not I_13305 (I231918,I231901);
not I_13306 (I231935,I225667);
nor I_13307 (I231952,I231935,I225679);
and I_13308 (I231969,I231952,I225688);
or I_13309 (I231986,I231969,I225682);
DFFARX1 I_13310  ( .D(I231986), .CLK(I5694_clk), .RSTB(I231757_rst), .Q(I232003) );
nor I_13311 (I232020,I232003,I231856);
nor I_13312 (I232037,I232003,I231918);
nand I_13313 (I231743,I231808,I232037);
nand I_13314 (I232068,I231774,I225667);
nand I_13315 (I232085,I232068,I232003);
and I_13316 (I232102,I232068,I232085);
DFFARX1 I_13317  ( .D(I232102), .CLK(I5694_clk), .RSTB(I231757_rst), .Q(I231725) );
DFFARX1 I_13318  ( .D(I232068), .CLK(I5694_clk), .RSTB(I231757_rst), .Q(I232133) );
and I_13319 (I231722,I231901,I232133);
DFFARX1 I_13320  ( .D(I225697), .CLK(I5694_clk), .RSTB(I231757_rst), .Q(I232164) );
not I_13321 (I232181,I232164);
nor I_13322 (I232198,I231856,I232181);
and I_13323 (I232215,I232164,I232198);
nand I_13324 (I231737,I232164,I231918);
DFFARX1 I_13325  ( .D(I232164), .CLK(I5694_clk), .RSTB(I231757_rst), .Q(I232246) );
not I_13326 (I231734,I232246);
DFFARX1 I_13327  ( .D(I225685), .CLK(I5694_clk), .RSTB(I231757_rst), .Q(I232277) );
not I_13328 (I232294,I232277);
or I_13329 (I232311,I232294,I232215);
DFFARX1 I_13330  ( .D(I232311), .CLK(I5694_clk), .RSTB(I231757_rst), .Q(I231740) );
nand I_13331 (I231749,I232294,I232020);
DFFARX1 I_13332  ( .D(I232294), .CLK(I5694_clk), .RSTB(I231757_rst), .Q(I231719) );
not I_13333 (I232403_rst,I5701);
not I_13334 (I232420,I214292);
nor I_13335 (I232437,I214277,I214304);
nand I_13336 (I232454,I232437,I214280);
DFFARX1 I_13337  ( .D(I232454), .CLK(I5694_clk), .RSTB(I232403_rst), .Q(I232377) );
nor I_13338 (I232485,I232420,I214277);
nand I_13339 (I232502,I232485,I214295);
not I_13340 (I232392,I232502);
DFFARX1 I_13341  ( .D(I232502), .CLK(I5694_clk), .RSTB(I232403_rst), .Q(I232374) );
not I_13342 (I232547,I214277);
not I_13343 (I232564,I232547);
not I_13344 (I232581,I214307);
nor I_13345 (I232598,I232581,I214289);
and I_13346 (I232615,I232598,I214298);
or I_13347 (I232632,I232615,I214283);
DFFARX1 I_13348  ( .D(I232632), .CLK(I5694_clk), .RSTB(I232403_rst), .Q(I232649) );
nor I_13349 (I232666,I232649,I232502);
nor I_13350 (I232683,I232649,I232564);
nand I_13351 (I232389,I232454,I232683);
nand I_13352 (I232714,I232420,I214307);
nand I_13353 (I232731,I232714,I232649);
and I_13354 (I232748,I232714,I232731);
DFFARX1 I_13355  ( .D(I232748), .CLK(I5694_clk), .RSTB(I232403_rst), .Q(I232371) );
DFFARX1 I_13356  ( .D(I232714), .CLK(I5694_clk), .RSTB(I232403_rst), .Q(I232779) );
and I_13357 (I232368,I232547,I232779);
DFFARX1 I_13358  ( .D(I214286), .CLK(I5694_clk), .RSTB(I232403_rst), .Q(I232810) );
not I_13359 (I232827,I232810);
nor I_13360 (I232844,I232502,I232827);
and I_13361 (I232861,I232810,I232844);
nand I_13362 (I232383,I232810,I232564);
DFFARX1 I_13363  ( .D(I232810), .CLK(I5694_clk), .RSTB(I232403_rst), .Q(I232892) );
not I_13364 (I232380,I232892);
DFFARX1 I_13365  ( .D(I214301), .CLK(I5694_clk), .RSTB(I232403_rst), .Q(I232923) );
not I_13366 (I232940,I232923);
or I_13367 (I232957,I232940,I232861);
DFFARX1 I_13368  ( .D(I232957), .CLK(I5694_clk), .RSTB(I232403_rst), .Q(I232386) );
nand I_13369 (I232395,I232940,I232666);
DFFARX1 I_13370  ( .D(I232940), .CLK(I5694_clk), .RSTB(I232403_rst), .Q(I232365) );
not I_13371 (I233049_rst,I5701);
not I_13372 (I233066,I181467);
nor I_13373 (I233083,I181497,I181476);
nand I_13374 (I233100,I233083,I181488);
DFFARX1 I_13375  ( .D(I233100), .CLK(I5694_clk), .RSTB(I233049_rst), .Q(I233023) );
nor I_13376 (I233131,I233066,I181497);
nand I_13377 (I233148,I233131,I181470);
not I_13378 (I233038,I233148);
DFFARX1 I_13379  ( .D(I233148), .CLK(I5694_clk), .RSTB(I233049_rst), .Q(I233020) );
not I_13380 (I233193,I181497);
not I_13381 (I233210,I233193);
not I_13382 (I233227,I181473);
nor I_13383 (I233244,I233227,I181491);
and I_13384 (I233261,I233244,I181482);
or I_13385 (I233278,I233261,I181479);
DFFARX1 I_13386  ( .D(I233278), .CLK(I5694_clk), .RSTB(I233049_rst), .Q(I233295) );
nor I_13387 (I233312,I233295,I233148);
nor I_13388 (I233329,I233295,I233210);
nand I_13389 (I233035,I233100,I233329);
nand I_13390 (I233360,I233066,I181473);
nand I_13391 (I233377,I233360,I233295);
and I_13392 (I233394,I233360,I233377);
DFFARX1 I_13393  ( .D(I233394), .CLK(I5694_clk), .RSTB(I233049_rst), .Q(I233017) );
DFFARX1 I_13394  ( .D(I233360), .CLK(I5694_clk), .RSTB(I233049_rst), .Q(I233425) );
and I_13395 (I233014,I233193,I233425);
DFFARX1 I_13396  ( .D(I181485), .CLK(I5694_clk), .RSTB(I233049_rst), .Q(I233456) );
not I_13397 (I233473,I233456);
nor I_13398 (I233490,I233148,I233473);
and I_13399 (I233507,I233456,I233490);
nand I_13400 (I233029,I233456,I233210);
DFFARX1 I_13401  ( .D(I233456), .CLK(I5694_clk), .RSTB(I233049_rst), .Q(I233538) );
not I_13402 (I233026,I233538);
DFFARX1 I_13403  ( .D(I181494), .CLK(I5694_clk), .RSTB(I233049_rst), .Q(I233569) );
not I_13404 (I233586,I233569);
or I_13405 (I233603,I233586,I233507);
DFFARX1 I_13406  ( .D(I233603), .CLK(I5694_clk), .RSTB(I233049_rst), .Q(I233032) );
nand I_13407 (I233041,I233586,I233312);
DFFARX1 I_13408  ( .D(I233586), .CLK(I5694_clk), .RSTB(I233049_rst), .Q(I233011) );
not I_13409 (I233695_rst,I5701);
not I_13410 (I233712,I193861);
nor I_13411 (I233729,I193873,I193855);
nand I_13412 (I233746,I233729,I193870);
DFFARX1 I_13413  ( .D(I233746), .CLK(I5694_clk), .RSTB(I233695_rst), .Q(I233669) );
nor I_13414 (I233777,I233712,I193873);
nand I_13415 (I233794,I233777,I193858);
not I_13416 (I233684,I233794);
DFFARX1 I_13417  ( .D(I233794), .CLK(I5694_clk), .RSTB(I233695_rst), .Q(I233666) );
not I_13418 (I233839,I193873);
not I_13419 (I233856,I233839);
not I_13420 (I233873,I193867);
nor I_13421 (I233890,I233873,I193846);
and I_13422 (I233907,I233890,I193849);
or I_13423 (I233924,I233907,I193852);
DFFARX1 I_13424  ( .D(I233924), .CLK(I5694_clk), .RSTB(I233695_rst), .Q(I233941) );
nor I_13425 (I233958,I233941,I233794);
nor I_13426 (I233975,I233941,I233856);
nand I_13427 (I233681,I233746,I233975);
nand I_13428 (I234006,I233712,I193867);
nand I_13429 (I234023,I234006,I233941);
and I_13430 (I234040,I234006,I234023);
DFFARX1 I_13431  ( .D(I234040), .CLK(I5694_clk), .RSTB(I233695_rst), .Q(I233663) );
DFFARX1 I_13432  ( .D(I234006), .CLK(I5694_clk), .RSTB(I233695_rst), .Q(I234071) );
and I_13433 (I233660,I233839,I234071);
DFFARX1 I_13434  ( .D(I193843), .CLK(I5694_clk), .RSTB(I233695_rst), .Q(I234102) );
not I_13435 (I234119,I234102);
nor I_13436 (I234136,I233794,I234119);
and I_13437 (I234153,I234102,I234136);
nand I_13438 (I233675,I234102,I233856);
DFFARX1 I_13439  ( .D(I234102), .CLK(I5694_clk), .RSTB(I233695_rst), .Q(I234184) );
not I_13440 (I233672,I234184);
DFFARX1 I_13441  ( .D(I193864), .CLK(I5694_clk), .RSTB(I233695_rst), .Q(I234215) );
not I_13442 (I234232,I234215);
or I_13443 (I234249,I234232,I234153);
DFFARX1 I_13444  ( .D(I234249), .CLK(I5694_clk), .RSTB(I233695_rst), .Q(I233678) );
nand I_13445 (I233687,I234232,I233958);
DFFARX1 I_13446  ( .D(I234232), .CLK(I5694_clk), .RSTB(I233695_rst), .Q(I233657) );
not I_13447 (I234341_rst,I5701);
not I_13448 (I234358,I197737);
nor I_13449 (I234375,I197719,I197734);
nand I_13450 (I234392,I234375,I197743);
DFFARX1 I_13451  ( .D(I234392), .CLK(I5694_clk), .RSTB(I234341_rst), .Q(I234315) );
nor I_13452 (I234423,I234358,I197719);
nand I_13453 (I234440,I234423,I197746);
not I_13454 (I234330,I234440);
DFFARX1 I_13455  ( .D(I234440), .CLK(I5694_clk), .RSTB(I234341_rst), .Q(I234312) );
not I_13456 (I234485,I197719);
not I_13457 (I234502,I234485);
not I_13458 (I234519,I197749);
nor I_13459 (I234536,I234519,I197725);
and I_13460 (I234553,I234536,I197728);
or I_13461 (I234570,I234553,I197722);
DFFARX1 I_13462  ( .D(I234570), .CLK(I5694_clk), .RSTB(I234341_rst), .Q(I234587) );
nor I_13463 (I234604,I234587,I234440);
nor I_13464 (I234621,I234587,I234502);
nand I_13465 (I234327,I234392,I234621);
nand I_13466 (I234652,I234358,I197749);
nand I_13467 (I234669,I234652,I234587);
and I_13468 (I234686,I234652,I234669);
DFFARX1 I_13469  ( .D(I234686), .CLK(I5694_clk), .RSTB(I234341_rst), .Q(I234309) );
DFFARX1 I_13470  ( .D(I234652), .CLK(I5694_clk), .RSTB(I234341_rst), .Q(I234717) );
and I_13471 (I234306,I234485,I234717);
DFFARX1 I_13472  ( .D(I197731), .CLK(I5694_clk), .RSTB(I234341_rst), .Q(I234748) );
not I_13473 (I234765,I234748);
nor I_13474 (I234782,I234440,I234765);
and I_13475 (I234799,I234748,I234782);
nand I_13476 (I234321,I234748,I234502);
DFFARX1 I_13477  ( .D(I234748), .CLK(I5694_clk), .RSTB(I234341_rst), .Q(I234830) );
not I_13478 (I234318,I234830);
DFFARX1 I_13479  ( .D(I197740), .CLK(I5694_clk), .RSTB(I234341_rst), .Q(I234861) );
not I_13480 (I234878,I234861);
or I_13481 (I234895,I234878,I234799);
DFFARX1 I_13482  ( .D(I234895), .CLK(I5694_clk), .RSTB(I234341_rst), .Q(I234324) );
nand I_13483 (I234333,I234878,I234604);
DFFARX1 I_13484  ( .D(I234878), .CLK(I5694_clk), .RSTB(I234341_rst), .Q(I234303) );
not I_13485 (I234987_rst,I5701);
not I_13486 (I235004,I196445);
nor I_13487 (I235021,I196457,I196439);
nand I_13488 (I235038,I235021,I196454);
DFFARX1 I_13489  ( .D(I235038), .CLK(I5694_clk), .RSTB(I234987_rst), .Q(I234961) );
nor I_13490 (I235069,I235004,I196457);
nand I_13491 (I235086,I235069,I196442);
not I_13492 (I234976,I235086);
DFFARX1 I_13493  ( .D(I235086), .CLK(I5694_clk), .RSTB(I234987_rst), .Q(I234958) );
not I_13494 (I235131,I196457);
not I_13495 (I235148,I235131);
not I_13496 (I235165,I196451);
nor I_13497 (I235182,I235165,I196430);
and I_13498 (I235199,I235182,I196433);
or I_13499 (I235216,I235199,I196436);
DFFARX1 I_13500  ( .D(I235216), .CLK(I5694_clk), .RSTB(I234987_rst), .Q(I235233) );
nor I_13501 (I235250,I235233,I235086);
nor I_13502 (I235267,I235233,I235148);
nand I_13503 (I234973,I235038,I235267);
nand I_13504 (I235298,I235004,I196451);
nand I_13505 (I235315,I235298,I235233);
and I_13506 (I235332,I235298,I235315);
DFFARX1 I_13507  ( .D(I235332), .CLK(I5694_clk), .RSTB(I234987_rst), .Q(I234955) );
DFFARX1 I_13508  ( .D(I235298), .CLK(I5694_clk), .RSTB(I234987_rst), .Q(I235363) );
and I_13509 (I234952,I235131,I235363);
DFFARX1 I_13510  ( .D(I196427), .CLK(I5694_clk), .RSTB(I234987_rst), .Q(I235394) );
not I_13511 (I235411,I235394);
nor I_13512 (I235428,I235086,I235411);
and I_13513 (I235445,I235394,I235428);
nand I_13514 (I234967,I235394,I235148);
DFFARX1 I_13515  ( .D(I235394), .CLK(I5694_clk), .RSTB(I234987_rst), .Q(I235476) );
not I_13516 (I234964,I235476);
DFFARX1 I_13517  ( .D(I196448), .CLK(I5694_clk), .RSTB(I234987_rst), .Q(I235507) );
not I_13518 (I235524,I235507);
or I_13519 (I235541,I235524,I235445);
DFFARX1 I_13520  ( .D(I235541), .CLK(I5694_clk), .RSTB(I234987_rst), .Q(I234970) );
nand I_13521 (I234979,I235524,I235250);
DFFARX1 I_13522  ( .D(I235524), .CLK(I5694_clk), .RSTB(I234987_rst), .Q(I234949) );
not I_13523 (I235633_rst,I5701);
not I_13524 (I235650,I222786);
nor I_13525 (I235667,I222783,I222780);
nand I_13526 (I235684,I235667,I222801);
DFFARX1 I_13527  ( .D(I235684), .CLK(I5694_clk), .RSTB(I235633_rst), .Q(I235607) );
nor I_13528 (I235715,I235650,I222783);
nand I_13529 (I235732,I235715,I222804);
not I_13530 (I235622,I235732);
DFFARX1 I_13531  ( .D(I235732), .CLK(I5694_clk), .RSTB(I235633_rst), .Q(I235604) );
not I_13532 (I235777,I222783);
not I_13533 (I235794,I235777);
not I_13534 (I235811,I222777);
nor I_13535 (I235828,I235811,I222789);
and I_13536 (I235845,I235828,I222798);
or I_13537 (I235862,I235845,I222792);
DFFARX1 I_13538  ( .D(I235862), .CLK(I5694_clk), .RSTB(I235633_rst), .Q(I235879) );
nor I_13539 (I235896,I235879,I235732);
nor I_13540 (I235913,I235879,I235794);
nand I_13541 (I235619,I235684,I235913);
nand I_13542 (I235944,I235650,I222777);
nand I_13543 (I235961,I235944,I235879);
and I_13544 (I235978,I235944,I235961);
DFFARX1 I_13545  ( .D(I235978), .CLK(I5694_clk), .RSTB(I235633_rst), .Q(I235601) );
DFFARX1 I_13546  ( .D(I235944), .CLK(I5694_clk), .RSTB(I235633_rst), .Q(I236009) );
and I_13547 (I235598,I235777,I236009);
DFFARX1 I_13548  ( .D(I222807), .CLK(I5694_clk), .RSTB(I235633_rst), .Q(I236040) );
not I_13549 (I236057,I236040);
nor I_13550 (I236074,I235732,I236057);
and I_13551 (I236091,I236040,I236074);
nand I_13552 (I235613,I236040,I235794);
DFFARX1 I_13553  ( .D(I236040), .CLK(I5694_clk), .RSTB(I235633_rst), .Q(I236122) );
not I_13554 (I235610,I236122);
DFFARX1 I_13555  ( .D(I222795), .CLK(I5694_clk), .RSTB(I235633_rst), .Q(I236153) );
not I_13556 (I236170,I236153);
or I_13557 (I236187,I236170,I236091);
DFFARX1 I_13558  ( .D(I236187), .CLK(I5694_clk), .RSTB(I235633_rst), .Q(I235616) );
nand I_13559 (I235625,I236170,I235896);
DFFARX1 I_13560  ( .D(I236170), .CLK(I5694_clk), .RSTB(I235633_rst), .Q(I235595) );
not I_13561 (I236279_rst,I5701);
not I_13562 (I236296,I210734);
nor I_13563 (I236313,I210710,I210716);
nand I_13564 (I236330,I236313,I210719);
DFFARX1 I_13565  ( .D(I236330), .CLK(I5694_clk), .RSTB(I236279_rst), .Q(I236253) );
nor I_13566 (I236361,I236296,I210710);
nand I_13567 (I236378,I236361,I210728);
not I_13568 (I23626_rst8,I236378);
DFFARX1 I_13569  ( .D(I236378), .CLK(I5694_clk), .RSTB(I236279_rst), .Q(I236250) );
not I_13570 (I236423,I210710);
not I_13571 (I236440,I236423);
not I_13572 (I236457,I210707);
nor I_13573 (I236474,I236457,I210722);
and I_13574 (I236491,I236474,I210713);
or I_13575 (I236508,I236491,I210725);
DFFARX1 I_13576  ( .D(I236508), .CLK(I5694_clk), .RSTB(I236279_rst), .Q(I236525) );
nor I_13577 (I236542,I236525,I236378);
nor I_13578 (I236559,I236525,I236440);
nand I_13579 (I23626_rst5,I236330,I236559);
nand I_13580 (I236590,I236296,I210707);
nand I_13581 (I236607,I236590,I236525);
and I_13582 (I236624,I236590,I236607);
DFFARX1 I_13583  ( .D(I236624), .CLK(I5694_clk), .RSTB(I236279_rst), .Q(I236247) );
DFFARX1 I_13584  ( .D(I236590), .CLK(I5694_clk), .RSTB(I236279_rst), .Q(I236655) );
and I_13585 (I236244,I236423,I236655);
DFFARX1 I_13586  ( .D(I210737), .CLK(I5694_clk), .RSTB(I236279_rst), .Q(I236686) );
not I_13587 (I236703,I236686);
nor I_13588 (I236720,I236378,I236703);
and I_13589 (I236737,I236686,I236720);
nand I_13590 (I236259,I236686,I236440);
DFFARX1 I_13591  ( .D(I236686), .CLK(I5694_clk), .RSTB(I236279_rst), .Q(I236768) );
not I_13592 (I236256,I236768);
DFFARX1 I_13593  ( .D(I210731), .CLK(I5694_clk), .RSTB(I236279_rst), .Q(I236799) );
not I_13594 (I236816,I236799);
or I_13595 (I236833,I236816,I236737);
DFFARX1 I_13596  ( .D(I236833), .CLK(I5694_clk), .RSTB(I236279_rst), .Q(I23626_rst2) );
nand I_13597 (I236271,I236816,I236542);
DFFARX1 I_13598  ( .D(I236816), .CLK(I5694_clk), .RSTB(I236279_rst), .Q(I236241) );
not I_13599 (I236925_rst,I5701);
not I_13600 (I236942,I217859);
nor I_13601 (I236959,I217865,I217877);
nand I_13602 (I236976,I236959,I217868);
DFFARX1 I_13603  ( .D(I236976), .CLK(I5694_clk), .RSTB(I236925_rst), .Q(I236896) );
nor I_13604 (I237007,I236942,I217865);
nand I_13605 (I237024,I237007,I217847);
nand I_13606 (I237041,I237024,I236976);
not I_13607 (I237058,I217865);
not I_13608 (I237075,I217862);
nor I_13609 (I237092,I237075,I217850);
and I_13610 (I237109,I237092,I217871);
or I_13611 (I237126,I237109,I217853);
DFFARX1 I_13612  ( .D(I237126), .CLK(I5694_clk), .RSTB(I236925_rst), .Q(I237143) );
nor I_13613 (I237160,I237143,I237024);
nand I_13614 (I236911,I237058,I237160);
not I_13615 (I236908,I237143);
and I_13616 (I237205,I237143,I237041);
DFFARX1 I_13617  ( .D(I237205), .CLK(I5694_clk), .RSTB(I236925_rst), .Q(I236893) );
DFFARX1 I_13618  ( .D(I237143), .CLK(I5694_clk), .RSTB(I236925_rst), .Q(I237236) );
and I_13619 (I236890,I237058,I237236);
nand I_13620 (I237267,I236942,I217862);
not I_13621 (I237284,I237267);
nor I_13622 (I237301,I237143,I237284);
DFFARX1 I_13623  ( .D(I217874), .CLK(I5694_clk), .RSTB(I236925_rst), .Q(I237318) );
nand I_13624 (I237335,I237318,I237267);
and I_13625 (I237352,I237058,I237335);
DFFARX1 I_13626  ( .D(I237352), .CLK(I5694_clk), .RSTB(I236925_rst), .Q(I236917) );
not I_13627 (I237383,I237318);
nand I_13628 (I236905,I237318,I237301);
nand I_13629 (I236899,I237318,I237284);
DFFARX1 I_13630  ( .D(I217856), .CLK(I5694_clk), .RSTB(I236925_rst), .Q(I237428) );
not I_13631 (I237445,I237428);
nor I_13632 (I236914,I237318,I237445);
nor I_13633 (I237476,I237445,I237383);
and I_13634 (I237493,I237024,I237476);
or I_13635 (I237510,I237267,I237493);
DFFARX1 I_13636  ( .D(I237510), .CLK(I5694_clk), .RSTB(I236925_rst), .Q(I236902) );
DFFARX1 I_13637  ( .D(I237445), .CLK(I5694_clk), .RSTB(I236925_rst), .Q(I236887) );
not I_13638 (I237588_rst,I5701);
not I_13639 (I237605,I183252);
nor I_13640 (I237622,I183261,I183273);
nand I_13641 (I237639,I237622,I183264);
DFFARX1 I_13642  ( .D(I237639), .CLK(I5694_clk), .RSTB(I237588_rst), .Q(I237559) );
nor I_13643 (I237670,I237605,I183261);
nand I_13644 (I237687,I237670,I183276);
nand I_13645 (I237704,I237687,I237639);
not I_13646 (I237721,I183261);
not I_13647 (I237738,I183282);
nor I_13648 (I237755,I237738,I183258);
and I_13649 (I237772,I237755,I183267);
or I_13650 (I237789,I237772,I183255);
DFFARX1 I_13651  ( .D(I237789), .CLK(I5694_clk), .RSTB(I237588_rst), .Q(I237806) );
nor I_13652 (I237823,I237806,I237687);
nand I_13653 (I237574,I237721,I237823);
not I_13654 (I237571,I237806);
and I_13655 (I237868,I237806,I237704);
DFFARX1 I_13656  ( .D(I237868), .CLK(I5694_clk), .RSTB(I237588_rst), .Q(I237556) );
DFFARX1 I_13657  ( .D(I237806), .CLK(I5694_clk), .RSTB(I237588_rst), .Q(I237899) );
and I_13658 (I237553,I237721,I237899);
nand I_13659 (I237930,I237605,I183282);
not I_13660 (I237947,I237930);
nor I_13661 (I237964,I237806,I237947);
DFFARX1 I_13662  ( .D(I183279), .CLK(I5694_clk), .RSTB(I237588_rst), .Q(I237981) );
nand I_13663 (I237998,I237981,I237930);
and I_13664 (I238015,I237721,I237998);
DFFARX1 I_13665  ( .D(I238015), .CLK(I5694_clk), .RSTB(I237588_rst), .Q(I237580) );
not I_13666 (I238046,I237981);
nand I_13667 (I237568,I237981,I237964);
nand I_13668 (I237562,I237981,I237947);
DFFARX1 I_13669  ( .D(I183270), .CLK(I5694_clk), .RSTB(I237588_rst), .Q(I238091) );
not I_13670 (I238108,I238091);
nor I_13671 (I237577,I237981,I238108);
nor I_13672 (I238139,I238108,I238046);
and I_13673 (I238156,I237687,I238139);
or I_13674 (I238173,I237930,I238156);
DFFARX1 I_13675  ( .D(I238173), .CLK(I5694_clk), .RSTB(I237588_rst), .Q(I237565) );
DFFARX1 I_13676  ( .D(I238108), .CLK(I5694_clk), .RSTB(I237588_rst), .Q(I237550) );
not I_13677 (I238251_rst,I5701);
not I_13678 (I238268,I219746);
nor I_13679 (I238285,I219752,I219764);
nand I_13680 (I238302,I238285,I219755);
DFFARX1 I_13681  ( .D(I238302), .CLK(I5694_clk), .RSTB(I238251_rst), .Q(I238222) );
nor I_13682 (I238333,I238268,I219752);
nand I_13683 (I238350,I238333,I219734);
nand I_13684 (I238367,I238350,I238302);
not I_13685 (I238384,I219752);
not I_13686 (I238401,I219749);
nor I_13687 (I238418,I238401,I219737);
and I_13688 (I238435,I238418,I219758);
or I_13689 (I238452,I238435,I219740);
DFFARX1 I_13690  ( .D(I238452), .CLK(I5694_clk), .RSTB(I238251_rst), .Q(I238469) );
nor I_13691 (I238486,I238469,I238350);
nand I_13692 (I238237,I238384,I238486);
not I_13693 (I238234,I238469);
and I_13694 (I238531,I238469,I238367);
DFFARX1 I_13695  ( .D(I238531), .CLK(I5694_clk), .RSTB(I238251_rst), .Q(I238219) );
DFFARX1 I_13696  ( .D(I238469), .CLK(I5694_clk), .RSTB(I238251_rst), .Q(I238562) );
and I_13697 (I238216,I238384,I238562);
nand I_13698 (I238593,I238268,I219749);
not I_13699 (I238610,I238593);
nor I_13700 (I238627,I238469,I238610);
DFFARX1 I_13701  ( .D(I219761), .CLK(I5694_clk), .RSTB(I238251_rst), .Q(I238644) );
nand I_13702 (I238661,I238644,I238593);
and I_13703 (I238678,I238384,I238661);
DFFARX1 I_13704  ( .D(I238678), .CLK(I5694_clk), .RSTB(I238251_rst), .Q(I238243) );
not I_13705 (I238709,I238644);
nand I_13706 (I238231,I238644,I238627);
nand I_13707 (I238225,I238644,I238610);
DFFARX1 I_13708  ( .D(I219743), .CLK(I5694_clk), .RSTB(I238251_rst), .Q(I238754) );
not I_13709 (I238771,I238754);
nor I_13710 (I238240,I238644,I238771);
nor I_13711 (I238802,I238771,I238709);
and I_13712 (I238819,I238350,I238802);
or I_13713 (I238836,I238593,I238819);
DFFARX1 I_13714  ( .D(I238836), .CLK(I5694_clk), .RSTB(I238251_rst), .Q(I238228) );
DFFARX1 I_13715  ( .D(I238771), .CLK(I5694_clk), .RSTB(I238251_rst), .Q(I238213) );
not I_13716 (I238914_rst,I5701);
not I_13717 (I238931,I224535);
nor I_13718 (I238948,I224514,I224526);
nand I_13719 (I238965,I238948,I224520);
DFFARX1 I_13720  ( .D(I238965), .CLK(I5694_clk), .RSTB(I238914_rst), .Q(I238885) );
nor I_13721 (I238996,I238931,I224514);
nand I_13722 (I239013,I238996,I224541);
nand I_13723 (I239030,I239013,I238965);
not I_13724 (I239047,I224514);
not I_13725 (I239064,I224517);
nor I_13726 (I239081,I239064,I224529);
and I_13727 (I239098,I239081,I224532);
or I_13728 (I239115,I239098,I224538);
DFFARX1 I_13729  ( .D(I239115), .CLK(I5694_clk), .RSTB(I238914_rst), .Q(I239132) );
nor I_13730 (I239149,I239132,I239013);
nand I_13731 (I238900,I239047,I239149);
not I_13732 (I238897,I239132);
and I_13733 (I239194,I239132,I239030);
DFFARX1 I_13734  ( .D(I239194), .CLK(I5694_clk), .RSTB(I238914_rst), .Q(I238882) );
DFFARX1 I_13735  ( .D(I239132), .CLK(I5694_clk), .RSTB(I238914_rst), .Q(I239225) );
and I_13736 (I238879,I239047,I239225);
nand I_13737 (I239256,I238931,I224517);
not I_13738 (I239273,I239256);
nor I_13739 (I239290,I239132,I239273);
DFFARX1 I_13740  ( .D(I224511), .CLK(I5694_clk), .RSTB(I238914_rst), .Q(I239307) );
nand I_13741 (I239324,I239307,I239256);
and I_13742 (I239341,I239047,I239324);
DFFARX1 I_13743  ( .D(I239341), .CLK(I5694_clk), .RSTB(I238914_rst), .Q(I238906) );
not I_13744 (I239372,I239307);
nand I_13745 (I238894,I239307,I239290);
nand I_13746 (I238888,I239307,I239273);
DFFARX1 I_13747  ( .D(I224523), .CLK(I5694_clk), .RSTB(I238914_rst), .Q(I239417) );
not I_13748 (I239434,I239417);
nor I_13749 (I238903,I239307,I239434);
nor I_13750 (I239465,I239434,I239372);
and I_13751 (I239482,I239013,I239465);
or I_13752 (I239499,I239256,I239482);
DFFARX1 I_13753  ( .D(I239499), .CLK(I5694_clk), .RSTB(I238914_rst), .Q(I238891) );
DFFARX1 I_13754  ( .D(I239434), .CLK(I5694_clk), .RSTB(I238914_rst), .Q(I238876) );
not I_13755 (I239577_rst,I5701);
not I_13756 (I239594,I180896);
nor I_13757 (I239611,I180878,I180872);
nand I_13758 (I239628,I239611,I180875);
DFFARX1 I_13759  ( .D(I239628), .CLK(I5694_clk), .RSTB(I239577_rst), .Q(I239548) );
nor I_13760 (I239659,I239594,I180878);
nand I_13761 (I239676,I239659,I180884);
nand I_13762 (I239693,I239676,I239628);
not I_13763 (I239710,I180878);
not I_13764 (I239727,I180893);
nor I_13765 (I239744,I239727,I180881);
and I_13766 (I239761,I239744,I180887);
or I_13767 (I239778,I239761,I180902);
DFFARX1 I_13768  ( .D(I239778), .CLK(I5694_clk), .RSTB(I239577_rst), .Q(I239795) );
nor I_13769 (I239812,I239795,I239676);
nand I_13770 (I239563,I239710,I239812);
not I_13771 (I239560,I239795);
and I_13772 (I239857,I239795,I239693);
DFFARX1 I_13773  ( .D(I239857), .CLK(I5694_clk), .RSTB(I239577_rst), .Q(I239545) );
DFFARX1 I_13774  ( .D(I239795), .CLK(I5694_clk), .RSTB(I239577_rst), .Q(I239888) );
and I_13775 (I239542,I239710,I239888);
nand I_13776 (I239919,I239594,I180893);
not I_13777 (I239936,I239919);
nor I_13778 (I239953,I239795,I239936);
DFFARX1 I_13779  ( .D(I180890), .CLK(I5694_clk), .RSTB(I239577_rst), .Q(I239970) );
nand I_13780 (I239987,I239970,I239919);
and I_13781 (I240004,I239710,I239987);
DFFARX1 I_13782  ( .D(I240004), .CLK(I5694_clk), .RSTB(I239577_rst), .Q(I239569) );
not I_13783 (I240035,I239970);
nand I_13784 (I239557,I239970,I239953);
nand I_13785 (I239551,I239970,I239936);
DFFARX1 I_13786  ( .D(I180899), .CLK(I5694_clk), .RSTB(I239577_rst), .Q(I240080) );
not I_13787 (I240097,I240080);
nor I_13788 (I239566,I239970,I240097);
nor I_13789 (I240128,I240097,I240035);
and I_13790 (I240145,I239676,I240128);
or I_13791 (I240162,I239919,I240145);
DFFARX1 I_13792  ( .D(I240162), .CLK(I5694_clk), .RSTB(I239577_rst), .Q(I239554) );
DFFARX1 I_13793  ( .D(I240097), .CLK(I5694_clk), .RSTB(I239577_rst), .Q(I239539) );
not I_13794 (I240240_rst,I5701);
or I_13795 (I240257,I199570,I199555);
or I_13796 (I240274,I199564,I199570);
DFFARX1 I_13797  ( .D(I240274), .CLK(I5694_clk), .RSTB(I240240_rst), .Q(I240214) );
nor I_13798 (I240305,I199576,I199585);
not I_13799 (I240322,I240305);
not I_13800 (I240339,I199576);
and I_13801 (I240356,I240339,I199573);
nor I_13802 (I240373,I240356,I199555);
nor I_13803 (I240390,I199582,I199558);
DFFARX1 I_13804  ( .D(I240390), .CLK(I5694_clk), .RSTB(I240240_rst), .Q(I240407) );
nand I_13805 (I240424,I240407,I240257);
and I_13806 (I240441,I240373,I240424);
DFFARX1 I_13807  ( .D(I240441), .CLK(I5694_clk), .RSTB(I240240_rst), .Q(I240208) );
nor I_13808 (I240472,I199582,I199564);
DFFARX1 I_13809  ( .D(I240472), .CLK(I5694_clk), .RSTB(I240240_rst), .Q(I240489) );
and I_13810 (I240205,I240305,I240489);
DFFARX1 I_13811  ( .D(I199567), .CLK(I5694_clk), .RSTB(I240240_rst), .Q(I240520) );
and I_13812 (I240537,I240520,I199561);
DFFARX1 I_13813  ( .D(I240537), .CLK(I5694_clk), .RSTB(I240240_rst), .Q(I240554) );
not I_13814 (I240217,I240554);
DFFARX1 I_13815  ( .D(I240537), .CLK(I5694_clk), .RSTB(I240240_rst), .Q(I240202) );
DFFARX1 I_13816  ( .D(I199579), .CLK(I5694_clk), .RSTB(I240240_rst), .Q(I240599) );
not I_13817 (I240616,I240599);
nor I_13818 (I240633,I240274,I240616);
and I_13819 (I240650,I240537,I240633);
or I_13820 (I240667,I240257,I240650);
DFFARX1 I_13821  ( .D(I240667), .CLK(I5694_clk), .RSTB(I240240_rst), .Q(I240223) );
nor I_13822 (I240698,I240599,I240407);
nand I_13823 (I240232,I240373,I240698);
nor I_13824 (I240729,I240599,I240322);
nand I_13825 (I240226,I240472,I240729);
not I_13826 (I240229,I240599);
nand I_13827 (I240220,I240599,I240322);
DFFARX1 I_13828  ( .D(I240599), .CLK(I5694_clk), .RSTB(I240240_rst), .Q(I240211) );
not I_13829 (I240835_rst,I5701);
or I_13830 (I240852,I227949,I227958);
or I_13831 (I240869,I227952,I227949);
DFFARX1 I_13832  ( .D(I240869), .CLK(I5694_clk), .RSTB(I240835_rst), .Q(I240809) );
nor I_13833 (I240900,I227928,I227931);
not I_13834 (I240917,I240900);
not I_13835 (I240934,I227928);
and I_13836 (I240951,I240934,I227940);
nor I_13837 (I240968,I240951,I227958);
nor I_13838 (I240985,I227946,I227937);
DFFARX1 I_13839  ( .D(I240985), .CLK(I5694_clk), .RSTB(I240835_rst), .Q(I241002) );
nand I_13840 (I241019,I241002,I240852);
and I_13841 (I241036,I240968,I241019);
DFFARX1 I_13842  ( .D(I241036), .CLK(I5694_clk), .RSTB(I240835_rst), .Q(I240803) );
nor I_13843 (I241067,I227946,I227952);
DFFARX1 I_13844  ( .D(I241067), .CLK(I5694_clk), .RSTB(I240835_rst), .Q(I241084) );
and I_13845 (I240800,I240900,I241084);
DFFARX1 I_13846  ( .D(I227943), .CLK(I5694_clk), .RSTB(I240835_rst), .Q(I241115) );
and I_13847 (I241132,I241115,I227934);
DFFARX1 I_13848  ( .D(I241132), .CLK(I5694_clk), .RSTB(I240835_rst), .Q(I241149) );
not I_13849 (I240812,I241149);
DFFARX1 I_13850  ( .D(I241132), .CLK(I5694_clk), .RSTB(I240835_rst), .Q(I240797) );
DFFARX1 I_13851  ( .D(I227955), .CLK(I5694_clk), .RSTB(I240835_rst), .Q(I241194) );
not I_13852 (I241211,I241194);
nor I_13853 (I241228,I240869,I241211);
and I_13854 (I241245,I241132,I241228);
or I_13855 (I241262,I240852,I241245);
DFFARX1 I_13856  ( .D(I241262), .CLK(I5694_clk), .RSTB(I240835_rst), .Q(I240818) );
nor I_13857 (I241293,I241194,I241002);
nand I_13858 (I240827,I240968,I241293);
nor I_13859 (I241324,I241194,I240917);
nand I_13860 (I240821,I241067,I241324);
not I_13861 (I240824,I241194);
nand I_13862 (I240815,I241194,I240917);
DFFARX1 I_13863  ( .D(I241194), .CLK(I5694_clk), .RSTB(I240835_rst), .Q(I240806) );
not I_13864 (I241430_rst,I5701);
or I_13865 (I241447,I184578,I184593);
or I_13866 (I241464,I184581,I184578);
DFFARX1 I_13867  ( .D(I241464), .CLK(I5694_clk), .RSTB(I241430_rst), .Q(I241404) );
nor I_13868 (I241495,I184584,I184599);
not I_13869 (I241512,I241495);
not I_13870 (I241529,I184584);
and I_13871 (I241546,I241529,I184587);
nor I_13872 (I241563,I241546,I184593);
nor I_13873 (I241580,I184590,I184608);
DFFARX1 I_13874  ( .D(I241580), .CLK(I5694_clk), .RSTB(I241430_rst), .Q(I241597) );
nand I_13875 (I241614,I241597,I241447);
and I_13876 (I241631,I241563,I241614);
DFFARX1 I_13877  ( .D(I241631), .CLK(I5694_clk), .RSTB(I241430_rst), .Q(I241398) );
nor I_13878 (I241662,I184590,I184581);
DFFARX1 I_13879  ( .D(I241662), .CLK(I5694_clk), .RSTB(I241430_rst), .Q(I241679) );
and I_13880 (I241395,I241495,I241679);
DFFARX1 I_13881  ( .D(I184605), .CLK(I5694_clk), .RSTB(I241430_rst), .Q(I241710) );
and I_13882 (I241727,I241710,I184596);
DFFARX1 I_13883  ( .D(I241727), .CLK(I5694_clk), .RSTB(I241430_rst), .Q(I241744) );
not I_13884 (I241407,I241744);
DFFARX1 I_13885  ( .D(I241727), .CLK(I5694_clk), .RSTB(I241430_rst), .Q(I241392) );
DFFARX1 I_13886  ( .D(I184602), .CLK(I5694_clk), .RSTB(I241430_rst), .Q(I241789) );
not I_13887 (I241806,I241789);
nor I_13888 (I241823,I241464,I241806);
and I_13889 (I241840,I241727,I241823);
or I_13890 (I241857,I241447,I241840);
DFFARX1 I_13891  ( .D(I241857), .CLK(I5694_clk), .RSTB(I241430_rst), .Q(I241413) );
nor I_13892 (I241888,I241789,I241597);
nand I_13893 (I241422,I241563,I241888);
nor I_13894 (I241919,I241789,I241512);
nand I_13895 (I241416,I241662,I241919);
not I_13896 (I241419,I241789);
nand I_13897 (I241410,I241789,I241512);
DFFARX1 I_13898  ( .D(I241789), .CLK(I5694_clk), .RSTB(I241430_rst), .Q(I241401) );
not I_13899 (I242025_rst,I5701);
or I_13900 (I24204_rst2,I192534,I192549);
or I_13901 (I242059,I192537,I192534);
DFFARX1 I_13902  ( .D(I242059), .CLK(I5694_clk), .RSTB(I242025_rst), .Q(I241999) );
nor I_13903 (I242090,I192540,I192555);
not I_13904 (I242107,I242090);
not I_13905 (I242124,I192540);
and I_13906 (I242141,I242124,I192543);
nor I_13907 (I242158,I242141,I192549);
nor I_13908 (I242175,I192546,I192564);
DFFARX1 I_13909  ( .D(I242175), .CLK(I5694_clk), .RSTB(I242025_rst), .Q(I242192) );
nand I_13910 (I242209,I242192,I24204_rst2);
and I_13911 (I242226,I242158,I242209);
DFFARX1 I_13912  ( .D(I242226), .CLK(I5694_clk), .RSTB(I242025_rst), .Q(I241993) );
nor I_13913 (I242257,I192546,I192537);
DFFARX1 I_13914  ( .D(I242257), .CLK(I5694_clk), .RSTB(I242025_rst), .Q(I242274) );
and I_13915 (I241990,I242090,I242274);
DFFARX1 I_13916  ( .D(I192561), .CLK(I5694_clk), .RSTB(I242025_rst), .Q(I242305) );
and I_13917 (I242322,I242305,I192552);
DFFARX1 I_13918  ( .D(I242322), .CLK(I5694_clk), .RSTB(I242025_rst), .Q(I242339) );
not I_13919 (I242002,I242339);
DFFARX1 I_13920  ( .D(I242322), .CLK(I5694_clk), .RSTB(I242025_rst), .Q(I241987) );
DFFARX1 I_13921  ( .D(I192558), .CLK(I5694_clk), .RSTB(I242025_rst), .Q(I242384) );
not I_13922 (I242401,I242384);
nor I_13923 (I242418,I242059,I242401);
and I_13924 (I242435,I242322,I242418);
or I_13925 (I242452,I24204_rst2,I242435);
DFFARX1 I_13926  ( .D(I242452), .CLK(I5694_clk), .RSTB(I242025_rst), .Q(I242008) );
nor I_13927 (I242483,I242384,I242192);
nand I_13928 (I242017,I242158,I242483);
nor I_13929 (I242514,I242384,I242107);
nand I_13930 (I242011,I242257,I242514);
not I_13931 (I242014,I242384);
nand I_13932 (I242005,I242384,I242107);
DFFARX1 I_13933  ( .D(I242384), .CLK(I5694_clk), .RSTB(I242025_rst), .Q(I241996) );
not I_13934 (I242620_rst,I5701);
or I_13935 (I242637,I211903,I211915);
not I_13936 (I242603,I242637);
DFFARX1 I_13937  ( .D(I242637), .CLK(I5694_clk), .RSTB(I242620_rst), .Q(I242582) );
or I_13938 (I242682,I211927,I211903);
nor I_13939 (I242699,I211921,I211906);
nor I_13940 (I242716,I242699,I242637);
not I_13941 (I242733,I211921);
and I_13942 (I242750,I242733,I211918);
nor I_13943 (I242767,I242750,I211915);
DFFARX1 I_13944  ( .D(I242767), .CLK(I5694_clk), .RSTB(I242620_rst), .Q(I242784) );
nor I_13945 (I242801,I211912,I211909);
DFFARX1 I_13946  ( .D(I242801), .CLK(I5694_clk), .RSTB(I242620_rst), .Q(I242818) );
nor I_13947 (I242609,I242818,I242767);
not I_13948 (I242849,I242818);
nor I_13949 (I242866,I211912,I211927);
nand I_13950 (I242883,I242767,I242866);
and I_13951 (I242900,I242682,I242883);
DFFARX1 I_13952  ( .D(I242900), .CLK(I5694_clk), .RSTB(I242620_rst), .Q(I242612) );
DFFARX1 I_13953  ( .D(I211924), .CLK(I5694_clk), .RSTB(I242620_rst), .Q(I242931) );
and I_13954 (I242948,I242931,I211897);
nor I_13955 (I242965,I242948,I242849);
and I_13956 (I242982,I242866,I242965);
or I_13957 (I242999,I242699,I242982);
DFFARX1 I_13958  ( .D(I242999), .CLK(I5694_clk), .RSTB(I242620_rst), .Q(I242597) );
not I_13959 (I243030,I242948);
nor I_13960 (I243047,I242637,I243030);
nand I_13961 (I242600,I242682,I243047);
nand I_13962 (I242594,I242818,I243030);
DFFARX1 I_13963  ( .D(I242948), .CLK(I5694_clk), .RSTB(I242620_rst), .Q(I242588) );
DFFARX1 I_13964  ( .D(I211900), .CLK(I5694_clk), .RSTB(I242620_rst), .Q(I243106) );
nand I_13965 (I242606,I243106,I242716);
DFFARX1 I_13966  ( .D(I243106), .CLK(I5694_clk), .RSTB(I242620_rst), .Q(I243137) );
not I_13967 (I242591,I243137);
and I_13968 (I242585,I243106,I242784);
not I_13969 (I243215_rst,I5701);
or I_13970 (I243232,I204213,I204243);
not I_13971 (I243198,I243232);
DFFARX1 I_13972  ( .D(I243232), .CLK(I5694_clk), .RSTB(I243215_rst), .Q(I243177) );
or I_13973 (I243277,I204222,I204213);
nor I_13974 (I243294,I204228,I204225);
nor I_13975 (I243311,I243294,I243232);
not I_13976 (I243328,I204228);
and I_13977 (I243345,I243328,I204234);
nor I_13978 (I243362,I243345,I204243);
DFFARX1 I_13979  ( .D(I243362), .CLK(I5694_clk), .RSTB(I243215_rst), .Q(I243379) );
nor I_13980 (I243396,I204219,I204237);
DFFARX1 I_13981  ( .D(I243396), .CLK(I5694_clk), .RSTB(I243215_rst), .Q(I243413) );
nor I_13982 (I243204,I243413,I243362);
not I_13983 (I243444,I243413);
nor I_13984 (I243461,I204219,I204222);
nand I_13985 (I243478,I243362,I243461);
and I_13986 (I243495,I243277,I243478);
DFFARX1 I_13987  ( .D(I243495), .CLK(I5694_clk), .RSTB(I243215_rst), .Q(I243207) );
DFFARX1 I_13988  ( .D(I204240), .CLK(I5694_clk), .RSTB(I243215_rst), .Q(I243526) );
and I_13989 (I243543,I243526,I204231);
nor I_13990 (I243560,I243543,I243444);
and I_13991 (I243577,I243461,I243560);
or I_13992 (I243594,I243294,I243577);
DFFARX1 I_13993  ( .D(I243594), .CLK(I5694_clk), .RSTB(I243215_rst), .Q(I243192) );
not I_13994 (I243625,I243543);
nor I_13995 (I243642,I243232,I243625);
nand I_13996 (I243195,I243277,I243642);
nand I_13997 (I243189,I243413,I243625);
DFFARX1 I_13998  ( .D(I243543), .CLK(I5694_clk), .RSTB(I243215_rst), .Q(I243183) );
DFFARX1 I_13999  ( .D(I204216), .CLK(I5694_clk), .RSTB(I243215_rst), .Q(I243701) );
nand I_14000 (I243201,I243701,I243311);
DFFARX1 I_14001  ( .D(I243701), .CLK(I5694_clk), .RSTB(I243215_rst), .Q(I243732) );
not I_14002 (I243186,I243732);
and I_14003 (I243180,I243701,I243379);
not I_14004 (I243810_rst,I5701);
not I_14005 (I243827,I218482);
nor I_14006 (I243844,I218500,I218491);
nand I_14007 (I243861,I243844,I218497);
nor I_14008 (I243878,I243827,I218500);
nand I_14009 (I243895,I243878,I218503);
not I_14010 (I243912,I243895);
not I_14011 (I243929,I218500);
nor I_14012 (I243799,I243895,I243929);
not I_14013 (I243960,I243929);
nand I_14014 (I243784,I243895,I243960);
not I_14015 (I243991,I218479);
nor I_14016 (I244008,I243991,I218494);
and I_14017 (I244025,I244008,I218476);
or I_14018 (I244042,I244025,I218485);
DFFARX1 I_14019  ( .D(I244042), .CLK(I5694_clk), .RSTB(I243810_rst), .Q(I244059) );
nor I_14020 (I244076,I244059,I243912);
DFFARX1 I_14021  ( .D(I244059), .CLK(I5694_clk), .RSTB(I243810_rst), .Q(I244093) );
not I_14022 (I243781,I244093);
nand I_14023 (I244124,I243827,I218479);
and I_14024 (I244141,I244124,I244076);
DFFARX1 I_14025  ( .D(I244124), .CLK(I5694_clk), .RSTB(I243810_rst), .Q(I243778) );
DFFARX1 I_14026  ( .D(I218488), .CLK(I5694_clk), .RSTB(I243810_rst), .Q(I244172) );
nor I_14027 (I244189,I244172,I243895);
nand I_14028 (I243796,I244059,I244189);
nor I_14029 (I244220,I244172,I243960);
not I_14030 (I243793,I244172);
nand I_14031 (I244251,I244172,I243861);
and I_14032 (I244268,I243929,I244251);
DFFARX1 I_14033  ( .D(I244268), .CLK(I5694_clk), .RSTB(I243810_rst), .Q(I243772) );
DFFARX1 I_14034  ( .D(I244172), .CLK(I5694_clk), .RSTB(I243810_rst), .Q(I243775) );
DFFARX1 I_14035  ( .D(I218506), .CLK(I5694_clk), .RSTB(I243810_rst), .Q(I244313) );
not I_14036 (I244330,I244313);
nand I_14037 (I244347,I244330,I243895);
and I_14038 (I244364,I244124,I244347);
DFFARX1 I_14039  ( .D(I244364), .CLK(I5694_clk), .RSTB(I243810_rst), .Q(I243802) );
or I_14040 (I244395,I244330,I244141);
DFFARX1 I_14041  ( .D(I244395), .CLK(I5694_clk), .RSTB(I243810_rst), .Q(I243787) );
nand I_14042 (I243790,I244330,I244220);
not I_14043 (I244473_rst,I5701);
not I_14044 (I244490,I223367);
nor I_14045 (I244507,I223358,I223364);
nand I_14046 (I244524,I244507,I223376);
nor I_14047 (I244541,I244490,I223358);
nand I_14048 (I244558,I244541,I223361);
not I_14049 (I244575,I244558);
not I_14050 (I244592,I223358);
nor I_14051 (I244462,I244558,I244592);
not I_14052 (I244623,I244592);
nand I_14053 (I244447,I244558,I244623);
not I_14054 (I244654,I223385);
nor I_14055 (I244671,I244654,I223379);
and I_14056 (I244688,I244671,I223370);
or I_14057 (I244705,I244688,I223355);
DFFARX1 I_14058  ( .D(I244705), .CLK(I5694_clk), .RSTB(I244473_rst), .Q(I244722) );
nor I_14059 (I244739,I244722,I244575);
DFFARX1 I_14060  ( .D(I244722), .CLK(I5694_clk), .RSTB(I244473_rst), .Q(I244756) );
not I_14061 (I244444,I244756);
nand I_14062 (I244787,I244490,I223385);
and I_14063 (I244804,I244787,I244739);
DFFARX1 I_14064  ( .D(I244787), .CLK(I5694_clk), .RSTB(I244473_rst), .Q(I244441) );
DFFARX1 I_14065  ( .D(I223373), .CLK(I5694_clk), .RSTB(I244473_rst), .Q(I244835) );
nor I_14066 (I244852,I244835,I244558);
nand I_14067 (I244459,I244722,I244852);
nor I_14068 (I244883,I244835,I244623);
not I_14069 (I244456,I244835);
nand I_14070 (I244914,I244835,I244524);
and I_14071 (I244931,I244592,I244914);
DFFARX1 I_14072  ( .D(I244931), .CLK(I5694_clk), .RSTB(I244473_rst), .Q(I244435) );
DFFARX1 I_14073  ( .D(I244835), .CLK(I5694_clk), .RSTB(I244473_rst), .Q(I244438) );
DFFARX1 I_14074  ( .D(I223382), .CLK(I5694_clk), .RSTB(I244473_rst), .Q(I244976) );
not I_14075 (I244993,I244976);
nand I_14076 (I245010,I244993,I244558);
and I_14077 (I245027,I244787,I245010);
DFFARX1 I_14078  ( .D(I245027), .CLK(I5694_clk), .RSTB(I244473_rst), .Q(I244465) );
or I_14079 (I245058,I244993,I244804);
DFFARX1 I_14080  ( .D(I245058), .CLK(I5694_clk), .RSTB(I244473_rst), .Q(I244450) );
nand I_14081 (I244453,I244993,I244883);
not I_14082 (I245136_rst,I5701);
not I_14083 (I245153,I236890);
nor I_14084 (I245170,I236896,I236902);
nand I_14085 (I245187,I245170,I236905);
nor I_14086 (I245204,I245153,I236896);
nand I_14087 (I245221,I245204,I236887);
not I_14088 (I245238,I245221);
not I_14089 (I245255,I236896);
nor I_14090 (I245125,I245221,I245255);
not I_14091 (I245286,I245255);
nand I_14092 (I245110,I245221,I245286);
not I_14093 (I245317,I236899);
nor I_14094 (I245334,I245317,I236893);
and I_14095 (I245351,I245334,I236908);
or I_14096 (I245368,I245351,I236914);
DFFARX1 I_14097  ( .D(I245368), .CLK(I5694_clk), .RSTB(I245136_rst), .Q(I245385) );
nor I_14098 (I245402,I245385,I245238);
DFFARX1 I_14099  ( .D(I245385), .CLK(I5694_clk), .RSTB(I245136_rst), .Q(I245419) );
not I_14100 (I245107,I245419);
nand I_14101 (I245450,I245153,I236899);
and I_14102 (I245467,I245450,I245402);
DFFARX1 I_14103  ( .D(I245450), .CLK(I5694_clk), .RSTB(I245136_rst), .Q(I245104) );
DFFARX1 I_14104  ( .D(I236911), .CLK(I5694_clk), .RSTB(I245136_rst), .Q(I245498) );
nor I_14105 (I245515,I245498,I245221);
nand I_14106 (I245122,I245385,I245515);
nor I_14107 (I245546,I245498,I245286);
not I_14108 (I245119,I245498);
nand I_14109 (I245577,I245498,I245187);
and I_14110 (I245594,I245255,I245577);
DFFARX1 I_14111  ( .D(I245594), .CLK(I5694_clk), .RSTB(I245136_rst), .Q(I245098) );
DFFARX1 I_14112  ( .D(I245498), .CLK(I5694_clk), .RSTB(I245136_rst), .Q(I245101) );
DFFARX1 I_14113  ( .D(I236917), .CLK(I5694_clk), .RSTB(I245136_rst), .Q(I245639) );
not I_14114 (I245656,I245639);
nand I_14115 (I245673,I245656,I245221);
and I_14116 (I245690,I245450,I245673);
DFFARX1 I_14117  ( .D(I245690), .CLK(I5694_clk), .RSTB(I245136_rst), .Q(I245128) );
or I_14118 (I245721,I245656,I245467);
DFFARX1 I_14119  ( .D(I245721), .CLK(I5694_clk), .RSTB(I245136_rst), .Q(I245113) );
nand I_14120 (I245116,I245656,I245546);
not I_14121 (I245799_rst,I5701);
not I_14122 (I245816,I217270);
nor I_14123 (I245833,I217267,I217258);
nand I_14124 (I245850,I245833,I217261);
nor I_14125 (I245867,I245816,I217267);
nand I_14126 (I245884,I245867,I217255);
not I_14127 (I245901,I245884);
not I_14128 (I245918,I217267);
nor I_14129 (I245788,I245884,I245918);
not I_14130 (I245949,I245918);
nand I_14131 (I245773,I245884,I245949);
not I_14132 (I245980,I217276);
nor I_14133 (I245997,I245980,I217279);
and I_14134 (I246014,I245997,I217264);
or I_14135 (I246031,I246014,I217252);
DFFARX1 I_14136  ( .D(I246031), .CLK(I5694_clk), .RSTB(I245799_rst), .Q(I246048) );
nor I_14137 (I246065,I246048,I245901);
DFFARX1 I_14138  ( .D(I246048), .CLK(I5694_clk), .RSTB(I245799_rst), .Q(I246082) );
not I_14139 (I245770,I246082);
nand I_14140 (I246113,I245816,I217276);
and I_14141 (I246130,I246113,I246065);
DFFARX1 I_14142  ( .D(I246113), .CLK(I5694_clk), .RSTB(I245799_rst), .Q(I245767) );
DFFARX1 I_14143  ( .D(I217273), .CLK(I5694_clk), .RSTB(I245799_rst), .Q(I246161) );
nor I_14144 (I246178,I246161,I245884);
nand I_14145 (I245785,I246048,I246178);
nor I_14146 (I246209,I246161,I245949);
not I_14147 (I245782,I246161);
nand I_14148 (I246240,I246161,I245850);
and I_14149 (I246257,I245918,I246240);
DFFARX1 I_14150  ( .D(I246257), .CLK(I5694_clk), .RSTB(I245799_rst), .Q(I245761) );
DFFARX1 I_14151  ( .D(I246161), .CLK(I5694_clk), .RSTB(I245799_rst), .Q(I245764) );
DFFARX1 I_14152  ( .D(I217282), .CLK(I5694_clk), .RSTB(I245799_rst), .Q(I246302) );
not I_14153 (I246319,I246302);
nand I_14154 (I246336,I246319,I245884);
and I_14155 (I246353,I246113,I246336);
DFFARX1 I_14156  ( .D(I246353), .CLK(I5694_clk), .RSTB(I245799_rst), .Q(I245791) );
or I_14157 (I246384,I246319,I246130);
DFFARX1 I_14158  ( .D(I246384), .CLK(I5694_clk), .RSTB(I245799_rst), .Q(I245776) );
nand I_14159 (I245779,I246319,I246209);
not I_14160 (I246462_rst,I5701);
not I_14161 (I246479,I198949);
nor I_14162 (I246496,I198952,I198958);
nand I_14163 (I246513,I246496,I198964);
nor I_14164 (I246530,I246479,I198952);
nand I_14165 (I246547,I246530,I198943);
not I_14166 (I246564,I246547);
not I_14167 (I246581,I198952);
nor I_14168 (I246451,I246547,I246581);
not I_14169 (I246612,I246581);
nand I_14170 (I246436,I246547,I246612);
not I_14171 (I246643,I198955);
nor I_14172 (I246660,I246643,I198970);
and I_14173 (I246677,I246660,I198973);
or I_14174 (I246694,I246677,I198946);
DFFARX1 I_14175  ( .D(I246694), .CLK(I5694_clk), .RSTB(I246462_rst), .Q(I246711) );
nor I_14176 (I246728,I246711,I246564);
DFFARX1 I_14177  ( .D(I246711), .CLK(I5694_clk), .RSTB(I246462_rst), .Q(I246745) );
not I_14178 (I246433,I246745);
nand I_14179 (I246776,I246479,I198955);
and I_14180 (I246793,I246776,I246728);
DFFARX1 I_14181  ( .D(I246776), .CLK(I5694_clk), .RSTB(I246462_rst), .Q(I246430) );
DFFARX1 I_14182  ( .D(I198967), .CLK(I5694_clk), .RSTB(I246462_rst), .Q(I246824) );
nor I_14183 (I246841,I246824,I246547);
nand I_14184 (I246448,I246711,I246841);
nor I_14185 (I246872,I246824,I246612);
not I_14186 (I246445,I246824);
nand I_14187 (I246903,I246824,I246513);
and I_14188 (I246920,I246581,I246903);
DFFARX1 I_14189  ( .D(I246920), .CLK(I5694_clk), .RSTB(I246462_rst), .Q(I246424) );
DFFARX1 I_14190  ( .D(I246824), .CLK(I5694_clk), .RSTB(I246462_rst), .Q(I246427) );
DFFARX1 I_14191  ( .D(I198961), .CLK(I5694_clk), .RSTB(I246462_rst), .Q(I246965) );
not I_14192 (I246982,I246965);
nand I_14193 (I246999,I246982,I246547);
and I_14194 (I247016,I246776,I246999);
DFFARX1 I_14195  ( .D(I247016), .CLK(I5694_clk), .RSTB(I246462_rst), .Q(I246454) );
or I_14196 (I247047,I246982,I246793);
DFFARX1 I_14197  ( .D(I247047), .CLK(I5694_clk), .RSTB(I246462_rst), .Q(I246439) );
nand I_14198 (I246442,I246982,I246872);
not I_14199 (I247125_rst,I5701);
not I_14200 (I247142,I202494);
nor I_14201 (I247159,I202506,I202488);
nand I_14202 (I247176,I247159,I202509);
nor I_14203 (I247193,I247142,I202506);
nand I_14204 (I247210,I247193,I202500);
not I_14205 (I247227,I247210);
not I_14206 (I247244,I202506);
nor I_14207 (I247114,I247210,I247244);
not I_14208 (I247275,I247244);
nand I_14209 (I247099,I247210,I247275);
not I_14210 (I247306,I202491);
nor I_14211 (I247323,I247306,I202485);
and I_14212 (I247340,I247323,I202497);
or I_14213 (I247357,I247340,I202482);
DFFARX1 I_14214  ( .D(I247357), .CLK(I5694_clk), .RSTB(I247125_rst), .Q(I247374) );
nor I_14215 (I247391,I247374,I247227);
DFFARX1 I_14216  ( .D(I247374), .CLK(I5694_clk), .RSTB(I247125_rst), .Q(I247408) );
not I_14217 (I247096,I247408);
nand I_14218 (I247439,I247142,I202491);
and I_14219 (I247456,I247439,I247391);
DFFARX1 I_14220  ( .D(I247439), .CLK(I5694_clk), .RSTB(I247125_rst), .Q(I247093) );
DFFARX1 I_14221  ( .D(I202479), .CLK(I5694_clk), .RSTB(I247125_rst), .Q(I247487) );
nor I_14222 (I247504,I247487,I247210);
nand I_14223 (I247111,I247374,I247504);
nor I_14224 (I247535,I247487,I247275);
not I_14225 (I247108,I247487);
nand I_14226 (I247566,I247487,I247176);
and I_14227 (I247583,I247244,I247566);
DFFARX1 I_14228  ( .D(I247583), .CLK(I5694_clk), .RSTB(I247125_rst), .Q(I247087) );
DFFARX1 I_14229  ( .D(I247487), .CLK(I5694_clk), .RSTB(I247125_rst), .Q(I247090) );
DFFARX1 I_14230  ( .D(I202503), .CLK(I5694_clk), .RSTB(I247125_rst), .Q(I247628) );
not I_14231 (I247645,I247628);
nand I_14232 (I247662,I247645,I247210);
and I_14233 (I247679,I247439,I247662);
DFFARX1 I_14234  ( .D(I247679), .CLK(I5694_clk), .RSTB(I247125_rst), .Q(I247117) );
or I_14235 (I247710,I247645,I247456);
DFFARX1 I_14236  ( .D(I247710), .CLK(I5694_clk), .RSTB(I247125_rst), .Q(I247102) );
nand I_14237 (I247105,I247645,I247535);
not I_14238 (I247788_rst,I5701);
not I_14239 (I247805,I229787);
nor I_14240 (I24782_rst2,I229784,I229808);
nand I_14241 (I247839,I24782_rst2,I229805);
nor I_14242 (I247856,I247805,I229784);
nand I_14243 (I247873,I247856,I229811);
not I_14244 (I247890,I247873);
not I_14245 (I247907,I229784);
nor I_14246 (I247777,I247873,I247907);
not I_14247 (I247938,I247907);
nand I_14248 (I247762,I247873,I247938);
not I_14249 (I247969,I229802);
nor I_14250 (I247986,I247969,I229793);
and I_14251 (I248003,I247986,I229790);
or I_14252 (I248020,I248003,I229799);
DFFARX1 I_14253  ( .D(I248020), .CLK(I5694_clk), .RSTB(I247788_rst), .Q(I248037) );
nor I_14254 (I248054,I248037,I247890);
DFFARX1 I_14255  ( .D(I248037), .CLK(I5694_clk), .RSTB(I247788_rst), .Q(I248071) );
not I_14256 (I247759,I248071);
nand I_14257 (I248102,I247805,I229802);
and I_14258 (I248119,I248102,I248054);
DFFARX1 I_14259  ( .D(I248102), .CLK(I5694_clk), .RSTB(I247788_rst), .Q(I247756) );
DFFARX1 I_14260  ( .D(I229781), .CLK(I5694_clk), .RSTB(I247788_rst), .Q(I248150) );
nor I_14261 (I248167,I248150,I247873);
nand I_14262 (I247774,I248037,I248167);
nor I_14263 (I248198,I248150,I247938);
not I_14264 (I247771,I248150);
nand I_14265 (I248229,I248150,I247839);
and I_14266 (I248246,I247907,I248229);
DFFARX1 I_14267  ( .D(I248246), .CLK(I5694_clk), .RSTB(I247788_rst), .Q(I247750) );
DFFARX1 I_14268  ( .D(I248150), .CLK(I5694_clk), .RSTB(I247788_rst), .Q(I247753) );
DFFARX1 I_14269  ( .D(I229796), .CLK(I5694_clk), .RSTB(I247788_rst), .Q(I248291) );
not I_14270 (I248308,I248291);
nand I_14271 (I248325,I248308,I247873);
and I_14272 (I248342,I248102,I248325);
DFFARX1 I_14273  ( .D(I248342), .CLK(I5694_clk), .RSTB(I247788_rst), .Q(I247780) );
or I_14274 (I248373,I248308,I248119);
DFFARX1 I_14275  ( .D(I248373), .CLK(I5694_clk), .RSTB(I247788_rst), .Q(I247765) );
nand I_14276 (I247768,I248308,I248198);
not I_14277 (I248451_rst,I5701);
not I_14278 (I248468,I205384);
nor I_14279 (I248485,I205396,I205378);
nand I_14280 (I248502,I248485,I205399);
nor I_14281 (I248519,I248468,I205396);
nand I_14282 (I248536,I248519,I205390);
not I_14283 (I248553,I248536);
not I_14284 (I248570,I205396);
nor I_14285 (I248440,I248536,I248570);
not I_14286 (I248601,I248570);
nand I_14287 (I248425,I248536,I248601);
not I_14288 (I248632,I205381);
nor I_14289 (I248649,I248632,I205375);
and I_14290 (I248666,I248649,I205387);
or I_14291 (I248683,I248666,I205372);
DFFARX1 I_14292  ( .D(I248683), .CLK(I5694_clk), .RSTB(I248451_rst), .Q(I248700) );
nor I_14293 (I248717,I248700,I248553);
DFFARX1 I_14294  ( .D(I248700), .CLK(I5694_clk), .RSTB(I248451_rst), .Q(I248734) );
not I_14295 (I248422,I248734);
nand I_14296 (I248765,I248468,I205381);
and I_14297 (I248782,I248765,I248717);
DFFARX1 I_14298  ( .D(I248765), .CLK(I5694_clk), .RSTB(I248451_rst), .Q(I248419) );
DFFARX1 I_14299  ( .D(I205369), .CLK(I5694_clk), .RSTB(I248451_rst), .Q(I248813) );
nor I_14300 (I248830,I248813,I248536);
nand I_14301 (I248437,I248700,I248830);
nor I_14302 (I248861,I248813,I248601);
not I_14303 (I248434,I248813);
nand I_14304 (I248892,I248813,I248502);
and I_14305 (I248909,I248570,I248892);
DFFARX1 I_14306  ( .D(I248909), .CLK(I5694_clk), .RSTB(I248451_rst), .Q(I248413) );
DFFARX1 I_14307  ( .D(I248813), .CLK(I5694_clk), .RSTB(I248451_rst), .Q(I248416) );
DFFARX1 I_14308  ( .D(I205393), .CLK(I5694_clk), .RSTB(I248451_rst), .Q(I248954) );
not I_14309 (I248971,I248954);
nand I_14310 (I248988,I248971,I248536);
and I_14311 (I249005,I248765,I248988);
DFFARX1 I_14312  ( .D(I249005), .CLK(I5694_clk), .RSTB(I248451_rst), .Q(I248443) );
or I_14313 (I249036,I248971,I248782);
DFFARX1 I_14314  ( .D(I249036), .CLK(I5694_clk), .RSTB(I248451_rst), .Q(I248428) );
nand I_14315 (I248431,I248971,I248861);
not I_14316 (I249114_rst,I5701);
not I_14317 (I249131,I220998);
nor I_14318 (I249148,I221016,I221007);
nand I_14319 (I249165,I249148,I221013);
nor I_14320 (I249182,I249131,I221016);
nand I_14321 (I249199,I249182,I221019);
not I_14322 (I249216,I249199);
not I_14323 (I249233,I221016);
nor I_14324 (I249103,I249199,I249233);
not I_14325 (I249264,I249233);
nand I_14326 (I249088,I249199,I249264);
not I_14327 (I249295,I220995);
nor I_14328 (I249312,I249295,I221010);
and I_14329 (I249329,I249312,I220992);
or I_14330 (I249346,I249329,I221001);
DFFARX1 I_14331  ( .D(I249346), .CLK(I5694_clk), .RSTB(I249114_rst), .Q(I249363) );
nor I_14332 (I249380,I249363,I249216);
DFFARX1 I_14333  ( .D(I249363), .CLK(I5694_clk), .RSTB(I249114_rst), .Q(I249397) );
not I_14334 (I249085,I249397);
nand I_14335 (I249428,I249131,I220995);
and I_14336 (I249445,I249428,I249380);
DFFARX1 I_14337  ( .D(I249428), .CLK(I5694_clk), .RSTB(I249114_rst), .Q(I249082) );
DFFARX1 I_14338  ( .D(I221004), .CLK(I5694_clk), .RSTB(I249114_rst), .Q(I249476) );
nor I_14339 (I249493,I249476,I249199);
nand I_14340 (I249100,I249363,I249493);
nor I_14341 (I249524,I249476,I249264);
not I_14342 (I249097,I249476);
nand I_14343 (I249555,I249476,I249165);
and I_14344 (I249572,I249233,I249555);
DFFARX1 I_14345  ( .D(I249572), .CLK(I5694_clk), .RSTB(I249114_rst), .Q(I249076) );
DFFARX1 I_14346  ( .D(I249476), .CLK(I5694_clk), .RSTB(I249114_rst), .Q(I249079) );
DFFARX1 I_14347  ( .D(I221022), .CLK(I5694_clk), .RSTB(I249114_rst), .Q(I249617) );
not I_14348 (I249634,I249617);
nand I_14349 (I249651,I249634,I249199);
and I_14350 (I249668,I249428,I249651);
DFFARX1 I_14351  ( .D(I249668), .CLK(I5694_clk), .RSTB(I249114_rst), .Q(I249106) );
or I_14352 (I249699,I249634,I249445);
DFFARX1 I_14353  ( .D(I249699), .CLK(I5694_clk), .RSTB(I249114_rst), .Q(I249091) );
nand I_14354 (I249094,I249634,I249524);
not I_14355 (I249777_rst,I5701);
not I_14356 (I249794,I201338);
nor I_14357 (I249811,I201350,I201332);
nand I_14358 (I249828,I249811,I201353);
nor I_14359 (I249845,I249794,I201350);
nand I_14360 (I249862,I249845,I201344);
not I_14361 (I249879,I249862);
not I_14362 (I249896,I201350);
nor I_14363 (I249766,I249862,I249896);
not I_14364 (I249927,I249896);
nand I_14365 (I249751,I249862,I249927);
not I_14366 (I249958,I201335);
nor I_14367 (I249975,I249958,I201329);
and I_14368 (I249992,I249975,I201341);
or I_14369 (I250009,I249992,I201326);
DFFARX1 I_14370  ( .D(I250009), .CLK(I5694_clk), .RSTB(I249777_rst), .Q(I250026) );
nor I_14371 (I250043,I250026,I249879);
DFFARX1 I_14372  ( .D(I250026), .CLK(I5694_clk), .RSTB(I249777_rst), .Q(I250060) );
not I_14373 (I249748,I250060);
nand I_14374 (I250091,I249794,I201335);
and I_14375 (I250108,I250091,I250043);
DFFARX1 I_14376  ( .D(I250091), .CLK(I5694_clk), .RSTB(I249777_rst), .Q(I249745) );
DFFARX1 I_14377  ( .D(I201323), .CLK(I5694_clk), .RSTB(I249777_rst), .Q(I250139) );
nor I_14378 (I250156,I250139,I249862);
nand I_14379 (I249763,I250026,I250156);
nor I_14380 (I250187,I250139,I249927);
not I_14381 (I249760,I250139);
nand I_14382 (I250218,I250139,I249828);
and I_14383 (I250235,I249896,I250218);
DFFARX1 I_14384  ( .D(I250235), .CLK(I5694_clk), .RSTB(I249777_rst), .Q(I249739) );
DFFARX1 I_14385  ( .D(I250139), .CLK(I5694_clk), .RSTB(I249777_rst), .Q(I249742) );
DFFARX1 I_14386  ( .D(I201347), .CLK(I5694_clk), .RSTB(I249777_rst), .Q(I250280) );
not I_14387 (I250297,I250280);
nand I_14388 (I250314,I250297,I249862);
and I_14389 (I250331,I250091,I250314);
DFFARX1 I_14390  ( .D(I250331), .CLK(I5694_clk), .RSTB(I249777_rst), .Q(I249769) );
or I_14391 (I250362,I250297,I250108);
DFFARX1 I_14392  ( .D(I250362), .CLK(I5694_clk), .RSTB(I249777_rst), .Q(I249754) );
nand I_14393 (I249757,I250297,I250187);
not I_14394 (I250440_rst,I5701);
not I_14395 (I250457,I220369);
nor I_14396 (I250474,I220387,I220378);
nand I_14397 (I250491,I250474,I220384);
nor I_14398 (I250508,I250457,I220387);
nand I_14399 (I250525,I250508,I220390);
not I_14400 (I250542,I250525);
not I_14401 (I250559,I220387);
nor I_14402 (I250429,I250525,I250559);
not I_14403 (I250590,I250559);
nand I_14404 (I250414,I250525,I250590);
not I_14405 (I250621,I220366);
nor I_14406 (I250638,I250621,I220381);
and I_14407 (I250655,I250638,I220363);
or I_14408 (I250672,I250655,I220372);
DFFARX1 I_14409  ( .D(I250672), .CLK(I5694_clk), .RSTB(I250440_rst), .Q(I250689) );
nor I_14410 (I250706,I250689,I250542);
DFFARX1 I_14411  ( .D(I250689), .CLK(I5694_clk), .RSTB(I250440_rst), .Q(I250723) );
not I_14412 (I250411,I250723);
nand I_14413 (I250754,I250457,I220366);
and I_14414 (I250771,I250754,I250706);
DFFARX1 I_14415  ( .D(I250754), .CLK(I5694_clk), .RSTB(I250440_rst), .Q(I250408) );
DFFARX1 I_14416  ( .D(I220375), .CLK(I5694_clk), .RSTB(I250440_rst), .Q(I250802) );
nor I_14417 (I250819,I250802,I250525);
nand I_14418 (I250426,I250689,I250819);
nor I_14419 (I250850,I250802,I250590);
not I_14420 (I250423,I250802);
nand I_14421 (I250881,I250802,I250491);
and I_14422 (I250898,I250559,I250881);
DFFARX1 I_14423  ( .D(I250898), .CLK(I5694_clk), .RSTB(I250440_rst), .Q(I250402) );
DFFARX1 I_14424  ( .D(I250802), .CLK(I5694_clk), .RSTB(I250440_rst), .Q(I250405) );
DFFARX1 I_14425  ( .D(I220393), .CLK(I5694_clk), .RSTB(I250440_rst), .Q(I250943) );
not I_14426 (I250960,I250943);
nand I_14427 (I250977,I250960,I250525);
and I_14428 (I250994,I250754,I250977);
DFFARX1 I_14429  ( .D(I250994), .CLK(I5694_clk), .RSTB(I250440_rst), .Q(I250432) );
or I_14430 (I251025,I250960,I250771);
DFFARX1 I_14431  ( .D(I251025), .CLK(I5694_clk), .RSTB(I250440_rst), .Q(I250417) );
nand I_14432 (I250420,I250960,I250850);
not I_14433 (I251103_rst,I5701);
not I_14434 (I251120,I225101);
nor I_14435 (I251137,I225092,I225098);
nand I_14436 (I251154,I251137,I225110);
nor I_14437 (I251171,I251120,I225092);
nand I_14438 (I251188,I251171,I225095);
not I_14439 (I251205,I251188);
not I_14440 (I251222,I225092);
nor I_14441 (I251092,I251188,I251222);
not I_14442 (I251253,I251222);
nand I_14443 (I251077,I251188,I251253);
not I_14444 (I251284,I225119);
nor I_14445 (I251301,I251284,I225113);
and I_14446 (I251318,I251301,I225104);
or I_14447 (I251335,I251318,I225089);
DFFARX1 I_14448  ( .D(I251335), .CLK(I5694_clk), .RSTB(I251103_rst), .Q(I251352) );
nor I_14449 (I251369,I251352,I251205);
DFFARX1 I_14450  ( .D(I251352), .CLK(I5694_clk), .RSTB(I251103_rst), .Q(I251386) );
not I_14451 (I251074,I251386);
nand I_14452 (I251417,I251120,I225119);
and I_14453 (I251434,I251417,I251369);
DFFARX1 I_14454  ( .D(I251417), .CLK(I5694_clk), .RSTB(I251103_rst), .Q(I251071) );
DFFARX1 I_14455  ( .D(I225107), .CLK(I5694_clk), .RSTB(I251103_rst), .Q(I251465) );
nor I_14456 (I251482,I251465,I251188);
nand I_14457 (I251089,I251352,I251482);
nor I_14458 (I251513,I251465,I251253);
not I_14459 (I251086,I251465);
nand I_14460 (I251544,I251465,I251154);
and I_14461 (I251561,I251222,I251544);
DFFARX1 I_14462  ( .D(I251561), .CLK(I5694_clk), .RSTB(I251103_rst), .Q(I251065) );
DFFARX1 I_14463  ( .D(I251465), .CLK(I5694_clk), .RSTB(I251103_rst), .Q(I251068) );
DFFARX1 I_14464  ( .D(I225116), .CLK(I5694_clk), .RSTB(I251103_rst), .Q(I251606) );
not I_14465 (I251623,I251606);
nand I_14466 (I251640,I251623,I251188);
and I_14467 (I251657,I251417,I251640);
DFFARX1 I_14468  ( .D(I251657), .CLK(I5694_clk), .RSTB(I251103_rst), .Q(I251095) );
or I_14469 (I251688,I251623,I251434);
DFFARX1 I_14470  ( .D(I251688), .CLK(I5694_clk), .RSTB(I251103_rst), .Q(I251080) );
nand I_14471 (I251083,I251623,I251513);
not I_14472 (I251766_rst,I5701);
not I_14473 (I251783,I194501);
nor I_14474 (I251800,I194498,I194516);
nand I_14475 (I251817,I251800,I194519);
nor I_14476 (I251834,I251783,I194498);
nand I_14477 (I251851,I251834,I194504);
not I_14478 (I251868,I251851);
not I_14479 (I251885,I194498);
nor I_14480 (I251755,I251851,I251885);
not I_14481 (I251916,I251885);
nand I_14482 (I251740,I251851,I251916);
not I_14483 (I251947,I194513);
nor I_14484 (I251964,I251947,I194495);
and I_14485 (I251981,I251964,I194489);
or I_14486 (I251998,I251981,I194507);
DFFARX1 I_14487  ( .D(I251998), .CLK(I5694_clk), .RSTB(I251766_rst), .Q(I252015) );
nor I_14488 (I252032,I252015,I251868);
DFFARX1 I_14489  ( .D(I252015), .CLK(I5694_clk), .RSTB(I251766_rst), .Q(I252049) );
not I_14490 (I251737,I252049);
nand I_14491 (I252080,I251783,I194513);
and I_14492 (I252097,I252080,I252032);
DFFARX1 I_14493  ( .D(I252080), .CLK(I5694_clk), .RSTB(I251766_rst), .Q(I251734) );
DFFARX1 I_14494  ( .D(I194492), .CLK(I5694_clk), .RSTB(I251766_rst), .Q(I252128) );
nor I_14495 (I252145,I252128,I251851);
nand I_14496 (I251752,I252015,I252145);
nor I_14497 (I252176,I252128,I251916);
not I_14498 (I251749,I252128);
nand I_14499 (I252207,I252128,I251817);
and I_14500 (I252224,I251885,I252207);
DFFARX1 I_14501  ( .D(I252224), .CLK(I5694_clk), .RSTB(I251766_rst), .Q(I251728) );
DFFARX1 I_14502  ( .D(I252128), .CLK(I5694_clk), .RSTB(I251766_rst), .Q(I251731) );
DFFARX1 I_14503  ( .D(I194510), .CLK(I5694_clk), .RSTB(I251766_rst), .Q(I252269) );
not I_14504 (I252286,I252269);
nand I_14505 (I252303,I252286,I251851);
and I_14506 (I252320,I252080,I252303);
DFFARX1 I_14507  ( .D(I252320), .CLK(I5694_clk), .RSTB(I251766_rst), .Q(I251758) );
or I_14508 (I252351,I252286,I252097);
DFFARX1 I_14509  ( .D(I252351), .CLK(I5694_clk), .RSTB(I251766_rst), .Q(I251743) );
nand I_14510 (I251746,I252286,I252176);
not I_14511 (I252429_rst,I5701);
not I_14512 (I252446,I234324);
nor I_14513 (I252463,I234315,I234306);
nand I_14514 (I252480,I252463,I234321);
nor I_14515 (I252497,I252446,I234315);
nand I_14516 (I252514,I252497,I234318);
DFFARX1 I_14517  ( .D(I252514), .CLK(I5694_clk), .RSTB(I252429_rst), .Q(I252531) );
not I_14518 (I252400,I252531);
not I_14519 (I252562,I234315);
not I_14520 (I252579,I252562);
not I_14521 (I252596,I234327);
nor I_14522 (I252613,I252596,I234312);
and I_14523 (I252630,I252613,I234330);
or I_14524 (I252647,I252630,I234303);
DFFARX1 I_14525  ( .D(I252647), .CLK(I5694_clk), .RSTB(I252429_rst), .Q(I252664) );
DFFARX1 I_14526  ( .D(I252664), .CLK(I5694_clk), .RSTB(I252429_rst), .Q(I252397) );
DFFARX1 I_14527  ( .D(I252664), .CLK(I5694_clk), .RSTB(I252429_rst), .Q(I252695) );
DFFARX1 I_14528  ( .D(I252664), .CLK(I5694_clk), .RSTB(I252429_rst), .Q(I252391) );
nand I_14529 (I252726,I252446,I234327);
nand I_14530 (I252743,I252726,I252480);
and I_14531 (I252760,I252562,I252743);
DFFARX1 I_14532  ( .D(I252760), .CLK(I5694_clk), .RSTB(I252429_rst), .Q(I252421) );
and I_14533 (I252394,I252726,I252695);
DFFARX1 I_14534  ( .D(I234333), .CLK(I5694_clk), .RSTB(I252429_rst), .Q(I252805) );
nor I_14535 (I252418,I252805,I252726);
nor I_14536 (I252836,I252805,I252480);
nand I_14537 (I252415,I252514,I252836);
not I_14538 (I252412,I252805);
DFFARX1 I_14539  ( .D(I234309), .CLK(I5694_clk), .RSTB(I252429_rst), .Q(I252881) );
not I_14540 (I252898,I252881);
nor I_14541 (I252915,I252898,I252579);
and I_14542 (I252932,I252805,I252915);
or I_14543 (I252949,I252726,I252932);
DFFARX1 I_14544  ( .D(I252949), .CLK(I5694_clk), .RSTB(I252429_rst), .Q(I252406) );
not I_14545 (I252980,I252898);
nor I_14546 (I252997,I252805,I252980);
nand I_14547 (I252409,I252898,I252997);
nand I_14548 (I252403,I252562,I252980);
not I_14549 (I253075_rst,I5701);
not I_14550 (I253092,I207745);
nor I_14551 (I253109,I207733,I207724);
nand I_14552 (I253126,I253109,I207736);
nor I_14553 (I253143,I253092,I207733);
nand I_14554 (I253160,I253143,I207742);
DFFARX1 I_14555  ( .D(I253160), .CLK(I5694_clk), .RSTB(I253075_rst), .Q(I253177) );
not I_14556 (I253046,I253177);
not I_14557 (I253208,I207733);
not I_14558 (I253225,I253208);
not I_14559 (I253242,I207718);
nor I_14560 (I253259,I253242,I207739);
and I_14561 (I253276,I253259,I207730);
or I_14562 (I253293,I253276,I207727);
DFFARX1 I_14563  ( .D(I253293), .CLK(I5694_clk), .RSTB(I253075_rst), .Q(I253310) );
DFFARX1 I_14564  ( .D(I253310), .CLK(I5694_clk), .RSTB(I253075_rst), .Q(I253043) );
DFFARX1 I_14565  ( .D(I253310), .CLK(I5694_clk), .RSTB(I253075_rst), .Q(I253341) );
DFFARX1 I_14566  ( .D(I253310), .CLK(I5694_clk), .RSTB(I253075_rst), .Q(I253037) );
nand I_14567 (I253372,I253092,I207718);
nand I_14568 (I253389,I253372,I253126);
and I_14569 (I253406,I253208,I253389);
DFFARX1 I_14570  ( .D(I253406), .CLK(I5694_clk), .RSTB(I253075_rst), .Q(I253067) );
and I_14571 (I253040,I253372,I253341);
DFFARX1 I_14572  ( .D(I207715), .CLK(I5694_clk), .RSTB(I253075_rst), .Q(I253451) );
nor I_14573 (I253064,I253451,I253372);
nor I_14574 (I253482,I253451,I253126);
nand I_14575 (I253061,I253160,I253482);
not I_14576 (I253058,I253451);
DFFARX1 I_14577  ( .D(I207721), .CLK(I5694_clk), .RSTB(I253075_rst), .Q(I253527) );
not I_14578 (I253544,I253527);
nor I_14579 (I253561,I253544,I253225);
and I_14580 (I253578,I253451,I253561);
or I_14581 (I253595,I253372,I253578);
DFFARX1 I_14582  ( .D(I253595), .CLK(I5694_clk), .RSTB(I253075_rst), .Q(I253052) );
not I_14583 (I253626,I253544);
nor I_14584 (I253643,I253451,I253626);
nand I_14585 (I253055,I253544,I253643);
nand I_14586 (I253049,I253208,I253626);
not I_14587 (I253721_rst,I5701);
not I_14588 (I253738,I247774);
nor I_14589 (I253755,I247753,I247765);
nand I_14590 (I253772,I253755,I247768);
nor I_14591 (I253789,I253738,I247753);
nand I_14592 (I253806,I253789,I247750);
DFFARX1 I_14593  ( .D(I253806), .CLK(I5694_clk), .RSTB(I253721_rst), .Q(I253823) );
not I_14594 (I253692,I253823);
not I_14595 (I253854,I247753);
not I_14596 (I253871,I253854);
not I_14597 (I253888,I247771);
nor I_14598 (I253905,I253888,I247762);
and I_14599 (I253922,I253905,I247756);
or I_14600 (I253939,I253922,I247780);
DFFARX1 I_14601  ( .D(I253939), .CLK(I5694_clk), .RSTB(I253721_rst), .Q(I253956) );
DFFARX1 I_14602  ( .D(I253956), .CLK(I5694_clk), .RSTB(I253721_rst), .Q(I253689) );
DFFARX1 I_14603  ( .D(I253956), .CLK(I5694_clk), .RSTB(I253721_rst), .Q(I253987) );
DFFARX1 I_14604  ( .D(I253956), .CLK(I5694_clk), .RSTB(I253721_rst), .Q(I253683) );
nand I_14605 (I254018,I253738,I247771);
nand I_14606 (I254035,I254018,I253772);
and I_14607 (I254052,I253854,I254035);
DFFARX1 I_14608  ( .D(I254052), .CLK(I5694_clk), .RSTB(I253721_rst), .Q(I253713) );
and I_14609 (I253686,I254018,I253987);
DFFARX1 I_14610  ( .D(I247777), .CLK(I5694_clk), .RSTB(I253721_rst), .Q(I254097) );
nor I_14611 (I253710,I254097,I254018);
nor I_14612 (I254128,I254097,I253772);
nand I_14613 (I253707,I253806,I254128);
not I_14614 (I253704,I254097);
DFFARX1 I_14615  ( .D(I247759), .CLK(I5694_clk), .RSTB(I253721_rst), .Q(I254173) );
not I_14616 (I254190,I254173);
nor I_14617 (I254207,I254190,I253871);
and I_14618 (I254224,I254097,I254207);
or I_14619 (I254241,I254018,I254224);
DFFARX1 I_14620  ( .D(I254241), .CLK(I5694_clk), .RSTB(I253721_rst), .Q(I253698) );
not I_14621 (I254272,I254190);
nor I_14622 (I254289,I254097,I254272);
nand I_14623 (I253701,I254190,I254289);
nand I_14624 (I253695,I253854,I254272);
not I_14625 (I254367_rst,I5701);
not I_14626 (I254384,I216080);
nor I_14627 (I254401,I216068,I216077);
nand I_14628 (I254418,I254401,I216092);
nor I_14629 (I254435,I254384,I216068);
nand I_14630 (I254452,I254435,I216074);
DFFARX1 I_14631  ( .D(I254452), .CLK(I5694_clk), .RSTB(I254367_rst), .Q(I254469) );
not I_14632 (I254338,I254469);
not I_14633 (I254500,I216068);
not I_14634 (I254517,I254500);
not I_14635 (I254534,I216062);
nor I_14636 (I254551,I254534,I216083);
and I_14637 (I254568,I254551,I216065);
or I_14638 (I254585,I254568,I216071);
DFFARX1 I_14639  ( .D(I254585), .CLK(I5694_clk), .RSTB(I254367_rst), .Q(I254602) );
DFFARX1 I_14640  ( .D(I254602), .CLK(I5694_clk), .RSTB(I254367_rst), .Q(I254335) );
DFFARX1 I_14641  ( .D(I254602), .CLK(I5694_clk), .RSTB(I254367_rst), .Q(I254633) );
DFFARX1 I_14642  ( .D(I254602), .CLK(I5694_clk), .RSTB(I254367_rst), .Q(I254329) );
nand I_14643 (I254664,I254384,I216062);
nand I_14644 (I254681,I254664,I254418);
and I_14645 (I254698,I254500,I254681);
DFFARX1 I_14646  ( .D(I254698), .CLK(I5694_clk), .RSTB(I254367_rst), .Q(I254359) );
and I_14647 (I254332,I254664,I254633);
DFFARX1 I_14648  ( .D(I216089), .CLK(I5694_clk), .RSTB(I254367_rst), .Q(I254743) );
nor I_14649 (I254356,I254743,I254664);
nor I_14650 (I254774,I254743,I254418);
nand I_14651 (I254353,I254452,I254774);
not I_14652 (I254350,I254743);
DFFARX1 I_14653  ( .D(I216086), .CLK(I5694_clk), .RSTB(I254367_rst), .Q(I254819) );
not I_14654 (I254836,I254819);
nor I_14655 (I254853,I254836,I254517);
and I_14656 (I254870,I254743,I254853);
or I_14657 (I254887,I254664,I254870);
DFFARX1 I_14658  ( .D(I254887), .CLK(I5694_clk), .RSTB(I254367_rst), .Q(I254344) );
not I_14659 (I254918,I254836);
nor I_14660 (I254935,I254743,I254918);
nand I_14661 (I254347,I254836,I254935);
nand I_14662 (I254341,I254500,I254918);
not I_14663 (I255013_rst,I5701);
not I_14664 (I255030,I229156);
nor I_14665 (I255047,I229147,I229138);
nand I_14666 (I255064,I255047,I229153);
nor I_14667 (I255081,I255030,I229147);
nand I_14668 (I255098,I255081,I229150);
DFFARX1 I_14669  ( .D(I255098), .CLK(I5694_clk), .RSTB(I255013_rst), .Q(I255115) );
not I_14670 (I254984,I255115);
not I_14671 (I255146,I229147);
not I_14672 (I255163,I255146);
not I_14673 (I255180,I229159);
nor I_14674 (I255197,I255180,I229144);
and I_14675 (I255214,I255197,I229162);
or I_14676 (I255231,I255214,I229135);
DFFARX1 I_14677  ( .D(I255231), .CLK(I5694_clk), .RSTB(I255013_rst), .Q(I255248) );
DFFARX1 I_14678  ( .D(I255248), .CLK(I5694_clk), .RSTB(I255013_rst), .Q(I254981) );
DFFARX1 I_14679  ( .D(I255248), .CLK(I5694_clk), .RSTB(I255013_rst), .Q(I255279) );
DFFARX1 I_14680  ( .D(I255248), .CLK(I5694_clk), .RSTB(I255013_rst), .Q(I254975) );
nand I_14681 (I255310,I255030,I229159);
nand I_14682 (I255327,I255310,I255064);
and I_14683 (I255344,I255146,I255327);
DFFARX1 I_14684  ( .D(I255344), .CLK(I5694_clk), .RSTB(I255013_rst), .Q(I255005) );
and I_14685 (I254978,I255310,I255279);
DFFARX1 I_14686  ( .D(I229165), .CLK(I5694_clk), .RSTB(I255013_rst), .Q(I255389) );
nor I_14687 (I255002,I255389,I255310);
nor I_14688 (I255420,I255389,I255064);
nand I_14689 (I254999,I255098,I255420);
not I_14690 (I254996,I255389);
DFFARX1 I_14691  ( .D(I229141), .CLK(I5694_clk), .RSTB(I255013_rst), .Q(I255465) );
not I_14692 (I255482,I255465);
nor I_14693 (I255499,I255482,I255163);
and I_14694 (I255516,I255389,I255499);
or I_14695 (I255533,I255310,I255516);
DFFARX1 I_14696  ( .D(I255533), .CLK(I5694_clk), .RSTB(I255013_rst), .Q(I254990) );
not I_14697 (I255564,I255482);
nor I_14698 (I255581,I255389,I255564);
nand I_14699 (I254993,I255482,I255581);
nand I_14700 (I254987,I255146,I255564);
not I_14701 (I255659_rst,I5701);
not I_14702 (I255676,I207133);
nor I_14703 (I255693,I207121,I207112);
nand I_14704 (I255710,I255693,I207124);
nor I_14705 (I255727,I255676,I207121);
nand I_14706 (I255744,I255727,I207130);
DFFARX1 I_14707  ( .D(I255744), .CLK(I5694_clk), .RSTB(I255659_rst), .Q(I255761) );
not I_14708 (I255630,I255761);
not I_14709 (I255792,I207121);
not I_14710 (I255809,I255792);
not I_14711 (I255826,I207106);
nor I_14712 (I255843,I255826,I207127);
and I_14713 (I255860,I255843,I207118);
or I_14714 (I255877,I255860,I207115);
DFFARX1 I_14715  ( .D(I255877), .CLK(I5694_clk), .RSTB(I255659_rst), .Q(I255894) );
DFFARX1 I_14716  ( .D(I255894), .CLK(I5694_clk), .RSTB(I255659_rst), .Q(I255627) );
DFFARX1 I_14717  ( .D(I255894), .CLK(I5694_clk), .RSTB(I255659_rst), .Q(I255925) );
DFFARX1 I_14718  ( .D(I255894), .CLK(I5694_clk), .RSTB(I255659_rst), .Q(I255621) );
nand I_14719 (I255956,I255676,I207106);
nand I_14720 (I255973,I255956,I255710);
and I_14721 (I255990,I255792,I255973);
DFFARX1 I_14722  ( .D(I255990), .CLK(I5694_clk), .RSTB(I255659_rst), .Q(I255651) );
and I_14723 (I255624,I255956,I255925);
DFFARX1 I_14724  ( .D(I207103), .CLK(I5694_clk), .RSTB(I255659_rst), .Q(I256035) );
nor I_14725 (I255648,I256035,I255956);
nor I_14726 (I256066,I256035,I255710);
nand I_14727 (I255645,I255744,I256066);
not I_14728 (I255642,I256035);
DFFARX1 I_14729  ( .D(I207109), .CLK(I5694_clk), .RSTB(I255659_rst), .Q(I256111) );
not I_14730 (I256128,I256111);
nor I_14731 (I256145,I256128,I255809);
and I_14732 (I256162,I256035,I256145);
or I_14733 (I256179,I255956,I256162);
DFFARX1 I_14734  ( .D(I256179), .CLK(I5694_clk), .RSTB(I255659_rst), .Q(I255636) );
not I_14735 (I256210,I256128);
nor I_14736 (I256227,I256035,I256210);
nand I_14737 (I255639,I256128,I256227);
nand I_14738 (I255633,I255792,I256210);
not I_14739 (I256305_rst,I5701);
not I_14740 (I256322,I200760);
nor I_14741 (I256339,I200763,I200745);
nand I_14742 (I256356,I256339,I200772);
nor I_14743 (I256373,I256322,I200763);
nand I_14744 (I256390,I256373,I200751);
DFFARX1 I_14745  ( .D(I256390), .CLK(I5694_clk), .RSTB(I256305_rst), .Q(I256407) );
not I_14746 (I256276,I256407);
not I_14747 (I256438,I200763);
not I_14748 (I256455,I256438);
not I_14749 (I256472,I200757);
nor I_14750 (I256489,I256472,I200769);
and I_14751 (I256506,I256489,I200775);
or I_14752 (I256523,I256506,I200754);
DFFARX1 I_14753  ( .D(I256523), .CLK(I5694_clk), .RSTB(I256305_rst), .Q(I256540) );
DFFARX1 I_14754  ( .D(I256540), .CLK(I5694_clk), .RSTB(I256305_rst), .Q(I256273) );
DFFARX1 I_14755  ( .D(I256540), .CLK(I5694_clk), .RSTB(I256305_rst), .Q(I256571) );
DFFARX1 I_14756  ( .D(I256540), .CLK(I5694_clk), .RSTB(I256305_rst), .Q(I256267) );
nand I_14757 (I256602,I256322,I200757);
nand I_14758 (I256619,I256602,I256356);
and I_14759 (I256636,I256438,I256619);
DFFARX1 I_14760  ( .D(I256636), .CLK(I5694_clk), .RSTB(I256305_rst), .Q(I256297) );
and I_14761 (I256270,I256602,I256571);
DFFARX1 I_14762  ( .D(I200766), .CLK(I5694_clk), .RSTB(I256305_rst), .Q(I256681) );
nor I_14763 (I256294,I256681,I256602);
nor I_14764 (I256712,I256681,I256356);
nand I_14765 (I256291,I256390,I256712);
not I_14766 (I256288,I256681);
DFFARX1 I_14767  ( .D(I200748), .CLK(I5694_clk), .RSTB(I256305_rst), .Q(I256757) );
not I_14768 (I256774,I256757);
nor I_14769 (I256791,I256774,I256455);
and I_14770 (I256808,I256681,I256791);
or I_14771 (I256825,I256602,I256808);
DFFARX1 I_14772  ( .D(I256825), .CLK(I5694_clk), .RSTB(I256305_rst), .Q(I256282) );
not I_14773 (I256856,I256774);
nor I_14774 (I256873,I256681,I256856);
nand I_14775 (I256285,I256774,I256873);
nand I_14776 (I256279,I256438,I256856);
not I_14777 (I256951_rst,I5701);
not I_14778 (I256968,I208957);
nor I_14779 (I256985,I208963,I208948);
nand I_14780 (I257002,I256985,I208942);
nor I_14781 (I257019,I256968,I208963);
nand I_14782 (I257036,I257019,I208969);
DFFARX1 I_14783  ( .D(I257036), .CLK(I5694_clk), .RSTB(I256951_rst), .Q(I257053) );
not I_14784 (I256922,I257053);
not I_14785 (I257084,I208963);
not I_14786 (I257101,I257084);
not I_14787 (I257118,I208954);
nor I_14788 (I257135,I257118,I208960);
and I_14789 (I257152,I257135,I208966);
or I_14790 (I257169,I257152,I208939);
DFFARX1 I_14791  ( .D(I257169), .CLK(I5694_clk), .RSTB(I256951_rst), .Q(I257186) );
DFFARX1 I_14792  ( .D(I257186), .CLK(I5694_clk), .RSTB(I256951_rst), .Q(I256919) );
DFFARX1 I_14793  ( .D(I257186), .CLK(I5694_clk), .RSTB(I256951_rst), .Q(I257217) );
DFFARX1 I_14794  ( .D(I257186), .CLK(I5694_clk), .RSTB(I256951_rst), .Q(I256913) );
nand I_14795 (I257248,I256968,I208954);
nand I_14796 (I257265,I257248,I257002);
and I_14797 (I257282,I257084,I257265);
DFFARX1 I_14798  ( .D(I257282), .CLK(I5694_clk), .RSTB(I256951_rst), .Q(I256943) );
and I_14799 (I256916,I257248,I257217);
DFFARX1 I_14800  ( .D(I208945), .CLK(I5694_clk), .RSTB(I256951_rst), .Q(I257327) );
nor I_14801 (I256940,I257327,I257248);
nor I_14802 (I257358,I257327,I257002);
nand I_14803 (I256937,I257036,I257358);
not I_14804 (I256934,I257327);
DFFARX1 I_14805  ( .D(I208951), .CLK(I5694_clk), .RSTB(I256951_rst), .Q(I257403) );
not I_14806 (I257420,I257403);
nor I_14807 (I257437,I257420,I257101);
and I_14808 (I257454,I257327,I257437);
or I_14809 (I257471,I257248,I257454);
DFFARX1 I_14810  ( .D(I257471), .CLK(I5694_clk), .RSTB(I256951_rst), .Q(I256928) );
not I_14811 (I257502,I257420);
nor I_14812 (I257519,I257327,I257502);
nand I_14813 (I256931,I257420,I257519);
nand I_14814 (I256925,I257084,I257502);
not I_14815 (I257597_rst,I5701);
not I_14816 (I257614,I228510);
nor I_14817 (I257631,I228501,I228492);
nand I_14818 (I257648,I257631,I228507);
nor I_14819 (I257665,I257614,I228501);
nand I_14820 (I257682,I257665,I228504);
DFFARX1 I_14821  ( .D(I257682), .CLK(I5694_clk), .RSTB(I257597_rst), .Q(I257699) );
not I_14822 (I257568,I257699);
not I_14823 (I257730,I228501);
not I_14824 (I257747,I257730);
not I_14825 (I257764,I228513);
nor I_14826 (I257781,I257764,I228498);
and I_14827 (I257798,I257781,I228516);
or I_14828 (I257815,I257798,I228489);
DFFARX1 I_14829  ( .D(I257815), .CLK(I5694_clk), .RSTB(I257597_rst), .Q(I257832) );
DFFARX1 I_14830  ( .D(I257832), .CLK(I5694_clk), .RSTB(I257597_rst), .Q(I257565) );
DFFARX1 I_14831  ( .D(I257832), .CLK(I5694_clk), .RSTB(I257597_rst), .Q(I257863) );
DFFARX1 I_14832  ( .D(I257832), .CLK(I5694_clk), .RSTB(I257597_rst), .Q(I257559) );
nand I_14833 (I257894,I257614,I228513);
nand I_14834 (I257911,I257894,I257648);
and I_14835 (I257928,I257730,I257911);
DFFARX1 I_14836  ( .D(I257928), .CLK(I5694_clk), .RSTB(I257597_rst), .Q(I257589) );
and I_14837 (I257562,I257894,I257863);
DFFARX1 I_14838  ( .D(I228519), .CLK(I5694_clk), .RSTB(I257597_rst), .Q(I257973) );
nor I_14839 (I257586,I257973,I257894);
nor I_14840 (I258004,I257973,I257648);
nand I_14841 (I257583,I257682,I258004);
not I_14842 (I257580,I257973);
DFFARX1 I_14843  ( .D(I228495), .CLK(I5694_clk), .RSTB(I257597_rst), .Q(I258049) );
not I_14844 (I258066,I258049);
nor I_14845 (I258083,I258066,I257747);
and I_14846 (I258100,I257973,I258083);
or I_14847 (I258117,I257894,I258100);
DFFARX1 I_14848  ( .D(I258117), .CLK(I5694_clk), .RSTB(I257597_rst), .Q(I257574) );
not I_14849 (I258148,I258066);
nor I_14850 (I258165,I257973,I258148);
nand I_14851 (I257577,I258066,I258165);
nand I_14852 (I257571,I257730,I258148);
not I_14853 (I258243_rst,I5701);
not I_14854 (I258260,I230448);
nor I_14855 (I258277,I230439,I230430);
nand I_14856 (I258294,I258277,I230445);
nor I_14857 (I258311,I258260,I230439);
nand I_14858 (I258328,I258311,I230442);
DFFARX1 I_14859  ( .D(I258328), .CLK(I5694_clk), .RSTB(I258243_rst), .Q(I258345) );
not I_14860 (I258214,I258345);
not I_14861 (I258376,I230439);
not I_14862 (I258393,I258376);
not I_14863 (I258410,I230451);
nor I_14864 (I258427,I258410,I230436);
and I_14865 (I258444,I258427,I230454);
or I_14866 (I258461,I258444,I230427);
DFFARX1 I_14867  ( .D(I258461), .CLK(I5694_clk), .RSTB(I258243_rst), .Q(I258478) );
DFFARX1 I_14868  ( .D(I258478), .CLK(I5694_clk), .RSTB(I258243_rst), .Q(I258211) );
DFFARX1 I_14869  ( .D(I258478), .CLK(I5694_clk), .RSTB(I258243_rst), .Q(I258509) );
DFFARX1 I_14870  ( .D(I258478), .CLK(I5694_clk), .RSTB(I258243_rst), .Q(I258205) );
nand I_14871 (I258540,I258260,I230451);
nand I_14872 (I258557,I258540,I258294);
and I_14873 (I258574,I258376,I258557);
DFFARX1 I_14874  ( .D(I258574), .CLK(I5694_clk), .RSTB(I258243_rst), .Q(I258235) );
and I_14875 (I258208,I258540,I258509);
DFFARX1 I_14876  ( .D(I230457), .CLK(I5694_clk), .RSTB(I258243_rst), .Q(I258619) );
nor I_14877 (I258232,I258619,I258540);
nor I_14878 (I258650,I258619,I258294);
nand I_14879 (I258229,I258328,I258650);
not I_14880 (I258226,I258619);
DFFARX1 I_14881  ( .D(I230433), .CLK(I5694_clk), .RSTB(I258243_rst), .Q(I258695) );
not I_14882 (I258712,I258695);
nor I_14883 (I258729,I258712,I258393);
and I_14884 (I258746,I258619,I258729);
or I_14885 (I258763,I258540,I258746);
DFFARX1 I_14886  ( .D(I258763), .CLK(I5694_clk), .RSTB(I258243_rst), .Q(I258220) );
not I_14887 (I258794,I258712);
nor I_14888 (I258811,I258619,I258794);
nand I_14889 (I258223,I258712,I258811);
nand I_14890 (I258217,I258376,I258794);
not I_14891 (I258889_rst,I5701);
or I_14892 (I258906,I216663,I216684);
or I_14893 (I258923,I216669,I216663);
nor I_14894 (I258940,I216672,I216660);
DFFARX1 I_14895  ( .D(I258940), .CLK(I5694_clk), .RSTB(I258889_rst), .Q(I258957) );
DFFARX1 I_14896  ( .D(I258940), .CLK(I5694_clk), .RSTB(I258889_rst), .Q(I258851) );
not I_14897 (I258988,I216672);
and I_14898 (I259005,I258988,I216678);
nor I_14899 (I259022,I259005,I216684);
nor I_14900 (I259039,I216666,I216681);
DFFARX1 I_14901  ( .D(I259039), .CLK(I5694_clk), .RSTB(I258889_rst), .Q(I259056) );
not I_14902 (I259073,I259056);
DFFARX1 I_14903  ( .D(I259056), .CLK(I5694_clk), .RSTB(I258889_rst), .Q(I258860) );
nor I_14904 (I259104,I216666,I216669);
and I_14905 (I258854,I259104,I258957);
DFFARX1 I_14906  ( .D(I216657), .CLK(I5694_clk), .RSTB(I258889_rst), .Q(I259135) );
and I_14907 (I259152,I259135,I216687);
nand I_14908 (I259169,I259152,I258923);
and I_14909 (I259186,I259056,I259169);
DFFARX1 I_14910  ( .D(I259186), .CLK(I5694_clk), .RSTB(I258889_rst), .Q(I258881) );
nor I_14911 (I258878,I259152,I259022);
not I_14912 (I259231,I259152);
nor I_14913 (I259248,I258906,I259231);
nor I_14914 (I259265,I259152,I259104);
nand I_14915 (I258875,I258923,I259265);
nor I_14916 (I259296,I259152,I259073);
not I_14917 (I258872,I259152);
nand I_14918 (I258863,I259152,I259073);
DFFARX1 I_14919  ( .D(I216675), .CLK(I5694_clk), .RSTB(I258889_rst), .Q(I259341) );
and I_14920 (I259358,I259341,I259248);
or I_14921 (I259375,I258906,I259358);
DFFARX1 I_14922  ( .D(I259375), .CLK(I5694_clk), .RSTB(I258889_rst), .Q(I258866) );
nand I_14923 (I258869,I259341,I259296);
nand I_14924 (I259420,I259341,I259022);
and I_14925 (I259437,I258940,I259420);
DFFARX1 I_14926  ( .D(I259437), .CLK(I5694_clk), .RSTB(I258889_rst), .Q(I258857) );
not I_14927 (I259501_rst,I5701);
nand I_14928 (I259518,I242011,I241996);
and I_14929 (I259535,I259518,I242005);
DFFARX1 I_14930  ( .D(I259535), .CLK(I5694_clk), .RSTB(I259501_rst), .Q(I259552) );
not I_14931 (I259569,I259552);
DFFARX1 I_14932  ( .D(I259552), .CLK(I5694_clk), .RSTB(I259501_rst), .Q(I259469) );
nor I_14933 (I259600,I242014,I241996);
DFFARX1 I_14934  ( .D(I241993), .CLK(I5694_clk), .RSTB(I259501_rst), .Q(I259617) );
DFFARX1 I_14935  ( .D(I259617), .CLK(I5694_clk), .RSTB(I259501_rst), .Q(I259634) );
not I_14936 (I259472,I259634);
DFFARX1 I_14937  ( .D(I259617), .CLK(I5694_clk), .RSTB(I259501_rst), .Q(I259665) );
and I_14938 (I259466,I259552,I259665);
nand I_14939 (I259696,I242017,I241990);
and I_14940 (I259713,I259696,I242008);
DFFARX1 I_14941  ( .D(I259713), .CLK(I5694_clk), .RSTB(I259501_rst), .Q(I259730) );
nor I_14942 (I259747,I259730,I259569);
not I_14943 (I259764,I259730);
nand I_14944 (I259475,I259552,I259764);
DFFARX1 I_14945  ( .D(I242002), .CLK(I5694_clk), .RSTB(I259501_rst), .Q(I259795) );
and I_14946 (I259812,I259795,I241987);
nor I_14947 (I259829,I259812,I259730);
nor I_14948 (I259846,I259812,I259764);
nand I_14949 (I259481,I259600,I259846);
not I_14950 (I259484,I259812);
DFFARX1 I_14951  ( .D(I259812), .CLK(I5694_clk), .RSTB(I259501_rst), .Q(I259463) );
DFFARX1 I_14952  ( .D(I241999), .CLK(I5694_clk), .RSTB(I259501_rst), .Q(I259905) );
nand I_14953 (I259922,I259905,I259617);
and I_14954 (I259939,I259600,I259922);
DFFARX1 I_14955  ( .D(I259939), .CLK(I5694_clk), .RSTB(I259501_rst), .Q(I259493) );
nor I_14956 (I259490,I259905,I259812);
and I_14957 (I259984,I259905,I259747);
or I_14958 (I260001,I259600,I259984);
DFFARX1 I_14959  ( .D(I260001), .CLK(I5694_clk), .RSTB(I259501_rst), .Q(I259478) );
nand I_14960 (I259487,I259905,I259829);
not I_14961 (I260079_rst,I5701);
nand I_14962 (I260096,I211329,I211317);
and I_14963 (I260113,I260096,I211311);
DFFARX1 I_14964  ( .D(I260113), .CLK(I5694_clk), .RSTB(I260079_rst), .Q(I260130) );
not I_14965 (I260147,I260130);
DFFARX1 I_14966  ( .D(I260130), .CLK(I5694_clk), .RSTB(I260079_rst), .Q(I260047) );
nor I_14967 (I260178,I211308,I211317);
DFFARX1 I_14968  ( .D(I211302), .CLK(I5694_clk), .RSTB(I260079_rst), .Q(I260195) );
DFFARX1 I_14969  ( .D(I260195), .CLK(I5694_clk), .RSTB(I260079_rst), .Q(I260212) );
not I_14970 (I260050,I260212);
DFFARX1 I_14971  ( .D(I260195), .CLK(I5694_clk), .RSTB(I260079_rst), .Q(I260243) );
and I_14972 (I260044,I260130,I260243);
nand I_14973 (I260274,I211305,I211320);
and I_14974 (I260291,I260274,I211332);
DFFARX1 I_14975  ( .D(I260291), .CLK(I5694_clk), .RSTB(I260079_rst), .Q(I260308) );
nor I_14976 (I260325,I260308,I260147);
not I_14977 (I260342,I260308);
nand I_14978 (I260053,I260130,I260342);
DFFARX1 I_14979  ( .D(I211323), .CLK(I5694_clk), .RSTB(I260079_rst), .Q(I260373) );
and I_14980 (I260390,I260373,I211314);
nor I_14981 (I260407,I260390,I260308);
nor I_14982 (I260424,I260390,I260342);
nand I_14983 (I260059,I260178,I260424);
not I_14984 (I260062,I260390);
DFFARX1 I_14985  ( .D(I260390), .CLK(I5694_clk), .RSTB(I260079_rst), .Q(I260041) );
DFFARX1 I_14986  ( .D(I211326), .CLK(I5694_clk), .RSTB(I260079_rst), .Q(I260483) );
nand I_14987 (I260500,I260483,I260195);
and I_14988 (I260517,I260178,I260500);
DFFARX1 I_14989  ( .D(I260517), .CLK(I5694_clk), .RSTB(I260079_rst), .Q(I260071) );
nor I_14990 (I260068,I260483,I260390);
and I_14991 (I260562,I260483,I260325);
or I_14992 (I260579,I260178,I260562);
DFFARX1 I_14993  ( .D(I260579), .CLK(I5694_clk), .RSTB(I260079_rst), .Q(I260056) );
nand I_14994 (I260065,I260483,I260407);
not I_14995 (I260657_rst,I5701);
nand I_14996 (I260674,I247090,I247117);
and I_14997 (I260691,I260674,I247105);
DFFARX1 I_14998  ( .D(I260691), .CLK(I5694_clk), .RSTB(I260657_rst), .Q(I260708) );
not I_14999 (I260725,I260708);
DFFARX1 I_15000  ( .D(I260708), .CLK(I5694_clk), .RSTB(I260657_rst), .Q(I260625) );
nor I_15001 (I260756,I247093,I247117);
DFFARX1 I_15002  ( .D(I247108), .CLK(I5694_clk), .RSTB(I260657_rst), .Q(I260773) );
DFFARX1 I_15003  ( .D(I260773), .CLK(I5694_clk), .RSTB(I260657_rst), .Q(I260790) );
not I_15004 (I260628,I260790);
DFFARX1 I_15005  ( .D(I260773), .CLK(I5694_clk), .RSTB(I260657_rst), .Q(I260821) );
and I_15006 (I260622,I260708,I260821);
nand I_15007 (I260852,I247102,I247099);
and I_15008 (I260869,I260852,I247096);
DFFARX1 I_15009  ( .D(I260869), .CLK(I5694_clk), .RSTB(I260657_rst), .Q(I260886) );
nor I_15010 (I260903,I260886,I260725);
not I_15011 (I260920,I260886);
nand I_15012 (I260631,I260708,I260920);
DFFARX1 I_15013  ( .D(I247111), .CLK(I5694_clk), .RSTB(I260657_rst), .Q(I260951) );
and I_15014 (I260968,I260951,I247087);
nor I_15015 (I260985,I260968,I260886);
nor I_15016 (I261002,I260968,I260920);
nand I_15017 (I260637,I260756,I261002);
not I_15018 (I260640,I260968);
DFFARX1 I_15019  ( .D(I260968), .CLK(I5694_clk), .RSTB(I260657_rst), .Q(I260619) );
DFFARX1 I_15020  ( .D(I247114), .CLK(I5694_clk), .RSTB(I260657_rst), .Q(I261061) );
nand I_15021 (I261078,I261061,I260773);
and I_15022 (I261095,I260756,I261078);
DFFARX1 I_15023  ( .D(I261095), .CLK(I5694_clk), .RSTB(I260657_rst), .Q(I260649) );
nor I_15024 (I260646,I261061,I260968);
and I_15025 (I261140,I261061,I260903);
or I_15026 (I261157,I260756,I261140);
DFFARX1 I_15027  ( .D(I261157), .CLK(I5694_clk), .RSTB(I260657_rst), .Q(I260634) );
nand I_15028 (I260643,I261061,I260985);
not I_15029 (I261235_rst,I5701);
nand I_15030 (I261252,I241416,I241401);
and I_15031 (I261269,I261252,I241410);
DFFARX1 I_15032  ( .D(I261269), .CLK(I5694_clk), .RSTB(I261235_rst), .Q(I261286) );
not I_15033 (I261303,I261286);
DFFARX1 I_15034  ( .D(I261286), .CLK(I5694_clk), .RSTB(I261235_rst), .Q(I261203) );
nor I_15035 (I261334,I241419,I241401);
DFFARX1 I_15036  ( .D(I241398), .CLK(I5694_clk), .RSTB(I261235_rst), .Q(I261351) );
DFFARX1 I_15037  ( .D(I261351), .CLK(I5694_clk), .RSTB(I261235_rst), .Q(I261368) );
not I_15038 (I261206,I261368);
DFFARX1 I_15039  ( .D(I261351), .CLK(I5694_clk), .RSTB(I261235_rst), .Q(I261399) );
and I_15040 (I261200,I261286,I261399);
nand I_15041 (I261430,I241422,I241395);
and I_15042 (I261447,I261430,I241413);
DFFARX1 I_15043  ( .D(I261447), .CLK(I5694_clk), .RSTB(I261235_rst), .Q(I261464) );
nor I_15044 (I261481,I261464,I261303);
not I_15045 (I261498,I261464);
nand I_15046 (I261209,I261286,I261498);
DFFARX1 I_15047  ( .D(I241407), .CLK(I5694_clk), .RSTB(I261235_rst), .Q(I261529) );
and I_15048 (I261546,I261529,I241392);
nor I_15049 (I261563,I261546,I261464);
nor I_15050 (I261580,I261546,I261498);
nand I_15051 (I261215,I261334,I261580);
not I_15052 (I261218,I261546);
DFFARX1 I_15053  ( .D(I261546), .CLK(I5694_clk), .RSTB(I261235_rst), .Q(I261197) );
DFFARX1 I_15054  ( .D(I241404), .CLK(I5694_clk), .RSTB(I261235_rst), .Q(I261639) );
nand I_15055 (I261656,I261639,I261351);
and I_15056 (I261673,I261334,I261656);
DFFARX1 I_15057  ( .D(I261673), .CLK(I5694_clk), .RSTB(I261235_rst), .Q(I261227) );
nor I_15058 (I261224,I261639,I261546);
and I_15059 (I261718,I261639,I261481);
or I_15060 (I261735,I261334,I261718);
DFFARX1 I_15061  ( .D(I261735), .CLK(I5694_clk), .RSTB(I261235_rst), .Q(I261212) );
nand I_15062 (I261221,I261639,I261563);
not I_15063 (I261813_rst,I5701);
nand I_15064 (I261830,I250405,I250432);
and I_15065 (I261847,I261830,I250420);
DFFARX1 I_15066  ( .D(I261847), .CLK(I5694_clk), .RSTB(I261813_rst), .Q(I261864) );
not I_15067 (I261881,I261864);
DFFARX1 I_15068  ( .D(I261864), .CLK(I5694_clk), .RSTB(I261813_rst), .Q(I261781) );
nor I_15069 (I261912,I250408,I250432);
DFFARX1 I_15070  ( .D(I250423), .CLK(I5694_clk), .RSTB(I261813_rst), .Q(I261929) );
DFFARX1 I_15071  ( .D(I261929), .CLK(I5694_clk), .RSTB(I261813_rst), .Q(I261946) );
not I_15072 (I261784,I261946);
DFFARX1 I_15073  ( .D(I261929), .CLK(I5694_clk), .RSTB(I261813_rst), .Q(I261977) );
and I_15074 (I261778,I261864,I261977);
nand I_15075 (I262008,I250417,I250414);
and I_15076 (I262025,I262008,I250411);
DFFARX1 I_15077  ( .D(I262025), .CLK(I5694_clk), .RSTB(I261813_rst), .Q(I262042) );
nor I_15078 (I262059,I262042,I261881);
not I_15079 (I262076,I262042);
nand I_15080 (I261787,I261864,I262076);
DFFARX1 I_15081  ( .D(I250426), .CLK(I5694_clk), .RSTB(I261813_rst), .Q(I262107) );
and I_15082 (I262124,I262107,I250402);
nor I_15083 (I262141,I262124,I262042);
nor I_15084 (I262158,I262124,I262076);
nand I_15085 (I261793,I261912,I262158);
not I_15086 (I261796,I262124);
DFFARX1 I_15087  ( .D(I262124), .CLK(I5694_clk), .RSTB(I261813_rst), .Q(I261775) );
DFFARX1 I_15088  ( .D(I250429), .CLK(I5694_clk), .RSTB(I261813_rst), .Q(I262217) );
nand I_15089 (I262234,I262217,I261929);
and I_15090 (I262251,I261912,I262234);
DFFARX1 I_15091  ( .D(I262251), .CLK(I5694_clk), .RSTB(I261813_rst), .Q(I261805) );
nor I_15092 (I261802,I262217,I262124);
and I_15093 (I262296,I262217,I262059);
or I_15094 (I262313,I261912,I262296);
DFFARX1 I_15095  ( .D(I262313), .CLK(I5694_clk), .RSTB(I261813_rst), .Q(I261790) );
nand I_15096 (I261799,I262217,I262141);
not I_15097 (I262391_rst,I5701);
nand I_15098 (I262408,I23626_rst2,I236244);
and I_15099 (I262425,I262408,I236256);
DFFARX1 I_15100  ( .D(I262425), .CLK(I5694_clk), .RSTB(I262391_rst), .Q(I262442) );
not I_15101 (I262459,I262442);
DFFARX1 I_15102  ( .D(I262442), .CLK(I5694_clk), .RSTB(I262391_rst), .Q(I262359) );
nor I_15103 (I262490,I236259,I236244);
DFFARX1 I_15104  ( .D(I23626_rst8), .CLK(I5694_clk), .RSTB(I262391_rst), .Q(I262507) );
DFFARX1 I_15105  ( .D(I262507), .CLK(I5694_clk), .RSTB(I262391_rst), .Q(I262524) );
not I_15106 (I262362,I262524);
DFFARX1 I_15107  ( .D(I262507), .CLK(I5694_clk), .RSTB(I262391_rst), .Q(I262555) );
and I_15108 (I262356,I262442,I262555);
nand I_15109 (I262586,I236247,I236271);
and I_15110 (I262603,I262586,I236250);
DFFARX1 I_15111  ( .D(I262603), .CLK(I5694_clk), .RSTB(I262391_rst), .Q(I262620) );
nor I_15112 (I262637,I262620,I262459);
not I_15113 (I262654,I262620);
nand I_15114 (I262365,I262442,I262654);
DFFARX1 I_15115  ( .D(I236253), .CLK(I5694_clk), .RSTB(I262391_rst), .Q(I262685) );
and I_15116 (I262702,I262685,I23626_rst5);
nor I_15117 (I262719,I262702,I262620);
nor I_15118 (I262736,I262702,I262654);
nand I_15119 (I262371,I262490,I262736);
not I_15120 (I262374,I262702);
DFFARX1 I_15121  ( .D(I262702), .CLK(I5694_clk), .RSTB(I262391_rst), .Q(I262353) );
DFFARX1 I_15122  ( .D(I236241), .CLK(I5694_clk), .RSTB(I262391_rst), .Q(I262795) );
nand I_15123 (I262812,I262795,I262507);
and I_15124 (I262829,I262490,I262812);
DFFARX1 I_15125  ( .D(I262829), .CLK(I5694_clk), .RSTB(I262391_rst), .Q(I262383) );
nor I_15126 (I262380,I262795,I262702);
and I_15127 (I262874,I262795,I262637);
or I_15128 (I262891,I262490,I262874);
DFFARX1 I_15129  ( .D(I262891), .CLK(I5694_clk), .RSTB(I262391_rst), .Q(I262368) );
nand I_15130 (I262377,I262795,I262719);
not I_15131 (I262969_rst,I5701);
nand I_15132 (I262986,I256928,I256925);
and I_15133 (I263003,I262986,I256937);
DFFARX1 I_15134  ( .D(I263003), .CLK(I5694_clk), .RSTB(I262969_rst), .Q(I263020) );
not I_15135 (I263037,I263020);
DFFARX1 I_15136  ( .D(I263020), .CLK(I5694_clk), .RSTB(I262969_rst), .Q(I262937) );
nor I_15137 (I263068,I256934,I256925);
DFFARX1 I_15138  ( .D(I256940), .CLK(I5694_clk), .RSTB(I262969_rst), .Q(I263085) );
DFFARX1 I_15139  ( .D(I263085), .CLK(I5694_clk), .RSTB(I262969_rst), .Q(I263102) );
not I_15140 (I262940,I263102);
DFFARX1 I_15141  ( .D(I263085), .CLK(I5694_clk), .RSTB(I262969_rst), .Q(I263133) );
and I_15142 (I262934,I263020,I263133);
nand I_15143 (I263164,I256916,I256919);
and I_15144 (I263181,I263164,I256943);
DFFARX1 I_15145  ( .D(I263181), .CLK(I5694_clk), .RSTB(I262969_rst), .Q(I263198) );
nor I_15146 (I263215,I263198,I263037);
not I_15147 (I263232,I263198);
nand I_15148 (I262943,I263020,I263232);
DFFARX1 I_15149  ( .D(I256922), .CLK(I5694_clk), .RSTB(I262969_rst), .Q(I263263) );
and I_15150 (I263280,I263263,I256913);
nor I_15151 (I263297,I263280,I263198);
nor I_15152 (I263314,I263280,I263232);
nand I_15153 (I262949,I263068,I263314);
not I_15154 (I262952,I263280);
DFFARX1 I_15155  ( .D(I263280), .CLK(I5694_clk), .RSTB(I262969_rst), .Q(I262931) );
DFFARX1 I_15156  ( .D(I256931), .CLK(I5694_clk), .RSTB(I262969_rst), .Q(I263373) );
nand I_15157 (I263390,I263373,I263085);
and I_15158 (I263407,I263068,I263390);
DFFARX1 I_15159  ( .D(I263407), .CLK(I5694_clk), .RSTB(I262969_rst), .Q(I262961) );
nor I_15160 (I262958,I263373,I263280);
and I_15161 (I263452,I263373,I263215);
or I_15162 (I263469,I263068,I263452);
DFFARX1 I_15163  ( .D(I263469), .CLK(I5694_clk), .RSTB(I262969_rst), .Q(I262946) );
nand I_15164 (I262955,I263373,I263297);
not I_15165 (I263547_rst,I5701);
nand I_15166 (I263564,I215476,I215473);
and I_15167 (I263581,I263564,I215467);
DFFARX1 I_15168  ( .D(I263581), .CLK(I5694_clk), .RSTB(I263547_rst), .Q(I263598) );
not I_15169 (I263615,I263598);
DFFARX1 I_15170  ( .D(I263598), .CLK(I5694_clk), .RSTB(I263547_rst), .Q(I263515) );
nor I_15171 (I263646,I215488,I215473);
DFFARX1 I_15172  ( .D(I215491), .CLK(I5694_clk), .RSTB(I263547_rst), .Q(I263663) );
DFFARX1 I_15173  ( .D(I263663), .CLK(I5694_clk), .RSTB(I263547_rst), .Q(I263680) );
not I_15174 (I263518,I263680);
DFFARX1 I_15175  ( .D(I263663), .CLK(I5694_clk), .RSTB(I263547_rst), .Q(I263711) );
and I_15176 (I263512,I263598,I263711);
nand I_15177 (I263742,I215494,I215485);
and I_15178 (I263759,I263742,I215497);
DFFARX1 I_15179  ( .D(I263759), .CLK(I5694_clk), .RSTB(I263547_rst), .Q(I263776) );
nor I_15180 (I263793,I263776,I263615);
not I_15181 (I263810,I263776);
nand I_15182 (I263521,I263598,I263810);
DFFARX1 I_15183  ( .D(I215470), .CLK(I5694_clk), .RSTB(I263547_rst), .Q(I263841) );
and I_15184 (I263858,I263841,I215479);
nor I_15185 (I263875,I263858,I263776);
nor I_15186 (I263892,I263858,I263810);
nand I_15187 (I263527,I263646,I263892);
not I_15188 (I263530,I263858);
DFFARX1 I_15189  ( .D(I263858), .CLK(I5694_clk), .RSTB(I263547_rst), .Q(I263509) );
DFFARX1 I_15190  ( .D(I215482), .CLK(I5694_clk), .RSTB(I263547_rst), .Q(I263951) );
nand I_15191 (I263968,I263951,I263663);
and I_15192 (I263985,I263646,I263968);
DFFARX1 I_15193  ( .D(I263985), .CLK(I5694_clk), .RSTB(I263547_rst), .Q(I263539) );
nor I_15194 (I263536,I263951,I263858);
and I_15195 (I264030,I263951,I263793);
or I_15196 (I264047,I263646,I264030);
DFFARX1 I_15197  ( .D(I264047), .CLK(I5694_clk), .RSTB(I263547_rst), .Q(I263524) );
nand I_15198 (I263533,I263951,I263875);
not I_15199 (I264125_rst,I5701);
nand I_15200 (I264142,I237577,I237556);
and I_15201 (I264159,I264142,I237553);
DFFARX1 I_15202  ( .D(I264159), .CLK(I5694_clk), .RSTB(I264125_rst), .Q(I264176) );
not I_15203 (I264193,I264176);
DFFARX1 I_15204  ( .D(I264176), .CLK(I5694_clk), .RSTB(I264125_rst), .Q(I264093) );
nor I_15205 (I264224,I237562,I237556);
DFFARX1 I_15206  ( .D(I237550), .CLK(I5694_clk), .RSTB(I264125_rst), .Q(I264241) );
DFFARX1 I_15207  ( .D(I264241), .CLK(I5694_clk), .RSTB(I264125_rst), .Q(I264258) );
not I_15208 (I264096,I264258);
DFFARX1 I_15209  ( .D(I264241), .CLK(I5694_clk), .RSTB(I264125_rst), .Q(I264289) );
and I_15210 (I264090,I264176,I264289);
nand I_15211 (I264320,I237580,I237571);
and I_15212 (I264337,I264320,I237568);
DFFARX1 I_15213  ( .D(I264337), .CLK(I5694_clk), .RSTB(I264125_rst), .Q(I264354) );
nor I_15214 (I264371,I264354,I264193);
not I_15215 (I264388,I264354);
nand I_15216 (I264099,I264176,I264388);
DFFARX1 I_15217  ( .D(I237565), .CLK(I5694_clk), .RSTB(I264125_rst), .Q(I264419) );
and I_15218 (I264436,I264419,I237574);
nor I_15219 (I264453,I264436,I264354);
nor I_15220 (I264470,I264436,I264388);
nand I_15221 (I264105,I264224,I264470);
not I_15222 (I264108,I264436);
DFFARX1 I_15223  ( .D(I264436), .CLK(I5694_clk), .RSTB(I264125_rst), .Q(I264087) );
DFFARX1 I_15224  ( .D(I237559), .CLK(I5694_clk), .RSTB(I264125_rst), .Q(I264529) );
nand I_15225 (I264546,I264529,I264241);
and I_15226 (I264563,I264224,I264546);
DFFARX1 I_15227  ( .D(I264563), .CLK(I5694_clk), .RSTB(I264125_rst), .Q(I264117) );
nor I_15228 (I264114,I264529,I264436);
and I_15229 (I264608,I264529,I264371);
or I_15230 (I264625,I264224,I264608);
DFFARX1 I_15231  ( .D(I264625), .CLK(I5694_clk), .RSTB(I264125_rst), .Q(I264102) );
nand I_15232 (I264111,I264529,I264453);
not I_15233 (I264703_rst,I5701);
nand I_15234 (I264720,I254990,I254987);
and I_15235 (I264737,I264720,I254999);
DFFARX1 I_15236  ( .D(I264737), .CLK(I5694_clk), .RSTB(I264703_rst), .Q(I264754) );
not I_15237 (I264771,I264754);
DFFARX1 I_15238  ( .D(I264754), .CLK(I5694_clk), .RSTB(I264703_rst), .Q(I264671) );
nor I_15239 (I264802,I254996,I254987);
DFFARX1 I_15240  ( .D(I255002), .CLK(I5694_clk), .RSTB(I264703_rst), .Q(I264819) );
DFFARX1 I_15241  ( .D(I264819), .CLK(I5694_clk), .RSTB(I264703_rst), .Q(I264836) );
not I_15242 (I264674,I264836);
DFFARX1 I_15243  ( .D(I264819), .CLK(I5694_clk), .RSTB(I264703_rst), .Q(I264867) );
and I_15244 (I264668,I264754,I264867);
nand I_15245 (I264898,I254978,I254981);
and I_15246 (I264915,I264898,I255005);
DFFARX1 I_15247  ( .D(I264915), .CLK(I5694_clk), .RSTB(I264703_rst), .Q(I264932) );
nor I_15248 (I264949,I264932,I264771);
not I_15249 (I264966,I264932);
nand I_15250 (I264677,I264754,I264966);
DFFARX1 I_15251  ( .D(I254984), .CLK(I5694_clk), .RSTB(I264703_rst), .Q(I264997) );
and I_15252 (I265014,I264997,I254975);
nor I_15253 (I265031,I265014,I264932);
nor I_15254 (I265048,I265014,I264966);
nand I_15255 (I264683,I264802,I265048);
not I_15256 (I264686,I265014);
DFFARX1 I_15257  ( .D(I265014), .CLK(I5694_clk), .RSTB(I264703_rst), .Q(I264665) );
DFFARX1 I_15258  ( .D(I254993), .CLK(I5694_clk), .RSTB(I264703_rst), .Q(I265107) );
nand I_15259 (I265124,I265107,I264819);
and I_15260 (I265141,I264802,I265124);
DFFARX1 I_15261  ( .D(I265141), .CLK(I5694_clk), .RSTB(I264703_rst), .Q(I264695) );
nor I_15262 (I264692,I265107,I265014);
and I_15263 (I265186,I265107,I264949);
or I_15264 (I265203,I264802,I265186);
DFFARX1 I_15265  ( .D(I265203), .CLK(I5694_clk), .RSTB(I264703_rst), .Q(I264680) );
nand I_15266 (I264689,I265107,I265031);
not I_15267 (I265281_rst,I5701);
nand I_15268 (I265298,I226821,I226836);
and I_15269 (I265315,I265298,I226824);
DFFARX1 I_15270  ( .D(I265315), .CLK(I5694_clk), .RSTB(I265281_rst), .Q(I265332) );
not I_15271 (I265349,I265332);
DFFARX1 I_15272  ( .D(I265332), .CLK(I5694_clk), .RSTB(I265281_rst), .Q(I265249) );
nor I_15273 (I265380,I226833,I226836);
DFFARX1 I_15274  ( .D(I226818), .CLK(I5694_clk), .RSTB(I265281_rst), .Q(I265397) );
DFFARX1 I_15275  ( .D(I265397), .CLK(I5694_clk), .RSTB(I265281_rst), .Q(I265414) );
not I_15276 (I265252,I265414);
DFFARX1 I_15277  ( .D(I265397), .CLK(I5694_clk), .RSTB(I265281_rst), .Q(I265445) );
and I_15278 (I265246,I265332,I265445);
nand I_15279 (I265476,I226809,I226806);
and I_15280 (I265493,I265476,I226812);
DFFARX1 I_15281  ( .D(I265493), .CLK(I5694_clk), .RSTB(I265281_rst), .Q(I265510) );
nor I_15282 (I265527,I265510,I265349);
not I_15283 (I265544,I265510);
nand I_15284 (I265255,I265332,I265544);
DFFARX1 I_15285  ( .D(I226815), .CLK(I5694_clk), .RSTB(I265281_rst), .Q(I265575) );
and I_15286 (I265592,I265575,I226827);
nor I_15287 (I265609,I265592,I265510);
nor I_15288 (I265626,I265592,I265544);
nand I_15289 (I265261,I265380,I265626);
not I_15290 (I265264,I265592);
DFFARX1 I_15291  ( .D(I265592), .CLK(I5694_clk), .RSTB(I265281_rst), .Q(I265243) );
DFFARX1 I_15292  ( .D(I226830), .CLK(I5694_clk), .RSTB(I265281_rst), .Q(I265685) );
nand I_15293 (I265702,I265685,I265397);
and I_15294 (I265719,I265380,I265702);
DFFARX1 I_15295  ( .D(I265719), .CLK(I5694_clk), .RSTB(I265281_rst), .Q(I265273) );
nor I_15296 (I265270,I265685,I265592);
and I_15297 (I265764,I265685,I265527);
or I_15298 (I265781,I265380,I265764);
DFFARX1 I_15299  ( .D(I265781), .CLK(I5694_clk), .RSTB(I265281_rst), .Q(I265258) );
nand I_15300 (I265267,I265685,I265609);
not I_15301 (I265859_rst,I5701);
nand I_15302 (I265876,I231740,I231722);
and I_15303 (I265893,I265876,I231734);
DFFARX1 I_15304  ( .D(I265893), .CLK(I5694_clk), .RSTB(I265859_rst), .Q(I265910) );
not I_15305 (I265927,I265910);
DFFARX1 I_15306  ( .D(I265910), .CLK(I5694_clk), .RSTB(I265859_rst), .Q(I265827) );
nor I_15307 (I265958,I231737,I231722);
DFFARX1 I_15308  ( .D(I231746), .CLK(I5694_clk), .RSTB(I265859_rst), .Q(I265975) );
DFFARX1 I_15309  ( .D(I265975), .CLK(I5694_clk), .RSTB(I265859_rst), .Q(I265992) );
not I_15310 (I265830,I265992);
DFFARX1 I_15311  ( .D(I265975), .CLK(I5694_clk), .RSTB(I265859_rst), .Q(I266023) );
and I_15312 (I265824,I265910,I266023);
nand I_15313 (I266054,I231725,I231749);
and I_15314 (I266071,I266054,I231728);
DFFARX1 I_15315  ( .D(I266071), .CLK(I5694_clk), .RSTB(I265859_rst), .Q(I266088) );
nor I_15316 (I266105,I266088,I265927);
not I_15317 (I266122,I266088);
nand I_15318 (I265833,I265910,I266122);
DFFARX1 I_15319  ( .D(I231731), .CLK(I5694_clk), .RSTB(I265859_rst), .Q(I266153) );
and I_15320 (I266170,I266153,I231743);
nor I_15321 (I266187,I266170,I266088);
nor I_15322 (I266204,I266170,I266122);
nand I_15323 (I265839,I265958,I266204);
not I_15324 (I26584_rst2,I266170);
DFFARX1 I_15325  ( .D(I266170), .CLK(I5694_clk), .RSTB(I265859_rst), .Q(I265821) );
DFFARX1 I_15326  ( .D(I231719), .CLK(I5694_clk), .RSTB(I265859_rst), .Q(I266263) );
nand I_15327 (I266280,I266263,I265975);
and I_15328 (I266297,I265958,I266280);
DFFARX1 I_15329  ( .D(I266297), .CLK(I5694_clk), .RSTB(I265859_rst), .Q(I265851) );
nor I_15330 (I26584_rst8,I266263,I266170);
and I_15331 (I266342,I266263,I266105);
or I_15332 (I266359,I265958,I266342);
DFFARX1 I_15333  ( .D(I266359), .CLK(I5694_clk), .RSTB(I265859_rst), .Q(I265836) );
nand I_15334 (I26584_rst5,I266263,I266187);
not I_15335 (I266437_rst,I5701);
nand I_15336 (I266454,I213709,I213697);
and I_15337 (I266471,I266454,I213691);
DFFARX1 I_15338  ( .D(I266471), .CLK(I5694_clk), .RSTB(I266437_rst), .Q(I266488) );
not I_15339 (I266505,I266488);
DFFARX1 I_15340  ( .D(I266488), .CLK(I5694_clk), .RSTB(I266437_rst), .Q(I266405) );
nor I_15341 (I266536,I213688,I213697);
DFFARX1 I_15342  ( .D(I213682), .CLK(I5694_clk), .RSTB(I266437_rst), .Q(I266553) );
DFFARX1 I_15343  ( .D(I266553), .CLK(I5694_clk), .RSTB(I266437_rst), .Q(I266570) );
not I_15344 (I266408,I266570);
DFFARX1 I_15345  ( .D(I266553), .CLK(I5694_clk), .RSTB(I266437_rst), .Q(I266601) );
and I_15346 (I266402,I266488,I266601);
nand I_15347 (I266632,I213685,I213700);
and I_15348 (I266649,I266632,I213712);
DFFARX1 I_15349  ( .D(I266649), .CLK(I5694_clk), .RSTB(I266437_rst), .Q(I266666) );
nor I_15350 (I266683,I266666,I266505);
not I_15351 (I266700,I266666);
nand I_15352 (I266411,I266488,I266700);
DFFARX1 I_15353  ( .D(I213703), .CLK(I5694_clk), .RSTB(I266437_rst), .Q(I266731) );
and I_15354 (I266748,I266731,I213694);
nor I_15355 (I266765,I266748,I266666);
nor I_15356 (I266782,I266748,I266700);
nand I_15357 (I266417,I266536,I266782);
not I_15358 (I266420,I266748);
DFFARX1 I_15359  ( .D(I266748), .CLK(I5694_clk), .RSTB(I266437_rst), .Q(I266399) );
DFFARX1 I_15360  ( .D(I213706), .CLK(I5694_clk), .RSTB(I266437_rst), .Q(I266841) );
nand I_15361 (I266858,I266841,I266553);
and I_15362 (I266875,I266536,I266858);
DFFARX1 I_15363  ( .D(I266875), .CLK(I5694_clk), .RSTB(I266437_rst), .Q(I266429) );
nor I_15364 (I266426,I266841,I266748);
and I_15365 (I266920,I266841,I266683);
or I_15366 (I266937,I266536,I266920);
DFFARX1 I_15367  ( .D(I266937), .CLK(I5694_clk), .RSTB(I266437_rst), .Q(I266414) );
nand I_15368 (I266423,I266841,I266765);
not I_15369 (I267015_rst,I5701);
nand I_15370 (I267032,I239557,I239569);
and I_15371 (I267049,I267032,I239548);
DFFARX1 I_15372  ( .D(I267049), .CLK(I5694_clk), .RSTB(I267015_rst), .Q(I267066) );
nor I_15373 (I267083,I239539,I239569);
nor I_15374 (I267100,I267083,I267066);
not I_15375 (I266998,I267083);
DFFARX1 I_15376  ( .D(I239551), .CLK(I5694_clk), .RSTB(I267015_rst), .Q(I267131) );
not I_15377 (I267148,I267131);
nor I_15378 (I267165,I267083,I267148);
nand I_15379 (I267001,I267131,I267100);
DFFARX1 I_15380  ( .D(I267131), .CLK(I5694_clk), .RSTB(I267015_rst), .Q(I266983) );
nand I_15381 (I267210,I239566,I239554);
and I_15382 (I267227,I267210,I239542);
DFFARX1 I_15383  ( .D(I267227), .CLK(I5694_clk), .RSTB(I267015_rst), .Q(I267244) );
nor I_15384 (I267004,I267244,I267066);
nand I_15385 (I266995,I267244,I267165);
DFFARX1 I_15386  ( .D(I239560), .CLK(I5694_clk), .RSTB(I267015_rst), .Q(I267289) );
and I_15387 (I267306,I267289,I239545);
DFFARX1 I_15388  ( .D(I267306), .CLK(I5694_clk), .RSTB(I267015_rst), .Q(I267323) );
not I_15389 (I266986,I267323);
nand I_15390 (I267354,I267306,I267244);
and I_15391 (I267371,I267066,I267354);
DFFARX1 I_15392  ( .D(I267371), .CLK(I5694_clk), .RSTB(I267015_rst), .Q(I266977) );
DFFARX1 I_15393  ( .D(I239563), .CLK(I5694_clk), .RSTB(I267015_rst), .Q(I267402) );
nand I_15394 (I267419,I267402,I267066);
and I_15395 (I267436,I267244,I267419);
DFFARX1 I_15396  ( .D(I267436), .CLK(I5694_clk), .RSTB(I267015_rst), .Q(I267007) );
not I_15397 (I267467,I267402);
nor I_15398 (I267484,I267083,I267467);
and I_15399 (I267501,I267402,I267484);
or I_15400 (I267518,I267306,I267501);
DFFARX1 I_15401  ( .D(I267518), .CLK(I5694_clk), .RSTB(I267015_rst), .Q(I266992) );
nand I_15402 (I266989,I267402,I267148);
DFFARX1 I_15403  ( .D(I267402), .CLK(I5694_clk), .RSTB(I267015_rst), .Q(I266980) );
not I_15404 (I267610_rst,I5701);
nand I_15405 (I267627,I261224,I261227);
and I_15406 (I267644,I267627,I261221);
DFFARX1 I_15407  ( .D(I267644), .CLK(I5694_clk), .RSTB(I267610_rst), .Q(I267661) );
nor I_15408 (I267678,I261218,I261227);
nor I_15409 (I267695,I267678,I267661);
not I_15410 (I267593,I267678);
DFFARX1 I_15411  ( .D(I261200), .CLK(I5694_clk), .RSTB(I267610_rst), .Q(I267726) );
not I_15412 (I267743,I267726);
nor I_15413 (I267760,I267678,I267743);
nand I_15414 (I267596,I267726,I267695);
DFFARX1 I_15415  ( .D(I267726), .CLK(I5694_clk), .RSTB(I267610_rst), .Q(I267578) );
nand I_15416 (I267805,I261209,I261206);
and I_15417 (I267822,I267805,I261215);
DFFARX1 I_15418  ( .D(I267822), .CLK(I5694_clk), .RSTB(I267610_rst), .Q(I267839) );
nor I_15419 (I267599,I267839,I267661);
nand I_15420 (I267590,I267839,I267760);
DFFARX1 I_15421  ( .D(I261197), .CLK(I5694_clk), .RSTB(I267610_rst), .Q(I267884) );
and I_15422 (I267901,I267884,I261212);
DFFARX1 I_15423  ( .D(I267901), .CLK(I5694_clk), .RSTB(I267610_rst), .Q(I267918) );
not I_15424 (I267581,I267918);
nand I_15425 (I267949,I267901,I267839);
and I_15426 (I267966,I267661,I267949);
DFFARX1 I_15427  ( .D(I267966), .CLK(I5694_clk), .RSTB(I267610_rst), .Q(I267572) );
DFFARX1 I_15428  ( .D(I261203), .CLK(I5694_clk), .RSTB(I267610_rst), .Q(I267997) );
nand I_15429 (I268014,I267997,I267661);
and I_15430 (I268031,I267839,I268014);
DFFARX1 I_15431  ( .D(I268031), .CLK(I5694_clk), .RSTB(I267610_rst), .Q(I267602) );
not I_15432 (I268062,I267997);
nor I_15433 (I268079,I267678,I268062);
and I_15434 (I268096,I267997,I268079);
or I_15435 (I268113,I267901,I268096);
DFFARX1 I_15436  ( .D(I268113), .CLK(I5694_clk), .RSTB(I267610_rst), .Q(I267587) );
nand I_15437 (I267584,I267997,I267743);
DFFARX1 I_15438  ( .D(I267997), .CLK(I5694_clk), .RSTB(I267610_rst), .Q(I267575) );
not I_15439 (I268205_rst,I5701);
nand I_15440 (I268222,I253055,I253067);
and I_15441 (I268239,I268222,I253049);
DFFARX1 I_15442  ( .D(I268239), .CLK(I5694_clk), .RSTB(I268205_rst), .Q(I268256) );
nor I_15443 (I268273,I253061,I253067);
nor I_15444 (I268290,I268273,I268256);
not I_15445 (I268188,I268273);
DFFARX1 I_15446  ( .D(I253046), .CLK(I5694_clk), .RSTB(I268205_rst), .Q(I268321) );
not I_15447 (I268338,I268321);
nor I_15448 (I268355,I268273,I268338);
nand I_15449 (I268191,I268321,I268290);
DFFARX1 I_15450  ( .D(I268321), .CLK(I5694_clk), .RSTB(I268205_rst), .Q(I268173) );
nand I_15451 (I268400,I253037,I253052);
and I_15452 (I268417,I268400,I253043);
DFFARX1 I_15453  ( .D(I268417), .CLK(I5694_clk), .RSTB(I268205_rst), .Q(I268434) );
nor I_15454 (I268194,I268434,I268256);
nand I_15455 (I268185,I268434,I268355);
DFFARX1 I_15456  ( .D(I253064), .CLK(I5694_clk), .RSTB(I268205_rst), .Q(I268479) );
and I_15457 (I268496,I268479,I253058);
DFFARX1 I_15458  ( .D(I268496), .CLK(I5694_clk), .RSTB(I268205_rst), .Q(I268513) );
not I_15459 (I268176,I268513);
nand I_15460 (I268544,I268496,I268434);
and I_15461 (I268561,I268256,I268544);
DFFARX1 I_15462  ( .D(I268561), .CLK(I5694_clk), .RSTB(I268205_rst), .Q(I268167) );
DFFARX1 I_15463  ( .D(I253040), .CLK(I5694_clk), .RSTB(I268205_rst), .Q(I268592) );
nand I_15464 (I268609,I268592,I268256);
and I_15465 (I268626,I268434,I268609);
DFFARX1 I_15466  ( .D(I268626), .CLK(I5694_clk), .RSTB(I268205_rst), .Q(I268197) );
not I_15467 (I268657,I268592);
nor I_15468 (I268674,I268273,I268657);
and I_15469 (I268691,I268592,I268674);
or I_15470 (I268708,I268496,I268691);
DFFARX1 I_15471  ( .D(I268708), .CLK(I5694_clk), .RSTB(I268205_rst), .Q(I268182) );
nand I_15472 (I268179,I268592,I268338);
DFFARX1 I_15473  ( .D(I268592), .CLK(I5694_clk), .RSTB(I268205_rst), .Q(I268170) );
not I_15474 (I268800_rst,I5701);
nand I_15475 (I268817,I238894,I238906);
and I_15476 (I268834,I268817,I238885);
DFFARX1 I_15477  ( .D(I268834), .CLK(I5694_clk), .RSTB(I268800_rst), .Q(I268851) );
nor I_15478 (I268868,I238876,I238906);
nor I_15479 (I268885,I268868,I268851);
not I_15480 (I268783,I268868);
DFFARX1 I_15481  ( .D(I238888), .CLK(I5694_clk), .RSTB(I268800_rst), .Q(I268916) );
not I_15482 (I268933,I268916);
nor I_15483 (I268950,I268868,I268933);
nand I_15484 (I268786,I268916,I268885);
DFFARX1 I_15485  ( .D(I268916), .CLK(I5694_clk), .RSTB(I268800_rst), .Q(I268768) );
nand I_15486 (I268995,I238903,I238891);
and I_15487 (I269012,I268995,I238879);
DFFARX1 I_15488  ( .D(I269012), .CLK(I5694_clk), .RSTB(I268800_rst), .Q(I269029) );
nor I_15489 (I268789,I269029,I268851);
nand I_15490 (I268780,I269029,I268950);
DFFARX1 I_15491  ( .D(I238897), .CLK(I5694_clk), .RSTB(I268800_rst), .Q(I269074) );
and I_15492 (I269091,I269074,I238882);
DFFARX1 I_15493  ( .D(I269091), .CLK(I5694_clk), .RSTB(I268800_rst), .Q(I269108) );
not I_15494 (I268771,I269108);
nand I_15495 (I269139,I269091,I269029);
and I_15496 (I269156,I268851,I269139);
DFFARX1 I_15497  ( .D(I269156), .CLK(I5694_clk), .RSTB(I268800_rst), .Q(I268762) );
DFFARX1 I_15498  ( .D(I238900), .CLK(I5694_clk), .RSTB(I268800_rst), .Q(I269187) );
nand I_15499 (I269204,I269187,I268851);
and I_15500 (I269221,I269029,I269204);
DFFARX1 I_15501  ( .D(I269221), .CLK(I5694_clk), .RSTB(I268800_rst), .Q(I268792) );
not I_15502 (I269252,I269187);
nor I_15503 (I269269,I268868,I269252);
and I_15504 (I269286,I269187,I269269);
or I_15505 (I269303,I269091,I269286);
DFFARX1 I_15506  ( .D(I269303), .CLK(I5694_clk), .RSTB(I268800_rst), .Q(I268777) );
nand I_15507 (I268774,I269187,I268933);
DFFARX1 I_15508  ( .D(I269187), .CLK(I5694_clk), .RSTB(I268800_rst), .Q(I268765) );
not I_15509 (I269395_rst,I5701);
nand I_15510 (I269412,I245116,I245122);
and I_15511 (I269429,I269412,I245104);
DFFARX1 I_15512  ( .D(I269429), .CLK(I5694_clk), .RSTB(I269395_rst), .Q(I269446) );
nor I_15513 (I269463,I245098,I245122);
nor I_15514 (I269480,I269463,I269446);
not I_15515 (I269378,I269463);
DFFARX1 I_15516  ( .D(I245128), .CLK(I5694_clk), .RSTB(I269395_rst), .Q(I269511) );
not I_15517 (I269528,I269511);
nor I_15518 (I269545,I269463,I269528);
nand I_15519 (I269381,I269511,I269480);
DFFARX1 I_15520  ( .D(I269511), .CLK(I5694_clk), .RSTB(I269395_rst), .Q(I269363) );
nand I_15521 (I269590,I245119,I245110);
and I_15522 (I269607,I269590,I245113);
DFFARX1 I_15523  ( .D(I269607), .CLK(I5694_clk), .RSTB(I269395_rst), .Q(I269624) );
nor I_15524 (I269384,I269624,I269446);
nand I_15525 (I269375,I269624,I269545);
DFFARX1 I_15526  ( .D(I245125), .CLK(I5694_clk), .RSTB(I269395_rst), .Q(I269669) );
and I_15527 (I269686,I269669,I245101);
DFFARX1 I_15528  ( .D(I269686), .CLK(I5694_clk), .RSTB(I269395_rst), .Q(I269703) );
not I_15529 (I269366,I269703);
nand I_15530 (I269734,I269686,I269624);
and I_15531 (I269751,I269446,I269734);
DFFARX1 I_15532  ( .D(I269751), .CLK(I5694_clk), .RSTB(I269395_rst), .Q(I269357) );
DFFARX1 I_15533  ( .D(I245107), .CLK(I5694_clk), .RSTB(I269395_rst), .Q(I269782) );
nand I_15534 (I269799,I269782,I269446);
and I_15535 (I269816,I269624,I269799);
DFFARX1 I_15536  ( .D(I269816), .CLK(I5694_clk), .RSTB(I269395_rst), .Q(I269387) );
not I_15537 (I269847,I269782);
nor I_15538 (I269864,I269463,I269847);
and I_15539 (I269881,I269782,I269864);
or I_15540 (I269898,I269686,I269881);
DFFARX1 I_15541  ( .D(I269898), .CLK(I5694_clk), .RSTB(I269395_rst), .Q(I269372) );
nand I_15542 (I269369,I269782,I269528);
DFFARX1 I_15543  ( .D(I269782), .CLK(I5694_clk), .RSTB(I269395_rst), .Q(I269360) );
not I_15544 (I269990_rst,I5701);
nand I_15545 (I270007,I264692,I264695);
and I_15546 (I270024,I270007,I264689);
DFFARX1 I_15547  ( .D(I270024), .CLK(I5694_clk), .RSTB(I269990_rst), .Q(I270041) );
nor I_15548 (I270058,I264686,I264695);
nor I_15549 (I270075,I270058,I270041);
not I_15550 (I269973,I270058);
DFFARX1 I_15551  ( .D(I264668), .CLK(I5694_clk), .RSTB(I269990_rst), .Q(I270106) );
not I_15552 (I270123,I270106);
nor I_15553 (I270140,I270058,I270123);
nand I_15554 (I269976,I270106,I270075);
DFFARX1 I_15555  ( .D(I270106), .CLK(I5694_clk), .RSTB(I269990_rst), .Q(I269958) );
nand I_15556 (I270185,I264677,I264674);
and I_15557 (I270202,I270185,I264683);
DFFARX1 I_15558  ( .D(I270202), .CLK(I5694_clk), .RSTB(I269990_rst), .Q(I270219) );
nor I_15559 (I269979,I270219,I270041);
nand I_15560 (I269970,I270219,I270140);
DFFARX1 I_15561  ( .D(I264665), .CLK(I5694_clk), .RSTB(I269990_rst), .Q(I270264) );
and I_15562 (I270281,I270264,I264680);
DFFARX1 I_15563  ( .D(I270281), .CLK(I5694_clk), .RSTB(I269990_rst), .Q(I270298) );
not I_15564 (I269961,I270298);
nand I_15565 (I270329,I270281,I270219);
and I_15566 (I270346,I270041,I270329);
DFFARX1 I_15567  ( .D(I270346), .CLK(I5694_clk), .RSTB(I269990_rst), .Q(I269952) );
DFFARX1 I_15568  ( .D(I264671), .CLK(I5694_clk), .RSTB(I269990_rst), .Q(I270377) );
nand I_15569 (I270394,I270377,I270041);
and I_15570 (I270411,I270219,I270394);
DFFARX1 I_15571  ( .D(I270411), .CLK(I5694_clk), .RSTB(I269990_rst), .Q(I269982) );
not I_15572 (I270442,I270377);
nor I_15573 (I270459,I270058,I270442);
and I_15574 (I270476,I270377,I270459);
or I_15575 (I270493,I270281,I270476);
DFFARX1 I_15576  ( .D(I270493), .CLK(I5694_clk), .RSTB(I269990_rst), .Q(I269967) );
nand I_15577 (I269964,I270377,I270123);
DFFARX1 I_15578  ( .D(I270377), .CLK(I5694_clk), .RSTB(I269990_rst), .Q(I269955) );
not I_15579 (I270585_rst,I5701);
nand I_15580 (I270602,I219123,I219114);
and I_15581 (I270619,I270602,I219132);
DFFARX1 I_15582  ( .D(I270619), .CLK(I5694_clk), .RSTB(I270585_rst), .Q(I270636) );
nor I_15583 (I270653,I219129,I219114);
nor I_15584 (I270670,I270653,I270636);
not I_15585 (I270568,I270653);
DFFARX1 I_15586  ( .D(I219111), .CLK(I5694_clk), .RSTB(I270585_rst), .Q(I270701) );
not I_15587 (I270718,I270701);
nor I_15588 (I270735,I270653,I270718);
nand I_15589 (I270571,I270701,I270670);
DFFARX1 I_15590  ( .D(I270701), .CLK(I5694_clk), .RSTB(I270585_rst), .Q(I270553) );
nand I_15591 (I270780,I219120,I219135);
and I_15592 (I270797,I270780,I219126);
DFFARX1 I_15593  ( .D(I270797), .CLK(I5694_clk), .RSTB(I270585_rst), .Q(I270814) );
nor I_15594 (I270574,I270814,I270636);
nand I_15595 (I270565,I270814,I270735);
DFFARX1 I_15596  ( .D(I219108), .CLK(I5694_clk), .RSTB(I270585_rst), .Q(I270859) );
and I_15597 (I270876,I270859,I219117);
DFFARX1 I_15598  ( .D(I270876), .CLK(I5694_clk), .RSTB(I270585_rst), .Q(I270893) );
not I_15599 (I270556,I270893);
nand I_15600 (I270924,I270876,I270814);
and I_15601 (I270941,I270636,I270924);
DFFARX1 I_15602  ( .D(I270941), .CLK(I5694_clk), .RSTB(I270585_rst), .Q(I270547) );
DFFARX1 I_15603  ( .D(I219105), .CLK(I5694_clk), .RSTB(I270585_rst), .Q(I270972) );
nand I_15604 (I270989,I270972,I270636);
and I_15605 (I271006,I270814,I270989);
DFFARX1 I_15606  ( .D(I271006), .CLK(I5694_clk), .RSTB(I270585_rst), .Q(I270577) );
not I_15607 (I271037,I270972);
nor I_15608 (I271054,I270653,I271037);
and I_15609 (I271071,I270972,I271054);
or I_15610 (I271088,I270876,I271071);
DFFARX1 I_15611  ( .D(I271088), .CLK(I5694_clk), .RSTB(I270585_rst), .Q(I270562) );
nand I_15612 (I270559,I270972,I270718);
DFFARX1 I_15613  ( .D(I270972), .CLK(I5694_clk), .RSTB(I270585_rst), .Q(I270550) );
not I_15614 (I271180_rst,I5701);
nand I_15615 (I271197,I227370,I227376);
and I_15616 (I271214,I271197,I227373);
DFFARX1 I_15617  ( .D(I271214), .CLK(I5694_clk), .RSTB(I271180_rst), .Q(I271231) );
nor I_15618 (I271248,I227397,I227376);
nor I_15619 (I271265,I271248,I271231);
not I_15620 (I271163,I271248);
DFFARX1 I_15621  ( .D(I227388), .CLK(I5694_clk), .RSTB(I271180_rst), .Q(I271296) );
not I_15622 (I271313,I271296);
nor I_15623 (I271330,I271248,I271313);
nand I_15624 (I271166,I271296,I271265);
DFFARX1 I_15625  ( .D(I271296), .CLK(I5694_clk), .RSTB(I271180_rst), .Q(I271148) );
nand I_15626 (I271375,I227391,I227394);
and I_15627 (I271392,I271375,I227367);
DFFARX1 I_15628  ( .D(I271392), .CLK(I5694_clk), .RSTB(I271180_rst), .Q(I271409) );
nor I_15629 (I271169,I271409,I271231);
nand I_15630 (I271160,I271409,I271330);
DFFARX1 I_15631  ( .D(I227385), .CLK(I5694_clk), .RSTB(I271180_rst), .Q(I271454) );
and I_15632 (I271471,I271454,I227379);
DFFARX1 I_15633  ( .D(I271471), .CLK(I5694_clk), .RSTB(I271180_rst), .Q(I271488) );
not I_15634 (I271151,I271488);
nand I_15635 (I271519,I271471,I271409);
and I_15636 (I271536,I271231,I271519);
DFFARX1 I_15637  ( .D(I271536), .CLK(I5694_clk), .RSTB(I271180_rst), .Q(I271142) );
DFFARX1 I_15638  ( .D(I227382), .CLK(I5694_clk), .RSTB(I271180_rst), .Q(I271567) );
nand I_15639 (I271584,I271567,I271231);
and I_15640 (I271601,I271409,I271584);
DFFARX1 I_15641  ( .D(I271601), .CLK(I5694_clk), .RSTB(I271180_rst), .Q(I271172) );
not I_15642 (I271632,I271567);
nor I_15643 (I271649,I271248,I271632);
and I_15644 (I271666,I271567,I271649);
or I_15645 (I271683,I271471,I271666);
DFFARX1 I_15646  ( .D(I271683), .CLK(I5694_clk), .RSTB(I271180_rst), .Q(I271157) );
nand I_15647 (I271154,I271567,I271313);
DFFARX1 I_15648  ( .D(I271567), .CLK(I5694_clk), .RSTB(I271180_rst), .Q(I271145) );
not I_15649 (I271775_rst,I5701);
nand I_15650 (I271792,I240812,I240809);
and I_15651 (I271809,I271792,I240806);
DFFARX1 I_15652  ( .D(I271809), .CLK(I5694_clk), .RSTB(I271775_rst), .Q(I271826) );
nor I_15653 (I271843,I240797,I240809);
nor I_15654 (I271860,I271843,I271826);
not I_15655 (I271758,I271843);
DFFARX1 I_15656  ( .D(I240815), .CLK(I5694_clk), .RSTB(I271775_rst), .Q(I271891) );
not I_15657 (I271908,I271891);
nor I_15658 (I271925,I271843,I271908);
nand I_15659 (I271761,I271891,I271860);
DFFARX1 I_15660  ( .D(I271891), .CLK(I5694_clk), .RSTB(I271775_rst), .Q(I271743) );
nand I_15661 (I271970,I240800,I240824);
and I_15662 (I271987,I271970,I240803);
DFFARX1 I_15663  ( .D(I271987), .CLK(I5694_clk), .RSTB(I271775_rst), .Q(I272004) );
nor I_15664 (I271764,I272004,I271826);
nand I_15665 (I271755,I272004,I271925);
DFFARX1 I_15666  ( .D(I240821), .CLK(I5694_clk), .RSTB(I271775_rst), .Q(I272049) );
and I_15667 (I272066,I272049,I240818);
DFFARX1 I_15668  ( .D(I272066), .CLK(I5694_clk), .RSTB(I271775_rst), .Q(I272083) );
not I_15669 (I271746,I272083);
nand I_15670 (I272114,I272066,I272004);
and I_15671 (I272131,I271826,I272114);
DFFARX1 I_15672  ( .D(I272131), .CLK(I5694_clk), .RSTB(I271775_rst), .Q(I271737) );
DFFARX1 I_15673  ( .D(I240827), .CLK(I5694_clk), .RSTB(I271775_rst), .Q(I272162) );
nand I_15674 (I272179,I272162,I271826);
and I_15675 (I272196,I272004,I272179);
DFFARX1 I_15676  ( .D(I272196), .CLK(I5694_clk), .RSTB(I271775_rst), .Q(I271767) );
not I_15677 (I272227,I272162);
nor I_15678 (I272244,I271843,I272227);
and I_15679 (I272261,I272162,I272244);
or I_15680 (I272278,I272066,I272261);
DFFARX1 I_15681  ( .D(I272278), .CLK(I5694_clk), .RSTB(I271775_rst), .Q(I271752) );
nand I_15682 (I271749,I272162,I271908);
DFFARX1 I_15683  ( .D(I272162), .CLK(I5694_clk), .RSTB(I271775_rst), .Q(I271740) );
not I_15684 (I272370_rst,I5701);
nand I_15685 (I272387,I243186,I243189);
and I_15686 (I272404,I272387,I243180);
DFFARX1 I_15687  ( .D(I272404), .CLK(I5694_clk), .RSTB(I272370_rst), .Q(I272421) );
nor I_15688 (I272438,I243204,I243189);
nor I_15689 (I272455,I272438,I272421);
not I_15690 (I272353,I272438);
DFFARX1 I_15691  ( .D(I243183), .CLK(I5694_clk), .RSTB(I272370_rst), .Q(I272486) );
not I_15692 (I272503,I272486);
nor I_15693 (I272520,I272438,I272503);
nand I_15694 (I272356,I272486,I272455);
DFFARX1 I_15695  ( .D(I272486), .CLK(I5694_clk), .RSTB(I272370_rst), .Q(I272338) );
nand I_15696 (I272565,I243201,I243192);
and I_15697 (I272582,I272565,I243177);
DFFARX1 I_15698  ( .D(I272582), .CLK(I5694_clk), .RSTB(I272370_rst), .Q(I272599) );
nor I_15699 (I272359,I272599,I272421);
nand I_15700 (I272350,I272599,I272520);
DFFARX1 I_15701  ( .D(I243207), .CLK(I5694_clk), .RSTB(I272370_rst), .Q(I272644) );
and I_15702 (I272661,I272644,I243198);
DFFARX1 I_15703  ( .D(I272661), .CLK(I5694_clk), .RSTB(I272370_rst), .Q(I272678) );
not I_15704 (I272341,I272678);
nand I_15705 (I272709,I272661,I272599);
and I_15706 (I272726,I272421,I272709);
DFFARX1 I_15707  ( .D(I272726), .CLK(I5694_clk), .RSTB(I272370_rst), .Q(I272332) );
DFFARX1 I_15708  ( .D(I243195), .CLK(I5694_clk), .RSTB(I272370_rst), .Q(I272757) );
nand I_15709 (I272774,I272757,I272421);
and I_15710 (I272791,I272599,I272774);
DFFARX1 I_15711  ( .D(I272791), .CLK(I5694_clk), .RSTB(I272370_rst), .Q(I272362) );
not I_15712 (I272822,I272757);
nor I_15713 (I272839,I272438,I272822);
and I_15714 (I272856,I272757,I272839);
or I_15715 (I272873,I272661,I272856);
DFFARX1 I_15716  ( .D(I272873), .CLK(I5694_clk), .RSTB(I272370_rst), .Q(I272347) );
nand I_15717 (I272344,I272757,I272503);
DFFARX1 I_15718  ( .D(I272757), .CLK(I5694_clk), .RSTB(I272370_rst), .Q(I272335) );
not I_15719 (I272965_rst,I5701);
nand I_15720 (I272982,I26584_rst8,I265851);
and I_15721 (I272999,I272982,I26584_rst5);
DFFARX1 I_15722  ( .D(I272999), .CLK(I5694_clk), .RSTB(I272965_rst), .Q(I273016) );
nor I_15723 (I273033,I26584_rst2,I265851);
nor I_15724 (I273050,I273033,I273016);
not I_15725 (I272948,I273033);
DFFARX1 I_15726  ( .D(I265824), .CLK(I5694_clk), .RSTB(I272965_rst), .Q(I273081) );
not I_15727 (I273098,I273081);
nor I_15728 (I273115,I273033,I273098);
nand I_15729 (I272951,I273081,I273050);
DFFARX1 I_15730  ( .D(I273081), .CLK(I5694_clk), .RSTB(I272965_rst), .Q(I272933) );
nand I_15731 (I273160,I265833,I265830);
and I_15732 (I273177,I273160,I265839);
DFFARX1 I_15733  ( .D(I273177), .CLK(I5694_clk), .RSTB(I272965_rst), .Q(I273194) );
nor I_15734 (I272954,I273194,I273016);
nand I_15735 (I272945,I273194,I273115);
DFFARX1 I_15736  ( .D(I265821), .CLK(I5694_clk), .RSTB(I272965_rst), .Q(I273239) );
and I_15737 (I273256,I273239,I265836);
DFFARX1 I_15738  ( .D(I273256), .CLK(I5694_clk), .RSTB(I272965_rst), .Q(I273273) );
not I_15739 (I272936,I273273);
nand I_15740 (I273304,I273256,I273194);
and I_15741 (I273321,I273016,I273304);
DFFARX1 I_15742  ( .D(I273321), .CLK(I5694_clk), .RSTB(I272965_rst), .Q(I272927) );
DFFARX1 I_15743  ( .D(I265827), .CLK(I5694_clk), .RSTB(I272965_rst), .Q(I273352) );
nand I_15744 (I273369,I273352,I273016);
and I_15745 (I273386,I273194,I273369);
DFFARX1 I_15746  ( .D(I273386), .CLK(I5694_clk), .RSTB(I272965_rst), .Q(I272957) );
not I_15747 (I273417,I273352);
nor I_15748 (I273434,I273033,I273417);
and I_15749 (I273451,I273352,I273434);
or I_15750 (I273468,I273256,I273451);
DFFARX1 I_15751  ( .D(I273468), .CLK(I5694_clk), .RSTB(I272965_rst), .Q(I272942) );
nand I_15752 (I272939,I273352,I273098);
DFFARX1 I_15753  ( .D(I273352), .CLK(I5694_clk), .RSTB(I272965_rst), .Q(I272930) );
not I_15754 (I273560_rst,I5701);
nand I_15755 (I273577,I260068,I260071);
and I_15756 (I273594,I273577,I260065);
DFFARX1 I_15757  ( .D(I273594), .CLK(I5694_clk), .RSTB(I273560_rst), .Q(I273611) );
nor I_15758 (I273628,I260062,I260071);
nor I_15759 (I273645,I273628,I273611);
not I_15760 (I273543,I273628);
DFFARX1 I_15761  ( .D(I260044), .CLK(I5694_clk), .RSTB(I273560_rst), .Q(I273676) );
not I_15762 (I273693,I273676);
nor I_15763 (I273710,I273628,I273693);
nand I_15764 (I273546,I273676,I273645);
DFFARX1 I_15765  ( .D(I273676), .CLK(I5694_clk), .RSTB(I273560_rst), .Q(I273528) );
nand I_15766 (I273755,I260053,I260050);
and I_15767 (I273772,I273755,I260059);
DFFARX1 I_15768  ( .D(I273772), .CLK(I5694_clk), .RSTB(I273560_rst), .Q(I273789) );
nor I_15769 (I273549,I273789,I273611);
nand I_15770 (I273540,I273789,I273710);
DFFARX1 I_15771  ( .D(I260041), .CLK(I5694_clk), .RSTB(I273560_rst), .Q(I273834) );
and I_15772 (I273851,I273834,I260056);
DFFARX1 I_15773  ( .D(I273851), .CLK(I5694_clk), .RSTB(I273560_rst), .Q(I273868) );
not I_15774 (I273531,I273868);
nand I_15775 (I273899,I273851,I273789);
and I_15776 (I273916,I273611,I273899);
DFFARX1 I_15777  ( .D(I273916), .CLK(I5694_clk), .RSTB(I273560_rst), .Q(I273522) );
DFFARX1 I_15778  ( .D(I260047), .CLK(I5694_clk), .RSTB(I273560_rst), .Q(I273947) );
nand I_15779 (I273964,I273947,I273611);
and I_15780 (I273981,I273789,I273964);
DFFARX1 I_15781  ( .D(I273981), .CLK(I5694_clk), .RSTB(I273560_rst), .Q(I273552) );
not I_15782 (I274012,I273947);
nor I_15783 (I274029,I273628,I274012);
and I_15784 (I274046,I273947,I274029);
or I_15785 (I274063,I273851,I274046);
DFFARX1 I_15786  ( .D(I274063), .CLK(I5694_clk), .RSTB(I273560_rst), .Q(I273537) );
nand I_15787 (I273534,I273947,I273693);
DFFARX1 I_15788  ( .D(I273947), .CLK(I5694_clk), .RSTB(I273560_rst), .Q(I273525) );
not I_15789 (I274155_rst,I5701);
nand I_15790 (I274172,I232374,I232386);
and I_15791 (I274189,I274172,I232395);
DFFARX1 I_15792  ( .D(I274189), .CLK(I5694_clk), .RSTB(I274155_rst), .Q(I274206) );
nor I_15793 (I274223,I232389,I232386);
nor I_15794 (I274240,I274223,I274206);
not I_15795 (I274138,I274223);
DFFARX1 I_15796  ( .D(I232383), .CLK(I5694_clk), .RSTB(I274155_rst), .Q(I274271) );
not I_15797 (I274288,I274271);
nor I_15798 (I274305,I274223,I274288);
nand I_15799 (I274141,I274271,I274240);
DFFARX1 I_15800  ( .D(I274271), .CLK(I5694_clk), .RSTB(I274155_rst), .Q(I274123) );
nand I_15801 (I274350,I232380,I232377);
and I_15802 (I274367,I274350,I232368);
DFFARX1 I_15803  ( .D(I274367), .CLK(I5694_clk), .RSTB(I274155_rst), .Q(I274384) );
nor I_15804 (I274144,I274384,I274206);
nand I_15805 (I274135,I274384,I274305);
DFFARX1 I_15806  ( .D(I232392), .CLK(I5694_clk), .RSTB(I274155_rst), .Q(I274429) );
and I_15807 (I274446,I274429,I232371);
DFFARX1 I_15808  ( .D(I274446), .CLK(I5694_clk), .RSTB(I274155_rst), .Q(I274463) );
not I_15809 (I274126,I274463);
nand I_15810 (I274494,I274446,I274384);
and I_15811 (I274511,I274206,I274494);
DFFARX1 I_15812  ( .D(I274511), .CLK(I5694_clk), .RSTB(I274155_rst), .Q(I274117) );
DFFARX1 I_15813  ( .D(I232365), .CLK(I5694_clk), .RSTB(I274155_rst), .Q(I274542) );
nand I_15814 (I274559,I274542,I274206);
and I_15815 (I274576,I274384,I274559);
DFFARX1 I_15816  ( .D(I274576), .CLK(I5694_clk), .RSTB(I274155_rst), .Q(I274147) );
not I_15817 (I274607,I274542);
nor I_15818 (I274624,I274223,I274607);
and I_15819 (I274641,I274542,I274624);
or I_15820 (I274658,I274446,I274641);
DFFARX1 I_15821  ( .D(I274658), .CLK(I5694_clk), .RSTB(I274155_rst), .Q(I274132) );
nand I_15822 (I274129,I274542,I274288);
DFFARX1 I_15823  ( .D(I274542), .CLK(I5694_clk), .RSTB(I274155_rst), .Q(I274120) );
not I_15824 (I274750_rst,I5701);
nand I_15825 (I274767,I242591,I242594);
and I_15826 (I274784,I274767,I242585);
DFFARX1 I_15827  ( .D(I274784), .CLK(I5694_clk), .RSTB(I274750_rst), .Q(I274801) );
nor I_15828 (I274818,I242609,I242594);
nor I_15829 (I274835,I274818,I274801);
not I_15830 (I274733,I274818);
DFFARX1 I_15831  ( .D(I242588), .CLK(I5694_clk), .RSTB(I274750_rst), .Q(I274866) );
not I_15832 (I274883,I274866);
nor I_15833 (I274900,I274818,I274883);
nand I_15834 (I274736,I274866,I274835);
DFFARX1 I_15835  ( .D(I274866), .CLK(I5694_clk), .RSTB(I274750_rst), .Q(I274718) );
nand I_15836 (I274945,I242606,I242597);
and I_15837 (I274962,I274945,I242582);
DFFARX1 I_15838  ( .D(I274962), .CLK(I5694_clk), .RSTB(I274750_rst), .Q(I274979) );
nor I_15839 (I274739,I274979,I274801);
nand I_15840 (I274730,I274979,I274900);
DFFARX1 I_15841  ( .D(I242612), .CLK(I5694_clk), .RSTB(I274750_rst), .Q(I275024) );
and I_15842 (I275041,I275024,I242603);
DFFARX1 I_15843  ( .D(I275041), .CLK(I5694_clk), .RSTB(I274750_rst), .Q(I275058) );
not I_15844 (I274721,I275058);
nand I_15845 (I275089,I275041,I274979);
and I_15846 (I275106,I274801,I275089);
DFFARX1 I_15847  ( .D(I275106), .CLK(I5694_clk), .RSTB(I274750_rst), .Q(I274712) );
DFFARX1 I_15848  ( .D(I242600), .CLK(I5694_clk), .RSTB(I274750_rst), .Q(I275137) );
nand I_15849 (I275154,I275137,I274801);
and I_15850 (I275171,I274979,I275154);
DFFARX1 I_15851  ( .D(I275171), .CLK(I5694_clk), .RSTB(I274750_rst), .Q(I274742) );
not I_15852 (I275202,I275137);
nor I_15853 (I275219,I274818,I275202);
and I_15854 (I275236,I275137,I275219);
or I_15855 (I275253,I275041,I275236);
DFFARX1 I_15856  ( .D(I275253), .CLK(I5694_clk), .RSTB(I274750_rst), .Q(I274727) );
nand I_15857 (I274724,I275137,I274883);
DFFARX1 I_15858  ( .D(I275137), .CLK(I5694_clk), .RSTB(I274750_rst), .Q(I274715) );
not I_15859 (I275345_rst,I5701);
nand I_15860 (I275362,I268777,I268762);
and I_15861 (I275379,I275362,I268768);
DFFARX1 I_15862  ( .D(I275379), .CLK(I5694_clk), .RSTB(I275345_rst), .Q(I275396) );
nor I_15863 (I275413,I268771,I268762);
DFFARX1 I_15864  ( .D(I268783), .CLK(I5694_clk), .RSTB(I275345_rst), .Q(I275430) );
nand I_15865 (I275447,I275430,I275413);
DFFARX1 I_15866  ( .D(I275430), .CLK(I5694_clk), .RSTB(I275345_rst), .Q(I275316) );
nand I_15867 (I275478,I268774,I268765);
and I_15868 (I275495,I275478,I268792);
DFFARX1 I_15869  ( .D(I275495), .CLK(I5694_clk), .RSTB(I275345_rst), .Q(I275512) );
not I_15870 (I275529,I275512);
nor I_15871 (I275546,I275396,I275529);
and I_15872 (I275563,I275413,I275546);
and I_15873 (I275580,I275512,I275447);
DFFARX1 I_15874  ( .D(I275580), .CLK(I5694_clk), .RSTB(I275345_rst), .Q(I275313) );
DFFARX1 I_15875  ( .D(I275512), .CLK(I5694_clk), .RSTB(I275345_rst), .Q(I275307) );
DFFARX1 I_15876  ( .D(I268780), .CLK(I5694_clk), .RSTB(I275345_rst), .Q(I275625) );
and I_15877 (I275642,I275625,I268786);
nand I_15878 (I275659,I275642,I275512);
nor I_15879 (I275334,I275642,I275413);
not I_15880 (I275690,I275642);
nor I_15881 (I275707,I275396,I275690);
nand I_15882 (I275325,I275430,I275707);
nand I_15883 (I275319,I275512,I275690);
or I_15884 (I275752,I275642,I275563);
DFFARX1 I_15885  ( .D(I275752), .CLK(I5694_clk), .RSTB(I275345_rst), .Q(I275322) );
DFFARX1 I_15886  ( .D(I268789), .CLK(I5694_clk), .RSTB(I275345_rst), .Q(I275783) );
and I_15887 (I275800,I275783,I275659);
DFFARX1 I_15888  ( .D(I275800), .CLK(I5694_clk), .RSTB(I275345_rst), .Q(I275337) );
nor I_15889 (I275831,I275783,I275396);
nand I_15890 (I275331,I275642,I275831);
not I_15891 (I275328,I275783);
DFFARX1 I_15892  ( .D(I275783), .CLK(I5694_clk), .RSTB(I275345_rst), .Q(I275876) );
and I_15893 (I275310,I275783,I275876);
not I_15894 (I275940_rst,I5701);
nand I_15895 (I275957,I226248,I226263);
and I_15896 (I275974,I275957,I226269);
DFFARX1 I_15897  ( .D(I275974), .CLK(I5694_clk), .RSTB(I275940_rst), .Q(I275991) );
nor I_15898 (I276008,I226257,I226263);
DFFARX1 I_15899  ( .D(I226245), .CLK(I5694_clk), .RSTB(I275940_rst), .Q(I276025) );
nand I_15900 (I276042,I276025,I276008);
DFFARX1 I_15901  ( .D(I276025), .CLK(I5694_clk), .RSTB(I275940_rst), .Q(I275911) );
nand I_15902 (I276073,I226251,I226254);
and I_15903 (I276090,I276073,I226260);
DFFARX1 I_15904  ( .D(I276090), .CLK(I5694_clk), .RSTB(I275940_rst), .Q(I276107) );
not I_15905 (I276124,I276107);
nor I_15906 (I276141,I275991,I276124);
and I_15907 (I276158,I276008,I276141);
and I_15908 (I276175,I276107,I276042);
DFFARX1 I_15909  ( .D(I276175), .CLK(I5694_clk), .RSTB(I275940_rst), .Q(I275908) );
DFFARX1 I_15910  ( .D(I276107), .CLK(I5694_clk), .RSTB(I275940_rst), .Q(I275902) );
DFFARX1 I_15911  ( .D(I226266), .CLK(I5694_clk), .RSTB(I275940_rst), .Q(I276220) );
and I_15912 (I276237,I276220,I226275);
nand I_15913 (I276254,I276237,I276107);
nor I_15914 (I275929,I276237,I276008);
not I_15915 (I276285,I276237);
nor I_15916 (I276302,I275991,I276285);
nand I_15917 (I275920,I276025,I276302);
nand I_15918 (I275914,I276107,I276285);
or I_15919 (I276347,I276237,I276158);
DFFARX1 I_15920  ( .D(I276347), .CLK(I5694_clk), .RSTB(I275940_rst), .Q(I275917) );
DFFARX1 I_15921  ( .D(I226272), .CLK(I5694_clk), .RSTB(I275940_rst), .Q(I276378) );
and I_15922 (I276395,I276378,I276254);
DFFARX1 I_15923  ( .D(I276395), .CLK(I5694_clk), .RSTB(I275940_rst), .Q(I275932) );
nor I_15924 (I276426,I276378,I275991);
nand I_15925 (I275926,I276237,I276426);
not I_15926 (I275923,I276378);
DFFARX1 I_15927  ( .D(I276378), .CLK(I5694_clk), .RSTB(I275940_rst), .Q(I276471) );
and I_15928 (I275905,I276378,I276471);
not I_15929 (I276535_rst,I5701);
nand I_15930 (I276552,I221621,I221624);
and I_15931 (I276569,I276552,I221633);
DFFARX1 I_15932  ( .D(I276569), .CLK(I5694_clk), .RSTB(I276535_rst), .Q(I276586) );
nor I_15933 (I276603,I221627,I221624);
DFFARX1 I_15934  ( .D(I221648), .CLK(I5694_clk), .RSTB(I276535_rst), .Q(I276620) );
nand I_15935 (I276637,I276620,I276603);
DFFARX1 I_15936  ( .D(I276620), .CLK(I5694_clk), .RSTB(I276535_rst), .Q(I276506) );
nand I_15937 (I276668,I221645,I221651);
and I_15938 (I276685,I276668,I221636);
DFFARX1 I_15939  ( .D(I276685), .CLK(I5694_clk), .RSTB(I276535_rst), .Q(I276702) );
not I_15940 (I276719,I276702);
nor I_15941 (I276736,I276586,I276719);
and I_15942 (I276753,I276603,I276736);
and I_15943 (I276770,I276702,I276637);
DFFARX1 I_15944  ( .D(I276770), .CLK(I5694_clk), .RSTB(I276535_rst), .Q(I276503) );
DFFARX1 I_15945  ( .D(I276702), .CLK(I5694_clk), .RSTB(I276535_rst), .Q(I276497) );
DFFARX1 I_15946  ( .D(I221639), .CLK(I5694_clk), .RSTB(I276535_rst), .Q(I276815) );
and I_15947 (I276832,I276815,I221642);
nand I_15948 (I276849,I276832,I276702);
nor I_15949 (I276524,I276832,I276603);
not I_15950 (I276880,I276832);
nor I_15951 (I276897,I276586,I276880);
nand I_15952 (I276515,I276620,I276897);
nand I_15953 (I276509,I276702,I276880);
or I_15954 (I276942,I276832,I276753);
DFFARX1 I_15955  ( .D(I276942), .CLK(I5694_clk), .RSTB(I276535_rst), .Q(I276512) );
DFFARX1 I_15956  ( .D(I221630), .CLK(I5694_clk), .RSTB(I276535_rst), .Q(I276973) );
and I_15957 (I276990,I276973,I276849);
DFFARX1 I_15958  ( .D(I276990), .CLK(I5694_clk), .RSTB(I276535_rst), .Q(I276527) );
nor I_15959 (I277021,I276973,I276586);
nand I_15960 (I276521,I276832,I277021);
not I_15961 (I276518,I276973);
DFFARX1 I_15962  ( .D(I276973), .CLK(I5694_clk), .RSTB(I276535_rst), .Q(I277066) );
and I_15963 (I276500,I276973,I277066);
not I_15964 (I277130_rst,I5701);
nand I_15965 (I277147,I251095,I251065);
and I_15966 (I277164,I277147,I251083);
DFFARX1 I_15967  ( .D(I277164), .CLK(I5694_clk), .RSTB(I277130_rst), .Q(I277181) );
nor I_15968 (I277198,I251077,I251065);
DFFARX1 I_15969  ( .D(I251074), .CLK(I5694_clk), .RSTB(I277130_rst), .Q(I277215) );
nand I_15970 (I277232,I277215,I277198);
DFFARX1 I_15971  ( .D(I277215), .CLK(I5694_clk), .RSTB(I277130_rst), .Q(I277101) );
nand I_15972 (I277263,I251068,I251071);
and I_15973 (I277280,I277263,I251089);
DFFARX1 I_15974  ( .D(I277280), .CLK(I5694_clk), .RSTB(I277130_rst), .Q(I277297) );
not I_15975 (I277314,I277297);
nor I_15976 (I277331,I277181,I277314);
and I_15977 (I277348,I277198,I277331);
and I_15978 (I277365,I277297,I277232);
DFFARX1 I_15979  ( .D(I277365), .CLK(I5694_clk), .RSTB(I277130_rst), .Q(I277098) );
DFFARX1 I_15980  ( .D(I277297), .CLK(I5694_clk), .RSTB(I277130_rst), .Q(I277092) );
DFFARX1 I_15981  ( .D(I251092), .CLK(I5694_clk), .RSTB(I277130_rst), .Q(I277410) );
and I_15982 (I277427,I277410,I251086);
nand I_15983 (I277444,I277427,I277297);
nor I_15984 (I277119,I277427,I277198);
not I_15985 (I277475,I277427);
nor I_15986 (I277492,I277181,I277475);
nand I_15987 (I277110,I277215,I277492);
nand I_15988 (I277104,I277297,I277475);
or I_15989 (I277537,I277427,I277348);
DFFARX1 I_15990  ( .D(I277537), .CLK(I5694_clk), .RSTB(I277130_rst), .Q(I277107) );
DFFARX1 I_15991  ( .D(I251080), .CLK(I5694_clk), .RSTB(I277130_rst), .Q(I277568) );
and I_15992 (I277585,I277568,I277444);
DFFARX1 I_15993  ( .D(I277585), .CLK(I5694_clk), .RSTB(I277130_rst), .Q(I277122) );
nor I_15994 (I277616,I277568,I277181);
nand I_15995 (I277116,I277427,I277616);
not I_15996 (I277113,I277568);
DFFARX1 I_15997  ( .D(I277568), .CLK(I5694_clk), .RSTB(I277130_rst), .Q(I277661) );
and I_15998 (I277095,I277568,I277661);
not I_15999 (I277725_rst,I5701);
nand I_16000 (I277742,I251758,I251728);
and I_16001 (I277759,I277742,I251746);
DFFARX1 I_16002  ( .D(I277759), .CLK(I5694_clk), .RSTB(I277725_rst), .Q(I277776) );
nor I_16003 (I277793,I251740,I251728);
DFFARX1 I_16004  ( .D(I251737), .CLK(I5694_clk), .RSTB(I277725_rst), .Q(I277810) );
nand I_16005 (I277827,I277810,I277793);
DFFARX1 I_16006  ( .D(I277810), .CLK(I5694_clk), .RSTB(I277725_rst), .Q(I277696) );
nand I_16007 (I277858,I251731,I251734);
and I_16008 (I277875,I277858,I251752);
DFFARX1 I_16009  ( .D(I277875), .CLK(I5694_clk), .RSTB(I277725_rst), .Q(I277892) );
not I_16010 (I277909,I277892);
nor I_16011 (I277926,I277776,I277909);
and I_16012 (I277943,I277793,I277926);
and I_16013 (I277960,I277892,I277827);
DFFARX1 I_16014  ( .D(I277960), .CLK(I5694_clk), .RSTB(I277725_rst), .Q(I277693) );
DFFARX1 I_16015  ( .D(I277892), .CLK(I5694_clk), .RSTB(I277725_rst), .Q(I277687) );
DFFARX1 I_16016  ( .D(I251755), .CLK(I5694_clk), .RSTB(I277725_rst), .Q(I278005) );
and I_16017 (I278022,I278005,I251749);
nand I_16018 (I278039,I278022,I277892);
nor I_16019 (I277714,I278022,I277793);
not I_16020 (I278070,I278022);
nor I_16021 (I278087,I277776,I278070);
nand I_16022 (I277705,I277810,I278087);
nand I_16023 (I277699,I277892,I278070);
or I_16024 (I278132,I278022,I277943);
DFFARX1 I_16025  ( .D(I278132), .CLK(I5694_clk), .RSTB(I277725_rst), .Q(I277702) );
DFFARX1 I_16026  ( .D(I251743), .CLK(I5694_clk), .RSTB(I277725_rst), .Q(I278163) );
and I_16027 (I278180,I278163,I278039);
DFFARX1 I_16028  ( .D(I278180), .CLK(I5694_clk), .RSTB(I277725_rst), .Q(I277717) );
nor I_16029 (I278211,I278163,I277776);
nand I_16030 (I277711,I278022,I278211);
not I_16031 (I277708,I278163);
DFFARX1 I_16032  ( .D(I278163), .CLK(I5694_clk), .RSTB(I277725_rst), .Q(I278256) );
and I_16033 (I277690,I278163,I278256);
not I_16034 (I278320_rst,I5701);
nand I_16035 (I278337,I222199,I222202);
and I_16036 (I278354,I278337,I222211);
DFFARX1 I_16037  ( .D(I278354), .CLK(I5694_clk), .RSTB(I278320_rst), .Q(I278371) );
nor I_16038 (I278388,I222205,I222202);
DFFARX1 I_16039  ( .D(I222226), .CLK(I5694_clk), .RSTB(I278320_rst), .Q(I278405) );
nand I_16040 (I278422,I278405,I278388);
DFFARX1 I_16041  ( .D(I278405), .CLK(I5694_clk), .RSTB(I278320_rst), .Q(I278291) );
nand I_16042 (I278453,I222223,I222229);
and I_16043 (I278470,I278453,I222214);
DFFARX1 I_16044  ( .D(I278470), .CLK(I5694_clk), .RSTB(I278320_rst), .Q(I278487) );
not I_16045 (I278504,I278487);
nor I_16046 (I278521,I278371,I278504);
and I_16047 (I278538,I278388,I278521);
and I_16048 (I278555,I278487,I278422);
DFFARX1 I_16049  ( .D(I278555), .CLK(I5694_clk), .RSTB(I278320_rst), .Q(I278288) );
DFFARX1 I_16050  ( .D(I278487), .CLK(I5694_clk), .RSTB(I278320_rst), .Q(I278282) );
DFFARX1 I_16051  ( .D(I222217), .CLK(I5694_clk), .RSTB(I278320_rst), .Q(I278600) );
and I_16052 (I278617,I278600,I222220);
nand I_16053 (I278634,I278617,I278487);
nor I_16054 (I278309,I278617,I278388);
not I_16055 (I278665,I278617);
nor I_16056 (I278682,I278371,I278665);
nand I_16057 (I278300,I278405,I278682);
nand I_16058 (I278294,I278487,I278665);
or I_16059 (I278727,I278617,I278538);
DFFARX1 I_16060  ( .D(I278727), .CLK(I5694_clk), .RSTB(I278320_rst), .Q(I278297) );
DFFARX1 I_16061  ( .D(I222208), .CLK(I5694_clk), .RSTB(I278320_rst), .Q(I278758) );
and I_16062 (I278775,I278758,I278634);
DFFARX1 I_16063  ( .D(I278775), .CLK(I5694_clk), .RSTB(I278320_rst), .Q(I278312) );
nor I_16064 (I278806,I278758,I278371);
nand I_16065 (I278306,I278617,I278806);
not I_16066 (I278303,I278758);
DFFARX1 I_16067  ( .D(I278758), .CLK(I5694_clk), .RSTB(I278320_rst), .Q(I278851) );
and I_16068 (I278285,I278758,I278851);
not I_16069 (I278915_rst,I5701);
not I_16070 (I278932,I238225);
nor I_16071 (I278949,I238216,I238240);
nand I_16072 (I278966,I278949,I238243);
nor I_16073 (I278983,I278932,I238216);
nand I_16074 (I279000,I278983,I238234);
not I_16075 (I279017,I238216);
not I_16076 (I279034,I279017);
not I_16077 (I279051,I238228);
nor I_16078 (I279068,I279051,I238222);
and I_16079 (I279085,I279068,I238231);
or I_16080 (I279102,I279085,I238219);
DFFARX1 I_16081  ( .D(I279102), .CLK(I5694_clk), .RSTB(I278915_rst), .Q(I279119) );
nand I_16082 (I279136,I278932,I238228);
or I_16083 (I278904,I279136,I279119);
not I_16084 (I279167,I279136);
nor I_16085 (I279184,I279119,I279167);
and I_16086 (I279201,I279017,I279184);
nand I_16087 (I278877,I279136,I279034);
DFFARX1 I_16088  ( .D(I238213), .CLK(I5694_clk), .RSTB(I278915_rst), .Q(I279232) );
or I_16089 (I278898,I279232,I279119);
nor I_16090 (I279263,I279232,I279000);
nor I_16091 (I279280,I279232,I279034);
nand I_16092 (I278883,I278966,I279280);
or I_16093 (I279311,I279232,I279201);
DFFARX1 I_16094  ( .D(I279311), .CLK(I5694_clk), .RSTB(I278915_rst), .Q(I278880) );
not I_16095 (I278886,I279232);
DFFARX1 I_16096  ( .D(I238237), .CLK(I5694_clk), .RSTB(I278915_rst), .Q(I279356) );
not I_16097 (I279373,I279356);
nor I_16098 (I279390,I279373,I278966);
DFFARX1 I_16099  ( .D(I279390), .CLK(I5694_clk), .RSTB(I278915_rst), .Q(I278892) );
nor I_16100 (I278907,I279232,I279373);
nor I_16101 (I278895,I279373,I279136);
not I_16102 (I279449,I279373);
and I_16103 (I279466,I279000,I279449);
nor I_16104 (I278901,I279136,I279466);
nand I_16105 (I278889,I279373,I279263);
not I_16106 (I279544_rst,I5701);
not I_16107 (I279561,I223939);
nor I_16108 (I279578,I223963,I223948);
nand I_16109 (I279595,I279578,I223933);
nor I_16110 (I279612,I279561,I223963);
nand I_16111 (I279629,I279612,I223960);
not I_16112 (I279646,I223963);
not I_16113 (I279663,I279646);
not I_16114 (I279680,I223942);
nor I_16115 (I279697,I279680,I223936);
and I_16116 (I279714,I279697,I223957);
or I_16117 (I279731,I279714,I223945);
DFFARX1 I_16118  ( .D(I279731), .CLK(I5694_clk), .RSTB(I279544_rst), .Q(I279748) );
nand I_16119 (I279765,I279561,I223942);
or I_16120 (I279533,I279765,I279748);
not I_16121 (I279796,I279765);
nor I_16122 (I279813,I279748,I279796);
and I_16123 (I279830,I279646,I279813);
nand I_16124 (I279506,I279765,I279663);
DFFARX1 I_16125  ( .D(I223954), .CLK(I5694_clk), .RSTB(I279544_rst), .Q(I279861) );
or I_16126 (I279527,I279861,I279748);
nor I_16127 (I279892,I279861,I279629);
nor I_16128 (I279909,I279861,I279663);
nand I_16129 (I279512,I279595,I279909);
or I_16130 (I279940,I279861,I279830);
DFFARX1 I_16131  ( .D(I279940), .CLK(I5694_clk), .RSTB(I279544_rst), .Q(I279509) );
not I_16132 (I279515,I279861);
DFFARX1 I_16133  ( .D(I223951), .CLK(I5694_clk), .RSTB(I279544_rst), .Q(I279985) );
not I_16134 (I280002,I279985);
nor I_16135 (I280019,I280002,I279595);
DFFARX1 I_16136  ( .D(I280019), .CLK(I5694_clk), .RSTB(I279544_rst), .Q(I279521) );
nor I_16137 (I279536,I279861,I280002);
nor I_16138 (I279524,I280002,I279765);
not I_16139 (I280078,I280002);
and I_16140 (I280095,I279629,I280078);
nor I_16141 (I279530,I279765,I280095);
nand I_16142 (I279518,I280002,I279892);
not I_16143 (I280173_rst,I5701);
not I_16144 (I280190,I233663);
nor I_16145 (I280207,I233681,I233660);
nand I_16146 (I280224,I280207,I233678);
nor I_16147 (I280241,I280190,I233681);
nand I_16148 (I280258,I280241,I233672);
not I_16149 (I280275,I233681);
not I_16150 (I280292,I280275);
not I_16151 (I280309,I233675);
nor I_16152 (I280326,I280309,I233669);
and I_16153 (I280343,I280326,I233666);
or I_16154 (I280360,I280343,I233657);
DFFARX1 I_16155  ( .D(I280360), .CLK(I5694_clk), .RSTB(I280173_rst), .Q(I280377) );
nand I_16156 (I280394,I280190,I233675);
or I_16157 (I280162,I280394,I280377);
not I_16158 (I280425,I280394);
nor I_16159 (I280442,I280377,I280425);
and I_16160 (I280459,I280275,I280442);
nand I_16161 (I280135,I280394,I280292);
DFFARX1 I_16162  ( .D(I233687), .CLK(I5694_clk), .RSTB(I280173_rst), .Q(I280490) );
or I_16163 (I280156,I280490,I280377);
nor I_16164 (I280521,I280490,I280258);
nor I_16165 (I280538,I280490,I280292);
nand I_16166 (I280141,I280224,I280538);
or I_16167 (I280569,I280490,I280459);
DFFARX1 I_16168  ( .D(I280569), .CLK(I5694_clk), .RSTB(I280173_rst), .Q(I280138) );
not I_16169 (I280144,I280490);
DFFARX1 I_16170  ( .D(I233684), .CLK(I5694_clk), .RSTB(I280173_rst), .Q(I280614) );
not I_16171 (I280631,I280614);
nor I_16172 (I280648,I280631,I280224);
DFFARX1 I_16173  ( .D(I280648), .CLK(I5694_clk), .RSTB(I280173_rst), .Q(I280150) );
nor I_16174 (I280165,I280490,I280631);
nor I_16175 (I280153,I280631,I280394);
not I_16176 (I280707,I280631);
and I_16177 (I280724,I280258,I280707);
nor I_16178 (I280159,I280394,I280724);
nand I_16179 (I280147,I280631,I280521);
not I_16180 (I280802_rst,I5701);
not I_16181 (I280819,I264117);
nor I_16182 (I280836,I264090,I264108);
nand I_16183 (I280853,I280836,I264093);
nor I_16184 (I280870,I280819,I264090);
nand I_16185 (I280887,I280870,I264111);
not I_16186 (I280904,I264090);
not I_16187 (I280921,I280904);
not I_16188 (I280938,I264087);
nor I_16189 (I280955,I280938,I264114);
and I_16190 (I280972,I280955,I264105);
or I_16191 (I280989,I280972,I264096);
DFFARX1 I_16192  ( .D(I280989), .CLK(I5694_clk), .RSTB(I280802_rst), .Q(I281006) );
nand I_16193 (I281023,I280819,I264087);
or I_16194 (I280791,I281023,I281006);
not I_16195 (I281054,I281023);
nor I_16196 (I281071,I281006,I281054);
and I_16197 (I281088,I280904,I281071);
nand I_16198 (I280764,I281023,I280921);
DFFARX1 I_16199  ( .D(I264099), .CLK(I5694_clk), .RSTB(I280802_rst), .Q(I281119) );
or I_16200 (I280785,I281119,I281006);
nor I_16201 (I281150,I281119,I280887);
nor I_16202 (I281167,I281119,I280921);
nand I_16203 (I280770,I280853,I281167);
or I_16204 (I281198,I281119,I281088);
DFFARX1 I_16205  ( .D(I281198), .CLK(I5694_clk), .RSTB(I280802_rst), .Q(I280767) );
not I_16206 (I280773,I281119);
DFFARX1 I_16207  ( .D(I264102), .CLK(I5694_clk), .RSTB(I280802_rst), .Q(I281243) );
not I_16208 (I281260,I281243);
nor I_16209 (I281277,I281260,I280853);
DFFARX1 I_16210  ( .D(I281277), .CLK(I5694_clk), .RSTB(I280802_rst), .Q(I280779) );
nor I_16211 (I280794,I281119,I281260);
nor I_16212 (I280782,I281260,I281023);
not I_16213 (I281336,I281260);
and I_16214 (I281353,I280887,I281336);
nor I_16215 (I280788,I281023,I281353);
nand I_16216 (I280776,I281260,I281150);
not I_16217 (I281431_rst,I5701);
not I_16218 (I281448,I231079);
nor I_16219 (I281465,I231097,I231076);
nand I_16220 (I281482,I281465,I231094);
nor I_16221 (I281499,I281448,I231097);
nand I_16222 (I281516,I281499,I231088);
not I_16223 (I281533,I231097);
not I_16224 (I281550,I281533);
not I_16225 (I281567,I231091);
nor I_16226 (I281584,I281567,I231085);
and I_16227 (I281601,I281584,I231082);
or I_16228 (I281618,I281601,I231073);
DFFARX1 I_16229  ( .D(I281618), .CLK(I5694_clk), .RSTB(I281431_rst), .Q(I281635) );
nand I_16230 (I281652,I281448,I231091);
or I_16231 (I281420,I281652,I281635);
not I_16232 (I281683,I281652);
nor I_16233 (I281700,I281635,I281683);
and I_16234 (I281717,I281533,I281700);
nand I_16235 (I281393,I281652,I281550);
DFFARX1 I_16236  ( .D(I231103), .CLK(I5694_clk), .RSTB(I281431_rst), .Q(I281748) );
or I_16237 (I281414,I281748,I281635);
nor I_16238 (I281779,I281748,I281516);
nor I_16239 (I281796,I281748,I281550);
nand I_16240 (I281399,I281482,I281796);
or I_16241 (I281827,I281748,I281717);
DFFARX1 I_16242  ( .D(I281827), .CLK(I5694_clk), .RSTB(I281431_rst), .Q(I281396) );
not I_16243 (I281402,I281748);
DFFARX1 I_16244  ( .D(I231100), .CLK(I5694_clk), .RSTB(I281431_rst), .Q(I281872) );
not I_16245 (I281889,I281872);
nor I_16246 (I281906,I281889,I281482);
DFFARX1 I_16247  ( .D(I281906), .CLK(I5694_clk), .RSTB(I281431_rst), .Q(I281408) );
nor I_16248 (I281423,I281748,I281889);
nor I_16249 (I281411,I281889,I281652);
not I_16250 (I281965,I281889);
and I_16251 (I281982,I281516,I281965);
nor I_16252 (I281417,I281652,I281982);
nand I_16253 (I281405,I281889,I281779);
not I_16254 (I282060_rst,I5701);
not I_16255 (I282077,I269958);
nor I_16256 (I282094,I269976,I269955);
nand I_16257 (I282111,I282094,I269979);
nor I_16258 (I282128,I282077,I269976);
nand I_16259 (I282145,I282128,I269973);
not I_16260 (I282162,I269976);
not I_16261 (I282179,I282162);
not I_16262 (I282196,I269964);
nor I_16263 (I282213,I282196,I269952);
and I_16264 (I282230,I282213,I269970);
or I_16265 (I282247,I282230,I269982);
DFFARX1 I_16266  ( .D(I282247), .CLK(I5694_clk), .RSTB(I282060_rst), .Q(I282264) );
nand I_16267 (I282281,I282077,I269964);
or I_16268 (I282049,I282281,I282264);
not I_16269 (I282312,I282281);
nor I_16270 (I282329,I282264,I282312);
and I_16271 (I282346,I282162,I282329);
nand I_16272 (I282022,I282281,I282179);
DFFARX1 I_16273  ( .D(I269961), .CLK(I5694_clk), .RSTB(I282060_rst), .Q(I282377) );
or I_16274 (I282043,I282377,I282264);
nor I_16275 (I282408,I282377,I282145);
nor I_16276 (I282425,I282377,I282179);
nand I_16277 (I282028,I282111,I282425);
or I_16278 (I282456,I282377,I282346);
DFFARX1 I_16279  ( .D(I282456), .CLK(I5694_clk), .RSTB(I282060_rst), .Q(I282025) );
not I_16280 (I282031,I282377);
DFFARX1 I_16281  ( .D(I269967), .CLK(I5694_clk), .RSTB(I282060_rst), .Q(I282501) );
not I_16282 (I282518,I282501);
nor I_16283 (I282535,I282518,I282111);
DFFARX1 I_16284  ( .D(I282535), .CLK(I5694_clk), .RSTB(I282060_rst), .Q(I282037) );
nor I_16285 (I282052,I282377,I282518);
nor I_16286 (I282040,I282518,I282281);
not I_16287 (I282594,I282518);
and I_16288 (I282611,I282145,I282594);
nor I_16289 (I282046,I282281,I282611);
nand I_16290 (I282034,I282518,I282408);
not I_16291 (I282689_rst,I5701);
not I_16292 (I282706,I249094);
nor I_16293 (I282723,I249100,I249079);
nand I_16294 (I282740,I282723,I249085);
nor I_16295 (I282757,I282706,I249100);
nand I_16296 (I282774,I282757,I249091);
not I_16297 (I282791,I249100);
not I_16298 (I282808,I282791);
not I_16299 (I282825,I249088);
nor I_16300 (I282842,I282825,I249106);
and I_16301 (I282859,I282842,I249097);
or I_16302 (I282876,I282859,I249076);
DFFARX1 I_16303  ( .D(I282876), .CLK(I5694_clk), .RSTB(I282689_rst), .Q(I282893) );
nand I_16304 (I282910,I282706,I249088);
or I_16305 (I282678,I282910,I282893);
not I_16306 (I282941,I282910);
nor I_16307 (I282958,I282893,I282941);
and I_16308 (I282975,I282791,I282958);
nand I_16309 (I282651,I282910,I282808);
DFFARX1 I_16310  ( .D(I249103), .CLK(I5694_clk), .RSTB(I282689_rst), .Q(I283006) );
or I_16311 (I282672,I283006,I282893);
nor I_16312 (I283037,I283006,I282774);
nor I_16313 (I283054,I283006,I282808);
nand I_16314 (I282657,I282740,I283054);
or I_16315 (I283085,I283006,I282975);
DFFARX1 I_16316  ( .D(I283085), .CLK(I5694_clk), .RSTB(I282689_rst), .Q(I282654) );
not I_16317 (I282660,I283006);
DFFARX1 I_16318  ( .D(I249082), .CLK(I5694_clk), .RSTB(I282689_rst), .Q(I283130) );
not I_16319 (I283147,I283130);
nor I_16320 (I283164,I283147,I282740);
DFFARX1 I_16321  ( .D(I283164), .CLK(I5694_clk), .RSTB(I282689_rst), .Q(I282666) );
nor I_16322 (I282681,I283006,I283147);
nor I_16323 (I282669,I283147,I282910);
not I_16324 (I283223,I283147);
and I_16325 (I283240,I282774,I283223);
nor I_16326 (I282675,I282910,I283240);
nand I_16327 (I282663,I283147,I283037);
not I_16328 (I283318_rst,I5701);
not I_16329 (I283335,I278291);
nor I_16330 (I283352,I278294,I278303);
nand I_16331 (I283369,I283352,I278288);
nor I_16332 (I283386,I283335,I278294);
nand I_16333 (I283403,I283386,I278297);
not I_16334 (I283420,I278294);
not I_16335 (I283437,I283420);
not I_16336 (I283454,I278312);
nor I_16337 (I283471,I283454,I278300);
and I_16338 (I283488,I283471,I278285);
or I_16339 (I283505,I283488,I278282);
DFFARX1 I_16340  ( .D(I283505), .CLK(I5694_clk), .RSTB(I283318_rst), .Q(I28352_rst2) );
nand I_16341 (I283539,I283335,I278312);
or I_16342 (I283307,I283539,I28352_rst2);
not I_16343 (I283570,I283539);
nor I_16344 (I283587,I28352_rst2,I283570);
and I_16345 (I283604,I283420,I283587);
nand I_16346 (I283280,I283539,I283437);
DFFARX1 I_16347  ( .D(I278306), .CLK(I5694_clk), .RSTB(I283318_rst), .Q(I283635) );
or I_16348 (I283301,I283635,I28352_rst2);
nor I_16349 (I283666,I283635,I283403);
nor I_16350 (I283683,I283635,I283437);
nand I_16351 (I283286,I283369,I283683);
or I_16352 (I283714,I283635,I283604);
DFFARX1 I_16353  ( .D(I283714), .CLK(I5694_clk), .RSTB(I283318_rst), .Q(I283283) );
not I_16354 (I283289,I283635);
DFFARX1 I_16355  ( .D(I278309), .CLK(I5694_clk), .RSTB(I283318_rst), .Q(I283759) );
not I_16356 (I283776,I283759);
nor I_16357 (I283793,I283776,I283369);
DFFARX1 I_16358  ( .D(I283793), .CLK(I5694_clk), .RSTB(I283318_rst), .Q(I283295) );
nor I_16359 (I283310,I283635,I283776);
nor I_16360 (I283298,I283776,I283539);
not I_16361 (I283852,I283776);
and I_16362 (I283869,I283403,I283852);
nor I_16363 (I283304,I283539,I283869);
nand I_16364 (I283292,I283776,I283666);
not I_16365 (I283947_rst,I5701);
not I_16366 (I283964,I258223);
nor I_16367 (I283981,I258232,I258235);
nand I_16368 (I283998,I283981,I258220);
nor I_16369 (I284015,I283964,I258232);
nand I_16370 (I284032,I284015,I258217);
not I_16371 (I284049,I258232);
not I_16372 (I284066,I284049);
not I_16373 (I284083,I258205);
nor I_16374 (I284100,I284083,I258211);
and I_16375 (I284117,I284100,I258208);
or I_16376 (I284134,I284117,I258229);
DFFARX1 I_16377  ( .D(I284134), .CLK(I5694_clk), .RSTB(I283947_rst), .Q(I284151) );
nand I_16378 (I284168,I283964,I258205);
or I_16379 (I283936,I284168,I284151);
not I_16380 (I284199,I284168);
nor I_16381 (I284216,I284151,I284199);
and I_16382 (I284233,I284049,I284216);
nand I_16383 (I283909,I284168,I284066);
DFFARX1 I_16384  ( .D(I258214), .CLK(I5694_clk), .RSTB(I283947_rst), .Q(I284264) );
or I_16385 (I283930,I284264,I284151);
nor I_16386 (I284295,I284264,I284032);
nor I_16387 (I284312,I284264,I284066);
nand I_16388 (I283915,I283998,I284312);
or I_16389 (I284343,I284264,I284233);
DFFARX1 I_16390  ( .D(I284343), .CLK(I5694_clk), .RSTB(I283947_rst), .Q(I283912) );
not I_16391 (I283918,I284264);
DFFARX1 I_16392  ( .D(I258226), .CLK(I5694_clk), .RSTB(I283947_rst), .Q(I284388) );
not I_16393 (I284405,I284388);
nor I_16394 (I284422,I284405,I283998);
DFFARX1 I_16395  ( .D(I284422), .CLK(I5694_clk), .RSTB(I283947_rst), .Q(I283924) );
nor I_16396 (I283939,I284264,I284405);
nor I_16397 (I283927,I284405,I284168);
not I_16398 (I284481,I284405);
and I_16399 (I284498,I284032,I284481);
nor I_16400 (I283933,I284168,I284498);
nand I_16401 (I283921,I284405,I284295);
not I_16402 (I284576_rst,I5701);
not I_16403 (I284593,I266429);
nor I_16404 (I284610,I266402,I266420);
nand I_16405 (I284627,I284610,I266405);
nor I_16406 (I284644,I284593,I266402);
nand I_16407 (I284661,I284644,I266423);
not I_16408 (I284678,I266402);
not I_16409 (I284695,I284678);
not I_16410 (I284712,I266399);
nor I_16411 (I284729,I284712,I266426);
and I_16412 (I284746,I284729,I266417);
or I_16413 (I284763,I284746,I266408);
DFFARX1 I_16414  ( .D(I284763), .CLK(I5694_clk), .RSTB(I284576_rst), .Q(I284780) );
nand I_16415 (I284797,I284593,I266399);
or I_16416 (I284565,I284797,I284780);
not I_16417 (I284828,I284797);
nor I_16418 (I284845,I284780,I284828);
and I_16419 (I284862,I284678,I284845);
nand I_16420 (I284538,I284797,I284695);
DFFARX1 I_16421  ( .D(I266411), .CLK(I5694_clk), .RSTB(I284576_rst), .Q(I284893) );
or I_16422 (I284559,I284893,I284780);
nor I_16423 (I284924,I284893,I284661);
nor I_16424 (I284941,I284893,I284695);
nand I_16425 (I284544,I284627,I284941);
or I_16426 (I284972,I284893,I284862);
DFFARX1 I_16427  ( .D(I284972), .CLK(I5694_clk), .RSTB(I284576_rst), .Q(I284541) );
not I_16428 (I284547,I284893);
DFFARX1 I_16429  ( .D(I266414), .CLK(I5694_clk), .RSTB(I284576_rst), .Q(I285017) );
not I_16430 (I285034,I285017);
nor I_16431 (I285051,I285034,I284627);
DFFARX1 I_16432  ( .D(I285051), .CLK(I5694_clk), .RSTB(I284576_rst), .Q(I284553) );
nor I_16433 (I284568,I284893,I285034);
nor I_16434 (I284556,I285034,I284797);
not I_16435 (I285110,I285034);
and I_16436 (I285127,I284661,I285110);
nor I_16437 (I284562,I284797,I285127);
nand I_16438 (I284550,I285034,I284924);
not I_16439 (I285205_rst,I5701);
not I_16440 (I285222,I252409);
nor I_16441 (I285239,I252418,I252421);
nand I_16442 (I285256,I285239,I252406);
nor I_16443 (I285273,I285222,I252418);
nand I_16444 (I285290,I285273,I252403);
not I_16445 (I285307,I252418);
not I_16446 (I285324,I285307);
not I_16447 (I285341,I252391);
nor I_16448 (I285358,I285341,I252397);
and I_16449 (I285375,I285358,I252394);
or I_16450 (I285392,I285375,I252415);
DFFARX1 I_16451  ( .D(I285392), .CLK(I5694_clk), .RSTB(I285205_rst), .Q(I285409) );
nand I_16452 (I285426,I285222,I252391);
or I_16453 (I285194,I285426,I285409);
not I_16454 (I285457,I285426);
nor I_16455 (I285474,I285409,I285457);
and I_16456 (I285491,I285307,I285474);
nand I_16457 (I285167,I285426,I285324);
DFFARX1 I_16458  ( .D(I252400), .CLK(I5694_clk), .RSTB(I285205_rst), .Q(I285522) );
or I_16459 (I285188,I285522,I285409);
nor I_16460 (I285553,I285522,I285290);
nor I_16461 (I285570,I285522,I285324);
nand I_16462 (I285173,I285256,I285570);
or I_16463 (I285601,I285522,I285491);
DFFARX1 I_16464  ( .D(I285601), .CLK(I5694_clk), .RSTB(I285205_rst), .Q(I285170) );
not I_16465 (I285176,I285522);
DFFARX1 I_16466  ( .D(I252412), .CLK(I5694_clk), .RSTB(I285205_rst), .Q(I285646) );
not I_16467 (I285663,I285646);
nor I_16468 (I285680,I285663,I285256);
DFFARX1 I_16469  ( .D(I285680), .CLK(I5694_clk), .RSTB(I285205_rst), .Q(I285182) );
nor I_16470 (I285197,I285522,I285663);
nor I_16471 (I285185,I285663,I285426);
not I_16472 (I285739,I285663);
and I_16473 (I285756,I285290,I285739);
nor I_16474 (I285191,I285426,I285756);
nand I_16475 (I285179,I285663,I285553);
not I_16476 (I285834_rst,I5701);
nand I_16477 (I285851,I240211,I240208);
and I_16478 (I285868,I285851,I240220);
DFFARX1 I_16479  ( .D(I285868), .CLK(I5694_clk), .RSTB(I285834_rst), .Q(I285885) );
not I_16480 (I285823,I285885);
DFFARX1 I_16481  ( .D(I285885), .CLK(I5694_clk), .RSTB(I285834_rst), .Q(I285916) );
not I_16482 (I285811,I285916);
nor I_16483 (I285947,I240223,I240208);
not I_16484 (I285964,I285947);
nor I_16485 (I285981,I285885,I285964);
DFFARX1 I_16486  ( .D(I240229), .CLK(I5694_clk), .RSTB(I285834_rst), .Q(I285998) );
not I_16487 (I286015,I285998);
nand I_16488 (I285814,I285998,I285964);
DFFARX1 I_16489  ( .D(I285998), .CLK(I5694_clk), .RSTB(I285834_rst), .Q(I286046) );
and I_16490 (I285799,I285885,I286046);
nand I_16491 (I286077,I240202,I240205);
and I_16492 (I286094,I286077,I240214);
DFFARX1 I_16493  ( .D(I286094), .CLK(I5694_clk), .RSTB(I285834_rst), .Q(I286111) );
nor I_16494 (I286128,I286111,I286015);
and I_16495 (I286145,I285947,I286128);
nor I_16496 (I286162,I286111,I285885);
DFFARX1 I_16497  ( .D(I286111), .CLK(I5694_clk), .RSTB(I285834_rst), .Q(I285805) );
DFFARX1 I_16498  ( .D(I240232), .CLK(I5694_clk), .RSTB(I285834_rst), .Q(I286193) );
and I_16499 (I286210,I286193,I240226);
or I_16500 (I286227,I286210,I286145);
DFFARX1 I_16501  ( .D(I286227), .CLK(I5694_clk), .RSTB(I285834_rst), .Q(I285817) );
nand I_16502 (I285826,I286210,I286162);
DFFARX1 I_16503  ( .D(I286210), .CLK(I5694_clk), .RSTB(I285834_rst), .Q(I285796) );
DFFARX1 I_16504  ( .D(I240217), .CLK(I5694_clk), .RSTB(I285834_rst), .Q(I286286) );
nand I_16505 (I285820,I286286,I285981);
DFFARX1 I_16506  ( .D(I286286), .CLK(I5694_clk), .RSTB(I285834_rst), .Q(I285808) );
nand I_16507 (I286331,I286286,I285947);
and I_16508 (I286348,I285998,I286331);
DFFARX1 I_16509  ( .D(I286348), .CLK(I5694_clk), .RSTB(I285834_rst), .Q(I285802) );
not I_16510 (I286412_rst,I5701);
nand I_16511 (I286429,I279509,I279527);
and I_16512 (I286446,I286429,I279524);
DFFARX1 I_16513  ( .D(I286446), .CLK(I5694_clk), .RSTB(I286412_rst), .Q(I286463) );
not I_16514 (I286401,I286463);
DFFARX1 I_16515  ( .D(I286463), .CLK(I5694_clk), .RSTB(I286412_rst), .Q(I286494) );
not I_16516 (I286389,I286494);
nor I_16517 (I286525,I279530,I279527);
not I_16518 (I286542,I286525);
nor I_16519 (I286559,I286463,I286542);
DFFARX1 I_16520  ( .D(I279533), .CLK(I5694_clk), .RSTB(I286412_rst), .Q(I286576) );
not I_16521 (I286593,I286576);
nand I_16522 (I286392,I286576,I286542);
DFFARX1 I_16523  ( .D(I286576), .CLK(I5694_clk), .RSTB(I286412_rst), .Q(I286624) );
and I_16524 (I286377,I286463,I286624);
nand I_16525 (I286655,I279518,I279512);
and I_16526 (I286672,I286655,I279515);
DFFARX1 I_16527  ( .D(I286672), .CLK(I5694_clk), .RSTB(I286412_rst), .Q(I286689) );
nor I_16528 (I286706,I286689,I286593);
and I_16529 (I286723,I286525,I286706);
nor I_16530 (I286740,I286689,I286463);
DFFARX1 I_16531  ( .D(I286689), .CLK(I5694_clk), .RSTB(I286412_rst), .Q(I286383) );
DFFARX1 I_16532  ( .D(I279521), .CLK(I5694_clk), .RSTB(I286412_rst), .Q(I286771) );
and I_16533 (I286788,I286771,I279506);
or I_16534 (I286805,I286788,I286723);
DFFARX1 I_16535  ( .D(I286805), .CLK(I5694_clk), .RSTB(I286412_rst), .Q(I286395) );
nand I_16536 (I286404,I286788,I286740);
DFFARX1 I_16537  ( .D(I286788), .CLK(I5694_clk), .RSTB(I286412_rst), .Q(I286374) );
DFFARX1 I_16538  ( .D(I279536), .CLK(I5694_clk), .RSTB(I286412_rst), .Q(I286864) );
nand I_16539 (I286398,I286864,I286559);
DFFARX1 I_16540  ( .D(I286864), .CLK(I5694_clk), .RSTB(I286412_rst), .Q(I286386) );
nand I_16541 (I286909,I286864,I286525);
and I_16542 (I286926,I286576,I286909);
DFFARX1 I_16543  ( .D(I286926), .CLK(I5694_clk), .RSTB(I286412_rst), .Q(I286380) );
not I_16544 (I286990_rst,I5701);
nand I_16545 (I287007,I268188,I268170);
and I_16546 (I287024,I287007,I268185);
DFFARX1 I_16547  ( .D(I287024), .CLK(I5694_clk), .RSTB(I286990_rst), .Q(I287041) );
not I_16548 (I286979,I287041);
DFFARX1 I_16549  ( .D(I287041), .CLK(I5694_clk), .RSTB(I286990_rst), .Q(I287072) );
not I_16550 (I286967,I287072);
nor I_16551 (I287103,I268176,I268170);
not I_16552 (I287120,I287103);
nor I_16553 (I287137,I287041,I287120);
DFFARX1 I_16554  ( .D(I268191), .CLK(I5694_clk), .RSTB(I286990_rst), .Q(I287154) );
not I_16555 (I287171,I287154);
nand I_16556 (I286970,I287154,I287120);
DFFARX1 I_16557  ( .D(I287154), .CLK(I5694_clk), .RSTB(I286990_rst), .Q(I287202) );
and I_16558 (I286955,I287041,I287202);
nand I_16559 (I287233,I268167,I268173);
and I_16560 (I287250,I287233,I268179);
DFFARX1 I_16561  ( .D(I287250), .CLK(I5694_clk), .RSTB(I286990_rst), .Q(I287267) );
nor I_16562 (I287284,I287267,I287171);
and I_16563 (I287301,I287103,I287284);
nor I_16564 (I287318,I287267,I287041);
DFFARX1 I_16565  ( .D(I287267), .CLK(I5694_clk), .RSTB(I286990_rst), .Q(I286961) );
DFFARX1 I_16566  ( .D(I268194), .CLK(I5694_clk), .RSTB(I286990_rst), .Q(I287349) );
and I_16567 (I287366,I287349,I268182);
or I_16568 (I287383,I287366,I287301);
DFFARX1 I_16569  ( .D(I287383), .CLK(I5694_clk), .RSTB(I286990_rst), .Q(I286973) );
nand I_16570 (I286982,I287366,I287318);
DFFARX1 I_16571  ( .D(I287366), .CLK(I5694_clk), .RSTB(I286990_rst), .Q(I286952) );
DFFARX1 I_16572  ( .D(I268197), .CLK(I5694_clk), .RSTB(I286990_rst), .Q(I287442) );
nand I_16573 (I286976,I287442,I287137);
DFFARX1 I_16574  ( .D(I287442), .CLK(I5694_clk), .RSTB(I286990_rst), .Q(I286964) );
nand I_16575 (I287487,I287442,I287103);
and I_16576 (I287504,I287154,I287487);
DFFARX1 I_16577  ( .D(I287504), .CLK(I5694_clk), .RSTB(I286990_rst), .Q(I286958) );
not I_16578 (I287568_rst,I5701);
nand I_16579 (I287585,I234970,I234955);
and I_16580 (I287602,I287585,I234949);
DFFARX1 I_16581  ( .D(I287602), .CLK(I5694_clk), .RSTB(I287568_rst), .Q(I287619) );
not I_16582 (I287557,I287619);
DFFARX1 I_16583  ( .D(I287619), .CLK(I5694_clk), .RSTB(I287568_rst), .Q(I287650) );
not I_16584 (I287545,I287650);
nor I_16585 (I287681,I234976,I234955);
not I_16586 (I287698,I287681);
nor I_16587 (I287715,I287619,I287698);
DFFARX1 I_16588  ( .D(I234979), .CLK(I5694_clk), .RSTB(I287568_rst), .Q(I287732) );
not I_16589 (I287749,I287732);
nand I_16590 (I287548,I287732,I287698);
DFFARX1 I_16591  ( .D(I287732), .CLK(I5694_clk), .RSTB(I287568_rst), .Q(I287780) );
and I_16592 (I287533,I287619,I287780);
nand I_16593 (I287811,I234961,I234964);
and I_16594 (I287828,I287811,I234967);
DFFARX1 I_16595  ( .D(I287828), .CLK(I5694_clk), .RSTB(I287568_rst), .Q(I287845) );
nor I_16596 (I287862,I287845,I287749);
and I_16597 (I287879,I287681,I287862);
nor I_16598 (I287896,I287845,I287619);
DFFARX1 I_16599  ( .D(I287845), .CLK(I5694_clk), .RSTB(I287568_rst), .Q(I287539) );
DFFARX1 I_16600  ( .D(I234973), .CLK(I5694_clk), .RSTB(I287568_rst), .Q(I287927) );
and I_16601 (I287944,I287927,I234958);
or I_16602 (I287961,I287944,I287879);
DFFARX1 I_16603  ( .D(I287961), .CLK(I5694_clk), .RSTB(I287568_rst), .Q(I287551) );
nand I_16604 (I287560,I287944,I287896);
DFFARX1 I_16605  ( .D(I287944), .CLK(I5694_clk), .RSTB(I287568_rst), .Q(I287530) );
DFFARX1 I_16606  ( .D(I234952), .CLK(I5694_clk), .RSTB(I287568_rst), .Q(I288020) );
nand I_16607 (I287554,I288020,I287715);
DFFARX1 I_16608  ( .D(I288020), .CLK(I5694_clk), .RSTB(I287568_rst), .Q(I287542) );
nand I_16609 (I288065,I288020,I287681);
and I_16610 (I288082,I287732,I288065);
DFFARX1 I_16611  ( .D(I288082), .CLK(I5694_clk), .RSTB(I287568_rst), .Q(I287536) );
not I_16612 (I288146_rst,I5701);
nand I_16613 (I288163,I243781,I243778);
and I_16614 (I288180,I288163,I243802);
DFFARX1 I_16615  ( .D(I288180), .CLK(I5694_clk), .RSTB(I288146_rst), .Q(I288197) );
not I_16616 (I288135,I288197);
DFFARX1 I_16617  ( .D(I288197), .CLK(I5694_clk), .RSTB(I288146_rst), .Q(I288228) );
not I_16618 (I288123,I288228);
nor I_16619 (I288259,I243784,I243778);
not I_16620 (I288276,I288259);
nor I_16621 (I288293,I288197,I288276);
DFFARX1 I_16622  ( .D(I243799), .CLK(I5694_clk), .RSTB(I288146_rst), .Q(I288310) );
not I_16623 (I288327,I288310);
nand I_16624 (I288126,I288310,I288276);
DFFARX1 I_16625  ( .D(I288310), .CLK(I5694_clk), .RSTB(I288146_rst), .Q(I288358) );
and I_16626 (I288111,I288197,I288358);
nand I_16627 (I288389,I243787,I243772);
and I_16628 (I288406,I288389,I243790);
DFFARX1 I_16629  ( .D(I288406), .CLK(I5694_clk), .RSTB(I288146_rst), .Q(I288423) );
nor I_16630 (I288440,I288423,I288327);
and I_16631 (I288457,I288259,I288440);
nor I_16632 (I288474,I288423,I288197);
DFFARX1 I_16633  ( .D(I288423), .CLK(I5694_clk), .RSTB(I288146_rst), .Q(I288117) );
DFFARX1 I_16634  ( .D(I243793), .CLK(I5694_clk), .RSTB(I288146_rst), .Q(I288505) );
and I_16635 (I288522,I288505,I243796);
or I_16636 (I288539,I288522,I288457);
DFFARX1 I_16637  ( .D(I288539), .CLK(I5694_clk), .RSTB(I288146_rst), .Q(I288129) );
nand I_16638 (I288138,I288522,I288474);
DFFARX1 I_16639  ( .D(I288522), .CLK(I5694_clk), .RSTB(I288146_rst), .Q(I288108) );
DFFARX1 I_16640  ( .D(I243775), .CLK(I5694_clk), .RSTB(I288146_rst), .Q(I288598) );
nand I_16641 (I288132,I288598,I288293);
DFFARX1 I_16642  ( .D(I288598), .CLK(I5694_clk), .RSTB(I288146_rst), .Q(I288120) );
nand I_16643 (I288643,I288598,I288259);
and I_16644 (I288660,I288310,I288643);
DFFARX1 I_16645  ( .D(I288660), .CLK(I5694_clk), .RSTB(I288146_rst), .Q(I288114) );
not I_16646 (I288724_rst,I5701);
nand I_16647 (I288741,I259475,I259472);
and I_16648 (I288758,I288741,I259466);
DFFARX1 I_16649  ( .D(I288758), .CLK(I5694_clk), .RSTB(I288724_rst), .Q(I288775) );
not I_16650 (I288792,I288775);
nor I_16651 (I288809,I259478,I259472);
or I_16652 (I288707,I288809,I288775);
not I_16653 (I288695,I288809);
DFFARX1 I_16654  ( .D(I259490), .CLK(I5694_clk), .RSTB(I288724_rst), .Q(I288854) );
nor I_16655 (I288871,I288854,I288809);
nand I_16656 (I288888,I259481,I259463);
and I_16657 (I288905,I288888,I259493);
DFFARX1 I_16658  ( .D(I288905), .CLK(I5694_clk), .RSTB(I288724_rst), .Q(I288922) );
nor I_16659 (I288704,I288922,I288775);
not I_16660 (I288953,I288922);
nor I_16661 (I288970,I288854,I288953);
DFFARX1 I_16662  ( .D(I259469), .CLK(I5694_clk), .RSTB(I288724_rst), .Q(I288987) );
and I_16663 (I289004,I288987,I259487);
or I_16664 (I288713,I289004,I288809);
nand I_16665 (I288692,I289004,I288970);
DFFARX1 I_16666  ( .D(I259484), .CLK(I5694_clk), .RSTB(I288724_rst), .Q(I289049) );
and I_16667 (I289066,I289049,I288792);
nor I_16668 (I288710,I289004,I289066);
nor I_16669 (I289097,I289049,I288854);
DFFARX1 I_16670  ( .D(I289097), .CLK(I5694_clk), .RSTB(I288724_rst), .Q(I288701) );
nor I_16671 (I288716,I289049,I288775);
not I_16672 (I289142,I289049);
nor I_16673 (I289159,I288922,I289142);
and I_16674 (I289176,I288809,I289159);
or I_16675 (I289193,I289004,I289176);
DFFARX1 I_16676  ( .D(I289193), .CLK(I5694_clk), .RSTB(I288724_rst), .Q(I288689) );
nand I_16677 (I288698,I289049,I288871);
nand I_16678 (I288686,I289049,I288953);
not I_16679 (I289285_rst,I5701);
nand I_16680 (I289302,I245785,I245776);
and I_16681 (I289319,I289302,I245791);
DFFARX1 I_16682  ( .D(I289319), .CLK(I5694_clk), .RSTB(I289285_rst), .Q(I289336) );
not I_16683 (I289353,I289336);
nor I_16684 (I289370,I245761,I245776);
or I_16685 (I289268,I289370,I289336);
not I_16686 (I289256,I289370);
DFFARX1 I_16687  ( .D(I245764), .CLK(I5694_clk), .RSTB(I289285_rst), .Q(I289415) );
nor I_16688 (I289432,I289415,I289370);
nand I_16689 (I289449,I245782,I245779);
and I_16690 (I289466,I289449,I245767);
DFFARX1 I_16691  ( .D(I289466), .CLK(I5694_clk), .RSTB(I289285_rst), .Q(I289483) );
nor I_16692 (I289265,I289483,I289336);
not I_16693 (I289514,I289483);
nor I_16694 (I289531,I289415,I289514);
DFFARX1 I_16695  ( .D(I245788), .CLK(I5694_clk), .RSTB(I289285_rst), .Q(I289548) );
and I_16696 (I289565,I289548,I245773);
or I_16697 (I289274,I289565,I289370);
nand I_16698 (I289253,I289565,I289531);
DFFARX1 I_16699  ( .D(I245770), .CLK(I5694_clk), .RSTB(I289285_rst), .Q(I289610) );
and I_16700 (I289627,I289610,I289353);
nor I_16701 (I289271,I289565,I289627);
nor I_16702 (I289658,I289610,I289415);
DFFARX1 I_16703  ( .D(I289658), .CLK(I5694_clk), .RSTB(I289285_rst), .Q(I289262) );
nor I_16704 (I289277,I289610,I289336);
not I_16705 (I289703,I289610);
nor I_16706 (I289720,I289483,I289703);
and I_16707 (I289737,I289370,I289720);
or I_16708 (I289754,I289565,I289737);
DFFARX1 I_16709  ( .D(I289754), .CLK(I5694_clk), .RSTB(I289285_rst), .Q(I289250) );
nand I_16710 (I289259,I289610,I289432);
nand I_16711 (I289247,I289610,I289514);
not I_16712 (I289846_rst,I5701);
nand I_16713 (I289863,I261787,I261784);
and I_16714 (I289880,I289863,I261778);
DFFARX1 I_16715  ( .D(I289880), .CLK(I5694_clk), .RSTB(I289846_rst), .Q(I289897) );
not I_16716 (I289914,I289897);
nor I_16717 (I289931,I261790,I261784);
or I_16718 (I289829,I289931,I289897);
not I_16719 (I289817,I289931);
DFFARX1 I_16720  ( .D(I261802), .CLK(I5694_clk), .RSTB(I289846_rst), .Q(I289976) );
nor I_16721 (I289993,I289976,I289931);
nand I_16722 (I290010,I261793,I261775);
and I_16723 (I290027,I290010,I261805);
DFFARX1 I_16724  ( .D(I290027), .CLK(I5694_clk), .RSTB(I289846_rst), .Q(I290044) );
nor I_16725 (I289826,I290044,I289897);
not I_16726 (I290075,I290044);
nor I_16727 (I290092,I289976,I290075);
DFFARX1 I_16728  ( .D(I261781), .CLK(I5694_clk), .RSTB(I289846_rst), .Q(I290109) );
and I_16729 (I290126,I290109,I261799);
or I_16730 (I289835,I290126,I289931);
nand I_16731 (I289814,I290126,I290092);
DFFARX1 I_16732  ( .D(I261796), .CLK(I5694_clk), .RSTB(I289846_rst), .Q(I290171) );
and I_16733 (I290188,I290171,I289914);
nor I_16734 (I289832,I290126,I290188);
nor I_16735 (I290219,I290171,I289976);
DFFARX1 I_16736  ( .D(I290219), .CLK(I5694_clk), .RSTB(I289846_rst), .Q(I289823) );
nor I_16737 (I289838,I290171,I289897);
not I_16738 (I290264,I290171);
nor I_16739 (I290281,I290044,I290264);
and I_16740 (I290298,I289931,I290281);
or I_16741 (I290315,I290126,I290298);
DFFARX1 I_16742  ( .D(I290315), .CLK(I5694_clk), .RSTB(I289846_rst), .Q(I289811) );
nand I_16743 (I289820,I290171,I289993);
nand I_16744 (I289808,I290171,I290075);
not I_16745 (I290407_rst,I5701);
nand I_16746 (I290424,I257589,I257580);
and I_16747 (I290441,I290424,I257583);
DFFARX1 I_16748  ( .D(I290441), .CLK(I5694_clk), .RSTB(I290407_rst), .Q(I290458) );
not I_16749 (I290475,I290458);
nor I_16750 (I290492,I257559,I257580);
or I_16751 (I290390,I290492,I290458);
not I_16752 (I290378,I290492);
DFFARX1 I_16753  ( .D(I257574), .CLK(I5694_clk), .RSTB(I290407_rst), .Q(I290537) );
nor I_16754 (I290554,I290537,I290492);
nand I_16755 (I290571,I257562,I257577);
and I_16756 (I290588,I290571,I257571);
DFFARX1 I_16757  ( .D(I290588), .CLK(I5694_clk), .RSTB(I290407_rst), .Q(I290605) );
nor I_16758 (I290387,I290605,I290458);
not I_16759 (I290636,I290605);
nor I_16760 (I290653,I290537,I290636);
DFFARX1 I_16761  ( .D(I257586), .CLK(I5694_clk), .RSTB(I290407_rst), .Q(I290670) );
and I_16762 (I290687,I290670,I257565);
or I_16763 (I290396,I290687,I290492);
nand I_16764 (I290375,I290687,I290653);
DFFARX1 I_16765  ( .D(I257568), .CLK(I5694_clk), .RSTB(I290407_rst), .Q(I290732) );
and I_16766 (I290749,I290732,I290475);
nor I_16767 (I290393,I290687,I290749);
nor I_16768 (I290780,I290732,I290537);
DFFARX1 I_16769  ( .D(I290780), .CLK(I5694_clk), .RSTB(I290407_rst), .Q(I290384) );
nor I_16770 (I290399,I290732,I290458);
not I_16771 (I290825,I290732);
nor I_16772 (I290842,I290605,I290825);
and I_16773 (I290859,I290492,I290842);
or I_16774 (I290876,I290687,I290859);
DFFARX1 I_16775  ( .D(I290876), .CLK(I5694_clk), .RSTB(I290407_rst), .Q(I290372) );
nand I_16776 (I290381,I290732,I290554);
nand I_16777 (I290369,I290732,I290636);
not I_16778 (I290968_rst,I5701);
nand I_16779 (I290985,I235616,I235619);
and I_16780 (I291002,I290985,I235601);
DFFARX1 I_16781  ( .D(I291002), .CLK(I5694_clk), .RSTB(I290968_rst), .Q(I291019) );
not I_16782 (I291036,I291019);
nor I_16783 (I291053,I235598,I235619);
or I_16784 (I290951,I291053,I291019);
not I_16785 (I290939,I291053);
DFFARX1 I_16786  ( .D(I235622), .CLK(I5694_clk), .RSTB(I290968_rst), .Q(I291098) );
nor I_16787 (I291115,I291098,I291053);
nand I_16788 (I291132,I235607,I235613);
and I_16789 (I291149,I291132,I235625);
DFFARX1 I_16790  ( .D(I291149), .CLK(I5694_clk), .RSTB(I290968_rst), .Q(I291166) );
nor I_16791 (I290948,I291166,I291019);
not I_16792 (I291197,I291166);
nor I_16793 (I291214,I291098,I291197);
DFFARX1 I_16794  ( .D(I235604), .CLK(I5694_clk), .RSTB(I290968_rst), .Q(I291231) );
and I_16795 (I291248,I291231,I235595);
or I_16796 (I290957,I291248,I291053);
nand I_16797 (I290936,I291248,I291214);
DFFARX1 I_16798  ( .D(I235610), .CLK(I5694_clk), .RSTB(I290968_rst), .Q(I291293) );
and I_16799 (I291310,I291293,I291036);
nor I_16800 (I290954,I291248,I291310);
nor I_16801 (I291341,I291293,I291098);
DFFARX1 I_16802  ( .D(I291341), .CLK(I5694_clk), .RSTB(I290968_rst), .Q(I290945) );
nor I_16803 (I290960,I291293,I291019);
not I_16804 (I291386,I291293);
nor I_16805 (I291403,I291166,I291386);
and I_16806 (I291420,I291053,I291403);
or I_16807 (I291437,I291248,I291420);
DFFARX1 I_16808  ( .D(I291437), .CLK(I5694_clk), .RSTB(I290968_rst), .Q(I290933) );
nand I_16809 (I290942,I291293,I291115);
nand I_16810 (I290930,I291293,I291197);
not I_16811 (I291529_rst,I5701);
nand I_16812 (I291546,I233032,I233035);
and I_16813 (I291563,I291546,I233017);
DFFARX1 I_16814  ( .D(I291563), .CLK(I5694_clk), .RSTB(I291529_rst), .Q(I291580) );
not I_16815 (I291597,I291580);
nor I_16816 (I291614,I233014,I233035);
or I_16817 (I291512,I291614,I291580);
not I_16818 (I291500,I291614);
DFFARX1 I_16819  ( .D(I233038), .CLK(I5694_clk), .RSTB(I291529_rst), .Q(I291659) );
nor I_16820 (I291676,I291659,I291614);
nand I_16821 (I291693,I233023,I233029);
and I_16822 (I291710,I291693,I233041);
DFFARX1 I_16823  ( .D(I291710), .CLK(I5694_clk), .RSTB(I291529_rst), .Q(I291727) );
nor I_16824 (I291509,I291727,I291580);
not I_16825 (I291758,I291727);
nor I_16826 (I291775,I291659,I291758);
DFFARX1 I_16827  ( .D(I233020), .CLK(I5694_clk), .RSTB(I291529_rst), .Q(I291792) );
and I_16828 (I291809,I291792,I233011);
or I_16829 (I291518,I291809,I291614);
nand I_16830 (I291497,I291809,I291775);
DFFARX1 I_16831  ( .D(I233026), .CLK(I5694_clk), .RSTB(I291529_rst), .Q(I291854) );
and I_16832 (I291871,I291854,I291597);
nor I_16833 (I291515,I291809,I291871);
nor I_16834 (I291902,I291854,I291659);
DFFARX1 I_16835  ( .D(I291902), .CLK(I5694_clk), .RSTB(I291529_rst), .Q(I291506) );
nor I_16836 (I291521,I291854,I291580);
not I_16837 (I291947,I291854);
nor I_16838 (I291964,I291727,I291947);
and I_16839 (I291981,I291614,I291964);
or I_16840 (I291998,I291809,I291981);
DFFARX1 I_16841  ( .D(I291998), .CLK(I5694_clk), .RSTB(I291529_rst), .Q(I291494) );
nand I_16842 (I291503,I291854,I291676);
nand I_16843 (I291491,I291854,I291758);
not I_16844 (I292090_rst,I5701);
nand I_16845 (I292107,I262365,I262362);
and I_16846 (I292124,I292107,I262356);
DFFARX1 I_16847  ( .D(I292124), .CLK(I5694_clk), .RSTB(I292090_rst), .Q(I292141) );
not I_16848 (I292158,I292141);
nor I_16849 (I292175,I262368,I262362);
or I_16850 (I292073,I292175,I292141);
not I_16851 (I292061,I292175);
DFFARX1 I_16852  ( .D(I262380), .CLK(I5694_clk), .RSTB(I292090_rst), .Q(I292220) );
nor I_16853 (I292237,I292220,I292175);
nand I_16854 (I292254,I262371,I262353);
and I_16855 (I292271,I292254,I262383);
DFFARX1 I_16856  ( .D(I292271), .CLK(I5694_clk), .RSTB(I292090_rst), .Q(I292288) );
nor I_16857 (I292070,I292288,I292141);
not I_16858 (I292319,I292288);
nor I_16859 (I292336,I292220,I292319);
DFFARX1 I_16860  ( .D(I262359), .CLK(I5694_clk), .RSTB(I292090_rst), .Q(I292353) );
and I_16861 (I292370,I292353,I262377);
or I_16862 (I292079,I292370,I292175);
nand I_16863 (I292058,I292370,I292336);
DFFARX1 I_16864  ( .D(I262374), .CLK(I5694_clk), .RSTB(I292090_rst), .Q(I292415) );
and I_16865 (I292432,I292415,I292158);
nor I_16866 (I292076,I292370,I292432);
nor I_16867 (I292463,I292415,I292220);
DFFARX1 I_16868  ( .D(I292463), .CLK(I5694_clk), .RSTB(I292090_rst), .Q(I292067) );
nor I_16869 (I292082,I292415,I292141);
not I_16870 (I292508,I292415);
nor I_16871 (I292525,I292288,I292508);
and I_16872 (I292542,I292175,I292525);
or I_16873 (I292559,I292370,I292542);
DFFARX1 I_16874  ( .D(I292559), .CLK(I5694_clk), .RSTB(I292090_rst), .Q(I292055) );
nand I_16875 (I292064,I292415,I292237);
nand I_16876 (I292052,I292415,I292319);
not I_16877 (I292651_rst,I5701);
nand I_16878 (I292668,I262943,I262940);
and I_16879 (I292685,I292668,I262934);
DFFARX1 I_16880  ( .D(I292685), .CLK(I5694_clk), .RSTB(I292651_rst), .Q(I292702) );
not I_16881 (I292719,I292702);
nor I_16882 (I292736,I262946,I262940);
or I_16883 (I292634,I292736,I292702);
not I_16884 (I292622,I292736);
DFFARX1 I_16885  ( .D(I262958), .CLK(I5694_clk), .RSTB(I292651_rst), .Q(I292781) );
nor I_16886 (I292798,I292781,I292736);
nand I_16887 (I292815,I262949,I262931);
and I_16888 (I292832,I292815,I262961);
DFFARX1 I_16889  ( .D(I292832), .CLK(I5694_clk), .RSTB(I292651_rst), .Q(I292849) );
nor I_16890 (I292631,I292849,I292702);
not I_16891 (I292880,I292849);
nor I_16892 (I292897,I292781,I292880);
DFFARX1 I_16893  ( .D(I262937), .CLK(I5694_clk), .RSTB(I292651_rst), .Q(I292914) );
and I_16894 (I292931,I292914,I262955);
or I_16895 (I292640,I292931,I292736);
nand I_16896 (I292619,I292931,I292897);
DFFARX1 I_16897  ( .D(I262952), .CLK(I5694_clk), .RSTB(I292651_rst), .Q(I292976) );
and I_16898 (I292993,I292976,I292719);
nor I_16899 (I292637,I292931,I292993);
nor I_16900 (I293024,I292976,I292781);
DFFARX1 I_16901  ( .D(I293024), .CLK(I5694_clk), .RSTB(I292651_rst), .Q(I292628) );
nor I_16902 (I292643,I292976,I292702);
not I_16903 (I293069,I292976);
nor I_16904 (I293086,I292849,I293069);
and I_16905 (I293103,I292736,I293086);
or I_16906 (I293120,I292931,I293103);
DFFARX1 I_16907  ( .D(I293120), .CLK(I5694_clk), .RSTB(I292651_rst), .Q(I292616) );
nand I_16908 (I292625,I292976,I292798);
nand I_16909 (I292613,I292976,I292880);
not I_16910 (I293212_rst,I5701);
nand I_16911 (I293229,I266980,I266983);
and I_16912 (I293246,I293229,I266995);
DFFARX1 I_16913  ( .D(I293246), .CLK(I5694_clk), .RSTB(I293212_rst), .Q(I293263) );
not I_16914 (I293280,I293263);
nor I_16915 (I293297,I266989,I266983);
or I_16916 (I293195,I293297,I293263);
not I_16917 (I293183,I293297);
DFFARX1 I_16918  ( .D(I266992), .CLK(I5694_clk), .RSTB(I293212_rst), .Q(I293342) );
nor I_16919 (I293359,I293342,I293297);
nand I_16920 (I293376,I266986,I267004);
and I_16921 (I293393,I293376,I267007);
DFFARX1 I_16922  ( .D(I293393), .CLK(I5694_clk), .RSTB(I293212_rst), .Q(I293410) );
nor I_16923 (I293192,I293410,I293263);
not I_16924 (I293441,I293410);
nor I_16925 (I293458,I293342,I293441);
DFFARX1 I_16926  ( .D(I266977), .CLK(I5694_clk), .RSTB(I293212_rst), .Q(I293475) );
and I_16927 (I293492,I293475,I266998);
or I_16928 (I293201,I293492,I293297);
nand I_16929 (I293180,I293492,I293458);
DFFARX1 I_16930  ( .D(I267001), .CLK(I5694_clk), .RSTB(I293212_rst), .Q(I293537) );
and I_16931 (I293554,I293537,I293280);
nor I_16932 (I293198,I293492,I293554);
nor I_16933 (I293585,I293537,I293342);
DFFARX1 I_16934  ( .D(I293585), .CLK(I5694_clk), .RSTB(I293212_rst), .Q(I293189) );
nor I_16935 (I293204,I293537,I293263);
not I_16936 (I293630,I293537);
nor I_16937 (I293647,I293410,I293630);
and I_16938 (I293664,I293297,I293647);
or I_16939 (I293681,I293492,I293664);
DFFARX1 I_16940  ( .D(I293681), .CLK(I5694_clk), .RSTB(I293212_rst), .Q(I293177) );
nand I_16941 (I293186,I293537,I293359);
nand I_16942 (I293174,I293537,I293441);
not I_16943 (I293773_rst,I5701);
not I_16944 (I293790,I244453);
nor I_16945 (I293807,I244450,I244438);
nand I_16946 (I293824,I293807,I244441);
DFFARX1 I_16947  ( .D(I293824), .CLK(I5694_clk), .RSTB(I293773_rst), .Q(I293747) );
nor I_16948 (I293855,I293790,I244450);
nand I_16949 (I293872,I293855,I244447);
not I_16950 (I293762,I293872);
DFFARX1 I_16951  ( .D(I293872), .CLK(I5694_clk), .RSTB(I293773_rst), .Q(I293744) );
not I_16952 (I293917,I244450);
not I_16953 (I293934,I293917);
not I_16954 (I293951,I244459);
nor I_16955 (I293968,I293951,I244435);
and I_16956 (I293985,I293968,I244456);
or I_16957 (I294002,I293985,I244444);
DFFARX1 I_16958  ( .D(I294002), .CLK(I5694_clk), .RSTB(I293773_rst), .Q(I294019) );
nor I_16959 (I294036,I294019,I293872);
nor I_16960 (I294053,I294019,I293934);
nand I_16961 (I293759,I293824,I294053);
nand I_16962 (I294084,I293790,I244459);
nand I_16963 (I294101,I294084,I294019);
and I_16964 (I294118,I294084,I294101);
DFFARX1 I_16965  ( .D(I294118), .CLK(I5694_clk), .RSTB(I293773_rst), .Q(I293741) );
DFFARX1 I_16966  ( .D(I294084), .CLK(I5694_clk), .RSTB(I293773_rst), .Q(I294149) );
and I_16967 (I293738,I293917,I294149);
DFFARX1 I_16968  ( .D(I244465), .CLK(I5694_clk), .RSTB(I293773_rst), .Q(I294180) );
not I_16969 (I294197,I294180);
nor I_16970 (I294214,I293872,I294197);
and I_16971 (I294231,I294180,I294214);
nand I_16972 (I293753,I294180,I293934);
DFFARX1 I_16973  ( .D(I294180), .CLK(I5694_clk), .RSTB(I293773_rst), .Q(I294262) );
not I_16974 (I293750,I294262);
DFFARX1 I_16975  ( .D(I244462), .CLK(I5694_clk), .RSTB(I293773_rst), .Q(I294293) );
not I_16976 (I294310,I294293);
or I_16977 (I294327,I294310,I294231);
DFFARX1 I_16978  ( .D(I294327), .CLK(I5694_clk), .RSTB(I293773_rst), .Q(I293756) );
nand I_16979 (I293765,I294310,I294036);
DFFARX1 I_16980  ( .D(I294310), .CLK(I5694_clk), .RSTB(I293773_rst), .Q(I293735) );
not I_16981 (I294419_rst,I5701);
not I_16982 (I294436,I253701);
nor I_16983 (I294453,I253713,I253695);
nand I_16984 (I294470,I294453,I253710);
DFFARX1 I_16985  ( .D(I294470), .CLK(I5694_clk), .RSTB(I294419_rst), .Q(I294393) );
nor I_16986 (I294501,I294436,I253713);
nand I_16987 (I294518,I294501,I253698);
not I_16988 (I294408,I294518);
DFFARX1 I_16989  ( .D(I294518), .CLK(I5694_clk), .RSTB(I294419_rst), .Q(I294390) );
not I_16990 (I294563,I253713);
not I_16991 (I294580,I294563);
not I_16992 (I294597,I253707);
nor I_16993 (I294614,I294597,I253686);
and I_16994 (I294631,I294614,I253689);
or I_16995 (I294648,I294631,I253692);
DFFARX1 I_16996  ( .D(I294648), .CLK(I5694_clk), .RSTB(I294419_rst), .Q(I294665) );
nor I_16997 (I294682,I294665,I294518);
nor I_16998 (I294699,I294665,I294580);
nand I_16999 (I294405,I294470,I294699);
nand I_17000 (I294730,I294436,I253707);
nand I_17001 (I294747,I294730,I294665);
and I_17002 (I294764,I294730,I294747);
DFFARX1 I_17003  ( .D(I294764), .CLK(I5694_clk), .RSTB(I294419_rst), .Q(I294387) );
DFFARX1 I_17004  ( .D(I294730), .CLK(I5694_clk), .RSTB(I294419_rst), .Q(I294795) );
and I_17005 (I294384,I294563,I294795);
DFFARX1 I_17006  ( .D(I253683), .CLK(I5694_clk), .RSTB(I294419_rst), .Q(I294826) );
not I_17007 (I294843,I294826);
nor I_17008 (I294860,I294518,I294843);
and I_17009 (I294877,I294826,I294860);
nand I_17010 (I294399,I294826,I294580);
DFFARX1 I_17011  ( .D(I294826), .CLK(I5694_clk), .RSTB(I294419_rst), .Q(I294908) );
not I_17012 (I294396,I294908);
DFFARX1 I_17013  ( .D(I253704), .CLK(I5694_clk), .RSTB(I294419_rst), .Q(I294939) );
not I_17014 (I294956,I294939);
or I_17015 (I294973,I294956,I294877);
DFFARX1 I_17016  ( .D(I294973), .CLK(I5694_clk), .RSTB(I294419_rst), .Q(I294402) );
nand I_17017 (I294411,I294956,I294682);
DFFARX1 I_17018  ( .D(I294956), .CLK(I5694_clk), .RSTB(I294419_rst), .Q(I294381) );
not I_17019 (I295065_rst,I5701);
not I_17020 (I295082,I285167);
nor I_17021 (I295099,I285182,I285197);
nand I_17022 (I295116,I295099,I285185);
DFFARX1 I_17023  ( .D(I295116), .CLK(I5694_clk), .RSTB(I295065_rst), .Q(I295039) );
nor I_17024 (I295147,I295082,I285182);
nand I_17025 (I295164,I295147,I285188);
not I_17026 (I295054,I295164);
DFFARX1 I_17027  ( .D(I295164), .CLK(I5694_clk), .RSTB(I295065_rst), .Q(I295036) );
not I_17028 (I295209,I285182);
not I_17029 (I295226,I295209);
not I_17030 (I295243,I285194);
nor I_17031 (I295260,I295243,I285191);
and I_17032 (I295277,I295260,I285170);
or I_17033 (I295294,I295277,I285179);
DFFARX1 I_17034  ( .D(I295294), .CLK(I5694_clk), .RSTB(I295065_rst), .Q(I295311) );
nor I_17035 (I295328,I295311,I295164);
nor I_17036 (I295345,I295311,I295226);
nand I_17037 (I295051,I295116,I295345);
nand I_17038 (I295376,I295082,I285194);
nand I_17039 (I295393,I295376,I295311);
and I_17040 (I295410,I295376,I295393);
DFFARX1 I_17041  ( .D(I295410), .CLK(I5694_clk), .RSTB(I295065_rst), .Q(I295033) );
DFFARX1 I_17042  ( .D(I295376), .CLK(I5694_clk), .RSTB(I295065_rst), .Q(I295441) );
and I_17043 (I295030,I295209,I295441);
DFFARX1 I_17044  ( .D(I285176), .CLK(I5694_clk), .RSTB(I295065_rst), .Q(I295472) );
not I_17045 (I295489,I295472);
nor I_17046 (I295506,I295164,I295489);
and I_17047 (I295523,I295472,I295506);
nand I_17048 (I295045,I295472,I295226);
DFFARX1 I_17049  ( .D(I295472), .CLK(I5694_clk), .RSTB(I295065_rst), .Q(I295554) );
not I_17050 (I295042,I295554);
DFFARX1 I_17051  ( .D(I285173), .CLK(I5694_clk), .RSTB(I295065_rst), .Q(I295585) );
not I_17052 (I295602,I295585);
or I_17053 (I295619,I295602,I295523);
DFFARX1 I_17054  ( .D(I295619), .CLK(I5694_clk), .RSTB(I295065_rst), .Q(I295048) );
nand I_17055 (I295057,I295602,I295328);
DFFARX1 I_17056  ( .D(I295602), .CLK(I5694_clk), .RSTB(I295065_rst), .Q(I295027) );
not I_17057 (I295711_rst,I5701);
not I_17058 (I295728,I272359);
nor I_17059 (I295745,I272335,I272341);
nand I_17060 (I295762,I295745,I272344);
DFFARX1 I_17061  ( .D(I295762), .CLK(I5694_clk), .RSTB(I295711_rst), .Q(I295685) );
nor I_17062 (I295793,I295728,I272335);
nand I_17063 (I295810,I295793,I272353);
not I_17064 (I295700,I295810);
DFFARX1 I_17065  ( .D(I295810), .CLK(I5694_clk), .RSTB(I295711_rst), .Q(I295682) );
not I_17066 (I295855,I272335);
not I_17067 (I295872,I295855);
not I_17068 (I295889,I272332);
nor I_17069 (I295906,I295889,I272347);
and I_17070 (I295923,I295906,I272338);
or I_17071 (I295940,I295923,I272350);
DFFARX1 I_17072  ( .D(I295940), .CLK(I5694_clk), .RSTB(I295711_rst), .Q(I295957) );
nor I_17073 (I295974,I295957,I295810);
nor I_17074 (I295991,I295957,I295872);
nand I_17075 (I295697,I295762,I295991);
nand I_17076 (I296022,I295728,I272332);
nand I_17077 (I296039,I296022,I295957);
and I_17078 (I296056,I296022,I296039);
DFFARX1 I_17079  ( .D(I296056), .CLK(I5694_clk), .RSTB(I295711_rst), .Q(I295679) );
DFFARX1 I_17080  ( .D(I296022), .CLK(I5694_clk), .RSTB(I295711_rst), .Q(I296087) );
and I_17081 (I295676,I295855,I296087);
DFFARX1 I_17082  ( .D(I272362), .CLK(I5694_clk), .RSTB(I295711_rst), .Q(I296118) );
not I_17083 (I296135,I296118);
nor I_17084 (I296152,I295810,I296135);
and I_17085 (I296169,I296118,I296152);
nand I_17086 (I295691,I296118,I295872);
DFFARX1 I_17087  ( .D(I296118), .CLK(I5694_clk), .RSTB(I295711_rst), .Q(I296200) );
not I_17088 (I295688,I296200);
DFFARX1 I_17089  ( .D(I272356), .CLK(I5694_clk), .RSTB(I295711_rst), .Q(I296231) );
not I_17090 (I296248,I296231);
or I_17091 (I296265,I296248,I296169);
DFFARX1 I_17092  ( .D(I296265), .CLK(I5694_clk), .RSTB(I295711_rst), .Q(I295694) );
nand I_17093 (I295703,I296248,I295974);
DFFARX1 I_17094  ( .D(I296248), .CLK(I5694_clk), .RSTB(I295711_rst), .Q(I295673) );
not I_17095 (I296357_rst,I5701);
not I_17096 (I296374,I256285);
nor I_17097 (I296391,I256297,I256279);
nand I_17098 (I296408,I296391,I256294);
DFFARX1 I_17099  ( .D(I296408), .CLK(I5694_clk), .RSTB(I296357_rst), .Q(I296331) );
nor I_17100 (I296439,I296374,I256297);
nand I_17101 (I296456,I296439,I256282);
not I_17102 (I296346,I296456);
DFFARX1 I_17103  ( .D(I296456), .CLK(I5694_clk), .RSTB(I296357_rst), .Q(I296328) );
not I_17104 (I296501,I256297);
not I_17105 (I296518,I296501);
not I_17106 (I296535,I256291);
nor I_17107 (I296552,I296535,I256270);
and I_17108 (I296569,I296552,I256273);
or I_17109 (I296586,I296569,I256276);
DFFARX1 I_17110  ( .D(I296586), .CLK(I5694_clk), .RSTB(I296357_rst), .Q(I296603) );
nor I_17111 (I296620,I296603,I296456);
nor I_17112 (I296637,I296603,I296518);
nand I_17113 (I296343,I296408,I296637);
nand I_17114 (I296668,I296374,I256291);
nand I_17115 (I296685,I296668,I296603);
and I_17116 (I296702,I296668,I296685);
DFFARX1 I_17117  ( .D(I296702), .CLK(I5694_clk), .RSTB(I296357_rst), .Q(I296325) );
DFFARX1 I_17118  ( .D(I296668), .CLK(I5694_clk), .RSTB(I296357_rst), .Q(I296733) );
and I_17119 (I296322,I296501,I296733);
DFFARX1 I_17120  ( .D(I256267), .CLK(I5694_clk), .RSTB(I296357_rst), .Q(I296764) );
not I_17121 (I296781,I296764);
nor I_17122 (I296798,I296456,I296781);
and I_17123 (I296815,I296764,I296798);
nand I_17124 (I296337,I296764,I296518);
DFFARX1 I_17125  ( .D(I296764), .CLK(I5694_clk), .RSTB(I296357_rst), .Q(I296846) );
not I_17126 (I296334,I296846);
DFFARX1 I_17127  ( .D(I256288), .CLK(I5694_clk), .RSTB(I296357_rst), .Q(I296877) );
not I_17128 (I296894,I296877);
or I_17129 (I296911,I296894,I296815);
DFFARX1 I_17130  ( .D(I296911), .CLK(I5694_clk), .RSTB(I296357_rst), .Q(I296340) );
nand I_17131 (I296349,I296894,I296620);
DFFARX1 I_17132  ( .D(I296894), .CLK(I5694_clk), .RSTB(I296357_rst), .Q(I296319) );
not I_17133 (I297003_rst,I5701);
not I_17134 (I297020,I271169);
nor I_17135 (I297037,I271145,I271151);
nand I_17136 (I297054,I297037,I271154);
DFFARX1 I_17137  ( .D(I297054), .CLK(I5694_clk), .RSTB(I297003_rst), .Q(I296977) );
nor I_17138 (I297085,I297020,I271145);
nand I_17139 (I297102,I297085,I271163);
not I_17140 (I296992,I297102);
DFFARX1 I_17141  ( .D(I297102), .CLK(I5694_clk), .RSTB(I297003_rst), .Q(I296974) );
not I_17142 (I297147,I271145);
not I_17143 (I297164,I297147);
not I_17144 (I297181,I271142);
nor I_17145 (I297198,I297181,I271157);
and I_17146 (I297215,I297198,I271148);
or I_17147 (I297232,I297215,I271160);
DFFARX1 I_17148  ( .D(I297232), .CLK(I5694_clk), .RSTB(I297003_rst), .Q(I297249) );
nor I_17149 (I297266,I297249,I297102);
nor I_17150 (I297283,I297249,I297164);
nand I_17151 (I296989,I297054,I297283);
nand I_17152 (I297314,I297020,I271142);
nand I_17153 (I297331,I297314,I297249);
and I_17154 (I297348,I297314,I297331);
DFFARX1 I_17155  ( .D(I297348), .CLK(I5694_clk), .RSTB(I297003_rst), .Q(I296971) );
DFFARX1 I_17156  ( .D(I297314), .CLK(I5694_clk), .RSTB(I297003_rst), .Q(I297379) );
and I_17157 (I296968,I297147,I297379);
DFFARX1 I_17158  ( .D(I271172), .CLK(I5694_clk), .RSTB(I297003_rst), .Q(I297410) );
not I_17159 (I297427,I297410);
nor I_17160 (I297444,I297102,I297427);
and I_17161 (I297461,I297410,I297444);
nand I_17162 (I296983,I297410,I297164);
DFFARX1 I_17163  ( .D(I297410), .CLK(I5694_clk), .RSTB(I297003_rst), .Q(I297492) );
not I_17164 (I296980,I297492);
DFFARX1 I_17165  ( .D(I271166), .CLK(I5694_clk), .RSTB(I297003_rst), .Q(I297523) );
not I_17166 (I297540,I297523);
or I_17167 (I297557,I297540,I297461);
DFFARX1 I_17168  ( .D(I297557), .CLK(I5694_clk), .RSTB(I297003_rst), .Q(I296986) );
nand I_17169 (I296995,I297540,I297266);
DFFARX1 I_17170  ( .D(I297540), .CLK(I5694_clk), .RSTB(I297003_rst), .Q(I296965) );
not I_17171 (I297649_rst,I5701);
not I_17172 (I297666,I274144);
nor I_17173 (I297683,I274120,I274126);
nand I_17174 (I297700,I297683,I274129);
DFFARX1 I_17175  ( .D(I297700), .CLK(I5694_clk), .RSTB(I297649_rst), .Q(I297623) );
nor I_17176 (I297731,I297666,I274120);
nand I_17177 (I297748,I297731,I274138);
not I_17178 (I297638,I297748);
DFFARX1 I_17179  ( .D(I297748), .CLK(I5694_clk), .RSTB(I297649_rst), .Q(I297620) );
not I_17180 (I297793,I274120);
not I_17181 (I297810,I297793);
not I_17182 (I297827,I274117);
nor I_17183 (I297844,I297827,I274132);
and I_17184 (I297861,I297844,I274123);
or I_17185 (I297878,I297861,I274135);
DFFARX1 I_17186  ( .D(I297878), .CLK(I5694_clk), .RSTB(I297649_rst), .Q(I297895) );
nor I_17187 (I297912,I297895,I297748);
nor I_17188 (I297929,I297895,I297810);
nand I_17189 (I297635,I297700,I297929);
nand I_17190 (I297960,I297666,I274117);
nand I_17191 (I297977,I297960,I297895);
and I_17192 (I297994,I297960,I297977);
DFFARX1 I_17193  ( .D(I297994), .CLK(I5694_clk), .RSTB(I297649_rst), .Q(I297617) );
DFFARX1 I_17194  ( .D(I297960), .CLK(I5694_clk), .RSTB(I297649_rst), .Q(I298025) );
and I_17195 (I297614,I297793,I298025);
DFFARX1 I_17196  ( .D(I274147), .CLK(I5694_clk), .RSTB(I297649_rst), .Q(I298056) );
not I_17197 (I298073,I298056);
nor I_17198 (I298090,I297748,I298073);
and I_17199 (I298107,I298056,I298090);
nand I_17200 (I297629,I298056,I297810);
DFFARX1 I_17201  ( .D(I298056), .CLK(I5694_clk), .RSTB(I297649_rst), .Q(I298138) );
not I_17202 (I297626,I298138);
DFFARX1 I_17203  ( .D(I274141), .CLK(I5694_clk), .RSTB(I297649_rst), .Q(I298169) );
not I_17204 (I298186,I298169);
or I_17205 (I298203,I298186,I298107);
DFFARX1 I_17206  ( .D(I298203), .CLK(I5694_clk), .RSTB(I297649_rst), .Q(I297632) );
nand I_17207 (I297641,I298186,I297912);
DFFARX1 I_17208  ( .D(I298186), .CLK(I5694_clk), .RSTB(I297649_rst), .Q(I297611) );
not I_17209 (I298295_rst,I5701);
not I_17210 (I298312,I288689);
nor I_17211 (I298329,I288701,I288686);
nand I_17212 (I298346,I298329,I288698);
DFFARX1 I_17213  ( .D(I298346), .CLK(I5694_clk), .RSTB(I298295_rst), .Q(I298269) );
nor I_17214 (I298377,I298312,I288701);
nand I_17215 (I298394,I298377,I288716);
not I_17216 (I298284,I298394);
DFFARX1 I_17217  ( .D(I298394), .CLK(I5694_clk), .RSTB(I298295_rst), .Q(I298266) );
not I_17218 (I298439,I288701);
not I_17219 (I298456,I298439);
not I_17220 (I298473,I288692);
nor I_17221 (I298490,I298473,I288704);
and I_17222 (I298507,I298490,I288695);
or I_17223 (I298524,I298507,I288710);
DFFARX1 I_17224  ( .D(I298524), .CLK(I5694_clk), .RSTB(I298295_rst), .Q(I298541) );
nor I_17225 (I298558,I298541,I298394);
nor I_17226 (I298575,I298541,I298456);
nand I_17227 (I298281,I298346,I298575);
nand I_17228 (I298606,I298312,I288692);
nand I_17229 (I298623,I298606,I298541);
and I_17230 (I298640,I298606,I298623);
DFFARX1 I_17231  ( .D(I298640), .CLK(I5694_clk), .RSTB(I298295_rst), .Q(I298263) );
DFFARX1 I_17232  ( .D(I298606), .CLK(I5694_clk), .RSTB(I298295_rst), .Q(I298671) );
and I_17233 (I298260,I298439,I298671);
DFFARX1 I_17234  ( .D(I288713), .CLK(I5694_clk), .RSTB(I298295_rst), .Q(I298702) );
not I_17235 (I298719,I298702);
nor I_17236 (I298736,I298394,I298719);
and I_17237 (I298753,I298702,I298736);
nand I_17238 (I298275,I298702,I298456);
DFFARX1 I_17239  ( .D(I298702), .CLK(I5694_clk), .RSTB(I298295_rst), .Q(I298784) );
not I_17240 (I298272,I298784);
DFFARX1 I_17241  ( .D(I288707), .CLK(I5694_clk), .RSTB(I298295_rst), .Q(I298815) );
not I_17242 (I298832,I298815);
or I_17243 (I298849,I298832,I298753);
DFFARX1 I_17244  ( .D(I298849), .CLK(I5694_clk), .RSTB(I298295_rst), .Q(I298278) );
nand I_17245 (I298287,I298832,I298558);
DFFARX1 I_17246  ( .D(I298832), .CLK(I5694_clk), .RSTB(I298295_rst), .Q(I298257) );
not I_17247 (I298941_rst,I5701);
not I_17248 (I298958,I255639);
nor I_17249 (I298975,I255651,I255633);
nand I_17250 (I298992,I298975,I255648);
DFFARX1 I_17251  ( .D(I298992), .CLK(I5694_clk), .RSTB(I298941_rst), .Q(I298915) );
nor I_17252 (I299023,I298958,I255651);
nand I_17253 (I299040,I299023,I255636);
not I_17254 (I298930,I299040);
DFFARX1 I_17255  ( .D(I299040), .CLK(I5694_clk), .RSTB(I298941_rst), .Q(I298912) );
not I_17256 (I299085,I255651);
not I_17257 (I299102,I299085);
not I_17258 (I299119,I255645);
nor I_17259 (I299136,I299119,I255624);
and I_17260 (I299153,I299136,I255627);
or I_17261 (I299170,I299153,I255630);
DFFARX1 I_17262  ( .D(I299170), .CLK(I5694_clk), .RSTB(I298941_rst), .Q(I299187) );
nor I_17263 (I299204,I299187,I299040);
nor I_17264 (I299221,I299187,I299102);
nand I_17265 (I298927,I298992,I299221);
nand I_17266 (I299252,I298958,I255645);
nand I_17267 (I299269,I299252,I299187);
and I_17268 (I299286,I299252,I299269);
DFFARX1 I_17269  ( .D(I299286), .CLK(I5694_clk), .RSTB(I298941_rst), .Q(I298909) );
DFFARX1 I_17270  ( .D(I299252), .CLK(I5694_clk), .RSTB(I298941_rst), .Q(I299317) );
and I_17271 (I298906,I299085,I299317);
DFFARX1 I_17272  ( .D(I255621), .CLK(I5694_clk), .RSTB(I298941_rst), .Q(I299348) );
not I_17273 (I299365,I299348);
nor I_17274 (I299382,I299040,I299365);
and I_17275 (I299399,I299348,I299382);
nand I_17276 (I298921,I299348,I299102);
DFFARX1 I_17277  ( .D(I299348), .CLK(I5694_clk), .RSTB(I298941_rst), .Q(I299430) );
not I_17278 (I298918,I299430);
DFFARX1 I_17279  ( .D(I255642), .CLK(I5694_clk), .RSTB(I298941_rst), .Q(I299461) );
not I_17280 (I299478,I299461);
or I_17281 (I299495,I299478,I299399);
DFFARX1 I_17282  ( .D(I299495), .CLK(I5694_clk), .RSTB(I298941_rst), .Q(I298924) );
nand I_17283 (I298933,I299478,I299204);
DFFARX1 I_17284  ( .D(I299478), .CLK(I5694_clk), .RSTB(I298941_rst), .Q(I298903) );
not I_17285 (I299587_rst,I5701);
not I_17286 (I299604,I277107);
nor I_17287 (I299621,I277092,I277119);
nand I_17288 (I299638,I299621,I277095);
DFFARX1 I_17289  ( .D(I299638), .CLK(I5694_clk), .RSTB(I299587_rst), .Q(I299561) );
nor I_17290 (I299669,I299604,I277092);
nand I_17291 (I299686,I299669,I277110);
not I_17292 (I299576,I299686);
DFFARX1 I_17293  ( .D(I299686), .CLK(I5694_clk), .RSTB(I299587_rst), .Q(I299558) );
not I_17294 (I299731,I277092);
not I_17295 (I299748,I299731);
not I_17296 (I299765,I277122);
nor I_17297 (I299782,I299765,I277104);
and I_17298 (I299799,I299782,I277113);
or I_17299 (I299816,I299799,I277098);
DFFARX1 I_17300  ( .D(I299816), .CLK(I5694_clk), .RSTB(I299587_rst), .Q(I299833) );
nor I_17301 (I299850,I299833,I299686);
nor I_17302 (I299867,I299833,I299748);
nand I_17303 (I299573,I299638,I299867);
nand I_17304 (I299898,I299604,I277122);
nand I_17305 (I299915,I299898,I299833);
and I_17306 (I299932,I299898,I299915);
DFFARX1 I_17307  ( .D(I299932), .CLK(I5694_clk), .RSTB(I299587_rst), .Q(I299555) );
DFFARX1 I_17308  ( .D(I299898), .CLK(I5694_clk), .RSTB(I299587_rst), .Q(I299963) );
and I_17309 (I299552,I299731,I299963);
DFFARX1 I_17310  ( .D(I277101), .CLK(I5694_clk), .RSTB(I299587_rst), .Q(I299994) );
not I_17311 (I300011,I299994);
nor I_17312 (I300028,I299686,I300011);
and I_17313 (I300045,I299994,I300028);
nand I_17314 (I299567,I299994,I299748);
DFFARX1 I_17315  ( .D(I299994), .CLK(I5694_clk), .RSTB(I299587_rst), .Q(I300076) );
not I_17316 (I299564,I300076);
DFFARX1 I_17317  ( .D(I277116), .CLK(I5694_clk), .RSTB(I299587_rst), .Q(I300107) );
not I_17318 (I300124,I300107);
or I_17319 (I300141,I300124,I300045);
DFFARX1 I_17320  ( .D(I300141), .CLK(I5694_clk), .RSTB(I299587_rst), .Q(I299570) );
nand I_17321 (I299579,I300124,I299850);
DFFARX1 I_17322  ( .D(I300124), .CLK(I5694_clk), .RSTB(I299587_rst), .Q(I299549) );
not I_17323 (I300233_rst,I5701);
not I_17324 (I300250,I280764);
nor I_17325 (I300267,I280779,I280794);
nand I_17326 (I300284,I300267,I280782);
DFFARX1 I_17327  ( .D(I300284), .CLK(I5694_clk), .RSTB(I300233_rst), .Q(I300207) );
nor I_17328 (I300315,I300250,I280779);
nand I_17329 (I300332,I300315,I280785);
not I_17330 (I300222,I300332);
DFFARX1 I_17331  ( .D(I300332), .CLK(I5694_clk), .RSTB(I300233_rst), .Q(I300204) );
not I_17332 (I300377,I280779);
not I_17333 (I300394,I300377);
not I_17334 (I300411,I280791);
nor I_17335 (I300428,I300411,I280788);
and I_17336 (I300445,I300428,I280767);
or I_17337 (I300462,I300445,I280776);
DFFARX1 I_17338  ( .D(I300462), .CLK(I5694_clk), .RSTB(I300233_rst), .Q(I300479) );
nor I_17339 (I300496,I300479,I300332);
nor I_17340 (I300513,I300479,I300394);
nand I_17341 (I300219,I300284,I300513);
nand I_17342 (I300544,I300250,I280791);
nand I_17343 (I300561,I300544,I300479);
and I_17344 (I300578,I300544,I300561);
DFFARX1 I_17345  ( .D(I300578), .CLK(I5694_clk), .RSTB(I300233_rst), .Q(I300201) );
DFFARX1 I_17346  ( .D(I300544), .CLK(I5694_clk), .RSTB(I300233_rst), .Q(I300609) );
and I_17347 (I300198,I300377,I300609);
DFFARX1 I_17348  ( .D(I280773), .CLK(I5694_clk), .RSTB(I300233_rst), .Q(I300640) );
not I_17349 (I300657,I300640);
nor I_17350 (I300674,I300332,I300657);
and I_17351 (I300691,I300640,I300674);
nand I_17352 (I300213,I300640,I300394);
DFFARX1 I_17353  ( .D(I300640), .CLK(I5694_clk), .RSTB(I300233_rst), .Q(I300722) );
not I_17354 (I300210,I300722);
DFFARX1 I_17355  ( .D(I280770), .CLK(I5694_clk), .RSTB(I300233_rst), .Q(I300753) );
not I_17356 (I300770,I300753);
or I_17357 (I300787,I300770,I300691);
DFFARX1 I_17358  ( .D(I300787), .CLK(I5694_clk), .RSTB(I300233_rst), .Q(I300216) );
nand I_17359 (I300225,I300770,I300496);
DFFARX1 I_17360  ( .D(I300770), .CLK(I5694_clk), .RSTB(I300233_rst), .Q(I300195) );
not I_17361 (I300879_rst,I5701);
not I_17362 (I300896,I275908);
nor I_17363 (I300913,I275923,I275905);
nand I_17364 (I300930,I300913,I275917);
DFFARX1 I_17365  ( .D(I300930), .CLK(I5694_clk), .RSTB(I300879_rst), .Q(I300850) );
nor I_17366 (I300961,I300896,I275923);
nand I_17367 (I300978,I300961,I275914);
nand I_17368 (I300995,I300978,I300930);
not I_17369 (I301012,I275923);
not I_17370 (I301029,I275932);
nor I_17371 (I301046,I301029,I275902);
and I_17372 (I301063,I301046,I275911);
or I_17373 (I301080,I301063,I275929);
DFFARX1 I_17374  ( .D(I301080), .CLK(I5694_clk), .RSTB(I300879_rst), .Q(I301097) );
nor I_17375 (I301114,I301097,I300978);
nand I_17376 (I300865,I301012,I301114);
not I_17377 (I300862,I301097);
and I_17378 (I301159,I301097,I300995);
DFFARX1 I_17379  ( .D(I301159), .CLK(I5694_clk), .RSTB(I300879_rst), .Q(I300847) );
DFFARX1 I_17380  ( .D(I301097), .CLK(I5694_clk), .RSTB(I300879_rst), .Q(I301190) );
and I_17381 (I300844,I301012,I301190);
nand I_17382 (I301221,I300896,I275932);
not I_17383 (I301238,I301221);
nor I_17384 (I301255,I301097,I301238);
DFFARX1 I_17385  ( .D(I275920), .CLK(I5694_clk), .RSTB(I300879_rst), .Q(I301272) );
nand I_17386 (I301289,I301272,I301221);
and I_17387 (I301306,I301012,I301289);
DFFARX1 I_17388  ( .D(I301306), .CLK(I5694_clk), .RSTB(I300879_rst), .Q(I300871) );
not I_17389 (I301337,I301272);
nand I_17390 (I300859,I301272,I301255);
nand I_17391 (I300853,I301272,I301238);
DFFARX1 I_17392  ( .D(I275926), .CLK(I5694_clk), .RSTB(I300879_rst), .Q(I301382) );
not I_17393 (I301399,I301382);
nor I_17394 (I300868,I301272,I301399);
nor I_17395 (I301430,I301399,I301337);
and I_17396 (I301447,I300978,I301430);
or I_17397 (I301464,I301221,I301447);
DFFARX1 I_17398  ( .D(I301464), .CLK(I5694_clk), .RSTB(I300879_rst), .Q(I300856) );
DFFARX1 I_17399  ( .D(I301399), .CLK(I5694_clk), .RSTB(I300879_rst), .Q(I300841) );
not I_17400 (I301542_rst,I5701);
not I_17401 (I301559,I246424);
nor I_17402 (I301576,I246433,I246445);
nand I_17403 (I301593,I301576,I246436);
DFFARX1 I_17404  ( .D(I301593), .CLK(I5694_clk), .RSTB(I301542_rst), .Q(I301513) );
nor I_17405 (I301624,I301559,I246433);
nand I_17406 (I301641,I301624,I246448);
nand I_17407 (I301658,I301641,I301593);
not I_17408 (I301675,I246433);
not I_17409 (I301692,I246454);
nor I_17410 (I301709,I301692,I246430);
and I_17411 (I301726,I301709,I246439);
or I_17412 (I301743,I301726,I246427);
DFFARX1 I_17413  ( .D(I301743), .CLK(I5694_clk), .RSTB(I301542_rst), .Q(I301760) );
nor I_17414 (I301777,I301760,I301641);
nand I_17415 (I301528,I301675,I301777);
not I_17416 (I301525,I301760);
and I_17417 (I301822,I301760,I301658);
DFFARX1 I_17418  ( .D(I301822), .CLK(I5694_clk), .RSTB(I301542_rst), .Q(I301510) );
DFFARX1 I_17419  ( .D(I301760), .CLK(I5694_clk), .RSTB(I301542_rst), .Q(I301853) );
and I_17420 (I301507,I301675,I301853);
nand I_17421 (I301884,I301559,I246454);
not I_17422 (I301901,I301884);
nor I_17423 (I301918,I301760,I301901);
DFFARX1 I_17424  ( .D(I246451), .CLK(I5694_clk), .RSTB(I301542_rst), .Q(I301935) );
nand I_17425 (I301952,I301935,I301884);
and I_17426 (I301969,I301675,I301952);
DFFARX1 I_17427  ( .D(I301969), .CLK(I5694_clk), .RSTB(I301542_rst), .Q(I301534) );
not I_17428 (I302000,I301935);
nand I_17429 (I301522,I301935,I301918);
nand I_17430 (I301516,I301935,I301901);
DFFARX1 I_17431  ( .D(I246442), .CLK(I5694_clk), .RSTB(I301542_rst), .Q(I302045) );
not I_17432 (I302062,I302045);
nor I_17433 (I301531,I301935,I302062);
nor I_17434 (I302093,I302062,I302000);
and I_17435 (I302110,I301641,I302093);
or I_17436 (I302127,I301884,I302110);
DFFARX1 I_17437  ( .D(I302127), .CLK(I5694_clk), .RSTB(I301542_rst), .Q(I301519) );
DFFARX1 I_17438  ( .D(I302062), .CLK(I5694_clk), .RSTB(I301542_rst), .Q(I301504) );
not I_17439 (I302205_rst,I5701);
not I_17440 (I302222,I293750);
nor I_17441 (I302239,I293738,I293762);
nand I_17442 (I302256,I302239,I293747);
DFFARX1 I_17443  ( .D(I302256), .CLK(I5694_clk), .RSTB(I302205_rst), .Q(I302176) );
nor I_17444 (I302287,I302222,I293738);
nand I_17445 (I302304,I302287,I293765);
nand I_17446 (I302321,I302304,I302256);
not I_17447 (I302338,I293738);
not I_17448 (I302355,I293735);
nor I_17449 (I302372,I302355,I293744);
and I_17450 (I302389,I302372,I293759);
or I_17451 (I302406,I302389,I293741);
DFFARX1 I_17452  ( .D(I302406), .CLK(I5694_clk), .RSTB(I302205_rst), .Q(I302423) );
nor I_17453 (I302440,I302423,I302304);
nand I_17454 (I302191,I302338,I302440);
not I_17455 (I302188,I302423);
and I_17456 (I302485,I302423,I302321);
DFFARX1 I_17457  ( .D(I302485), .CLK(I5694_clk), .RSTB(I302205_rst), .Q(I302173) );
DFFARX1 I_17458  ( .D(I302423), .CLK(I5694_clk), .RSTB(I302205_rst), .Q(I302516) );
and I_17459 (I302170,I302338,I302516);
nand I_17460 (I302547,I302222,I293735);
not I_17461 (I302564,I302547);
nor I_17462 (I302581,I302423,I302564);
DFFARX1 I_17463  ( .D(I293756), .CLK(I5694_clk), .RSTB(I302205_rst), .Q(I302598) );
nand I_17464 (I302615,I302598,I302547);
and I_17465 (I302632,I302338,I302615);
DFFARX1 I_17466  ( .D(I302632), .CLK(I5694_clk), .RSTB(I302205_rst), .Q(I302197) );
not I_17467 (I302663,I302598);
nand I_17468 (I302185,I302598,I302581);
nand I_17469 (I302179,I302598,I302564);
DFFARX1 I_17470  ( .D(I293753), .CLK(I5694_clk), .RSTB(I302205_rst), .Q(I302708) );
not I_17471 (I302725,I302708);
nor I_17472 (I302194,I302598,I302725);
nor I_17473 (I302756,I302725,I302663);
and I_17474 (I302773,I302304,I302756);
or I_17475 (I302790,I302547,I302773);
DFFARX1 I_17476  ( .D(I302790), .CLK(I5694_clk), .RSTB(I302205_rst), .Q(I302182) );
DFFARX1 I_17477  ( .D(I302725), .CLK(I5694_clk), .RSTB(I302205_rst), .Q(I302167) );
not I_17478 (I302868_rst,I5701);
not I_17479 (I302885,I249739);
nor I_17480 (I302902,I249748,I249760);
nand I_17481 (I302919,I302902,I249751);
DFFARX1 I_17482  ( .D(I302919), .CLK(I5694_clk), .RSTB(I302868_rst), .Q(I302839) );
nor I_17483 (I302950,I302885,I249748);
nand I_17484 (I302967,I302950,I249763);
nand I_17485 (I302984,I302967,I302919);
not I_17486 (I303001,I249748);
not I_17487 (I303018,I249769);
nor I_17488 (I303035,I303018,I249745);
and I_17489 (I303052,I303035,I249754);
or I_17490 (I303069,I303052,I249742);
DFFARX1 I_17491  ( .D(I303069), .CLK(I5694_clk), .RSTB(I302868_rst), .Q(I303086) );
nor I_17492 (I303103,I303086,I302967);
nand I_17493 (I302854,I303001,I303103);
not I_17494 (I302851,I303086);
and I_17495 (I303148,I303086,I302984);
DFFARX1 I_17496  ( .D(I303148), .CLK(I5694_clk), .RSTB(I302868_rst), .Q(I302836) );
DFFARX1 I_17497  ( .D(I303086), .CLK(I5694_clk), .RSTB(I302868_rst), .Q(I303179) );
and I_17498 (I302833,I303001,I303179);
nand I_17499 (I303210,I302885,I249769);
not I_17500 (I303227,I303210);
nor I_17501 (I303244,I303086,I303227);
DFFARX1 I_17502  ( .D(I249766), .CLK(I5694_clk), .RSTB(I302868_rst), .Q(I303261) );
nand I_17503 (I303278,I303261,I303210);
and I_17504 (I303295,I303001,I303278);
DFFARX1 I_17505  ( .D(I303295), .CLK(I5694_clk), .RSTB(I302868_rst), .Q(I302860) );
not I_17506 (I303326,I303261);
nand I_17507 (I302848,I303261,I303244);
nand I_17508 (I302842,I303261,I303227);
DFFARX1 I_17509  ( .D(I249757), .CLK(I5694_clk), .RSTB(I302868_rst), .Q(I303371) );
not I_17510 (I303388,I303371);
nor I_17511 (I302857,I303261,I303388);
nor I_17512 (I303419,I303388,I303326);
and I_17513 (I303436,I302967,I303419);
or I_17514 (I303453,I303210,I303436);
DFFARX1 I_17515  ( .D(I303453), .CLK(I5694_clk), .RSTB(I302868_rst), .Q(I302845) );
DFFARX1 I_17516  ( .D(I303388), .CLK(I5694_clk), .RSTB(I302868_rst), .Q(I302830) );
not I_17517 (I303531_rst,I5701);
not I_17518 (I303548,I286976);
nor I_17519 (I303565,I286955,I286967);
nand I_17520 (I303582,I303565,I286961);
DFFARX1 I_17521  ( .D(I303582), .CLK(I5694_clk), .RSTB(I303531_rst), .Q(I303502) );
nor I_17522 (I303613,I303548,I286955);
nand I_17523 (I303630,I303613,I286982);
nand I_17524 (I303647,I303630,I303582);
not I_17525 (I303664,I286955);
not I_17526 (I303681,I286958);
nor I_17527 (I303698,I303681,I286970);
and I_17528 (I303715,I303698,I286973);
or I_17529 (I303732,I303715,I286979);
DFFARX1 I_17530  ( .D(I303732), .CLK(I5694_clk), .RSTB(I303531_rst), .Q(I303749) );
nor I_17531 (I303766,I303749,I303630);
nand I_17532 (I303517,I303664,I303766);
not I_17533 (I303514,I303749);
and I_17534 (I303811,I303749,I303647);
DFFARX1 I_17535  ( .D(I303811), .CLK(I5694_clk), .RSTB(I303531_rst), .Q(I303499) );
DFFARX1 I_17536  ( .D(I303749), .CLK(I5694_clk), .RSTB(I303531_rst), .Q(I303842) );
and I_17537 (I303496,I303664,I303842);
nand I_17538 (I303873,I303548,I286958);
not I_17539 (I303890,I303873);
nor I_17540 (I303907,I303749,I303890);
DFFARX1 I_17541  ( .D(I286952), .CLK(I5694_clk), .RSTB(I303531_rst), .Q(I303924) );
nand I_17542 (I303941,I303924,I303873);
and I_17543 (I303958,I303664,I303941);
DFFARX1 I_17544  ( .D(I303958), .CLK(I5694_clk), .RSTB(I303531_rst), .Q(I303523) );
not I_17545 (I303989,I303924);
nand I_17546 (I303511,I303924,I303907);
nand I_17547 (I303505,I303924,I303890);
DFFARX1 I_17548  ( .D(I286964), .CLK(I5694_clk), .RSTB(I303531_rst), .Q(I304034) );
not I_17549 (I304051,I304034);
nor I_17550 (I303520,I303924,I304051);
nor I_17551 (I304082,I304051,I303989);
and I_17552 (I304099,I303630,I304082);
or I_17553 (I304116,I303873,I304099);
DFFARX1 I_17554  ( .D(I304116), .CLK(I5694_clk), .RSTB(I303531_rst), .Q(I303508) );
DFFARX1 I_17555  ( .D(I304051), .CLK(I5694_clk), .RSTB(I303531_rst), .Q(I303493) );
not I_17556 (I304194_rst,I5701);
or I_17557 (I304211,I289268,I289277);
or I_17558 (I304228,I289271,I289268);
DFFARX1 I_17559  ( .D(I304228), .CLK(I5694_clk), .RSTB(I304194_rst), .Q(I304168) );
nor I_17560 (I304259,I289247,I289250);
not I_17561 (I304276,I304259);
not I_17562 (I304293,I289247);
and I_17563 (I304310,I304293,I289259);
nor I_17564 (I304327,I304310,I289277);
nor I_17565 (I304344,I289265,I289256);
DFFARX1 I_17566  ( .D(I304344), .CLK(I5694_clk), .RSTB(I304194_rst), .Q(I304361) );
nand I_17567 (I304378,I304361,I304211);
and I_17568 (I304395,I304327,I304378);
DFFARX1 I_17569  ( .D(I304395), .CLK(I5694_clk), .RSTB(I304194_rst), .Q(I304162) );
nor I_17570 (I304426,I289265,I289271);
DFFARX1 I_17571  ( .D(I304426), .CLK(I5694_clk), .RSTB(I304194_rst), .Q(I304443) );
and I_17572 (I304159,I304259,I304443);
DFFARX1 I_17573  ( .D(I289262), .CLK(I5694_clk), .RSTB(I304194_rst), .Q(I304474) );
and I_17574 (I304491,I304474,I289253);
DFFARX1 I_17575  ( .D(I304491), .CLK(I5694_clk), .RSTB(I304194_rst), .Q(I304508) );
not I_17576 (I304171,I304508);
DFFARX1 I_17577  ( .D(I304491), .CLK(I5694_clk), .RSTB(I304194_rst), .Q(I304156) );
DFFARX1 I_17578  ( .D(I289274), .CLK(I5694_clk), .RSTB(I304194_rst), .Q(I304553) );
not I_17579 (I304570,I304553);
nor I_17580 (I304587,I304228,I304570);
and I_17581 (I304604,I304491,I304587);
or I_17582 (I304621,I304211,I304604);
DFFARX1 I_17583  ( .D(I304621), .CLK(I5694_clk), .RSTB(I304194_rst), .Q(I304177) );
nor I_17584 (I304652,I304553,I304361);
nand I_17585 (I304186,I304327,I304652);
nor I_17586 (I304683,I304553,I304276);
nand I_17587 (I304180,I304426,I304683);
not I_17588 (I304183,I304553);
nand I_17589 (I304174,I304553,I304276);
DFFARX1 I_17590  ( .D(I304553), .CLK(I5694_clk), .RSTB(I304194_rst), .Q(I304165) );
not I_17591 (I304789_rst,I5701);
or I_17592 (I304806,I298278,I298272);
or I_17593 (I304823,I298266,I298278);
DFFARX1 I_17594  ( .D(I304823), .CLK(I5694_clk), .RSTB(I304789_rst), .Q(I304763) );
nor I_17595 (I304854,I298284,I298275);
not I_17596 (I304871,I304854);
not I_17597 (I304888,I298284);
and I_17598 (I304905,I304888,I298281);
nor I_17599 (I304922,I304905,I298272);
nor I_17600 (I304939,I298257,I298263);
DFFARX1 I_17601  ( .D(I304939), .CLK(I5694_clk), .RSTB(I304789_rst), .Q(I304956) );
nand I_17602 (I304973,I304956,I304806);
and I_17603 (I304990,I304922,I304973);
DFFARX1 I_17604  ( .D(I304990), .CLK(I5694_clk), .RSTB(I304789_rst), .Q(I304757) );
nor I_17605 (I305021,I298257,I298266);
DFFARX1 I_17606  ( .D(I305021), .CLK(I5694_clk), .RSTB(I304789_rst), .Q(I305038) );
and I_17607 (I304754,I304854,I305038);
DFFARX1 I_17608  ( .D(I298269), .CLK(I5694_clk), .RSTB(I304789_rst), .Q(I305069) );
and I_17609 (I305086,I305069,I298287);
DFFARX1 I_17610  ( .D(I305086), .CLK(I5694_clk), .RSTB(I304789_rst), .Q(I305103) );
not I_17611 (I304766,I305103);
DFFARX1 I_17612  ( .D(I305086), .CLK(I5694_clk), .RSTB(I304789_rst), .Q(I304751) );
DFFARX1 I_17613  ( .D(I298260), .CLK(I5694_clk), .RSTB(I304789_rst), .Q(I305148) );
not I_17614 (I305165,I305148);
nor I_17615 (I305182,I304823,I305165);
and I_17616 (I305199,I305086,I305182);
or I_17617 (I305216,I304806,I305199);
DFFARX1 I_17618  ( .D(I305216), .CLK(I5694_clk), .RSTB(I304789_rst), .Q(I304772) );
nor I_17619 (I305247,I305148,I304956);
nand I_17620 (I304781,I304922,I305247);
nor I_17621 (I305278,I305148,I304871);
nand I_17622 (I304775,I305021,I305278);
not I_17623 (I304778,I305148);
nand I_17624 (I304769,I305148,I304871);
DFFARX1 I_17625  ( .D(I305148), .CLK(I5694_clk), .RSTB(I304789_rst), .Q(I304760) );
not I_17626 (I305384_rst,I5701);
or I_17627 (I305401,I269372,I269357);
or I_17628 (I305418,I269378,I269372);
DFFARX1 I_17629  ( .D(I305418), .CLK(I5694_clk), .RSTB(I305384_rst), .Q(I305358) );
nor I_17630 (I305449,I269384,I269366);
not I_17631 (I305466,I305449);
not I_17632 (I305483,I269384);
and I_17633 (I305500,I305483,I269363);
nor I_17634 (I305517,I305500,I269357);
nor I_17635 (I305534,I269360,I269369);
DFFARX1 I_17636  ( .D(I305534), .CLK(I5694_clk), .RSTB(I305384_rst), .Q(I305551) );
nand I_17637 (I305568,I305551,I305401);
and I_17638 (I305585,I305517,I305568);
DFFARX1 I_17639  ( .D(I305585), .CLK(I5694_clk), .RSTB(I305384_rst), .Q(I305352) );
nor I_17640 (I305616,I269360,I269378);
DFFARX1 I_17641  ( .D(I305616), .CLK(I5694_clk), .RSTB(I305384_rst), .Q(I305633) );
and I_17642 (I305349,I305449,I305633);
DFFARX1 I_17643  ( .D(I269387), .CLK(I5694_clk), .RSTB(I305384_rst), .Q(I305664) );
and I_17644 (I305681,I305664,I269375);
DFFARX1 I_17645  ( .D(I305681), .CLK(I5694_clk), .RSTB(I305384_rst), .Q(I305698) );
not I_17646 (I305361,I305698);
DFFARX1 I_17647  ( .D(I305681), .CLK(I5694_clk), .RSTB(I305384_rst), .Q(I305346) );
DFFARX1 I_17648  ( .D(I269381), .CLK(I5694_clk), .RSTB(I305384_rst), .Q(I305743) );
not I_17649 (I305760,I305743);
nor I_17650 (I305777,I305418,I305760);
and I_17651 (I305794,I305681,I305777);
or I_17652 (I305811,I305401,I305794);
DFFARX1 I_17653  ( .D(I305811), .CLK(I5694_clk), .RSTB(I305384_rst), .Q(I305367) );
nor I_17654 (I305842,I305743,I305551);
nand I_17655 (I305376,I305517,I305842);
nor I_17656 (I305873,I305743,I305466);
nand I_17657 (I305370,I305616,I305873);
not I_17658 (I305373,I305743);
nand I_17659 (I305364,I305743,I305466);
DFFARX1 I_17660  ( .D(I305743), .CLK(I5694_clk), .RSTB(I305384_rst), .Q(I305355) );
not I_17661 (I305979_rst,I5701);
or I_17662 (I305996,I290951,I290960);
or I_17663 (I306013,I290954,I290951);
DFFARX1 I_17664  ( .D(I306013), .CLK(I5694_clk), .RSTB(I305979_rst), .Q(I305953) );
nor I_17665 (I306044,I290930,I290933);
not I_17666 (I306061,I306044);
not I_17667 (I306078,I290930);
and I_17668 (I306095,I306078,I290942);
nor I_17669 (I306112,I306095,I290960);
nor I_17670 (I306129,I290948,I290939);
DFFARX1 I_17671  ( .D(I306129), .CLK(I5694_clk), .RSTB(I305979_rst), .Q(I306146) );
nand I_17672 (I306163,I306146,I305996);
and I_17673 (I306180,I306112,I306163);
DFFARX1 I_17674  ( .D(I306180), .CLK(I5694_clk), .RSTB(I305979_rst), .Q(I305947) );
nor I_17675 (I306211,I290948,I290954);
DFFARX1 I_17676  ( .D(I306211), .CLK(I5694_clk), .RSTB(I305979_rst), .Q(I306228) );
and I_17677 (I305944,I306044,I306228);
DFFARX1 I_17678  ( .D(I290945), .CLK(I5694_clk), .RSTB(I305979_rst), .Q(I306259) );
and I_17679 (I306276,I306259,I290936);
DFFARX1 I_17680  ( .D(I306276), .CLK(I5694_clk), .RSTB(I305979_rst), .Q(I306293) );
not I_17681 (I305956,I306293);
DFFARX1 I_17682  ( .D(I306276), .CLK(I5694_clk), .RSTB(I305979_rst), .Q(I305941) );
DFFARX1 I_17683  ( .D(I290957), .CLK(I5694_clk), .RSTB(I305979_rst), .Q(I306338) );
not I_17684 (I306355,I306338);
nor I_17685 (I306372,I306013,I306355);
and I_17686 (I306389,I306276,I306372);
or I_17687 (I306406,I305996,I306389);
DFFARX1 I_17688  ( .D(I306406), .CLK(I5694_clk), .RSTB(I305979_rst), .Q(I305962) );
nor I_17689 (I306437,I306338,I306146);
nand I_17690 (I305971,I306112,I306437);
nor I_17691 (I306468,I306338,I306061);
nand I_17692 (I305965,I306211,I306468);
not I_17693 (I305968,I306338);
nand I_17694 (I305959,I306338,I306061);
DFFARX1 I_17695  ( .D(I306338), .CLK(I5694_clk), .RSTB(I305979_rst), .Q(I305950) );
not I_17696 (I306574_rst,I5701);
or I_17697 (I306591,I267587,I267572);
or I_17698 (I306608,I267593,I267587);
DFFARX1 I_17699  ( .D(I306608), .CLK(I5694_clk), .RSTB(I306574_rst), .Q(I306548) );
nor I_17700 (I306639,I267599,I267581);
not I_17701 (I306656,I306639);
not I_17702 (I306673,I267599);
and I_17703 (I306690,I306673,I267578);
nor I_17704 (I306707,I306690,I267572);
nor I_17705 (I306724,I267575,I267584);
DFFARX1 I_17706  ( .D(I306724), .CLK(I5694_clk), .RSTB(I306574_rst), .Q(I306741) );
nand I_17707 (I306758,I306741,I306591);
and I_17708 (I306775,I306707,I306758);
DFFARX1 I_17709  ( .D(I306775), .CLK(I5694_clk), .RSTB(I306574_rst), .Q(I306542) );
nor I_17710 (I306806,I267575,I267593);
DFFARX1 I_17711  ( .D(I306806), .CLK(I5694_clk), .RSTB(I306574_rst), .Q(I306823) );
and I_17712 (I306539,I306639,I306823);
DFFARX1 I_17713  ( .D(I267602), .CLK(I5694_clk), .RSTB(I306574_rst), .Q(I306854) );
and I_17714 (I306871,I306854,I267590);
DFFARX1 I_17715  ( .D(I306871), .CLK(I5694_clk), .RSTB(I306574_rst), .Q(I306888) );
not I_17716 (I306551,I306888);
DFFARX1 I_17717  ( .D(I306871), .CLK(I5694_clk), .RSTB(I306574_rst), .Q(I306536) );
DFFARX1 I_17718  ( .D(I267596), .CLK(I5694_clk), .RSTB(I306574_rst), .Q(I306933) );
not I_17719 (I306950,I306933);
nor I_17720 (I306967,I306608,I306950);
and I_17721 (I306984,I306871,I306967);
or I_17722 (I307001,I306591,I306984);
DFFARX1 I_17723  ( .D(I307001), .CLK(I5694_clk), .RSTB(I306574_rst), .Q(I306557) );
nor I_17724 (I307032,I306933,I306741);
nand I_17725 (I306566,I306707,I307032);
nor I_17726 (I307063,I306933,I306656);
nand I_17727 (I306560,I306806,I307063);
not I_17728 (I306563,I306933);
nand I_17729 (I306554,I306933,I306656);
DFFARX1 I_17730  ( .D(I306933), .CLK(I5694_clk), .RSTB(I306574_rst), .Q(I306545) );
not I_17731 (I307169_rst,I5701);
or I_17732 (I307186,I248413,I248428);
or I_17733 (I307203,I248416,I248413);
DFFARX1 I_17734  ( .D(I307203), .CLK(I5694_clk), .RSTB(I307169_rst), .Q(I307143) );
nor I_17735 (I307234,I248419,I248434);
not I_17736 (I307251,I307234);
not I_17737 (I307268,I248419);
and I_17738 (I307285,I307268,I248422);
nor I_17739 (I307302,I307285,I248428);
nor I_17740 (I307319,I248425,I248443);
DFFARX1 I_17741  ( .D(I307319), .CLK(I5694_clk), .RSTB(I307169_rst), .Q(I307336) );
nand I_17742 (I307353,I307336,I307186);
and I_17743 (I307370,I307302,I307353);
DFFARX1 I_17744  ( .D(I307370), .CLK(I5694_clk), .RSTB(I307169_rst), .Q(I307137) );
nor I_17745 (I307401,I248425,I248416);
DFFARX1 I_17746  ( .D(I307401), .CLK(I5694_clk), .RSTB(I307169_rst), .Q(I307418) );
and I_17747 (I307134,I307234,I307418);
DFFARX1 I_17748  ( .D(I248440), .CLK(I5694_clk), .RSTB(I307169_rst), .Q(I307449) );
and I_17749 (I307466,I307449,I248431);
DFFARX1 I_17750  ( .D(I307466), .CLK(I5694_clk), .RSTB(I307169_rst), .Q(I307483) );
not I_17751 (I307146,I307483);
DFFARX1 I_17752  ( .D(I307466), .CLK(I5694_clk), .RSTB(I307169_rst), .Q(I307131) );
DFFARX1 I_17753  ( .D(I248437), .CLK(I5694_clk), .RSTB(I307169_rst), .Q(I307528) );
not I_17754 (I307545,I307528);
nor I_17755 (I307562,I307203,I307545);
and I_17756 (I307579,I307466,I307562);
or I_17757 (I307596,I307186,I307579);
DFFARX1 I_17758  ( .D(I307596), .CLK(I5694_clk), .RSTB(I307169_rst), .Q(I307152) );
nor I_17759 (I307627,I307528,I307336);
nand I_17760 (I307161,I307302,I307627);
nor I_17761 (I307658,I307528,I307251);
nand I_17762 (I307155,I307401,I307658);
not I_17763 (I307158,I307528);
nand I_17764 (I307149,I307528,I307251);
DFFARX1 I_17765  ( .D(I307528), .CLK(I5694_clk), .RSTB(I307169_rst), .Q(I307140) );
not I_17766 (I307764_rst,I5701);
or I_17767 (I307781,I272933,I272945);
not I_17768 (I307747,I307781);
DFFARX1 I_17769  ( .D(I307781), .CLK(I5694_clk), .RSTB(I307764_rst), .Q(I307726) );
or I_17770 (I307826,I272957,I272933);
nor I_17771 (I307843,I272951,I272936);
nor I_17772 (I307860,I307843,I307781);
not I_17773 (I307877,I272951);
and I_17774 (I307894,I307877,I272948);
nor I_17775 (I307911,I307894,I272945);
DFFARX1 I_17776  ( .D(I307911), .CLK(I5694_clk), .RSTB(I307764_rst), .Q(I307928) );
nor I_17777 (I307945,I272942,I272939);
DFFARX1 I_17778  ( .D(I307945), .CLK(I5694_clk), .RSTB(I307764_rst), .Q(I307962) );
nor I_17779 (I307753,I307962,I307911);
not I_17780 (I307993,I307962);
nor I_17781 (I308010,I272942,I272957);
nand I_17782 (I308027,I307911,I308010);
and I_17783 (I308044,I307826,I308027);
DFFARX1 I_17784  ( .D(I308044), .CLK(I5694_clk), .RSTB(I307764_rst), .Q(I307756) );
DFFARX1 I_17785  ( .D(I272954), .CLK(I5694_clk), .RSTB(I307764_rst), .Q(I308075) );
and I_17786 (I308092,I308075,I272927);
nor I_17787 (I308109,I308092,I307993);
and I_17788 (I308126,I308010,I308109);
or I_17789 (I308143,I307843,I308126);
DFFARX1 I_17790  ( .D(I308143), .CLK(I5694_clk), .RSTB(I307764_rst), .Q(I307741) );
not I_17791 (I308174,I308092);
nor I_17792 (I308191,I307781,I308174);
nand I_17793 (I307744,I307826,I308191);
nand I_17794 (I307738,I307962,I308174);
DFFARX1 I_17795  ( .D(I308092), .CLK(I5694_clk), .RSTB(I307764_rst), .Q(I307732) );
DFFARX1 I_17796  ( .D(I272930), .CLK(I5694_clk), .RSTB(I307764_rst), .Q(I308250) );
nand I_17797 (I307750,I308250,I307860);
DFFARX1 I_17798  ( .D(I308250), .CLK(I5694_clk), .RSTB(I307764_rst), .Q(I308281) );
not I_17799 (I307735,I308281);
and I_17800 (I307729,I308250,I307928);
not I_17801 (I308359_rst,I5701);
or I_17802 (I308376,I283915,I283924);
not I_17803 (I308342,I308376);
DFFARX1 I_17804  ( .D(I308376), .CLK(I5694_clk), .RSTB(I308359_rst), .Q(I308321) );
or I_17805 (I308421,I283933,I283915);
nor I_17806 (I308438,I283927,I283921);
nor I_17807 (I308455,I308438,I308376);
not I_17808 (I308472,I283927);
and I_17809 (I308489,I308472,I283930);
nor I_17810 (I308506,I308489,I283924);
DFFARX1 I_17811  ( .D(I308506), .CLK(I5694_clk), .RSTB(I308359_rst), .Q(I308523) );
nor I_17812 (I308540,I283918,I283936);
DFFARX1 I_17813  ( .D(I308540), .CLK(I5694_clk), .RSTB(I308359_rst), .Q(I308557) );
nor I_17814 (I308348,I308557,I308506);
not I_17815 (I308588,I308557);
nor I_17816 (I308605,I283918,I283933);
nand I_17817 (I308622,I308506,I308605);
and I_17818 (I308639,I308421,I308622);
DFFARX1 I_17819  ( .D(I308639), .CLK(I5694_clk), .RSTB(I308359_rst), .Q(I308351) );
DFFARX1 I_17820  ( .D(I283939), .CLK(I5694_clk), .RSTB(I308359_rst), .Q(I308670) );
and I_17821 (I308687,I308670,I283912);
nor I_17822 (I308704,I308687,I308588);
and I_17823 (I308721,I308605,I308704);
or I_17824 (I308738,I308438,I308721);
DFFARX1 I_17825  ( .D(I308738), .CLK(I5694_clk), .RSTB(I308359_rst), .Q(I308336) );
not I_17826 (I308769,I308687);
nor I_17827 (I308786,I308376,I308769);
nand I_17828 (I308339,I308421,I308786);
nand I_17829 (I308333,I308557,I308769);
DFFARX1 I_17830  ( .D(I308687), .CLK(I5694_clk), .RSTB(I308359_rst), .Q(I308327) );
DFFARX1 I_17831  ( .D(I283909), .CLK(I5694_clk), .RSTB(I308359_rst), .Q(I308845) );
nand I_17832 (I308345,I308845,I308455);
DFFARX1 I_17833  ( .D(I308845), .CLK(I5694_clk), .RSTB(I308359_rst), .Q(I308876) );
not I_17834 (I308330,I308876);
and I_17835 (I308324,I308845,I308523);
not I_17836 (I308954_rst,I5701);
not I_17837 (I308971,I287542);
nor I_17838 (I308988,I287533,I287539);
nand I_17839 (I309005,I308988,I287551);
nor I_17840 (I309022,I308971,I287533);
nand I_17841 (I309039,I309022,I287536);
not I_17842 (I309056,I309039);
not I_17843 (I309073,I287533);
nor I_17844 (I308943,I309039,I309073);
not I_17845 (I309104,I309073);
nand I_17846 (I308928,I309039,I309104);
not I_17847 (I309135,I287560);
nor I_17848 (I309152,I309135,I287554);
and I_17849 (I309169,I309152,I287545);
or I_17850 (I309186,I309169,I287530);
DFFARX1 I_17851  ( .D(I309186), .CLK(I5694_clk), .RSTB(I308954_rst), .Q(I309203) );
nor I_17852 (I309220,I309203,I309056);
DFFARX1 I_17853  ( .D(I309203), .CLK(I5694_clk), .RSTB(I308954_rst), .Q(I309237) );
not I_17854 (I308925,I309237);
nand I_17855 (I309268,I308971,I287560);
and I_17856 (I309285,I309268,I309220);
DFFARX1 I_17857  ( .D(I309268), .CLK(I5694_clk), .RSTB(I308954_rst), .Q(I308922) );
DFFARX1 I_17858  ( .D(I287548), .CLK(I5694_clk), .RSTB(I308954_rst), .Q(I309316) );
nor I_17859 (I309333,I309316,I309039);
nand I_17860 (I308940,I309203,I309333);
nor I_17861 (I309364,I309316,I309104);
not I_17862 (I308937,I309316);
nand I_17863 (I309395,I309316,I309005);
and I_17864 (I309412,I309073,I309395);
DFFARX1 I_17865  ( .D(I309412), .CLK(I5694_clk), .RSTB(I308954_rst), .Q(I308916) );
DFFARX1 I_17866  ( .D(I309316), .CLK(I5694_clk), .RSTB(I308954_rst), .Q(I308919) );
DFFARX1 I_17867  ( .D(I287557), .CLK(I5694_clk), .RSTB(I308954_rst), .Q(I309457) );
not I_17868 (I309474,I309457);
nand I_17869 (I309491,I309474,I309039);
and I_17870 (I309508,I309268,I309491);
DFFARX1 I_17871  ( .D(I309508), .CLK(I5694_clk), .RSTB(I308954_rst), .Q(I308946) );
or I_17872 (I309539,I309474,I309285);
DFFARX1 I_17873  ( .D(I309539), .CLK(I5694_clk), .RSTB(I308954_rst), .Q(I308931) );
nand I_17874 (I308934,I309474,I309364);
not I_17875 (I309617_rst,I5701);
not I_17876 (I309634,I298909);
nor I_17877 (I309651,I298906,I298930);
nand I_17878 (I309668,I309651,I298927);
nor I_17879 (I309685,I309634,I298906);
nand I_17880 (I309702,I309685,I298933);
not I_17881 (I309719,I309702);
not I_17882 (I309736,I298906);
nor I_17883 (I309606,I309702,I309736);
not I_17884 (I309767,I309736);
nand I_17885 (I309591,I309702,I309767);
not I_17886 (I309798,I298924);
nor I_17887 (I309815,I309798,I298915);
and I_17888 (I309832,I309815,I298912);
or I_17889 (I309849,I309832,I298921);
DFFARX1 I_17890  ( .D(I309849), .CLK(I5694_clk), .RSTB(I309617_rst), .Q(I309866) );
nor I_17891 (I309883,I309866,I309719);
DFFARX1 I_17892  ( .D(I309866), .CLK(I5694_clk), .RSTB(I309617_rst), .Q(I309900) );
not I_17893 (I309588,I309900);
nand I_17894 (I309931,I309634,I298924);
and I_17895 (I309948,I309931,I309883);
DFFARX1 I_17896  ( .D(I309931), .CLK(I5694_clk), .RSTB(I309617_rst), .Q(I309585) );
DFFARX1 I_17897  ( .D(I298903), .CLK(I5694_clk), .RSTB(I309617_rst), .Q(I309979) );
nor I_17898 (I309996,I309979,I309702);
nand I_17899 (I309603,I309866,I309996);
nor I_17900 (I310027,I309979,I309767);
not I_17901 (I309600,I309979);
nand I_17902 (I310058,I309979,I309668);
and I_17903 (I310075,I309736,I310058);
DFFARX1 I_17904  ( .D(I310075), .CLK(I5694_clk), .RSTB(I309617_rst), .Q(I309579) );
DFFARX1 I_17905  ( .D(I309979), .CLK(I5694_clk), .RSTB(I309617_rst), .Q(I309582) );
DFFARX1 I_17906  ( .D(I298918), .CLK(I5694_clk), .RSTB(I309617_rst), .Q(I310120) );
not I_17907 (I310137,I310120);
nand I_17908 (I310154,I310137,I309702);
and I_17909 (I310171,I309931,I310154);
DFFARX1 I_17910  ( .D(I310171), .CLK(I5694_clk), .RSTB(I309617_rst), .Q(I309609) );
or I_17911 (I310202,I310137,I309948);
DFFARX1 I_17912  ( .D(I310202), .CLK(I5694_clk), .RSTB(I309617_rst), .Q(I309594) );
nand I_17913 (I309597,I310137,I310027);
not I_17914 (I310280_rst,I5701);
not I_17915 (I310297,I302170);
nor I_17916 (I310314,I302176,I302182);
nand I_17917 (I310331,I310314,I302185);
nor I_17918 (I310348,I310297,I302176);
nand I_17919 (I310365,I310348,I302167);
not I_17920 (I310382,I310365);
not I_17921 (I310399,I302176);
nor I_17922 (I310269,I310365,I310399);
not I_17923 (I310430,I310399);
nand I_17924 (I310254,I310365,I310430);
not I_17925 (I310461,I302179);
nor I_17926 (I310478,I310461,I302173);
and I_17927 (I310495,I310478,I302188);
or I_17928 (I310512,I310495,I302194);
DFFARX1 I_17929  ( .D(I310512), .CLK(I5694_clk), .RSTB(I310280_rst), .Q(I310529) );
nor I_17930 (I310546,I310529,I310382);
DFFARX1 I_17931  ( .D(I310529), .CLK(I5694_clk), .RSTB(I310280_rst), .Q(I310563) );
not I_17932 (I310251,I310563);
nand I_17933 (I310594,I310297,I302179);
and I_17934 (I310611,I310594,I310546);
DFFARX1 I_17935  ( .D(I310594), .CLK(I5694_clk), .RSTB(I310280_rst), .Q(I310248) );
DFFARX1 I_17936  ( .D(I302191), .CLK(I5694_clk), .RSTB(I310280_rst), .Q(I310642) );
nor I_17937 (I310659,I310642,I310365);
nand I_17938 (I310266,I310529,I310659);
nor I_17939 (I310690,I310642,I310430);
not I_17940 (I310263,I310642);
nand I_17941 (I310721,I310642,I310331);
and I_17942 (I310738,I310399,I310721);
DFFARX1 I_17943  ( .D(I310738), .CLK(I5694_clk), .RSTB(I310280_rst), .Q(I310242) );
DFFARX1 I_17944  ( .D(I310642), .CLK(I5694_clk), .RSTB(I310280_rst), .Q(I310245) );
DFFARX1 I_17945  ( .D(I302197), .CLK(I5694_clk), .RSTB(I310280_rst), .Q(I310783) );
not I_17946 (I310800,I310783);
nand I_17947 (I310817,I310800,I310365);
and I_17948 (I310834,I310594,I310817);
DFFARX1 I_17949  ( .D(I310834), .CLK(I5694_clk), .RSTB(I310280_rst), .Q(I310272) );
or I_17950 (I310865,I310800,I310611);
DFFARX1 I_17951  ( .D(I310865), .CLK(I5694_clk), .RSTB(I310280_rst), .Q(I310257) );
nand I_17952 (I310260,I310800,I310690);
not I_17953 (I310943_rst,I5701);
not I_17954 (I310960,I282657);
nor I_17955 (I310977,I282675,I282666);
nand I_17956 (I310994,I310977,I282672);
nor I_17957 (I311011,I310960,I282675);
nand I_17958 (I311028,I311011,I282678);
not I_17959 (I311045,I311028);
not I_17960 (I311062,I282675);
nor I_17961 (I310932,I311028,I311062);
not I_17962 (I311093,I311062);
nand I_17963 (I310917,I311028,I311093);
not I_17964 (I311124,I282654);
nor I_17965 (I311141,I311124,I282669);
and I_17966 (I311158,I311141,I282651);
or I_17967 (I311175,I311158,I282660);
DFFARX1 I_17968  ( .D(I311175), .CLK(I5694_clk), .RSTB(I310943_rst), .Q(I311192) );
nor I_17969 (I311209,I311192,I311045);
DFFARX1 I_17970  ( .D(I311192), .CLK(I5694_clk), .RSTB(I310943_rst), .Q(I311226) );
not I_17971 (I310914,I311226);
nand I_17972 (I311257,I310960,I282654);
and I_17973 (I311274,I311257,I311209);
DFFARX1 I_17974  ( .D(I311257), .CLK(I5694_clk), .RSTB(I310943_rst), .Q(I310911) );
DFFARX1 I_17975  ( .D(I282663), .CLK(I5694_clk), .RSTB(I310943_rst), .Q(I311305) );
nor I_17976 (I311322,I311305,I311028);
nand I_17977 (I310929,I311192,I311322);
nor I_17978 (I311353,I311305,I311093);
not I_17979 (I310926,I311305);
nand I_17980 (I311384,I311305,I310994);
and I_17981 (I311401,I311062,I311384);
DFFARX1 I_17982  ( .D(I311401), .CLK(I5694_clk), .RSTB(I310943_rst), .Q(I310905) );
DFFARX1 I_17983  ( .D(I311305), .CLK(I5694_clk), .RSTB(I310943_rst), .Q(I310908) );
DFFARX1 I_17984  ( .D(I282681), .CLK(I5694_clk), .RSTB(I310943_rst), .Q(I311446) );
not I_17985 (I311463,I311446);
nand I_17986 (I311480,I311463,I311028);
and I_17987 (I311497,I311257,I311480);
DFFARX1 I_17988  ( .D(I311497), .CLK(I5694_clk), .RSTB(I310943_rst), .Q(I310935) );
or I_17989 (I311528,I311463,I311274);
DFFARX1 I_17990  ( .D(I311528), .CLK(I5694_clk), .RSTB(I310943_rst), .Q(I310920) );
nand I_17991 (I310923,I311463,I311353);
not I_17992 (I311606_rst,I5701);
not I_17993 (I311623,I305959);
nor I_17994 (I311640,I305953,I305944);
nand I_17995 (I311657,I311640,I305956);
nor I_17996 (I311674,I311623,I305953);
nand I_17997 (I311691,I311674,I305971);
not I_17998 (I311708,I311691);
not I_17999 (I311725,I305953);
nor I_18000 (I311595,I311691,I311725);
not I_18001 (I311756,I311725);
nand I_18002 (I311580,I311691,I311756);
not I_18003 (I311787,I305947);
nor I_18004 (I311804,I311787,I305941);
and I_18005 (I311821,I311804,I305968);
or I_18006 (I311838,I311821,I305965);
DFFARX1 I_18007  ( .D(I311838), .CLK(I5694_clk), .RSTB(I311606_rst), .Q(I311855) );
nor I_18008 (I311872,I311855,I311708);
DFFARX1 I_18009  ( .D(I311855), .CLK(I5694_clk), .RSTB(I311606_rst), .Q(I311889) );
not I_18010 (I311577,I311889);
nand I_18011 (I311920,I311623,I305947);
and I_18012 (I311937,I311920,I311872);
DFFARX1 I_18013  ( .D(I311920), .CLK(I5694_clk), .RSTB(I311606_rst), .Q(I311574) );
DFFARX1 I_18014  ( .D(I305962), .CLK(I5694_clk), .RSTB(I311606_rst), .Q(I311968) );
nor I_18015 (I311985,I311968,I311691);
nand I_18016 (I311592,I311855,I311985);
nor I_18017 (I312016,I311968,I311756);
not I_18018 (I311589,I311968);
nand I_18019 (I312047,I311968,I311657);
and I_18020 (I312064,I311725,I312047);
DFFARX1 I_18021  ( .D(I312064), .CLK(I5694_clk), .RSTB(I311606_rst), .Q(I311568) );
DFFARX1 I_18022  ( .D(I311968), .CLK(I5694_clk), .RSTB(I311606_rst), .Q(I311571) );
DFFARX1 I_18023  ( .D(I305950), .CLK(I5694_clk), .RSTB(I311606_rst), .Q(I312109) );
not I_18024 (I312126,I312109);
nand I_18025 (I312143,I312126,I311691);
and I_18026 (I312160,I311920,I312143);
DFFARX1 I_18027  ( .D(I312160), .CLK(I5694_clk), .RSTB(I311606_rst), .Q(I311598) );
or I_18028 (I312191,I312126,I311937);
DFFARX1 I_18029  ( .D(I312191), .CLK(I5694_clk), .RSTB(I311606_rst), .Q(I311583) );
nand I_18030 (I311586,I312126,I312016);
not I_18031 (I312269_rst,I5701);
not I_18032 (I312286,I293192);
nor I_18033 (I312303,I293198,I293201);
nand I_18034 (I312320,I312303,I293177);
nor I_18035 (I312337,I312286,I293198);
nand I_18036 (I312354,I312337,I293186);
not I_18037 (I312371,I312354);
not I_18038 (I312388,I293198);
nor I_18039 (I312258,I312354,I312388);
not I_18040 (I312419,I312388);
nand I_18041 (I312243,I312354,I312419);
not I_18042 (I312450,I293180);
nor I_18043 (I312467,I312450,I293204);
and I_18044 (I312484,I312467,I293174);
or I_18045 (I312501,I312484,I293183);
DFFARX1 I_18046  ( .D(I312501), .CLK(I5694_clk), .RSTB(I312269_rst), .Q(I312518) );
nor I_18047 (I312535,I312518,I312371);
DFFARX1 I_18048  ( .D(I312518), .CLK(I5694_clk), .RSTB(I312269_rst), .Q(I312552) );
not I_18049 (I312240,I312552);
nand I_18050 (I312583,I312286,I293180);
and I_18051 (I312600,I312583,I312535);
DFFARX1 I_18052  ( .D(I312583), .CLK(I5694_clk), .RSTB(I312269_rst), .Q(I312237) );
DFFARX1 I_18053  ( .D(I293189), .CLK(I5694_clk), .RSTB(I312269_rst), .Q(I312631) );
nor I_18054 (I312648,I312631,I312354);
nand I_18055 (I312255,I312518,I312648);
nor I_18056 (I312679,I312631,I312419);
not I_18057 (I312252,I312631);
nand I_18058 (I312710,I312631,I312320);
and I_18059 (I312727,I312388,I312710);
DFFARX1 I_18060  ( .D(I312727), .CLK(I5694_clk), .RSTB(I312269_rst), .Q(I312231) );
DFFARX1 I_18061  ( .D(I312631), .CLK(I5694_clk), .RSTB(I312269_rst), .Q(I312234) );
DFFARX1 I_18062  ( .D(I293195), .CLK(I5694_clk), .RSTB(I312269_rst), .Q(I312772) );
not I_18063 (I312789,I312772);
nand I_18064 (I312806,I312789,I312354);
and I_18065 (I312823,I312583,I312806);
DFFARX1 I_18066  ( .D(I312823), .CLK(I5694_clk), .RSTB(I312269_rst), .Q(I312261) );
or I_18067 (I312854,I312789,I312600);
DFFARX1 I_18068  ( .D(I312854), .CLK(I5694_clk), .RSTB(I312269_rst), .Q(I312246) );
nand I_18069 (I312249,I312789,I312679);
not I_18070 (I312932_rst,I5701);
not I_18071 (I312949,I303496);
nor I_18072 (I312966,I303502,I303508);
nand I_18073 (I312983,I312966,I303511);
nor I_18074 (I313000,I312949,I303502);
nand I_18075 (I313017,I313000,I303493);
not I_18076 (I313034,I313017);
not I_18077 (I313051,I303502);
nor I_18078 (I312921,I313017,I313051);
not I_18079 (I313082,I313051);
nand I_18080 (I312906,I313017,I313082);
not I_18081 (I313113,I303505);
nor I_18082 (I313130,I313113,I303499);
and I_18083 (I313147,I313130,I303514);
or I_18084 (I313164,I313147,I303520);
DFFARX1 I_18085  ( .D(I313164), .CLK(I5694_clk), .RSTB(I312932_rst), .Q(I313181) );
nor I_18086 (I313198,I313181,I313034);
DFFARX1 I_18087  ( .D(I313181), .CLK(I5694_clk), .RSTB(I312932_rst), .Q(I313215) );
not I_18088 (I312903,I313215);
nand I_18089 (I313246,I312949,I303505);
and I_18090 (I313263,I313246,I313198);
DFFARX1 I_18091  ( .D(I313246), .CLK(I5694_clk), .RSTB(I312932_rst), .Q(I312900) );
DFFARX1 I_18092  ( .D(I303517), .CLK(I5694_clk), .RSTB(I312932_rst), .Q(I313294) );
nor I_18093 (I313311,I313294,I313017);
nand I_18094 (I312918,I313181,I313311);
nor I_18095 (I313342,I313294,I313082);
not I_18096 (I312915,I313294);
nand I_18097 (I313373,I313294,I312983);
and I_18098 (I313390,I313051,I313373);
DFFARX1 I_18099  ( .D(I313390), .CLK(I5694_clk), .RSTB(I312932_rst), .Q(I312894) );
DFFARX1 I_18100  ( .D(I313294), .CLK(I5694_clk), .RSTB(I312932_rst), .Q(I312897) );
DFFARX1 I_18101  ( .D(I303523), .CLK(I5694_clk), .RSTB(I312932_rst), .Q(I313435) );
not I_18102 (I313452,I313435);
nand I_18103 (I313469,I313452,I313017);
and I_18104 (I313486,I313246,I313469);
DFFARX1 I_18105  ( .D(I313486), .CLK(I5694_clk), .RSTB(I312932_rst), .Q(I312924) );
or I_18106 (I313517,I313452,I313263);
DFFARX1 I_18107  ( .D(I313517), .CLK(I5694_clk), .RSTB(I312932_rst), .Q(I312909) );
nand I_18108 (I312912,I313452,I313342);
not I_18109 (I313595_rst,I5701);
not I_18110 (I31361_rst2,I254341);
nor I_18111 (I313629,I254338,I254356);
nand I_18112 (I313646,I313629,I254359);
nor I_18113 (I313663,I31361_rst2,I254338);
nand I_18114 (I313680,I313663,I254344);
not I_18115 (I313697,I313680);
not I_18116 (I313714,I254338);
nor I_18117 (I313584,I313680,I313714);
not I_18118 (I313745,I313714);
nand I_18119 (I313569,I313680,I313745);
not I_18120 (I313776,I254353);
nor I_18121 (I313793,I313776,I254335);
and I_18122 (I313810,I313793,I254329);
or I_18123 (I313827,I313810,I254347);
DFFARX1 I_18124  ( .D(I313827), .CLK(I5694_clk), .RSTB(I313595_rst), .Q(I313844) );
nor I_18125 (I313861,I313844,I313697);
DFFARX1 I_18126  ( .D(I313844), .CLK(I5694_clk), .RSTB(I313595_rst), .Q(I313878) );
not I_18127 (I313566,I313878);
nand I_18128 (I313909,I31361_rst2,I254353);
and I_18129 (I313926,I313909,I313861);
DFFARX1 I_18130  ( .D(I313909), .CLK(I5694_clk), .RSTB(I313595_rst), .Q(I313563) );
DFFARX1 I_18131  ( .D(I254332), .CLK(I5694_clk), .RSTB(I313595_rst), .Q(I313957) );
nor I_18132 (I313974,I313957,I313680);
nand I_18133 (I313581,I313844,I313974);
nor I_18134 (I314005,I313957,I313745);
not I_18135 (I313578,I313957);
nand I_18136 (I314036,I313957,I313646);
and I_18137 (I314053,I313714,I314036);
DFFARX1 I_18138  ( .D(I314053), .CLK(I5694_clk), .RSTB(I313595_rst), .Q(I313557) );
DFFARX1 I_18139  ( .D(I313957), .CLK(I5694_clk), .RSTB(I313595_rst), .Q(I313560) );
DFFARX1 I_18140  ( .D(I254350), .CLK(I5694_clk), .RSTB(I313595_rst), .Q(I314098) );
not I_18141 (I314115,I314098);
nand I_18142 (I314132,I314115,I313680);
and I_18143 (I314149,I313909,I314132);
DFFARX1 I_18144  ( .D(I314149), .CLK(I5694_clk), .RSTB(I313595_rst), .Q(I313587) );
or I_18145 (I314180,I314115,I313926);
DFFARX1 I_18146  ( .D(I314180), .CLK(I5694_clk), .RSTB(I313595_rst), .Q(I313572) );
nand I_18147 (I313575,I314115,I314005);
not I_18148 (I314258_rst,I5701);
not I_18149 (I314275,I263524);
nor I_18150 (I314292,I263536,I263518);
nand I_18151 (I314309,I314292,I263539);
nor I_18152 (I314326,I314275,I263536);
nand I_18153 (I314343,I314326,I263530);
not I_18154 (I314360,I314343);
not I_18155 (I314377,I263536);
nor I_18156 (I314247,I314343,I314377);
not I_18157 (I314408,I314377);
nand I_18158 (I314232,I314343,I314408);
not I_18159 (I314439,I263521);
nor I_18160 (I314456,I314439,I263515);
and I_18161 (I314473,I314456,I263527);
or I_18162 (I314490,I314473,I263512);
DFFARX1 I_18163  ( .D(I314490), .CLK(I5694_clk), .RSTB(I314258_rst), .Q(I314507) );
nor I_18164 (I314524,I314507,I314360);
DFFARX1 I_18165  ( .D(I314507), .CLK(I5694_clk), .RSTB(I314258_rst), .Q(I314541) );
not I_18166 (I314229,I314541);
nand I_18167 (I314572,I314275,I263521);
and I_18168 (I314589,I314572,I314524);
DFFARX1 I_18169  ( .D(I314572), .CLK(I5694_clk), .RSTB(I314258_rst), .Q(I314226) );
DFFARX1 I_18170  ( .D(I263509), .CLK(I5694_clk), .RSTB(I314258_rst), .Q(I314620) );
nor I_18171 (I314637,I314620,I314343);
nand I_18172 (I314244,I314507,I314637);
nor I_18173 (I314668,I314620,I314408);
not I_18174 (I314241,I314620);
nand I_18175 (I314699,I314620,I314309);
and I_18176 (I314716,I314377,I314699);
DFFARX1 I_18177  ( .D(I314716), .CLK(I5694_clk), .RSTB(I314258_rst), .Q(I314220) );
DFFARX1 I_18178  ( .D(I314620), .CLK(I5694_clk), .RSTB(I314258_rst), .Q(I314223) );
DFFARX1 I_18179  ( .D(I263533), .CLK(I5694_clk), .RSTB(I314258_rst), .Q(I314761) );
not I_18180 (I314778,I314761);
nand I_18181 (I314795,I314778,I314343);
and I_18182 (I314812,I314572,I314795);
DFFARX1 I_18183  ( .D(I314812), .CLK(I5694_clk), .RSTB(I314258_rst), .Q(I314250) );
or I_18184 (I314843,I314778,I314589);
DFFARX1 I_18185  ( .D(I314843), .CLK(I5694_clk), .RSTB(I314258_rst), .Q(I314235) );
nand I_18186 (I314238,I314778,I314668);
not I_18187 (I314921_rst,I5701);
not I_18188 (I314938,I304174);
nor I_18189 (I314955,I304168,I304159);
nand I_18190 (I314972,I314955,I304171);
nor I_18191 (I314989,I314938,I304168);
nand I_18192 (I315006,I314989,I304186);
not I_18193 (I315023,I315006);
not I_18194 (I315040,I304168);
nor I_18195 (I314910,I315006,I315040);
not I_18196 (I315071,I315040);
nand I_18197 (I314895,I315006,I315071);
not I_18198 (I315102,I304162);
nor I_18199 (I315119,I315102,I304156);
and I_18200 (I315136,I315119,I304183);
or I_18201 (I315153,I315136,I304180);
DFFARX1 I_18202  ( .D(I315153), .CLK(I5694_clk), .RSTB(I314921_rst), .Q(I315170) );
nor I_18203 (I315187,I315170,I315023);
DFFARX1 I_18204  ( .D(I315170), .CLK(I5694_clk), .RSTB(I314921_rst), .Q(I315204) );
not I_18205 (I314892,I315204);
nand I_18206 (I315235,I314938,I304162);
and I_18207 (I315252,I315235,I315187);
DFFARX1 I_18208  ( .D(I315235), .CLK(I5694_clk), .RSTB(I314921_rst), .Q(I314889) );
DFFARX1 I_18209  ( .D(I304177), .CLK(I5694_clk), .RSTB(I314921_rst), .Q(I315283) );
nor I_18210 (I315300,I315283,I315006);
nand I_18211 (I314907,I315170,I315300);
nor I_18212 (I315331,I315283,I315071);
not I_18213 (I314904,I315283);
nand I_18214 (I315362,I315283,I314972);
and I_18215 (I315379,I315040,I315362);
DFFARX1 I_18216  ( .D(I315379), .CLK(I5694_clk), .RSTB(I314921_rst), .Q(I314883) );
DFFARX1 I_18217  ( .D(I315283), .CLK(I5694_clk), .RSTB(I314921_rst), .Q(I314886) );
DFFARX1 I_18218  ( .D(I304165), .CLK(I5694_clk), .RSTB(I314921_rst), .Q(I315424) );
not I_18219 (I315441,I315424);
nand I_18220 (I315458,I315441,I315006);
and I_18221 (I315475,I315235,I315458);
DFFARX1 I_18222  ( .D(I315475), .CLK(I5694_clk), .RSTB(I314921_rst), .Q(I314913) );
or I_18223 (I315506,I315441,I315252);
DFFARX1 I_18224  ( .D(I315506), .CLK(I5694_clk), .RSTB(I314921_rst), .Q(I314898) );
nand I_18225 (I314901,I315441,I315331);
not I_18226 (I315584_rst,I5701);
not I_18227 (I315601,I291509);
nor I_18228 (I315618,I291515,I291518);
nand I_18229 (I315635,I315618,I291494);
nor I_18230 (I315652,I315601,I291515);
nand I_18231 (I315669,I315652,I291503);
not I_18232 (I315686,I315669);
not I_18233 (I315703,I291515);
nor I_18234 (I315573,I315669,I315703);
not I_18235 (I315734,I315703);
nand I_18236 (I315558,I315669,I315734);
not I_18237 (I315765,I291497);
nor I_18238 (I315782,I315765,I291521);
and I_18239 (I315799,I315782,I291491);
or I_18240 (I315816,I315799,I291500);
DFFARX1 I_18241  ( .D(I315816), .CLK(I5694_clk), .RSTB(I315584_rst), .Q(I315833) );
nor I_18242 (I315850,I315833,I315686);
DFFARX1 I_18243  ( .D(I315833), .CLK(I5694_clk), .RSTB(I315584_rst), .Q(I315867) );
not I_18244 (I315555,I315867);
nand I_18245 (I315898,I315601,I291497);
and I_18246 (I315915,I315898,I315850);
DFFARX1 I_18247  ( .D(I315898), .CLK(I5694_clk), .RSTB(I315584_rst), .Q(I315552) );
DFFARX1 I_18248  ( .D(I291506), .CLK(I5694_clk), .RSTB(I315584_rst), .Q(I315946) );
nor I_18249 (I315963,I315946,I315669);
nand I_18250 (I315570,I315833,I315963);
nor I_18251 (I315994,I315946,I315734);
not I_18252 (I315567,I315946);
nand I_18253 (I316025,I315946,I315635);
and I_18254 (I316042,I315703,I316025);
DFFARX1 I_18255  ( .D(I316042), .CLK(I5694_clk), .RSTB(I315584_rst), .Q(I315546) );
DFFARX1 I_18256  ( .D(I315946), .CLK(I5694_clk), .RSTB(I315584_rst), .Q(I315549) );
DFFARX1 I_18257  ( .D(I291512), .CLK(I5694_clk), .RSTB(I315584_rst), .Q(I316087) );
not I_18258 (I316104,I316087);
nand I_18259 (I316121,I316104,I315669);
and I_18260 (I316138,I315898,I316121);
DFFARX1 I_18261  ( .D(I316138), .CLK(I5694_clk), .RSTB(I315584_rst), .Q(I315576) );
or I_18262 (I316169,I316104,I315915);
DFFARX1 I_18263  ( .D(I316169), .CLK(I5694_clk), .RSTB(I315584_rst), .Q(I315561) );
nand I_18264 (I315564,I316104,I315994);
not I_18265 (I316247_rst,I5701);
not I_18266 (I316264,I285814);
nor I_18267 (I316281,I285799,I285805);
nand I_18268 (I316298,I316281,I285802);
nor I_18269 (I316315,I316264,I285799);
nand I_18270 (I316332,I316315,I285811);
DFFARX1 I_18271  ( .D(I316332), .CLK(I5694_clk), .RSTB(I316247_rst), .Q(I316349) );
not I_18272 (I316218,I316349);
not I_18273 (I316380,I285799);
not I_18274 (I316397,I316380);
not I_18275 (I316414,I285826);
nor I_18276 (I316431,I316414,I285820);
and I_18277 (I316448,I316431,I285817);
or I_18278 (I316465,I316448,I285796);
DFFARX1 I_18279  ( .D(I316465), .CLK(I5694_clk), .RSTB(I316247_rst), .Q(I316482) );
DFFARX1 I_18280  ( .D(I316482), .CLK(I5694_clk), .RSTB(I316247_rst), .Q(I316215) );
DFFARX1 I_18281  ( .D(I316482), .CLK(I5694_clk), .RSTB(I316247_rst), .Q(I316513) );
DFFARX1 I_18282  ( .D(I316482), .CLK(I5694_clk), .RSTB(I316247_rst), .Q(I316209) );
nand I_18283 (I316544,I316264,I285826);
nand I_18284 (I316561,I316544,I316298);
and I_18285 (I316578,I316380,I316561);
DFFARX1 I_18286  ( .D(I316578), .CLK(I5694_clk), .RSTB(I316247_rst), .Q(I316239) );
and I_18287 (I316212,I316544,I316513);
DFFARX1 I_18288  ( .D(I285823), .CLK(I5694_clk), .RSTB(I316247_rst), .Q(I316623) );
nor I_18289 (I316236,I316623,I316544);
nor I_18290 (I316654,I316623,I316298);
nand I_18291 (I316233,I316332,I316654);
not I_18292 (I316230,I316623);
DFFARX1 I_18293  ( .D(I285808), .CLK(I5694_clk), .RSTB(I316247_rst), .Q(I316699) );
not I_18294 (I316716,I316699);
nor I_18295 (I316733,I316716,I316397);
and I_18296 (I316750,I316623,I316733);
or I_18297 (I316767,I316544,I316750);
DFFARX1 I_18298  ( .D(I316767), .CLK(I5694_clk), .RSTB(I316247_rst), .Q(I316224) );
not I_18299 (I316798,I316716);
nor I_18300 (I316815,I316623,I316798);
nand I_18301 (I316227,I316716,I316815);
nand I_18302 (I316221,I316380,I316798);
not I_18303 (I316893_rst,I5701);
not I_18304 (I316910,I284559);
nor I_18305 (I316927,I284556,I284541);
nand I_18306 (I316944,I316927,I284550);
nor I_18307 (I316961,I316910,I284556);
nand I_18308 (I316978,I316961,I284565);
DFFARX1 I_18309  ( .D(I316978), .CLK(I5694_clk), .RSTB(I316893_rst), .Q(I316995) );
not I_18310 (I316864,I316995);
not I_18311 (I317026,I284556);
not I_18312 (I317043,I317026);
not I_18313 (I317060,I284538);
nor I_18314 (I317077,I317060,I284544);
and I_18315 (I317094,I317077,I284568);
or I_18316 (I317111,I317094,I284562);
DFFARX1 I_18317  ( .D(I317111), .CLK(I5694_clk), .RSTB(I316893_rst), .Q(I317128) );
DFFARX1 I_18318  ( .D(I317128), .CLK(I5694_clk), .RSTB(I316893_rst), .Q(I316861) );
DFFARX1 I_18319  ( .D(I317128), .CLK(I5694_clk), .RSTB(I316893_rst), .Q(I317159) );
DFFARX1 I_18320  ( .D(I317128), .CLK(I5694_clk), .RSTB(I316893_rst), .Q(I316855) );
nand I_18321 (I317190,I316910,I284538);
nand I_18322 (I317207,I317190,I316944);
and I_18323 (I317224,I317026,I317207);
DFFARX1 I_18324  ( .D(I317224), .CLK(I5694_clk), .RSTB(I316893_rst), .Q(I316885) );
and I_18325 (I316858,I317190,I317159);
DFFARX1 I_18326  ( .D(I284547), .CLK(I5694_clk), .RSTB(I316893_rst), .Q(I317269) );
nor I_18327 (I316882,I317269,I317190);
nor I_18328 (I317300,I317269,I316944);
nand I_18329 (I316879,I316978,I317300);
not I_18330 (I316876,I317269);
DFFARX1 I_18331  ( .D(I284553), .CLK(I5694_clk), .RSTB(I316893_rst), .Q(I317345) );
not I_18332 (I317362,I317345);
nor I_18333 (I317379,I317362,I317043);
and I_18334 (I317396,I317269,I317379);
or I_18335 (I317413,I317190,I317396);
DFFARX1 I_18336  ( .D(I317413), .CLK(I5694_clk), .RSTB(I316893_rst), .Q(I316870) );
not I_18337 (I317444,I317362);
nor I_18338 (I317461,I317269,I317444);
nand I_18339 (I316873,I317362,I317461);
nand I_18340 (I316867,I317026,I317444);
not I_18341 (I317539_rst,I5701);
not I_18342 (I317556,I265258);
nor I_18343 (I317573,I265261,I265243);
nand I_18344 (I317590,I317573,I265270);
nor I_18345 (I317607,I317556,I265261);
nand I_18346 (I317624,I317607,I265249);
DFFARX1 I_18347  ( .D(I317624), .CLK(I5694_clk), .RSTB(I317539_rst), .Q(I317641) );
not I_18348 (I317510,I317641);
not I_18349 (I317672,I265261);
not I_18350 (I317689,I317672);
not I_18351 (I317706,I265255);
nor I_18352 (I317723,I317706,I265267);
and I_18353 (I317740,I317723,I265273);
or I_18354 (I317757,I317740,I265252);
DFFARX1 I_18355  ( .D(I317757), .CLK(I5694_clk), .RSTB(I317539_rst), .Q(I317774) );
DFFARX1 I_18356  ( .D(I317774), .CLK(I5694_clk), .RSTB(I317539_rst), .Q(I317507) );
DFFARX1 I_18357  ( .D(I317774), .CLK(I5694_clk), .RSTB(I317539_rst), .Q(I317805) );
DFFARX1 I_18358  ( .D(I317774), .CLK(I5694_clk), .RSTB(I317539_rst), .Q(I317501) );
nand I_18359 (I317836,I317556,I265255);
nand I_18360 (I317853,I317836,I317590);
and I_18361 (I317870,I317672,I317853);
DFFARX1 I_18362  ( .D(I317870), .CLK(I5694_clk), .RSTB(I317539_rst), .Q(I317531) );
and I_18363 (I317504,I317836,I317805);
DFFARX1 I_18364  ( .D(I265264), .CLK(I5694_clk), .RSTB(I317539_rst), .Q(I317915) );
nor I_18365 (I317528,I317915,I317836);
nor I_18366 (I317946,I317915,I317590);
nand I_18367 (I317525,I317624,I317946);
not I_18368 (I317522,I317915);
DFFARX1 I_18369  ( .D(I265246), .CLK(I5694_clk), .RSTB(I317539_rst), .Q(I317991) );
not I_18370 (I318008,I317991);
nor I_18371 (I318025,I318008,I317689);
and I_18372 (I318042,I317915,I318025);
or I_18373 (I318059,I317836,I318042);
DFFARX1 I_18374  ( .D(I318059), .CLK(I5694_clk), .RSTB(I317539_rst), .Q(I317516) );
not I_18375 (I318090,I318008);
nor I_18376 (I318107,I317915,I318090);
nand I_18377 (I317519,I318008,I318107);
nand I_18378 (I317513,I317672,I318090);
not I_18379 (I318185_rst,I5701);
not I_18380 (I318202,I258869);
nor I_18381 (I318219,I258878,I258863);
nand I_18382 (I318236,I318219,I258851);
nor I_18383 (I318253,I318202,I258878);
nand I_18384 (I318270,I318253,I258854);
DFFARX1 I_18385  ( .D(I318270), .CLK(I5694_clk), .RSTB(I318185_rst), .Q(I318287) );
not I_18386 (I318156,I318287);
not I_18387 (I318318,I258878);
not I_18388 (I318335,I318318);
not I_18389 (I318352,I258866);
nor I_18390 (I318369,I318352,I258860);
and I_18391 (I318386,I318369,I258857);
or I_18392 (I318403,I318386,I258872);
DFFARX1 I_18393  ( .D(I318403), .CLK(I5694_clk), .RSTB(I318185_rst), .Q(I318420) );
DFFARX1 I_18394  ( .D(I318420), .CLK(I5694_clk), .RSTB(I318185_rst), .Q(I318153) );
DFFARX1 I_18395  ( .D(I318420), .CLK(I5694_clk), .RSTB(I318185_rst), .Q(I318451) );
DFFARX1 I_18396  ( .D(I318420), .CLK(I5694_clk), .RSTB(I318185_rst), .Q(I318147) );
nand I_18397 (I318482,I318202,I258866);
nand I_18398 (I318499,I318482,I318236);
and I_18399 (I318516,I318318,I318499);
DFFARX1 I_18400  ( .D(I318516), .CLK(I5694_clk), .RSTB(I318185_rst), .Q(I318177) );
and I_18401 (I318150,I318482,I318451);
DFFARX1 I_18402  ( .D(I258881), .CLK(I5694_clk), .RSTB(I318185_rst), .Q(I318561) );
nor I_18403 (I318174,I318561,I318482);
nor I_18404 (I318592,I318561,I318236);
nand I_18405 (I318171,I318270,I318592);
not I_18406 (I318168,I318561);
DFFARX1 I_18407  ( .D(I258875), .CLK(I5694_clk), .RSTB(I318185_rst), .Q(I318637) );
not I_18408 (I318654,I318637);
nor I_18409 (I318671,I318654,I318335);
and I_18410 (I318688,I318561,I318671);
or I_18411 (I318705,I318482,I318688);
DFFARX1 I_18412  ( .D(I318705), .CLK(I5694_clk), .RSTB(I318185_rst), .Q(I318162) );
not I_18413 (I318736,I318654);
nor I_18414 (I318753,I318561,I318736);
nand I_18415 (I318165,I318654,I318753);
nand I_18416 (I318159,I318318,I318736);
not I_18417 (I318831_rst,I5701);
not I_18418 (I318848,I290378);
nor I_18419 (I318865,I290393,I290387);
nand I_18420 (I318882,I318865,I290396);
nor I_18421 (I318899,I318848,I290393);
nand I_18422 (I318916,I318899,I290372);
DFFARX1 I_18423  ( .D(I318916), .CLK(I5694_clk), .RSTB(I318831_rst), .Q(I318933) );
not I_18424 (I318802,I318933);
not I_18425 (I318964,I290393);
not I_18426 (I318981,I318964);
not I_18427 (I318998,I290369);
nor I_18428 (I319015,I318998,I290384);
and I_18429 (I319032,I319015,I290390);
or I_18430 (I319049,I319032,I290399);
DFFARX1 I_18431  ( .D(I319049), .CLK(I5694_clk), .RSTB(I318831_rst), .Q(I319066) );
DFFARX1 I_18432  ( .D(I319066), .CLK(I5694_clk), .RSTB(I318831_rst), .Q(I318799) );
DFFARX1 I_18433  ( .D(I319066), .CLK(I5694_clk), .RSTB(I318831_rst), .Q(I319097) );
DFFARX1 I_18434  ( .D(I319066), .CLK(I5694_clk), .RSTB(I318831_rst), .Q(I318793) );
nand I_18435 (I319128,I318848,I290369);
nand I_18436 (I319145,I319128,I318882);
and I_18437 (I319162,I318964,I319145);
DFFARX1 I_18438  ( .D(I319162), .CLK(I5694_clk), .RSTB(I318831_rst), .Q(I318823) );
and I_18439 (I318796,I319128,I319097);
DFFARX1 I_18440  ( .D(I290381), .CLK(I5694_clk), .RSTB(I318831_rst), .Q(I319207) );
nor I_18441 (I318820,I319207,I319128);
nor I_18442 (I319238,I319207,I318882);
nand I_18443 (I318817,I318916,I319238);
not I_18444 (I318814,I319207);
DFFARX1 I_18445  ( .D(I290375), .CLK(I5694_clk), .RSTB(I318831_rst), .Q(I319283) );
not I_18446 (I319300,I319283);
nor I_18447 (I319317,I319300,I318981);
and I_18448 (I319334,I319207,I319317);
or I_18449 (I319351,I319128,I319334);
DFFARX1 I_18450  ( .D(I319351), .CLK(I5694_clk), .RSTB(I318831_rst), .Q(I318808) );
not I_18451 (I319382,I319300);
nor I_18452 (I319399,I319207,I319382);
nand I_18453 (I318811,I319300,I319399);
nand I_18454 (I318805,I318964,I319382);
not I_18455 (I319477_rst,I5701);
not I_18456 (I319494,I275325);
nor I_18457 (I319511,I275313,I275322);
nand I_18458 (I319528,I319511,I275337);
nor I_18459 (I319545,I319494,I275313);
nand I_18460 (I319562,I319545,I275319);
DFFARX1 I_18461  ( .D(I319562), .CLK(I5694_clk), .RSTB(I319477_rst), .Q(I319579) );
not I_18462 (I319448,I319579);
not I_18463 (I319610,I275313);
not I_18464 (I319627,I319610);
not I_18465 (I319644,I275307);
nor I_18466 (I319661,I319644,I275328);
and I_18467 (I319678,I319661,I275310);
or I_18468 (I319695,I319678,I275316);
DFFARX1 I_18469  ( .D(I319695), .CLK(I5694_clk), .RSTB(I319477_rst), .Q(I319712) );
DFFARX1 I_18470  ( .D(I319712), .CLK(I5694_clk), .RSTB(I319477_rst), .Q(I319445) );
DFFARX1 I_18471  ( .D(I319712), .CLK(I5694_clk), .RSTB(I319477_rst), .Q(I319743) );
DFFARX1 I_18472  ( .D(I319712), .CLK(I5694_clk), .RSTB(I319477_rst), .Q(I319439) );
nand I_18473 (I319774,I319494,I275307);
nand I_18474 (I319791,I319774,I319528);
and I_18475 (I319808,I319610,I319791);
DFFARX1 I_18476  ( .D(I319808), .CLK(I5694_clk), .RSTB(I319477_rst), .Q(I319469) );
and I_18477 (I319442,I319774,I319743);
DFFARX1 I_18478  ( .D(I275334), .CLK(I5694_clk), .RSTB(I319477_rst), .Q(I319853) );
nor I_18479 (I319466,I319853,I319774);
nor I_18480 (I319884,I319853,I319528);
nand I_18481 (I319463,I319562,I319884);
not I_18482 (I319460,I319853);
DFFARX1 I_18483  ( .D(I275331), .CLK(I5694_clk), .RSTB(I319477_rst), .Q(I319929) );
not I_18484 (I319946,I319929);
nor I_18485 (I319963,I319946,I319627);
and I_18486 (I319980,I319853,I319963);
or I_18487 (I319997,I319774,I319980);
DFFARX1 I_18488  ( .D(I319997), .CLK(I5694_clk), .RSTB(I319477_rst), .Q(I319454) );
not I_18489 (I320028,I319946);
nor I_18490 (I320045,I319853,I320028);
nand I_18491 (I319457,I319946,I320045);
nand I_18492 (I319451,I319610,I320028);
not I_18493 (I320123_rst,I5701);
not I_18494 (I320140,I278898);
nor I_18495 (I320157,I278895,I278880);
nand I_18496 (I320174,I320157,I278889);
nor I_18497 (I320191,I320140,I278895);
nand I_18498 (I320208,I320191,I278904);
DFFARX1 I_18499  ( .D(I320208), .CLK(I5694_clk), .RSTB(I320123_rst), .Q(I320225) );
not I_18500 (I320094,I320225);
not I_18501 (I320256,I278895);
not I_18502 (I320273,I320256);
not I_18503 (I320290,I278877);
nor I_18504 (I320307,I320290,I278883);
and I_18505 (I320324,I320307,I278907);
or I_18506 (I320341,I320324,I278901);
DFFARX1 I_18507  ( .D(I320341), .CLK(I5694_clk), .RSTB(I320123_rst), .Q(I320358) );
DFFARX1 I_18508  ( .D(I320358), .CLK(I5694_clk), .RSTB(I320123_rst), .Q(I320091) );
DFFARX1 I_18509  ( .D(I320358), .CLK(I5694_clk), .RSTB(I320123_rst), .Q(I320389) );
DFFARX1 I_18510  ( .D(I320358), .CLK(I5694_clk), .RSTB(I320123_rst), .Q(I320085) );
nand I_18511 (I320420,I320140,I278877);
nand I_18512 (I320437,I320420,I320174);
and I_18513 (I320454,I320256,I320437);
DFFARX1 I_18514  ( .D(I320454), .CLK(I5694_clk), .RSTB(I320123_rst), .Q(I320115) );
and I_18515 (I320088,I320420,I320389);
DFFARX1 I_18516  ( .D(I278886), .CLK(I5694_clk), .RSTB(I320123_rst), .Q(I320499) );
nor I_18517 (I320112,I320499,I320420);
nor I_18518 (I320530,I320499,I320174);
nand I_18519 (I320109,I320208,I320530);
not I_18520 (I320106,I320499);
DFFARX1 I_18521  ( .D(I278892), .CLK(I5694_clk), .RSTB(I320123_rst), .Q(I320575) );
not I_18522 (I320592,I320575);
nor I_18523 (I320609,I320592,I320273);
and I_18524 (I320626,I320499,I320609);
or I_18525 (I320643,I320420,I320626);
DFFARX1 I_18526  ( .D(I320643), .CLK(I5694_clk), .RSTB(I320123_rst), .Q(I320100) );
not I_18527 (I320674,I320592);
nor I_18528 (I320691,I320499,I320674);
nand I_18529 (I320103,I320592,I320691);
nand I_18530 (I320097,I320256,I320674);
not I_18531 (I320769_rst,I5701);
or I_18532 (I320786,I317516,I317528);
or I_18533 (I320803,I317510,I317516);
nor I_18534 (I320820,I317531,I317507);
DFFARX1 I_18535  ( .D(I320820), .CLK(I5694_clk), .RSTB(I320769_rst), .Q(I320837) );
DFFARX1 I_18536  ( .D(I320820), .CLK(I5694_clk), .RSTB(I320769_rst), .Q(I320731) );
not I_18537 (I320868,I317531);
and I_18538 (I320885,I320868,I317522);
nor I_18539 (I320902,I320885,I317528);
nor I_18540 (I320919,I317501,I317519);
DFFARX1 I_18541  ( .D(I320919), .CLK(I5694_clk), .RSTB(I320769_rst), .Q(I320936) );
not I_18542 (I320953,I320936);
DFFARX1 I_18543  ( .D(I320936), .CLK(I5694_clk), .RSTB(I320769_rst), .Q(I320740) );
nor I_18544 (I320984,I317501,I317510);
and I_18545 (I320734,I320984,I320837);
DFFARX1 I_18546  ( .D(I317525), .CLK(I5694_clk), .RSTB(I320769_rst), .Q(I321015) );
and I_18547 (I321032,I321015,I317504);
nand I_18548 (I321049,I321032,I320803);
and I_18549 (I321066,I320936,I321049);
DFFARX1 I_18550  ( .D(I321066), .CLK(I5694_clk), .RSTB(I320769_rst), .Q(I320761) );
nor I_18551 (I320758,I321032,I320902);
not I_18552 (I321111,I321032);
nor I_18553 (I321128,I320786,I321111);
nor I_18554 (I321145,I321032,I320984);
nand I_18555 (I320755,I320803,I321145);
nor I_18556 (I321176,I321032,I320953);
not I_18557 (I320752,I321032);
nand I_18558 (I320743,I321032,I320953);
DFFARX1 I_18559  ( .D(I317513), .CLK(I5694_clk), .RSTB(I320769_rst), .Q(I321221) );
and I_18560 (I321238,I321221,I321128);
or I_18561 (I321255,I320786,I321238);
DFFARX1 I_18562  ( .D(I321255), .CLK(I5694_clk), .RSTB(I320769_rst), .Q(I320746) );
nand I_18563 (I320749,I321221,I321176);
nand I_18564 (I321300,I321221,I320902);
and I_18565 (I321317,I320820,I321300);
DFFARX1 I_18566  ( .D(I321317), .CLK(I5694_clk), .RSTB(I320769_rst), .Q(I320737) );
not I_18567 (I321381_rst,I5701);
nand I_18568 (I321398,I274739,I274727);
and I_18569 (I321415,I321398,I274721);
DFFARX1 I_18570  ( .D(I321415), .CLK(I5694_clk), .RSTB(I321381_rst), .Q(I321432) );
not I_18571 (I321449,I321432);
DFFARX1 I_18572  ( .D(I321432), .CLK(I5694_clk), .RSTB(I321381_rst), .Q(I321349) );
nor I_18573 (I321480,I274718,I274727);
DFFARX1 I_18574  ( .D(I274712), .CLK(I5694_clk), .RSTB(I321381_rst), .Q(I321497) );
DFFARX1 I_18575  ( .D(I321497), .CLK(I5694_clk), .RSTB(I321381_rst), .Q(I321514) );
not I_18576 (I321352,I321514);
DFFARX1 I_18577  ( .D(I321497), .CLK(I5694_clk), .RSTB(I321381_rst), .Q(I321545) );
and I_18578 (I321346,I321432,I321545);
nand I_18579 (I321576,I274715,I274730);
and I_18580 (I321593,I321576,I274742);
DFFARX1 I_18581  ( .D(I321593), .CLK(I5694_clk), .RSTB(I321381_rst), .Q(I321610) );
nor I_18582 (I321627,I321610,I321449);
not I_18583 (I321644,I321610);
nand I_18584 (I321355,I321432,I321644);
DFFARX1 I_18585  ( .D(I274733), .CLK(I5694_clk), .RSTB(I321381_rst), .Q(I321675) );
and I_18586 (I321692,I321675,I274724);
nor I_18587 (I321709,I321692,I321610);
nor I_18588 (I321726,I321692,I321644);
nand I_18589 (I321361,I321480,I321726);
not I_18590 (I321364,I321692);
DFFARX1 I_18591  ( .D(I321692), .CLK(I5694_clk), .RSTB(I321381_rst), .Q(I321343) );
DFFARX1 I_18592  ( .D(I274736), .CLK(I5694_clk), .RSTB(I321381_rst), .Q(I321785) );
nand I_18593 (I321802,I321785,I321497);
and I_18594 (I321819,I321480,I321802);
DFFARX1 I_18595  ( .D(I321819), .CLK(I5694_clk), .RSTB(I321381_rst), .Q(I321373) );
nor I_18596 (I321370,I321785,I321692);
and I_18597 (I321864,I321785,I321627);
or I_18598 (I321881,I321480,I321864);
DFFARX1 I_18599  ( .D(I321881), .CLK(I5694_clk), .RSTB(I321381_rst), .Q(I321358) );
nand I_18600 (I321367,I321785,I321709);
not I_18601 (I321959_rst,I5701);
nand I_18602 (I321976,I320100,I320097);
and I_18603 (I321993,I321976,I320109);
DFFARX1 I_18604  ( .D(I321993), .CLK(I5694_clk), .RSTB(I321959_rst), .Q(I322010) );
not I_18605 (I322027,I322010);
DFFARX1 I_18606  ( .D(I322010), .CLK(I5694_clk), .RSTB(I321959_rst), .Q(I321927) );
nor I_18607 (I322058,I320106,I320097);
DFFARX1 I_18608  ( .D(I320112), .CLK(I5694_clk), .RSTB(I321959_rst), .Q(I322075) );
DFFARX1 I_18609  ( .D(I322075), .CLK(I5694_clk), .RSTB(I321959_rst), .Q(I322092) );
not I_18610 (I321930,I322092);
DFFARX1 I_18611  ( .D(I322075), .CLK(I5694_clk), .RSTB(I321959_rst), .Q(I322123) );
and I_18612 (I321924,I322010,I322123);
nand I_18613 (I322154,I320088,I320091);
and I_18614 (I322171,I322154,I320115);
DFFARX1 I_18615  ( .D(I322171), .CLK(I5694_clk), .RSTB(I321959_rst), .Q(I322188) );
nor I_18616 (I322205,I322188,I322027);
not I_18617 (I322222,I322188);
nand I_18618 (I321933,I322010,I322222);
DFFARX1 I_18619  ( .D(I320094), .CLK(I5694_clk), .RSTB(I321959_rst), .Q(I322253) );
and I_18620 (I322270,I322253,I320085);
nor I_18621 (I322287,I322270,I322188);
nor I_18622 (I322304,I322270,I322222);
nand I_18623 (I321939,I322058,I322304);
not I_18624 (I321942,I322270);
DFFARX1 I_18625  ( .D(I322270), .CLK(I5694_clk), .RSTB(I321959_rst), .Q(I321921) );
DFFARX1 I_18626  ( .D(I320103), .CLK(I5694_clk), .RSTB(I321959_rst), .Q(I322363) );
nand I_18627 (I322380,I322363,I322075);
and I_18628 (I322397,I322058,I322380);
DFFARX1 I_18629  ( .D(I322397), .CLK(I5694_clk), .RSTB(I321959_rst), .Q(I321951) );
nor I_18630 (I321948,I322363,I322270);
and I_18631 (I322442,I322363,I322205);
or I_18632 (I322459,I322058,I322442);
DFFARX1 I_18633  ( .D(I322459), .CLK(I5694_clk), .RSTB(I321959_rst), .Q(I321936) );
nand I_18634 (I321945,I322363,I322287);
not I_18635 (I322537_rst,I5701);
nand I_18636 (I322554,I308919,I308946);
and I_18637 (I322571,I322554,I308934);
DFFARX1 I_18638  ( .D(I322571), .CLK(I5694_clk), .RSTB(I322537_rst), .Q(I322588) );
not I_18639 (I322605,I322588);
DFFARX1 I_18640  ( .D(I322588), .CLK(I5694_clk), .RSTB(I322537_rst), .Q(I322505) );
nor I_18641 (I322636,I308922,I308946);
DFFARX1 I_18642  ( .D(I308937), .CLK(I5694_clk), .RSTB(I322537_rst), .Q(I322653) );
DFFARX1 I_18643  ( .D(I322653), .CLK(I5694_clk), .RSTB(I322537_rst), .Q(I322670) );
not I_18644 (I322508,I322670);
DFFARX1 I_18645  ( .D(I322653), .CLK(I5694_clk), .RSTB(I322537_rst), .Q(I322701) );
and I_18646 (I322502,I322588,I322701);
nand I_18647 (I322732,I308931,I308928);
and I_18648 (I322749,I322732,I308925);
DFFARX1 I_18649  ( .D(I322749), .CLK(I5694_clk), .RSTB(I322537_rst), .Q(I322766) );
nor I_18650 (I322783,I322766,I322605);
not I_18651 (I322800,I322766);
nand I_18652 (I322511,I322588,I322800);
DFFARX1 I_18653  ( .D(I308940), .CLK(I5694_clk), .RSTB(I322537_rst), .Q(I322831) );
and I_18654 (I322848,I322831,I308916);
nor I_18655 (I322865,I322848,I322766);
nor I_18656 (I322882,I322848,I322800);
nand I_18657 (I322517,I322636,I322882);
not I_18658 (I322520,I322848);
DFFARX1 I_18659  ( .D(I322848), .CLK(I5694_clk), .RSTB(I322537_rst), .Q(I322499) );
DFFARX1 I_18660  ( .D(I308943), .CLK(I5694_clk), .RSTB(I322537_rst), .Q(I322941) );
nand I_18661 (I322958,I322941,I322653);
and I_18662 (I322975,I322636,I322958);
DFFARX1 I_18663  ( .D(I322975), .CLK(I5694_clk), .RSTB(I322537_rst), .Q(I322529) );
nor I_18664 (I322526,I322941,I322848);
and I_18665 (I323020,I322941,I322783);
or I_18666 (I323037,I322636,I323020);
DFFARX1 I_18667  ( .D(I323037), .CLK(I5694_clk), .RSTB(I322537_rst), .Q(I322514) );
nand I_18668 (I322523,I322941,I322865);
not I_18669 (I323115_rst,I5701);
nand I_18670 (I323132,I316870,I316867);
and I_18671 (I323149,I323132,I316879);
DFFARX1 I_18672  ( .D(I323149), .CLK(I5694_clk), .RSTB(I323115_rst), .Q(I323166) );
not I_18673 (I323183,I323166);
DFFARX1 I_18674  ( .D(I323166), .CLK(I5694_clk), .RSTB(I323115_rst), .Q(I323083) );
nor I_18675 (I323214,I316876,I316867);
DFFARX1 I_18676  ( .D(I316882), .CLK(I5694_clk), .RSTB(I323115_rst), .Q(I323231) );
DFFARX1 I_18677  ( .D(I323231), .CLK(I5694_clk), .RSTB(I323115_rst), .Q(I323248) );
not I_18678 (I323086,I323248);
DFFARX1 I_18679  ( .D(I323231), .CLK(I5694_clk), .RSTB(I323115_rst), .Q(I323279) );
and I_18680 (I323080,I323166,I323279);
nand I_18681 (I323310,I316858,I316861);
and I_18682 (I323327,I323310,I316885);
DFFARX1 I_18683  ( .D(I323327), .CLK(I5694_clk), .RSTB(I323115_rst), .Q(I323344) );
nor I_18684 (I323361,I323344,I323183);
not I_18685 (I323378,I323344);
nand I_18686 (I323089,I323166,I323378);
DFFARX1 I_18687  ( .D(I316864), .CLK(I5694_clk), .RSTB(I323115_rst), .Q(I323409) );
and I_18688 (I323426,I323409,I316855);
nor I_18689 (I323443,I323426,I323344);
nor I_18690 (I323460,I323426,I323378);
nand I_18691 (I323095,I323214,I323460);
not I_18692 (I323098,I323426);
DFFARX1 I_18693  ( .D(I323426), .CLK(I5694_clk), .RSTB(I323115_rst), .Q(I323077) );
DFFARX1 I_18694  ( .D(I316873), .CLK(I5694_clk), .RSTB(I323115_rst), .Q(I323519) );
nand I_18695 (I323536,I323519,I323231);
and I_18696 (I323553,I323214,I323536);
DFFARX1 I_18697  ( .D(I323553), .CLK(I5694_clk), .RSTB(I323115_rst), .Q(I323107) );
nor I_18698 (I323104,I323519,I323426);
and I_18699 (I323598,I323519,I323361);
or I_18700 (I323615,I323214,I323598);
DFFARX1 I_18701  ( .D(I323615), .CLK(I5694_clk), .RSTB(I323115_rst), .Q(I323092) );
nand I_18702 (I323101,I323519,I323443);
not I_18703 (I323693_rst,I5701);
nand I_18704 (I323710,I271764,I271752);
and I_18705 (I323727,I323710,I271746);
DFFARX1 I_18706  ( .D(I323727), .CLK(I5694_clk), .RSTB(I323693_rst), .Q(I323744) );
not I_18707 (I323761,I323744);
DFFARX1 I_18708  ( .D(I323744), .CLK(I5694_clk), .RSTB(I323693_rst), .Q(I323661) );
nor I_18709 (I323792,I271743,I271752);
DFFARX1 I_18710  ( .D(I271737), .CLK(I5694_clk), .RSTB(I323693_rst), .Q(I323809) );
DFFARX1 I_18711  ( .D(I323809), .CLK(I5694_clk), .RSTB(I323693_rst), .Q(I323826) );
not I_18712 (I323664,I323826);
DFFARX1 I_18713  ( .D(I323809), .CLK(I5694_clk), .RSTB(I323693_rst), .Q(I323857) );
and I_18714 (I323658,I323744,I323857);
nand I_18715 (I323888,I271740,I271755);
and I_18716 (I323905,I323888,I271767);
DFFARX1 I_18717  ( .D(I323905), .CLK(I5694_clk), .RSTB(I323693_rst), .Q(I323922) );
nor I_18718 (I323939,I323922,I323761);
not I_18719 (I323956,I323922);
nand I_18720 (I323667,I323744,I323956);
DFFARX1 I_18721  ( .D(I271758), .CLK(I5694_clk), .RSTB(I323693_rst), .Q(I323987) );
and I_18722 (I324004,I323987,I271749);
nor I_18723 (I324021,I324004,I323922);
nor I_18724 (I324038,I324004,I323956);
nand I_18725 (I323673,I323792,I324038);
not I_18726 (I323676,I324004);
DFFARX1 I_18727  ( .D(I324004), .CLK(I5694_clk), .RSTB(I323693_rst), .Q(I323655) );
DFFARX1 I_18728  ( .D(I271761), .CLK(I5694_clk), .RSTB(I323693_rst), .Q(I324097) );
nand I_18729 (I324114,I324097,I323809);
and I_18730 (I324131,I323792,I324114);
DFFARX1 I_18731  ( .D(I324131), .CLK(I5694_clk), .RSTB(I323693_rst), .Q(I323685) );
nor I_18732 (I323682,I324097,I324004);
and I_18733 (I324176,I324097,I323939);
or I_18734 (I324193,I323792,I324176);
DFFARX1 I_18735  ( .D(I324193), .CLK(I5694_clk), .RSTB(I323693_rst), .Q(I323670) );
nand I_18736 (I323679,I324097,I324021);
not I_18737 (I324271_rst,I5701);
nand I_18738 (I324288,I310245,I310272);
and I_18739 (I324305,I324288,I310260);
DFFARX1 I_18740  ( .D(I324305), .CLK(I5694_clk), .RSTB(I324271_rst), .Q(I324322) );
not I_18741 (I324339,I324322);
DFFARX1 I_18742  ( .D(I324322), .CLK(I5694_clk), .RSTB(I324271_rst), .Q(I324239) );
nor I_18743 (I324370,I310248,I310272);
DFFARX1 I_18744  ( .D(I310263), .CLK(I5694_clk), .RSTB(I324271_rst), .Q(I324387) );
DFFARX1 I_18745  ( .D(I324387), .CLK(I5694_clk), .RSTB(I324271_rst), .Q(I324404) );
not I_18746 (I324242,I324404);
DFFARX1 I_18747  ( .D(I324387), .CLK(I5694_clk), .RSTB(I324271_rst), .Q(I324435) );
and I_18748 (I324236,I324322,I324435);
nand I_18749 (I324466,I310257,I310254);
and I_18750 (I324483,I324466,I310251);
DFFARX1 I_18751  ( .D(I324483), .CLK(I5694_clk), .RSTB(I324271_rst), .Q(I324500) );
nor I_18752 (I324517,I324500,I324339);
not I_18753 (I324534,I324500);
nand I_18754 (I324245,I324322,I324534);
DFFARX1 I_18755  ( .D(I310266), .CLK(I5694_clk), .RSTB(I324271_rst), .Q(I324565) );
and I_18756 (I324582,I324565,I310242);
nor I_18757 (I324599,I324582,I324500);
nor I_18758 (I324616,I324582,I324534);
nand I_18759 (I324251,I324370,I324616);
not I_18760 (I324254,I324582);
DFFARX1 I_18761  ( .D(I324582), .CLK(I5694_clk), .RSTB(I324271_rst), .Q(I324233) );
DFFARX1 I_18762  ( .D(I310269), .CLK(I5694_clk), .RSTB(I324271_rst), .Q(I324675) );
nand I_18763 (I324692,I324675,I324387);
and I_18764 (I324709,I324370,I324692);
DFFARX1 I_18765  ( .D(I324709), .CLK(I5694_clk), .RSTB(I324271_rst), .Q(I324263) );
nor I_18766 (I324260,I324675,I324582);
and I_18767 (I324754,I324675,I324517);
or I_18768 (I324771,I324370,I324754);
DFFARX1 I_18769  ( .D(I324771), .CLK(I5694_clk), .RSTB(I324271_rst), .Q(I324248) );
nand I_18770 (I324257,I324675,I324599);
not I_18771 (I324849_rst,I5701);
nand I_18772 (I324866,I299570,I299552);
and I_18773 (I324883,I324866,I299564);
DFFARX1 I_18774  ( .D(I324883), .CLK(I5694_clk), .RSTB(I324849_rst), .Q(I324900) );
not I_18775 (I324917,I324900);
DFFARX1 I_18776  ( .D(I324900), .CLK(I5694_clk), .RSTB(I324849_rst), .Q(I324817) );
nor I_18777 (I324948,I299567,I299552);
DFFARX1 I_18778  ( .D(I299576), .CLK(I5694_clk), .RSTB(I324849_rst), .Q(I324965) );
DFFARX1 I_18779  ( .D(I324965), .CLK(I5694_clk), .RSTB(I324849_rst), .Q(I324982) );
not I_18780 (I324820,I324982);
DFFARX1 I_18781  ( .D(I324965), .CLK(I5694_clk), .RSTB(I324849_rst), .Q(I325013) );
and I_18782 (I324814,I324900,I325013);
nand I_18783 (I325044,I299555,I299579);
and I_18784 (I325061,I325044,I299558);
DFFARX1 I_18785  ( .D(I325061), .CLK(I5694_clk), .RSTB(I324849_rst), .Q(I325078) );
nor I_18786 (I325095,I325078,I324917);
not I_18787 (I325112,I325078);
nand I_18788 (I324823,I324900,I325112);
DFFARX1 I_18789  ( .D(I299561), .CLK(I5694_clk), .RSTB(I324849_rst), .Q(I325143) );
and I_18790 (I325160,I325143,I299573);
nor I_18791 (I325177,I325160,I325078);
nor I_18792 (I325194,I325160,I325112);
nand I_18793 (I324829,I324948,I325194);
not I_18794 (I324832,I325160);
DFFARX1 I_18795  ( .D(I325160), .CLK(I5694_clk), .RSTB(I324849_rst), .Q(I324811) );
DFFARX1 I_18796  ( .D(I299549), .CLK(I5694_clk), .RSTB(I324849_rst), .Q(I325253) );
nand I_18797 (I325270,I325253,I324965);
and I_18798 (I325287,I324948,I325270);
DFFARX1 I_18799  ( .D(I325287), .CLK(I5694_clk), .RSTB(I324849_rst), .Q(I324841) );
nor I_18800 (I324838,I325253,I325160);
and I_18801 (I325332,I325253,I325095);
or I_18802 (I325349,I324948,I325332);
DFFARX1 I_18803  ( .D(I325349), .CLK(I5694_clk), .RSTB(I324849_rst), .Q(I324826) );
nand I_18804 (I324835,I325253,I325177);
not I_18805 (I325427_rst,I5701);
nand I_18806 (I325444,I312897,I312924);
and I_18807 (I325461,I325444,I312912);
DFFARX1 I_18808  ( .D(I325461), .CLK(I5694_clk), .RSTB(I325427_rst), .Q(I325478) );
not I_18809 (I325495,I325478);
DFFARX1 I_18810  ( .D(I325478), .CLK(I5694_clk), .RSTB(I325427_rst), .Q(I325395) );
nor I_18811 (I325526,I312900,I312924);
DFFARX1 I_18812  ( .D(I312915), .CLK(I5694_clk), .RSTB(I325427_rst), .Q(I325543) );
DFFARX1 I_18813  ( .D(I325543), .CLK(I5694_clk), .RSTB(I325427_rst), .Q(I325560) );
not I_18814 (I325398,I325560);
DFFARX1 I_18815  ( .D(I325543), .CLK(I5694_clk), .RSTB(I325427_rst), .Q(I325591) );
and I_18816 (I325392,I325478,I325591);
nand I_18817 (I325622,I312909,I312906);
and I_18818 (I325639,I325622,I312903);
DFFARX1 I_18819  ( .D(I325639), .CLK(I5694_clk), .RSTB(I325427_rst), .Q(I325656) );
nor I_18820 (I325673,I325656,I325495);
not I_18821 (I325690,I325656);
nand I_18822 (I325401,I325478,I325690);
DFFARX1 I_18823  ( .D(I312918), .CLK(I5694_clk), .RSTB(I325427_rst), .Q(I325721) );
and I_18824 (I325738,I325721,I312894);
nor I_18825 (I325755,I325738,I325656);
nor I_18826 (I325772,I325738,I325690);
nand I_18827 (I325407,I325526,I325772);
not I_18828 (I325410,I325738);
DFFARX1 I_18829  ( .D(I325738), .CLK(I5694_clk), .RSTB(I325427_rst), .Q(I325389) );
DFFARX1 I_18830  ( .D(I312921), .CLK(I5694_clk), .RSTB(I325427_rst), .Q(I325831) );
nand I_18831 (I325848,I325831,I325543);
and I_18832 (I325865,I325526,I325848);
DFFARX1 I_18833  ( .D(I325865), .CLK(I5694_clk), .RSTB(I325427_rst), .Q(I325419) );
nor I_18834 (I325416,I325831,I325738);
and I_18835 (I325910,I325831,I325673);
or I_18836 (I325927,I325526,I325910);
DFFARX1 I_18837  ( .D(I325927), .CLK(I5694_clk), .RSTB(I325427_rst), .Q(I325404) );
nand I_18838 (I325413,I325831,I325755);
not I_18839 (I326005_rst,I5701);
nand I_18840 (I326022,I277702,I277693);
and I_18841 (I326039,I326022,I277711);
DFFARX1 I_18842  ( .D(I326039), .CLK(I5694_clk), .RSTB(I326005_rst), .Q(I326056) );
nor I_18843 (I326073,I277690,I277693);
nor I_18844 (I326090,I326073,I326056);
not I_18845 (I325988,I326073);
DFFARX1 I_18846  ( .D(I277699), .CLK(I5694_clk), .RSTB(I326005_rst), .Q(I326121) );
not I_18847 (I326138,I326121);
nor I_18848 (I326155,I326073,I326138);
nand I_18849 (I325991,I326121,I326090);
DFFARX1 I_18850  ( .D(I326121), .CLK(I5694_clk), .RSTB(I326005_rst), .Q(I325973) );
nand I_18851 (I326200,I277714,I277696);
and I_18852 (I326217,I326200,I277717);
DFFARX1 I_18853  ( .D(I326217), .CLK(I5694_clk), .RSTB(I326005_rst), .Q(I326234) );
nor I_18854 (I325994,I326234,I326056);
nand I_18855 (I325985,I326234,I326155);
DFFARX1 I_18856  ( .D(I277705), .CLK(I5694_clk), .RSTB(I326005_rst), .Q(I326279) );
and I_18857 (I326296,I326279,I277687);
DFFARX1 I_18858  ( .D(I326296), .CLK(I5694_clk), .RSTB(I326005_rst), .Q(I326313) );
not I_18859 (I325976,I326313);
nand I_18860 (I326344,I326296,I326234);
and I_18861 (I326361,I326056,I326344);
DFFARX1 I_18862  ( .D(I326361), .CLK(I5694_clk), .RSTB(I326005_rst), .Q(I325967) );
DFFARX1 I_18863  ( .D(I277708), .CLK(I5694_clk), .RSTB(I326005_rst), .Q(I326392) );
nand I_18864 (I326409,I326392,I326056);
and I_18865 (I326426,I326234,I326409);
DFFARX1 I_18866  ( .D(I326426), .CLK(I5694_clk), .RSTB(I326005_rst), .Q(I325997) );
not I_18867 (I326457,I326392);
nor I_18868 (I326474,I326073,I326457);
and I_18869 (I326491,I326392,I326474);
or I_18870 (I326508,I326296,I326491);
DFFARX1 I_18871  ( .D(I326508), .CLK(I5694_clk), .RSTB(I326005_rst), .Q(I325982) );
nand I_18872 (I325979,I326392,I326138);
DFFARX1 I_18873  ( .D(I326392), .CLK(I5694_clk), .RSTB(I326005_rst), .Q(I325970) );
not I_18874 (I326600_rst,I5701);
nand I_18875 (I326617,I280153,I280144);
and I_18876 (I326634,I326617,I280162);
DFFARX1 I_18877  ( .D(I326634), .CLK(I5694_clk), .RSTB(I326600_rst), .Q(I326651) );
nor I_18878 (I326668,I280159,I280144);
nor I_18879 (I326685,I326668,I326651);
not I_18880 (I326583,I326668);
DFFARX1 I_18881  ( .D(I280141), .CLK(I5694_clk), .RSTB(I326600_rst), .Q(I326716) );
not I_18882 (I326733,I326716);
nor I_18883 (I326750,I326668,I326733);
nand I_18884 (I326586,I326716,I326685);
DFFARX1 I_18885  ( .D(I326716), .CLK(I5694_clk), .RSTB(I326600_rst), .Q(I326568) );
nand I_18886 (I326795,I280150,I280165);
and I_18887 (I326812,I326795,I280156);
DFFARX1 I_18888  ( .D(I326812), .CLK(I5694_clk), .RSTB(I326600_rst), .Q(I326829) );
nor I_18889 (I326589,I326829,I326651);
nand I_18890 (I326580,I326829,I326750);
DFFARX1 I_18891  ( .D(I280138), .CLK(I5694_clk), .RSTB(I326600_rst), .Q(I326874) );
and I_18892 (I326891,I326874,I280147);
DFFARX1 I_18893  ( .D(I326891), .CLK(I5694_clk), .RSTB(I326600_rst), .Q(I326908) );
not I_18894 (I326571,I326908);
nand I_18895 (I326939,I326891,I326829);
and I_18896 (I326956,I326651,I326939);
DFFARX1 I_18897  ( .D(I326956), .CLK(I5694_clk), .RSTB(I326600_rst), .Q(I326562) );
DFFARX1 I_18898  ( .D(I280135), .CLK(I5694_clk), .RSTB(I326600_rst), .Q(I326987) );
nand I_18899 (I327004,I326987,I326651);
and I_18900 (I327021,I326829,I327004);
DFFARX1 I_18901  ( .D(I327021), .CLK(I5694_clk), .RSTB(I326600_rst), .Q(I326592) );
not I_18902 (I327052,I326987);
nor I_18903 (I327069,I326668,I327052);
and I_18904 (I327086,I326987,I327069);
or I_18905 (I327103,I326891,I327086);
DFFARX1 I_18906  ( .D(I327103), .CLK(I5694_clk), .RSTB(I326600_rst), .Q(I326577) );
nand I_18907 (I326574,I326987,I326733);
DFFARX1 I_18908  ( .D(I326987), .CLK(I5694_clk), .RSTB(I326600_rst), .Q(I326565) );
not I_18909 (I327195_rst,I5701);
nand I_18910 (I327212,I276512,I276503);
and I_18911 (I327229,I327212,I276521);
DFFARX1 I_18912  ( .D(I327229), .CLK(I5694_clk), .RSTB(I327195_rst), .Q(I327246) );
nor I_18913 (I327263,I276500,I276503);
nor I_18914 (I327280,I327263,I327246);
not I_18915 (I327178,I327263);
DFFARX1 I_18916  ( .D(I276509), .CLK(I5694_clk), .RSTB(I327195_rst), .Q(I327311) );
not I_18917 (I327328,I327311);
nor I_18918 (I327345,I327263,I327328);
nand I_18919 (I327181,I327311,I327280);
DFFARX1 I_18920  ( .D(I327311), .CLK(I5694_clk), .RSTB(I327195_rst), .Q(I327163) );
nand I_18921 (I327390,I276524,I276506);
and I_18922 (I327407,I327390,I276527);
DFFARX1 I_18923  ( .D(I327407), .CLK(I5694_clk), .RSTB(I327195_rst), .Q(I327424) );
nor I_18924 (I327184,I327424,I327246);
nand I_18925 (I327175,I327424,I327345);
DFFARX1 I_18926  ( .D(I276515), .CLK(I5694_clk), .RSTB(I327195_rst), .Q(I327469) );
and I_18927 (I327486,I327469,I276497);
DFFARX1 I_18928  ( .D(I327486), .CLK(I5694_clk), .RSTB(I327195_rst), .Q(I327503) );
not I_18929 (I327166,I327503);
nand I_18930 (I327534,I327486,I327424);
and I_18931 (I327551,I327246,I327534);
DFFARX1 I_18932  ( .D(I327551), .CLK(I5694_clk), .RSTB(I327195_rst), .Q(I327157) );
DFFARX1 I_18933  ( .D(I276518), .CLK(I5694_clk), .RSTB(I327195_rst), .Q(I327582) );
nand I_18934 (I327599,I327582,I327246);
and I_18935 (I327616,I327424,I327599);
DFFARX1 I_18936  ( .D(I327616), .CLK(I5694_clk), .RSTB(I327195_rst), .Q(I327187) );
not I_18937 (I327647,I327582);
nor I_18938 (I327664,I327263,I327647);
and I_18939 (I327681,I327582,I327664);
or I_18940 (I327698,I327486,I327681);
DFFARX1 I_18941  ( .D(I327698), .CLK(I5694_clk), .RSTB(I327195_rst), .Q(I327172) );
nand I_18942 (I327169,I327582,I327328);
DFFARX1 I_18943  ( .D(I327582), .CLK(I5694_clk), .RSTB(I327195_rst), .Q(I327160) );
not I_18944 (I327790_rst,I5701);
nand I_18945 (I327807,I296328,I296340);
and I_18946 (I327824,I327807,I296349);
DFFARX1 I_18947  ( .D(I327824), .CLK(I5694_clk), .RSTB(I327790_rst), .Q(I327841) );
nor I_18948 (I327858,I296343,I296340);
nor I_18949 (I327875,I327858,I327841);
not I_18950 (I327773,I327858);
DFFARX1 I_18951  ( .D(I296337), .CLK(I5694_clk), .RSTB(I327790_rst), .Q(I327906) );
not I_18952 (I327923,I327906);
nor I_18953 (I327940,I327858,I327923);
nand I_18954 (I327776,I327906,I327875);
DFFARX1 I_18955  ( .D(I327906), .CLK(I5694_clk), .RSTB(I327790_rst), .Q(I327758) );
nand I_18956 (I327985,I296334,I296331);
and I_18957 (I328002,I327985,I296322);
DFFARX1 I_18958  ( .D(I328002), .CLK(I5694_clk), .RSTB(I327790_rst), .Q(I328019) );
nor I_18959 (I327779,I328019,I327841);
nand I_18960 (I327770,I328019,I327940);
DFFARX1 I_18961  ( .D(I296346), .CLK(I5694_clk), .RSTB(I327790_rst), .Q(I328064) );
and I_18962 (I328081,I328064,I296325);
DFFARX1 I_18963  ( .D(I328081), .CLK(I5694_clk), .RSTB(I327790_rst), .Q(I328098) );
not I_18964 (I327761,I328098);
nand I_18965 (I328129,I328081,I328019);
and I_18966 (I328146,I327841,I328129);
DFFARX1 I_18967  ( .D(I328146), .CLK(I5694_clk), .RSTB(I327790_rst), .Q(I327752) );
DFFARX1 I_18968  ( .D(I296319), .CLK(I5694_clk), .RSTB(I327790_rst), .Q(I328177) );
nand I_18969 (I328194,I328177,I327841);
and I_18970 (I328211,I328019,I328194);
DFFARX1 I_18971  ( .D(I328211), .CLK(I5694_clk), .RSTB(I327790_rst), .Q(I327782) );
not I_18972 (I328242,I328177);
nor I_18973 (I328259,I327858,I328242);
and I_18974 (I328276,I328177,I328259);
or I_18975 (I328293,I328081,I328276);
DFFARX1 I_18976  ( .D(I328293), .CLK(I5694_clk), .RSTB(I327790_rst), .Q(I327767) );
nand I_18977 (I327764,I328177,I327923);
DFFARX1 I_18978  ( .D(I328177), .CLK(I5694_clk), .RSTB(I327790_rst), .Q(I327755) );
not I_18979 (I328385_rst,I5701);
nand I_18980 (I328402,I324260,I324263);
and I_18981 (I328419,I328402,I324257);
DFFARX1 I_18982  ( .D(I328419), .CLK(I5694_clk), .RSTB(I328385_rst), .Q(I328436) );
nor I_18983 (I328453,I324254,I324263);
nor I_18984 (I328470,I328453,I328436);
not I_18985 (I328368,I328453);
DFFARX1 I_18986  ( .D(I324236), .CLK(I5694_clk), .RSTB(I328385_rst), .Q(I328501) );
not I_18987 (I328518,I328501);
nor I_18988 (I328535,I328453,I328518);
nand I_18989 (I328371,I328501,I328470);
DFFARX1 I_18990  ( .D(I328501), .CLK(I5694_clk), .RSTB(I328385_rst), .Q(I328353) );
nand I_18991 (I328580,I324245,I324242);
and I_18992 (I328597,I328580,I324251);
DFFARX1 I_18993  ( .D(I328597), .CLK(I5694_clk), .RSTB(I328385_rst), .Q(I328614) );
nor I_18994 (I328374,I328614,I328436);
nand I_18995 (I328365,I328614,I328535);
DFFARX1 I_18996  ( .D(I324233), .CLK(I5694_clk), .RSTB(I328385_rst), .Q(I328659) );
and I_18997 (I328676,I328659,I324248);
DFFARX1 I_18998  ( .D(I328676), .CLK(I5694_clk), .RSTB(I328385_rst), .Q(I328693) );
not I_18999 (I328356,I328693);
nand I_19000 (I328724,I328676,I328614);
and I_19001 (I328741,I328436,I328724);
DFFARX1 I_19002  ( .D(I328741), .CLK(I5694_clk), .RSTB(I328385_rst), .Q(I328347) );
DFFARX1 I_19003  ( .D(I324239), .CLK(I5694_clk), .RSTB(I328385_rst), .Q(I328772) );
nand I_19004 (I328789,I328772,I328436);
and I_19005 (I328806,I328614,I328789);
DFFARX1 I_19006  ( .D(I328806), .CLK(I5694_clk), .RSTB(I328385_rst), .Q(I328377) );
not I_19007 (I328837,I328772);
nor I_19008 (I328854,I328453,I328837);
and I_19009 (I328871,I328772,I328854);
or I_19010 (I328888,I328676,I328871);
DFFARX1 I_19011  ( .D(I328888), .CLK(I5694_clk), .RSTB(I328385_rst), .Q(I328362) );
nand I_19012 (I328359,I328772,I328518);
DFFARX1 I_19013  ( .D(I328772), .CLK(I5694_clk), .RSTB(I328385_rst), .Q(I328350) );
not I_19014 (I328980_rst,I5701);
nand I_19015 (I328997,I292616,I292622);
and I_19016 (I329014,I328997,I292619);
DFFARX1 I_19017  ( .D(I329014), .CLK(I5694_clk), .RSTB(I328980_rst), .Q(I329031) );
nor I_19018 (I329048,I292643,I292622);
nor I_19019 (I329065,I329048,I329031);
not I_19020 (I328963,I329048);
DFFARX1 I_19021  ( .D(I292634), .CLK(I5694_clk), .RSTB(I328980_rst), .Q(I329096) );
not I_19022 (I329113,I329096);
nor I_19023 (I329130,I329048,I329113);
nand I_19024 (I328966,I329096,I329065);
DFFARX1 I_19025  ( .D(I329096), .CLK(I5694_clk), .RSTB(I328980_rst), .Q(I328948) );
nand I_19026 (I329175,I292637,I292640);
and I_19027 (I329192,I329175,I292613);
DFFARX1 I_19028  ( .D(I329192), .CLK(I5694_clk), .RSTB(I328980_rst), .Q(I329209) );
nor I_19029 (I328969,I329209,I329031);
nand I_19030 (I328960,I329209,I329130);
DFFARX1 I_19031  ( .D(I292631), .CLK(I5694_clk), .RSTB(I328980_rst), .Q(I329254) );
and I_19032 (I329271,I329254,I292625);
DFFARX1 I_19033  ( .D(I329271), .CLK(I5694_clk), .RSTB(I328980_rst), .Q(I329288) );
not I_19034 (I328951,I329288);
nand I_19035 (I329319,I329271,I329209);
and I_19036 (I329336,I329031,I329319);
DFFARX1 I_19037  ( .D(I329336), .CLK(I5694_clk), .RSTB(I328980_rst), .Q(I328942) );
DFFARX1 I_19038  ( .D(I292628), .CLK(I5694_clk), .RSTB(I328980_rst), .Q(I329367) );
nand I_19039 (I329384,I329367,I329031);
and I_19040 (I329401,I329209,I329384);
DFFARX1 I_19041  ( .D(I329401), .CLK(I5694_clk), .RSTB(I328980_rst), .Q(I328972) );
not I_19042 (I329432,I329367);
nor I_19043 (I329449,I329048,I329432);
and I_19044 (I329466,I329367,I329449);
or I_19045 (I329483,I329271,I329466);
DFFARX1 I_19046  ( .D(I329483), .CLK(I5694_clk), .RSTB(I328980_rst), .Q(I328957) );
nand I_19047 (I328954,I329367,I329113);
DFFARX1 I_19048  ( .D(I329367), .CLK(I5694_clk), .RSTB(I328980_rst), .Q(I328945) );
not I_19049 (I329575_rst,I5701);
nand I_19050 (I329592,I281411,I281402);
and I_19051 (I329609,I329592,I281420);
DFFARX1 I_19052  ( .D(I329609), .CLK(I5694_clk), .RSTB(I329575_rst), .Q(I329626) );
nor I_19053 (I329643,I281417,I281402);
nor I_19054 (I329660,I329643,I329626);
not I_19055 (I329558,I329643);
DFFARX1 I_19056  ( .D(I281399), .CLK(I5694_clk), .RSTB(I329575_rst), .Q(I329691) );
not I_19057 (I329708,I329691);
nor I_19058 (I329725,I329643,I329708);
nand I_19059 (I329561,I329691,I329660);
DFFARX1 I_19060  ( .D(I329691), .CLK(I5694_clk), .RSTB(I329575_rst), .Q(I329543) );
nand I_19061 (I329770,I281408,I281423);
and I_19062 (I329787,I329770,I281414);
DFFARX1 I_19063  ( .D(I329787), .CLK(I5694_clk), .RSTB(I329575_rst), .Q(I329804) );
nor I_19064 (I329564,I329804,I329626);
nand I_19065 (I329555,I329804,I329725);
DFFARX1 I_19066  ( .D(I281396), .CLK(I5694_clk), .RSTB(I329575_rst), .Q(I329849) );
and I_19067 (I329866,I329849,I281405);
DFFARX1 I_19068  ( .D(I329866), .CLK(I5694_clk), .RSTB(I329575_rst), .Q(I329883) );
not I_19069 (I329546,I329883);
nand I_19070 (I329914,I329866,I329804);
and I_19071 (I329931,I329626,I329914);
DFFARX1 I_19072  ( .D(I329931), .CLK(I5694_clk), .RSTB(I329575_rst), .Q(I329537) );
DFFARX1 I_19073  ( .D(I281393), .CLK(I5694_clk), .RSTB(I329575_rst), .Q(I329962) );
nand I_19074 (I329979,I329962,I329626);
and I_19075 (I329996,I329804,I329979);
DFFARX1 I_19076  ( .D(I329996), .CLK(I5694_clk), .RSTB(I329575_rst), .Q(I329567) );
not I_19077 (I330027,I329962);
nor I_19078 (I330044,I329643,I330027);
and I_19079 (I330061,I329962,I330044);
or I_19080 (I330078,I329866,I330061);
DFFARX1 I_19081  ( .D(I330078), .CLK(I5694_clk), .RSTB(I329575_rst), .Q(I329552) );
nand I_19082 (I329549,I329962,I329708);
DFFARX1 I_19083  ( .D(I329962), .CLK(I5694_clk), .RSTB(I329575_rst), .Q(I329540) );
not I_19084 (I330170_rst,I5701);
nand I_19085 (I330187,I300204,I300216);
and I_19086 (I330204,I330187,I300225);
DFFARX1 I_19087  ( .D(I330204), .CLK(I5694_clk), .RSTB(I330170_rst), .Q(I330221) );
nor I_19088 (I330238,I300219,I300216);
nor I_19089 (I330255,I330238,I330221);
not I_19090 (I330153,I330238);
DFFARX1 I_19091  ( .D(I300213), .CLK(I5694_clk), .RSTB(I330170_rst), .Q(I330286) );
not I_19092 (I330303,I330286);
nor I_19093 (I330320,I330238,I330303);
nand I_19094 (I330156,I330286,I330255);
DFFARX1 I_19095  ( .D(I330286), .CLK(I5694_clk), .RSTB(I330170_rst), .Q(I330138) );
nand I_19096 (I330365,I300210,I300207);
and I_19097 (I330382,I330365,I300198);
DFFARX1 I_19098  ( .D(I330382), .CLK(I5694_clk), .RSTB(I330170_rst), .Q(I330399) );
nor I_19099 (I330159,I330399,I330221);
nand I_19100 (I330150,I330399,I330320);
DFFARX1 I_19101  ( .D(I300222), .CLK(I5694_clk), .RSTB(I330170_rst), .Q(I330444) );
and I_19102 (I330461,I330444,I300201);
DFFARX1 I_19103  ( .D(I330461), .CLK(I5694_clk), .RSTB(I330170_rst), .Q(I330478) );
not I_19104 (I330141,I330478);
nand I_19105 (I330509,I330461,I330399);
and I_19106 (I330526,I330221,I330509);
DFFARX1 I_19107  ( .D(I330526), .CLK(I5694_clk), .RSTB(I330170_rst), .Q(I330132) );
DFFARX1 I_19108  ( .D(I300195), .CLK(I5694_clk), .RSTB(I330170_rst), .Q(I330557) );
nand I_19109 (I330574,I330557,I330221);
and I_19110 (I330591,I330399,I330574);
DFFARX1 I_19111  ( .D(I330591), .CLK(I5694_clk), .RSTB(I330170_rst), .Q(I330162) );
not I_19112 (I330622,I330557);
nor I_19113 (I330639,I330238,I330622);
and I_19114 (I330656,I330557,I330639);
or I_19115 (I330673,I330461,I330656);
DFFARX1 I_19116  ( .D(I330673), .CLK(I5694_clk), .RSTB(I330170_rst), .Q(I330147) );
nand I_19117 (I330144,I330557,I330303);
DFFARX1 I_19118  ( .D(I330557), .CLK(I5694_clk), .RSTB(I330170_rst), .Q(I330135) );
not I_19119 (I330765_rst,I5701);
nand I_19120 (I330782,I283310,I283298);
and I_19121 (I330799,I330782,I283283);
DFFARX1 I_19122  ( .D(I330799), .CLK(I5694_clk), .RSTB(I330765_rst), .Q(I330816) );
nor I_19123 (I330833,I283295,I283298);
DFFARX1 I_19124  ( .D(I283307), .CLK(I5694_clk), .RSTB(I330765_rst), .Q(I330850) );
nand I_19125 (I330867,I330850,I330833);
DFFARX1 I_19126  ( .D(I330850), .CLK(I5694_clk), .RSTB(I330765_rst), .Q(I330736) );
nand I_19127 (I330898,I283280,I283304);
and I_19128 (I330915,I330898,I283289);
DFFARX1 I_19129  ( .D(I330915), .CLK(I5694_clk), .RSTB(I330765_rst), .Q(I330932) );
not I_19130 (I330949,I330932);
nor I_19131 (I330966,I330816,I330949);
and I_19132 (I330983,I330833,I330966);
and I_19133 (I331000,I330932,I330867);
DFFARX1 I_19134  ( .D(I331000), .CLK(I5694_clk), .RSTB(I330765_rst), .Q(I330733) );
DFFARX1 I_19135  ( .D(I330932), .CLK(I5694_clk), .RSTB(I330765_rst), .Q(I330727) );
DFFARX1 I_19136  ( .D(I283292), .CLK(I5694_clk), .RSTB(I330765_rst), .Q(I331045) );
and I_19137 (I331062,I331045,I283301);
nand I_19138 (I331079,I331062,I330932);
nor I_19139 (I330754,I331062,I330833);
not I_19140 (I331110,I331062);
nor I_19141 (I331127,I330816,I331110);
nand I_19142 (I330745,I330850,I331127);
nand I_19143 (I330739,I330932,I331110);
or I_19144 (I331172,I331062,I330983);
DFFARX1 I_19145  ( .D(I331172), .CLK(I5694_clk), .RSTB(I330765_rst), .Q(I330742) );
DFFARX1 I_19146  ( .D(I283286), .CLK(I5694_clk), .RSTB(I330765_rst), .Q(I331203) );
and I_19147 (I331220,I331203,I331079);
DFFARX1 I_19148  ( .D(I331220), .CLK(I5694_clk), .RSTB(I330765_rst), .Q(I330757) );
nor I_19149 (I331251,I331203,I330816);
nand I_19150 (I330751,I331062,I331251);
not I_19151 (I330748,I331203);
DFFARX1 I_19152  ( .D(I331203), .CLK(I5694_clk), .RSTB(I330765_rst), .Q(I331296) );
and I_19153 (I330730,I331203,I331296);
not I_19154 (I331360_rst,I5701);
nand I_19155 (I331377,I321355,I321370);
and I_19156 (I331394,I331377,I321367);
DFFARX1 I_19157  ( .D(I331394), .CLK(I5694_clk), .RSTB(I331360_rst), .Q(I331411) );
nor I_19158 (I331428,I321343,I321370);
DFFARX1 I_19159  ( .D(I321361), .CLK(I5694_clk), .RSTB(I331360_rst), .Q(I331445) );
nand I_19160 (I331462,I331445,I331428);
DFFARX1 I_19161  ( .D(I331445), .CLK(I5694_clk), .RSTB(I331360_rst), .Q(I331331) );
nand I_19162 (I331493,I321364,I321352);
and I_19163 (I331510,I331493,I321358);
DFFARX1 I_19164  ( .D(I331510), .CLK(I5694_clk), .RSTB(I331360_rst), .Q(I331527) );
not I_19165 (I331544,I331527);
nor I_19166 (I331561,I331411,I331544);
and I_19167 (I331578,I331428,I331561);
and I_19168 (I331595,I331527,I331462);
DFFARX1 I_19169  ( .D(I331595), .CLK(I5694_clk), .RSTB(I331360_rst), .Q(I331328) );
DFFARX1 I_19170  ( .D(I331527), .CLK(I5694_clk), .RSTB(I331360_rst), .Q(I331322) );
DFFARX1 I_19171  ( .D(I321349), .CLK(I5694_clk), .RSTB(I331360_rst), .Q(I331640) );
and I_19172 (I331657,I331640,I321373);
nand I_19173 (I331674,I331657,I331527);
nor I_19174 (I331349,I331657,I331428);
not I_19175 (I331705,I331657);
nor I_19176 (I331722,I331411,I331705);
nand I_19177 (I331340,I331445,I331722);
nand I_19178 (I331334,I331527,I331705);
or I_19179 (I331767,I331657,I331578);
DFFARX1 I_19180  ( .D(I331767), .CLK(I5694_clk), .RSTB(I331360_rst), .Q(I331337) );
DFFARX1 I_19181  ( .D(I321346), .CLK(I5694_clk), .RSTB(I331360_rst), .Q(I331798) );
and I_19182 (I331815,I331798,I331674);
DFFARX1 I_19183  ( .D(I331815), .CLK(I5694_clk), .RSTB(I331360_rst), .Q(I331352) );
nor I_19184 (I331846,I331798,I331411);
nand I_19185 (I331346,I331657,I331846);
not I_19186 (I331343,I331798);
DFFARX1 I_19187  ( .D(I331798), .CLK(I5694_clk), .RSTB(I331360_rst), .Q(I331891) );
and I_19188 (I331325,I331798,I331891);
not I_19189 (I331955_rst,I5701);
nand I_19190 (I331972,I288108,I288111);
and I_19191 (I331989,I331972,I288120);
DFFARX1 I_19192  ( .D(I331989), .CLK(I5694_clk), .RSTB(I331955_rst), .Q(I332006) );
nor I_19193 (I332023,I288114,I288111);
DFFARX1 I_19194  ( .D(I288135), .CLK(I5694_clk), .RSTB(I331955_rst), .Q(I332040) );
nand I_19195 (I332057,I332040,I332023);
DFFARX1 I_19196  ( .D(I332040), .CLK(I5694_clk), .RSTB(I331955_rst), .Q(I331926) );
nand I_19197 (I332088,I288132,I288138);
and I_19198 (I332105,I332088,I288123);
DFFARX1 I_19199  ( .D(I332105), .CLK(I5694_clk), .RSTB(I331955_rst), .Q(I332122) );
not I_19200 (I332139,I332122);
nor I_19201 (I332156,I332006,I332139);
and I_19202 (I332173,I332023,I332156);
and I_19203 (I332190,I332122,I332057);
DFFARX1 I_19204  ( .D(I332190), .CLK(I5694_clk), .RSTB(I331955_rst), .Q(I331923) );
DFFARX1 I_19205  ( .D(I332122), .CLK(I5694_clk), .RSTB(I331955_rst), .Q(I331917) );
DFFARX1 I_19206  ( .D(I288126), .CLK(I5694_clk), .RSTB(I331955_rst), .Q(I332235) );
and I_19207 (I332252,I332235,I288129);
nand I_19208 (I332269,I332252,I332122);
nor I_19209 (I331944,I332252,I332023);
not I_19210 (I332300,I332252);
nor I_19211 (I332317,I332006,I332300);
nand I_19212 (I331935,I332040,I332317);
nand I_19213 (I331929,I332122,I332300);
or I_19214 (I332362,I332252,I332173);
DFFARX1 I_19215  ( .D(I332362), .CLK(I5694_clk), .RSTB(I331955_rst), .Q(I331932) );
DFFARX1 I_19216  ( .D(I288117), .CLK(I5694_clk), .RSTB(I331955_rst), .Q(I332393) );
and I_19217 (I332410,I332393,I332269);
DFFARX1 I_19218  ( .D(I332410), .CLK(I5694_clk), .RSTB(I331955_rst), .Q(I331947) );
nor I_19219 (I332441,I332393,I332006);
nand I_19220 (I331941,I332252,I332441);
not I_19221 (I331938,I332393);
DFFARX1 I_19222  ( .D(I332393), .CLK(I5694_clk), .RSTB(I331955_rst), .Q(I33248_rst6) );
and I_19223 (I331920,I332393,I33248_rst6);
not I_19224 (I332550_rst,I5701);
not I_19225 (I332567,I295679);
nor I_19226 (I332584,I295697,I295676);
nand I_19227 (I332601,I332584,I295694);
nor I_19228 (I332618,I332567,I295697);
nand I_19229 (I332635,I332618,I295688);
not I_19230 (I332652,I295697);
not I_19231 (I332669,I332652);
not I_19232 (I332686,I295691);
nor I_19233 (I332703,I332686,I295685);
and I_19234 (I332720,I332703,I295682);
or I_19235 (I332737,I332720,I295673);
DFFARX1 I_19236  ( .D(I332737), .CLK(I5694_clk), .RSTB(I332550_rst), .Q(I332754) );
nand I_19237 (I332771,I332567,I295691);
or I_19238 (I332539,I332771,I332754);
not I_19239 (I332802,I332771);
nor I_19240 (I332819,I332754,I332802);
and I_19241 (I332836,I332652,I332819);
nand I_19242 (I332512,I332771,I332669);
DFFARX1 I_19243  ( .D(I295703), .CLK(I5694_clk), .RSTB(I332550_rst), .Q(I332867) );
or I_19244 (I332533,I332867,I332754);
nor I_19245 (I332898,I332867,I332635);
nor I_19246 (I332915,I332867,I332669);
nand I_19247 (I332518,I332601,I332915);
or I_19248 (I332946,I332867,I332836);
DFFARX1 I_19249  ( .D(I332946), .CLK(I5694_clk), .RSTB(I332550_rst), .Q(I332515) );
not I_19250 (I332521,I332867);
DFFARX1 I_19251  ( .D(I295700), .CLK(I5694_clk), .RSTB(I332550_rst), .Q(I332991) );
not I_19252 (I333008,I332991);
nor I_19253 (I333025,I333008,I332601);
DFFARX1 I_19254  ( .D(I333025), .CLK(I5694_clk), .RSTB(I332550_rst), .Q(I332527) );
nor I_19255 (I332542,I332867,I333008);
nor I_19256 (I332530,I333008,I332771);
not I_19257 (I333084,I333008);
and I_19258 (I333101,I332635,I333084);
nor I_19259 (I332536,I332771,I333101);
nand I_19260 (I332524,I333008,I332898);
not I_19261 (I333179_rst,I5701);
not I_19262 (I333196,I314238);
nor I_19263 (I333213,I314244,I314223);
nand I_19264 (I333230,I333213,I314229);
nor I_19265 (I333247,I333196,I314244);
nand I_19266 (I333264,I333247,I314235);
not I_19267 (I333281,I314244);
not I_19268 (I333298,I333281);
not I_19269 (I333315,I314232);
nor I_19270 (I333332,I333315,I314250);
and I_19271 (I333349,I333332,I314241);
or I_19272 (I333366,I333349,I314220);
DFFARX1 I_19273  ( .D(I333366), .CLK(I5694_clk), .RSTB(I333179_rst), .Q(I333383) );
nand I_19274 (I333400,I333196,I314232);
or I_19275 (I333168,I333400,I333383);
not I_19276 (I333431,I333400);
nor I_19277 (I333448,I333383,I333431);
and I_19278 (I333465,I333281,I333448);
nand I_19279 (I333141,I333400,I333298);
DFFARX1 I_19280  ( .D(I314247), .CLK(I5694_clk), .RSTB(I333179_rst), .Q(I333496) );
or I_19281 (I333162,I333496,I333383);
nor I_19282 (I333527,I333496,I333264);
nor I_19283 (I333544,I333496,I333298);
nand I_19284 (I333147,I333230,I333544);
or I_19285 (I333575,I333496,I333465);
DFFARX1 I_19286  ( .D(I333575), .CLK(I5694_clk), .RSTB(I333179_rst), .Q(I333144) );
not I_19287 (I333150,I333496);
DFFARX1 I_19288  ( .D(I314226), .CLK(I5694_clk), .RSTB(I333179_rst), .Q(I333620) );
not I_19289 (I333637,I333620);
nor I_19290 (I333654,I333637,I333230);
DFFARX1 I_19291  ( .D(I333654), .CLK(I5694_clk), .RSTB(I333179_rst), .Q(I333156) );
nor I_19292 (I333171,I333496,I333637);
nor I_19293 (I333159,I333637,I333400);
not I_19294 (I333713,I333637);
and I_19295 (I333730,I333264,I333713);
nor I_19296 (I333165,I333400,I333730);
nand I_19297 (I333153,I333637,I333527);
not I_19298 (I333808_rst,I5701);
not I_19299 (I333825,I311586);
nor I_19300 (I333842,I311592,I311571);
nand I_19301 (I333859,I333842,I311577);
nor I_19302 (I333876,I333825,I311592);
nand I_19303 (I333893,I333876,I311583);
not I_19304 (I333910,I311592);
not I_19305 (I333927,I333910);
not I_19306 (I333944,I311580);
nor I_19307 (I333961,I333944,I311598);
and I_19308 (I333978,I333961,I311589);
or I_19309 (I333995,I333978,I311568);
DFFARX1 I_19310  ( .D(I333995), .CLK(I5694_clk), .RSTB(I333808_rst), .Q(I334012) );
nand I_19311 (I334029,I333825,I311580);
or I_19312 (I333797,I334029,I334012);
not I_19313 (I334060,I334029);
nor I_19314 (I334077,I334012,I334060);
and I_19315 (I334094,I333910,I334077);
nand I_19316 (I333770,I334029,I333927);
DFFARX1 I_19317  ( .D(I311595), .CLK(I5694_clk), .RSTB(I333808_rst), .Q(I334125) );
or I_19318 (I333791,I334125,I334012);
nor I_19319 (I334156,I334125,I333893);
nor I_19320 (I334173,I334125,I333927);
nand I_19321 (I333776,I333859,I334173);
or I_19322 (I334204,I334125,I334094);
DFFARX1 I_19323  ( .D(I334204), .CLK(I5694_clk), .RSTB(I333808_rst), .Q(I333773) );
not I_19324 (I333779,I334125);
DFFARX1 I_19325  ( .D(I311574), .CLK(I5694_clk), .RSTB(I333808_rst), .Q(I334249) );
not I_19326 (I334266,I334249);
nor I_19327 (I334283,I334266,I333859);
DFFARX1 I_19328  ( .D(I334283), .CLK(I5694_clk), .RSTB(I333808_rst), .Q(I333785) );
nor I_19329 (I333800,I334125,I334266);
nor I_19330 (I333788,I334266,I334029);
not I_19331 (I334342,I334266);
and I_19332 (I334359,I333893,I334342);
nor I_19333 (I333794,I334029,I334359);
nand I_19334 (I333782,I334266,I334156);
not I_19335 (I334437_rst,I5701);
not I_19336 (I334454,I297617);
nor I_19337 (I334471,I297635,I297614);
nand I_19338 (I334488,I334471,I297632);
nor I_19339 (I334505,I334454,I297635);
nand I_19340 (I334522,I334505,I297626);
not I_19341 (I334539,I297635);
not I_19342 (I334556,I334539);
not I_19343 (I334573,I297629);
nor I_19344 (I334590,I334573,I297623);
and I_19345 (I334607,I334590,I297620);
or I_19346 (I334624,I334607,I297611);
DFFARX1 I_19347  ( .D(I334624), .CLK(I5694_clk), .RSTB(I334437_rst), .Q(I334641) );
nand I_19348 (I334658,I334454,I297629);
or I_19349 (I334426,I334658,I334641);
not I_19350 (I334689,I334658);
nor I_19351 (I334706,I334641,I334689);
and I_19352 (I334723,I334539,I334706);
nand I_19353 (I334399,I334658,I334556);
DFFARX1 I_19354  ( .D(I297641), .CLK(I5694_clk), .RSTB(I334437_rst), .Q(I334754) );
or I_19355 (I334420,I334754,I334641);
nor I_19356 (I334785,I334754,I334522);
nor I_19357 (I334802,I334754,I334556);
nand I_19358 (I334405,I334488,I334802);
or I_19359 (I334833,I334754,I334723);
DFFARX1 I_19360  ( .D(I334833), .CLK(I5694_clk), .RSTB(I334437_rst), .Q(I334402) );
not I_19361 (I334408,I334754);
DFFARX1 I_19362  ( .D(I297638), .CLK(I5694_clk), .RSTB(I334437_rst), .Q(I334878) );
not I_19363 (I334895,I334878);
nor I_19364 (I334912,I334895,I334488);
DFFARX1 I_19365  ( .D(I334912), .CLK(I5694_clk), .RSTB(I334437_rst), .Q(I334414) );
nor I_19366 (I334429,I334754,I334895);
nor I_19367 (I334417,I334895,I334658);
not I_19368 (I334971,I334895);
and I_19369 (I334988,I334522,I334971);
nor I_19370 (I334423,I334658,I334988);
nand I_19371 (I334411,I334895,I334785);
not I_19372 (I335066_rst,I5701);
not I_19373 (I335083,I292055);
nor I_19374 (I335100,I292058,I292067);
nand I_19375 (I335117,I335100,I292082);
nor I_19376 (I335134,I335083,I292058);
nand I_19377 (I335151,I335134,I292061);
not I_19378 (I335168,I292058);
not I_19379 (I335185,I335168);
not I_19380 (I335202,I292052);
nor I_19381 (I335219,I335202,I292076);
and I_19382 (I335236,I335219,I292064);
or I_19383 (I335253,I335236,I292070);
DFFARX1 I_19384  ( .D(I335253), .CLK(I5694_clk), .RSTB(I335066_rst), .Q(I335270) );
nand I_19385 (I335287,I335083,I292052);
or I_19386 (I335055,I335287,I335270);
not I_19387 (I335318,I335287);
nor I_19388 (I335335,I335270,I335318);
and I_19389 (I335352,I335168,I335335);
nand I_19390 (I335028,I335287,I335185);
DFFARX1 I_19391  ( .D(I292073), .CLK(I5694_clk), .RSTB(I335066_rst), .Q(I335383) );
or I_19392 (I335049,I335383,I335270);
nor I_19393 (I335414,I335383,I335151);
nor I_19394 (I335431,I335383,I335185);
nand I_19395 (I335034,I335117,I335431);
or I_19396 (I335462,I335383,I335352);
DFFARX1 I_19397  ( .D(I335462), .CLK(I5694_clk), .RSTB(I335066_rst), .Q(I335031) );
not I_19398 (I335037,I335383);
DFFARX1 I_19399  ( .D(I292079), .CLK(I5694_clk), .RSTB(I335066_rst), .Q(I335507) );
not I_19400 (I335524,I335507);
nor I_19401 (I335541,I335524,I335117);
DFFARX1 I_19402  ( .D(I335541), .CLK(I5694_clk), .RSTB(I335066_rst), .Q(I335043) );
nor I_19403 (I335058,I335383,I335524);
nor I_19404 (I335046,I335524,I335287);
not I_19405 (I335600,I335524);
and I_19406 (I335617,I335151,I335600);
nor I_19407 (I335052,I335287,I335617);
nand I_19408 (I335040,I335524,I335414);
not I_19409 (I335695_rst,I5701);
not I_19410 (I335712,I313575);
nor I_19411 (I335729,I313581,I313560);
nand I_19412 (I335746,I335729,I313566);
nor I_19413 (I335763,I335712,I313581);
nand I_19414 (I335780,I335763,I313572);
not I_19415 (I335797,I313581);
not I_19416 (I335814,I335797);
not I_19417 (I335831,I313569);
nor I_19418 (I335848,I335831,I313587);
and I_19419 (I335865,I335848,I313578);
or I_19420 (I335882,I335865,I313557);
DFFARX1 I_19421  ( .D(I335882), .CLK(I5694_clk), .RSTB(I335695_rst), .Q(I335899) );
nand I_19422 (I335916,I335712,I313569);
or I_19423 (I335684,I335916,I335899);
not I_19424 (I335947,I335916);
nor I_19425 (I335964,I335899,I335947);
and I_19426 (I335981,I335797,I335964);
nand I_19427 (I335657,I335916,I335814);
DFFARX1 I_19428  ( .D(I313584), .CLK(I5694_clk), .RSTB(I335695_rst), .Q(I336012) );
or I_19429 (I335678,I336012,I335899);
nor I_19430 (I336043,I336012,I335780);
nor I_19431 (I336060,I336012,I335814);
nand I_19432 (I335663,I335746,I336060);
or I_19433 (I336091,I336012,I335981);
DFFARX1 I_19434  ( .D(I336091), .CLK(I5694_clk), .RSTB(I335695_rst), .Q(I335660) );
not I_19435 (I335666,I336012);
DFFARX1 I_19436  ( .D(I313563), .CLK(I5694_clk), .RSTB(I335695_rst), .Q(I336136) );
not I_19437 (I336153,I336136);
nor I_19438 (I336170,I336153,I335746);
DFFARX1 I_19439  ( .D(I336170), .CLK(I5694_clk), .RSTB(I335695_rst), .Q(I335672) );
nor I_19440 (I335687,I336012,I336153);
nor I_19441 (I335675,I336153,I335916);
not I_19442 (I336229,I336153);
and I_19443 (I336246,I335780,I336229);
nor I_19444 (I335681,I335916,I336246);
nand I_19445 (I335669,I336153,I336043);
not I_19446 (I336324_rst,I5701);
not I_19447 (I336341,I286380);
nor I_19448 (I336358,I286404,I286389);
nand I_19449 (I336375,I336358,I286374);
nor I_19450 (I336392,I336341,I286404);
nand I_19451 (I336409,I336392,I286401);
not I_19452 (I336426,I286404);
not I_19453 (I336443,I336426);
not I_19454 (I336460,I286383);
nor I_19455 (I336477,I336460,I286377);
and I_19456 (I336494,I336477,I286398);
or I_19457 (I336511,I336494,I286386);
DFFARX1 I_19458  ( .D(I336511), .CLK(I5694_clk), .RSTB(I336324_rst), .Q(I336528) );
nand I_19459 (I336545,I336341,I286383);
or I_19460 (I336313,I336545,I336528);
not I_19461 (I336576,I336545);
nor I_19462 (I336593,I336528,I336576);
and I_19463 (I336610,I336426,I336593);
nand I_19464 (I336286,I336545,I336443);
DFFARX1 I_19465  ( .D(I286395), .CLK(I5694_clk), .RSTB(I336324_rst), .Q(I336641) );
or I_19466 (I336307,I336641,I336528);
nor I_19467 (I336672,I336641,I336409);
nor I_19468 (I336689,I336641,I336443);
nand I_19469 (I336292,I336375,I336689);
or I_19470 (I336720,I336641,I336610);
DFFARX1 I_19471  ( .D(I336720), .CLK(I5694_clk), .RSTB(I336324_rst), .Q(I336289) );
not I_19472 (I336295,I336641);
DFFARX1 I_19473  ( .D(I286392), .CLK(I5694_clk), .RSTB(I336324_rst), .Q(I336765) );
not I_19474 (I336782,I336765);
nor I_19475 (I336799,I336782,I336375);
DFFARX1 I_19476  ( .D(I336799), .CLK(I5694_clk), .RSTB(I336324_rst), .Q(I336301) );
nor I_19477 (I336316,I336641,I336782);
nor I_19478 (I336304,I336782,I336545);
not I_19479 (I336858,I336782);
and I_19480 (I336875,I336409,I336858);
nor I_19481 (I336310,I336545,I336875);
nand I_19482 (I336298,I336782,I336672);
not I_19483 (I336953_rst,I5701);
not I_19484 (I336970,I301516);
nor I_19485 (I336987,I301507,I301531);
nand I_19486 (I337004,I336987,I301534);
nor I_19487 (I337021,I336970,I301507);
nand I_19488 (I337038,I337021,I301525);
not I_19489 (I337055,I301507);
not I_19490 (I337072,I337055);
not I_19491 (I337089,I301519);
nor I_19492 (I337106,I337089,I301513);
and I_19493 (I337123,I337106,I301522);
or I_19494 (I337140,I337123,I301510);
DFFARX1 I_19495  ( .D(I337140), .CLK(I5694_clk), .RSTB(I336953_rst), .Q(I337157) );
nand I_19496 (I337174,I336970,I301519);
or I_19497 (I336942,I337174,I337157);
not I_19498 (I337205,I337174);
nor I_19499 (I337222,I337157,I337205);
and I_19500 (I337239,I337055,I337222);
nand I_19501 (I336915,I337174,I337072);
DFFARX1 I_19502  ( .D(I301504), .CLK(I5694_clk), .RSTB(I336953_rst), .Q(I337270) );
or I_19503 (I336936,I337270,I337157);
nor I_19504 (I337301,I337270,I337038);
nor I_19505 (I337318,I337270,I337072);
nand I_19506 (I336921,I337004,I337318);
or I_19507 (I337349,I337270,I337239);
DFFARX1 I_19508  ( .D(I337349), .CLK(I5694_clk), .RSTB(I336953_rst), .Q(I336918) );
not I_19509 (I336924,I337270);
DFFARX1 I_19510  ( .D(I301528), .CLK(I5694_clk), .RSTB(I336953_rst), .Q(I337394) );
not I_19511 (I337411,I337394);
nor I_19512 (I337428,I337411,I337004);
DFFARX1 I_19513  ( .D(I337428), .CLK(I5694_clk), .RSTB(I336953_rst), .Q(I336930) );
nor I_19514 (I336945,I337270,I337411);
nor I_19515 (I336933,I337411,I337174);
not I_19516 (I337487,I337411);
and I_19517 (I337504,I337038,I337487);
nor I_19518 (I336939,I337174,I337504);
nand I_19519 (I336927,I337411,I337301);
not I_19520 (I337582_rst,I5701);
nand I_19521 (I337599,I320752,I320749);
and I_19522 (I337616,I337599,I320731);
DFFARX1 I_19523  ( .D(I337616), .CLK(I5694_clk), .RSTB(I337582_rst), .Q(I337633) );
not I_19524 (I337571,I337633);
DFFARX1 I_19525  ( .D(I337633), .CLK(I5694_clk), .RSTB(I337582_rst), .Q(I337664) );
not I_19526 (I337559,I337664);
nor I_19527 (I337695,I320761,I320749);
not I_19528 (I337712,I337695);
nor I_19529 (I337729,I337633,I337712);
DFFARX1 I_19530  ( .D(I320737), .CLK(I5694_clk), .RSTB(I337582_rst), .Q(I337746) );
not I_19531 (I337763,I337746);
nand I_19532 (I337562,I337746,I337712);
DFFARX1 I_19533  ( .D(I337746), .CLK(I5694_clk), .RSTB(I337582_rst), .Q(I337794) );
and I_19534 (I337547,I337633,I337794);
nand I_19535 (I337825,I320758,I320755);
and I_19536 (I337842,I337825,I320740);
DFFARX1 I_19537  ( .D(I337842), .CLK(I5694_clk), .RSTB(I337582_rst), .Q(I337859) );
nor I_19538 (I337876,I337859,I337763);
and I_19539 (I337893,I337695,I337876);
nor I_19540 (I337910,I337859,I337633);
DFFARX1 I_19541  ( .D(I337859), .CLK(I5694_clk), .RSTB(I337582_rst), .Q(I337553) );
DFFARX1 I_19542  ( .D(I320743), .CLK(I5694_clk), .RSTB(I337582_rst), .Q(I337941) );
and I_19543 (I337958,I337941,I320746);
or I_19544 (I337975,I337958,I337893);
DFFARX1 I_19545  ( .D(I337975), .CLK(I5694_clk), .RSTB(I337582_rst), .Q(I337565) );
nand I_19546 (I337574,I337958,I337910);
DFFARX1 I_19547  ( .D(I337958), .CLK(I5694_clk), .RSTB(I337582_rst), .Q(I337544) );
DFFARX1 I_19548  ( .D(I320734), .CLK(I5694_clk), .RSTB(I337582_rst), .Q(I338034) );
nand I_19549 (I337568,I338034,I337729);
DFFARX1 I_19550  ( .D(I338034), .CLK(I5694_clk), .RSTB(I337582_rst), .Q(I337556) );
nand I_19551 (I338079,I338034,I337695);
and I_19552 (I338096,I337746,I338079);
DFFARX1 I_19553  ( .D(I338096), .CLK(I5694_clk), .RSTB(I337582_rst), .Q(I337550) );
not I_19554 (I338160_rst,I5701);
nand I_19555 (I338177,I333144,I333162);
and I_19556 (I338194,I338177,I333159);
DFFARX1 I_19557  ( .D(I338194), .CLK(I5694_clk), .RSTB(I338160_rst), .Q(I338211) );
not I_19558 (I338149,I338211);
DFFARX1 I_19559  ( .D(I338211), .CLK(I5694_clk), .RSTB(I338160_rst), .Q(I338242) );
not I_19560 (I338137,I338242);
nor I_19561 (I338273,I333165,I333162);
not I_19562 (I338290,I338273);
nor I_19563 (I338307,I338211,I338290);
DFFARX1 I_19564  ( .D(I333168), .CLK(I5694_clk), .RSTB(I338160_rst), .Q(I338324) );
not I_19565 (I338341,I338324);
nand I_19566 (I338140,I338324,I338290);
DFFARX1 I_19567  ( .D(I338324), .CLK(I5694_clk), .RSTB(I338160_rst), .Q(I338372) );
and I_19568 (I338125,I338211,I338372);
nand I_19569 (I338403,I333153,I333147);
and I_19570 (I338420,I338403,I333150);
DFFARX1 I_19571  ( .D(I338420), .CLK(I5694_clk), .RSTB(I338160_rst), .Q(I338437) );
nor I_19572 (I338454,I338437,I338341);
and I_19573 (I338471,I338273,I338454);
nor I_19574 (I338488,I338437,I338211);
DFFARX1 I_19575  ( .D(I338437), .CLK(I5694_clk), .RSTB(I338160_rst), .Q(I338131) );
DFFARX1 I_19576  ( .D(I333156), .CLK(I5694_clk), .RSTB(I338160_rst), .Q(I338519) );
and I_19577 (I338536,I338519,I333141);
or I_19578 (I338553,I338536,I338471);
DFFARX1 I_19579  ( .D(I338553), .CLK(I5694_clk), .RSTB(I338160_rst), .Q(I338143) );
nand I_19580 (I338152,I338536,I338488);
DFFARX1 I_19581  ( .D(I338536), .CLK(I5694_clk), .RSTB(I338160_rst), .Q(I338122) );
DFFARX1 I_19582  ( .D(I333171), .CLK(I5694_clk), .RSTB(I338160_rst), .Q(I338612) );
nand I_19583 (I338146,I338612,I338307);
DFFARX1 I_19584  ( .D(I338612), .CLK(I5694_clk), .RSTB(I338160_rst), .Q(I338134) );
nand I_19585 (I338657,I338612,I338273);
and I_19586 (I338674,I338324,I338657);
DFFARX1 I_19587  ( .D(I338674), .CLK(I5694_clk), .RSTB(I338160_rst), .Q(I338128) );
not I_19588 (I338738_rst,I5701);
nand I_19589 (I338755,I294402,I294387);
and I_19590 (I33877_rst2,I338755,I294381);
DFFARX1 I_19591  ( .D(I33877_rst2), .CLK(I5694_clk), .RSTB(I338738_rst), .Q(I338789) );
not I_19592 (I338727,I338789);
DFFARX1 I_19593  ( .D(I338789), .CLK(I5694_clk), .RSTB(I338738_rst), .Q(I338820) );
not I_19594 (I338715,I338820);
nor I_19595 (I338851,I294408,I294387);
not I_19596 (I338868,I338851);
nor I_19597 (I338885,I338789,I338868);
DFFARX1 I_19598  ( .D(I294411), .CLK(I5694_clk), .RSTB(I338738_rst), .Q(I338902) );
not I_19599 (I338919,I338902);
nand I_19600 (I338718,I338902,I338868);
DFFARX1 I_19601  ( .D(I338902), .CLK(I5694_clk), .RSTB(I338738_rst), .Q(I338950) );
and I_19602 (I338703,I338789,I338950);
nand I_19603 (I338981,I294393,I294396);
and I_19604 (I338998,I338981,I294399);
DFFARX1 I_19605  ( .D(I338998), .CLK(I5694_clk), .RSTB(I338738_rst), .Q(I339015) );
nor I_19606 (I339032,I339015,I338919);
and I_19607 (I339049,I338851,I339032);
nor I_19608 (I339066,I339015,I338789);
DFFARX1 I_19609  ( .D(I339015), .CLK(I5694_clk), .RSTB(I338738_rst), .Q(I338709) );
DFFARX1 I_19610  ( .D(I294405), .CLK(I5694_clk), .RSTB(I338738_rst), .Q(I339097) );
and I_19611 (I339114,I339097,I294390);
or I_19612 (I339131,I339114,I339049);
DFFARX1 I_19613  ( .D(I339131), .CLK(I5694_clk), .RSTB(I338738_rst), .Q(I338721) );
nand I_19614 (I338730,I339114,I339066);
DFFARX1 I_19615  ( .D(I339114), .CLK(I5694_clk), .RSTB(I338738_rst), .Q(I338700) );
DFFARX1 I_19616  ( .D(I294384), .CLK(I5694_clk), .RSTB(I338738_rst), .Q(I339190) );
nand I_19617 (I338724,I339190,I338885);
DFFARX1 I_19618  ( .D(I339190), .CLK(I5694_clk), .RSTB(I338738_rst), .Q(I338712) );
nand I_19619 (I339235,I339190,I338851);
and I_19620 (I339252,I338902,I339235);
DFFARX1 I_19621  ( .D(I339252), .CLK(I5694_clk), .RSTB(I338738_rst), .Q(I338706) );
not I_19622 (I339316_rst,I5701);
nand I_19623 (I339333,I336286,I336289);
and I_19624 (I339350,I339333,I336295);
DFFARX1 I_19625  ( .D(I339350), .CLK(I5694_clk), .RSTB(I339316_rst), .Q(I339367) );
not I_19626 (I339384,I339367);
nor I_19627 (I339401,I336307,I336289);
or I_19628 (I339299,I339401,I339367);
not I_19629 (I339287,I339401);
DFFARX1 I_19630  ( .D(I336316), .CLK(I5694_clk), .RSTB(I339316_rst), .Q(I339446) );
nor I_19631 (I339463,I339446,I339401);
nand I_19632 (I339480,I336304,I336301);
and I_19633 (I339497,I339480,I336313);
DFFARX1 I_19634  ( .D(I339497), .CLK(I5694_clk), .RSTB(I339316_rst), .Q(I339514) );
nor I_19635 (I339296,I339514,I339367);
not I_19636 (I339545,I339514);
nor I_19637 (I339562,I339446,I339545);
DFFARX1 I_19638  ( .D(I336310), .CLK(I5694_clk), .RSTB(I339316_rst), .Q(I339579) );
and I_19639 (I339596,I339579,I336298);
or I_19640 (I339305,I339596,I339401);
nand I_19641 (I339284,I339596,I339562);
DFFARX1 I_19642  ( .D(I336292), .CLK(I5694_clk), .RSTB(I339316_rst), .Q(I339641) );
and I_19643 (I339658,I339641,I339384);
nor I_19644 (I339302,I339596,I339658);
nor I_19645 (I339689,I339641,I339446);
DFFARX1 I_19646  ( .D(I339689), .CLK(I5694_clk), .RSTB(I339316_rst), .Q(I339293) );
nor I_19647 (I339308,I339641,I339367);
not I_19648 (I339734,I339641);
nor I_19649 (I339751,I339514,I339734);
and I_19650 (I339768,I339401,I339751);
or I_19651 (I339785,I339596,I339768);
DFFARX1 I_19652  ( .D(I339785), .CLK(I5694_clk), .RSTB(I339316_rst), .Q(I339281) );
nand I_19653 (I339290,I339641,I339463);
nand I_19654 (I339278,I339641,I339545);
not I_19655 (I339877_rst,I5701);
nand I_19656 (I339894,I296986,I296989);
and I_19657 (I339911,I339894,I296971);
DFFARX1 I_19658  ( .D(I339911), .CLK(I5694_clk), .RSTB(I339877_rst), .Q(I339928) );
not I_19659 (I339945,I339928);
nor I_19660 (I339962,I296968,I296989);
or I_19661 (I339860,I339962,I339928);
not I_19662 (I339848,I339962);
DFFARX1 I_19663  ( .D(I296992), .CLK(I5694_clk), .RSTB(I339877_rst), .Q(I340007) );
nor I_19664 (I340024,I340007,I339962);
nand I_19665 (I340041,I296977,I296983);
and I_19666 (I340058,I340041,I296995);
DFFARX1 I_19667  ( .D(I340058), .CLK(I5694_clk), .RSTB(I339877_rst), .Q(I340075) );
nor I_19668 (I339857,I340075,I339928);
not I_19669 (I340106,I340075);
nor I_19670 (I340123,I340007,I340106);
DFFARX1 I_19671  ( .D(I296974), .CLK(I5694_clk), .RSTB(I339877_rst), .Q(I340140) );
and I_19672 (I340157,I340140,I296965);
or I_19673 (I339866,I340157,I339962);
nand I_19674 (I339845,I340157,I340123);
DFFARX1 I_19675  ( .D(I296980), .CLK(I5694_clk), .RSTB(I339877_rst), .Q(I340202) );
and I_19676 (I340219,I340202,I339945);
nor I_19677 (I339863,I340157,I340219);
nor I_19678 (I340250,I340202,I340007);
DFFARX1 I_19679  ( .D(I340250), .CLK(I5694_clk), .RSTB(I339877_rst), .Q(I339854) );
nor I_19680 (I339869,I340202,I339928);
not I_19681 (I340295,I340202);
nor I_19682 (I340312,I340075,I340295);
and I_19683 (I340329,I339962,I340312);
or I_19684 (I340346,I340157,I340329);
DFFARX1 I_19685  ( .D(I340346), .CLK(I5694_clk), .RSTB(I339877_rst), .Q(I339842) );
nand I_19686 (I339851,I340202,I340024);
nand I_19687 (I339839,I340202,I340106);
not I_19688 (I340438_rst,I5701);
nand I_19689 (I340455,I314907,I314898);
and I_19690 (I340472,I340455,I314913);
DFFARX1 I_19691  ( .D(I340472), .CLK(I5694_clk), .RSTB(I340438_rst), .Q(I340489) );
not I_19692 (I340506,I340489);
nor I_19693 (I340523,I314883,I314898);
or I_19694 (I340421,I340523,I340489);
not I_19695 (I340409,I340523);
DFFARX1 I_19696  ( .D(I314886), .CLK(I5694_clk), .RSTB(I340438_rst), .Q(I340568) );
nor I_19697 (I340585,I340568,I340523);
nand I_19698 (I340602,I314904,I314901);
and I_19699 (I340619,I340602,I314889);
DFFARX1 I_19700  ( .D(I340619), .CLK(I5694_clk), .RSTB(I340438_rst), .Q(I340636) );
nor I_19701 (I340418,I340636,I340489);
not I_19702 (I340667,I340636);
nor I_19703 (I340684,I340568,I340667);
DFFARX1 I_19704  ( .D(I314910), .CLK(I5694_clk), .RSTB(I340438_rst), .Q(I340701) );
and I_19705 (I340718,I340701,I314895);
or I_19706 (I340427,I340718,I340523);
nand I_19707 (I340406,I340718,I340684);
DFFARX1 I_19708  ( .D(I314892), .CLK(I5694_clk), .RSTB(I340438_rst), .Q(I340763) );
and I_19709 (I340780,I340763,I340506);
nor I_19710 (I340424,I340718,I340780);
nor I_19711 (I340811,I340763,I340568);
DFFARX1 I_19712  ( .D(I340811), .CLK(I5694_clk), .RSTB(I340438_rst), .Q(I340415) );
nor I_19713 (I340430,I340763,I340489);
not I_19714 (I340856,I340763);
nor I_19715 (I340873,I340636,I340856);
and I_19716 (I340890,I340523,I340873);
or I_19717 (I340907,I340718,I340890);
DFFARX1 I_19718  ( .D(I340907), .CLK(I5694_clk), .RSTB(I340438_rst), .Q(I340403) );
nand I_19719 (I340412,I340763,I340585);
nand I_19720 (I340400,I340763,I340667);
not I_19721 (I340999_rst,I5701);
nand I_19722 (I341016,I300850,I300847);
and I_19723 (I341033,I341016,I300844);
DFFARX1 I_19724  ( .D(I341033), .CLK(I5694_clk), .RSTB(I340999_rst), .Q(I341050) );
not I_19725 (I341067,I341050);
nor I_19726 (I341084,I300868,I300847);
or I_19727 (I340982,I341084,I341050);
not I_19728 (I340970,I341084);
DFFARX1 I_19729  ( .D(I300862), .CLK(I5694_clk), .RSTB(I340999_rst), .Q(I341129) );
nor I_19730 (I341146,I341129,I341084);
nand I_19731 (I341163,I300841,I300853);
and I_19732 (I341180,I341163,I300856);
DFFARX1 I_19733  ( .D(I341180), .CLK(I5694_clk), .RSTB(I340999_rst), .Q(I341197) );
nor I_19734 (I340979,I341197,I341050);
not I_19735 (I341228,I341197);
nor I_19736 (I341245,I341129,I341228);
DFFARX1 I_19737  ( .D(I300865), .CLK(I5694_clk), .RSTB(I340999_rst), .Q(I341262) );
and I_19738 (I341279,I341262,I300871);
or I_19739 (I340988,I341279,I341084);
nand I_19740 (I340967,I341279,I341245);
DFFARX1 I_19741  ( .D(I300859), .CLK(I5694_clk), .RSTB(I340999_rst), .Q(I341324) );
and I_19742 (I341341,I341324,I341067);
nor I_19743 (I340985,I341279,I341341);
nor I_19744 (I341372,I341324,I341129);
DFFARX1 I_19745  ( .D(I341372), .CLK(I5694_clk), .RSTB(I340999_rst), .Q(I340976) );
nor I_19746 (I340991,I341324,I341050);
not I_19747 (I341417,I341324);
nor I_19748 (I341434,I341197,I341417);
and I_19749 (I341451,I341084,I341434);
or I_19750 (I341468,I341279,I341451);
DFFARX1 I_19751  ( .D(I341468), .CLK(I5694_clk), .RSTB(I340999_rst), .Q(I340964) );
nand I_19752 (I340973,I341324,I341146);
nand I_19753 (I340961,I341324,I341228);
not I_19754 (I341560_rst,I5701);
nand I_19755 (I341577,I322511,I322508);
and I_19756 (I341594,I341577,I322502);
DFFARX1 I_19757  ( .D(I341594), .CLK(I5694_clk), .RSTB(I341560_rst), .Q(I341611) );
not I_19758 (I341628,I341611);
nor I_19759 (I341645,I322514,I322508);
or I_19760 (I341543,I341645,I341611);
not I_19761 (I341531,I341645);
DFFARX1 I_19762  ( .D(I322526), .CLK(I5694_clk), .RSTB(I341560_rst), .Q(I341690) );
nor I_19763 (I341707,I341690,I341645);
nand I_19764 (I341724,I322517,I322499);
and I_19765 (I341741,I341724,I322529);
DFFARX1 I_19766  ( .D(I341741), .CLK(I5694_clk), .RSTB(I341560_rst), .Q(I341758) );
nor I_19767 (I341540,I341758,I341611);
not I_19768 (I341789,I341758);
nor I_19769 (I341806,I341690,I341789);
DFFARX1 I_19770  ( .D(I322505), .CLK(I5694_clk), .RSTB(I341560_rst), .Q(I341823) );
and I_19771 (I341840,I341823,I322523);
or I_19772 (I341549,I341840,I341645);
nand I_19773 (I341528,I341840,I341806);
DFFARX1 I_19774  ( .D(I322520), .CLK(I5694_clk), .RSTB(I341560_rst), .Q(I341885) );
and I_19775 (I341902,I341885,I341628);
nor I_19776 (I341546,I341840,I341902);
nor I_19777 (I341933,I341885,I341690);
DFFARX1 I_19778  ( .D(I341933), .CLK(I5694_clk), .RSTB(I341560_rst), .Q(I341537) );
nor I_19779 (I341552,I341885,I341611);
not I_19780 (I341978,I341885);
nor I_19781 (I341995,I341758,I341978);
and I_19782 (I342012,I341645,I341995);
or I_19783 (I342029,I341840,I342012);
DFFARX1 I_19784  ( .D(I342029), .CLK(I5694_clk), .RSTB(I341560_rst), .Q(I341525) );
nand I_19785 (I341534,I341885,I341707);
nand I_19786 (I341522,I341885,I341789);
not I_19787 (I342121_rst,I5701);
not I_19788 (I342138,I302848);
nor I_19789 (I342155,I302836,I302842);
nand I_19790 (I342172,I342155,I302851);
DFFARX1 I_19791  ( .D(I342172), .CLK(I5694_clk), .RSTB(I342121_rst), .Q(I342095) );
nor I_19792 (I342203,I342138,I302836);
nand I_19793 (I342220,I342203,I302839);
not I_19794 (I342110,I342220);
DFFARX1 I_19795  ( .D(I342220), .CLK(I5694_clk), .RSTB(I342121_rst), .Q(I342092) );
not I_19796 (I342265,I302836);
not I_19797 (I342282,I342265);
not I_19798 (I342299,I302860);
nor I_19799 (I342316,I342299,I302833);
and I_19800 (I342333,I342316,I302854);
or I_19801 (I342350,I342333,I302845);
DFFARX1 I_19802  ( .D(I342350), .CLK(I5694_clk), .RSTB(I342121_rst), .Q(I342367) );
nor I_19803 (I342384,I342367,I342220);
nor I_19804 (I342401,I342367,I342282);
nand I_19805 (I342107,I342172,I342401);
nand I_19806 (I342432,I342138,I302860);
nand I_19807 (I342449,I342432,I342367);
and I_19808 (I342466,I342432,I342449);
DFFARX1 I_19809  ( .D(I342466), .CLK(I5694_clk), .RSTB(I342121_rst), .Q(I342089) );
DFFARX1 I_19810  ( .D(I342432), .CLK(I5694_clk), .RSTB(I342121_rst), .Q(I342497) );
and I_19811 (I342086,I342265,I342497);
DFFARX1 I_19812  ( .D(I302830), .CLK(I5694_clk), .RSTB(I342121_rst), .Q(I342528) );
not I_19813 (I342545,I342528);
nor I_19814 (I342562,I342220,I342545);
and I_19815 (I342579,I342528,I342562);
nand I_19816 (I342101,I342528,I342282);
DFFARX1 I_19817  ( .D(I342528), .CLK(I5694_clk), .RSTB(I342121_rst), .Q(I342610) );
not I_19818 (I342098,I342610);
DFFARX1 I_19819  ( .D(I302857), .CLK(I5694_clk), .RSTB(I342121_rst), .Q(I342641) );
not I_19820 (I342658,I342641);
or I_19821 (I342675,I342658,I342579);
DFFARX1 I_19822  ( .D(I342675), .CLK(I5694_clk), .RSTB(I342121_rst), .Q(I342104) );
nand I_19823 (I342113,I342658,I342384);
DFFARX1 I_19824  ( .D(I342658), .CLK(I5694_clk), .RSTB(I342121_rst), .Q(I342083) );
not I_19825 (I342767_rst,I5701);
not I_19826 (I342784,I339842);
nor I_19827 (I342801,I339854,I339839);
nand I_19828 (I342818,I342801,I339851);
DFFARX1 I_19829  ( .D(I342818), .CLK(I5694_clk), .RSTB(I342767_rst), .Q(I342741) );
nor I_19830 (I342849,I342784,I339854);
nand I_19831 (I342866,I342849,I339869);
not I_19832 (I342756,I342866);
DFFARX1 I_19833  ( .D(I342866), .CLK(I5694_clk), .RSTB(I342767_rst), .Q(I342738) );
not I_19834 (I342911,I339854);
not I_19835 (I342928,I342911);
not I_19836 (I342945,I339845);
nor I_19837 (I342962,I342945,I339857);
and I_19838 (I342979,I342962,I339848);
or I_19839 (I342996,I342979,I339863);
DFFARX1 I_19840  ( .D(I342996), .CLK(I5694_clk), .RSTB(I342767_rst), .Q(I343013) );
nor I_19841 (I343030,I343013,I342866);
nor I_19842 (I343047,I343013,I342928);
nand I_19843 (I342753,I342818,I343047);
nand I_19844 (I343078,I342784,I339845);
nand I_19845 (I343095,I343078,I343013);
and I_19846 (I343112,I343078,I343095);
DFFARX1 I_19847  ( .D(I343112), .CLK(I5694_clk), .RSTB(I342767_rst), .Q(I342735) );
DFFARX1 I_19848  ( .D(I343078), .CLK(I5694_clk), .RSTB(I342767_rst), .Q(I343143) );
and I_19849 (I342732,I342911,I343143);
DFFARX1 I_19850  ( .D(I339866), .CLK(I5694_clk), .RSTB(I342767_rst), .Q(I343174) );
not I_19851 (I343191,I343174);
nor I_19852 (I343208,I342866,I343191);
and I_19853 (I343225,I343174,I343208);
nand I_19854 (I342747,I343174,I342928);
DFFARX1 I_19855  ( .D(I343174), .CLK(I5694_clk), .RSTB(I342767_rst), .Q(I343256) );
not I_19856 (I342744,I343256);
DFFARX1 I_19857  ( .D(I339860), .CLK(I5694_clk), .RSTB(I342767_rst), .Q(I343287) );
not I_19858 (I343304,I343287);
or I_19859 (I343321,I343304,I343225);
DFFARX1 I_19860  ( .D(I343321), .CLK(I5694_clk), .RSTB(I342767_rst), .Q(I342750) );
nand I_19861 (I342759,I343304,I343030);
DFFARX1 I_19862  ( .D(I343304), .CLK(I5694_clk), .RSTB(I342767_rst), .Q(I342729) );
not I_19863 (I343413_rst,I5701);
not I_19864 (I343430,I316227);
nor I_19865 (I343447,I316239,I316221);
nand I_19866 (I343464,I343447,I316236);
DFFARX1 I_19867  ( .D(I343464), .CLK(I5694_clk), .RSTB(I343413_rst), .Q(I343387) );
nor I_19868 (I343495,I343430,I316239);
nand I_19869 (I343512,I343495,I316224);
not I_19870 (I343402,I343512);
DFFARX1 I_19871  ( .D(I343512), .CLK(I5694_clk), .RSTB(I343413_rst), .Q(I343384) );
not I_19872 (I343557,I316239);
not I_19873 (I343574,I343557);
not I_19874 (I343591,I316233);
nor I_19875 (I343608,I343591,I316212);
and I_19876 (I343625,I343608,I316215);
or I_19877 (I343642,I343625,I316218);
DFFARX1 I_19878  ( .D(I343642), .CLK(I5694_clk), .RSTB(I343413_rst), .Q(I343659) );
nor I_19879 (I343676,I343659,I343512);
nor I_19880 (I343693,I343659,I343574);
nand I_19881 (I343399,I343464,I343693);
nand I_19882 (I343724,I343430,I316233);
nand I_19883 (I343741,I343724,I343659);
and I_19884 (I343758,I343724,I343741);
DFFARX1 I_19885  ( .D(I343758), .CLK(I5694_clk), .RSTB(I343413_rst), .Q(I343381) );
DFFARX1 I_19886  ( .D(I343724), .CLK(I5694_clk), .RSTB(I343413_rst), .Q(I343789) );
and I_19887 (I343378,I343557,I343789);
DFFARX1 I_19888  ( .D(I316209), .CLK(I5694_clk), .RSTB(I343413_rst), .Q(I343820) );
not I_19889 (I343837,I343820);
nor I_19890 (I343854,I343512,I343837);
and I_19891 (I343871,I343820,I343854);
nand I_19892 (I343393,I343820,I343574);
DFFARX1 I_19893  ( .D(I343820), .CLK(I5694_clk), .RSTB(I343413_rst), .Q(I343902) );
not I_19894 (I343390,I343902);
DFFARX1 I_19895  ( .D(I316230), .CLK(I5694_clk), .RSTB(I343413_rst), .Q(I343933) );
not I_19896 (I343950,I343933);
or I_19897 (I343967,I343950,I343871);
DFFARX1 I_19898  ( .D(I343967), .CLK(I5694_clk), .RSTB(I343413_rst), .Q(I343396) );
nand I_19899 (I343405,I343950,I343676);
DFFARX1 I_19900  ( .D(I343950), .CLK(I5694_clk), .RSTB(I343413_rst), .Q(I343375) );
not I_19901 (I344059_rst,I5701);
not I_19902 (I344076,I312249);
nor I_19903 (I344093,I312246,I312234);
nand I_19904 (I344110,I344093,I312237);
DFFARX1 I_19905  ( .D(I344110), .CLK(I5694_clk), .RSTB(I344059_rst), .Q(I344033) );
nor I_19906 (I344141,I344076,I312246);
nand I_19907 (I344158,I344141,I312243);
not I_19908 (I344048,I344158);
DFFARX1 I_19909  ( .D(I344158), .CLK(I5694_clk), .RSTB(I344059_rst), .Q(I344030) );
not I_19910 (I344203,I312246);
not I_19911 (I344220,I344203);
not I_19912 (I344237,I312255);
nor I_19913 (I344254,I344237,I312231);
and I_19914 (I344271,I344254,I312252);
or I_19915 (I344288,I344271,I312240);
DFFARX1 I_19916  ( .D(I344288), .CLK(I5694_clk), .RSTB(I344059_rst), .Q(I344305) );
nor I_19917 (I344322,I344305,I344158);
nor I_19918 (I344339,I344305,I344220);
nand I_19919 (I344045,I344110,I344339);
nand I_19920 (I344370,I344076,I312255);
nand I_19921 (I344387,I344370,I344305);
and I_19922 (I344404,I344370,I344387);
DFFARX1 I_19923  ( .D(I344404), .CLK(I5694_clk), .RSTB(I344059_rst), .Q(I344027) );
DFFARX1 I_19924  ( .D(I344370), .CLK(I5694_clk), .RSTB(I344059_rst), .Q(I344435) );
and I_19925 (I344024,I344203,I344435);
DFFARX1 I_19926  ( .D(I312261), .CLK(I5694_clk), .RSTB(I344059_rst), .Q(I344466) );
not I_19927 (I344483,I344466);
nor I_19928 (I344500,I344158,I344483);
and I_19929 (I344517,I344466,I344500);
nand I_19930 (I344039,I344466,I344220);
DFFARX1 I_19931  ( .D(I344466), .CLK(I5694_clk), .RSTB(I344059_rst), .Q(I344548) );
not I_19932 (I344036,I344548);
DFFARX1 I_19933  ( .D(I312258), .CLK(I5694_clk), .RSTB(I344059_rst), .Q(I344579) );
not I_19934 (I344596,I344579);
or I_19935 (I344613,I344596,I344517);
DFFARX1 I_19936  ( .D(I344613), .CLK(I5694_clk), .RSTB(I344059_rst), .Q(I344042) );
nand I_19937 (I344051,I344596,I344322);
DFFARX1 I_19938  ( .D(I344596), .CLK(I5694_clk), .RSTB(I344059_rst), .Q(I344021) );
not I_19939 (I344705_rst,I5701);
not I_19940 (I344722,I325994);
nor I_19941 (I344739,I325970,I325976);
nand I_19942 (I344756,I344739,I325979);
DFFARX1 I_19943  ( .D(I344756), .CLK(I5694_clk), .RSTB(I344705_rst), .Q(I344679) );
nor I_19944 (I344787,I344722,I325970);
nand I_19945 (I344804,I344787,I325988);
not I_19946 (I344694,I344804);
DFFARX1 I_19947  ( .D(I344804), .CLK(I5694_clk), .RSTB(I344705_rst), .Q(I344676) );
not I_19948 (I344849,I325970);
not I_19949 (I344866,I344849);
not I_19950 (I344883,I325967);
nor I_19951 (I344900,I344883,I325982);
and I_19952 (I344917,I344900,I325973);
or I_19953 (I344934,I344917,I325985);
DFFARX1 I_19954  ( .D(I344934), .CLK(I5694_clk), .RSTB(I344705_rst), .Q(I344951) );
nor I_19955 (I344968,I344951,I344804);
nor I_19956 (I344985,I344951,I344866);
nand I_19957 (I344691,I344756,I344985);
nand I_19958 (I345016,I344722,I325967);
nand I_19959 (I345033,I345016,I344951);
and I_19960 (I345050,I345016,I345033);
DFFARX1 I_19961  ( .D(I345050), .CLK(I5694_clk), .RSTB(I344705_rst), .Q(I344673) );
DFFARX1 I_19962  ( .D(I345016), .CLK(I5694_clk), .RSTB(I344705_rst), .Q(I345081) );
and I_19963 (I344670,I344849,I345081);
DFFARX1 I_19964  ( .D(I325997), .CLK(I5694_clk), .RSTB(I344705_rst), .Q(I345112) );
not I_19965 (I345129,I345112);
nor I_19966 (I345146,I344804,I345129);
and I_19967 (I345163,I345112,I345146);
nand I_19968 (I344685,I345112,I344866);
DFFARX1 I_19969  ( .D(I345112), .CLK(I5694_clk), .RSTB(I344705_rst), .Q(I345194) );
not I_19970 (I344682,I345194);
DFFARX1 I_19971  ( .D(I325991), .CLK(I5694_clk), .RSTB(I344705_rst), .Q(I345225) );
not I_19972 (I345242,I345225);
or I_19973 (I345259,I345242,I345163);
DFFARX1 I_19974  ( .D(I345259), .CLK(I5694_clk), .RSTB(I344705_rst), .Q(I344688) );
nand I_19975 (I344697,I345242,I344968);
DFFARX1 I_19976  ( .D(I345242), .CLK(I5694_clk), .RSTB(I344705_rst), .Q(I344667) );
not I_19977 (I345351_rst,I5701);
not I_19978 (I345368,I334399);
nor I_19979 (I345385,I334414,I334429);
nand I_19980 (I345402,I345385,I334417);
DFFARX1 I_19981  ( .D(I345402), .CLK(I5694_clk), .RSTB(I345351_rst), .Q(I345325) );
nor I_19982 (I345433,I345368,I334414);
nand I_19983 (I345450,I345433,I334420);
not I_19984 (I345340,I345450);
DFFARX1 I_19985  ( .D(I345450), .CLK(I5694_clk), .RSTB(I345351_rst), .Q(I345322) );
not I_19986 (I345495,I334414);
not I_19987 (I345512,I345495);
not I_19988 (I345529,I334426);
nor I_19989 (I345546,I345529,I334423);
and I_19990 (I345563,I345546,I334402);
or I_19991 (I345580,I345563,I334411);
DFFARX1 I_19992  ( .D(I345580), .CLK(I5694_clk), .RSTB(I345351_rst), .Q(I345597) );
nor I_19993 (I345614,I345597,I345450);
nor I_19994 (I345631,I345597,I345512);
nand I_19995 (I345337,I345402,I345631);
nand I_19996 (I345662,I345368,I334426);
nand I_19997 (I345679,I345662,I345597);
and I_19998 (I345696,I345662,I345679);
DFFARX1 I_19999  ( .D(I345696), .CLK(I5694_clk), .RSTB(I345351_rst), .Q(I345319) );
DFFARX1 I_20000  ( .D(I345662), .CLK(I5694_clk), .RSTB(I345351_rst), .Q(I345727) );
and I_20001 (I345316,I345495,I345727);
DFFARX1 I_20002  ( .D(I334408), .CLK(I5694_clk), .RSTB(I345351_rst), .Q(I345758) );
not I_20003 (I345775,I345758);
nor I_20004 (I345792,I345450,I345775);
and I_20005 (I345809,I345758,I345792);
nand I_20006 (I345331,I345758,I345512);
DFFARX1 I_20007  ( .D(I345758), .CLK(I5694_clk), .RSTB(I345351_rst), .Q(I345840) );
not I_20008 (I345328,I345840);
DFFARX1 I_20009  ( .D(I334405), .CLK(I5694_clk), .RSTB(I345351_rst), .Q(I345871) );
not I_20010 (I345888,I345871);
or I_20011 (I345905,I345888,I345809);
DFFARX1 I_20012  ( .D(I345905), .CLK(I5694_clk), .RSTB(I345351_rst), .Q(I345334) );
nand I_20013 (I345343,I345888,I345614);
DFFARX1 I_20014  ( .D(I345888), .CLK(I5694_clk), .RSTB(I345351_rst), .Q(I345313) );
not I_20015 (I345997_rst,I5701);
not I_20016 (I346014,I327779);
nor I_20017 (I346031,I327755,I327761);
nand I_20018 (I346048,I346031,I327764);
DFFARX1 I_20019  ( .D(I346048), .CLK(I5694_clk), .RSTB(I345997_rst), .Q(I345971) );
nor I_20020 (I346079,I346014,I327755);
nand I_20021 (I346096,I346079,I327773);
not I_20022 (I345986,I346096);
DFFARX1 I_20023  ( .D(I346096), .CLK(I5694_clk), .RSTB(I345997_rst), .Q(I345968) );
not I_20024 (I346141,I327755);
not I_20025 (I346158,I346141);
not I_20026 (I346175,I327752);
nor I_20027 (I346192,I346175,I327767);
and I_20028 (I346209,I346192,I327758);
or I_20029 (I346226,I346209,I327770);
DFFARX1 I_20030  ( .D(I346226), .CLK(I5694_clk), .RSTB(I345997_rst), .Q(I346243) );
nor I_20031 (I346260,I346243,I346096);
nor I_20032 (I346277,I346243,I346158);
nand I_20033 (I345983,I346048,I346277);
nand I_20034 (I346308,I346014,I327752);
nand I_20035 (I346325,I346308,I346243);
and I_20036 (I346342,I346308,I346325);
DFFARX1 I_20037  ( .D(I346342), .CLK(I5694_clk), .RSTB(I345997_rst), .Q(I345965) );
DFFARX1 I_20038  ( .D(I346308), .CLK(I5694_clk), .RSTB(I345997_rst), .Q(I346373) );
and I_20039 (I345962,I346141,I346373);
DFFARX1 I_20040  ( .D(I327782), .CLK(I5694_clk), .RSTB(I345997_rst), .Q(I346404) );
not I_20041 (I346421,I346404);
nor I_20042 (I346438,I346096,I346421);
and I_20043 (I346455,I346404,I346438);
nand I_20044 (I345977,I346404,I346158);
DFFARX1 I_20045  ( .D(I346404), .CLK(I5694_clk), .RSTB(I345997_rst), .Q(I346486) );
not I_20046 (I345974,I346486);
DFFARX1 I_20047  ( .D(I327776), .CLK(I5694_clk), .RSTB(I345997_rst), .Q(I346517) );
not I_20048 (I346534,I346517);
or I_20049 (I346551,I346534,I346455);
DFFARX1 I_20050  ( .D(I346551), .CLK(I5694_clk), .RSTB(I345997_rst), .Q(I345980) );
nand I_20051 (I345989,I346534,I346260);
DFFARX1 I_20052  ( .D(I346534), .CLK(I5694_clk), .RSTB(I345997_rst), .Q(I345959) );
not I_20053 (I346643_rst,I5701);
not I_20054 (I346660,I326589);
nor I_20055 (I346677,I326565,I326571);
nand I_20056 (I346694,I346677,I326574);
DFFARX1 I_20057  ( .D(I346694), .CLK(I5694_clk), .RSTB(I346643_rst), .Q(I346617) );
nor I_20058 (I346725,I346660,I326565);
nand I_20059 (I346742,I346725,I326583);
not I_20060 (I346632,I346742);
DFFARX1 I_20061  ( .D(I346742), .CLK(I5694_clk), .RSTB(I346643_rst), .Q(I346614) );
not I_20062 (I346787,I326565);
not I_20063 (I346804,I346787);
not I_20064 (I346821,I326562);
nor I_20065 (I346838,I346821,I326577);
and I_20066 (I346855,I346838,I326568);
or I_20067 (I346872,I346855,I326580);
DFFARX1 I_20068  ( .D(I346872), .CLK(I5694_clk), .RSTB(I346643_rst), .Q(I346889) );
nor I_20069 (I346906,I346889,I346742);
nor I_20070 (I346923,I346889,I346804);
nand I_20071 (I346629,I346694,I346923);
nand I_20072 (I346954,I346660,I326562);
nand I_20073 (I346971,I346954,I346889);
and I_20074 (I346988,I346954,I346971);
DFFARX1 I_20075  ( .D(I346988), .CLK(I5694_clk), .RSTB(I346643_rst), .Q(I346611) );
DFFARX1 I_20076  ( .D(I346954), .CLK(I5694_clk), .RSTB(I346643_rst), .Q(I347019) );
and I_20077 (I346608,I346787,I347019);
DFFARX1 I_20078  ( .D(I326592), .CLK(I5694_clk), .RSTB(I346643_rst), .Q(I347050) );
not I_20079 (I347067,I347050);
nor I_20080 (I347084,I346742,I347067);
and I_20081 (I347101,I347050,I347084);
nand I_20082 (I346623,I347050,I346804);
DFFARX1 I_20083  ( .D(I347050), .CLK(I5694_clk), .RSTB(I346643_rst), .Q(I347132) );
not I_20084 (I346620,I347132);
DFFARX1 I_20085  ( .D(I326586), .CLK(I5694_clk), .RSTB(I346643_rst), .Q(I347163) );
not I_20086 (I347180,I347163);
or I_20087 (I347197,I347180,I347101);
DFFARX1 I_20088  ( .D(I347197), .CLK(I5694_clk), .RSTB(I346643_rst), .Q(I346626) );
nand I_20089 (I346635,I347180,I346906);
DFFARX1 I_20090  ( .D(I347180), .CLK(I5694_clk), .RSTB(I346643_rst), .Q(I346605) );
not I_20091 (I347289_rst,I5701);
not I_20092 (I347306,I308327);
nor I_20093 (I347323,I308348,I308321);
nand I_20094 (I347340,I347323,I308336);
DFFARX1 I_20095  ( .D(I347340), .CLK(I5694_clk), .RSTB(I347289_rst), .Q(I347263) );
nor I_20096 (I347371,I347306,I308348);
nand I_20097 (I347388,I347371,I308351);
not I_20098 (I347278,I347388);
DFFARX1 I_20099  ( .D(I347388), .CLK(I5694_clk), .RSTB(I347289_rst), .Q(I347260) );
not I_20100 (I347433,I308348);
not I_20101 (I347450,I347433);
not I_20102 (I347467,I308324);
nor I_20103 (I347484,I347467,I308342);
and I_20104 (I347501,I347484,I308330);
or I_20105 (I347518,I347501,I308333);
DFFARX1 I_20106  ( .D(I347518), .CLK(I5694_clk), .RSTB(I347289_rst), .Q(I347535) );
nor I_20107 (I347552,I347535,I347388);
nor I_20108 (I347569,I347535,I347450);
nand I_20109 (I347275,I347340,I347569);
nand I_20110 (I347600,I347306,I308324);
nand I_20111 (I347617,I347600,I347535);
and I_20112 (I347634,I347600,I347617);
DFFARX1 I_20113  ( .D(I347634), .CLK(I5694_clk), .RSTB(I347289_rst), .Q(I347257) );
DFFARX1 I_20114  ( .D(I347600), .CLK(I5694_clk), .RSTB(I347289_rst), .Q(I347665) );
and I_20115 (I347254,I347433,I347665);
DFFARX1 I_20116  ( .D(I308345), .CLK(I5694_clk), .RSTB(I347289_rst), .Q(I347696) );
not I_20117 (I347713,I347696);
nor I_20118 (I347730,I347388,I347713);
and I_20119 (I347747,I347696,I347730);
nand I_20120 (I347269,I347696,I347450);
DFFARX1 I_20121  ( .D(I347696), .CLK(I5694_clk), .RSTB(I347289_rst), .Q(I347778) );
not I_20122 (I347266,I347778);
DFFARX1 I_20123  ( .D(I308339), .CLK(I5694_clk), .RSTB(I347289_rst), .Q(I347809) );
not I_20124 (I347826,I347809);
or I_20125 (I347843,I347826,I347747);
DFFARX1 I_20126  ( .D(I347843), .CLK(I5694_clk), .RSTB(I347289_rst), .Q(I347272) );
nand I_20127 (I347281,I347826,I347552);
DFFARX1 I_20128  ( .D(I347826), .CLK(I5694_clk), .RSTB(I347289_rst), .Q(I347251) );
not I_20129 (I347935_rst,I5701);
not I_20130 (I347952,I339281);
nor I_20131 (I347969,I339293,I339278);
nand I_20132 (I347986,I347969,I339290);
DFFARX1 I_20133  ( .D(I347986), .CLK(I5694_clk), .RSTB(I347935_rst), .Q(I347909) );
nor I_20134 (I348017,I347952,I339293);
nand I_20135 (I348034,I348017,I339308);
not I_20136 (I347924,I348034);
DFFARX1 I_20137  ( .D(I348034), .CLK(I5694_clk), .RSTB(I347935_rst), .Q(I347906) );
not I_20138 (I348079,I339293);
not I_20139 (I348096,I348079);
not I_20140 (I348113,I339284);
nor I_20141 (I348130,I348113,I339296);
and I_20142 (I348147,I348130,I339287);
or I_20143 (I348164,I348147,I339302);
DFFARX1 I_20144  ( .D(I348164), .CLK(I5694_clk), .RSTB(I347935_rst), .Q(I348181) );
nor I_20145 (I348198,I348181,I348034);
nor I_20146 (I348215,I348181,I348096);
nand I_20147 (I347921,I347986,I348215);
nand I_20148 (I348246,I347952,I339284);
nand I_20149 (I348263,I348246,I348181);
and I_20150 (I348280,I348246,I348263);
DFFARX1 I_20151  ( .D(I348280), .CLK(I5694_clk), .RSTB(I347935_rst), .Q(I347903) );
DFFARX1 I_20152  ( .D(I348246), .CLK(I5694_clk), .RSTB(I347935_rst), .Q(I348311) );
and I_20153 (I347900,I348079,I348311);
DFFARX1 I_20154  ( .D(I339305), .CLK(I5694_clk), .RSTB(I347935_rst), .Q(I348342) );
not I_20155 (I348359,I348342);
nor I_20156 (I348376,I348034,I348359);
and I_20157 (I348393,I348342,I348376);
nand I_20158 (I347915,I348342,I348096);
DFFARX1 I_20159  ( .D(I348342), .CLK(I5694_clk), .RSTB(I347935_rst), .Q(I348424) );
not I_20160 (I347912,I348424);
DFFARX1 I_20161  ( .D(I339299), .CLK(I5694_clk), .RSTB(I347935_rst), .Q(I348455) );
not I_20162 (I348472,I348455);
or I_20163 (I348489,I348472,I348393);
DFFARX1 I_20164  ( .D(I348489), .CLK(I5694_clk), .RSTB(I347935_rst), .Q(I347918) );
nand I_20165 (I347927,I348472,I348198);
DFFARX1 I_20166  ( .D(I348472), .CLK(I5694_clk), .RSTB(I347935_rst), .Q(I347897) );
not I_20167 (I348581_rst,I5701);
not I_20168 (I348598,I307131);
nor I_20169 (I348615,I307161,I307140);
nand I_20170 (I348632,I348615,I307152);
DFFARX1 I_20171  ( .D(I348632), .CLK(I5694_clk), .RSTB(I348581_rst), .Q(I348555) );
nor I_20172 (I348663,I348598,I307161);
nand I_20173 (I348680,I348663,I307134);
not I_20174 (I348570,I348680);
DFFARX1 I_20175  ( .D(I348680), .CLK(I5694_clk), .RSTB(I348581_rst), .Q(I348552) );
not I_20176 (I348725,I307161);
not I_20177 (I348742,I348725);
not I_20178 (I348759,I307137);
nor I_20179 (I348776,I348759,I307155);
and I_20180 (I348793,I348776,I307146);
or I_20181 (I348810,I348793,I307143);
DFFARX1 I_20182  ( .D(I348810), .CLK(I5694_clk), .RSTB(I348581_rst), .Q(I348827) );
nor I_20183 (I348844,I348827,I348680);
nor I_20184 (I348861,I348827,I348742);
nand I_20185 (I348567,I348632,I348861);
nand I_20186 (I348892,I348598,I307137);
nand I_20187 (I348909,I348892,I348827);
and I_20188 (I348926,I348892,I348909);
DFFARX1 I_20189  ( .D(I348926), .CLK(I5694_clk), .RSTB(I348581_rst), .Q(I348549) );
DFFARX1 I_20190  ( .D(I348892), .CLK(I5694_clk), .RSTB(I348581_rst), .Q(I348957) );
and I_20191 (I348546,I348725,I348957);
DFFARX1 I_20192  ( .D(I307149), .CLK(I5694_clk), .RSTB(I348581_rst), .Q(I348988) );
not I_20193 (I349005,I348988);
nor I_20194 (I349022,I348680,I349005);
and I_20195 (I349039,I348988,I349022);
nand I_20196 (I348561,I348988,I348742);
DFFARX1 I_20197  ( .D(I348988), .CLK(I5694_clk), .RSTB(I348581_rst), .Q(I349070) );
not I_20198 (I348558,I349070);
DFFARX1 I_20199  ( .D(I307158), .CLK(I5694_clk), .RSTB(I348581_rst), .Q(I349101) );
not I_20200 (I349118,I349101);
or I_20201 (I349135,I349118,I349039);
DFFARX1 I_20202  ( .D(I349135), .CLK(I5694_clk), .RSTB(I348581_rst), .Q(I348564) );
nand I_20203 (I348573,I349118,I348844);
DFFARX1 I_20204  ( .D(I349118), .CLK(I5694_clk), .RSTB(I348581_rst), .Q(I348543) );
not I_20205 (I349227_rst,I5701);
not I_20206 (I349244,I347266);
nor I_20207 (I349261,I347254,I347278);
nand I_20208 (I349278,I349261,I347263);
DFFARX1 I_20209  ( .D(I349278), .CLK(I5694_clk), .RSTB(I349227_rst), .Q(I349198) );
nor I_20210 (I349309,I349244,I347254);
nand I_20211 (I349326,I349309,I347281);
nand I_20212 (I349343,I349326,I349278);
not I_20213 (I349360,I347254);
not I_20214 (I349377,I347251);
nor I_20215 (I349394,I349377,I347260);
and I_20216 (I349411,I349394,I347275);
or I_20217 (I349428,I349411,I347257);
DFFARX1 I_20218  ( .D(I349428), .CLK(I5694_clk), .RSTB(I349227_rst), .Q(I349445) );
nor I_20219 (I349462,I349445,I349326);
nand I_20220 (I349213,I349360,I349462);
not I_20221 (I349210,I349445);
and I_20222 (I349507,I349445,I349343);
DFFARX1 I_20223  ( .D(I349507), .CLK(I5694_clk), .RSTB(I349227_rst), .Q(I349195) );
DFFARX1 I_20224  ( .D(I349445), .CLK(I5694_clk), .RSTB(I349227_rst), .Q(I349538) );
and I_20225 (I349192,I349360,I349538);
nand I_20226 (I349569,I349244,I347251);
not I_20227 (I349586,I349569);
nor I_20228 (I349603,I349445,I349586);
DFFARX1 I_20229  ( .D(I347272), .CLK(I5694_clk), .RSTB(I349227_rst), .Q(I349620) );
nand I_20230 (I349637,I349620,I349569);
and I_20231 (I349654,I349360,I349637);
DFFARX1 I_20232  ( .D(I349654), .CLK(I5694_clk), .RSTB(I349227_rst), .Q(I349219) );
not I_20233 (I349685,I349620);
nand I_20234 (I349207,I349620,I349603);
nand I_20235 (I349201,I349620,I349586);
DFFARX1 I_20236  ( .D(I347269), .CLK(I5694_clk), .RSTB(I349227_rst), .Q(I349730) );
not I_20237 (I349747,I349730);
nor I_20238 (I349216,I349620,I349747);
nor I_20239 (I349778,I349747,I349685);
and I_20240 (I349795,I349326,I349778);
or I_20241 (I349812,I349569,I349795);
DFFARX1 I_20242  ( .D(I349812), .CLK(I5694_clk), .RSTB(I349227_rst), .Q(I349204) );
DFFARX1 I_20243  ( .D(I349747), .CLK(I5694_clk), .RSTB(I349227_rst), .Q(I349189) );
not I_20244 (I349890_rst,I5701);
not I_20245 (I349907,I330733);
nor I_20246 (I349924,I330748,I330730);
nand I_20247 (I349941,I349924,I330742);
DFFARX1 I_20248  ( .D(I349941), .CLK(I5694_clk), .RSTB(I349890_rst), .Q(I349861) );
nor I_20249 (I349972,I349907,I330748);
nand I_20250 (I349989,I349972,I330739);
nand I_20251 (I350006,I349989,I349941);
not I_20252 (I350023,I330748);
not I_20253 (I350040,I330757);
nor I_20254 (I350057,I350040,I330727);
and I_20255 (I350074,I350057,I330736);
or I_20256 (I350091,I350074,I330754);
DFFARX1 I_20257  ( .D(I350091), .CLK(I5694_clk), .RSTB(I349890_rst), .Q(I350108) );
nor I_20258 (I350125,I350108,I349989);
nand I_20259 (I349876,I350023,I350125);
not I_20260 (I349873,I350108);
and I_20261 (I350170,I350108,I350006);
DFFARX1 I_20262  ( .D(I350170), .CLK(I5694_clk), .RSTB(I349890_rst), .Q(I349858) );
DFFARX1 I_20263  ( .D(I350108), .CLK(I5694_clk), .RSTB(I349890_rst), .Q(I350201) );
and I_20264 (I349855,I350023,I350201);
nand I_20265 (I350232,I349907,I330757);
not I_20266 (I350249,I350232);
nor I_20267 (I350266,I350108,I350249);
DFFARX1 I_20268  ( .D(I330745), .CLK(I5694_clk), .RSTB(I349890_rst), .Q(I350283) );
nand I_20269 (I350300,I350283,I350232);
and I_20270 (I350317,I350023,I350300);
DFFARX1 I_20271  ( .D(I350317), .CLK(I5694_clk), .RSTB(I349890_rst), .Q(I349882) );
not I_20272 (I350348,I350283);
nand I_20273 (I349870,I350283,I350266);
nand I_20274 (I349864,I350283,I350249);
DFFARX1 I_20275  ( .D(I330751), .CLK(I5694_clk), .RSTB(I349890_rst), .Q(I350393) );
not I_20276 (I350410,I350393);
nor I_20277 (I349879,I350283,I350410);
nor I_20278 (I350441,I350410,I350348);
and I_20279 (I350458,I349989,I350441);
or I_20280 (I350475,I350232,I350458);
DFFARX1 I_20281  ( .D(I350475), .CLK(I5694_clk), .RSTB(I349890_rst), .Q(I349867) );
DFFARX1 I_20282  ( .D(I350410), .CLK(I5694_clk), .RSTB(I349890_rst), .Q(I349852) );
not I_20283 (I350553_rst,I5701);
not I_20284 (I350570,I309579);
nor I_20285 (I350587,I309588,I309600);
nand I_20286 (I350604,I350587,I309591);
DFFARX1 I_20287  ( .D(I350604), .CLK(I5694_clk), .RSTB(I350553_rst), .Q(I350524) );
nor I_20288 (I350635,I350570,I309588);
nand I_20289 (I350652,I350635,I309603);
nand I_20290 (I350669,I350652,I350604);
not I_20291 (I350686,I309588);
not I_20292 (I350703,I309609);
nor I_20293 (I350720,I350703,I309585);
and I_20294 (I350737,I350720,I309594);
or I_20295 (I350754,I350737,I309582);
DFFARX1 I_20296  ( .D(I350754), .CLK(I5694_clk), .RSTB(I350553_rst), .Q(I350771) );
nor I_20297 (I350788,I350771,I350652);
nand I_20298 (I350539,I350686,I350788);
not I_20299 (I350536,I350771);
and I_20300 (I350833,I350771,I350669);
DFFARX1 I_20301  ( .D(I350833), .CLK(I5694_clk), .RSTB(I350553_rst), .Q(I350521) );
DFFARX1 I_20302  ( .D(I350771), .CLK(I5694_clk), .RSTB(I350553_rst), .Q(I350864) );
and I_20303 (I350518,I350686,I350864);
nand I_20304 (I350895,I350570,I309609);
not I_20305 (I350912,I350895);
nor I_20306 (I350929,I350771,I350912);
DFFARX1 I_20307  ( .D(I309606), .CLK(I5694_clk), .RSTB(I350553_rst), .Q(I350946) );
nand I_20308 (I350963,I350946,I350895);
and I_20309 (I350980,I350686,I350963);
DFFARX1 I_20310  ( .D(I350980), .CLK(I5694_clk), .RSTB(I350553_rst), .Q(I350545) );
not I_20311 (I351011,I350946);
nand I_20312 (I350533,I350946,I350929);
nand I_20313 (I350527,I350946,I350912);
DFFARX1 I_20314  ( .D(I309597), .CLK(I5694_clk), .RSTB(I350553_rst), .Q(I351056) );
not I_20315 (I351073,I351056);
nor I_20316 (I350542,I350946,I351073);
nor I_20317 (I351104,I351073,I351011);
and I_20318 (I351121,I350652,I351104);
or I_20319 (I351138,I350895,I351121);
DFFARX1 I_20320  ( .D(I351138), .CLK(I5694_clk), .RSTB(I350553_rst), .Q(I350530) );
DFFARX1 I_20321  ( .D(I351073), .CLK(I5694_clk), .RSTB(I350553_rst), .Q(I350515) );
not I_20322 (I351216_rst,I5701);
or I_20323 (I351233,I338122,I338140);
or I_20324 (I351250,I338125,I338122);
DFFARX1 I_20325  ( .D(I351250), .CLK(I5694_clk), .RSTB(I351216_rst), .Q(I351190) );
nor I_20326 (I351281,I338134,I338137);
not I_20327 (I351298,I351281);
not I_20328 (I351315,I338134);
and I_20329 (I351332,I351315,I338143);
nor I_20330 (I351349,I351332,I338140);
nor I_20331 (I351366,I338149,I338128);
DFFARX1 I_20332  ( .D(I351366), .CLK(I5694_clk), .RSTB(I351216_rst), .Q(I351383) );
nand I_20333 (I351400,I351383,I351233);
and I_20334 (I351417,I351349,I351400);
DFFARX1 I_20335  ( .D(I351417), .CLK(I5694_clk), .RSTB(I351216_rst), .Q(I351184) );
nor I_20336 (I351448,I338149,I338125);
DFFARX1 I_20337  ( .D(I351448), .CLK(I5694_clk), .RSTB(I351216_rst), .Q(I351465) );
and I_20338 (I351181,I351281,I351465);
DFFARX1 I_20339  ( .D(I338152), .CLK(I5694_clk), .RSTB(I351216_rst), .Q(I351496) );
and I_20340 (I351513,I351496,I338146);
DFFARX1 I_20341  ( .D(I351513), .CLK(I5694_clk), .RSTB(I351216_rst), .Q(I351530) );
not I_20342 (I351193,I351530);
DFFARX1 I_20343  ( .D(I351513), .CLK(I5694_clk), .RSTB(I351216_rst), .Q(I351178) );
DFFARX1 I_20344  ( .D(I338131), .CLK(I5694_clk), .RSTB(I351216_rst), .Q(I351575) );
not I_20345 (I351592,I351575);
nor I_20346 (I351609,I351250,I351592);
and I_20347 (I351626,I351513,I351609);
or I_20348 (I351643,I351233,I351626);
DFFARX1 I_20349  ( .D(I351643), .CLK(I5694_clk), .RSTB(I351216_rst), .Q(I351199) );
nor I_20350 (I351674,I351575,I351383);
nand I_20351 (I351208,I351349,I351674);
nor I_20352 (I351705,I351575,I351298);
nand I_20353 (I351202,I351448,I351705);
not I_20354 (I351205,I351575);
nand I_20355 (I351196,I351575,I351298);
DFFARX1 I_20356  ( .D(I351575), .CLK(I5694_clk), .RSTB(I351216_rst), .Q(I351187) );
not I_20357 (I351811_rst,I5701);
or I_20358 (I351828,I315546,I315561);
or I_20359 (I351845,I315549,I315546);
DFFARX1 I_20360  ( .D(I351845), .CLK(I5694_clk), .RSTB(I351811_rst), .Q(I351785) );
nor I_20361 (I351876,I315552,I315567);
not I_20362 (I351893,I351876);
not I_20363 (I351910,I315552);
and I_20364 (I351927,I351910,I315555);
nor I_20365 (I351944,I351927,I315561);
nor I_20366 (I351961,I315558,I315576);
DFFARX1 I_20367  ( .D(I351961), .CLK(I5694_clk), .RSTB(I351811_rst), .Q(I351978) );
nand I_20368 (I351995,I351978,I351828);
and I_20369 (I352012,I351944,I351995);
DFFARX1 I_20370  ( .D(I352012), .CLK(I5694_clk), .RSTB(I351811_rst), .Q(I351779) );
nor I_20371 (I352043,I315558,I315549);
DFFARX1 I_20372  ( .D(I352043), .CLK(I5694_clk), .RSTB(I351811_rst), .Q(I352060) );
and I_20373 (I351776,I351876,I352060);
DFFARX1 I_20374  ( .D(I315573), .CLK(I5694_clk), .RSTB(I351811_rst), .Q(I352091) );
and I_20375 (I352108,I352091,I315564);
DFFARX1 I_20376  ( .D(I352108), .CLK(I5694_clk), .RSTB(I351811_rst), .Q(I352125) );
not I_20377 (I351788,I352125);
DFFARX1 I_20378  ( .D(I352108), .CLK(I5694_clk), .RSTB(I351811_rst), .Q(I351773) );
DFFARX1 I_20379  ( .D(I315570), .CLK(I5694_clk), .RSTB(I351811_rst), .Q(I352170) );
not I_20380 (I352187,I352170);
nor I_20381 (I352204,I351845,I352187);
and I_20382 (I352221,I352108,I352204);
or I_20383 (I352238,I351828,I352221);
DFFARX1 I_20384  ( .D(I352238), .CLK(I5694_clk), .RSTB(I351811_rst), .Q(I351794) );
nor I_20385 (I352269,I352170,I351978);
nand I_20386 (I351803,I351944,I352269);
nor I_20387 (I352300,I352170,I351893);
nand I_20388 (I351797,I352043,I352300);
not I_20389 (I351800,I352170);
nand I_20390 (I351791,I352170,I351893);
DFFARX1 I_20391  ( .D(I352170), .CLK(I5694_clk), .RSTB(I351811_rst), .Q(I351782) );
not I_20392 (I352406_rst,I5701);
or I_20393 (I352423,I343396,I343390);
or I_20394 (I352440,I343384,I343396);
DFFARX1 I_20395  ( .D(I352440), .CLK(I5694_clk), .RSTB(I352406_rst), .Q(I352380) );
nor I_20396 (I352471,I343402,I343393);
not I_20397 (I352488,I352471);
not I_20398 (I352505,I343402);
and I_20399 (I352522,I352505,I343399);
nor I_20400 (I352539,I352522,I343390);
nor I_20401 (I352556,I343375,I343381);
DFFARX1 I_20402  ( .D(I352556), .CLK(I5694_clk), .RSTB(I352406_rst), .Q(I352573) );
nand I_20403 (I352590,I352573,I352423);
and I_20404 (I352607,I352539,I352590);
DFFARX1 I_20405  ( .D(I352607), .CLK(I5694_clk), .RSTB(I352406_rst), .Q(I352374) );
nor I_20406 (I352638,I343375,I343384);
DFFARX1 I_20407  ( .D(I352638), .CLK(I5694_clk), .RSTB(I352406_rst), .Q(I352655) );
and I_20408 (I352371,I352471,I352655);
DFFARX1 I_20409  ( .D(I343387), .CLK(I5694_clk), .RSTB(I352406_rst), .Q(I352686) );
and I_20410 (I352703,I352686,I343405);
DFFARX1 I_20411  ( .D(I352703), .CLK(I5694_clk), .RSTB(I352406_rst), .Q(I352720) );
not I_20412 (I352383,I352720);
DFFARX1 I_20413  ( .D(I352703), .CLK(I5694_clk), .RSTB(I352406_rst), .Q(I352368) );
DFFARX1 I_20414  ( .D(I343378), .CLK(I5694_clk), .RSTB(I352406_rst), .Q(I352765) );
not I_20415 (I352782,I352765);
nor I_20416 (I352799,I352440,I352782);
and I_20417 (I352816,I352703,I352799);
or I_20418 (I352833,I352423,I352816);
DFFARX1 I_20419  ( .D(I352833), .CLK(I5694_clk), .RSTB(I352406_rst), .Q(I352389) );
nor I_20420 (I352864,I352765,I352573);
nand I_20421 (I352398,I352539,I352864);
nor I_20422 (I352895,I352765,I352488);
nand I_20423 (I352392,I352638,I352895);
not I_20424 (I352395,I352765);
nand I_20425 (I352386,I352765,I352488);
DFFARX1 I_20426  ( .D(I352765), .CLK(I5694_clk), .RSTB(I352406_rst), .Q(I352377) );
not I_20427 (I353001_rst,I5701);
not I_20428 (I353018,I331935);
nor I_20429 (I353035,I331932,I331923);
nand I_20430 (I353052,I353035,I331926);
nor I_20431 (I353069,I353018,I331932);
nand I_20432 (I353086,I353069,I331920);
not I_20433 (I353103,I353086);
not I_20434 (I353120,I331932);
nor I_20435 (I352990,I353086,I353120);
not I_20436 (I353151,I353120);
nand I_20437 (I352975,I353086,I353151);
not I_20438 (I353182,I331941);
nor I_20439 (I353199,I353182,I331944);
and I_20440 (I353216,I353199,I331929);
or I_20441 (I353233,I353216,I331917);
DFFARX1 I_20442  ( .D(I353233), .CLK(I5694_clk), .RSTB(I353001_rst), .Q(I353250) );
nor I_20443 (I353267,I353250,I353103);
DFFARX1 I_20444  ( .D(I353250), .CLK(I5694_clk), .RSTB(I353001_rst), .Q(I353284) );
not I_20445 (I352972,I353284);
nand I_20446 (I353315,I353018,I331941);
and I_20447 (I353332,I353315,I353267);
DFFARX1 I_20448  ( .D(I353315), .CLK(I5694_clk), .RSTB(I353001_rst), .Q(I352969) );
DFFARX1 I_20449  ( .D(I331938), .CLK(I5694_clk), .RSTB(I353001_rst), .Q(I353363) );
nor I_20450 (I353380,I353363,I353086);
nand I_20451 (I352987,I353250,I353380);
nor I_20452 (I353411,I353363,I353151);
not I_20453 (I352984,I353363);
nand I_20454 (I353442,I353363,I353052);
and I_20455 (I353459,I353120,I353442);
DFFARX1 I_20456  ( .D(I353459), .CLK(I5694_clk), .RSTB(I353001_rst), .Q(I352963) );
DFFARX1 I_20457  ( .D(I353363), .CLK(I5694_clk), .RSTB(I353001_rst), .Q(I352966) );
DFFARX1 I_20458  ( .D(I331947), .CLK(I5694_clk), .RSTB(I353001_rst), .Q(I353504) );
not I_20459 (I353521,I353504);
nand I_20460 (I353538,I353521,I353086);
and I_20461 (I353555,I353315,I353538);
DFFARX1 I_20462  ( .D(I353555), .CLK(I5694_clk), .RSTB(I353001_rst), .Q(I352993) );
or I_20463 (I353586,I353521,I353332);
DFFARX1 I_20464  ( .D(I353586), .CLK(I5694_clk), .RSTB(I353001_rst), .Q(I352978) );
nand I_20465 (I352981,I353521,I353411);
not I_20466 (I353664_rst,I5701);
not I_20467 (I353681,I323092);
nor I_20468 (I353698,I323104,I323086);
nand I_20469 (I353715,I353698,I323107);
nor I_20470 (I353732,I353681,I323104);
nand I_20471 (I353749,I353732,I323098);
not I_20472 (I353766,I353749);
not I_20473 (I353783,I323104);
nor I_20474 (I353653,I353749,I353783);
not I_20475 (I353814,I353783);
nand I_20476 (I353638,I353749,I353814);
not I_20477 (I353845,I323089);
nor I_20478 (I353862,I353845,I323083);
and I_20479 (I353879,I353862,I323095);
or I_20480 (I353896,I353879,I323080);
DFFARX1 I_20481  ( .D(I353896), .CLK(I5694_clk), .RSTB(I353664_rst), .Q(I353913) );
nor I_20482 (I353930,I353913,I353766);
DFFARX1 I_20483  ( .D(I353913), .CLK(I5694_clk), .RSTB(I353664_rst), .Q(I353947) );
not I_20484 (I353635,I353947);
nand I_20485 (I353978,I353681,I323089);
and I_20486 (I353995,I353978,I353930);
DFFARX1 I_20487  ( .D(I353978), .CLK(I5694_clk), .RSTB(I353664_rst), .Q(I353632) );
DFFARX1 I_20488  ( .D(I323077), .CLK(I5694_clk), .RSTB(I353664_rst), .Q(I354026) );
nor I_20489 (I354043,I354026,I353749);
nand I_20490 (I353650,I353913,I354043);
nor I_20491 (I354074,I354026,I353814);
not I_20492 (I353647,I354026);
nand I_20493 (I354105,I354026,I353715);
and I_20494 (I354122,I353783,I354105);
DFFARX1 I_20495  ( .D(I354122), .CLK(I5694_clk), .RSTB(I353664_rst), .Q(I353626) );
DFFARX1 I_20496  ( .D(I354026), .CLK(I5694_clk), .RSTB(I353664_rst), .Q(I353629) );
DFFARX1 I_20497  ( .D(I323101), .CLK(I5694_clk), .RSTB(I353664_rst), .Q(I354167) );
not I_20498 (I354184,I354167);
nand I_20499 (I354201,I354184,I353749);
and I_20500 (I354218,I353978,I354201);
DFFARX1 I_20501  ( .D(I354218), .CLK(I5694_clk), .RSTB(I353664_rst), .Q(I353656) );
or I_20502 (I354249,I354184,I353995);
DFFARX1 I_20503  ( .D(I354249), .CLK(I5694_clk), .RSTB(I353664_rst), .Q(I353641) );
nand I_20504 (I353644,I354184,I354074);
not I_20505 (I354327_rst,I5701);
not I_20506 (I354344,I351791);
nor I_20507 (I354361,I351785,I351776);
nand I_20508 (I354378,I354361,I351788);
nor I_20509 (I354395,I354344,I351785);
nand I_20510 (I354412,I354395,I351803);
not I_20511 (I354429,I354412);
not I_20512 (I354446,I351785);
nor I_20513 (I354316,I354412,I354446);
not I_20514 (I354477,I354446);
nand I_20515 (I354301,I354412,I354477);
not I_20516 (I354508,I351779);
nor I_20517 (I354525,I354508,I351773);
and I_20518 (I354542,I354525,I351800);
or I_20519 (I354559,I354542,I351797);
DFFARX1 I_20520  ( .D(I354559), .CLK(I5694_clk), .RSTB(I354327_rst), .Q(I354576) );
nor I_20521 (I354593,I354576,I354429);
DFFARX1 I_20522  ( .D(I354576), .CLK(I5694_clk), .RSTB(I354327_rst), .Q(I354610) );
not I_20523 (I354298,I354610);
nand I_20524 (I354641,I354344,I351779);
and I_20525 (I354658,I354641,I354593);
DFFARX1 I_20526  ( .D(I354641), .CLK(I5694_clk), .RSTB(I354327_rst), .Q(I354295) );
DFFARX1 I_20527  ( .D(I351794), .CLK(I5694_clk), .RSTB(I354327_rst), .Q(I354689) );
nor I_20528 (I354706,I354689,I354412);
nand I_20529 (I354313,I354576,I354706);
nor I_20530 (I354737,I354689,I354477);
not I_20531 (I354310,I354689);
nand I_20532 (I354768,I354689,I354378);
and I_20533 (I354785,I354446,I354768);
DFFARX1 I_20534  ( .D(I354785), .CLK(I5694_clk), .RSTB(I354327_rst), .Q(I354289) );
DFFARX1 I_20535  ( .D(I354689), .CLK(I5694_clk), .RSTB(I354327_rst), .Q(I354292) );
DFFARX1 I_20536  ( .D(I351782), .CLK(I5694_clk), .RSTB(I354327_rst), .Q(I354830) );
not I_20537 (I354847,I354830);
nand I_20538 (I354864,I354847,I354412);
and I_20539 (I354881,I354641,I354864);
DFFARX1 I_20540  ( .D(I354881), .CLK(I5694_clk), .RSTB(I354327_rst), .Q(I354319) );
or I_20541 (I354912,I354847,I354658);
DFFARX1 I_20542  ( .D(I354912), .CLK(I5694_clk), .RSTB(I354327_rst), .Q(I354304) );
nand I_20543 (I354307,I354847,I354737);
not I_20544 (I354990_rst,I5701);
not I_20545 (I355007,I318159);
nor I_20546 (I355024,I318156,I318174);
nand I_20547 (I355041,I355024,I318177);
nor I_20548 (I355058,I355007,I318156);
nand I_20549 (I355075,I355058,I318162);
not I_20550 (I355092,I355075);
not I_20551 (I355109,I318156);
nor I_20552 (I354979,I355075,I355109);
not I_20553 (I355140,I355109);
nand I_20554 (I354964,I355075,I355140);
not I_20555 (I355171,I318171);
nor I_20556 (I355188,I355171,I318153);
and I_20557 (I355205,I355188,I318147);
or I_20558 (I355222,I355205,I318165);
DFFARX1 I_20559  ( .D(I355222), .CLK(I5694_clk), .RSTB(I354990_rst), .Q(I355239) );
nor I_20560 (I355256,I355239,I355092);
DFFARX1 I_20561  ( .D(I355239), .CLK(I5694_clk), .RSTB(I354990_rst), .Q(I355273) );
not I_20562 (I354961,I355273);
nand I_20563 (I355304,I355007,I318171);
and I_20564 (I355321,I355304,I355256);
DFFARX1 I_20565  ( .D(I355304), .CLK(I5694_clk), .RSTB(I354990_rst), .Q(I354958) );
DFFARX1 I_20566  ( .D(I318150), .CLK(I5694_clk), .RSTB(I354990_rst), .Q(I355352) );
nor I_20567 (I355369,I355352,I355075);
nand I_20568 (I354976,I355239,I355369);
nor I_20569 (I355400,I355352,I355140);
not I_20570 (I354973,I355352);
nand I_20571 (I355431,I355352,I355041);
and I_20572 (I355448,I355109,I355431);
DFFARX1 I_20573  ( .D(I355448), .CLK(I5694_clk), .RSTB(I354990_rst), .Q(I354952) );
DFFARX1 I_20574  ( .D(I355352), .CLK(I5694_clk), .RSTB(I354990_rst), .Q(I354955) );
DFFARX1 I_20575  ( .D(I318168), .CLK(I5694_clk), .RSTB(I354990_rst), .Q(I355493) );
not I_20576 (I355510,I355493);
nand I_20577 (I355527,I355510,I355075);
and I_20578 (I355544,I355304,I355527);
DFFARX1 I_20579  ( .D(I355544), .CLK(I5694_clk), .RSTB(I354990_rst), .Q(I354982) );
or I_20580 (I355575,I355510,I355321);
DFFARX1 I_20581  ( .D(I355575), .CLK(I5694_clk), .RSTB(I354990_rst), .Q(I354967) );
nand I_20582 (I354970,I355510,I355400);
not I_20583 (I355653_rst,I5701);
not I_20584 (I355670,I321936);
nor I_20585 (I355687,I321948,I321930);
nand I_20586 (I355704,I355687,I321951);
nor I_20587 (I355721,I355670,I321948);
nand I_20588 (I355738,I355721,I321942);
not I_20589 (I355755,I355738);
not I_20590 (I355772,I321948);
nor I_20591 (I355642,I355738,I355772);
not I_20592 (I355803,I355772);
nand I_20593 (I355627,I355738,I355803);
not I_20594 (I355834,I321933);
nor I_20595 (I355851,I355834,I321927);
and I_20596 (I355868,I355851,I321939);
or I_20597 (I355885,I355868,I321924);
DFFARX1 I_20598  ( .D(I355885), .CLK(I5694_clk), .RSTB(I355653_rst), .Q(I355902) );
nor I_20599 (I355919,I355902,I355755);
DFFARX1 I_20600  ( .D(I355902), .CLK(I5694_clk), .RSTB(I355653_rst), .Q(I355936) );
not I_20601 (I355624,I355936);
nand I_20602 (I355967,I355670,I321933);
and I_20603 (I355984,I355967,I355919);
DFFARX1 I_20604  ( .D(I355967), .CLK(I5694_clk), .RSTB(I355653_rst), .Q(I355621) );
DFFARX1 I_20605  ( .D(I321921), .CLK(I5694_clk), .RSTB(I355653_rst), .Q(I356015) );
nor I_20606 (I356032,I356015,I355738);
nand I_20607 (I355639,I355902,I356032);
nor I_20608 (I356063,I356015,I355803);
not I_20609 (I355636,I356015);
nand I_20610 (I356094,I356015,I355704);
and I_20611 (I35611_rst1,I355772,I356094);
DFFARX1 I_20612  ( .D(I35611_rst1), .CLK(I5694_clk), .RSTB(I355653_rst), .Q(I355615) );
DFFARX1 I_20613  ( .D(I356015), .CLK(I5694_clk), .RSTB(I355653_rst), .Q(I355618) );
DFFARX1 I_20614  ( .D(I321945), .CLK(I5694_clk), .RSTB(I355653_rst), .Q(I356156) );
not I_20615 (I356173,I356156);
nand I_20616 (I356190,I356173,I355738);
and I_20617 (I356207,I355967,I356190);
DFFARX1 I_20618  ( .D(I356207), .CLK(I5694_clk), .RSTB(I355653_rst), .Q(I355645) );
or I_20619 (I356238,I356173,I355984);
DFFARX1 I_20620  ( .D(I356238), .CLK(I5694_clk), .RSTB(I355653_rst), .Q(I355630) );
nand I_20621 (I355633,I356173,I356063);
not I_20622 (I356316_rst,I5701);
not I_20623 (I356333,I351196);
nor I_20624 (I356350,I351190,I351181);
nand I_20625 (I356367,I356350,I351193);
nor I_20626 (I356384,I356333,I351190);
nand I_20627 (I356401,I356384,I351208);
not I_20628 (I356418,I356401);
not I_20629 (I356435,I351190);
nor I_20630 (I356305,I356401,I356435);
not I_20631 (I356466,I356435);
nand I_20632 (I356290,I356401,I356466);
not I_20633 (I356497,I351184);
nor I_20634 (I356514,I356497,I351178);
and I_20635 (I356531,I356514,I351205);
or I_20636 (I356548,I356531,I351202);
DFFARX1 I_20637  ( .D(I356548), .CLK(I5694_clk), .RSTB(I356316_rst), .Q(I356565) );
nor I_20638 (I356582,I356565,I356418);
DFFARX1 I_20639  ( .D(I356565), .CLK(I5694_clk), .RSTB(I356316_rst), .Q(I356599) );
not I_20640 (I356287,I356599);
nand I_20641 (I356630,I356333,I351184);
and I_20642 (I356647,I356630,I356582);
DFFARX1 I_20643  ( .D(I356630), .CLK(I5694_clk), .RSTB(I356316_rst), .Q(I356284) );
DFFARX1 I_20644  ( .D(I351199), .CLK(I5694_clk), .RSTB(I356316_rst), .Q(I356678) );
nor I_20645 (I356695,I356678,I356401);
nand I_20646 (I356302,I356565,I356695);
nor I_20647 (I356726,I356678,I356466);
not I_20648 (I356299,I356678);
nand I_20649 (I356757,I356678,I356367);
and I_20650 (I356774,I356435,I356757);
DFFARX1 I_20651  ( .D(I356774), .CLK(I5694_clk), .RSTB(I356316_rst), .Q(I356278) );
DFFARX1 I_20652  ( .D(I356678), .CLK(I5694_clk), .RSTB(I356316_rst), .Q(I356281) );
DFFARX1 I_20653  ( .D(I351187), .CLK(I5694_clk), .RSTB(I356316_rst), .Q(I356819) );
not I_20654 (I356836,I356819);
nand I_20655 (I356853,I356836,I356401);
and I_20656 (I356870,I356630,I356853);
DFFARX1 I_20657  ( .D(I356870), .CLK(I5694_clk), .RSTB(I356316_rst), .Q(I356308) );
or I_20658 (I356901,I356836,I356647);
DFFARX1 I_20659  ( .D(I356901), .CLK(I5694_clk), .RSTB(I356316_rst), .Q(I356293) );
nand I_20660 (I356296,I356836,I356726);
not I_20661 (I356979_rst,I5701);
not I_20662 (I356996,I329555);
nor I_20663 (I357013,I329564,I329546);
nand I_20664 (I357030,I357013,I329567);
nor I_20665 (I357047,I356996,I329564);
nand I_20666 (I357064,I357047,I329558);
not I_20667 (I357081,I357064);
not I_20668 (I357098,I329564);
nor I_20669 (I356968,I357064,I357098);
not I_20670 (I357129,I357098);
nand I_20671 (I356953,I357064,I357129);
not I_20672 (I357160,I329552);
nor I_20673 (I357177,I357160,I329543);
and I_20674 (I357194,I357177,I329540);
or I_20675 (I357211,I357194,I329537);
DFFARX1 I_20676  ( .D(I357211), .CLK(I5694_clk), .RSTB(I356979_rst), .Q(I357228) );
nor I_20677 (I357245,I357228,I357081);
DFFARX1 I_20678  ( .D(I357228), .CLK(I5694_clk), .RSTB(I356979_rst), .Q(I357262) );
not I_20679 (I356950,I357262);
nand I_20680 (I357293,I356996,I329552);
and I_20681 (I357310,I357293,I357245);
DFFARX1 I_20682  ( .D(I357293), .CLK(I5694_clk), .RSTB(I356979_rst), .Q(I356947) );
DFFARX1 I_20683  ( .D(I329561), .CLK(I5694_clk), .RSTB(I356979_rst), .Q(I357341) );
nor I_20684 (I357358,I357341,I357064);
nand I_20685 (I356965,I357228,I357358);
nor I_20686 (I357389,I357341,I357129);
not I_20687 (I356962,I357341);
nand I_20688 (I357420,I357341,I357030);
and I_20689 (I357437,I357098,I357420);
DFFARX1 I_20690  ( .D(I357437), .CLK(I5694_clk), .RSTB(I356979_rst), .Q(I356941) );
DFFARX1 I_20691  ( .D(I357341), .CLK(I5694_clk), .RSTB(I356979_rst), .Q(I356944) );
DFFARX1 I_20692  ( .D(I329549), .CLK(I5694_clk), .RSTB(I356979_rst), .Q(I357482) );
not I_20693 (I357499,I357482);
nand I_20694 (I357516,I357499,I357064);
and I_20695 (I357533,I357293,I357516);
DFFARX1 I_20696  ( .D(I357533), .CLK(I5694_clk), .RSTB(I356979_rst), .Q(I356971) );
or I_20697 (I357564,I357499,I357310);
DFFARX1 I_20698  ( .D(I357564), .CLK(I5694_clk), .RSTB(I356979_rst), .Q(I356956) );
nand I_20699 (I356959,I357499,I357389);
not I_20700 (I357642_rst,I5701);
not I_20701 (I357659,I323670);
nor I_20702 (I357676,I323682,I323664);
nand I_20703 (I357693,I357676,I323685);
nor I_20704 (I357710,I357659,I323682);
nand I_20705 (I357727,I357710,I323676);
not I_20706 (I357744,I357727);
not I_20707 (I357761,I323682);
nor I_20708 (I357631,I357727,I357761);
not I_20709 (I357792,I357761);
nand I_20710 (I357616,I357727,I357792);
not I_20711 (I357823,I323667);
nor I_20712 (I357840,I357823,I323661);
and I_20713 (I357857,I357840,I323673);
or I_20714 (I357874,I357857,I323658);
DFFARX1 I_20715  ( .D(I357874), .CLK(I5694_clk), .RSTB(I357642_rst), .Q(I357891) );
nor I_20716 (I357908,I357891,I357744);
DFFARX1 I_20717  ( .D(I357891), .CLK(I5694_clk), .RSTB(I357642_rst), .Q(I357925) );
not I_20718 (I357613,I357925);
nand I_20719 (I357956,I357659,I323667);
and I_20720 (I357973,I357956,I357908);
DFFARX1 I_20721  ( .D(I357956), .CLK(I5694_clk), .RSTB(I357642_rst), .Q(I357610) );
DFFARX1 I_20722  ( .D(I323655), .CLK(I5694_clk), .RSTB(I357642_rst), .Q(I358004) );
nor I_20723 (I358021,I358004,I357727);
nand I_20724 (I357628,I357891,I358021);
nor I_20725 (I358052,I358004,I357792);
not I_20726 (I357625,I358004);
nand I_20727 (I358083,I358004,I357693);
and I_20728 (I358100,I357761,I358083);
DFFARX1 I_20729  ( .D(I358100), .CLK(I5694_clk), .RSTB(I357642_rst), .Q(I357604) );
DFFARX1 I_20730  ( .D(I358004), .CLK(I5694_clk), .RSTB(I357642_rst), .Q(I357607) );
DFFARX1 I_20731  ( .D(I323679), .CLK(I5694_clk), .RSTB(I357642_rst), .Q(I358145) );
not I_20732 (I358162,I358145);
nand I_20733 (I358179,I358162,I357727);
and I_20734 (I358196,I357956,I358179);
DFFARX1 I_20735  ( .D(I358196), .CLK(I5694_clk), .RSTB(I357642_rst), .Q(I357634) );
or I_20736 (I358227,I358162,I357973);
DFFARX1 I_20737  ( .D(I358227), .CLK(I5694_clk), .RSTB(I357642_rst), .Q(I357619) );
nand I_20738 (I357622,I358162,I358052);
not I_20739 (I358305_rst,I5701);
not I_20740 (I358322,I328960);
nor I_20741 (I358339,I328969,I328951);
nand I_20742 (I358356,I358339,I328972);
nor I_20743 (I358373,I358322,I328969);
nand I_20744 (I358390,I358373,I328963);
not I_20745 (I358407,I358390);
not I_20746 (I358424,I328969);
nor I_20747 (I358294,I358390,I358424);
not I_20748 (I358455,I358424);
nand I_20749 (I358279,I358390,I358455);
not I_20750 (I358486,I328957);
nor I_20751 (I358503,I358486,I328948);
and I_20752 (I358520,I358503,I328945);
or I_20753 (I358537,I358520,I328942);
DFFARX1 I_20754  ( .D(I358537), .CLK(I5694_clk), .RSTB(I358305_rst), .Q(I358554) );
nor I_20755 (I358571,I358554,I358407);
DFFARX1 I_20756  ( .D(I358554), .CLK(I5694_clk), .RSTB(I358305_rst), .Q(I358588) );
not I_20757 (I358276,I358588);
nand I_20758 (I358619,I358322,I328957);
and I_20759 (I358636,I358619,I358571);
DFFARX1 I_20760  ( .D(I358619), .CLK(I5694_clk), .RSTB(I358305_rst), .Q(I358273) );
DFFARX1 I_20761  ( .D(I328966), .CLK(I5694_clk), .RSTB(I358305_rst), .Q(I358667) );
nor I_20762 (I358684,I358667,I358390);
nand I_20763 (I358291,I358554,I358684);
nor I_20764 (I358715,I358667,I358455);
not I_20765 (I358288,I358667);
nand I_20766 (I358746,I358667,I358356);
and I_20767 (I358763,I358424,I358746);
DFFARX1 I_20768  ( .D(I358763), .CLK(I5694_clk), .RSTB(I358305_rst), .Q(I358267) );
DFFARX1 I_20769  ( .D(I358667), .CLK(I5694_clk), .RSTB(I358305_rst), .Q(I358270) );
DFFARX1 I_20770  ( .D(I328954), .CLK(I5694_clk), .RSTB(I358305_rst), .Q(I358808) );
not I_20771 (I358825,I358808);
nand I_20772 (I358842,I358825,I358390);
and I_20773 (I358859,I358619,I358842);
DFFARX1 I_20774  ( .D(I358859), .CLK(I5694_clk), .RSTB(I358305_rst), .Q(I358297) );
or I_20775 (I358890,I358825,I358636);
DFFARX1 I_20776  ( .D(I358890), .CLK(I5694_clk), .RSTB(I358305_rst), .Q(I358282) );
nand I_20777 (I358285,I358825,I358715);
not I_20778 (I358968_rst,I5701);
not I_20779 (I358985,I335663);
nor I_20780 (I359002,I335681,I335672);
nand I_20781 (I359019,I359002,I335678);
nor I_20782 (I359036,I358985,I335681);
nand I_20783 (I359053,I359036,I335684);
not I_20784 (I359070,I359053);
not I_20785 (I359087,I335681);
nor I_20786 (I358957,I359053,I359087);
not I_20787 (I359118,I359087);
nand I_20788 (I358942,I359053,I359118);
not I_20789 (I359149,I335660);
nor I_20790 (I359166,I359149,I335675);
and I_20791 (I359183,I359166,I335657);
or I_20792 (I359200,I359183,I335666);
DFFARX1 I_20793  ( .D(I359200), .CLK(I5694_clk), .RSTB(I358968_rst), .Q(I359217) );
nor I_20794 (I359234,I359217,I359070);
DFFARX1 I_20795  ( .D(I359217), .CLK(I5694_clk), .RSTB(I358968_rst), .Q(I359251) );
not I_20796 (I358939,I359251);
nand I_20797 (I359282,I358985,I335660);
and I_20798 (I359299,I359282,I359234);
DFFARX1 I_20799  ( .D(I359282), .CLK(I5694_clk), .RSTB(I358968_rst), .Q(I358936) );
DFFARX1 I_20800  ( .D(I335669), .CLK(I5694_clk), .RSTB(I358968_rst), .Q(I359330) );
nor I_20801 (I359347,I359330,I359053);
nand I_20802 (I358954,I359217,I359347);
nor I_20803 (I359378,I359330,I359118);
not I_20804 (I358951,I359330);
nand I_20805 (I359409,I359330,I359019);
and I_20806 (I359426,I359087,I359409);
DFFARX1 I_20807  ( .D(I359426), .CLK(I5694_clk), .RSTB(I358968_rst), .Q(I358930) );
DFFARX1 I_20808  ( .D(I359330), .CLK(I5694_clk), .RSTB(I358968_rst), .Q(I358933) );
DFFARX1 I_20809  ( .D(I335687), .CLK(I5694_clk), .RSTB(I358968_rst), .Q(I359471) );
not I_20810 (I359488,I359471);
nand I_20811 (I359505,I359488,I359053);
and I_20812 (I359522,I359282,I359505);
DFFARX1 I_20813  ( .D(I359522), .CLK(I5694_clk), .RSTB(I358968_rst), .Q(I358960) );
or I_20814 (I359553,I359488,I359299);
DFFARX1 I_20815  ( .D(I359553), .CLK(I5694_clk), .RSTB(I358968_rst), .Q(I358945) );
nand I_20816 (I358948,I359488,I359378);
not I_20817 (I359631_rst,I5701);
not I_20818 (I359648,I345965);
nor I_20819 (I359665,I345962,I345986);
nand I_20820 (I359682,I359665,I345983);
nor I_20821 (I359699,I359648,I345962);
nand I_20822 (I359716,I359699,I345989);
not I_20823 (I359733,I359716);
not I_20824 (I359750,I345962);
nor I_20825 (I359620,I359716,I359750);
not I_20826 (I359781,I359750);
nand I_20827 (I359605,I359716,I359781);
not I_20828 (I359812,I345980);
nor I_20829 (I359829,I359812,I345971);
and I_20830 (I359846,I359829,I345968);
or I_20831 (I359863,I359846,I345977);
DFFARX1 I_20832  ( .D(I359863), .CLK(I5694_clk), .RSTB(I359631_rst), .Q(I359880) );
nor I_20833 (I359897,I359880,I359733);
DFFARX1 I_20834  ( .D(I359880), .CLK(I5694_clk), .RSTB(I359631_rst), .Q(I359914) );
not I_20835 (I359602,I359914);
nand I_20836 (I359945,I359648,I345980);
and I_20837 (I359962,I359945,I359897);
DFFARX1 I_20838  ( .D(I359945), .CLK(I5694_clk), .RSTB(I359631_rst), .Q(I359599) );
DFFARX1 I_20839  ( .D(I345959), .CLK(I5694_clk), .RSTB(I359631_rst), .Q(I359993) );
nor I_20840 (I360010,I359993,I359716);
nand I_20841 (I359617,I359880,I360010);
nor I_20842 (I360041,I359993,I359781);
not I_20843 (I359614,I359993);
nand I_20844 (I360072,I359993,I359682);
and I_20845 (I360089,I359750,I360072);
DFFARX1 I_20846  ( .D(I360089), .CLK(I5694_clk), .RSTB(I359631_rst), .Q(I359593) );
DFFARX1 I_20847  ( .D(I359993), .CLK(I5694_clk), .RSTB(I359631_rst), .Q(I359596) );
DFFARX1 I_20848  ( .D(I345974), .CLK(I5694_clk), .RSTB(I359631_rst), .Q(I360134) );
not I_20849 (I360151,I360134);
nand I_20850 (I360168,I360151,I359716);
and I_20851 (I360185,I359945,I360168);
DFFARX1 I_20852  ( .D(I360185), .CLK(I5694_clk), .RSTB(I359631_rst), .Q(I359623) );
or I_20853 (I360216,I360151,I359962);
DFFARX1 I_20854  ( .D(I360216), .CLK(I5694_clk), .RSTB(I359631_rst), .Q(I359608) );
nand I_20855 (I359611,I360151,I360041);
not I_20856 (I360294_rst,I5701);
not I_20857 (I360311,I328365);
nor I_20858 (I360328,I328374,I328356);
nand I_20859 (I360345,I360328,I328377);
nor I_20860 (I360362,I360311,I328374);
nand I_20861 (I360379,I360362,I328368);
not I_20862 (I360396,I360379);
not I_20863 (I360413,I328374);
nor I_20864 (I360283,I360379,I360413);
not I_20865 (I360444,I360413);
nand I_20866 (I360268,I360379,I360444);
not I_20867 (I360475,I328362);
nor I_20868 (I360492,I360475,I328353);
and I_20869 (I360509,I360492,I328350);
or I_20870 (I360526,I360509,I328347);
DFFARX1 I_20871  ( .D(I360526), .CLK(I5694_clk), .RSTB(I360294_rst), .Q(I360543) );
nor I_20872 (I360560,I360543,I360396);
DFFARX1 I_20873  ( .D(I360543), .CLK(I5694_clk), .RSTB(I360294_rst), .Q(I360577) );
not I_20874 (I360265,I360577);
nand I_20875 (I360608,I360311,I328362);
and I_20876 (I360625,I360608,I360560);
DFFARX1 I_20877  ( .D(I360608), .CLK(I5694_clk), .RSTB(I360294_rst), .Q(I360262) );
DFFARX1 I_20878  ( .D(I328371), .CLK(I5694_clk), .RSTB(I360294_rst), .Q(I360656) );
nor I_20879 (I360673,I360656,I360379);
nand I_20880 (I360280,I360543,I360673);
nor I_20881 (I360704,I360656,I360444);
not I_20882 (I360277,I360656);
nand I_20883 (I360735,I360656,I360345);
and I_20884 (I360752,I360413,I360735);
DFFARX1 I_20885  ( .D(I360752), .CLK(I5694_clk), .RSTB(I360294_rst), .Q(I360256) );
DFFARX1 I_20886  ( .D(I360656), .CLK(I5694_clk), .RSTB(I360294_rst), .Q(I360259) );
DFFARX1 I_20887  ( .D(I328359), .CLK(I5694_clk), .RSTB(I360294_rst), .Q(I360797) );
not I_20888 (I360814,I360797);
nand I_20889 (I360831,I360814,I360379);
and I_20890 (I360848,I360608,I360831);
DFFARX1 I_20891  ( .D(I360848), .CLK(I5694_clk), .RSTB(I360294_rst), .Q(I360286) );
or I_20892 (I360879,I360814,I360625);
DFFARX1 I_20893  ( .D(I360879), .CLK(I5694_clk), .RSTB(I360294_rst), .Q(I360271) );
nand I_20894 (I360274,I360814,I360704);
not I_20895 (I360957_rst,I5701);
not I_20896 (I360974,I319451);
nor I_20897 (I360991,I319448,I319466);
nand I_20898 (I361008,I360991,I319469);
nor I_20899 (I361025,I360974,I319448);
nand I_20900 (I361042,I361025,I319454);
not I_20901 (I361059,I361042);
not I_20902 (I361076,I319448);
nor I_20903 (I360946,I361042,I361076);
not I_20904 (I361107,I361076);
nand I_20905 (I360931,I361042,I361107);
not I_20906 (I361138,I319463);
nor I_20907 (I361155,I361138,I319445);
and I_20908 (I361172,I361155,I319439);
or I_20909 (I361189,I361172,I319457);
DFFARX1 I_20910  ( .D(I361189), .CLK(I5694_clk), .RSTB(I360957_rst), .Q(I361206) );
nor I_20911 (I361223,I361206,I361059);
DFFARX1 I_20912  ( .D(I361206), .CLK(I5694_clk), .RSTB(I360957_rst), .Q(I361240) );
not I_20913 (I360928,I361240);
nand I_20914 (I361271,I360974,I319463);
and I_20915 (I361288,I361271,I361223);
DFFARX1 I_20916  ( .D(I361271), .CLK(I5694_clk), .RSTB(I360957_rst), .Q(I360925) );
DFFARX1 I_20917  ( .D(I319442), .CLK(I5694_clk), .RSTB(I360957_rst), .Q(I361319) );
nor I_20918 (I361336,I361319,I361042);
nand I_20919 (I360943,I361206,I361336);
nor I_20920 (I361367,I361319,I361107);
not I_20921 (I360940,I361319);
nand I_20922 (I361398,I361319,I361008);
and I_20923 (I361415,I361076,I361398);
DFFARX1 I_20924  ( .D(I361415), .CLK(I5694_clk), .RSTB(I360957_rst), .Q(I360919) );
DFFARX1 I_20925  ( .D(I361319), .CLK(I5694_clk), .RSTB(I360957_rst), .Q(I360922) );
DFFARX1 I_20926  ( .D(I319460), .CLK(I5694_clk), .RSTB(I360957_rst), .Q(I361460) );
not I_20927 (I361477,I361460);
nand I_20928 (I361494,I361477,I361042);
and I_20929 (I361511,I361271,I361494);
DFFARX1 I_20930  ( .D(I361511), .CLK(I5694_clk), .RSTB(I360957_rst), .Q(I360949) );
or I_20931 (I361542,I361477,I361288);
DFFARX1 I_20932  ( .D(I361542), .CLK(I5694_clk), .RSTB(I360957_rst), .Q(I360934) );
nand I_20933 (I360937,I361477,I361367);
not I_20934 (I361620_rst,I5701);
not I_20935 (I361637,I344688);
nor I_20936 (I361654,I344679,I344670);
nand I_20937 (I361671,I361654,I344685);
nor I_20938 (I361688,I361637,I344679);
nand I_20939 (I361705,I361688,I344682);
DFFARX1 I_20940  ( .D(I361705), .CLK(I5694_clk), .RSTB(I361620_rst), .Q(I361722) );
not I_20941 (I361591,I361722);
not I_20942 (I361753,I344679);
not I_20943 (I361770,I361753);
not I_20944 (I361787,I344691);
nor I_20945 (I361804,I361787,I344676);
and I_20946 (I361821,I361804,I344694);
or I_20947 (I361838,I361821,I344667);
DFFARX1 I_20948  ( .D(I361838), .CLK(I5694_clk), .RSTB(I361620_rst), .Q(I361855) );
DFFARX1 I_20949  ( .D(I361855), .CLK(I5694_clk), .RSTB(I361620_rst), .Q(I361588) );
DFFARX1 I_20950  ( .D(I361855), .CLK(I5694_clk), .RSTB(I361620_rst), .Q(I361886) );
DFFARX1 I_20951  ( .D(I361855), .CLK(I5694_clk), .RSTB(I361620_rst), .Q(I361582) );
nand I_20952 (I361917,I361637,I344691);
nand I_20953 (I361934,I361917,I361671);
and I_20954 (I361951,I361753,I361934);
DFFARX1 I_20955  ( .D(I361951), .CLK(I5694_clk), .RSTB(I361620_rst), .Q(I361612) );
and I_20956 (I361585,I361917,I361886);
DFFARX1 I_20957  ( .D(I344697), .CLK(I5694_clk), .RSTB(I361620_rst), .Q(I361996) );
nor I_20958 (I361609,I361996,I361917);
nor I_20959 (I362027,I361996,I361671);
nand I_20960 (I361606,I361705,I362027);
not I_20961 (I361603,I361996);
DFFARX1 I_20962  ( .D(I344673), .CLK(I5694_clk), .RSTB(I361620_rst), .Q(I362072) );
not I_20963 (I362089,I362072);
nor I_20964 (I362106,I362089,I361770);
and I_20965 (I362123,I361996,I362106);
or I_20966 (I362140,I361917,I362123);
DFFARX1 I_20967  ( .D(I362140), .CLK(I5694_clk), .RSTB(I361620_rst), .Q(I361597) );
not I_20968 (I362171,I362089);
nor I_20969 (I362188,I361996,I362171);
nand I_20970 (I361600,I362089,I362188);
nand I_20971 (I361594,I361753,I362171);
not I_20972 (I362266_rst,I5701);
not I_20973 (I362283,I356965);
nor I_20974 (I362300,I356944,I356956);
nand I_20975 (I362317,I362300,I356959);
nor I_20976 (I362334,I362283,I356944);
nand I_20977 (I362351,I362334,I356941);
DFFARX1 I_20978  ( .D(I362351), .CLK(I5694_clk), .RSTB(I362266_rst), .Q(I362368) );
not I_20979 (I362237,I362368);
not I_20980 (I362399,I356944);
not I_20981 (I362416,I362399);
not I_20982 (I362433,I356962);
nor I_20983 (I362450,I362433,I356953);
and I_20984 (I362467,I362450,I356947);
or I_20985 (I362484,I362467,I356971);
DFFARX1 I_20986  ( .D(I362484), .CLK(I5694_clk), .RSTB(I362266_rst), .Q(I362501) );
DFFARX1 I_20987  ( .D(I362501), .CLK(I5694_clk), .RSTB(I362266_rst), .Q(I362234) );
DFFARX1 I_20988  ( .D(I362501), .CLK(I5694_clk), .RSTB(I362266_rst), .Q(I362532) );
DFFARX1 I_20989  ( .D(I362501), .CLK(I5694_clk), .RSTB(I362266_rst), .Q(I362228) );
nand I_20990 (I362563,I362283,I356962);
nand I_20991 (I362580,I362563,I362317);
and I_20992 (I362597,I362399,I362580);
DFFARX1 I_20993  ( .D(I362597), .CLK(I5694_clk), .RSTB(I362266_rst), .Q(I362258) );
and I_20994 (I362231,I362563,I362532);
DFFARX1 I_20995  ( .D(I356968), .CLK(I5694_clk), .RSTB(I362266_rst), .Q(I362642) );
nor I_20996 (I362255,I362642,I362563);
nor I_20997 (I362673,I362642,I362317);
nand I_20998 (I362252,I362351,I362673);
not I_20999 (I362249,I362642);
DFFARX1 I_21000  ( .D(I356950), .CLK(I5694_clk), .RSTB(I362266_rst), .Q(I362718) );
not I_21001 (I362735,I362718);
nor I_21002 (I362752,I362735,I362416);
and I_21003 (I362769,I362642,I362752);
or I_21004 (I362786,I362563,I362769);
DFFARX1 I_21005  ( .D(I362786), .CLK(I5694_clk), .RSTB(I362266_rst), .Q(I362243) );
not I_21006 (I362817,I362735);
nor I_21007 (I362834,I362642,I362817);
nand I_21008 (I362246,I362735,I362834);
nand I_21009 (I362240,I362399,I362817);
not I_21010 (I362912_rst,I5701);
not I_21011 (I362929,I358291);
nor I_21012 (I362946,I358270,I358282);
nand I_21013 (I362963,I362946,I358285);
nor I_21014 (I362980,I362929,I358270);
nand I_21015 (I362997,I362980,I358267);
DFFARX1 I_21016  ( .D(I362997), .CLK(I5694_clk), .RSTB(I362912_rst), .Q(I363014) );
not I_21017 (I362883,I363014);
not I_21018 (I363045,I358270);
not I_21019 (I363062,I363045);
not I_21020 (I363079,I358288);
nor I_21021 (I363096,I363079,I358279);
and I_21022 (I363113,I363096,I358273);
or I_21023 (I363130,I363113,I358297);
DFFARX1 I_21024  ( .D(I363130), .CLK(I5694_clk), .RSTB(I362912_rst), .Q(I363147) );
DFFARX1 I_21025  ( .D(I363147), .CLK(I5694_clk), .RSTB(I362912_rst), .Q(I362880) );
DFFARX1 I_21026  ( .D(I363147), .CLK(I5694_clk), .RSTB(I362912_rst), .Q(I363178) );
DFFARX1 I_21027  ( .D(I363147), .CLK(I5694_clk), .RSTB(I362912_rst), .Q(I362874) );
nand I_21028 (I363209,I362929,I358288);
nand I_21029 (I363226,I363209,I362963);
and I_21030 (I363243,I363045,I363226);
DFFARX1 I_21031  ( .D(I363243), .CLK(I5694_clk), .RSTB(I362912_rst), .Q(I362904) );
and I_21032 (I362877,I363209,I363178);
DFFARX1 I_21033  ( .D(I358294), .CLK(I5694_clk), .RSTB(I362912_rst), .Q(I363288) );
nor I_21034 (I362901,I363288,I363209);
nor I_21035 (I363319,I363288,I362963);
nand I_21036 (I362898,I362997,I363319);
not I_21037 (I362895,I363288);
DFFARX1 I_21038  ( .D(I358276), .CLK(I5694_clk), .RSTB(I362912_rst), .Q(I363364) );
not I_21039 (I363381,I363364);
nor I_21040 (I363398,I363381,I363062);
and I_21041 (I363415,I363288,I363398);
or I_21042 (I363432,I363209,I363415);
DFFARX1 I_21043  ( .D(I363432), .CLK(I5694_clk), .RSTB(I362912_rst), .Q(I362889) );
not I_21044 (I363463,I363381);
nor I_21045 (I363480,I363288,I363463);
nand I_21046 (I362892,I363381,I363480);
nand I_21047 (I362886,I363045,I363463);
not I_21048 (I363558_rst,I5701);
not I_21049 (I363575,I359617);
nor I_21050 (I363592,I359596,I359608);
nand I_21051 (I363609,I363592,I359611);
nor I_21052 (I363626,I363575,I359596);
nand I_21053 (I363643,I363626,I359593);
DFFARX1 I_21054  ( .D(I363643), .CLK(I5694_clk), .RSTB(I363558_rst), .Q(I363660) );
not I_21055 (I363529,I363660);
not I_21056 (I363691,I359596);
not I_21057 (I363708,I363691);
not I_21058 (I363725,I359614);
nor I_21059 (I363742,I363725,I359605);
and I_21060 (I363759,I363742,I359599);
or I_21061 (I363776,I363759,I359623);
DFFARX1 I_21062  ( .D(I363776), .CLK(I5694_clk), .RSTB(I363558_rst), .Q(I363793) );
DFFARX1 I_21063  ( .D(I363793), .CLK(I5694_clk), .RSTB(I363558_rst), .Q(I363526) );
DFFARX1 I_21064  ( .D(I363793), .CLK(I5694_clk), .RSTB(I363558_rst), .Q(I363824) );
DFFARX1 I_21065  ( .D(I363793), .CLK(I5694_clk), .RSTB(I363558_rst), .Q(I363520) );
nand I_21066 (I363855,I363575,I359614);
nand I_21067 (I363872,I363855,I363609);
and I_21068 (I363889,I363691,I363872);
DFFARX1 I_21069  ( .D(I363889), .CLK(I5694_clk), .RSTB(I363558_rst), .Q(I363550) );
and I_21070 (I363523,I363855,I363824);
DFFARX1 I_21071  ( .D(I359620), .CLK(I5694_clk), .RSTB(I363558_rst), .Q(I363934) );
nor I_21072 (I363547,I363934,I363855);
nor I_21073 (I363965,I363934,I363609);
nand I_21074 (I363544,I363643,I363965);
not I_21075 (I363541,I363934);
DFFARX1 I_21076  ( .D(I359602), .CLK(I5694_clk), .RSTB(I363558_rst), .Q(I364010) );
not I_21077 (I364027,I364010);
nor I_21078 (I364044,I364027,I363708);
and I_21079 (I364061,I363934,I364044);
or I_21080 (I364078,I363855,I364061);
DFFARX1 I_21081  ( .D(I364078), .CLK(I5694_clk), .RSTB(I363558_rst), .Q(I363535) );
not I_21082 (I364109,I364027);
nor I_21083 (I364126,I363934,I364109);
nand I_21084 (I363538,I364027,I364126);
nand I_21085 (I363532,I363691,I364109);
not I_21086 (I364204_rst,I5701);
or I_21087 (I364221,I327166,I327178);
or I_21088 (I364238,I327181,I327166);
nor I_21089 (I364255,I327163,I327157);
DFFARX1 I_21090  ( .D(I364255), .CLK(I5694_clk), .RSTB(I364204_rst), .Q(I364272) );
DFFARX1 I_21091  ( .D(I364255), .CLK(I5694_clk), .RSTB(I364204_rst), .Q(I364166) );
not I_21092 (I364303,I327163);
and I_21093 (I364320,I364303,I327169);
nor I_21094 (I364337,I364320,I327178);
nor I_21095 (I364354,I327172,I327175);
DFFARX1 I_21096  ( .D(I364354), .CLK(I5694_clk), .RSTB(I364204_rst), .Q(I364371) );
not I_21097 (I364388,I364371);
DFFARX1 I_21098  ( .D(I364371), .CLK(I5694_clk), .RSTB(I364204_rst), .Q(I364175) );
nor I_21099 (I364419,I327172,I327181);
and I_21100 (I364169,I364419,I364272);
DFFARX1 I_21101  ( .D(I327187), .CLK(I5694_clk), .RSTB(I364204_rst), .Q(I364450) );
and I_21102 (I364467,I364450,I327160);
nand I_21103 (I364484,I364467,I364238);
and I_21104 (I364501,I364371,I364484);
DFFARX1 I_21105  ( .D(I364501), .CLK(I5694_clk), .RSTB(I364204_rst), .Q(I364196) );
nor I_21106 (I364193,I364467,I364337);
not I_21107 (I364546,I364467);
nor I_21108 (I364563,I364221,I364546);
nor I_21109 (I364580,I364467,I364419);
nand I_21110 (I364190,I364238,I364580);
nor I_21111 (I364611,I364467,I364388);
not I_21112 (I364187,I364467);
nand I_21113 (I364178,I364467,I364388);
DFFARX1 I_21114  ( .D(I327184), .CLK(I5694_clk), .RSTB(I364204_rst), .Q(I364656) );
and I_21115 (I364673,I364656,I364563);
or I_21116 (I364690,I364221,I364673);
DFFARX1 I_21117  ( .D(I364690), .CLK(I5694_clk), .RSTB(I364204_rst), .Q(I364181) );
nand I_21118 (I364184,I364656,I364611);
nand I_21119 (I364735,I364656,I364337);
and I_21120 (I364752,I364255,I364735);
DFFARX1 I_21121  ( .D(I364752), .CLK(I5694_clk), .RSTB(I364204_rst), .Q(I364172) );
not I_21122 (I364816_rst,I5701);
nand I_21123 (I364833,I337559,I337571);
and I_21124 (I364850,I364833,I337544);
DFFARX1 I_21125  ( .D(I364850), .CLK(I5694_clk), .RSTB(I364816_rst), .Q(I364867) );
not I_21126 (I364884,I364867);
DFFARX1 I_21127  ( .D(I364867), .CLK(I5694_clk), .RSTB(I364816_rst), .Q(I364784) );
nor I_21128 (I364915,I337562,I337571);
DFFARX1 I_21129  ( .D(I337553), .CLK(I5694_clk), .RSTB(I364816_rst), .Q(I364932) );
DFFARX1 I_21130  ( .D(I364932), .CLK(I5694_clk), .RSTB(I364816_rst), .Q(I364949) );
not I_21131 (I364787,I364949);
DFFARX1 I_21132  ( .D(I364932), .CLK(I5694_clk), .RSTB(I364816_rst), .Q(I364980) );
and I_21133 (I364781,I364867,I364980);
nand I_21134 (I365011,I337550,I337556);
and I_21135 (I365028,I365011,I337568);
DFFARX1 I_21136  ( .D(I365028), .CLK(I5694_clk), .RSTB(I364816_rst), .Q(I365045) );
nor I_21137 (I365062,I365045,I364884);
not I_21138 (I365079,I365045);
nand I_21139 (I364790,I364867,I365079);
DFFARX1 I_21140  ( .D(I337574), .CLK(I5694_clk), .RSTB(I364816_rst), .Q(I365110) );
and I_21141 (I365127,I365110,I337565);
nor I_21142 (I365144,I365127,I365045);
nor I_21143 (I365161,I365127,I365079);
nand I_21144 (I364796,I364915,I365161);
not I_21145 (I364799,I365127);
DFFARX1 I_21146  ( .D(I365127), .CLK(I5694_clk), .RSTB(I364816_rst), .Q(I364778) );
DFFARX1 I_21147  ( .D(I337547), .CLK(I5694_clk), .RSTB(I364816_rst), .Q(I365220) );
nand I_21148 (I365237,I365220,I364932);
and I_21149 (I365254,I364915,I365237);
DFFARX1 I_21150  ( .D(I365254), .CLK(I5694_clk), .RSTB(I364816_rst), .Q(I364808) );
nor I_21151 (I364805,I365220,I365127);
and I_21152 (I365299,I365220,I365062);
or I_21153 (I365316,I364915,I365299);
DFFARX1 I_21154  ( .D(I365316), .CLK(I5694_clk), .RSTB(I364816_rst), .Q(I364793) );
nand I_21155 (I364802,I365220,I365144);
not I_21156 (I365394_rst,I5701);
nand I_21157 (I365411,I344042,I344024);
and I_21158 (I365428,I365411,I344036);
DFFARX1 I_21159  ( .D(I365428), .CLK(I5694_clk), .RSTB(I365394_rst), .Q(I365445) );
not I_21160 (I365462,I365445);
DFFARX1 I_21161  ( .D(I365445), .CLK(I5694_clk), .RSTB(I365394_rst), .Q(I365362) );
nor I_21162 (I365493,I344039,I344024);
DFFARX1 I_21163  ( .D(I344048), .CLK(I5694_clk), .RSTB(I365394_rst), .Q(I365510) );
DFFARX1 I_21164  ( .D(I365510), .CLK(I5694_clk), .RSTB(I365394_rst), .Q(I365527) );
not I_21165 (I365365,I365527);
DFFARX1 I_21166  ( .D(I365510), .CLK(I5694_clk), .RSTB(I365394_rst), .Q(I365558) );
and I_21167 (I365359,I365445,I365558);
nand I_21168 (I365589,I344027,I344051);
and I_21169 (I365606,I365589,I344030);
DFFARX1 I_21170  ( .D(I365606), .CLK(I5694_clk), .RSTB(I365394_rst), .Q(I365623) );
nor I_21171 (I365640,I365623,I365462);
not I_21172 (I365657,I365623);
nand I_21173 (I365368,I365445,I365657);
DFFARX1 I_21174  ( .D(I344033), .CLK(I5694_clk), .RSTB(I365394_rst), .Q(I365688) );
and I_21175 (I365705,I365688,I344045);
nor I_21176 (I365722,I365705,I365623);
nor I_21177 (I365739,I365705,I365657);
nand I_21178 (I365374,I365493,I365739);
not I_21179 (I365377,I365705);
DFFARX1 I_21180  ( .D(I365705), .CLK(I5694_clk), .RSTB(I365394_rst), .Q(I365356) );
DFFARX1 I_21181  ( .D(I344021), .CLK(I5694_clk), .RSTB(I365394_rst), .Q(I365798) );
nand I_21182 (I365815,I365798,I365510);
and I_21183 (I365832,I365493,I365815);
DFFARX1 I_21184  ( .D(I365832), .CLK(I5694_clk), .RSTB(I365394_rst), .Q(I365386) );
nor I_21185 (I365383,I365798,I365705);
and I_21186 (I365877,I365798,I365640);
or I_21187 (I365894,I365493,I365877);
DFFARX1 I_21188  ( .D(I365894), .CLK(I5694_clk), .RSTB(I365394_rst), .Q(I365371) );
nand I_21189 (I365380,I365798,I365722);
not I_21190 (I365972_rst,I5701);
or I_21191 (I365989,I338700,I338715);
or I_21192 (I366006,I338709,I338700);
nor I_21193 (I366023,I338706,I338703);
not I_21194 (I366040,I366023);
DFFARX1 I_21195  ( .D(I366023), .CLK(I5694_clk), .RSTB(I365972_rst), .Q(I365940) );
nand I_21196 (I366071,I366023,I365989);
not I_21197 (I366088,I338706);
and I_21198 (I366105,I366088,I338721);
nor I_21199 (I366122,I366105,I338715);
nor I_21200 (I366139,I338712,I338718);
DFFARX1 I_21201  ( .D(I366139), .CLK(I5694_clk), .RSTB(I365972_rst), .Q(I366156) );
nor I_21202 (I366173,I366156,I366040);
not I_21203 (I366190,I366156);
nand I_21204 (I365946,I366023,I366190);
DFFARX1 I_21205  ( .D(I366156), .CLK(I5694_clk), .RSTB(I365972_rst), .Q(I365937) );
nor I_21206 (I366235,I338712,I338709);
nand I_21207 (I366252,I366006,I366235);
nor I_21208 (I365961,I365989,I366235);
and I_21209 (I366283,I366235,I366173);
or I_21210 (I366300,I366122,I366283);
DFFARX1 I_21211  ( .D(I366300), .CLK(I5694_clk), .RSTB(I365972_rst), .Q(I365949) );
DFFARX1 I_21212  ( .D(I338730), .CLK(I5694_clk), .RSTB(I365972_rst), .Q(I366331) );
and I_21213 (I366348,I366331,I338727);
not I_21214 (I365955,I366348);
DFFARX1 I_21215  ( .D(I366348), .CLK(I5694_clk), .RSTB(I365972_rst), .Q(I366379) );
not I_21216 (I365943,I366379);
and I_21217 (I366410,I366348,I366071);
DFFARX1 I_21218  ( .D(I366410), .CLK(I5694_clk), .RSTB(I365972_rst), .Q(I365934) );
DFFARX1 I_21219  ( .D(I338724), .CLK(I5694_clk), .RSTB(I365972_rst), .Q(I366441) );
and I_21220 (I366458,I366441,I366252);
DFFARX1 I_21221  ( .D(I366458), .CLK(I5694_clk), .RSTB(I365972_rst), .Q(I365964) );
nor I_21222 (I366489,I366441,I366348);
nand I_21223 (I365958,I366122,I366489);
nor I_21224 (I366520,I366441,I366190);
nand I_21225 (I365952,I366006,I366520);
not I_21226 (I366584_rst,I5701);
or I_21227 (I366601,I358939,I358933);
or I_21228 (I366618,I358951,I358939);
nor I_21229 (I366635,I358930,I358957);
or I_21230 (I366573,I366635,I366601);
not I_21231 (I366666,I358930);
and I_21232 (I366683,I366666,I358954);
nor I_21233 (I366700,I366683,I358933);
not I_21234 (I366717,I366700);
nor I_21235 (I366734,I358945,I358960);
DFFARX1 I_21236  ( .D(I366734), .CLK(I5694_clk), .RSTB(I366584_rst), .Q(I366751) );
nor I_21237 (I366768,I366751,I366700);
nand I_21238 (I366558,I366601,I366768);
nor I_21239 (I366799,I366751,I366717);
not I_21240 (I366555,I366751);
nor I_21241 (I366830,I358945,I358951);
or I_21242 (I366567,I366601,I366830);
DFFARX1 I_21243  ( .D(I358942), .CLK(I5694_clk), .RSTB(I366584_rst), .Q(I366861) );
and I_21244 (I366878,I366861,I358948);
nor I_21245 (I366895,I366878,I366751);
DFFARX1 I_21246  ( .D(I366895), .CLK(I5694_clk), .RSTB(I366584_rst), .Q(I366561) );
nor I_21247 (I366576,I366878,I366830);
not I_21248 (I366940,I366878);
nor I_21249 (I366957,I366618,I366940);
nand I_21250 (I366546,I366878,I366717);
DFFARX1 I_21251  ( .D(I358936), .CLK(I5694_clk), .RSTB(I366584_rst), .Q(I366988) );
nor I_21252 (I366564,I366988,I366618);
not I_21253 (I367019,I366988);
and I_21254 (I367036,I366830,I367019);
nor I_21255 (I366570,I366635,I367036);
and I_21256 (I367067,I366988,I366957);
or I_21257 (I367084,I366635,I367067);
DFFARX1 I_21258  ( .D(I367084), .CLK(I5694_clk), .RSTB(I366584_rst), .Q(I366549) );
nand I_21259 (I366552,I366988,I366799);
not I_21260 (I367162_rst,I5701);
nand I_21261 (I367179,I364196,I364184);
and I_21262 (I367196,I367179,I364190);
DFFARX1 I_21263  ( .D(I367196), .CLK(I5694_clk), .RSTB(I367162_rst), .Q(I367213) );
nor I_21264 (I367230,I364181,I364184);
nor I_21265 (I367247,I367230,I367213);
not I_21266 (I367145,I367230);
DFFARX1 I_21267  ( .D(I364166), .CLK(I5694_clk), .RSTB(I367162_rst), .Q(I367278) );
not I_21268 (I367295,I367278);
nor I_21269 (I367312,I367230,I367295);
nand I_21270 (I367148,I367278,I367247);
DFFARX1 I_21271  ( .D(I367278), .CLK(I5694_clk), .RSTB(I367162_rst), .Q(I367130) );
nand I_21272 (I367357,I364175,I364193);
and I_21273 (I367374,I367357,I364187);
DFFARX1 I_21274  ( .D(I367374), .CLK(I5694_clk), .RSTB(I367162_rst), .Q(I367391) );
nor I_21275 (I367151,I367391,I367213);
nand I_21276 (I367142,I367391,I367312);
DFFARX1 I_21277  ( .D(I364178), .CLK(I5694_clk), .RSTB(I367162_rst), .Q(I367436) );
and I_21278 (I367453,I367436,I364172);
DFFARX1 I_21279  ( .D(I367453), .CLK(I5694_clk), .RSTB(I367162_rst), .Q(I367470) );
not I_21280 (I367133,I367470);
nand I_21281 (I367501,I367453,I367391);
and I_21282 (I367518,I367213,I367501);
DFFARX1 I_21283  ( .D(I367518), .CLK(I5694_clk), .RSTB(I367162_rst), .Q(I367124) );
DFFARX1 I_21284  ( .D(I364169), .CLK(I5694_clk), .RSTB(I367162_rst), .Q(I367549) );
nand I_21285 (I367566,I367549,I367213);
and I_21286 (I367583,I367391,I367566);
DFFARX1 I_21287  ( .D(I367583), .CLK(I5694_clk), .RSTB(I367162_rst), .Q(I367154) );
not I_21288 (I367614,I367549);
nor I_21289 (I367631,I367230,I367614);
and I_21290 (I367648,I367549,I367631);
or I_21291 (I367665,I367453,I367648);
DFFARX1 I_21292  ( .D(I367665), .CLK(I5694_clk), .RSTB(I367162_rst), .Q(I367139) );
nand I_21293 (I367136,I367549,I367295);
DFFARX1 I_21294  ( .D(I367549), .CLK(I5694_clk), .RSTB(I367162_rst), .Q(I367127) );
not I_21295 (I367757_rst,I5701);
nand I_21296 (I367774,I354307,I354313);
and I_21297 (I367791,I367774,I354295);
DFFARX1 I_21298  ( .D(I367791), .CLK(I5694_clk), .RSTB(I367757_rst), .Q(I367808) );
nor I_21299 (I367825,I354289,I354313);
nor I_21300 (I367842,I367825,I367808);
not I_21301 (I367740,I367825);
DFFARX1 I_21302  ( .D(I354319), .CLK(I5694_clk), .RSTB(I367757_rst), .Q(I367873) );
not I_21303 (I367890,I367873);
nor I_21304 (I367907,I367825,I367890);
nand I_21305 (I367743,I367873,I367842);
DFFARX1 I_21306  ( .D(I367873), .CLK(I5694_clk), .RSTB(I367757_rst), .Q(I367725) );
nand I_21307 (I367952,I354310,I354301);
and I_21308 (I367969,I367952,I354304);
DFFARX1 I_21309  ( .D(I367969), .CLK(I5694_clk), .RSTB(I367757_rst), .Q(I367986) );
nor I_21310 (I367746,I367986,I367808);
nand I_21311 (I367737,I367986,I367907);
DFFARX1 I_21312  ( .D(I354316), .CLK(I5694_clk), .RSTB(I367757_rst), .Q(I368031) );
and I_21313 (I368048,I368031,I354292);
DFFARX1 I_21314  ( .D(I368048), .CLK(I5694_clk), .RSTB(I367757_rst), .Q(I368065) );
not I_21315 (I367728,I368065);
nand I_21316 (I368096,I368048,I367986);
and I_21317 (I368113,I367808,I368096);
DFFARX1 I_21318  ( .D(I368113), .CLK(I5694_clk), .RSTB(I367757_rst), .Q(I367719) );
DFFARX1 I_21319  ( .D(I354298), .CLK(I5694_clk), .RSTB(I367757_rst), .Q(I368144) );
nand I_21320 (I368161,I368144,I367808);
and I_21321 (I368178,I367986,I368161);
DFFARX1 I_21322  ( .D(I368178), .CLK(I5694_clk), .RSTB(I367757_rst), .Q(I367749) );
not I_21323 (I368209,I368144);
nor I_21324 (I368226,I367825,I368209);
and I_21325 (I368243,I368144,I368226);
or I_21326 (I368260,I368048,I368243);
DFFARX1 I_21327  ( .D(I368260), .CLK(I5694_clk), .RSTB(I367757_rst), .Q(I367734) );
nand I_21328 (I367731,I368144,I367890);
DFFARX1 I_21329  ( .D(I368144), .CLK(I5694_clk), .RSTB(I367757_rst), .Q(I367722) );
not I_21330 (I368352_rst,I5701);
nand I_21331 (I368369,I332530,I332521);
and I_21332 (I368386,I368369,I332539);
DFFARX1 I_21333  ( .D(I368386), .CLK(I5694_clk), .RSTB(I368352_rst), .Q(I368403) );
nor I_21334 (I368420,I332536,I332521);
nor I_21335 (I368437,I368420,I368403);
not I_21336 (I368335,I368420);
DFFARX1 I_21337  ( .D(I332518), .CLK(I5694_clk), .RSTB(I368352_rst), .Q(I368468) );
not I_21338 (I368485,I368468);
nor I_21339 (I368502,I368420,I368485);
nand I_21340 (I368338,I368468,I368437);
DFFARX1 I_21341  ( .D(I368468), .CLK(I5694_clk), .RSTB(I368352_rst), .Q(I368320) );
nand I_21342 (I368547,I332527,I332542);
and I_21343 (I368564,I368547,I332533);
DFFARX1 I_21344  ( .D(I368564), .CLK(I5694_clk), .RSTB(I368352_rst), .Q(I368581) );
nor I_21345 (I368341,I368581,I368403);
nand I_21346 (I368332,I368581,I368502);
DFFARX1 I_21347  ( .D(I332515), .CLK(I5694_clk), .RSTB(I368352_rst), .Q(I368626) );
and I_21348 (I368643,I368626,I332524);
DFFARX1 I_21349  ( .D(I368643), .CLK(I5694_clk), .RSTB(I368352_rst), .Q(I368660) );
not I_21350 (I368323,I368660);
nand I_21351 (I368691,I368643,I368581);
and I_21352 (I368708,I368403,I368691);
DFFARX1 I_21353  ( .D(I368708), .CLK(I5694_clk), .RSTB(I368352_rst), .Q(I368314) );
DFFARX1 I_21354  ( .D(I332512), .CLK(I5694_clk), .RSTB(I368352_rst), .Q(I368739) );
nand I_21355 (I368756,I368739,I368403);
and I_21356 (I368773,I368581,I368756);
DFFARX1 I_21357  ( .D(I368773), .CLK(I5694_clk), .RSTB(I368352_rst), .Q(I368344) );
not I_21358 (I368804,I368739);
nor I_21359 (I368821,I368420,I368804);
and I_21360 (I368838,I368739,I368821);
or I_21361 (I368855,I368643,I368838);
DFFARX1 I_21362  ( .D(I368855), .CLK(I5694_clk), .RSTB(I368352_rst), .Q(I368329) );
nand I_21363 (I368326,I368739,I368485);
DFFARX1 I_21364  ( .D(I368739), .CLK(I5694_clk), .RSTB(I368352_rst), .Q(I368317) );
not I_21365 (I368947_rst,I5701);
nand I_21366 (I368964,I348552,I348564);
and I_21367 (I368981,I368964,I348573);
DFFARX1 I_21368  ( .D(I368981), .CLK(I5694_clk), .RSTB(I368947_rst), .Q(I368998) );
nor I_21369 (I369015,I348567,I348564);
nor I_21370 (I369032,I369015,I368998);
not I_21371 (I368930,I369015);
DFFARX1 I_21372  ( .D(I348561), .CLK(I5694_clk), .RSTB(I368947_rst), .Q(I369063) );
not I_21373 (I369080,I369063);
nor I_21374 (I369097,I369015,I369080);
nand I_21375 (I368933,I369063,I369032);
DFFARX1 I_21376  ( .D(I369063), .CLK(I5694_clk), .RSTB(I368947_rst), .Q(I368915) );
nand I_21377 (I369142,I348558,I348555);
and I_21378 (I369159,I369142,I348546);
DFFARX1 I_21379  ( .D(I369159), .CLK(I5694_clk), .RSTB(I368947_rst), .Q(I369176) );
nor I_21380 (I368936,I369176,I368998);
nand I_21381 (I368927,I369176,I369097);
DFFARX1 I_21382  ( .D(I348570), .CLK(I5694_clk), .RSTB(I368947_rst), .Q(I369221) );
and I_21383 (I369238,I369221,I348549);
DFFARX1 I_21384  ( .D(I369238), .CLK(I5694_clk), .RSTB(I368947_rst), .Q(I369255) );
not I_21385 (I368918,I369255);
nand I_21386 (I369286,I369238,I369176);
and I_21387 (I369303,I368998,I369286);
DFFARX1 I_21388  ( .D(I369303), .CLK(I5694_clk), .RSTB(I368947_rst), .Q(I368909) );
DFFARX1 I_21389  ( .D(I348543), .CLK(I5694_clk), .RSTB(I368947_rst), .Q(I369334) );
nand I_21390 (I369351,I369334,I368998);
and I_21391 (I369368,I369176,I369351);
DFFARX1 I_21392  ( .D(I369368), .CLK(I5694_clk), .RSTB(I368947_rst), .Q(I368939) );
not I_21393 (I369399,I369334);
nor I_21394 (I369416,I369015,I369399);
and I_21395 (I369433,I369334,I369416);
or I_21396 (I369450,I369238,I369433);
DFFARX1 I_21397  ( .D(I369450), .CLK(I5694_clk), .RSTB(I368947_rst), .Q(I368924) );
nand I_21398 (I368921,I369334,I369080);
DFFARX1 I_21399  ( .D(I369334), .CLK(I5694_clk), .RSTB(I368947_rst), .Q(I368912) );
not I_21400 (I369542_rst,I5701);
nand I_21401 (I369559,I361600,I361612);
and I_21402 (I369576,I369559,I361594);
DFFARX1 I_21403  ( .D(I369576), .CLK(I5694_clk), .RSTB(I369542_rst), .Q(I369593) );
nor I_21404 (I369610,I361606,I361612);
nor I_21405 (I369627,I369610,I369593);
not I_21406 (I369525,I369610);
DFFARX1 I_21407  ( .D(I361591), .CLK(I5694_clk), .RSTB(I369542_rst), .Q(I369658) );
not I_21408 (I369675,I369658);
nor I_21409 (I369692,I369610,I369675);
nand I_21410 (I369528,I369658,I369627);
DFFARX1 I_21411  ( .D(I369658), .CLK(I5694_clk), .RSTB(I369542_rst), .Q(I369510) );
nand I_21412 (I369737,I361582,I361597);
and I_21413 (I369754,I369737,I361588);
DFFARX1 I_21414  ( .D(I369754), .CLK(I5694_clk), .RSTB(I369542_rst), .Q(I369771) );
nor I_21415 (I369531,I369771,I369593);
nand I_21416 (I369522,I369771,I369692);
DFFARX1 I_21417  ( .D(I361609), .CLK(I5694_clk), .RSTB(I369542_rst), .Q(I369816) );
and I_21418 (I369833,I369816,I361603);
DFFARX1 I_21419  ( .D(I369833), .CLK(I5694_clk), .RSTB(I369542_rst), .Q(I369850) );
not I_21420 (I369513,I369850);
nand I_21421 (I369881,I369833,I369771);
and I_21422 (I369898,I369593,I369881);
DFFARX1 I_21423  ( .D(I369898), .CLK(I5694_clk), .RSTB(I369542_rst), .Q(I369504) );
DFFARX1 I_21424  ( .D(I361585), .CLK(I5694_clk), .RSTB(I369542_rst), .Q(I369929) );
nand I_21425 (I369946,I369929,I369593);
and I_21426 (I369963,I369771,I369946);
DFFARX1 I_21427  ( .D(I369963), .CLK(I5694_clk), .RSTB(I369542_rst), .Q(I369534) );
not I_21428 (I369994,I369929);
nor I_21429 (I370011,I369610,I369994);
and I_21430 (I370028,I369929,I370011);
or I_21431 (I370045,I369833,I370028);
DFFARX1 I_21432  ( .D(I370045), .CLK(I5694_clk), .RSTB(I369542_rst), .Q(I369519) );
nand I_21433 (I369516,I369929,I369675);
DFFARX1 I_21434  ( .D(I369929), .CLK(I5694_clk), .RSTB(I369542_rst), .Q(I369507) );
not I_21435 (I370137_rst,I5701);
nand I_21436 (I370154,I336945,I336933);
and I_21437 (I370171,I370154,I336918);
DFFARX1 I_21438  ( .D(I370171), .CLK(I5694_clk), .RSTB(I370137_rst), .Q(I370188) );
nor I_21439 (I370205,I336930,I336933);
DFFARX1 I_21440  ( .D(I336942), .CLK(I5694_clk), .RSTB(I370137_rst), .Q(I370222) );
nand I_21441 (I370239,I370222,I370205);
DFFARX1 I_21442  ( .D(I370222), .CLK(I5694_clk), .RSTB(I370137_rst), .Q(I370108) );
nand I_21443 (I370270,I336915,I336939);
and I_21444 (I370287,I370270,I336924);
DFFARX1 I_21445  ( .D(I370287), .CLK(I5694_clk), .RSTB(I370137_rst), .Q(I370304) );
not I_21446 (I370321,I370304);
nor I_21447 (I370338,I370188,I370321);
and I_21448 (I370355,I370205,I370338);
and I_21449 (I370372,I370304,I370239);
DFFARX1 I_21450  ( .D(I370372), .CLK(I5694_clk), .RSTB(I370137_rst), .Q(I370105) );
DFFARX1 I_21451  ( .D(I370304), .CLK(I5694_clk), .RSTB(I370137_rst), .Q(I370099) );
DFFARX1 I_21452  ( .D(I336927), .CLK(I5694_clk), .RSTB(I370137_rst), .Q(I370417) );
and I_21453 (I370434,I370417,I336936);
nand I_21454 (I370451,I370434,I370304);
nor I_21455 (I370126,I370434,I370205);
not I_21456 (I370482,I370434);
nor I_21457 (I370499,I370188,I370482);
nand I_21458 (I370117,I370222,I370499);
nand I_21459 (I370111,I370304,I370482);
or I_21460 (I370544,I370434,I370355);
DFFARX1 I_21461  ( .D(I370544), .CLK(I5694_clk), .RSTB(I370137_rst), .Q(I370114) );
DFFARX1 I_21462  ( .D(I336921), .CLK(I5694_clk), .RSTB(I370137_rst), .Q(I370575) );
and I_21463 (I370592,I370575,I370451);
DFFARX1 I_21464  ( .D(I370592), .CLK(I5694_clk), .RSTB(I370137_rst), .Q(I370129) );
nor I_21465 (I370623,I370575,I370188);
nand I_21466 (I370123,I370434,I370623);
not I_21467 (I370120,I370575);
DFFARX1 I_21468  ( .D(I370575), .CLK(I5694_clk), .RSTB(I370137_rst), .Q(I370668) );
and I_21469 (I370102,I370575,I370668);
not I_21470 (I370732_rst,I5701);
nand I_21471 (I370749,I335058,I335046);
and I_21472 (I370766,I370749,I335031);
DFFARX1 I_21473  ( .D(I370766), .CLK(I5694_clk), .RSTB(I370732_rst), .Q(I370783) );
nor I_21474 (I370800,I335043,I335046);
DFFARX1 I_21475  ( .D(I335055), .CLK(I5694_clk), .RSTB(I370732_rst), .Q(I370817) );
nand I_21476 (I370834,I370817,I370800);
DFFARX1 I_21477  ( .D(I370817), .CLK(I5694_clk), .RSTB(I370732_rst), .Q(I370703) );
nand I_21478 (I370865,I335028,I335052);
and I_21479 (I370882,I370865,I335037);
DFFARX1 I_21480  ( .D(I370882), .CLK(I5694_clk), .RSTB(I370732_rst), .Q(I370899) );
not I_21481 (I370916,I370899);
nor I_21482 (I370933,I370783,I370916);
and I_21483 (I370950,I370800,I370933);
and I_21484 (I370967,I370899,I370834);
DFFARX1 I_21485  ( .D(I370967), .CLK(I5694_clk), .RSTB(I370732_rst), .Q(I370700) );
DFFARX1 I_21486  ( .D(I370899), .CLK(I5694_clk), .RSTB(I370732_rst), .Q(I370694) );
DFFARX1 I_21487  ( .D(I335040), .CLK(I5694_clk), .RSTB(I370732_rst), .Q(I371012) );
and I_21488 (I371029,I371012,I335049);
nand I_21489 (I371046,I371029,I370899);
nor I_21490 (I370721,I371029,I370800);
not I_21491 (I371077,I371029);
nor I_21492 (I371094,I370783,I371077);
nand I_21493 (I370712,I370817,I371094);
nand I_21494 (I370706,I370899,I371077);
or I_21495 (I371139,I371029,I370950);
DFFARX1 I_21496  ( .D(I371139), .CLK(I5694_clk), .RSTB(I370732_rst), .Q(I370709) );
DFFARX1 I_21497  ( .D(I335034), .CLK(I5694_clk), .RSTB(I370732_rst), .Q(I371170) );
and I_21498 (I371187,I371170,I371046);
DFFARX1 I_21499  ( .D(I371187), .CLK(I5694_clk), .RSTB(I370732_rst), .Q(I370724) );
nor I_21500 (I371218,I371170,I370783);
nand I_21501 (I370718,I371029,I371218);
not I_21502 (I370715,I371170);
DFFARX1 I_21503  ( .D(I371170), .CLK(I5694_clk), .RSTB(I370732_rst), .Q(I371263) );
and I_21504 (I370697,I371170,I371263);
not I_21505 (I371327_rst,I5701);
not I_21506 (I371344,I342735);
nor I_21507 (I371361,I342753,I342732);
nand I_21508 (I371378,I371361,I342750);
nor I_21509 (I371395,I371344,I342753);
nand I_21510 (I371412,I371395,I342744);
not I_21511 (I371429,I342753);
not I_21512 (I371446,I371429);
not I_21513 (I371463,I342747);
nor I_21514 (I371480,I371463,I342741);
and I_21515 (I371497,I371480,I342738);
or I_21516 (I371514,I371497,I342729);
DFFARX1 I_21517  ( .D(I371514), .CLK(I5694_clk), .RSTB(I371327_rst), .Q(I371531) );
nand I_21518 (I371548,I371344,I342747);
or I_21519 (I371316,I371548,I371531);
not I_21520 (I371579,I371548);
nor I_21521 (I371596,I371531,I371579);
and I_21522 (I371613,I371429,I371596);
nand I_21523 (I371289,I371548,I371446);
DFFARX1 I_21524  ( .D(I342759), .CLK(I5694_clk), .RSTB(I371327_rst), .Q(I371644) );
or I_21525 (I371310,I371644,I371531);
nor I_21526 (I371675,I371644,I371412);
nor I_21527 (I371692,I371644,I371446);
nand I_21528 (I371295,I371378,I371692);
or I_21529 (I371723,I371644,I371613);
DFFARX1 I_21530  ( .D(I371723), .CLK(I5694_clk), .RSTB(I371327_rst), .Q(I371292) );
not I_21531 (I371298,I371644);
DFFARX1 I_21532  ( .D(I342756), .CLK(I5694_clk), .RSTB(I371327_rst), .Q(I371768) );
not I_21533 (I371785,I371768);
nor I_21534 (I371802,I371785,I371378);
DFFARX1 I_21535  ( .D(I371802), .CLK(I5694_clk), .RSTB(I371327_rst), .Q(I371304) );
nor I_21536 (I371319,I371644,I371785);
nor I_21537 (I371307,I371785,I371548);
not I_21538 (I371861,I371785);
and I_21539 (I371878,I371412,I371861);
nor I_21540 (I371313,I371548,I371878);
nand I_21541 (I371301,I371785,I371675);
not I_21542 (I371956_rst,I5701);
not I_21543 (I371973,I368915);
nor I_21544 (I371990,I368933,I368912);
nand I_21545 (I372007,I371990,I368936);
nor I_21546 (I372024,I371973,I368933);
nand I_21547 (I372041,I372024,I368930);
not I_21548 (I372058,I368933);
not I_21549 (I372075,I372058);
not I_21550 (I372092,I368921);
nor I_21551 (I372109,I372092,I368909);
and I_21552 (I372126,I372109,I368927);
or I_21553 (I372143,I372126,I368939);
DFFARX1 I_21554  ( .D(I372143), .CLK(I5694_clk), .RSTB(I371956_rst), .Q(I372160) );
nand I_21555 (I372177,I371973,I368921);
or I_21556 (I371945,I372177,I372160);
not I_21557 (I372208,I372177);
nor I_21558 (I372225,I372160,I372208);
and I_21559 (I372242,I372058,I372225);
nand I_21560 (I371918,I372177,I372075);
DFFARX1 I_21561  ( .D(I368918), .CLK(I5694_clk), .RSTB(I371956_rst), .Q(I372273) );
or I_21562 (I371939,I372273,I372160);
nor I_21563 (I372304,I372273,I372041);
nor I_21564 (I372321,I372273,I372075);
nand I_21565 (I371924,I372007,I372321);
or I_21566 (I372352,I372273,I372242);
DFFARX1 I_21567  ( .D(I372352), .CLK(I5694_clk), .RSTB(I371956_rst), .Q(I371921) );
not I_21568 (I371927,I372273);
DFFARX1 I_21569  ( .D(I368924), .CLK(I5694_clk), .RSTB(I371956_rst), .Q(I372397) );
not I_21570 (I372414,I372397);
nor I_21571 (I372431,I372414,I372007);
DFFARX1 I_21572  ( .D(I372431), .CLK(I5694_clk), .RSTB(I371956_rst), .Q(I371933) );
nor I_21573 (I371948,I372273,I372414);
nor I_21574 (I371936,I372414,I372177);
not I_21575 (I372490,I372414);
and I_21576 (I372507,I372041,I372490);
nor I_21577 (I371942,I372177,I372507);
nand I_21578 (I371930,I372414,I372304);
not I_21579 (I372585_rst,I5701);
not I_21580 (I372602,I342089);
nor I_21581 (I372619,I342107,I342086);
nand I_21582 (I372636,I372619,I342104);
nor I_21583 (I372653,I372602,I342107);
nand I_21584 (I372670,I372653,I342098);
not I_21585 (I372687,I342107);
not I_21586 (I372704,I372687);
not I_21587 (I372721,I342101);
nor I_21588 (I372738,I372721,I342095);
and I_21589 (I372755,I372738,I342092);
or I_21590 (I372772,I372755,I342083);
DFFARX1 I_21591  ( .D(I372772), .CLK(I5694_clk), .RSTB(I372585_rst), .Q(I372789) );
nand I_21592 (I372806,I372602,I342101);
or I_21593 (I372574,I372806,I372789);
not I_21594 (I372837,I372806);
nor I_21595 (I372854,I372789,I372837);
and I_21596 (I372871,I372687,I372854);
nand I_21597 (I372547,I372806,I372704);
DFFARX1 I_21598  ( .D(I342113), .CLK(I5694_clk), .RSTB(I372585_rst), .Q(I372902) );
or I_21599 (I372568,I372902,I372789);
nor I_21600 (I372933,I372902,I372670);
nor I_21601 (I372950,I372902,I372704);
nand I_21602 (I372553,I372636,I372950);
or I_21603 (I372981,I372902,I372871);
DFFARX1 I_21604  ( .D(I372981), .CLK(I5694_clk), .RSTB(I372585_rst), .Q(I372550) );
not I_21605 (I372556,I372902);
DFFARX1 I_21606  ( .D(I342110), .CLK(I5694_clk), .RSTB(I372585_rst), .Q(I373026) );
not I_21607 (I373043,I373026);
nor I_21608 (I373060,I373043,I372636);
DFFARX1 I_21609  ( .D(I373060), .CLK(I5694_clk), .RSTB(I372585_rst), .Q(I372562) );
nor I_21610 (I372577,I372902,I373043);
nor I_21611 (I372565,I373043,I372806);
not I_21612 (I373119,I373043);
and I_21613 (I373136,I372670,I373119);
nor I_21614 (I372571,I372806,I373136);
nand I_21615 (I372559,I373043,I372933);
not I_21616 (I373214_rst,I5701);
nand I_21617 (I373231,I341546,I341531);
and I_21618 (I373248,I373231,I341540);
DFFARX1 I_21619  ( .D(I373248), .CLK(I5694_clk), .RSTB(I373214_rst), .Q(I373265) );
not I_21620 (I373203,I373265);
DFFARX1 I_21621  ( .D(I373265), .CLK(I5694_clk), .RSTB(I373214_rst), .Q(I373296) );
not I_21622 (I373191,I373296);
nor I_21623 (I373327,I341552,I341531);
not I_21624 (I373344,I373327);
nor I_21625 (I373361,I373265,I373344);
DFFARX1 I_21626  ( .D(I341543), .CLK(I5694_clk), .RSTB(I373214_rst), .Q(I373378) );
not I_21627 (I373395,I373378);
nand I_21628 (I373194,I373378,I373344);
DFFARX1 I_21629  ( .D(I373378), .CLK(I5694_clk), .RSTB(I373214_rst), .Q(I373426) );
and I_21630 (I373179,I373265,I373426);
nand I_21631 (I37345_rst7,I341528,I341522);
and I_21632 (I373474,I37345_rst7,I341537);
DFFARX1 I_21633  ( .D(I373474), .CLK(I5694_clk), .RSTB(I373214_rst), .Q(I373491) );
nor I_21634 (I373508,I373491,I373395);
and I_21635 (I373525,I373327,I373508);
nor I_21636 (I373542,I373491,I373265);
DFFARX1 I_21637  ( .D(I373491), .CLK(I5694_clk), .RSTB(I373214_rst), .Q(I373185) );
DFFARX1 I_21638  ( .D(I341525), .CLK(I5694_clk), .RSTB(I373214_rst), .Q(I373573) );
and I_21639 (I373590,I373573,I341549);
or I_21640 (I373607,I373590,I373525);
DFFARX1 I_21641  ( .D(I373607), .CLK(I5694_clk), .RSTB(I373214_rst), .Q(I373197) );
nand I_21642 (I373206,I373590,I373542);
DFFARX1 I_21643  ( .D(I373590), .CLK(I5694_clk), .RSTB(I373214_rst), .Q(I373176) );
DFFARX1 I_21644  ( .D(I341534), .CLK(I5694_clk), .RSTB(I373214_rst), .Q(I373666) );
nand I_21645 (I373200,I373666,I373361);
DFFARX1 I_21646  ( .D(I373666), .CLK(I5694_clk), .RSTB(I373214_rst), .Q(I373188) );
nand I_21647 (I373711,I373666,I373327);
and I_21648 (I373728,I373378,I373711);
DFFARX1 I_21649  ( .D(I373728), .CLK(I5694_clk), .RSTB(I373214_rst), .Q(I373182) );
not I_21650 (I373792_rst,I5701);
nand I_21651 (I373809,I345334,I345319);
and I_21652 (I373826,I373809,I345313);
DFFARX1 I_21653  ( .D(I373826), .CLK(I5694_clk), .RSTB(I373792_rst), .Q(I373843) );
not I_21654 (I373781,I373843);
DFFARX1 I_21655  ( .D(I373843), .CLK(I5694_clk), .RSTB(I373792_rst), .Q(I373874) );
not I_21656 (I373769,I373874);
nor I_21657 (I373905,I345340,I345319);
not I_21658 (I373922,I373905);
nor I_21659 (I373939,I373843,I373922);
DFFARX1 I_21660  ( .D(I345343), .CLK(I5694_clk), .RSTB(I373792_rst), .Q(I373956) );
not I_21661 (I373973,I373956);
nand I_21662 (I373772,I373956,I373922);
DFFARX1 I_21663  ( .D(I373956), .CLK(I5694_clk), .RSTB(I373792_rst), .Q(I374004) );
and I_21664 (I373757,I373843,I374004);
nand I_21665 (I374035,I345325,I345328);
and I_21666 (I374052,I374035,I345331);
DFFARX1 I_21667  ( .D(I374052), .CLK(I5694_clk), .RSTB(I373792_rst), .Q(I374069) );
nor I_21668 (I374086,I374069,I373973);
and I_21669 (I374103,I373905,I374086);
nor I_21670 (I374120,I374069,I373843);
DFFARX1 I_21671  ( .D(I374069), .CLK(I5694_clk), .RSTB(I373792_rst), .Q(I373763) );
DFFARX1 I_21672  ( .D(I345337), .CLK(I5694_clk), .RSTB(I373792_rst), .Q(I374151) );
and I_21673 (I374168,I374151,I345322);
or I_21674 (I374185,I374168,I374103);
DFFARX1 I_21675  ( .D(I374185), .CLK(I5694_clk), .RSTB(I373792_rst), .Q(I373775) );
nand I_21676 (I373784,I374168,I374120);
DFFARX1 I_21677  ( .D(I374168), .CLK(I5694_clk), .RSTB(I373792_rst), .Q(I373754) );
DFFARX1 I_21678  ( .D(I345316), .CLK(I5694_clk), .RSTB(I373792_rst), .Q(I374244) );
nand I_21679 (I373778,I374244,I373939);
DFFARX1 I_21680  ( .D(I374244), .CLK(I5694_clk), .RSTB(I373792_rst), .Q(I373766) );
nand I_21681 (I374289,I374244,I373905);
and I_21682 (I374306,I373956,I374289);
DFFARX1 I_21683  ( .D(I374306), .CLK(I5694_clk), .RSTB(I373792_rst), .Q(I373760) );
not I_21684 (I374370_rst,I5701);
nand I_21685 (I374387,I349861,I349858);
and I_21686 (I374404,I374387,I349855);
DFFARX1 I_21687  ( .D(I374404), .CLK(I5694_clk), .RSTB(I374370_rst), .Q(I374421) );
not I_21688 (I374438,I374421);
nor I_21689 (I374455,I349879,I349858);
or I_21690 (I374353,I374455,I374421);
not I_21691 (I374341,I374455);
DFFARX1 I_21692  ( .D(I349873), .CLK(I5694_clk), .RSTB(I374370_rst), .Q(I374500) );
nor I_21693 (I374517,I374500,I374455);
nand I_21694 (I374534,I349852,I349864);
and I_21695 (I374551,I374534,I349867);
DFFARX1 I_21696  ( .D(I374551), .CLK(I5694_clk), .RSTB(I374370_rst), .Q(I374568) );
nor I_21697 (I374350,I374568,I374421);
not I_21698 (I374599,I374568);
nor I_21699 (I374616,I374500,I374599);
DFFARX1 I_21700  ( .D(I349876), .CLK(I5694_clk), .RSTB(I374370_rst), .Q(I374633) );
and I_21701 (I374650,I374633,I349882);
or I_21702 (I374359,I374650,I374455);
nand I_21703 (I374338,I374650,I374616);
DFFARX1 I_21704  ( .D(I349870), .CLK(I5694_clk), .RSTB(I374370_rst), .Q(I374695) );
and I_21705 (I374712,I374695,I374438);
nor I_21706 (I374356,I374650,I374712);
nor I_21707 (I374743,I374695,I374500);
DFFARX1 I_21708  ( .D(I374743), .CLK(I5694_clk), .RSTB(I374370_rst), .Q(I374347) );
nor I_21709 (I374362,I374695,I374421);
not I_21710 (I374788,I374695);
nor I_21711 (I374805,I374568,I374788);
and I_21712 (I374822,I374455,I374805);
or I_21713 (I374839,I374650,I374822);
DFFARX1 I_21714  ( .D(I374839), .CLK(I5694_clk), .RSTB(I374370_rst), .Q(I374335) );
nand I_21715 (I374344,I374695,I374517);
nand I_21716 (I374332,I374695,I374599);
not I_21717 (I374931_rst,I5701);
nand I_21718 (I374948,I370715,I370703);
and I_21719 (I374965,I374948,I370700);
DFFARX1 I_21720  ( .D(I374965), .CLK(I5694_clk), .RSTB(I374931_rst), .Q(I374982) );
not I_21721 (I374999,I374982);
nor I_21722 (I375016,I370721,I370703);
or I_21723 (I374914,I375016,I374982);
not I_21724 (I374902,I375016);
DFFARX1 I_21725  ( .D(I370724), .CLK(I5694_clk), .RSTB(I374931_rst), .Q(I375061) );
nor I_21726 (I375078,I375061,I375016);
nand I_21727 (I375095,I370694,I370712);
and I_21728 (I375112,I375095,I370709);
DFFARX1 I_21729  ( .D(I375112), .CLK(I5694_clk), .RSTB(I374931_rst), .Q(I375129) );
nor I_21730 (I374911,I375129,I374982);
not I_21731 (I375160,I375129);
nor I_21732 (I375177,I375061,I375160);
DFFARX1 I_21733  ( .D(I370718), .CLK(I5694_clk), .RSTB(I374931_rst), .Q(I375194) );
and I_21734 (I375211,I375194,I370706);
or I_21735 (I374920,I375211,I375016);
nand I_21736 (I374899,I375211,I375177);
DFFARX1 I_21737  ( .D(I370697), .CLK(I5694_clk), .RSTB(I374931_rst), .Q(I375256) );
and I_21738 (I375273,I375256,I374999);
nor I_21739 (I374917,I375211,I375273);
nor I_21740 (I375304,I375256,I375061);
DFFARX1 I_21741  ( .D(I375304), .CLK(I5694_clk), .RSTB(I374931_rst), .Q(I374908) );
nor I_21742 (I374923,I375256,I374982);
not I_21743 (I375349,I375256);
nor I_21744 (I375366,I375129,I375349);
and I_21745 (I375383,I375016,I375366);
or I_21746 (I375400,I375211,I375383);
DFFARX1 I_21747  ( .D(I375400), .CLK(I5694_clk), .RSTB(I374931_rst), .Q(I374896) );
nand I_21748 (I374905,I375256,I375078);
nand I_21749 (I374893,I375256,I375160);
not I_21750 (I375492_rst,I5701);
nand I_21751 (I375509,I355639,I355630);
and I_21752 (I375526,I375509,I355645);
DFFARX1 I_21753  ( .D(I375526), .CLK(I5694_clk), .RSTB(I375492_rst), .Q(I375543) );
not I_21754 (I375560,I375543);
nor I_21755 (I375577,I355615,I355630);
or I_21756 (I375475,I375577,I375543);
not I_21757 (I375463,I375577);
DFFARX1 I_21758  ( .D(I355618), .CLK(I5694_clk), .RSTB(I375492_rst), .Q(I375622) );
nor I_21759 (I375639,I375622,I375577);
nand I_21760 (I375656,I355636,I355633);
and I_21761 (I375673,I375656,I355621);
DFFARX1 I_21762  ( .D(I375673), .CLK(I5694_clk), .RSTB(I375492_rst), .Q(I375690) );
nor I_21763 (I375472,I375690,I375543);
not I_21764 (I375721,I375690);
nor I_21765 (I375738,I375622,I375721);
DFFARX1 I_21766  ( .D(I355642), .CLK(I5694_clk), .RSTB(I375492_rst), .Q(I375755) );
and I_21767 (I375772,I375755,I355627);
or I_21768 (I375481,I375772,I375577);
nand I_21769 (I375460,I375772,I375738);
DFFARX1 I_21770  ( .D(I355624), .CLK(I5694_clk), .RSTB(I375492_rst), .Q(I375817) );
and I_21771 (I375834,I375817,I375560);
nor I_21772 (I375478,I375772,I375834);
nor I_21773 (I375865,I375817,I375622);
DFFARX1 I_21774  ( .D(I375865), .CLK(I5694_clk), .RSTB(I375492_rst), .Q(I375469) );
nor I_21775 (I375484,I375817,I375543);
not I_21776 (I375910,I375817);
nor I_21777 (I375927,I375690,I375910);
and I_21778 (I375944,I375577,I375927);
or I_21779 (I375961,I375772,I375944);
DFFARX1 I_21780  ( .D(I375961), .CLK(I5694_clk), .RSTB(I375492_rst), .Q(I375457) );
nand I_21781 (I375466,I375817,I375639);
nand I_21782 (I375454,I375817,I375721);
not I_21783 (I376053_rst,I5701);
not I_21784 (I376070,I365371);
nor I_21785 (I376087,I365359,I365365);
nand I_21786 (I376104,I376087,I365356);
DFFARX1 I_21787  ( .D(I376104), .CLK(I5694_clk), .RSTB(I376053_rst), .Q(I376027) );
nor I_21788 (I376135,I376070,I365359);
nand I_21789 (I376152,I376135,I365362);
not I_21790 (I376042,I376152);
DFFARX1 I_21791  ( .D(I376152), .CLK(I5694_clk), .RSTB(I376053_rst), .Q(I376024) );
not I_21792 (I376197,I365359);
not I_21793 (I376214,I376197);
not I_21794 (I376231,I365374);
nor I_21795 (I376248,I376231,I365386);
and I_21796 (I376265,I376248,I365368);
or I_21797 (I376282,I376265,I365383);
DFFARX1 I_21798  ( .D(I376282), .CLK(I5694_clk), .RSTB(I376053_rst), .Q(I376299) );
nor I_21799 (I376316,I376299,I376152);
nor I_21800 (I376333,I376299,I376214);
nand I_21801 (I376039,I376104,I376333);
nand I_21802 (I376364,I376070,I365374);
nand I_21803 (I376381,I376364,I376299);
and I_21804 (I376398,I376364,I376381);
DFFARX1 I_21805  ( .D(I376398), .CLK(I5694_clk), .RSTB(I376053_rst), .Q(I376021) );
DFFARX1 I_21806  ( .D(I376364), .CLK(I5694_clk), .RSTB(I376053_rst), .Q(I376429) );
and I_21807 (I376018,I376197,I376429);
DFFARX1 I_21808  ( .D(I365377), .CLK(I5694_clk), .RSTB(I376053_rst), .Q(I376460) );
not I_21809 (I376477,I376460);
nor I_21810 (I376494,I376152,I376477);
and I_21811 (I376511,I376460,I376494);
nand I_21812 (I376033,I376460,I376214);
DFFARX1 I_21813  ( .D(I376460), .CLK(I5694_clk), .RSTB(I376053_rst), .Q(I376542) );
not I_21814 (I376030,I376542);
DFFARX1 I_21815  ( .D(I365380), .CLK(I5694_clk), .RSTB(I376053_rst), .Q(I376573) );
not I_21816 (I376590,I376573);
or I_21817 (I376607,I376590,I376511);
DFFARX1 I_21818  ( .D(I376607), .CLK(I5694_clk), .RSTB(I376053_rst), .Q(I376036) );
nand I_21819 (I376045,I376590,I376316);
DFFARX1 I_21820  ( .D(I376590), .CLK(I5694_clk), .RSTB(I376053_rst), .Q(I376015) );
not I_21821 (I376699_rst,I5701);
not I_21822 (I376716,I352963);
nor I_21823 (I376733,I352972,I352984);
nand I_21824 (I376750,I376733,I352975);
DFFARX1 I_21825  ( .D(I376750), .CLK(I5694_clk), .RSTB(I376699_rst), .Q(I376670) );
nor I_21826 (I376781,I376716,I352972);
nand I_21827 (I376798,I376781,I352987);
nand I_21828 (I376815,I376798,I376750);
not I_21829 (I376832,I352972);
not I_21830 (I376849,I352993);
nor I_21831 (I376866,I376849,I352969);
and I_21832 (I376883,I376866,I352978);
or I_21833 (I376900,I376883,I352966);
DFFARX1 I_21834  ( .D(I376900), .CLK(I5694_clk), .RSTB(I376699_rst), .Q(I376917) );
nor I_21835 (I376934,I376917,I376798);
nand I_21836 (I376685,I376832,I376934);
not I_21837 (I376682,I376917);
and I_21838 (I376979,I376917,I376815);
DFFARX1 I_21839  ( .D(I376979), .CLK(I5694_clk), .RSTB(I376699_rst), .Q(I376667) );
DFFARX1 I_21840  ( .D(I376917), .CLK(I5694_clk), .RSTB(I376699_rst), .Q(I377010) );
and I_21841 (I376664,I376832,I377010);
nand I_21842 (I377041,I376716,I352993);
not I_21843 (I377058,I377041);
nor I_21844 (I377075,I376917,I377058);
DFFARX1 I_21845  ( .D(I352990), .CLK(I5694_clk), .RSTB(I376699_rst), .Q(I377092) );
nand I_21846 (I377109,I377092,I377041);
and I_21847 (I377126,I376832,I377109);
DFFARX1 I_21848  ( .D(I377126), .CLK(I5694_clk), .RSTB(I376699_rst), .Q(I376691) );
not I_21849 (I377157,I377092);
nand I_21850 (I376679,I377092,I377075);
nand I_21851 (I376673,I377092,I377058);
DFFARX1 I_21852  ( .D(I352981), .CLK(I5694_clk), .RSTB(I376699_rst), .Q(I377202) );
not I_21853 (I377219,I377202);
nor I_21854 (I376688,I377092,I377219);
nor I_21855 (I377250,I377219,I377157);
and I_21856 (I377267,I376798,I377250);
or I_21857 (I377284,I377041,I377267);
DFFARX1 I_21858  ( .D(I377284), .CLK(I5694_clk), .RSTB(I376699_rst), .Q(I376676) );
DFFARX1 I_21859  ( .D(I377219), .CLK(I5694_clk), .RSTB(I376699_rst), .Q(I376661) );
not I_21860 (I377362_rst,I5701);
or I_21861 (I377379,I367734,I367719);
or I_21862 (I377396,I367740,I367734);
DFFARX1 I_21863  ( .D(I377396), .CLK(I5694_clk), .RSTB(I377362_rst), .Q(I377336) );
nor I_21864 (I377427,I367746,I367728);
not I_21865 (I377444,I377427);
not I_21866 (I377461,I367746);
and I_21867 (I377478,I377461,I367725);
nor I_21868 (I377495,I377478,I367719);
nor I_21869 (I377512,I367722,I367731);
DFFARX1 I_21870  ( .D(I377512), .CLK(I5694_clk), .RSTB(I377362_rst), .Q(I377529) );
nand I_21871 (I377546,I377529,I377379);
and I_21872 (I377563,I377495,I377546);
DFFARX1 I_21873  ( .D(I377563), .CLK(I5694_clk), .RSTB(I377362_rst), .Q(I377330) );
nor I_21874 (I377594,I367722,I367740);
DFFARX1 I_21875  ( .D(I377594), .CLK(I5694_clk), .RSTB(I377362_rst), .Q(I377611) );
and I_21876 (I377327,I377427,I377611);
DFFARX1 I_21877  ( .D(I367749), .CLK(I5694_clk), .RSTB(I377362_rst), .Q(I377642) );
and I_21878 (I377659,I377642,I367737);
DFFARX1 I_21879  ( .D(I377659), .CLK(I5694_clk), .RSTB(I377362_rst), .Q(I377676) );
not I_21880 (I377339,I377676);
DFFARX1 I_21881  ( .D(I377659), .CLK(I5694_clk), .RSTB(I377362_rst), .Q(I377324) );
DFFARX1 I_21882  ( .D(I367743), .CLK(I5694_clk), .RSTB(I377362_rst), .Q(I377721) );
not I_21883 (I377738,I377721);
nor I_21884 (I377755,I377396,I377738);
and I_21885 (I377772,I377659,I377755);
or I_21886 (I377789,I377379,I377772);
DFFARX1 I_21887  ( .D(I377789), .CLK(I5694_clk), .RSTB(I377362_rst), .Q(I377345) );
nor I_21888 (I377820,I377721,I377529);
nand I_21889 (I377354,I377495,I377820);
nor I_21890 (I377851,I377721,I377444);
nand I_21891 (I377348,I377594,I377851);
not I_21892 (I377351,I377721);
nand I_21893 (I377342,I377721,I377444);
DFFARX1 I_21894  ( .D(I377721), .CLK(I5694_clk), .RSTB(I377362_rst), .Q(I377333) );
not I_21895 (I377957_rst,I5701);
or I_21896 (I377974,I363538,I363535);
or I_21897 (I377991,I363520,I363538);
DFFARX1 I_21898  ( .D(I377991), .CLK(I5694_clk), .RSTB(I377957_rst), .Q(I377931) );
nor I_21899 (I378022,I363529,I363532);
not I_21900 (I378039,I378022);
not I_21901 (I378056,I363529);
and I_21902 (I378073,I378056,I363544);
nor I_21903 (I378090,I378073,I363535);
nor I_21904 (I378107,I363550,I363526);
DFFARX1 I_21905  ( .D(I378107), .CLK(I5694_clk), .RSTB(I377957_rst), .Q(I378124) );
nand I_21906 (I378141,I378124,I377974);
and I_21907 (I378158,I378090,I378141);
DFFARX1 I_21908  ( .D(I378158), .CLK(I5694_clk), .RSTB(I377957_rst), .Q(I377925) );
nor I_21909 (I378189,I363550,I363520);
DFFARX1 I_21910  ( .D(I378189), .CLK(I5694_clk), .RSTB(I377957_rst), .Q(I378206) );
and I_21911 (I377922,I378022,I378206);
DFFARX1 I_21912  ( .D(I363541), .CLK(I5694_clk), .RSTB(I377957_rst), .Q(I378237) );
and I_21913 (I378254,I378237,I363547);
DFFARX1 I_21914  ( .D(I378254), .CLK(I5694_clk), .RSTB(I377957_rst), .Q(I378271) );
not I_21915 (I377934,I378271);
DFFARX1 I_21916  ( .D(I378254), .CLK(I5694_clk), .RSTB(I377957_rst), .Q(I377919) );
DFFARX1 I_21917  ( .D(I363523), .CLK(I5694_clk), .RSTB(I377957_rst), .Q(I378316) );
not I_21918 (I378333,I378316);
nor I_21919 (I378350,I377991,I378333);
and I_21920 (I378367,I378254,I378350);
or I_21921 (I378384,I377974,I378367);
DFFARX1 I_21922  ( .D(I378384), .CLK(I5694_clk), .RSTB(I377957_rst), .Q(I377940) );
nor I_21923 (I378415,I378316,I378124);
nand I_21924 (I377949,I378090,I378415);
nor I_21925 (I378446,I378316,I378039);
nand I_21926 (I377943,I378189,I378446);
not I_21927 (I377946,I378316);
nand I_21928 (I377937,I378316,I378039);
DFFARX1 I_21929  ( .D(I378316), .CLK(I5694_clk), .RSTB(I377957_rst), .Q(I377928) );
not I_21930 (I378552_rst,I5701);
or I_21931 (I378569,I372553,I372562);
not I_21932 (I378535,I378569);
DFFARX1 I_21933  ( .D(I378569), .CLK(I5694_clk), .RSTB(I378552_rst), .Q(I378514) );
or I_21934 (I378614,I372571,I372553);
nor I_21935 (I378631,I372565,I372559);
nor I_21936 (I378648,I378631,I378569);
not I_21937 (I378665,I372565);
and I_21938 (I378682,I378665,I372568);
nor I_21939 (I378699,I378682,I372562);
DFFARX1 I_21940  ( .D(I378699), .CLK(I5694_clk), .RSTB(I378552_rst), .Q(I378716) );
nor I_21941 (I378733,I372556,I372574);
DFFARX1 I_21942  ( .D(I378733), .CLK(I5694_clk), .RSTB(I378552_rst), .Q(I378750) );
nor I_21943 (I378541,I378750,I378699);
not I_21944 (I378781,I378750);
nor I_21945 (I378798,I372556,I372571);
nand I_21946 (I378815,I378699,I378798);
and I_21947 (I378832,I378614,I378815);
DFFARX1 I_21948  ( .D(I378832), .CLK(I5694_clk), .RSTB(I378552_rst), .Q(I378544) );
DFFARX1 I_21949  ( .D(I372577), .CLK(I5694_clk), .RSTB(I378552_rst), .Q(I378863) );
and I_21950 (I378880,I378863,I372550);
nor I_21951 (I378897,I378880,I378781);
and I_21952 (I378914,I378798,I378897);
or I_21953 (I378931,I378631,I378914);
DFFARX1 I_21954  ( .D(I378931), .CLK(I5694_clk), .RSTB(I378552_rst), .Q(I378529) );
not I_21955 (I378962,I378880);
nor I_21956 (I378979,I378569,I378962);
nand I_21957 (I378532,I378614,I378979);
nand I_21958 (I378526,I378750,I378962);
DFFARX1 I_21959  ( .D(I378880), .CLK(I5694_clk), .RSTB(I378552_rst), .Q(I378520) );
DFFARX1 I_21960  ( .D(I372547), .CLK(I5694_clk), .RSTB(I378552_rst), .Q(I379038) );
nand I_21961 (I378538,I379038,I378648);
DFFARX1 I_21962  ( .D(I379038), .CLK(I5694_clk), .RSTB(I378552_rst), .Q(I37906_rst9) );
not I_21963 (I378523,I37906_rst9);
and I_21964 (I378517,I379038,I378716);
not I_21965 (I379147_rst,I5701);
not I_21966 (I379164,I377342);
nor I_21967 (I379181,I377336,I377327);
nand I_21968 (I379198,I379181,I377339);
nor I_21969 (I379215,I379164,I377336);
nand I_21970 (I379232,I379215,I377354);
not I_21971 (I379249,I379232);
not I_21972 (I379266,I377336);
nor I_21973 (I379136,I379232,I379266);
not I_21974 (I379297,I379266);
nand I_21975 (I379121,I379232,I379297);
not I_21976 (I379328,I377330);
nor I_21977 (I379345,I379328,I377324);
and I_21978 (I379362,I379345,I377351);
or I_21979 (I379379,I379362,I377348);
DFFARX1 I_21980  ( .D(I379379), .CLK(I5694_clk), .RSTB(I379147_rst), .Q(I379396) );
nor I_21981 (I379413,I379396,I379249);
DFFARX1 I_21982  ( .D(I379396), .CLK(I5694_clk), .RSTB(I379147_rst), .Q(I379430) );
not I_21983 (I379118,I379430);
nand I_21984 (I379461,I379164,I377330);
and I_21985 (I379478,I379461,I379413);
DFFARX1 I_21986  ( .D(I379461), .CLK(I5694_clk), .RSTB(I379147_rst), .Q(I379115) );
DFFARX1 I_21987  ( .D(I377345), .CLK(I5694_clk), .RSTB(I379147_rst), .Q(I379509) );
nor I_21988 (I379526,I379509,I379232);
nand I_21989 (I379133,I379396,I379526);
nor I_21990 (I379557,I379509,I379297);
not I_21991 (I379130,I379509);
nand I_21992 (I379588,I379509,I379198);
and I_21993 (I379605,I379266,I379588);
DFFARX1 I_21994  ( .D(I379605), .CLK(I5694_clk), .RSTB(I379147_rst), .Q(I379109) );
DFFARX1 I_21995  ( .D(I379509), .CLK(I5694_clk), .RSTB(I379147_rst), .Q(I379112) );
DFFARX1 I_21996  ( .D(I377333), .CLK(I5694_clk), .RSTB(I379147_rst), .Q(I379650) );
not I_21997 (I379667,I379650);
nand I_21998 (I379684,I379667,I379232);
and I_21999 (I379701,I379461,I379684);
DFFARX1 I_22000  ( .D(I379701), .CLK(I5694_clk), .RSTB(I379147_rst), .Q(I379139) );
or I_22001 (I379732,I379667,I379478);
DFFARX1 I_22002  ( .D(I379732), .CLK(I5694_clk), .RSTB(I379147_rst), .Q(I379124) );
nand I_22003 (I379127,I379667,I379557);
not I_22004 (I379810_rst,I5701);
not I_22005 (I379827,I370117);
nor I_22006 (I379844,I370114,I370105);
nand I_22007 (I379861,I379844,I370108);
nor I_22008 (I379878,I379827,I370114);
nand I_22009 (I379895,I379878,I370102);
not I_22010 (I379912,I379895);
not I_22011 (I379929,I370114);
nor I_22012 (I379799,I379895,I379929);
not I_22013 (I379960,I379929);
nand I_22014 (I379784,I379895,I379960);
not I_22015 (I379991,I370123);
nor I_22016 (I380008,I379991,I370126);
and I_22017 (I380025,I380008,I370111);
or I_22018 (I380042,I380025,I370099);
DFFARX1 I_22019  ( .D(I380042), .CLK(I5694_clk), .RSTB(I379810_rst), .Q(I380059) );
nor I_22020 (I380076,I380059,I379912);
DFFARX1 I_22021  ( .D(I380059), .CLK(I5694_clk), .RSTB(I379810_rst), .Q(I380093) );
not I_22022 (I379781,I380093);
nand I_22023 (I380124,I379827,I370123);
and I_22024 (I380141,I380124,I380076);
DFFARX1 I_22025  ( .D(I380124), .CLK(I5694_clk), .RSTB(I379810_rst), .Q(I379778) );
DFFARX1 I_22026  ( .D(I370120), .CLK(I5694_clk), .RSTB(I379810_rst), .Q(I380172) );
nor I_22027 (I380189,I380172,I379895);
nand I_22028 (I379796,I380059,I380189);
nor I_22029 (I380220,I380172,I379960);
not I_22030 (I379793,I380172);
nand I_22031 (I380251,I380172,I379861);
and I_22032 (I380268,I379929,I380251);
DFFARX1 I_22033  ( .D(I380268), .CLK(I5694_clk), .RSTB(I379810_rst), .Q(I379772) );
DFFARX1 I_22034  ( .D(I380172), .CLK(I5694_clk), .RSTB(I379810_rst), .Q(I379775) );
DFFARX1 I_22035  ( .D(I370129), .CLK(I5694_clk), .RSTB(I379810_rst), .Q(I380313) );
not I_22036 (I380330,I380313);
nand I_22037 (I380347,I380330,I379895);
and I_22038 (I380364,I380124,I380347);
DFFARX1 I_22039  ( .D(I380364), .CLK(I5694_clk), .RSTB(I379810_rst), .Q(I379802) );
or I_22040 (I380395,I380330,I380141);
DFFARX1 I_22041  ( .D(I380395), .CLK(I5694_clk), .RSTB(I379810_rst), .Q(I379787) );
nand I_22042 (I379790,I380330,I380220);
not I_22043 (I380473_rst,I5701);
nand I_22044 (I380490,I373191,I373203);
and I_22045 (I380507,I380490,I373176);
DFFARX1 I_22046  ( .D(I380507), .CLK(I5694_clk), .RSTB(I380473_rst), .Q(I380524) );
not I_22047 (I380541,I380524);
DFFARX1 I_22048  ( .D(I380524), .CLK(I5694_clk), .RSTB(I380473_rst), .Q(I380441) );
nor I_22049 (I380572,I373194,I373203);
DFFARX1 I_22050  ( .D(I373185), .CLK(I5694_clk), .RSTB(I380473_rst), .Q(I380589) );
DFFARX1 I_22051  ( .D(I380589), .CLK(I5694_clk), .RSTB(I380473_rst), .Q(I380606) );
not I_22052 (I380444,I380606);
DFFARX1 I_22053  ( .D(I380589), .CLK(I5694_clk), .RSTB(I380473_rst), .Q(I380637) );
and I_22054 (I380438,I380524,I380637);
nand I_22055 (I380668,I373182,I373188);
and I_22056 (I380685,I380668,I373200);
DFFARX1 I_22057  ( .D(I380685), .CLK(I5694_clk), .RSTB(I380473_rst), .Q(I380702) );
nor I_22058 (I380719,I380702,I380541);
not I_22059 (I380736,I380702);
nand I_22060 (I380447,I380524,I380736);
DFFARX1 I_22061  ( .D(I373206), .CLK(I5694_clk), .RSTB(I380473_rst), .Q(I380767) );
and I_22062 (I380784,I380767,I373197);
nor I_22063 (I380801,I380784,I380702);
nor I_22064 (I380818,I380784,I380736);
nand I_22065 (I380453,I380572,I380818);
not I_22066 (I380456,I380784);
DFFARX1 I_22067  ( .D(I380784), .CLK(I5694_clk), .RSTB(I380473_rst), .Q(I380435) );
DFFARX1 I_22068  ( .D(I373179), .CLK(I5694_clk), .RSTB(I380473_rst), .Q(I380877) );
nand I_22069 (I380894,I380877,I380589);
and I_22070 (I380911,I380572,I380894);
DFFARX1 I_22071  ( .D(I380911), .CLK(I5694_clk), .RSTB(I380473_rst), .Q(I380465) );
nor I_22072 (I380462,I380877,I380784);
and I_22073 (I380956,I380877,I380719);
or I_22074 (I380973,I380572,I380956);
DFFARX1 I_22075  ( .D(I380973), .CLK(I5694_clk), .RSTB(I380473_rst), .Q(I380450) );
nand I_22076 (I380459,I380877,I380801);
not I_22077 (I381051_rst,I5701);
nand I_22078 (I381068,I377943,I377928);
and I_22079 (I381085,I381068,I377937);
DFFARX1 I_22080  ( .D(I381085), .CLK(I5694_clk), .RSTB(I381051_rst), .Q(I381102) );
not I_22081 (I381119,I381102);
DFFARX1 I_22082  ( .D(I381102), .CLK(I5694_clk), .RSTB(I381051_rst), .Q(I381019) );
nor I_22083 (I381150,I377946,I377928);
DFFARX1 I_22084  ( .D(I377925), .CLK(I5694_clk), .RSTB(I381051_rst), .Q(I381167) );
DFFARX1 I_22085  ( .D(I381167), .CLK(I5694_clk), .RSTB(I381051_rst), .Q(I381184) );
not I_22086 (I381022,I381184);
DFFARX1 I_22087  ( .D(I381167), .CLK(I5694_clk), .RSTB(I381051_rst), .Q(I381215) );
and I_22088 (I381016,I381102,I381215);
nand I_22089 (I381246,I377949,I377922);
and I_22090 (I381263,I381246,I377940);
DFFARX1 I_22091  ( .D(I381263), .CLK(I5694_clk), .RSTB(I381051_rst), .Q(I381280) );
nor I_22092 (I381297,I381280,I381119);
not I_22093 (I381314,I381280);
nand I_22094 (I381025,I381102,I381314);
DFFARX1 I_22095  ( .D(I377934), .CLK(I5694_clk), .RSTB(I381051_rst), .Q(I381345) );
and I_22096 (I381362,I381345,I377919);
nor I_22097 (I381379,I381362,I381280);
nor I_22098 (I381396,I381362,I381314);
nand I_22099 (I381031,I381150,I381396);
not I_22100 (I381034,I381362);
DFFARX1 I_22101  ( .D(I381362), .CLK(I5694_clk), .RSTB(I381051_rst), .Q(I381013) );
DFFARX1 I_22102  ( .D(I377931), .CLK(I5694_clk), .RSTB(I381051_rst), .Q(I381455) );
nand I_22103 (I381472,I381455,I381167);
and I_22104 (I381489,I381150,I381472);
DFFARX1 I_22105  ( .D(I381489), .CLK(I5694_clk), .RSTB(I381051_rst), .Q(I381043) );
nor I_22106 (I381040,I381455,I381362);
and I_22107 (I381534,I381455,I381297);
or I_22108 (I381551,I381150,I381534);
DFFARX1 I_22109  ( .D(I381551), .CLK(I5694_clk), .RSTB(I381051_rst), .Q(I381028) );
nand I_22110 (I381037,I381455,I381379);
not I_22111 (I381629_rst,I5701);
nand I_22112 (I381646,I374347,I374362);
and I_22113 (I381663,I381646,I374350);
DFFARX1 I_22114  ( .D(I381663), .CLK(I5694_clk), .RSTB(I381629_rst), .Q(I381680) );
not I_22115 (I381697,I381680);
DFFARX1 I_22116  ( .D(I381680), .CLK(I5694_clk), .RSTB(I381629_rst), .Q(I381597) );
nor I_22117 (I381728,I374359,I374362);
DFFARX1 I_22118  ( .D(I374344), .CLK(I5694_clk), .RSTB(I381629_rst), .Q(I381745) );
DFFARX1 I_22119  ( .D(I381745), .CLK(I5694_clk), .RSTB(I381629_rst), .Q(I381762) );
not I_22120 (I381600,I381762);
DFFARX1 I_22121  ( .D(I381745), .CLK(I5694_clk), .RSTB(I381629_rst), .Q(I381793) );
and I_22122 (I381594,I381680,I381793);
nand I_22123 (I381824,I374335,I374332);
and I_22124 (I381841,I381824,I374338);
DFFARX1 I_22125  ( .D(I381841), .CLK(I5694_clk), .RSTB(I381629_rst), .Q(I381858) );
nor I_22126 (I381875,I381858,I381697);
not I_22127 (I381892,I381858);
nand I_22128 (I381603,I381680,I381892);
DFFARX1 I_22129  ( .D(I374341), .CLK(I5694_clk), .RSTB(I381629_rst), .Q(I381923) );
and I_22130 (I381940,I381923,I374353);
nor I_22131 (I381957,I381940,I381858);
nor I_22132 (I381974,I381940,I381892);
nand I_22133 (I381609,I381728,I381974);
not I_22134 (I381612,I381940);
DFFARX1 I_22135  ( .D(I381940), .CLK(I5694_clk), .RSTB(I381629_rst), .Q(I381591) );
DFFARX1 I_22136  ( .D(I374356), .CLK(I5694_clk), .RSTB(I381629_rst), .Q(I382033) );
nand I_22137 (I382050,I382033,I381745);
and I_22138 (I382067,I381728,I382050);
DFFARX1 I_22139  ( .D(I382067), .CLK(I5694_clk), .RSTB(I381629_rst), .Q(I381621) );
nor I_22140 (I381618,I382033,I381940);
and I_22141 (I382112,I382033,I381875);
or I_22142 (I382129,I381728,I382112);
DFFARX1 I_22143  ( .D(I382129), .CLK(I5694_clk), .RSTB(I381629_rst), .Q(I381606) );
nand I_22144 (I381615,I382033,I381957);
not I_22145 (I382207_rst,I5701);
nand I_22146 (I382224,I371936,I371927);
and I_22147 (I382241,I382224,I371945);
DFFARX1 I_22148  ( .D(I382241), .CLK(I5694_clk), .RSTB(I382207_rst), .Q(I382258) );
nor I_22149 (I382275,I371942,I371927);
nor I_22150 (I382292,I382275,I382258);
not I_22151 (I382190,I382275);
DFFARX1 I_22152  ( .D(I371924), .CLK(I5694_clk), .RSTB(I382207_rst), .Q(I382323) );
not I_22153 (I382340,I382323);
nor I_22154 (I382357,I382275,I382340);
nand I_22155 (I382193,I382323,I382292);
DFFARX1 I_22156  ( .D(I382323), .CLK(I5694_clk), .RSTB(I382207_rst), .Q(I382175) );
nand I_22157 (I382402,I371933,I371948);
and I_22158 (I382419,I382402,I371939);
DFFARX1 I_22159  ( .D(I382419), .CLK(I5694_clk), .RSTB(I382207_rst), .Q(I382436) );
nor I_22160 (I382196,I382436,I382258);
nand I_22161 (I382187,I382436,I382357);
DFFARX1 I_22162  ( .D(I371921), .CLK(I5694_clk), .RSTB(I382207_rst), .Q(I382481) );
and I_22163 (I382498,I382481,I371930);
DFFARX1 I_22164  ( .D(I382498), .CLK(I5694_clk), .RSTB(I382207_rst), .Q(I382515) );
not I_22165 (I382178,I382515);
nand I_22166 (I382546,I382498,I382436);
and I_22167 (I382563,I382258,I382546);
DFFARX1 I_22168  ( .D(I382563), .CLK(I5694_clk), .RSTB(I382207_rst), .Q(I382169) );
DFFARX1 I_22169  ( .D(I371918), .CLK(I5694_clk), .RSTB(I382207_rst), .Q(I382594) );
nand I_22170 (I382611,I382594,I382258);
and I_22171 (I382628,I382436,I382611);
DFFARX1 I_22172  ( .D(I382628), .CLK(I5694_clk), .RSTB(I382207_rst), .Q(I382199) );
not I_22173 (I382659,I382594);
nor I_22174 (I382676,I382275,I382659);
and I_22175 (I382693,I382594,I382676);
or I_22176 (I382710,I382498,I382693);
DFFARX1 I_22177  ( .D(I382710), .CLK(I5694_clk), .RSTB(I382207_rst), .Q(I382184) );
nand I_22178 (I382181,I382594,I382340);
DFFARX1 I_22179  ( .D(I382594), .CLK(I5694_clk), .RSTB(I382207_rst), .Q(I382172) );
not I_22180 (I382802_rst,I5701);
not I_22181 (I382819,I379790);
nor I_22182 (I382836,I379787,I379775);
nand I_22183 (I382853,I382836,I379778);
DFFARX1 I_22184  ( .D(I382853), .CLK(I5694_clk), .RSTB(I382802_rst), .Q(I382776) );
nor I_22185 (I382884,I382819,I379787);
nand I_22186 (I382901,I382884,I379784);
not I_22187 (I382791,I382901);
DFFARX1 I_22188  ( .D(I382901), .CLK(I5694_clk), .RSTB(I382802_rst), .Q(I382773) );
not I_22189 (I382946,I379787);
not I_22190 (I382963,I382946);
not I_22191 (I382980,I379796);
nor I_22192 (I382997,I382980,I379772);
and I_22193 (I383014,I382997,I379793);
or I_22194 (I383031,I383014,I379781);
DFFARX1 I_22195  ( .D(I383031), .CLK(I5694_clk), .RSTB(I382802_rst), .Q(I383048) );
nor I_22196 (I383065,I383048,I382901);
nor I_22197 (I383082,I383048,I382963);
nand I_22198 (I382788,I382853,I383082);
nand I_22199 (I383113,I382819,I379796);
nand I_22200 (I383130,I383113,I383048);
and I_22201 (I383147,I383113,I383130);
DFFARX1 I_22202  ( .D(I383147), .CLK(I5694_clk), .RSTB(I382802_rst), .Q(I382770) );
DFFARX1 I_22203  ( .D(I383113), .CLK(I5694_clk), .RSTB(I382802_rst), .Q(I383178) );
and I_22204 (I382767,I382946,I383178);
DFFARX1 I_22205  ( .D(I379802), .CLK(I5694_clk), .RSTB(I382802_rst), .Q(I383209) );
not I_22206 (I383226,I383209);
nor I_22207 (I383243,I382901,I383226);
and I_22208 (I383260,I383209,I383243);
nand I_22209 (I382782,I383209,I382963);
DFFARX1 I_22210  ( .D(I383209), .CLK(I5694_clk), .RSTB(I382802_rst), .Q(I383291) );
not I_22211 (I382779,I383291);
DFFARX1 I_22212  ( .D(I379799), .CLK(I5694_clk), .RSTB(I382802_rst), .Q(I383322) );
not I_22213 (I383339,I383322);
or I_22214 (I383356,I383339,I383260);
DFFARX1 I_22215  ( .D(I383356), .CLK(I5694_clk), .RSTB(I382802_rst), .Q(I382785) );
nand I_22216 (I382794,I383339,I383065);
DFFARX1 I_22217  ( .D(I383339), .CLK(I5694_clk), .RSTB(I382802_rst), .Q(I382764) );
not I_22218 (I383448_rst,I5701);
not I_22219 (I383465,I378520);
nor I_22220 (I383482,I378541,I378514);
nand I_22221 (I383499,I383482,I378529);
DFFARX1 I_22222  ( .D(I383499), .CLK(I5694_clk), .RSTB(I383448_rst), .Q(I383422) );
nor I_22223 (I383530,I383465,I378541);
nand I_22224 (I383547,I383530,I378544);
not I_22225 (I383437,I383547);
DFFARX1 I_22226  ( .D(I383547), .CLK(I5694_clk), .RSTB(I383448_rst), .Q(I383419) );
not I_22227 (I383592,I378541);
not I_22228 (I383609,I383592);
not I_22229 (I383626,I378517);
nor I_22230 (I383643,I383626,I378535);
and I_22231 (I383660,I383643,I378523);
or I_22232 (I383677,I383660,I378526);
DFFARX1 I_22233  ( .D(I383677), .CLK(I5694_clk), .RSTB(I383448_rst), .Q(I383694) );
nor I_22234 (I383711,I383694,I383547);
nor I_22235 (I383728,I383694,I383609);
nand I_22236 (I383434,I383499,I383728);
nand I_22237 (I383759,I383465,I378517);
nand I_22238 (I383776,I383759,I383694);
and I_22239 (I383793,I383759,I383776);
DFFARX1 I_22240  ( .D(I383793), .CLK(I5694_clk), .RSTB(I383448_rst), .Q(I383416) );
DFFARX1 I_22241  ( .D(I383759), .CLK(I5694_clk), .RSTB(I383448_rst), .Q(I383824) );
and I_22242 (I383413,I383592,I383824);
DFFARX1 I_22243  ( .D(I378538), .CLK(I5694_clk), .RSTB(I383448_rst), .Q(I383855) );
not I_22244 (I383872,I383855);
nor I_22245 (I383889,I383547,I383872);
and I_22246 (I383906,I383855,I383889);
nand I_22247 (I383428,I383855,I383609);
DFFARX1 I_22248  ( .D(I383855), .CLK(I5694_clk), .RSTB(I383448_rst), .Q(I383937) );
not I_22249 (I383425,I383937);
DFFARX1 I_22250  ( .D(I378532), .CLK(I5694_clk), .RSTB(I383448_rst), .Q(I383968) );
not I_22251 (I383985,I383968);
or I_22252 (I384002,I383985,I383906);
DFFARX1 I_22253  ( .D(I384002), .CLK(I5694_clk), .RSTB(I383448_rst), .Q(I383431) );
nand I_22254 (I383440,I383985,I383711);
DFFARX1 I_22255  ( .D(I383985), .CLK(I5694_clk), .RSTB(I383448_rst), .Q(I383410) );
not I_22256 (I384094_rst,I5701);
not I_22257 (I384111,I382770);
nor I_22258 (I384128,I382767,I382791);
nand I_22259 (I384145,I384128,I382788);
nor I_22260 (I384162,I384111,I382767);
nand I_22261 (I384179,I384162,I382794);
not I_22262 (I384196,I384179);
not I_22263 (I384213,I382767);
nor I_22264 (I384083,I384179,I384213);
not I_22265 (I384244,I384213);
nand I_22266 (I384068,I384179,I384244);
not I_22267 (I384275,I382785);
nor I_22268 (I384292,I384275,I382776);
and I_22269 (I384309,I384292,I382773);
or I_22270 (I384326,I384309,I382782);
DFFARX1 I_22271  ( .D(I384326), .CLK(I5694_clk), .RSTB(I384094_rst), .Q(I384343) );
nor I_22272 (I384360,I384343,I384196);
DFFARX1 I_22273  ( .D(I384343), .CLK(I5694_clk), .RSTB(I384094_rst), .Q(I384377) );
not I_22274 (I384065,I384377);
nand I_22275 (I384408,I384111,I382785);
and I_22276 (I384425,I384408,I384360);
DFFARX1 I_22277  ( .D(I384408), .CLK(I5694_clk), .RSTB(I384094_rst), .Q(I384062) );
DFFARX1 I_22278  ( .D(I382764), .CLK(I5694_clk), .RSTB(I384094_rst), .Q(I384456) );
nor I_22279 (I384473,I384456,I384179);
nand I_22280 (I384080,I384343,I384473);
nor I_22281 (I384504,I384456,I384244);
not I_22282 (I384077,I384456);
nand I_22283 (I384535,I384456,I384145);
and I_22284 (I384552,I384213,I384535);
DFFARX1 I_22285  ( .D(I384552), .CLK(I5694_clk), .RSTB(I384094_rst), .Q(I384056) );
DFFARX1 I_22286  ( .D(I384456), .CLK(I5694_clk), .RSTB(I384094_rst), .Q(I384059) );
DFFARX1 I_22287  ( .D(I382779), .CLK(I5694_clk), .RSTB(I384094_rst), .Q(I384597) );
not I_22288 (I384614,I384597);
nand I_22289 (I384631,I384614,I384179);
and I_22290 (I384648,I384408,I384631);
DFFARX1 I_22291  ( .D(I384648), .CLK(I5694_clk), .RSTB(I384094_rst), .Q(I384086) );
or I_22292 (I38467_rst9,I384614,I384425);
DFFARX1 I_22293  ( .D(I38467_rst9), .CLK(I5694_clk), .RSTB(I384094_rst), .Q(I384071) );
nand I_22294 (I384074,I384614,I384504);
endmodule


