module test_I7026(I1477,I3521,I3846,I1470,I5122,I7026);
input I1477,I3521,I3846,I1470,I5122;
output I7026;
wire I5416,I3380,I5070,I5249,I3356,I5105,I5481;
nand I_0(I5416,I5122,I3356);
nand I_1(I3380,I3521,I3846);
not I_2(I7026,I5070);
and I_3(I5070,I5249,I5481);
not I_4(I5249,I3380);
DFFARX1 I_5(I1470,,,I3356,);
not I_6(I5105,I1477);
DFFARX1 I_7(I5416,I1470,I5105,,,I5481,);
endmodule


