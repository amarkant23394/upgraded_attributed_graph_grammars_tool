module test_I11088(I9576,I1477,I1470,I9771,I11088);
input I9576,I1477,I1470,I9771;
output I11088;
wire I9477,I10647,I9833,I9491,I10698,I9816,I9480,I9468,I9960,I10681,I9943,I11009,I9621,I9456,I9864;
nor I_0(I9477,I9771,I9833);
not I_1(I10647,I1477);
and I_2(I9833,I9816);
not I_3(I9491,I1477);
nand I_4(I10698,I10681,I9456);
DFFARX1 I_5(I1470,I9491,,,I9816,);
or I_6(I9480,I9771,I9576);
DFFARX1 I_7(I9864,I1470,I9491,,,I9468,);
or I_8(I9960,I9771,I9943);
nor I_9(I10681,I9477,I9480);
and I_10(I9943,I9576);
DFFARX1 I_11(I9468,I1470,I10647,,,I11009,);
DFFARX1 I_12(I1470,I9491,,,I9621,);
DFFARX1 I_13(I9960,I1470,I9491,,,I9456,);
nand I_14(I11088,I11009,I10698);
nor I_15(I9864,I9816,I9621);
endmodule


