module tb_test_I5368;
reg [0:8] N;
reg CK, reset;
bit [0:0] output_single;
integer i,f;
test_I5368 U1 (N[0],N[1],N[2],N[3],N[4],N[5],N[6],N[7],N[8],CK, reset,output_single[0]);
initial 
begin
    CK = 0;
end
always #10 CK = ~CK;
initial
begin
  reset = 1;
  #5;
  reset = 0;
end
always @(posedge CK)
begin
f = $fopen("./trojan_detection_data/Simulated_Data_Output/Benchmark_testing1000/I5368.txt","w");
N = 9'b000000000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000000001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000000010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000000011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000000100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000000101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000000110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000000111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000001000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000001001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000001010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000001011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000001100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000001101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000001110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000001111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000010000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000010001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000010010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000010011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000010100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000010101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000010110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000010111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000011000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000011001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000011010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000011011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000011100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000011101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000011110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000011111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000100000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000100001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000100010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000100011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000100100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000100101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000100110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000100111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000101000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000101001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000101010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000101011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000101100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000101101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000101110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000101111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000110000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000110001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000110010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000110011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000110100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000110101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000110110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000110111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000111000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000111001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000111010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000111011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000111100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000111101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000111110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b000111111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001000000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001000001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001000010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001000011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001000100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001000101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001000110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001000111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001001000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001001001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001001010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001001011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001001100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001001101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001001110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001001111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001010000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001010001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001010010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001010011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001010100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001010101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001010110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001010111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001011000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001011001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001011010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001011011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001011100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001011101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001011110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001011111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001100000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001100001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001100010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001100011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001100100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001100101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001100110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001100111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001101000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001101001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001101010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001101011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001101100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001101101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001101110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001101111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001110000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001110001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001110010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001110011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001110100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001110101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001110110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001110111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001111000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001111001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001111010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001111011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001111100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001111101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001111110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b001111111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010000000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010000001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010000010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010000011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010000100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010000101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010000110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010000111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010001000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010001001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010001010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010001011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010001100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010001101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010001110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010001111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010010000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010010001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010010010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010010011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010010100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010010101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010010110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010010111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010011000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010011001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010011010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010011011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010011100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010011101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010011110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010011111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010100000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010100001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010100010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010100011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010100100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010100101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010100110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010100111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010101000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010101001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010101010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010101011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010101100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010101101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010101110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010101111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010110000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010110001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010110010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010110011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010110100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010110101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010110110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010110111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010111000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010111001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010111010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010111011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010111100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010111101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010111110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b010111111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011000000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011000001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011000010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011000011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011000100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011000101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011000110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011000111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011001000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011001001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011001010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011001011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011001100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011001101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011001110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011001111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011010000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011010001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011010010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011010011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011010100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011010101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011010110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011010111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011011000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011011001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011011010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011011011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011011100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011011101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011011110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011011111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011100000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011100001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011100010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011100011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011100100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011100101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011100110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011100111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011101000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011101001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011101010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011101011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011101100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011101101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011101110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011101111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011110000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011110001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011110010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011110011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011110100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011110101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011110110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011110111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011111000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011111001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011111010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011111011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011111100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011111101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011111110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b011111111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100000000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100000001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100000010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100000011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100000100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100000101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100000110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100000111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100001000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100001001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100001010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100001011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100001100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100001101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100001110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100001111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100010000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100010001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100010010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100010011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100010100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100010101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100010110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100010111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100011000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100011001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100011010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100011011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100011100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100011101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100011110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100011111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100100000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100100001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100100010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100100011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100100100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100100101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100100110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100100111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100101000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100101001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100101010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100101011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100101100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100101101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100101110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100101111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100110000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100110001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100110010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100110011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100110100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100110101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100110110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100110111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100111000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100111001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100111010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100111011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100111100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100111101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100111110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b100111111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101000000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101000001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101000010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101000011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101000100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101000101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101000110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101000111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101001000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101001001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101001010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101001011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101001100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101001101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101001110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101001111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101010000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101010001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101010010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101010011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101010100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101010101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101010110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101010111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101011000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101011001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101011010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101011011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101011100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101011101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101011110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101011111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101100000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101100001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101100010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101100011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101100100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101100101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101100110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101100111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101101000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101101001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101101010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101101011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101101100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101101101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101101110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101101111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101110000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101110001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101110010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101110011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101110100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101110101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101110110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101110111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101111000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101111001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101111010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101111011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101111100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101111101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101111110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b101111111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110000000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110000001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110000010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110000011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110000100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110000101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110000110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110000111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110001000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110001001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110001010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110001011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110001100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110001101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110001110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110001111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110010000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110010001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110010010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110010011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110010100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110010101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110010110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110010111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110011000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110011001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110011010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110011011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110011100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110011101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110011110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110011111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110100000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110100001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110100010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110100011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110100100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110100101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110100110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110100111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110101000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110101001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110101010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110101011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110101100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110101101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110101110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110101111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110110000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110110001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110110010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110110011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110110100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110110101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110110110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110110111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110111000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110111001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110111010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110111011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110111100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110111101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110111110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b110111111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111000000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111000001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111000010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111000011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111000100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111000101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111000110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111000111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111001000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111001001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111001010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111001011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111001100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111001101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111001110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111001111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111010000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111010001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111010010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111010011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111010100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111010101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111010110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111010111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111011000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111011001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111011010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111011011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111011100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111011101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111011110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111011111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111100000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111100001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111100010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111100011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111100100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111100101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111100110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111100111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111101000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111101001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111101010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111101011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111101100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111101101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111101110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111101111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111110000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111110001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111110010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111110011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111110100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111110101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111110110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111110111;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111111000;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111111001;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111111010;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111111011;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111111100;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111111101;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111111110;
#10
$fwrite(f,"%b %b\n",N,output_single);
N = 9'b111111111;
#10
$fwrite(f,"%b %b\n",N,output_single);
$fclose(f);
$finish;
end
endmodule