module test_I1733(I1367,I1439,I1207,I1733);
input I1367,I1439,I1207;
output I1733;
wire I1716,I1699;
nor I_0(I1716,I1699,I1367);
and I_1(I1733,I1716,I1439);
not I_2(I1699,I1207);
endmodule


