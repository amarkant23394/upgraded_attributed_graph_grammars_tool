module test_final(IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_5_r_11,blif_reset_net_5_r_11,N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11);
input IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_5_r_11,blif_reset_net_5_r_11;
output N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11;
wire N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_102_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13,n4_7_l_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13,n_102_5_r_11,N1372_10_r_11,n_431_5_r_11,n9_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11;
nor I_0(N1371_0_r_13,n59_13,n61_13);
nor I_1(N1508_0_r_13,n59_13,n60_13);
not I_2(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_3(n_431_5_r_13,blif_clk_net_5_r_11,n9_11,G78_5_r_13,);
nand I_4(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_5(n_102_5_r_13,IN_9_7_l_13,IN_10_7_l_13);
nand I_6(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_7(n1_13,blif_clk_net_5_r_11,n9_11,G42_7_r_13,);
nor I_8(n_572_7_r_13,n40_13,n41_13);
nand I_9(n_573_7_r_13,n37_13,n38_13);
nor I_10(n_549_7_r_13,n46_13,n47_13);
nand I_11(n_569_7_r_13,n37_13,n43_13);
nand I_12(n_452_7_r_13,n52_13,n53_13);
nor I_13(n4_7_l_13,G18_7_l_13,IN_1_7_l_13);
DFFARX1 I_14(n4_7_l_13,blif_clk_net_5_r_11,n9_11,n62_13,);
not I_15(n33_13,n62_13);
nand I_16(n_431_5_r_13,n54_13,n55_13);
not I_17(n1_13,n52_13);
nor I_18(n34_13,n35_13,n36_13);
nor I_19(n35_13,G15_7_l_13,n42_13);
nand I_20(n36_13,n50_13,n58_13);
nand I_21(n37_13,n44_13,n45_13);
or I_22(n38_13,IN_3_1_l_13,n39_13);
nand I_23(n39_13,IN_1_1_l_13,IN_2_1_l_13);
not I_24(n40_13,n36_13);
nor I_25(n41_13,IN_10_7_l_13,n35_13);
not I_26(n42_13,IN_4_7_l_13);
or I_27(n43_13,G18_7_l_13,IN_5_7_l_13);
not I_28(n44_13,G15_7_l_13);
not I_29(n45_13,IN_7_7_l_13);
nor I_30(n46_13,n39_13,n40_13);
nor I_31(n47_13,G18_7_l_13,IN_5_7_l_13);
nor I_32(n48_13,n50_13,n51_13);
nor I_33(n49_13,G15_7_l_13,IN_7_7_l_13);
not I_34(n50_13,n59_13);
not I_35(n51_13,n_102_5_r_13);
nand I_36(n52_13,n33_13,n39_13);
nand I_37(n53_13,IN_3_1_l_13,n33_13);
nor I_38(n54_13,IN_5_7_l_13,IN_9_7_l_13);
nand I_39(n55_13,n62_13,n56_13);
nor I_40(n56_13,n39_13,n57_13);
not I_41(n57_13,G18_7_l_13);
or I_42(n58_13,IN_3_10_l_13,IN_4_10_l_13);
nand I_43(n59_13,IN_1_10_l_13,IN_2_10_l_13);
nor I_44(n60_13,IN_5_7_l_13,n51_13);
nor I_45(n61_13,IN_3_1_l_13,n39_13);
not I_46(N1372_1_r_11,n53_11);
nor I_47(N1508_1_r_11,n39_11,n53_11);
nor I_48(N6147_2_r_11,n48_11,n49_11);
nor I_49(N6147_3_r_11,n44_11,n45_11);
nand I_50(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_51(n_431_5_r_11,blif_clk_net_5_r_11,n9_11,G78_5_r_11,);
nand I_52(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_53(n_102_5_r_11,n39_11);
nand I_54(n_547_5_r_11,n36_11,n37_11);
nor I_55(N1507_6_r_11,n52_11,n57_11);
nor I_56(N1508_6_r_11,n46_11,n51_11);
nor I_57(N1372_10_r_11,n43_11,n47_11);
nor I_58(N1508_10_r_11,n55_11,n56_11);
nand I_59(n_431_5_r_11,n40_11,n41_11);
not I_60(n9_11,blif_reset_net_5_r_11);
nor I_61(n36_11,n38_11,n39_11);
not I_62(n37_11,n40_11);
nor I_63(n38_11,n60_11,N1508_0_r_13);
nor I_64(n39_11,n54_11,n_573_7_r_13);
nand I_65(n40_11,N1371_0_r_13,n_429_or_0_5_r_13);
nand I_66(n41_11,n_102_5_r_11,n42_11);
and I_67(n42_11,n58_11,n_547_5_r_13);
not I_68(n43_11,n44_11);
nor I_69(n44_11,n40_11,G42_7_r_13);
nand I_70(n45_11,n46_11,n47_11);
not I_71(n46_11,n38_11);
nand I_72(n47_11,n59_11,n62_11);
and I_73(n48_11,n37_11,n47_11);
or I_74(n49_11,n44_11,n50_11);
nor I_75(n50_11,n60_11,n61_11);
or I_76(n51_11,n_102_5_r_11,n52_11);
nor I_77(n52_11,n42_11,n57_11);
nand I_78(n53_11,n37_11,n50_11);
or I_79(n54_11,n_576_5_r_13,N1508_0_r_13);
nor I_80(n55_11,n38_11,n42_11);
not I_81(n56_11,N1372_10_r_11);
and I_82(n57_11,n38_11,n50_11);
and I_83(n58_11,n59_11,n_572_7_r_13);
or I_84(n59_11,n63_11,G78_5_r_13);
not I_85(n60_11,n_569_7_r_13);
nor I_86(n61_11,N1371_0_r_13,n_452_7_r_13);
nand I_87(n62_11,n_429_or_0_5_r_13,n_549_7_r_13);
and I_88(n63_11,n_429_or_0_5_r_13,n_549_7_r_13);
endmodule


