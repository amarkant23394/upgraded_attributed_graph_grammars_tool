module test_I17205(I12605,I1477,I1470,I17205);
input I12605,I1477,I1470;
output I17205;
wire I14927,I16818,I14965,I15485,I15502;
DFFARX1 I_0(I15502,I1470,I14965,,,I14927,);
DFFARX1 I_1(I14927,I1470,I16818,,,I17205,);
not I_2(I16818,I1477);
not I_3(I14965,I1477);
DFFARX1 I_4(I12605,I1470,I14965,,,I15485,);
not I_5(I15502,I15485);
endmodule


