module test_I9114(I7026,I6975,I7427,I5097,I9114);
input I7026,I6975,I7427,I5097;
output I9114;
wire I8879,I7057,I7317,I6881,I9083,I6887,I6992;
not I_0(I8879,I6887);
not I_1(I7057,I7026);
nor I_2(I7317,I7057);
nand I_3(I6881,I6992,I7057);
nand I_4(I9083,I8879,I6881);
nand I_5(I6887,I7427,I7317);
nand I_6(I6992,I6975,I5097);
not I_7(I9114,I9083);
endmodule


