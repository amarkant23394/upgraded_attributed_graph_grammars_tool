module test_I17775(I1477,I13746,I1470,I13758,I15679,I17775);
input I1477,I13746,I1470,I13758,I15679;
output I17775;
wire I13752,I17413,I15696,I16052,I15585,I15611,I15959,I15928,I16069;
DFFARX1 I_0(I1470,,,I13752,);
not I_1(I17413,I1477);
nand I_2(I15696,I15679,I13758);
DFFARX1 I_3(I15585,I1470,I17413,,,I17775,);
DFFARX1 I_4(I13752,I1470,I15611,,,I16052,);
nand I_5(I15585,I16069,I15959);
not I_6(I15611,I1477);
nor I_7(I15959,I15928,I15696);
DFFARX1 I_8(I13746,I1470,I15611,,,I15928,);
not I_9(I16069,I16052);
endmodule


