module test_I3353(I1668,I1383,I1477,I1603,I1470,I1535,I1207,I3353);
input I1668,I1383,I1477,I1603,I1470,I1535,I1207;
output I3353;
wire I1518,I3388,I1486,I3620,I3637,I1880,I1501,I3453,I1832,I1492,I1483;
not I_0(I1518,I1477);
not I_1(I3388,I1477);
DFFARX1 I_2(I1832,I1470,I1518,,,I1486,);
nor I_3(I3620,I1492,I1483);
and I_4(I3353,I3453,I3637);
DFFARX1 I_5(I3620,I1470,I3388,,,I3637,);
DFFARX1 I_6(I1383,I1470,I1518,,,I1880,);
not I_7(I1501,I1880);
nor I_8(I3453,I1486,I1501);
nand I_9(I1832,I1535,I1207);
nand I_10(I1492,I1603,I1668);
DFFARX1 I_11(I1880,I1470,I1518,,,I1483,);
endmodule


