module test_I2345(I1477,I1470,I1375,I2345);
input I1477,I1470,I1375;
output I2345;
wire I2181;
not I_0(I2181,I1477);
DFFARX1 I_1(I1375,I1470,I2181,,,I2345,);
endmodule


