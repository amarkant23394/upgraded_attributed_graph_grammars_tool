module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_5_r_13,blif_reset_net_5_r_13,N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13);
input IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_5_r_13,blif_reset_net_5_r_13;
output N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13;
wire N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14,I_BUFF_1_9_r_14,N3_8_l_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14,n_102_5_r_13,n4_7_l_13,n9_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13;
nor I_0(N1371_0_r_14,n47_14,n30_14);
nor I_1(N1508_0_r_14,n30_14,n41_14);
nor I_2(N1507_6_r_14,n37_14,n44_14);
nor I_3(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_4(n4_7_r_14,blif_clk_net_5_r_13,n9_13,G42_7_r_14,);
nor I_5(n_572_7_r_14,n28_14,n29_14);
nand I_6(n_573_7_r_14,n26_14,n27_14);
nor I_7(n_549_7_r_14,n31_14,n32_14);
nand I_8(n_569_7_r_14,n26_14,n30_14);
nor I_9(n_452_7_r_14,n47_14,n28_14);
nor I_10(N6147_9_r_14,n36_14,n37_14);
nor I_11(N6134_9_r_14,n28_14,n36_14);
not I_12(I_BUFF_1_9_r_14,n26_14);
and I_13(N3_8_l_14,IN_6_8_l_14,n38_14);
DFFARX1 I_14(N3_8_l_14,blif_clk_net_5_r_13,n9_13,n47_14,);
nor I_15(n4_7_r_14,n47_14,n35_14);
nand I_16(n26_14,IN_1_10_l_14,IN_2_10_l_14);
not I_17(n27_14,n28_14);
nor I_18(n28_14,IN_2_0_l_14,n43_14);
not I_19(n29_14,n33_14);
not I_20(n30_14,n31_14);
nor I_21(n31_14,IN_1_3_l_14,n46_14);
and I_22(n32_14,n33_14,n34_14);
nand I_23(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_24(n34_14,n42_14,n43_14);
nor I_25(n35_14,IN_1_8_l_14,IN_3_8_l_14);
nor I_26(n36_14,n47_14,n34_14);
not I_27(n37_14,n35_14);
nand I_28(n38_14,IN_2_8_l_14,IN_3_8_l_14);
nand I_29(n39_14,n29_14,n40_14);
nand I_30(n40_14,n27_14,n37_14);
nor I_31(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_32(n42_14,IN_3_0_l_14,IN_4_0_l_14);
not I_33(n43_14,IN_1_0_l_14);
nor I_34(n44_14,n27_14,n33_14);
or I_35(n45_14,IN_3_10_l_14,IN_4_10_l_14);
or I_36(n46_14,IN_2_3_l_14,IN_3_3_l_14);
nor I_37(N1371_0_r_13,n59_13,n61_13);
nor I_38(N1508_0_r_13,n59_13,n60_13);
not I_39(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_40(n_431_5_r_13,blif_clk_net_5_r_13,n9_13,G78_5_r_13,);
nand I_41(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_42(n_102_5_r_13,n_572_7_r_14,N1371_0_r_14);
nand I_43(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_44(n1_13,blif_clk_net_5_r_13,n9_13,G42_7_r_13,);
nor I_45(n_572_7_r_13,n40_13,n41_13);
nand I_46(n_573_7_r_13,n37_13,n38_13);
nor I_47(n_549_7_r_13,n46_13,n47_13);
nand I_48(n_569_7_r_13,n37_13,n43_13);
nand I_49(n_452_7_r_13,n52_13,n53_13);
nor I_50(n4_7_l_13,G42_7_r_14,n_573_7_r_14);
not I_51(n9_13,blif_reset_net_5_r_13);
DFFARX1 I_52(n4_7_l_13,blif_clk_net_5_r_13,n9_13,n62_13,);
not I_53(n33_13,n62_13);
nand I_54(n_431_5_r_13,n54_13,n55_13);
not I_55(n1_13,n52_13);
nor I_56(n34_13,n35_13,n36_13);
nor I_57(n35_13,n42_13,N6134_9_r_14);
nand I_58(n36_13,n50_13,n58_13);
nand I_59(n37_13,n44_13,n45_13);
or I_60(n38_13,n39_13,N1508_0_r_14);
nand I_61(n39_13,N1371_0_r_14,N1507_6_r_14);
not I_62(n40_13,n36_13);
nor I_63(n41_13,n35_13,n_572_7_r_14);
not I_64(n42_13,n_569_7_r_14);
or I_65(n43_13,n_573_7_r_14,N6147_9_r_14);
not I_66(n44_13,N6134_9_r_14);
not I_67(n45_13,N1508_6_r_14);
nor I_68(n46_13,n39_13,n40_13);
nor I_69(n47_13,n_573_7_r_14,N6147_9_r_14);
nor I_70(n48_13,n50_13,n51_13);
nor I_71(n49_13,N1508_6_r_14,N6134_9_r_14);
not I_72(n50_13,n59_13);
not I_73(n51_13,n_102_5_r_13);
nand I_74(n52_13,n33_13,n39_13);
nand I_75(n53_13,n33_13,N1508_0_r_14);
nor I_76(n54_13,N6147_9_r_14,N1371_0_r_14);
nand I_77(n55_13,n62_13,n56_13);
nor I_78(n56_13,n39_13,n57_13);
not I_79(n57_13,n_573_7_r_14);
or I_80(n58_13,N1508_0_r_14,n_549_7_r_14);
nand I_81(n59_13,n_452_7_r_14,N1507_6_r_14);
nor I_82(n60_13,n51_13,N6147_9_r_14);
nor I_83(n61_13,n39_13,N1508_0_r_14);
endmodule


