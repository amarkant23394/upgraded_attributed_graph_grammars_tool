module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_5_r_7,blif_reset_net_5_r_7,N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7);
input IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_5_r_7,blif_reset_net_5_r_7;
output N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7;
wire N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_102_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1372_10_r_11,N1508_10_r_11,n_431_5_r_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11,n_102_5_r_7,n_452_7_r_7,n4_7_l_7,n6_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7;
not I_0(N1372_1_r_11,n53_11);
nor I_1(N1508_1_r_11,n39_11,n53_11);
nor I_2(N6147_2_r_11,n48_11,n49_11);
nor I_3(N6147_3_r_11,n44_11,n45_11);
nand I_4(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_5(n_431_5_r_11,blif_clk_net_5_r_7,n6_7,G78_5_r_11,);
nand I_6(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_7(n_102_5_r_11,n39_11);
nand I_8(n_547_5_r_11,n36_11,n37_11);
nor I_9(N1507_6_r_11,n52_11,n57_11);
nor I_10(N1508_6_r_11,n46_11,n51_11);
nor I_11(N1372_10_r_11,n43_11,n47_11);
nor I_12(N1508_10_r_11,n55_11,n56_11);
nand I_13(n_431_5_r_11,n40_11,n41_11);
nor I_14(n36_11,n38_11,n39_11);
not I_15(n37_11,n40_11);
nor I_16(n38_11,IN_2_0_l_11,n60_11);
nor I_17(n39_11,IN_1_3_l_11,n54_11);
nand I_18(n40_11,IN_1_1_l_11,IN_2_1_l_11);
nand I_19(n41_11,n_102_5_r_11,n42_11);
and I_20(n42_11,IN_2_6_l_11,n58_11);
not I_21(n43_11,n44_11);
nor I_22(n44_11,IN_3_1_l_11,n40_11);
nand I_23(n45_11,n46_11,n47_11);
not I_24(n46_11,n38_11);
nand I_25(n47_11,n59_11,n62_11);
and I_26(n48_11,n37_11,n47_11);
or I_27(n49_11,n44_11,n50_11);
nor I_28(n50_11,n60_11,n61_11);
or I_29(n51_11,n_102_5_r_11,n52_11);
nor I_30(n52_11,n42_11,n57_11);
nand I_31(n53_11,n37_11,n50_11);
or I_32(n54_11,IN_2_3_l_11,IN_3_3_l_11);
nor I_33(n55_11,n38_11,n42_11);
not I_34(n56_11,N1372_10_r_11);
and I_35(n57_11,n38_11,n50_11);
and I_36(n58_11,IN_1_6_l_11,n59_11);
or I_37(n59_11,IN_5_6_l_11,n63_11);
not I_38(n60_11,IN_1_0_l_11);
nor I_39(n61_11,IN_3_0_l_11,IN_4_0_l_11);
nand I_40(n62_11,IN_3_6_l_11,IN_4_6_l_11);
and I_41(n63_11,IN_3_6_l_11,IN_4_6_l_11);
nor I_42(N1371_0_r_7,n53_7,n52_7);
nor I_43(N1508_0_r_7,n51_7,n52_7);
nand I_44(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_45(n_431_5_r_7,blif_clk_net_5_r_7,n6_7,G78_5_r_7,);
nand I_46(n_576_5_r_7,n31_7,n32_7);
nor I_47(n_102_5_r_7,N1508_1_r_11,N1508_10_r_11);
nand I_48(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_49(n4_7_r_7,blif_clk_net_5_r_7,n6_7,G42_7_r_7,);
nor I_50(n_572_7_r_7,n54_7,n33_7);
nand I_51(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_52(n_549_7_r_7,n53_7,n36_7);
nand I_53(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_54(n_452_7_r_7,n_576_5_r_11,n_547_5_r_11);
nor I_55(n4_7_l_7,N1372_1_r_11,N6147_2_r_11);
not I_56(n6_7,blif_reset_net_5_r_7);
DFFARX1 I_57(n4_7_l_7,blif_clk_net_5_r_7,n6_7,n53_7,);
not I_58(n30_7,n53_7);
and I_59(N3_8_l_7,n50_7,N1372_1_r_11);
DFFARX1 I_60(N3_8_l_7,blif_clk_net_5_r_7,n6_7,n54_7,);
nand I_61(n_431_5_r_7,n40_7,n41_7);
nor I_62(n4_7_r_7,n54_7,n49_7);
and I_63(n31_7,n_102_5_r_7,n39_7);
not I_64(n32_7,N1372_1_r_11);
nor I_65(n33_7,n34_7,N1508_6_r_11);
and I_66(n34_7,n35_7,N6147_3_r_11);
not I_67(n35_7,n_429_or_0_5_r_11);
nor I_68(n36_7,n37_7,N1372_1_r_11);
or I_69(n37_7,n54_7,N1508_10_r_11);
or I_70(n38_7,N6147_2_r_11,N1507_6_r_11);
nor I_71(n39_7,n_452_7_r_7,N1508_1_r_11);
nand I_72(n40_7,n46_7,n47_7);
nand I_73(n41_7,n42_7,n43_7);
nor I_74(n42_7,n44_7,n45_7);
nor I_75(n43_7,N6147_2_r_11,N1507_6_r_11);
nor I_76(n44_7,n_429_or_0_5_r_11,G78_5_r_11);
nor I_77(n45_7,N1508_1_r_11,N1508_6_r_11);
nand I_78(n46_7,n35_7,N6147_3_r_11);
not I_79(n47_7,N1508_6_r_11);
or I_80(n48_7,n_452_7_r_7,N1508_1_r_11);
not I_81(n49_7,n_452_7_r_7);
nand I_82(n50_7,N6147_3_r_11,N1507_6_r_11);
and I_83(n51_7,n_452_7_r_7,n45_7);
not I_84(n52_7,n44_7);
endmodule


