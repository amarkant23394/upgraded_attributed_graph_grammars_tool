module test_I1954(I1376,I1263,I1294,I1639,I1301,I1954);
input I1376,I1263,I1294,I1639,I1301;
output I1954;
wire I1704,I1322,I1342,I1427,I1393,I1687;
nor I_0(I1704,I1393,I1687);
nand I_1(I1322,I1427,I1704);
not I_2(I1342,I1301);
DFFARX1 I_3(I1263,I1294,I1342,,,I1427,);
not I_4(I1954,I1322);
DFFARX1 I_5(I1376,I1294,I1342,,,I1393,);
not I_6(I1687,I1639);
endmodule


