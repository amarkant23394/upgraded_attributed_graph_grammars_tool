module test_final(IN_1_2_l_1,IN_2_2_l_1,G1_3_l_1,G2_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_5_3_l_1,IN_7_3_l_1,IN_8_3_l_1,IN_10_3_l_1,IN_11_3_l_1,blif_reset_net_0_r_4,blif_clk_net_0_r_4,ACVQN2_0_r_4,n_266_and_0_0_r_4,ACVQN1_2_r_4,P6_2_r_4,n_429_or_0_3_r_4,G78_3_r_4,n_576_3_r_4,n_102_3_r_4,n_547_3_r_4,n_42_5_r_4,G199_5_r_4);
input IN_1_2_l_1,IN_2_2_l_1,G1_3_l_1,G2_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_5_3_l_1,IN_7_3_l_1,IN_8_3_l_1,IN_10_3_l_1,IN_11_3_l_1,blif_reset_net_0_r_4,blif_clk_net_0_r_4;
output ACVQN2_0_r_4,n_266_and_0_0_r_4,ACVQN1_2_r_4,P6_2_r_4,n_429_or_0_3_r_4,G78_3_r_4,n_576_3_r_4,n_102_3_r_4,n_547_3_r_4,n_42_5_r_4,G199_5_r_4;
wire ACVQN2_0_r_1,n_266_and_0_0_r_1,G199_1_r_1,G214_1_r_1,ACVQN1_2_r_1,P6_2_r_1,n_429_or_0_3_r_1,G78_3_r_1,n_576_3_r_1,n_102_3_r_1,n_547_3_r_1,ACVQN1_2_l_1,P6_2_l_1,P6_internal_2_l_1,n_429_or_0_3_l_1,n12_3_l_1,n_431_3_l_1,G78_3_l_1,n_576_3_l_1,n11_3_l_1,n_102_3_l_1,n_547_3_l_1,n13_3_l_1,n14_3_l_1,n15_3_l_1,n16_3_l_1,ACVQN1_0_r_1,N1_1_r_1,n3_1_r_1,P6_internal_2_r_1,n12_3_r_1,n_431_3_r_1,n11_3_r_1,n13_3_r_1,n14_3_r_1,n15_3_r_1,n16_3_r_1,n1_0_r_4,ACVQN2_0_l_4,n_266_and_0_0_l_4,ACVQN1_0_l_4,n4_4_l_4,G42_4_l_4,n_87_4_l_4,n_572_4_l_4,n_573_4_l_4,n_549_4_l_4,n7_4_l_4,n_569_4_l_4,n_452_4_l_4,ACVQN1_0_r_4,P6_internal_2_r_4,n12_3_r_4,n_431_3_r_4,n11_3_r_4,n13_3_r_4,n14_3_r_4,n15_3_r_4,n16_3_r_4,N3_5_r_4,n3_5_r_4;
DFFARX1 I_0(P6_2_l_1,blif_clk_net_0_r_4,n1_0_r_4,ACVQN2_0_r_1,);
and I_1(n_266_and_0_0_r_1,n_102_3_l_1,ACVQN1_0_r_1);
DFFARX1 I_2(N1_1_r_1,blif_clk_net_0_r_4,n1_0_r_4,G199_1_r_1,);
DFFARX1 I_3(n_576_3_l_1,blif_clk_net_0_r_4,n1_0_r_4,G214_1_r_1,);
DFFARX1 I_4(n_547_3_l_1,blif_clk_net_0_r_4,n1_0_r_4,ACVQN1_2_r_1,);
not I_5(P6_2_r_1,P6_internal_2_r_1);
nand I_6(n_429_or_0_3_r_1,ACVQN1_2_l_1,n12_3_r_1);
DFFARX1 I_7(n_431_3_r_1,blif_clk_net_0_r_4,n1_0_r_4,G78_3_r_1,);
nand I_8(n_576_3_r_1,n_547_3_l_1,n11_3_r_1);
not I_9(n_102_3_r_1,n_576_3_l_1);
nand I_10(n_547_3_r_1,P6_2_l_1,n13_3_r_1);
DFFARX1 I_11(IN_2_2_l_1,blif_clk_net_0_r_4,n1_0_r_4,ACVQN1_2_l_1,);
not I_12(P6_2_l_1,P6_internal_2_l_1);
DFFARX1 I_13(IN_1_2_l_1,blif_clk_net_0_r_4,n1_0_r_4,P6_internal_2_l_1,);
nand I_14(n_429_or_0_3_l_1,G1_3_l_1,n12_3_l_1);
not I_15(n12_3_l_1,IN_5_3_l_1);
or I_16(n_431_3_l_1,IN_8_3_l_1,n14_3_l_1);
DFFARX1 I_17(n_431_3_l_1,blif_clk_net_0_r_4,n1_0_r_4,G78_3_l_1,);
nand I_18(n_576_3_l_1,IN_7_3_l_1,n11_3_l_1);
nor I_19(n11_3_l_1,G2_3_l_1,n12_3_l_1);
not I_20(n_102_3_l_1,G2_3_l_1);
nand I_21(n_547_3_l_1,IN_11_3_l_1,n13_3_l_1);
nor I_22(n13_3_l_1,G2_3_l_1,IN_10_3_l_1);
and I_23(n14_3_l_1,IN_2_3_l_1,n15_3_l_1);
nor I_24(n15_3_l_1,IN_4_3_l_1,n16_3_l_1);
not I_25(n16_3_l_1,G1_3_l_1);
DFFARX1 I_26(n_429_or_0_3_l_1,blif_clk_net_0_r_4,n1_0_r_4,ACVQN1_0_r_1,);
and I_27(N1_1_r_1,n_429_or_0_3_l_1,n3_1_r_1);
nand I_28(n3_1_r_1,n_429_or_0_3_l_1,G78_3_l_1);
DFFARX1 I_29(ACVQN1_2_l_1,blif_clk_net_0_r_4,n1_0_r_4,P6_internal_2_r_1,);
not I_30(n12_3_r_1,n_102_3_l_1);
or I_31(n_431_3_r_1,P6_2_l_1,n14_3_r_1);
nor I_32(n11_3_r_1,G78_3_l_1,n12_3_r_1);
nor I_33(n13_3_r_1,G78_3_l_1,n_576_3_l_1);
and I_34(n14_3_r_1,ACVQN1_2_l_1,n15_3_r_1);
nor I_35(n15_3_r_1,n_576_3_l_1,n16_3_r_1);
not I_36(n16_3_r_1,ACVQN1_2_l_1);
DFFARX1 I_37(n_569_4_l_4,blif_clk_net_0_r_4,n1_0_r_4,ACVQN2_0_r_4,);
and I_38(n_266_and_0_0_r_4,ACVQN2_0_l_4,ACVQN1_0_r_4);
DFFARX1 I_39(n_266_and_0_0_l_4,blif_clk_net_0_r_4,n1_0_r_4,ACVQN1_2_r_4,);
not I_40(P6_2_r_4,P6_internal_2_r_4);
nand I_41(n_429_or_0_3_r_4,G42_4_l_4,n12_3_r_4);
DFFARX1 I_42(n_431_3_r_4,blif_clk_net_0_r_4,n1_0_r_4,G78_3_r_4,);
nand I_43(n_576_3_r_4,n_573_4_l_4,n11_3_r_4);
not I_44(n_102_3_r_4,n_569_4_l_4);
nand I_45(n_547_3_r_4,ACVQN2_0_l_4,n13_3_r_4);
nor I_46(n_42_5_r_4,G42_4_l_4,n_549_4_l_4);
DFFARX1 I_47(N3_5_r_4,blif_clk_net_0_r_4,n1_0_r_4,G199_5_r_4,);
not I_48(n1_0_r_4,blif_reset_net_0_r_4);
DFFARX1 I_49(n_576_3_r_1,blif_clk_net_0_r_4,n1_0_r_4,ACVQN2_0_l_4,);
and I_50(n_266_and_0_0_l_4,ACVQN1_0_l_4,ACVQN1_2_r_1);
DFFARX1 I_51(G199_1_r_1,blif_clk_net_0_r_4,n1_0_r_4,ACVQN1_0_l_4,);
nor I_52(n4_4_l_4,n_266_and_0_0_r_1,n_547_3_r_1);
DFFARX1 I_53(n4_4_l_4,blif_clk_net_0_r_4,n1_0_r_4,G42_4_l_4,);
not I_54(n_87_4_l_4,n_102_3_r_1);
nor I_55(n_572_4_l_4,ACVQN2_0_r_1,n_102_3_r_1);
or I_56(n_573_4_l_4,G214_1_r_1,n_429_or_0_3_r_1);
nor I_57(n_549_4_l_4,n7_4_l_4,P6_2_r_1);
and I_58(n7_4_l_4,n_87_4_l_4,G78_3_r_1);
or I_59(n_569_4_l_4,P6_2_r_1,n_429_or_0_3_r_1);
nor I_60(n_452_4_l_4,n_266_and_0_0_r_1,G214_1_r_1);
DFFARX1 I_61(n_549_4_l_4,blif_clk_net_0_r_4,n1_0_r_4,ACVQN1_0_r_4,);
DFFARX1 I_62(ACVQN2_0_l_4,blif_clk_net_0_r_4,n1_0_r_4,P6_internal_2_r_4,);
not I_63(n12_3_r_4,n_266_and_0_0_l_4);
or I_64(n_431_3_r_4,n_572_4_l_4,n14_3_r_4);
nor I_65(n11_3_r_4,n_569_4_l_4,n12_3_r_4);
nor I_66(n13_3_r_4,n_572_4_l_4,n_569_4_l_4);
and I_67(n14_3_r_4,n_452_4_l_4,n15_3_r_4);
nor I_68(n15_3_r_4,n_266_and_0_0_l_4,n16_3_r_4);
not I_69(n16_3_r_4,G42_4_l_4);
and I_70(N3_5_r_4,n_573_4_l_4,n3_5_r_4);
nand I_71(n3_5_r_4,n_549_4_l_4,n_452_4_l_4);
endmodule


