module test_I17498(I13908,I1477,I15662,I15781,I16145,I15696,I1470,I15976,I17498);
input I13908,I1477,I15662,I15781,I16145,I15696,I1470,I15976;
output I17498;
wire I13749,I13743,I15600,I15832,I15815,I15579,I15611,I15597,I16162,I17430,I13767,I14162,I15628,I17481,I15798;
nand I_0(I13749,I14162,I13908);
DFFARX1 I_1(I1470,,,I13743,);
or I_2(I15600,I15832,I15815);
nand I_3(I15832,I15628,I13749);
DFFARX1 I_4(I15798,I1470,I15611,,,I15815,);
nand I_5(I15579,I15662,I15976);
not I_6(I15611,I1477);
nand I_7(I17498,I17481,I15600);
nor I_8(I15597,I15832,I16162);
and I_9(I16162,I15696,I16145);
not I_10(I17430,I15579);
DFFARX1 I_11(I1470,,,I13767,);
DFFARX1 I_12(I1470,,,I14162,);
not I_13(I15628,I13743);
nor I_14(I17481,I17430,I15597);
or I_15(I15798,I15781,I13767);
endmodule


