module test_I8208(I5728,I8233,I8428,I1477,I1470,I5881,I8208);
input I5728,I8233,I8428,I1477,I1470,I5881;
output I8208;
wire I8479,I8216,I8753,I8445,I5915,I5802,I8298,I5719,I5740,I5731,I8315,I8736,I8462;
nor I_0(I8479,I8462,I8315);
not I_1(I8216,I1477);
not I_2(I8753,I8736);
or I_3(I8445,I8428,I5728);
DFFARX1 I_4(I1470,,,I5915,);
DFFARX1 I_5(I1470,,,I5802,);
nor I_6(I8298,I8233,I5719);
DFFARX1 I_7(I1470,,,I5719,);
not I_8(I5740,I5802);
nand I_9(I5731,I5915,I5881);
nand I_10(I8315,I8298,I5740);
DFFARX1 I_11(I5731,I1470,I8216,,,I8736,);
DFFARX1 I_12(I8445,I1470,I8216,,,I8462,);
nand I_13(I8208,I8753,I8479);
endmodule


