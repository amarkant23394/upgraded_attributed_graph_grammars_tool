module test_I17387(I15628,I15579,I13749,I1470,I15611,I16162,I15798,I17387);
input I15628,I15579,I13749,I1470,I15611,I16162,I15798;
output I17387;
wire I17563,I17430,I15597,I15600,I17532,I15832,I15815,I17481,I17498;
not I_0(I17563,I17532);
not I_1(I17430,I15579);
nand I_2(I17387,I17498,I17563);
nor I_3(I15597,I15832,I16162);
or I_4(I15600,I15832,I15815);
not I_5(I17532,I15597);
nand I_6(I15832,I15628,I13749);
DFFARX1 I_7(I15798,I1470,I15611,,,I15815,);
nor I_8(I17481,I17430,I15597);
nand I_9(I17498,I17481,I15600);
endmodule


