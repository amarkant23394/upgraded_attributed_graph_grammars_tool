module test_I14930(I12718,I1477,I1470,I12964,I12653,I14930);
input I12718,I1477,I1470,I12964,I12653;
output I14930;
wire I12619,I12670,I12584,I12783,I15109,I14982,I12596,I15276,I12599,I12735,I14965,I15341;
not I_0(I12619,I1477);
DFFARX1 I_1(I12653,I1470,I12619,,,I12670,);
and I_2(I14930,I15109,I15341);
and I_3(I12584,I12670,I12783);
DFFARX1 I_4(I12735,I1470,I12619,,,I12783,);
not I_5(I15109,I12584);
not I_6(I14982,I12596);
DFFARX1 I_7(I1470,I12619,,,I12596,);
nand I_8(I15276,I14982,I12599);
nand I_9(I12599,I12718,I12964);
DFFARX1 I_10(I1470,I12619,,,I12735,);
not I_11(I14965,I1477);
DFFARX1 I_12(I15276,I1470,I14965,,,I15341,);
endmodule


