module test_I5105(I1477,I5105);
input I1477;
output I5105;
wire ;
not I_0(I5105,I1477);
endmodule


