module test_I10896(I8202,I8181,I9720,I1477,I1470,I10828,I10896);
input I8202,I8181,I9720,I1477,I1470,I10828;
output I10896;
wire I10879,I10647,I9462,I9576,I10862,I9816,I9483,I10845,I9453;
or I_0(I10879,I10862,I9462);
not I_1(I10647,I1477);
not I_2(I9462,I9576);
nor I_3(I9576,I8181,I8202);
and I_4(I10862,I10845,I9453);
DFFARX1 I_5(I1470,,,I9816,);
nor I_6(I9483,I9816);
nor I_7(I10845,I10828,I9483);
DFFARX1 I_8(I10879,I1470,I10647,,,I10896,);
nand I_9(I9453,I9816,I9720);
endmodule


