module test_I13296(I8830,I1477,I11830,I1470,I9258,I11395,I13296);
input I8830,I1477,I11830,I1470,I9258,I11395;
output I13296;
wire I8827,I11327,I11302,I11847,I11278,I8862,I11310,I11864,I11624;
DFFARX1 I_0(I9258,I1470,I8862,,,I8827,);
not I_1(I11327,I8830);
DFFARX1 I_2(I11864,I1470,I11310,,,I11302,);
nand I_3(I11847,I11830,I11395);
DFFARX1 I_4(I11624,I1470,I11310,,,I11278,);
not I_5(I8862,I1477);
nor I_6(I13296,I11278,I11302);
not I_7(I11310,I1477);
and I_8(I11864,I11624,I11847);
nand I_9(I11624,I11327,I8827);
endmodule


