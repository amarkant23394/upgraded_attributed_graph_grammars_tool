module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_7_r_1,n9_1,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
and I_35(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_36(N1508_0_r_1,n40_1,n44_1);
nor I_37(N1507_6_r_1,n43_1,n49_1);
nor I_38(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_39(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_40(n_572_7_r_1,n29_1,n30_1);
not I_41(n_573_7_r_1,n_452_7_r_1);
nor I_42(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_43(n_569_7_r_1,n30_1,n31_1);
nor I_44(n_452_7_r_1,n30_1,n32_1);
nor I_45(N6147_9_r_1,n35_1,n36_1);
nand I_46(N6134_9_r_1,n38_1,n39_1);
not I_47(I_BUFF_1_9_r_1,n40_1);
nor I_48(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_49(n9_1,blif_reset_net_7_r_1);
nor I_50(n29_1,n34_1,n_452_7_r_4);
nor I_51(n30_1,n33_1,n34_1);
nor I_52(n31_1,n54_1,G42_7_r_4);
not I_53(n32_1,n48_1);
nor I_54(n33_1,N6134_9_r_4,n_549_7_r_4);
not I_55(n34_1,N1371_0_r_4);
nor I_56(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_57(n36_1,n29_1);
not I_58(n37_1,n41_1);
nand I_59(n38_1,I_BUFF_1_9_r_1,N1371_0_r_4);
nand I_60(n39_1,n37_1,n40_1);
nand I_61(n40_1,N1507_6_r_4,n_549_7_r_4);
nand I_62(n41_1,n52_1,n_572_7_r_4);
or I_63(n42_1,n36_1,n43_1);
nor I_64(n43_1,n32_1,n49_1);
nand I_65(n44_1,n45_1,n46_1);
nand I_66(n45_1,n47_1,n48_1);
not I_67(n46_1,N1371_0_r_4);
not I_68(n47_1,n31_1);
nand I_69(n48_1,n50_1,G42_7_r_4);
nor I_70(n49_1,n41_1,n47_1);
and I_71(n50_1,n51_1,n_569_7_r_4);
nand I_72(n51_1,n52_1,n53_1);
nand I_73(n52_1,N1507_6_r_4,N1508_6_r_4);
not I_74(n53_1,n_572_7_r_4);
or I_75(n54_1,N1508_6_r_4,n_572_7_r_4);
nor I_76(n55_1,n29_1,N1371_0_r_4);
endmodule


