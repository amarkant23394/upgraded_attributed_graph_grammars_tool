module test_I3622(I2600,I1294,I2457,I1301,I3622);
input I2600,I1294,I2457,I1301;
output I3622;
wire I2668,I1914,I2651,I1937,I2039,I1908,I3246,I2702,I2572;
DFFARX1 I_0(I2572,I1294,I3246,,,I3622,);
nand I_1(I2668,I2651,I1914);
DFFARX1 I_2(I2457,I1294,I1937,,,I1914,);
nor I_3(I2651,I2600,I1908);
not I_4(I1937,I1301);
DFFARX1 I_5(I1294,I1937,,,I2039,);
not I_6(I1908,I2039);
not I_7(I3246,I1301);
not I_8(I2702,I1908);
nor I_9(I2572,I2668,I2702);
endmodule


