module test_I13775(I1477,I13775);
input I1477;
output I13775;
wire ;
not I_0(I13775,I1477);
endmodule


