module test_I6899(I5659,I1477,I1470,I5097,I6899);
input I5659,I1477,I1470,I5097;
output I6899;
wire I5105,I5073,I6992,I6975,I7461,I7427,I5088,I6907,I7410,I7221,I6924,I7444;
not I_0(I5105,I1477);
DFFARX1 I_1(I1470,I5105,,,I5073,);
nand I_2(I6992,I6975,I5097);
nor I_3(I6975,I6924);
and I_4(I7461,I7221,I7444);
not I_5(I7427,I7410);
DFFARX1 I_6(I5659,I1470,I5105,,,I5088,);
not I_7(I6907,I1477);
DFFARX1 I_8(I1470,I6907,,,I7410,);
nand I_9(I7221,I6924,I5088);
DFFARX1 I_10(I7461,I1470,I6907,,,I6899,);
not I_11(I6924,I5073);
nand I_12(I7444,I7427,I6992);
endmodule


