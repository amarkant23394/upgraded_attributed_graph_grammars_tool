module test_final(IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_8_r_6,blif_reset_net_8_r_6,N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_8_r_6,blif_reset_net_8_r_6;
output N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_573_7_r_12,n_549_7_r_12,n_569_7_r_12,n_452_7_r_12,N6147_9_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12,I_BUFF_1_9_r_6,N3_8_r_6,n9_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6;
nor I_0(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_1(N1508_0_r_12,n30_12,n37_12);
nor I_2(N1507_6_r_12,n25_12,n39_12);
nor I_3(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_4(n1_12,blif_clk_net_8_r_6,n9_6,G42_7_r_12,);
nor I_5(n_572_7_r_12,n23_12,n24_12);
nand I_6(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_7(n_549_7_r_12,n27_12,n28_12);
nand I_8(n_569_7_r_12,n25_12,n26_12);
nand I_9(n_452_7_r_12,IN_1_1_l_12,IN_2_1_l_12);
nand I_10(N6147_9_r_12,n30_12,n31_12);
nor I_11(N6134_9_r_12,n35_12,n36_12);
not I_12(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_13(n1_12,n_573_7_r_12);
not I_14(n23_12,n36_12);
nor I_15(n24_12,IN_3_1_l_12,n_452_7_r_12);
nand I_16(n25_12,n23_12,n40_12);
not I_17(n26_12,n35_12);
not I_18(n27_12,N6134_9_r_12);
nand I_19(n28_12,n26_12,n29_12);
not I_20(n29_12,n24_12);
nand I_21(n30_12,n33_12,n41_12);
nand I_22(n31_12,n32_12,n33_12);
nor I_23(n32_12,n26_12,n34_12);
nor I_24(n33_12,IN_1_2_l_12,IN_2_2_l_12);
nor I_25(n34_12,IN_5_2_l_12,n42_12);
nor I_26(n35_12,IN_1_3_l_12,n38_12);
nand I_27(n36_12,IN_1_10_l_12,IN_2_10_l_12);
nand I_28(n37_12,n23_12,n35_12);
or I_29(n38_12,IN_2_3_l_12,IN_3_3_l_12);
not I_30(n39_12,n30_12);
or I_31(n40_12,IN_3_10_l_12,IN_4_10_l_12);
nor I_32(n41_12,n34_12,n36_12);
nor I_33(n42_12,IN_3_2_l_12,IN_4_2_l_12);
nor I_34(N1371_0_r_6,n30_6,n33_6);
nor I_35(N1508_0_r_6,n33_6,n44_6);
not I_36(N1372_1_r_6,n41_6);
nor I_37(N1508_1_r_6,n40_6,n41_6);
nor I_38(N1507_6_r_6,n39_6,n45_6);
nor I_39(N1508_6_r_6,n37_6,n38_6);
nor I_40(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_41(N3_8_r_6,blif_clk_net_8_r_6,n9_6,G199_8_r_6,);
nor I_42(N6147_9_r_6,n32_6,n33_6);
nor I_43(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_44(I_BUFF_1_9_r_6,n37_6);
not I_45(N1372_10_r_6,n43_6);
nor I_46(N1508_10_r_6,n42_6,n43_6);
nor I_47(N3_8_r_6,n36_6,N1508_0_r_12);
not I_48(n9_6,blif_reset_net_8_r_6);
nor I_49(n30_6,n53_6,n_572_7_r_12);
not I_50(n31_6,n36_6);
nor I_51(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_52(n33_6,N1508_0_r_12);
not I_53(n34_6,n35_6);
nand I_54(n35_6,n49_6,N1508_0_r_12);
nand I_55(n36_6,n51_6,G42_7_r_12);
nand I_56(n37_6,n54_6,n_569_7_r_12);
or I_57(n38_6,n35_6,n39_6);
nor I_58(n39_6,n40_6,n45_6);
and I_59(n40_6,n46_6,n47_6);
nand I_60(n41_6,n30_6,n31_6);
nor I_61(n42_6,n34_6,n40_6);
nand I_62(n43_6,n30_6,N1508_0_r_12);
nor I_63(n44_6,n31_6,n40_6);
nor I_64(n45_6,n35_6,n36_6);
nor I_65(n46_6,N1371_0_r_12,n_572_7_r_12);
or I_66(n47_6,n48_6,G42_7_r_12);
nor I_67(n48_6,N1507_6_r_12,N6147_9_r_12);
and I_68(n49_6,n50_6,N1507_6_r_12);
nand I_69(n50_6,n51_6,n52_6);
nand I_70(n51_6,n_549_7_r_12,N1508_6_r_12);
not I_71(n52_6,G42_7_r_12);
nor I_72(n53_6,N1508_6_r_12,N1371_0_r_12);
or I_73(n54_6,N1508_6_r_12,N1371_0_r_12);
endmodule


