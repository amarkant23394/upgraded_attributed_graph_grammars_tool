module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_15,blif_reset_net_1_r_15,G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_15,blif_reset_net_1_r_15;
output G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15;
wire G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6,N3_2_l_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6,n_452_1_r_15,n4_1_l_15,n4_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15;
DFFARX1 I_0(n4_1_r_6,blif_clk_net_1_r_15,n4_15,G42_1_r_6,);
nor I_1(n_572_1_r_6,n27_6,n28_6);
nand I_2(n_573_1_r_6,n18_6,n19_6);
nor I_3(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_4(n_569_1_r_6,n19_6,n20_6);
nor I_5(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_6(N1_4_r_6,blif_clk_net_1_r_15,n4_15,G199_4_r_6,);
DFFARX1 I_7(n_42_2_l_6,blif_clk_net_1_r_15,n4_15,G214_4_r_6,);
DFFARX1 I_8(n_42_2_l_6,blif_clk_net_1_r_15,n4_15,ACVQN1_5_r_6,);
not I_9(P6_5_r_6,P6_5_r_internal_6);
and I_10(N3_2_l_6,IN_6_2_l_6,n23_6);
DFFARX1 I_11(N3_2_l_6,blif_clk_net_1_r_15,n4_15,n27_6,);
not I_12(n17_6,n27_6);
DFFARX1 I_13(IN_1_3_l_6,blif_clk_net_1_r_15,n4_15,n28_6,);
DFFARX1 I_14(IN_2_3_l_6,blif_clk_net_1_r_15,n4_15,n26_6,);
and I_15(N1_4_l_6,IN_6_4_l_6,n25_6);
DFFARX1 I_16(N1_4_l_6,blif_clk_net_1_r_15,n4_15,n29_6,);
not I_17(n18_6,n29_6);
DFFARX1 I_18(IN_3_4_l_6,blif_clk_net_1_r_15,n4_15,G214_4_l_6,);
not I_19(n12_6,G214_4_l_6);
nor I_20(n4_1_r_6,n28_6,n22_6);
nor I_21(N1_4_r_6,n12_6,n24_6);
nor I_22(n_42_2_l_6,IN_1_2_l_6,IN_3_2_l_6);
DFFARX1 I_23(G214_4_l_6,blif_clk_net_1_r_15,n4_15,P6_5_r_internal_6,);
nand I_24(n19_6,IN_4_3_l_6,n26_6);
not I_25(n20_6,n_42_2_l_6);
nor I_26(n21_6,n17_6,n28_6);
and I_27(n22_6,IN_4_3_l_6,n26_6);
nand I_28(n23_6,IN_2_2_l_6,IN_3_2_l_6);
nor I_29(n24_6,n17_6,n18_6);
nand I_30(n25_6,IN_1_4_l_6,IN_2_4_l_6);
DFFARX1 I_31(n_452_1_r_15,blif_clk_net_1_r_15,n4_15,G42_1_r_15,);
and I_32(n_572_1_r_15,n17_15,n19_15);
nand I_33(n_573_1_r_15,n15_15,n18_15);
nor I_34(n_549_1_r_15,n21_15,n22_15);
nand I_35(n_569_1_r_15,n15_15,n20_15);
nor I_36(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_37(G42_1_l_15,blif_clk_net_1_r_15,n4_15,ACVQN2_3_r_15,);
nor I_38(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_39(N1_4_r_15,blif_clk_net_1_r_15,n4_15,G199_4_r_15,);
DFFARX1 I_40(n_573_1_l_15,blif_clk_net_1_r_15,n4_15,G214_4_r_15,);
nor I_41(n4_1_l_15,G199_4_r_6,G214_4_r_6);
not I_42(n4_15,blif_reset_net_1_r_15);
DFFARX1 I_43(n4_1_l_15,blif_clk_net_1_r_15,n4_15,G42_1_l_15,);
not I_44(n15_15,G42_1_l_15);
DFFARX1 I_45(G42_1_r_6,blif_clk_net_1_r_15,n4_15,n17_internal_15,);
not I_46(n17_15,n17_internal_15);
DFFARX1 I_47(n_572_1_r_6,blif_clk_net_1_r_15,n4_15,n30_15,);
nor I_48(n_572_1_l_15,n_549_1_r_6,P6_5_r_6);
DFFARX1 I_49(n_572_1_l_15,blif_clk_net_1_r_15,n4_15,n14_internal_15,);
not I_50(n14_15,n14_internal_15);
nand I_51(N1_4_r_15,n25_15,n26_15);
or I_52(n_573_1_l_15,G42_1_r_6,n_452_1_r_6);
nor I_53(n18_15,G42_1_r_6,n_573_1_r_6);
nand I_54(n19_15,n27_15,n28_15);
nand I_55(n20_15,n30_15,n_569_1_r_6);
not I_56(n21_15,n20_15);
and I_57(n22_15,n17_15,n_572_1_l_15);
nor I_58(n23_15,n_452_1_r_6,G199_4_r_6);
or I_59(n24_15,G42_1_r_6,n_573_1_r_6);
or I_60(n25_15,n_573_1_l_15,G199_4_r_6);
nand I_61(n26_15,n19_15,n23_15);
not I_62(n27_15,n_573_1_r_6);
nand I_63(n28_15,n29_15,ACVQN1_5_r_6);
not I_64(n29_15,n_549_1_r_6);
endmodule


