module test_I7570_rst(I1477_rst,I7570_rst);
,I7570_rst);
input I1477_rst;
output I7570_rst;
wire ;
not I_0(I7570_rst,I1477_rst);
endmodule


