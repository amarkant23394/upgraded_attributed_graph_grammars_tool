module test_final(IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_5_r_13,blif_reset_net_5_r_13,N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13);
input IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_5_r_13,blif_reset_net_5_r_13;
output N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13;
wire N1371_0_r_8,N1508_0_r_8,N1372_1_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N1508_10_r_8,N3_8_l_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8,n_102_5_r_13,n4_7_l_13,n9_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13;
nor I_0(N1371_0_r_8,n46_8,n51_8);
not I_1(N1508_0_r_8,n46_8);
nor I_2(N1372_1_r_8,n37_8,n49_8);
and I_3(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_4(N1507_6_r_8,n47_8,n48_8);
nor I_5(N1508_6_r_8,n37_8,n38_8);
nor I_6(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_7(N3_8_r_8,blif_clk_net_5_r_13,n9_13,G199_8_r_8,);
nor I_8(N6147_9_r_8,n29_8,n30_8);
nor I_9(N6134_9_r_8,n30_8,n31_8);
not I_10(I_BUFF_1_9_r_8,n35_8);
nor I_11(N1372_10_r_8,n46_8,n49_8);
nor I_12(N1508_10_r_8,n40_8,n41_8);
and I_13(N3_8_l_8,IN_6_8_l_8,n36_8);
DFFARX1 I_14(N3_8_l_8,blif_clk_net_5_r_13,n9_13,n53_8,);
not I_15(n29_8,n53_8);
nor I_16(N3_8_r_8,n33_8,n34_8);
and I_17(n30_8,n32_8,n33_8);
nor I_18(n31_8,IN_1_8_l_8,IN_3_8_l_8);
nand I_19(n32_8,IN_2_6_l_8,n42_8);
or I_20(n33_8,IN_3_1_l_8,n46_8);
nor I_21(n34_8,n32_8,n35_8);
nand I_22(n35_8,IN_5_6_l_8,n44_8);
nand I_23(n36_8,IN_2_8_l_8,IN_3_8_l_8);
not I_24(n37_8,n31_8);
nand I_25(n38_8,N1508_0_r_8,n39_8);
nand I_26(n39_8,n33_8,n50_8);
and I_27(n40_8,n32_8,n35_8);
not I_28(n41_8,N1372_10_r_8);
and I_29(n42_8,IN_1_6_l_8,n43_8);
nand I_30(n43_8,n44_8,n45_8);
nand I_31(n44_8,IN_3_6_l_8,IN_4_6_l_8);
not I_32(n45_8,IN_5_6_l_8);
nand I_33(n46_8,IN_1_1_l_8,IN_2_1_l_8);
not I_34(n47_8,n39_8);
nor I_35(n48_8,n35_8,n49_8);
not I_36(n49_8,n51_8);
nand I_37(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_38(n51_8,IN_1_3_l_8,n52_8);
or I_39(n52_8,IN_2_3_l_8,IN_3_3_l_8);
nor I_40(N1371_0_r_13,n59_13,n61_13);
nor I_41(N1508_0_r_13,n59_13,n60_13);
not I_42(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_43(n_431_5_r_13,blif_clk_net_5_r_13,n9_13,G78_5_r_13,);
nand I_44(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_45(n_102_5_r_13,N1508_6_r_8,G199_8_r_8);
nand I_46(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_47(n1_13,blif_clk_net_5_r_13,n9_13,G42_7_r_13,);
nor I_48(n_572_7_r_13,n40_13,n41_13);
nand I_49(n_573_7_r_13,n37_13,n38_13);
nor I_50(n_549_7_r_13,n46_13,n47_13);
nand I_51(n_569_7_r_13,n37_13,n43_13);
nand I_52(n_452_7_r_13,n52_13,n53_13);
nor I_53(n4_7_l_13,N6134_9_r_8,N1508_10_r_8);
not I_54(n9_13,blif_reset_net_5_r_13);
DFFARX1 I_55(n4_7_l_13,blif_clk_net_5_r_13,n9_13,n62_13,);
not I_56(n33_13,n62_13);
nand I_57(n_431_5_r_13,n54_13,n55_13);
not I_58(n1_13,n52_13);
nor I_59(n34_13,n35_13,n36_13);
nor I_60(n35_13,n42_13,N1371_0_r_8);
nand I_61(n36_13,n50_13,n58_13);
nand I_62(n37_13,n44_13,n45_13);
or I_63(n38_13,n39_13,N1371_0_r_8);
nand I_64(n39_13,n_42_8_r_8,N1508_1_r_8);
not I_65(n40_13,n36_13);
nor I_66(n41_13,n35_13,N1508_6_r_8);
not I_67(n42_13,n_42_8_r_8);
or I_68(n43_13,N6147_9_r_8,N1508_10_r_8);
not I_69(n44_13,N1371_0_r_8);
not I_70(n45_13,N1507_6_r_8);
nor I_71(n46_13,n39_13,n40_13);
nor I_72(n47_13,N6147_9_r_8,N1508_10_r_8);
nor I_73(n48_13,n50_13,n51_13);
nor I_74(n49_13,N1507_6_r_8,N1371_0_r_8);
not I_75(n50_13,n59_13);
not I_76(n51_13,n_102_5_r_13);
nand I_77(n52_13,n33_13,n39_13);
nand I_78(n53_13,n33_13,N1371_0_r_8);
nor I_79(n54_13,N6147_9_r_8,G199_8_r_8);
nand I_80(n55_13,n62_13,n56_13);
nor I_81(n56_13,n39_13,n57_13);
not I_82(n57_13,N1508_10_r_8);
or I_83(n58_13,N1508_1_r_8,G199_8_r_8);
nand I_84(n59_13,N1507_6_r_8,N1508_6_r_8);
nor I_85(n60_13,n51_13,N6147_9_r_8);
nor I_86(n61_13,n39_13,N1371_0_r_8);
endmodule


