module test_final(IN_1_1_l_4,IN_2_1_l_4,IN_3_1_l_4,IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_3_l_4,IN_2_3_l_4,IN_3_3_l_4,blif_clk_net_5_r_3,blif_reset_net_5_r_3,N1371_0_r_3,N1508_0_r_3,N6147_3_r_3,n_429_or_0_5_r_3,G78_5_r_3,n_576_5_r_3,n_102_5_r_3,n_547_5_r_3,N1508_10_r_3);
input IN_1_1_l_4,IN_2_1_l_4,IN_3_1_l_4,IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_3_l_4,IN_2_3_l_4,IN_3_3_l_4,blif_clk_net_5_r_3,blif_reset_net_5_r_3;
output N1371_0_r_3,N1508_0_r_3,N6147_3_r_3,n_429_or_0_5_r_3,G78_5_r_3,n_576_5_r_3,n_102_5_r_3,n_547_5_r_3,N1508_10_r_3;
wire N1371_0_r_4,N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_102_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4,n_431_5_r_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,N1372_10_r_3,N3_8_l_3,n5_3,n39_3,n_431_5_r_3,n22_3,n23_3,n24_3,n25_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3;
nor I_0(N1371_0_r_4,n25_4,n29_4);
nor I_1(N1508_0_r_4,n25_4,n32_4);
nor I_2(N6147_2_r_4,n24_4,n31_4);
or I_3(n_429_or_0_5_r_4,n23_4,n30_4);
DFFARX1 I_4(n_431_5_r_4,blif_clk_net_5_r_3,n5_3,G78_5_r_4,);
nand I_5(n_576_5_r_4,n22_4,n23_4);
nand I_6(n_102_5_r_4,n34_4,n35_4);
nand I_7(n_547_5_r_4,n26_4,n27_4);
nor I_8(N1507_6_r_4,n27_4,n30_4);
nor I_9(N1508_6_r_4,n30_4,n33_4);
nand I_10(n_431_5_r_4,n_102_5_r_4,n28_4);
nor I_11(n22_4,n24_4,n25_4);
nor I_12(n23_4,IN_1_3_l_4,n37_4);
not I_13(n24_4,n_102_5_r_4);
nand I_14(n25_4,IN_1_1_l_4,IN_2_1_l_4);
nor I_15(n26_4,n23_4,n24_4);
not I_16(n27_4,n25_4);
nand I_17(n28_4,n23_4,n29_4);
nor I_18(n29_4,IN_3_1_l_4,n25_4);
not I_19(n30_4,n29_4);
nor I_20(n31_4,N1371_0_r_4,n32_4);
nor I_21(n32_4,n23_4,n29_4);
nand I_22(n33_4,n23_4,n24_4);
nor I_23(n34_4,IN_1_2_l_4,IN_2_2_l_4);
or I_24(n35_4,IN_5_2_l_4,n36_4);
nor I_25(n36_4,IN_3_2_l_4,IN_4_2_l_4);
or I_26(n37_4,IN_2_3_l_4,IN_3_3_l_4);
nor I_27(N1371_0_r_3,n39_3,n37_3);
nor I_28(N1508_0_r_3,n25_3,n37_3);
nor I_29(N6147_3_r_3,N1372_10_r_3,n33_3);
nand I_30(n_429_or_0_5_r_3,N1372_10_r_3,n30_3);
DFFARX1 I_31(n_431_5_r_3,blif_clk_net_5_r_3,n5_3,G78_5_r_3,);
nand I_32(n_576_5_r_3,n22_3,n23_3);
not I_33(n_102_5_r_3,n39_3);
nand I_34(n_547_5_r_3,n26_3,n27_3);
not I_35(N1372_10_r_3,n36_3);
nor I_36(N1508_10_r_3,n35_3,n36_3);
and I_37(N3_8_l_3,n34_3,N1508_0_r_4);
not I_38(n5_3,blif_reset_net_5_r_3);
DFFARX1 I_39(N3_8_l_3,blif_clk_net_5_r_3,n5_3,n39_3,);
nand I_40(n_431_5_r_3,n29_3,n30_3);
nor I_41(n22_3,n24_3,n25_3);
nor I_42(n23_3,n39_3,N1508_6_r_4);
not I_43(n24_3,n27_3);
nand I_44(n25_3,n_429_or_0_5_r_4,G78_5_r_4);
nor I_45(n26_3,n39_3,n28_3);
nor I_46(n27_3,N6147_2_r_4,N1507_6_r_4);
not I_47(n28_3,n37_3);
nand I_48(n29_3,N1372_10_r_3,n39_3);
nand I_49(n30_3,n31_3,n32_3);
not I_50(n31_3,n25_3);
not I_51(n32_3,N1508_6_r_4);
nand I_52(n33_3,n24_3,n25_3);
nand I_53(n34_3,n_576_5_r_4,N1507_6_r_4);
nor I_54(n35_3,n27_3,n31_3);
nand I_55(n36_3,n28_3,n38_3);
nand I_56(n37_3,n_547_5_r_4,n_429_or_0_5_r_4);
or I_57(n38_3,N1508_0_r_4,N6147_2_r_4);
endmodule


