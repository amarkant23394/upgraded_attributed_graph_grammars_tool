module test_I9576(I1477,I5898,I5716,I6265,I8445,I8233,I1470,I9576);
input I1477,I5898,I5716,I6265,I8445,I8233,I1470;
output I9576;
wire I8527,I8202,I8496,I8216,I5719,I8377,I8250,I5737,I8181,I8360,I5751,I6203,I8592,I8462,I8267,I5713;
nand I_0(I8527,I8233,I5713);
nand I_1(I8202,I8267,I8496);
nor I_2(I8496,I8462,I8377);
not I_3(I8216,I1477);
DFFARX1 I_4(I6265,I1470,I5751,,,I5719,);
not I_5(I8377,I8360);
nor I_6(I8250,I5719,I5716);
nand I_7(I5737,I6203,I5898);
and I_8(I8181,I8360,I8592);
not I_9(I8360,I5719);
not I_10(I5751,I1477);
DFFARX1 I_11(I1470,I5751,,,I6203,);
DFFARX1 I_12(I8527,I1470,I8216,,,I8592,);
DFFARX1 I_13(I8445,I1470,I8216,,,I8462,);
nor I_14(I9576,I8181,I8202);
nand I_15(I8267,I8250,I5737);
DFFARX1 I_16(I1470,I5751,,,I5713,);
endmodule


