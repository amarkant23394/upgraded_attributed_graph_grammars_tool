module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_8_r_8,blif_reset_net_8_r_8,N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_8_r_8,blif_reset_net_8_r_8;
output N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,N1508_0_r_8,N1372_1_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N3_8_l_8,n8_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_8_r_8,n8_8,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_8_r_8,n8_8,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
nor I_35(N1371_0_r_8,n46_8,n51_8);
not I_36(N1508_0_r_8,n46_8);
nor I_37(N1372_1_r_8,n37_8,n49_8);
and I_38(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_39(N1507_6_r_8,n47_8,n48_8);
nor I_40(N1508_6_r_8,n37_8,n38_8);
nor I_41(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_42(N3_8_r_8,blif_clk_net_8_r_8,n8_8,G199_8_r_8,);
nor I_43(N6147_9_r_8,n29_8,n30_8);
nor I_44(N6134_9_r_8,n30_8,n31_8);
not I_45(I_BUFF_1_9_r_8,n35_8);
nor I_46(N1372_10_r_8,n46_8,n49_8);
nor I_47(N1508_10_r_8,n40_8,n41_8);
and I_48(N3_8_l_8,n36_8,n_547_5_r_0);
not I_49(n8_8,blif_reset_net_8_r_8);
DFFARX1 I_50(N3_8_l_8,blif_clk_net_8_r_8,n8_8,n53_8,);
not I_51(n29_8,n53_8);
nor I_52(N3_8_r_8,n33_8,n34_8);
and I_53(n30_8,n32_8,n33_8);
nor I_54(n31_8,N1371_0_r_0,N1508_0_r_0);
nand I_55(n32_8,n42_8,n_429_or_0_5_r_0);
or I_56(n33_8,n46_8,n_572_7_r_0);
nor I_57(n34_8,n32_8,n35_8);
nand I_58(n35_8,n44_8,n_576_5_r_0);
nand I_59(n36_8,N1371_0_r_0,N1508_0_r_0);
not I_60(n37_8,n31_8);
nand I_61(n38_8,N1508_0_r_8,n39_8);
nand I_62(n39_8,n33_8,n50_8);
and I_63(n40_8,n32_8,n35_8);
not I_64(n41_8,N1372_10_r_8);
and I_65(n42_8,n43_8,n_569_7_r_0);
nand I_66(n43_8,n44_8,n45_8);
nand I_67(n44_8,G42_7_r_0,N1371_0_r_0);
not I_68(n45_8,n_576_5_r_0);
nand I_69(n46_8,G78_5_r_0,n_549_7_r_0);
not I_70(n47_8,n39_8);
nor I_71(n48_8,n35_8,n49_8);
not I_72(n49_8,n51_8);
nand I_73(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_74(n51_8,n52_8,n_573_7_r_0);
or I_75(n52_8,n_429_or_0_5_r_0,G78_5_r_0);
endmodule


