module test_final(IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_102_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7,n_452_7_r_7,n4_7_l_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
nor I_0(N1371_0_r_7,n53_7,n52_7);
nor I_1(N1508_0_r_7,n51_7,n52_7);
nand I_2(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_3(n_431_5_r_7,blif_clk_net_7_r_1,n9_1,G78_5_r_7,);
nand I_4(n_576_5_r_7,n31_7,n32_7);
nor I_5(n_102_5_r_7,IN_5_7_l_7,IN_9_7_l_7);
nand I_6(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_7(n4_7_r_7,blif_clk_net_7_r_1,n9_1,G42_7_r_7,);
nor I_8(n_572_7_r_7,n54_7,n33_7);
nand I_9(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_10(n_549_7_r_7,n53_7,n36_7);
nand I_11(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_12(n_452_7_r_7,IN_1_1_l_7,IN_2_1_l_7);
nor I_13(n4_7_l_7,G18_7_l_7,IN_1_7_l_7);
DFFARX1 I_14(n4_7_l_7,blif_clk_net_7_r_1,n9_1,n53_7,);
not I_15(n30_7,n53_7);
and I_16(N3_8_l_7,IN_6_8_l_7,n50_7);
DFFARX1 I_17(N3_8_l_7,blif_clk_net_7_r_1,n9_1,n54_7,);
nand I_18(n_431_5_r_7,n40_7,n41_7);
nor I_19(n4_7_r_7,n54_7,n49_7);
and I_20(n31_7,n_102_5_r_7,n39_7);
not I_21(n32_7,G18_7_l_7);
nor I_22(n33_7,IN_10_7_l_7,n34_7);
and I_23(n34_7,IN_4_7_l_7,n35_7);
not I_24(n35_7,G15_7_l_7);
nor I_25(n36_7,G18_7_l_7,n37_7);
or I_26(n37_7,IN_5_7_l_7,n54_7);
or I_27(n38_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_28(n39_7,IN_3_1_l_7,n_452_7_r_7);
nand I_29(n40_7,n46_7,n47_7);
nand I_30(n41_7,n42_7,n43_7);
nor I_31(n42_7,n44_7,n45_7);
nor I_32(n43_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_33(n44_7,G15_7_l_7,IN_7_7_l_7);
nor I_34(n45_7,IN_9_7_l_7,IN_10_7_l_7);
nand I_35(n46_7,IN_4_7_l_7,n35_7);
not I_36(n47_7,IN_10_7_l_7);
or I_37(n48_7,IN_3_1_l_7,n_452_7_r_7);
not I_38(n49_7,n_452_7_r_7);
nand I_39(n50_7,IN_2_8_l_7,IN_3_8_l_7);
and I_40(n51_7,n_452_7_r_7,n45_7);
not I_41(n52_7,n44_7);
and I_42(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_43(N1508_0_r_1,n40_1,n44_1);
nor I_44(N1507_6_r_1,n43_1,n49_1);
nor I_45(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_46(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_47(n_572_7_r_1,n29_1,n30_1);
not I_48(n_573_7_r_1,n_452_7_r_1);
nor I_49(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_50(n_569_7_r_1,n30_1,n31_1);
nor I_51(n_452_7_r_1,n30_1,n32_1);
nor I_52(N6147_9_r_1,n35_1,n36_1);
nand I_53(N6134_9_r_1,n38_1,n39_1);
not I_54(I_BUFF_1_9_r_1,n40_1);
nor I_55(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_56(n9_1,blif_reset_net_7_r_1);
nor I_57(n29_1,n34_1,G78_5_r_7);
nor I_58(n30_1,n33_1,n34_1);
nor I_59(n31_1,n54_1,n_572_7_r_7);
not I_60(n32_1,n48_1);
nor I_61(n33_1,N1371_0_r_7,N1508_0_r_7);
not I_62(n34_1,n_547_5_r_7);
nor I_63(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_64(n36_1,n29_1);
not I_65(n37_1,n41_1);
nand I_66(n38_1,I_BUFF_1_9_r_1,n_576_5_r_7);
nand I_67(n39_1,n37_1,n40_1);
nand I_68(n40_1,n_429_or_0_5_r_7,n_569_7_r_7);
nand I_69(n41_1,n52_1,G78_5_r_7);
or I_70(n42_1,n36_1,n43_1);
nor I_71(n43_1,n32_1,n49_1);
nand I_72(n44_1,n45_1,n46_1);
nand I_73(n45_1,n47_1,n48_1);
not I_74(n46_1,n_576_5_r_7);
not I_75(n47_1,n31_1);
nand I_76(n48_1,n50_1,n_573_7_r_7);
nor I_77(n49_1,n41_1,n47_1);
and I_78(n50_1,n51_1,n_549_7_r_7);
nand I_79(n51_1,n52_1,n53_1);
nand I_80(n52_1,G42_7_r_7,n_429_or_0_5_r_7);
not I_81(n53_1,G78_5_r_7);
or I_82(n54_1,N1371_0_r_7,N1508_0_r_7);
nor I_83(n55_1,n29_1,n_576_5_r_7);
endmodule


