module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_7_r_12,blif_reset_net_7_r_12,N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_7_r_12,blif_reset_net_7_r_12;
output N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12;
wire N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1372_4_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10,n_573_7_r_12,n_452_7_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n8_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12;
nor I_0(N1371_0_r_10,n37_10,n38_10);
nor I_1(N1508_0_r_10,n37_10,n58_10);
nand I_2(N6147_2_r_10,n39_10,n40_10);
not I_3(N6147_3_r_10,n39_10);
nor I_4(N1372_4_r_10,n46_10,n49_10);
nor I_5(N1508_4_r_10,n51_10,n52_10);
nor I_6(N1507_6_r_10,n49_10,n60_10);
nor I_7(N1508_6_r_10,n49_10,n50_10);
nor I_8(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_9(N3_8_r_10,blif_clk_net_7_r_12,n8_12,G199_8_r_10,);
nor I_10(N6147_9_r_10,n36_10,n37_10);
nor I_11(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_12(I_BUFF_1_9_r_10,n48_10);
nor I_13(N3_8_r_10,n44_10,n47_10);
not I_14(n35_10,n49_10);
nor I_15(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_16(n37_10,IN_1_9_l_10);
not I_17(n38_10,n46_10);
nand I_18(n39_10,n43_10,n44_10);
nand I_19(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_20(n41_10,IN_1_9_l_10,n42_10);
not I_21(n42_10,n44_10);
nor I_22(n43_10,IN_1_9_l_10,n45_10);
nand I_23(n44_10,IN_2_6_l_10,n54_10);
nor I_24(n45_10,IN_5_9_l_10,n59_10);
nand I_25(n46_10,IN_2_9_l_10,n61_10);
nor I_26(n47_10,n46_10,n48_10);
nand I_27(n48_10,n62_10,n63_10);
nand I_28(n49_10,IN_5_6_l_10,n56_10);
not I_29(n50_10,n45_10);
nor I_30(n51_10,n42_10,n53_10);
not I_31(n52_10,N1372_4_r_10);
nor I_32(n53_10,n48_10,n50_10);
and I_33(n54_10,IN_1_6_l_10,n55_10);
nand I_34(n55_10,n56_10,n57_10);
nand I_35(n56_10,IN_3_6_l_10,IN_4_6_l_10);
not I_36(n57_10,IN_5_6_l_10);
nor I_37(n58_10,n35_10,n45_10);
nor I_38(n59_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_39(n60_10,n37_10,n46_10);
or I_40(n61_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_41(n62_10,IN_1_2_l_10,IN_2_2_l_10);
or I_42(n63_10,IN_5_2_l_10,n64_10);
nor I_43(n64_10,IN_3_2_l_10,IN_4_2_l_10);
nor I_44(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_45(N1508_0_r_12,n30_12,n37_12);
nor I_46(N1507_6_r_12,n25_12,n39_12);
nor I_47(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_48(n1_12,blif_clk_net_7_r_12,n8_12,G42_7_r_12,);
nor I_49(n_572_7_r_12,n23_12,n24_12);
nand I_50(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_51(n_549_7_r_12,n27_12,n28_12);
nand I_52(n_569_7_r_12,n25_12,n26_12);
nand I_53(n_452_7_r_12,G199_8_r_10,N1508_0_r_10);
nand I_54(N6147_9_r_12,n30_12,n31_12);
nor I_55(N6134_9_r_12,n35_12,n36_12);
not I_56(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_57(n1_12,n_573_7_r_12);
not I_58(n8_12,blif_reset_net_7_r_12);
not I_59(n23_12,n36_12);
nor I_60(n24_12,n_452_7_r_12,N1371_0_r_10);
nand I_61(n25_12,n23_12,n40_12);
not I_62(n26_12,n35_12);
not I_63(n27_12,N6134_9_r_12);
nand I_64(n28_12,n26_12,n29_12);
not I_65(n29_12,n24_12);
nand I_66(n30_12,n33_12,n41_12);
nand I_67(n31_12,n32_12,n33_12);
nor I_68(n32_12,n26_12,n34_12);
nor I_69(n33_12,n_42_8_r_10,N1371_0_r_10);
nor I_70(n34_12,n42_12,N6134_9_r_10);
nor I_71(n35_12,n38_12,N1508_4_r_10);
nand I_72(n36_12,N1508_0_r_10,N1508_6_r_10);
nand I_73(n37_12,n23_12,n35_12);
or I_74(n38_12,N1507_6_r_10,N6147_2_r_10);
not I_75(n39_12,n30_12);
or I_76(n40_12,N6147_2_r_10,N6147_9_r_10);
nor I_77(n41_12,n34_12,n36_12);
nor I_78(n42_12,N6147_3_r_10,N1508_4_r_10);
endmodule


