module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_7_r_16,blif_reset_net_7_r_16,N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16);
input IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_7_r_16,blif_reset_net_7_r_16;
output N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16;
wire N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_102_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1372_10_r_11,N1508_10_r_11,n_431_5_r_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11,n_549_7_r_16,N3_8_l_16,n8_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16;
not I_0(N1372_1_r_11,n53_11);
nor I_1(N1508_1_r_11,n39_11,n53_11);
nor I_2(N6147_2_r_11,n48_11,n49_11);
nor I_3(N6147_3_r_11,n44_11,n45_11);
nand I_4(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_5(n_431_5_r_11,blif_clk_net_7_r_16,n8_16,G78_5_r_11,);
nand I_6(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_7(n_102_5_r_11,n39_11);
nand I_8(n_547_5_r_11,n36_11,n37_11);
nor I_9(N1507_6_r_11,n52_11,n57_11);
nor I_10(N1508_6_r_11,n46_11,n51_11);
nor I_11(N1372_10_r_11,n43_11,n47_11);
nor I_12(N1508_10_r_11,n55_11,n56_11);
nand I_13(n_431_5_r_11,n40_11,n41_11);
nor I_14(n36_11,n38_11,n39_11);
not I_15(n37_11,n40_11);
nor I_16(n38_11,IN_2_0_l_11,n60_11);
nor I_17(n39_11,IN_1_3_l_11,n54_11);
nand I_18(n40_11,IN_1_1_l_11,IN_2_1_l_11);
nand I_19(n41_11,n_102_5_r_11,n42_11);
and I_20(n42_11,IN_2_6_l_11,n58_11);
not I_21(n43_11,n44_11);
nor I_22(n44_11,IN_3_1_l_11,n40_11);
nand I_23(n45_11,n46_11,n47_11);
not I_24(n46_11,n38_11);
nand I_25(n47_11,n59_11,n62_11);
and I_26(n48_11,n37_11,n47_11);
or I_27(n49_11,n44_11,n50_11);
nor I_28(n50_11,n60_11,n61_11);
or I_29(n51_11,n_102_5_r_11,n52_11);
nor I_30(n52_11,n42_11,n57_11);
nand I_31(n53_11,n37_11,n50_11);
or I_32(n54_11,IN_2_3_l_11,IN_3_3_l_11);
nor I_33(n55_11,n38_11,n42_11);
not I_34(n56_11,N1372_10_r_11);
and I_35(n57_11,n38_11,n50_11);
and I_36(n58_11,IN_1_6_l_11,n59_11);
or I_37(n59_11,IN_5_6_l_11,n63_11);
not I_38(n60_11,IN_1_0_l_11);
nor I_39(n61_11,IN_3_0_l_11,IN_4_0_l_11);
nand I_40(n62_11,IN_3_6_l_11,IN_4_6_l_11);
and I_41(n63_11,IN_3_6_l_11,IN_4_6_l_11);
nor I_42(N1371_0_r_16,n35_16,n39_16);
nor I_43(N1508_0_r_16,n39_16,n46_16);
not I_44(N1372_1_r_16,n45_16);
nor I_45(N1508_1_r_16,n53_16,n45_16);
nor I_46(N6147_2_r_16,n37_16,n38_16);
nor I_47(N1507_6_r_16,n44_16,n49_16);
nor I_48(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_49(n4_7_r_16,blif_clk_net_7_r_16,n8_16,G42_7_r_16,);
nor I_50(n_572_7_r_16,n32_16,n33_16);
nand I_51(n_573_7_r_16,n30_16,n31_16);
nand I_52(n_549_7_r_16,n47_16,N6147_2_r_11);
nand I_53(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_54(n_452_7_r_16,n34_16,n35_16);
and I_55(N3_8_l_16,n41_16,N1507_6_r_11);
not I_56(n8_16,blif_reset_net_7_r_16);
DFFARX1 I_57(N3_8_l_16,blif_clk_net_7_r_16,n8_16,n53_16,);
not I_58(n29_16,n53_16);
nor I_59(n4_7_r_16,n35_16,n36_16);
nand I_60(n30_16,n_429_or_0_5_r_11,n_547_5_r_11);
not I_61(n31_16,n34_16);
nor I_62(n32_16,n30_16,N6147_3_r_11);
not I_63(n33_16,n_549_7_r_16);
nor I_64(n34_16,n48_16,N1508_1_r_11);
and I_65(n35_16,n50_16,n_576_5_r_11);
not I_66(n36_16,n30_16);
nor I_67(n37_16,n31_16,n40_16);
nand I_68(n38_16,n29_16,n39_16);
not I_69(n39_16,n32_16);
nor I_70(n40_16,N6147_2_r_11,N1508_6_r_11);
nand I_71(n41_16,G78_5_r_11,N1508_6_r_11);
nand I_72(n42_16,n35_16,n43_16);
not I_73(n43_16,n44_16);
nor I_74(n44_16,n32_16,n49_16);
nand I_75(n45_16,n36_16,n40_16);
nor I_76(n46_16,n33_16,n34_16);
nand I_77(n47_16,N1508_1_r_11,N1372_1_r_11);
or I_78(n48_16,N1372_1_r_11,N1508_10_r_11);
and I_79(n49_16,n35_16,n36_16);
and I_80(n50_16,n51_16,N6147_3_r_11);
nand I_81(n51_16,n47_16,n52_16);
not I_82(n52_16,N6147_2_r_11);
endmodule


