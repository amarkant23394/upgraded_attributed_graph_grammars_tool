module test_I9816(I1477,I5743,I1470,I9816);
input I1477,I5743,I1470;
output I9816;
wire I8216,I8623,I8705,I8193,I9491;
not I_0(I8216,I1477);
DFFARX1 I_1(I5743,I1470,I8216,,,I8623,);
DFFARX1 I_2(I8623,I1470,I8216,,,I8705,);
DFFARX1 I_3(I8193,I1470,I9491,,,I9816,);
not I_4(I8193,I8705);
not I_5(I9491,I1477);
endmodule


