module test_I5187(I1477,I3538,I3487,I1489,I1504,I1498,I1470,I2103,I5187);
input I1477,I3538,I3487,I1489,I1504,I1498,I1470,I2103;
output I5187;
wire I3521,I3504,I1495,I3747,I3685,I3388,I3668,I3846,I5122,I1518,I3380,I3350,I3555;
nor I_0(I3521,I3504,I1495);
and I_1(I3504,I3487,I1489);
DFFARX1 I_2(I2103,I1470,I1518,,,I1495,);
DFFARX1 I_3(I1504,I1470,I3388,,,I3747,);
and I_4(I3685,I3668,I1498);
not I_5(I3388,I1477);
DFFARX1 I_6(I1470,I3388,,,I3668,);
nor I_7(I3846,I3747,I3555);
not I_8(I5122,I3350);
not I_9(I1518,I1477);
nor I_10(I5187,I5122,I3380);
nand I_11(I3380,I3521,I3846);
DFFARX1 I_12(I3685,I1470,I3388,,,I3350,);
DFFARX1 I_13(I3538,I1470,I3388,,,I3555,);
endmodule


