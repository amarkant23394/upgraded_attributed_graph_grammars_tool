module test_I8862_rst(I1477_rst,I8862_rst);
,I8862_rst);
input I1477_rst;
output I8862_rst;
wire ;
not I_0(I8862_rst,I1477_rst);
endmodule


