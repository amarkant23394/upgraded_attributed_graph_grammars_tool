module test_I5351(I3374,I1477,I1470,I5283,I5351);
input I3374,I1477,I1470,I5283;
output I5351;
wire I3388,I3422,I3702,I3362,I1480,I1483,I5334,I3365,I5317,I5105,I5300;
not I_0(I3388,I1477);
or I_1(I3422,I1483,I1480);
DFFARX1 I_2(I1470,I3388,,,I3702,);
DFFARX1 I_3(I5334,I1470,I5105,,,I5351,);
DFFARX1 I_4(I3422,I1470,I3388,,,I3362,);
DFFARX1 I_5(I1470,,,I1480,);
DFFARX1 I_6(I1470,,,I1483,);
or I_7(I5334,I5317,I3362);
not I_8(I3365,I3702);
and I_9(I5317,I5300,I3365);
not I_10(I5105,I1477);
nor I_11(I5300,I5283,I3374);
endmodule


