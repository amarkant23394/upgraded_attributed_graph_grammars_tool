module test_I5563(I1504,I1477,I5122,I3380,I1470,I3453,I5563);
input I1504,I1477,I5122,I3380,I1470,I3453;
output I5563;
wire I3388,I3368,I3470,I5187,I5546,I5204,I3353,I3637,I5529,I5512,I3747,I5105;
not I_0(I3388,I1477);
nand I_1(I3368,I3747,I3470);
not I_2(I3470,I3453);
nor I_3(I5187,I5122,I3380);
nor I_4(I5546,I5204,I5529);
nand I_5(I5204,I5187,I3353);
and I_6(I3353,I3453,I3637);
DFFARX1 I_7(I1470,I3388,,,I3637,);
and I_8(I5563,I5512,I5546);
not I_9(I5529,I5512);
DFFARX1 I_10(I3368,I1470,I5105,,,I5512,);
DFFARX1 I_11(I1504,I1470,I3388,,,I3747,);
not I_12(I5105,I1477);
endmodule


