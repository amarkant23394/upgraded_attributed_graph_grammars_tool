module test_I3560(I2733,I2583,I1902,I1294,I3560);
input I2733,I2583,I1902,I1294;
output I3560;
wire I3263,I3168,I3280,I2945,I2563,I2548,I2962,I3297,I2832,I2560,I2993,I3543,I2569,I2566,I3086,I3103;
not I_0(I3263,I2569);
nand I_1(I3560,I3543,I3297);
or I_2(I3168,I3103);
nor I_3(I3280,I2548,I2560);
DFFARX1 I_4(I1902,I1294,I2583,,,I2945,);
nand I_5(I2563,I3103,I2993);
DFFARX1 I_6(I2945,I1294,I2583,,,I2548,);
nor I_7(I2962,I2945);
nand I_8(I3297,I3280,I2563);
DFFARX1 I_9(I1294,I2583,,,I2832,);
DFFARX1 I_10(I3168,I1294,I2583,,,I2560,);
nor I_11(I2993,I2945,I2733);
nand I_12(I3543,I3263,I2566);
nand I_13(I2569,I2832,I2962);
not I_14(I2566,I2945);
DFFARX1 I_15(I1294,I2583,,,I3086,);
not I_16(I3103,I3086);
endmodule


