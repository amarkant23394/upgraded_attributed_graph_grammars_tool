module test_final(IN_1_2_l_1,IN_2_2_l_1,IN_3_2_l_1,IN_6_2_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_1_4_l_1,IN_2_4_l_1,IN_3_4_l_1,IN_6_4_l_1,blif_clk_net_1_r_3,blif_reset_net_1_r_3,G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3);
input IN_1_2_l_1,IN_2_2_l_1,IN_3_2_l_1,IN_6_2_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_1_4_l_1,IN_2_4_l_1,IN_3_4_l_1,IN_6_4_l_1,blif_clk_net_1_r_3,blif_reset_net_1_r_3;
output G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3;
wire G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1,N3_2_l_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1,n4_1_l_3,n9_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3;
DFFARX1 I_0(n4_1_r_1,blif_clk_net_1_r_3,n9_3,G42_1_r_1,);
nor I_1(n_572_1_r_1,n26_1,n19_1);
nand I_2(n_573_1_r_1,n16_1,n18_1);
nor I_3(n_549_1_r_1,n20_1,n21_1);
nor I_4(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_5(G199_4_l_1,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_1,);
nor I_6(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_7(N1_4_r_1,blif_clk_net_1_r_3,n9_3,G199_4_r_1,);
DFFARX1 I_8(G199_4_l_1,blif_clk_net_1_r_3,n9_3,G214_4_r_1,);
and I_9(N3_2_l_1,IN_6_2_l_1,n23_1);
DFFARX1 I_10(N3_2_l_1,blif_clk_net_1_r_3,n9_3,n26_1,);
not I_11(n17_1,n26_1);
DFFARX1 I_12(IN_1_3_l_1,blif_clk_net_1_r_3,n9_3,n16_internal_1,);
not I_13(n16_1,n16_internal_1);
DFFARX1 I_14(IN_2_3_l_1,blif_clk_net_1_r_3,n9_3,ACVQN1_3_l_1,);
and I_15(N1_4_l_1,IN_6_4_l_1,n25_1);
DFFARX1 I_16(N1_4_l_1,blif_clk_net_1_r_3,n9_3,G199_4_l_1,);
DFFARX1 I_17(IN_3_4_l_1,blif_clk_net_1_r_3,n9_3,G214_4_l_1,);
nor I_18(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_19(G214_4_l_1,blif_clk_net_1_r_3,n9_3,n14_internal_1,);
not I_20(n14_1,n14_internal_1);
nor I_21(N1_4_r_1,n17_1,n24_1);
nand I_22(n18_1,IN_4_3_l_1,ACVQN1_3_l_1);
nor I_23(n19_1,IN_1_2_l_1,IN_3_2_l_1);
not I_24(n20_1,n18_1);
nor I_25(n21_1,n26_1,n22_1);
not I_26(n22_1,n19_1);
nand I_27(n23_1,IN_2_2_l_1,IN_3_2_l_1);
nor I_28(n24_1,n18_1,n22_1);
nand I_29(n25_1,IN_1_4_l_1,IN_2_4_l_1);
DFFARX1 I_30(n4_1_r_3,blif_clk_net_1_r_3,n9_3,G42_1_r_3,);
nor I_31(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_32(n_573_1_r_3,n26_3,n27_3);
nor I_33(n_549_1_r_3,n40_3,n32_3);
nand I_34(n_569_1_r_3,n27_3,n31_3);
and I_35(n_452_1_r_3,n26_3,n_549_1_r_1);
nor I_36(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_37(N3_2_r_3,blif_clk_net_1_r_3,n9_3,G199_2_r_3,);
DFFARX1 I_38(n_572_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_3,);
nor I_39(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_40(n4_1_l_3,n_549_1_r_1,n_572_1_r_1);
not I_41(n9_3,blif_reset_net_1_r_3);
DFFARX1 I_42(n4_1_l_3,blif_clk_net_1_r_3,n9_3,G42_1_l_3,);
not I_43(n22_3,G42_1_l_3);
DFFARX1 I_44(G42_1_r_1,blif_clk_net_1_r_3,n9_3,n40_3,);
DFFARX1 I_45(G42_1_r_1,blif_clk_net_1_r_3,n9_3,n25_internal_3,);
not I_46(n25_3,n25_internal_3);
nor I_47(n4_1_r_3,n40_3,n36_3);
nor I_48(N3_2_r_3,n26_3,n37_3);
nor I_49(n_572_1_l_3,n_572_1_r_1,G199_4_r_1);
DFFARX1 I_50(G42_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN1_3_r_3,);
nor I_51(n26_3,n_266_and_0_3_r_1,G214_4_r_1);
not I_52(n27_3,n_452_1_r_1);
nor I_53(n28_3,n29_3,n_452_1_r_1);
nor I_54(n29_3,n30_3,n_572_1_r_1);
not I_55(n30_3,n_573_1_r_1);
nor I_56(n31_3,n40_3,G214_4_r_1);
nor I_57(n32_3,n25_3,n33_3);
nand I_58(n33_3,n22_3,ACVQN2_3_r_1);
or I_59(n34_3,n_452_1_r_1,G214_4_r_1);
nand I_60(n35_3,ACVQN1_3_r_3,ACVQN2_3_r_1);
nor I_61(n36_3,n_549_1_r_1,n_266_and_0_3_r_1);
nor I_62(n37_3,n38_3,n39_3);
not I_63(n38_3,n_572_1_l_3);
nand I_64(n39_3,n27_3,n30_3);
endmodule


