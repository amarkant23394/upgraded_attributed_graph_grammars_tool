module test_final(IN_1_2_l_1,IN_2_2_l_1,IN_3_2_l_1,IN_6_2_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_1_4_l_1,IN_2_4_l_1,IN_3_4_l_1,IN_6_4_l_1,blif_clk_net_1_r_14,blif_reset_net_1_r_14,G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14);
input IN_1_2_l_1,IN_2_2_l_1,IN_3_2_l_1,IN_6_2_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_1_4_l_1,IN_2_4_l_1,IN_3_4_l_1,IN_6_4_l_1,blif_clk_net_1_r_14,blif_reset_net_1_r_14;
output G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14;
wire G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1,N3_2_l_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1,n_452_1_r_14,n4_1_l_14,n3_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14;
DFFARX1 I_0(n4_1_r_1,blif_clk_net_1_r_14,n3_14,G42_1_r_1,);
nor I_1(n_572_1_r_1,n26_1,n19_1);
nand I_2(n_573_1_r_1,n16_1,n18_1);
nor I_3(n_549_1_r_1,n20_1,n21_1);
nor I_4(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_5(G199_4_l_1,blif_clk_net_1_r_14,n3_14,ACVQN2_3_r_1,);
nor I_6(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_7(N1_4_r_1,blif_clk_net_1_r_14,n3_14,G199_4_r_1,);
DFFARX1 I_8(G199_4_l_1,blif_clk_net_1_r_14,n3_14,G214_4_r_1,);
and I_9(N3_2_l_1,IN_6_2_l_1,n23_1);
DFFARX1 I_10(N3_2_l_1,blif_clk_net_1_r_14,n3_14,n26_1,);
not I_11(n17_1,n26_1);
DFFARX1 I_12(IN_1_3_l_1,blif_clk_net_1_r_14,n3_14,n16_internal_1,);
not I_13(n16_1,n16_internal_1);
DFFARX1 I_14(IN_2_3_l_1,blif_clk_net_1_r_14,n3_14,ACVQN1_3_l_1,);
and I_15(N1_4_l_1,IN_6_4_l_1,n25_1);
DFFARX1 I_16(N1_4_l_1,blif_clk_net_1_r_14,n3_14,G199_4_l_1,);
DFFARX1 I_17(IN_3_4_l_1,blif_clk_net_1_r_14,n3_14,G214_4_l_1,);
nor I_18(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_19(G214_4_l_1,blif_clk_net_1_r_14,n3_14,n14_internal_1,);
not I_20(n14_1,n14_internal_1);
nor I_21(N1_4_r_1,n17_1,n24_1);
nand I_22(n18_1,IN_4_3_l_1,ACVQN1_3_l_1);
nor I_23(n19_1,IN_1_2_l_1,IN_3_2_l_1);
not I_24(n20_1,n18_1);
nor I_25(n21_1,n26_1,n22_1);
not I_26(n22_1,n19_1);
nand I_27(n23_1,IN_2_2_l_1,IN_3_2_l_1);
nor I_28(n24_1,n18_1,n22_1);
nand I_29(n25_1,IN_1_4_l_1,IN_2_4_l_1);
DFFARX1 I_30(n_452_1_r_14,blif_clk_net_1_r_14,n3_14,G42_1_r_14,);
and I_31(n_572_1_r_14,n18_14,n19_14);
nand I_32(n_573_1_r_14,n16_14,n17_14);
nor I_33(n_549_1_r_14,n20_14,n21_14);
or I_34(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_35(n_452_1_r_14,n23_14,n_549_1_r_1);
nor I_36(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_37(N3_2_r_14,blif_clk_net_1_r_14,n3_14,G199_2_r_14,);
DFFARX1 I_38(n_572_1_l_14,blif_clk_net_1_r_14,n3_14,ACVQN1_5_r_14,);
not I_39(P6_5_r_14,P6_5_r_internal_14);
nor I_40(n4_1_l_14,G42_1_r_1,n_572_1_r_1);
not I_41(n3_14,blif_reset_net_1_r_14);
DFFARX1 I_42(n4_1_l_14,blif_clk_net_1_r_14,n3_14,n15_internal_14,);
not I_43(n15_14,n15_internal_14);
DFFARX1 I_44(n_573_1_r_1,blif_clk_net_1_r_14,n3_14,ACVQN2_3_l_14,);
DFFARX1 I_45(n_573_1_r_1,blif_clk_net_1_r_14,n3_14,ACVQN1_3_l_14,);
and I_46(N3_2_r_14,n26_14,n27_14);
nor I_47(n_572_1_l_14,ACVQN2_3_r_1,G199_4_r_1);
DFFARX1 I_48(ACVQN2_3_l_14,blif_clk_net_1_r_14,n3_14,P6_5_r_internal_14,);
nor I_49(n16_14,n_549_1_r_1,G214_4_r_1);
not I_50(n17_14,n_572_1_l_14);
nor I_51(n18_14,n_266_and_0_3_r_1,G214_4_r_1);
nand I_52(n19_14,ACVQN1_3_l_14,n_572_1_r_1);
nor I_53(n20_14,n_266_and_0_3_r_1,n_572_1_r_1);
nor I_54(n21_14,n15_14,n22_14);
nand I_55(n22_14,n24_14,n25_14);
nand I_56(n23_14,n15_14,n24_14);
not I_57(n24_14,G214_4_r_1);
not I_58(n25_14,n_266_and_0_3_r_1);
nor I_59(n26_14,n20_14,n_549_1_r_1);
nand I_60(n27_14,n28_14,n_452_1_r_1);
not I_61(n28_14,ACVQN2_3_r_1);
endmodule


