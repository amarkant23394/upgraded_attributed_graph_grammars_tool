module test_final(IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_7_r_14,blif_reset_net_7_r_14,N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14);
input IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_7_r_14,blif_reset_net_7_r_14;
output N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14;
wire N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_573_7_r_12,n_549_7_r_12,n_569_7_r_12,n_452_7_r_12,N6147_9_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12,I_BUFF_1_9_r_14,N3_8_l_14,n8_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14;
nor I_0(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_1(N1508_0_r_12,n30_12,n37_12);
nor I_2(N1507_6_r_12,n25_12,n39_12);
nor I_3(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_4(n1_12,blif_clk_net_7_r_14,n8_14,G42_7_r_12,);
nor I_5(n_572_7_r_12,n23_12,n24_12);
nand I_6(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_7(n_549_7_r_12,n27_12,n28_12);
nand I_8(n_569_7_r_12,n25_12,n26_12);
nand I_9(n_452_7_r_12,IN_1_1_l_12,IN_2_1_l_12);
nand I_10(N6147_9_r_12,n30_12,n31_12);
nor I_11(N6134_9_r_12,n35_12,n36_12);
not I_12(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_13(n1_12,n_573_7_r_12);
not I_14(n23_12,n36_12);
nor I_15(n24_12,IN_3_1_l_12,n_452_7_r_12);
nand I_16(n25_12,n23_12,n40_12);
not I_17(n26_12,n35_12);
not I_18(n27_12,N6134_9_r_12);
nand I_19(n28_12,n26_12,n29_12);
not I_20(n29_12,n24_12);
nand I_21(n30_12,n33_12,n41_12);
nand I_22(n31_12,n32_12,n33_12);
nor I_23(n32_12,n26_12,n34_12);
nor I_24(n33_12,IN_1_2_l_12,IN_2_2_l_12);
nor I_25(n34_12,IN_5_2_l_12,n42_12);
nor I_26(n35_12,IN_1_3_l_12,n38_12);
nand I_27(n36_12,IN_1_10_l_12,IN_2_10_l_12);
nand I_28(n37_12,n23_12,n35_12);
or I_29(n38_12,IN_2_3_l_12,IN_3_3_l_12);
not I_30(n39_12,n30_12);
or I_31(n40_12,IN_3_10_l_12,IN_4_10_l_12);
nor I_32(n41_12,n34_12,n36_12);
nor I_33(n42_12,IN_3_2_l_12,IN_4_2_l_12);
nor I_34(N1371_0_r_14,n47_14,n30_14);
nor I_35(N1508_0_r_14,n30_14,n41_14);
nor I_36(N1507_6_r_14,n37_14,n44_14);
nor I_37(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_38(n4_7_r_14,blif_clk_net_7_r_14,n8_14,G42_7_r_14,);
nor I_39(n_572_7_r_14,n28_14,n29_14);
nand I_40(n_573_7_r_14,n26_14,n27_14);
nor I_41(n_549_7_r_14,n31_14,n32_14);
nand I_42(n_569_7_r_14,n26_14,n30_14);
nor I_43(n_452_7_r_14,n47_14,n28_14);
nor I_44(N6147_9_r_14,n36_14,n37_14);
nor I_45(N6134_9_r_14,n28_14,n36_14);
not I_46(I_BUFF_1_9_r_14,n26_14);
and I_47(N3_8_l_14,n38_14,n_549_7_r_12);
not I_48(n8_14,blif_reset_net_7_r_14);
DFFARX1 I_49(N3_8_l_14,blif_clk_net_7_r_14,n8_14,n47_14,);
nor I_50(n4_7_r_14,n47_14,n35_14);
nand I_51(n26_14,n_569_7_r_12,G42_7_r_12);
not I_52(n27_14,n28_14);
nor I_53(n28_14,n43_14,n_572_7_r_12);
not I_54(n29_14,n33_14);
not I_55(n30_14,n31_14);
nor I_56(n31_14,n46_14,N1371_0_r_12);
and I_57(n32_14,n33_14,n34_14);
nand I_58(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_59(n34_14,n42_14,n43_14);
nor I_60(n35_14,G42_7_r_12,N1371_0_r_12);
nor I_61(n36_14,n47_14,n34_14);
not I_62(n37_14,n35_14);
nand I_63(n38_14,N1508_6_r_12,G42_7_r_12);
nand I_64(n39_14,n29_14,n40_14);
nand I_65(n40_14,n27_14,n37_14);
nor I_66(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_67(n42_14,n_572_7_r_12,N1508_6_r_12);
not I_68(n43_14,N6147_9_r_12);
nor I_69(n44_14,n27_14,n33_14);
or I_70(n45_14,N1508_0_r_12,N1507_6_r_12);
or I_71(n46_14,N1507_6_r_12,n_549_7_r_12);
endmodule


