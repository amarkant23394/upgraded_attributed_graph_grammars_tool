module test_I14650(I13214,I11290,I1477,I1470,I14650);
input I13214,I11290,I1477,I1470;
output I14650;
wire I13231,I13197,I13165,I13248,I14370;
and I_0(I13231,I13214,I11290);
not I_1(I13197,I1477);
DFFARX1 I_2(I13248,I1470,I13197,,,I13165,);
DFFARX1 I_3(I13165,I1470,I14370,,,I14650,);
DFFARX1 I_4(I13231,I1470,I13197,,,I13248,);
not I_5(I14370,I1477);
endmodule


