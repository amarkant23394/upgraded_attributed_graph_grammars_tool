module test_I6312(I6510,I3975,I1477,I1470,I4263,I4068,I6312);
input I6510,I3975,I1477,I1470,I4263,I4068;
output I6312;
wire I6606,I3954,I6722,I6640,I6442,I6329,I6688,I3948,I6623,I6705,I3972;
DFFARX1 I_0(I1470,I6329,,,I6606,);
not I_1(I3954,I4068);
or I_2(I6722,I6705,I6640);
and I_3(I6640,I6442,I6623);
nor I_4(I6442,I3975,I3954);
not I_5(I6329,I1477);
DFFARX1 I_6(I3948,I1470,I6329,,,I6688,);
DFFARX1 I_7(I1470,,,I3948,);
nor I_8(I6623,I6606,I6510);
DFFARX1 I_9(I6722,I1470,I6329,,,I6312,);
and I_10(I6705,I6688,I3972);
or I_11(I3972,I4263,I4068);
endmodule


