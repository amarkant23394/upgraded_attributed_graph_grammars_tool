module test_I4917(I1477,I1470,I1239,I4917);
input I1477,I1470,I1239;
output I4917;
wire I2181,I4544,I4869,I2149,I4674,I2155,I2678,I2345,I2633,I2695;
nor I_0(I4917,I4869,I4674);
not I_1(I2181,I1477);
not I_2(I4544,I1477);
DFFARX1 I_3(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_4(I2695,I1470,I2181,,,I2149,);
DFFARX1 I_5(I2155,I1470,I4544,,,I4674,);
DFFARX1 I_6(I2633,I1470,I2181,,,I2155,);
nand I_7(I2678,I2633);
DFFARX1 I_8(I1470,I2181,,,I2345,);
DFFARX1 I_9(I1239,I1470,I2181,,,I2633,);
and I_10(I2695,I2345,I2678);
endmodule


