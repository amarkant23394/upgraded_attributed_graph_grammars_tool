module test_I15194(I10633,I1477,I10766,I10732,I12599,I12653,I1470,I13057,I15194);
input I10633,I1477,I10766,I10732,I12599,I12653,I1470,I13057;
output I15194;
wire I12670,I11105,I10647,I12930,I12848,I12611,I13023,I12608,I10636,I12593,I12619,I12913,I15177,I15143,I12882,I15160,I10609;
DFFARX1 I_0(I12653,I1470,I12619,,,I12670,);
and I_1(I11105,I10766);
not I_2(I10647,I1477);
and I_3(I12930,I12913,I10609);
DFFARX1 I_4(I1470,I12619,,,I12848,);
DFFARX1 I_5(I13057,I1470,I12619,,,I12611,);
DFFARX1 I_6(I10636,I1470,I12619,,,I13023,);
nor I_7(I12608,I13023,I12930);
or I_8(I15194,I15177,I12608);
nor I_9(I10636,I10732,I10766);
nand I_10(I12593,I12670,I12882);
not I_11(I12619,I1477);
DFFARX1 I_12(I10633,I1470,I12619,,,I12913,);
and I_13(I15177,I15160,I12593);
not I_14(I15143,I12599);
not I_15(I12882,I12848);
nor I_16(I15160,I15143,I12611);
DFFARX1 I_17(I11105,I1470,I10647,,,I10609,);
endmodule


