module test_I11950(I10032,I1477,I10041,I1470,I12442,I12123,I11950);
input I10032,I1477,I10041,I1470,I12442,I12123;
output I11950;
wire I12270,I10219,I12476,I10014,I12349,I12493,I11990,I11973,I10052,I12459;
nand I_0(I12270,I11990,I10014);
DFFARX1 I_1(I12493,I1470,I11973,,,I11950,);
DFFARX1 I_2(I1470,I10052,,,I10219,);
and I_3(I12476,I12349,I12459);
DFFARX1 I_4(I10219,I1470,I10052,,,I10014,);
DFFARX1 I_5(I10041,I1470,I11973,,,I12349,);
or I_6(I12493,I12270,I12476);
not I_7(I11990,I10032);
not I_8(I11973,I1477);
not I_9(I10052,I1477);
nor I_10(I12459,I12442,I12123);
endmodule


