module test_I6329_rst(I1477_rst,I6329_rst);
,I6329_rst);
input I1477_rst;
output I6329_rst;
wire ;
not I_0(I6329_rst,I1477_rst);
endmodule


