module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_7_r_2,blif_reset_net_7_r_2,N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2);
input IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_7_r_2,blif_reset_net_7_r_2;
output N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2;
wire N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_102_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1372_10_r_11,N1508_10_r_11,n_431_5_r_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11,n4_7_l_2,n10_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2;
not I_0(N1372_1_r_11,n53_11);
nor I_1(N1508_1_r_11,n39_11,n53_11);
nor I_2(N6147_2_r_11,n48_11,n49_11);
nor I_3(N6147_3_r_11,n44_11,n45_11);
nand I_4(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_5(n_431_5_r_11,blif_clk_net_7_r_2,n10_2,G78_5_r_11,);
nand I_6(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_7(n_102_5_r_11,n39_11);
nand I_8(n_547_5_r_11,n36_11,n37_11);
nor I_9(N1507_6_r_11,n52_11,n57_11);
nor I_10(N1508_6_r_11,n46_11,n51_11);
nor I_11(N1372_10_r_11,n43_11,n47_11);
nor I_12(N1508_10_r_11,n55_11,n56_11);
nand I_13(n_431_5_r_11,n40_11,n41_11);
nor I_14(n36_11,n38_11,n39_11);
not I_15(n37_11,n40_11);
nor I_16(n38_11,IN_2_0_l_11,n60_11);
nor I_17(n39_11,IN_1_3_l_11,n54_11);
nand I_18(n40_11,IN_1_1_l_11,IN_2_1_l_11);
nand I_19(n41_11,n_102_5_r_11,n42_11);
and I_20(n42_11,IN_2_6_l_11,n58_11);
not I_21(n43_11,n44_11);
nor I_22(n44_11,IN_3_1_l_11,n40_11);
nand I_23(n45_11,n46_11,n47_11);
not I_24(n46_11,n38_11);
nand I_25(n47_11,n59_11,n62_11);
and I_26(n48_11,n37_11,n47_11);
or I_27(n49_11,n44_11,n50_11);
nor I_28(n50_11,n60_11,n61_11);
or I_29(n51_11,n_102_5_r_11,n52_11);
nor I_30(n52_11,n42_11,n57_11);
nand I_31(n53_11,n37_11,n50_11);
or I_32(n54_11,IN_2_3_l_11,IN_3_3_l_11);
nor I_33(n55_11,n38_11,n42_11);
not I_34(n56_11,N1372_10_r_11);
and I_35(n57_11,n38_11,n50_11);
and I_36(n58_11,IN_1_6_l_11,n59_11);
or I_37(n59_11,IN_5_6_l_11,n63_11);
not I_38(n60_11,IN_1_0_l_11);
nor I_39(n61_11,IN_3_0_l_11,IN_4_0_l_11);
nand I_40(n62_11,IN_3_6_l_11,IN_4_6_l_11);
and I_41(n63_11,IN_3_6_l_11,IN_4_6_l_11);
nor I_42(N1371_0_r_2,n32_2,n35_2);
nor I_43(N1508_0_r_2,n32_2,n55_2);
not I_44(N1372_1_r_2,n54_2);
nor I_45(N1508_1_r_2,n59_2,n54_2);
nor I_46(N6147_2_r_2,n42_2,n43_2);
nor I_47(N1507_6_r_2,n40_2,n53_2);
nor I_48(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_49(n4_7_r_2,blif_clk_net_7_r_2,n10_2,G42_7_r_2,);
nor I_50(n_572_7_r_2,n36_2,n37_2);
or I_51(n_573_7_r_2,n34_2,n35_2);
nor I_52(n_549_7_r_2,n40_2,n41_2);
nand I_53(n_569_7_r_2,n38_2,n39_2);
nor I_54(n_452_7_r_2,n59_2,n35_2);
nor I_55(n4_7_l_2,N6147_2_r_11,n_576_5_r_11);
not I_56(n10_2,blif_reset_net_7_r_2);
DFFARX1 I_57(n4_7_l_2,blif_clk_net_7_r_2,n10_2,n59_2,);
not I_58(n33_2,n59_2);
and I_59(N3_8_l_2,n49_2,G78_5_r_11);
DFFARX1 I_60(N3_8_l_2,blif_clk_net_7_r_2,n10_2,n32_internal_2,);
not I_61(n32_2,n32_internal_2);
nor I_62(n4_7_r_2,n59_2,n36_2);
not I_63(n34_2,n39_2);
nor I_64(n35_2,N1508_6_r_11,N1372_1_r_11);
nor I_65(n36_2,n_576_5_r_11,N6147_2_r_11);
or I_66(n37_2,N1507_6_r_11,N1508_10_r_11);
not I_67(n38_2,n40_2);
nand I_68(n39_2,n45_2,n57_2);
nor I_69(n40_2,n47_2,N1372_1_r_11);
nor I_70(n41_2,n32_2,n36_2);
not I_71(n42_2,n53_2);
nand I_72(n43_2,n44_2,n45_2);
nand I_73(n44_2,n38_2,n46_2);
not I_74(n45_2,N1508_10_r_11);
nand I_75(n46_2,n47_2,n48_2);
nand I_76(n47_2,n_429_or_0_5_r_11,n_547_5_r_11);
or I_77(n48_2,N1508_1_r_11,N6147_3_r_11);
nand I_78(n49_2,N6147_3_r_11,N1508_6_r_11);
nand I_79(n50_2,n51_2,n52_2);
not I_80(n51_2,n47_2);
nand I_81(n52_2,n38_2,n53_2);
nor I_82(n53_2,N1507_6_r_11,N6147_2_r_11);
nand I_83(n54_2,n42_2,n56_2);
nor I_84(n55_2,n34_2,n56_2);
nor I_85(n56_2,N1508_1_r_11,N6147_3_r_11);
nand I_86(n57_2,n58_2,N1508_1_r_11);
not I_87(n58_2,N6147_3_r_11);
endmodule


