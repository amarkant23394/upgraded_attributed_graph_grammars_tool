module test_final(G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_3,blif_reset_net_1_r_3,G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3);
input G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_3,blif_reset_net_1_r_3;
output G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3;
wire G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4,n_431_0_l_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n4_1_l_3,n9_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3;
DFFARX1 I_0(n4_1_r_4,blif_clk_net_1_r_3,n9_3,G42_1_r_4,);
nor I_1(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_2(n_573_1_r_4,G2_0_l_4,n16_4);
nor I_3(n_549_1_r_4,n22_4,n23_4);
nand I_4(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_5(n19_4,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_4,);
nor I_6(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_7(n19_4,blif_clk_net_1_r_3,n9_3,ACVQN1_5_r_4,);
not I_8(P6_5_r_4,P6_5_r_internal_4);
or I_9(n_431_0_l_4,IN_8_0_l_4,n26_4);
DFFARX1 I_10(n_431_0_l_4,blif_clk_net_1_r_3,n9_3,G78_0_l_4,);
DFFARX1 I_11(IN_2_5_l_4,blif_clk_net_1_r_3,n9_3,ACVQN1_5_l_4,);
not I_12(n16_4,ACVQN1_5_l_4);
DFFARX1 I_13(IN_1_5_l_4,blif_clk_net_1_r_3,n9_3,n17_internal_4,);
not I_14(n17_4,n17_internal_4);
nor I_15(n4_1_r_4,n30_4,n31_4);
nand I_16(n19_4,G1_0_l_4,n33_4);
DFFARX1 I_17(G78_0_l_4,blif_clk_net_1_r_3,n9_3,n15_internal_4,);
not I_18(n15_4,n15_internal_4);
DFFARX1 I_19(ACVQN1_5_l_4,blif_clk_net_1_r_3,n9_3,P6_5_r_internal_4,);
and I_20(n20_4,IN_11_0_l_4,n16_4);
nor I_21(n21_4,G2_0_l_4,IN_10_0_l_4);
nand I_22(n22_4,G78_0_l_4,n25_4);
nand I_23(n23_4,IN_11_0_l_4,n24_4);
not I_24(n24_4,G2_0_l_4);
not I_25(n25_4,IN_10_0_l_4);
and I_26(n26_4,IN_2_0_l_4,n27_4);
nor I_27(n27_4,IN_4_0_l_4,n28_4);
not I_28(n28_4,G1_0_l_4);
not I_29(n29_4,n30_4);
nand I_30(n30_4,IN_7_0_l_4,n32_4);
nand I_31(n31_4,IN_11_0_l_4,n25_4);
nor I_32(n32_4,G2_0_l_4,n33_4);
not I_33(n33_4,IN_5_0_l_4);
DFFARX1 I_34(n4_1_r_3,blif_clk_net_1_r_3,n9_3,G42_1_r_3,);
nor I_35(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_36(n_573_1_r_3,n26_3,n27_3);
nor I_37(n_549_1_r_3,n40_3,n32_3);
nand I_38(n_569_1_r_3,n27_3,n31_3);
and I_39(n_452_1_r_3,n26_3,n_569_1_r_4);
nor I_40(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_41(N3_2_r_3,blif_clk_net_1_r_3,n9_3,G199_2_r_3,);
DFFARX1 I_42(n_572_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_3,);
nor I_43(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_44(n4_1_l_3,n_569_1_r_4,n_266_and_0_3_r_4);
not I_45(n9_3,blif_reset_net_1_r_3);
DFFARX1 I_46(n4_1_l_3,blif_clk_net_1_r_3,n9_3,G42_1_l_3,);
not I_47(n22_3,G42_1_l_3);
DFFARX1 I_48(n_573_1_r_4,blif_clk_net_1_r_3,n9_3,n40_3,);
DFFARX1 I_49(G42_1_r_4,blif_clk_net_1_r_3,n9_3,n25_internal_3,);
not I_50(n25_3,n25_internal_3);
nor I_51(n4_1_r_3,n40_3,n36_3);
nor I_52(N3_2_r_3,n26_3,n37_3);
nor I_53(n_572_1_l_3,ACVQN2_3_r_4,P6_5_r_4);
DFFARX1 I_54(G42_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN1_3_r_3,);
nor I_55(n26_3,n_549_1_r_4,n_572_1_r_4);
not I_56(n27_3,ACVQN1_5_r_4);
nor I_57(n28_3,n29_3,ACVQN1_5_r_4);
nor I_58(n29_3,n30_3,ACVQN2_3_r_4);
not I_59(n30_3,n_572_1_r_4);
nor I_60(n31_3,n40_3,n_549_1_r_4);
nor I_61(n32_3,n25_3,n33_3);
nand I_62(n33_3,n22_3,G42_1_r_4);
or I_63(n34_3,n_549_1_r_4,ACVQN1_5_r_4);
nand I_64(n35_3,ACVQN1_3_r_3,G42_1_r_4);
nor I_65(n36_3,n_569_1_r_4,n_572_1_r_4);
nor I_66(n37_3,n38_3,n39_3);
not I_67(n38_3,n_572_1_l_3);
nand I_68(n39_3,n27_3,n30_3);
endmodule


