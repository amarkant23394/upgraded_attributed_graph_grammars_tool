module test_I8839(I6893,I1477,I1470,I8839);
input I6893,I1477,I1470;
output I8839;
wire I9320,I7190,I8896,I6875,I8913,I6872,I9303,I8862,I9337,I6878;
not I_0(I9320,I9303);
DFFARX1 I_1(I1470,,,I7190,);
DFFARX1 I_2(I9337,I1470,I8862,,,I8839,);
nor I_3(I8896,I6893,I6872);
DFFARX1 I_4(I1470,,,I6875,);
nand I_5(I8913,I8896,I6878);
DFFARX1 I_6(I1470,,,I6872,);
DFFARX1 I_7(I6875,I1470,I8862,,,I9303,);
not I_8(I8862,I1477);
nor I_9(I9337,I9320,I8913);
not I_10(I6878,I7190);
endmodule


