module test_I16339(I14438,I1477,I14520,I1470,I16339);
input I14438,I1477,I14520,I1470;
output I16339;
wire I14338,I13361,I13162,I14537,I14472,I13248,I14455,I14353,I14808,I14605,I14370;
DFFARX1 I_0(I14605,I1470,I14370,,,I14338,);
DFFARX1 I_1(I1470,,,I13361,);
and I_2(I13162,I13248,I13361);
DFFARX1 I_3(I14520,I1470,I14370,,,I14537,);
nor I_4(I16339,I14353,I14338);
nand I_5(I14472,I14455,I14438);
DFFARX1 I_6(I1470,,,I13248,);
DFFARX1 I_7(I1470,I14370,,,I14455,);
not I_8(I14353,I14808);
DFFARX1 I_9(I13162,I1470,I14370,,,I14808,);
and I_10(I14605,I14537,I14472);
not I_11(I14370,I1477);
endmodule


