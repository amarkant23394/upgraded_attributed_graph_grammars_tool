module test_I7492(I5659,I7139,I1477,I6992,I1470,I7492);
input I5659,I7139,I1477,I6992,I1470;
output I7492;
wire I7173,I7009,I5073,I7156,I5594,I7238,I7427,I5088,I7410,I6907,I5082,I7221,I5105,I6924;
nor I_0(I7173,I7156,I7009);
not I_1(I7009,I6992);
DFFARX1 I_2(I1470,I5105,,,I5073,);
DFFARX1 I_3(I7139,I1470,I6907,,,I7156,);
DFFARX1 I_4(I1470,I5105,,,I5594,);
and I_5(I7238,I7221,I7173);
not I_6(I7427,I7410);
DFFARX1 I_7(I5659,I1470,I5105,,,I5088,);
DFFARX1 I_8(I5082,I1470,I6907,,,I7410,);
not I_9(I6907,I1477);
not I_10(I5082,I5594);
nand I_11(I7221,I6924,I5088);
not I_12(I5105,I1477);
not I_13(I6924,I5073);
or I_14(I7492,I7427,I7238);
endmodule


