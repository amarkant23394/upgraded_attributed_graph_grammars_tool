module test_I16435(I1477,I13296,I14404,I1470,I13508,I16435);
input I1477,I13296,I14404,I1470,I13508;
output I16435;
wire I14667,I13177,I14455,I14421,I14715,I14350,I13601,I13186,I14650,I13165,I14359,I14370,I13197,I13542,I13635,I13159,I14438,I13189,I14732;
and I_0(I14667,I14650,I13189);
nand I_1(I13177,I13296,I13542);
DFFARX1 I_2(I13177,I1470,I14370,,,I14455,);
DFFARX1 I_3(I14404,I1470,I14370,,,I14421,);
nand I_4(I16435,I14359,I14350);
not I_5(I14715,I14667);
nand I_6(I14350,I14455,I14732);
DFFARX1 I_7(I1470,I13197,,,I13601,);
nor I_8(I13186,I13601,I13508);
DFFARX1 I_9(I13165,I1470,I14370,,,I14650,);
DFFARX1 I_10(I1470,I13197,,,I13165,);
nor I_11(I14359,I14667,I14438);
not I_12(I14370,I1477);
not I_13(I13197,I1477);
nor I_14(I13542,I13508);
and I_15(I13635,I13296);
DFFARX1 I_16(I13508,I1470,I13197,,,I13159,);
nor I_17(I14438,I13159,I13186);
DFFARX1 I_18(I13635,I1470,I13197,,,I13189,);
nor I_19(I14732,I14421,I14715);
endmodule


