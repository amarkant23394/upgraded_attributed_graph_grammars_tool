module test_I8854(I1477,I5070,I1470,I7221,I5097,I8854);
input I1477,I5070,I1470,I7221,I5097;
output I8854;
wire I9320,I6875,I6992,I6975,I7026,I9303,I9179,I8862,I6907,I6896;
not I_0(I9320,I9303);
DFFARX1 I_1(I7221,I1470,I6907,,,I6875,);
nor I_2(I8854,I9179,I9320);
nand I_3(I6992,I6975,I5097);
nor I_4(I6975,I5070);
not I_5(I7026,I5070);
DFFARX1 I_6(I6875,I1470,I8862,,,I9303,);
DFFARX1 I_7(I6896,I1470,I8862,,,I9179,);
not I_8(I8862,I1477);
not I_9(I6907,I1477);
nor I_10(I6896,I6992,I7026);
endmodule


