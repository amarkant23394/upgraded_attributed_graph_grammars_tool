module test_final(IN_1_2_l_2,IN_2_2_l_2,G1_3_l_2,G2_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_5_3_l_2,IN_7_3_l_2,IN_8_3_l_2,IN_10_3_l_2,IN_11_3_l_2,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G199_1_r_9,G214_1_r_9,ACVQN1_2_r_9,P6_2_r_9,n_429_or_0_3_r_9,G78_3_r_9,n_576_3_r_9,n_102_3_r_9,n_547_3_r_9,n_42_5_r_9,G199_5_r_9);
input IN_1_2_l_2,IN_2_2_l_2,G1_3_l_2,G2_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_5_3_l_2,IN_7_3_l_2,IN_8_3_l_2,IN_10_3_l_2,IN_11_3_l_2,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G199_1_r_9,G214_1_r_9,ACVQN1_2_r_9,P6_2_r_9,n_429_or_0_3_r_9,G78_3_r_9,n_576_3_r_9,n_102_3_r_9,n_547_3_r_9,n_42_5_r_9,G199_5_r_9;
wire ACVQN2_0_r_2,n_266_and_0_0_r_2,G199_1_r_2,G214_1_r_2,n_429_or_0_3_r_2,G78_3_r_2,n_576_3_r_2,n_102_3_r_2,n_547_3_r_2,n_42_5_r_2,G199_5_r_2,ACVQN1_2_l_2,P6_2_l_2,P6_internal_2_l_2,n_429_or_0_3_l_2,n12_3_l_2,n_431_3_l_2,G78_3_l_2,n_576_3_l_2,n11_3_l_2,n_102_3_l_2,n_547_3_l_2,n13_3_l_2,n14_3_l_2,n15_3_l_2,n16_3_l_2,ACVQN1_0_r_2,N1_1_r_2,n3_1_r_2,n12_3_r_2,n_431_3_r_2,n11_3_r_2,n13_3_r_2,n14_3_r_2,n15_3_r_2,n16_3_r_2,N3_5_r_2,n3_5_r_2,n1_1_r_9,ACVQN2_0_l_9,n_266_and_0_0_l_9,ACVQN1_0_l_9,n4_4_l_9,G42_4_l_9,n_87_4_l_9,n_572_4_l_9,n_573_4_l_9,n_549_4_l_9,n7_4_l_9,n_569_4_l_9,n_452_4_l_9,N1_1_r_9,n3_1_r_9,P6_internal_2_r_9,n12_3_r_9,n_431_3_r_9,n11_3_r_9,n13_3_r_9,n14_3_r_9,n15_3_r_9,n16_3_r_9,N3_5_r_9,n3_5_r_9;
DFFARX1 I_0(P6_2_l_2,blif_clk_net_1_r_9,n1_1_r_9,ACVQN2_0_r_2,);
and I_1(n_266_and_0_0_r_2,n_102_3_l_2,ACVQN1_0_r_2);
DFFARX1 I_2(N1_1_r_2,blif_clk_net_1_r_9,n1_1_r_9,G199_1_r_2,);
DFFARX1 I_3(n_547_3_l_2,blif_clk_net_1_r_9,n1_1_r_9,G214_1_r_2,);
nand I_4(n_429_or_0_3_r_2,ACVQN1_2_l_2,n12_3_r_2);
DFFARX1 I_5(n_431_3_r_2,blif_clk_net_1_r_9,n1_1_r_9,G78_3_r_2,);
nand I_6(n_576_3_r_2,ACVQN1_2_l_2,n11_3_r_2);
not I_7(n_102_3_r_2,G78_3_l_2);
nand I_8(n_547_3_r_2,n_102_3_l_2,n13_3_r_2);
nor I_9(n_42_5_r_2,ACVQN1_2_l_2,P6_2_l_2);
DFFARX1 I_10(N3_5_r_2,blif_clk_net_1_r_9,n1_1_r_9,G199_5_r_2,);
DFFARX1 I_11(IN_2_2_l_2,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_2_l_2,);
not I_12(P6_2_l_2,P6_internal_2_l_2);
DFFARX1 I_13(IN_1_2_l_2,blif_clk_net_1_r_9,n1_1_r_9,P6_internal_2_l_2,);
nand I_14(n_429_or_0_3_l_2,G1_3_l_2,n12_3_l_2);
not I_15(n12_3_l_2,IN_5_3_l_2);
or I_16(n_431_3_l_2,IN_8_3_l_2,n14_3_l_2);
DFFARX1 I_17(n_431_3_l_2,blif_clk_net_1_r_9,n1_1_r_9,G78_3_l_2,);
nand I_18(n_576_3_l_2,IN_7_3_l_2,n11_3_l_2);
nor I_19(n11_3_l_2,G2_3_l_2,n12_3_l_2);
not I_20(n_102_3_l_2,G2_3_l_2);
nand I_21(n_547_3_l_2,IN_11_3_l_2,n13_3_l_2);
nor I_22(n13_3_l_2,G2_3_l_2,IN_10_3_l_2);
and I_23(n14_3_l_2,IN_2_3_l_2,n15_3_l_2);
nor I_24(n15_3_l_2,IN_4_3_l_2,n16_3_l_2);
not I_25(n16_3_l_2,G1_3_l_2);
DFFARX1 I_26(G78_3_l_2,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_0_r_2,);
and I_27(N1_1_r_2,G78_3_l_2,n3_1_r_2);
nand I_28(n3_1_r_2,n_576_3_l_2,n_547_3_l_2);
not I_29(n12_3_r_2,n_429_or_0_3_l_2);
or I_30(n_431_3_r_2,n_429_or_0_3_l_2,n14_3_r_2);
nor I_31(n11_3_r_2,G78_3_l_2,n12_3_r_2);
nor I_32(n13_3_r_2,G78_3_l_2,n_576_3_l_2);
and I_33(n14_3_r_2,n_576_3_l_2,n15_3_r_2);
nor I_34(n15_3_r_2,P6_2_l_2,n16_3_r_2);
not I_35(n16_3_r_2,ACVQN1_2_l_2);
and I_36(N3_5_r_2,n_102_3_l_2,n3_5_r_2);
nand I_37(n3_5_r_2,ACVQN1_2_l_2,n_429_or_0_3_l_2);
DFFARX1 I_38(N1_1_r_9,blif_clk_net_1_r_9,n1_1_r_9,G199_1_r_9,);
DFFARX1 I_39(G42_4_l_9,blif_clk_net_1_r_9,n1_1_r_9,G214_1_r_9,);
DFFARX1 I_40(n_572_4_l_9,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_2_r_9,);
not I_41(P6_2_r_9,P6_internal_2_r_9);
nand I_42(n_429_or_0_3_r_9,n_572_4_l_9,n12_3_r_9);
DFFARX1 I_43(n_431_3_r_9,blif_clk_net_1_r_9,n1_1_r_9,G78_3_r_9,);
nand I_44(n_576_3_r_9,n_573_4_l_9,n11_3_r_9);
not I_45(n_102_3_r_9,n_266_and_0_0_l_9);
nand I_46(n_547_3_r_9,n_549_4_l_9,n13_3_r_9);
nor I_47(n_42_5_r_9,n_569_4_l_9,n_452_4_l_9);
DFFARX1 I_48(N3_5_r_9,blif_clk_net_1_r_9,n1_1_r_9,G199_5_r_9,);
not I_49(n1_1_r_9,blif_reset_net_1_r_9);
DFFARX1 I_50(n_576_3_r_2,blif_clk_net_1_r_9,n1_1_r_9,ACVQN2_0_l_9,);
and I_51(n_266_and_0_0_l_9,ACVQN1_0_l_9,G78_3_r_2);
DFFARX1 I_52(G199_5_r_2,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_0_l_9,);
nor I_53(n4_4_l_9,G199_1_r_2,n_102_3_r_2);
DFFARX1 I_54(n4_4_l_9,blif_clk_net_1_r_9,n1_1_r_9,G42_4_l_9,);
not I_55(n_87_4_l_9,n_42_5_r_2);
nor I_56(n_572_4_l_9,n_266_and_0_0_r_2,n_42_5_r_2);
or I_57(n_573_4_l_9,G214_1_r_2,n_429_or_0_3_r_2);
nor I_58(n_549_4_l_9,n7_4_l_9,ACVQN2_0_r_2);
and I_59(n7_4_l_9,n_87_4_l_9,n_547_3_r_2);
or I_60(n_569_4_l_9,ACVQN2_0_r_2,G214_1_r_2);
nor I_61(n_452_4_l_9,n_429_or_0_3_r_2,n_102_3_r_2);
and I_62(N1_1_r_9,n_266_and_0_0_l_9,n3_1_r_9);
nand I_63(n3_1_r_9,n_572_4_l_9,n_569_4_l_9);
DFFARX1 I_64(n_266_and_0_0_l_9,blif_clk_net_1_r_9,n1_1_r_9,P6_internal_2_r_9,);
not I_65(n12_3_r_9,G42_4_l_9);
or I_66(n_431_3_r_9,n_549_4_l_9,n14_3_r_9);
nor I_67(n11_3_r_9,ACVQN2_0_l_9,n12_3_r_9);
nor I_68(n13_3_r_9,ACVQN2_0_l_9,n_266_and_0_0_l_9);
and I_69(n14_3_r_9,n_452_4_l_9,n15_3_r_9);
nor I_70(n15_3_r_9,G42_4_l_9,n16_3_r_9);
not I_71(n16_3_r_9,n_572_4_l_9);
and I_72(N3_5_r_9,ACVQN2_0_l_9,n3_5_r_9);
nand I_73(n3_5_r_9,n_573_4_l_9,n_452_4_l_9);
endmodule


