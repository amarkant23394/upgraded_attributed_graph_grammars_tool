module test_I5097(I1477,I5122,I3380,I1470,I3453,I5317,I5097);
input I1477,I5122,I3380,I1470,I3453,I5317;
output I5097;
wire I3747,I5105,I5351,I3362,I5187,I5334,I5625,I5368,I3353,I3637,I3377,I5204,I5642;
DFFARX1 I_0(I1470,,,I3747,);
not I_1(I5105,I1477);
DFFARX1 I_2(I5334,I1470,I5105,,,I5351,);
DFFARX1 I_3(I1470,,,I3362,);
nor I_4(I5187,I5122,I3380);
or I_5(I5334,I5317,I3362);
DFFARX1 I_6(I3377,I1470,I5105,,,I5625,);
nor I_7(I5368,I5351,I5204);
and I_8(I3353,I3453,I3637);
DFFARX1 I_9(I1470,,,I3637,);
not I_10(I3377,I3747);
nand I_11(I5097,I5642,I5368);
nand I_12(I5204,I5187,I3353);
not I_13(I5642,I5625);
endmodule


