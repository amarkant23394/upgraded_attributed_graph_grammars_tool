module test_I17871(I1477,I13749,I16069,I15696,I15628,I1470,I17871);
input I1477,I13749,I16069,I15696,I15628,I1470;
output I17871;
wire I17413,I17854,I15585,I15832,I17532,I15815,I15959,I15928,I15597,I15588,I17775,I16145,I16162,I17447,I15594,I17464;
not I_0(I17413,I1477);
nand I_1(I17854,I17775,I17464);
and I_2(I17871,I17532,I17854);
nand I_3(I15585,I16069,I15959);
nand I_4(I15832,I15628,I13749);
not I_5(I17532,I15597);
DFFARX1 I_6(I1470,,,I15815,);
nor I_7(I15959,I15928,I15696);
DFFARX1 I_8(I1470,,,I15928,);
nor I_9(I15597,I15832,I16162);
DFFARX1 I_10(I1470,,,I15588,);
DFFARX1 I_11(I15585,I1470,I17413,,,I17775,);
not I_12(I16145,I16069);
and I_13(I16162,I15696,I16145);
nor I_14(I17447,I15597,I15588);
or I_15(I15594,I15928,I15815);
nand I_16(I17464,I17447,I15594);
endmodule


