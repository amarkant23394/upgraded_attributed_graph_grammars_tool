module test_I3124(I1351,I1447,I1477,I1470,I3124);
input I1351,I1447,I1477,I1470;
output I3124;
wire I2878,I2759,I3076,I2861;
not I_0(I2878,I2861);
not I_1(I2759,I1477);
nor I_2(I3124,I3076,I2878);
DFFARX1 I_3(I1447,I1470,I2759,,,I3076,);
not I_4(I2861,I1351);
endmodule


