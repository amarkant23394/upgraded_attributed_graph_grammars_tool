module test_final(IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_5_r_13,blif_reset_net_5_r_13,N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13);
input IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_5_r_13,blif_reset_net_5_r_13;
output N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13;
wire N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_549_7_r_5,n_569_7_r_5,n_452_7_r_5,n4_7_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5,n_102_5_r_13,n4_7_l_13,n9_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13;
nor I_0(N1371_0_r_5,n28_5,n46_5);
nand I_1(N1508_0_r_5,n26_5,n43_5);
not I_2(N1372_1_r_5,n43_5);
nor I_3(N1508_1_r_5,n30_5,n43_5);
nor I_4(N6147_2_r_5,n29_5,n32_5);
nor I_5(N1507_6_r_5,n26_5,n44_5);
nor I_6(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_7(n4_7_r_5,blif_clk_net_5_r_13,n9_13,G42_7_r_5,);
and I_8(n_572_7_r_5,n27_5,n28_5);
nand I_9(n_573_7_r_5,n26_5,n27_5);
nand I_10(n_549_7_r_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_11(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_12(n_452_7_r_5,n29_5);
nor I_13(n4_7_r_5,n30_5,n31_5);
not I_14(n26_5,n35_5);
nand I_15(n27_5,n40_5,n41_5);
nand I_16(n28_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_17(n29_5,n27_5,n33_5);
nor I_18(n30_5,IN_1_3_l_5,n45_5);
not I_19(n31_5,n_549_7_r_5);
nor I_20(n32_5,n34_5,n35_5);
not I_21(n33_5,n30_5);
nor I_22(n34_5,n31_5,n36_5);
nor I_23(n35_5,IN_3_1_l_5,n28_5);
not I_24(n36_5,n28_5);
nand I_25(n37_5,n36_5,n38_5);
nand I_26(n38_5,n26_5,n39_5);
nand I_27(n39_5,n30_5,n31_5);
nor I_28(n40_5,IN_1_2_l_5,IN_2_2_l_5);
or I_29(n41_5,IN_5_2_l_5,n42_5);
nor I_30(n42_5,IN_3_2_l_5,IN_4_2_l_5);
nand I_31(n43_5,n36_5,n46_5);
nor I_32(n44_5,n_549_7_r_5,n33_5);
or I_33(n45_5,IN_2_3_l_5,IN_3_3_l_5);
and I_34(n46_5,n31_5,n47_5);
or I_35(n47_5,IN_3_10_l_5,IN_4_10_l_5);
nor I_36(N1371_0_r_13,n59_13,n61_13);
nor I_37(N1508_0_r_13,n59_13,n60_13);
not I_38(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_39(n_431_5_r_13,blif_clk_net_5_r_13,n9_13,G78_5_r_13,);
nand I_40(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_41(n_102_5_r_13,N6147_2_r_5,n_452_7_r_5);
nand I_42(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_43(n1_13,blif_clk_net_5_r_13,n9_13,G42_7_r_13,);
nor I_44(n_572_7_r_13,n40_13,n41_13);
nand I_45(n_573_7_r_13,n37_13,n38_13);
nor I_46(n_549_7_r_13,n46_13,n47_13);
nand I_47(n_569_7_r_13,n37_13,n43_13);
nand I_48(n_452_7_r_13,n52_13,n53_13);
nor I_49(n4_7_l_13,N1371_0_r_5,N1508_0_r_5);
not I_50(n9_13,blif_reset_net_5_r_13);
DFFARX1 I_51(n4_7_l_13,blif_clk_net_5_r_13,n9_13,n62_13,);
not I_52(n33_13,n62_13);
nand I_53(n_431_5_r_13,n54_13,n55_13);
not I_54(n1_13,n52_13);
nor I_55(n34_13,n35_13,n36_13);
nor I_56(n35_13,n42_13,N1508_6_r_5);
nand I_57(n36_13,n50_13,n58_13);
nand I_58(n37_13,n44_13,n45_13);
or I_59(n38_13,n39_13,N1372_1_r_5);
nand I_60(n39_13,N1508_0_r_5,n_573_7_r_5);
not I_61(n40_13,n36_13);
nor I_62(n41_13,n35_13,N6147_2_r_5);
not I_63(n42_13,N1508_1_r_5);
or I_64(n43_13,N1508_1_r_5,N1371_0_r_5);
not I_65(n44_13,N1508_6_r_5);
not I_66(n45_13,n_572_7_r_5);
nor I_67(n46_13,n39_13,n40_13);
nor I_68(n47_13,N1508_1_r_5,N1371_0_r_5);
nor I_69(n48_13,n50_13,n51_13);
nor I_70(n49_13,N1508_6_r_5,n_572_7_r_5);
not I_71(n50_13,n59_13);
not I_72(n51_13,n_102_5_r_13);
nand I_73(n52_13,n33_13,n39_13);
nand I_74(n53_13,n33_13,N1372_1_r_5);
nor I_75(n54_13,N1508_1_r_5,n_452_7_r_5);
nand I_76(n55_13,n62_13,n56_13);
nor I_77(n56_13,n39_13,n57_13);
not I_78(n57_13,N1371_0_r_5);
or I_79(n58_13,n_569_7_r_5,N1372_1_r_5);
nand I_80(n59_13,N1507_6_r_5,G42_7_r_5);
nor I_81(n60_13,n51_13,N1508_1_r_5);
nor I_82(n61_13,n39_13,N1372_1_r_5);
endmodule


