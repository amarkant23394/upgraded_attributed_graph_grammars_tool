module test_I11284(I8830,I9049,I8862,I6881,I8879,I1470,I9413,I11284);
input I8830,I9049,I8862,I6881,I8879,I1470,I9413;
output I11284;
wire I11378,I11429,I9066,I11395,I11460,I8848,I11327,I9083,I8851;
nor I_0(I11378,I11327,I8848);
not I_1(I11429,I8848);
DFFARX1 I_2(I9049,I1470,I8862,,,I9066,);
nand I_3(I11395,I11378,I8851);
nand I_4(I11284,I11395,I11460);
not I_5(I11460,I11429);
nor I_6(I8848,I9083,I9413);
not I_7(I11327,I8830);
nand I_8(I9083,I8879,I6881);
or I_9(I8851,I9083,I9066);
endmodule


