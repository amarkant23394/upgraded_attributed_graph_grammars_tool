module test_I12075(I10349,I10032,I1477,I1470,I10202,I12075);
input I10349,I10032,I1477,I1470,I10202;
output I12075;
wire I10219,I12041,I10052,I10020,I10397,I12058,I11990,I11973,I10287,I10026;
DFFARX1 I_0(I10202,I1470,I10052,,,I10219,);
nor I_1(I12041,I11990,I10020);
not I_2(I10052,I1477);
DFFARX1 I_3(I10287,I1470,I10052,,,I10020,);
not I_4(I10397,I10349);
nand I_5(I12058,I12041,I10026);
not I_6(I11990,I10032);
not I_7(I11973,I1477);
and I_8(I10287,I10219);
DFFARX1 I_9(I12058,I1470,I11973,,,I12075,);
nand I_10(I10026,I10219,I10397);
endmodule


