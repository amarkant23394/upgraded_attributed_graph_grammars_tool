module test_final(IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_1_8_l_0,IN_2_8_l_0,IN_3_8_l_0,IN_6_8_l_0,IN_1_10_l_0,IN_2_10_l_0,IN_3_10_l_0,IN_4_10_l_0,blif_clk_net_5_r_5,blif_reset_net_5_r_5,N1371_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1508_6_r_5);
input IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_1_8_l_0,IN_2_8_l_0,IN_3_8_l_0,IN_6_8_l_0,IN_1_10_l_0,IN_2_10_l_0,IN_3_10_l_0,IN_4_10_l_0,blif_clk_net_5_r_5,blif_reset_net_5_r_5;
output N1371_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1508_6_r_5;
wire N1371_0_r_0,N1508_0_r_0,N6147_2_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,N1507_6_r_0,N1508_6_r_0,N3_8_l_0,n40_0,n4_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,N1508_0_r_5,N1507_6_r_5,n_431_5_r_5,n6_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5;
nor I_0(N1371_0_r_0,n24_0,n25_0);
not I_1(N1508_0_r_0,n25_0);
nor I_2(N6147_2_r_0,n28_0,n29_0);
nand I_3(n_429_or_0_5_r_0,n4_0,n25_0);
DFFARX1 I_4(n4_0,blif_clk_net_5_r_5,n6_5,G78_5_r_0,);
nand I_5(n_576_5_r_0,n23_0,n24_0);
not I_6(n_102_5_r_0,n40_0);
nand I_7(n_547_5_r_0,n26_0,n27_0);
nor I_8(N1507_6_r_0,n_102_5_r_0,n37_0);
nor I_9(N1508_6_r_0,n25_0,n33_0);
and I_10(N3_8_l_0,IN_6_8_l_0,n32_0);
DFFARX1 I_11(N3_8_l_0,blif_clk_net_5_r_5,n6_5,n40_0,);
not I_12(n4_0,n31_0);
nor I_13(n23_0,n40_0,n25_0);
and I_14(n24_0,n4_0,n39_0);
nand I_15(n25_0,IN_1_1_l_0,IN_2_1_l_0);
nor I_16(n26_0,n40_0,n24_0);
nor I_17(n27_0,IN_1_8_l_0,IN_3_8_l_0);
nor I_18(n28_0,IN_3_1_l_0,n25_0);
nand I_19(n29_0,n_102_5_r_0,n30_0);
nand I_20(n30_0,n27_0,n31_0);
nand I_21(n31_0,IN_1_10_l_0,IN_2_10_l_0);
nand I_22(n32_0,IN_2_8_l_0,IN_3_8_l_0);
nand I_23(n33_0,n34_0,n35_0);
nand I_24(n34_0,n_102_5_r_0,n36_0);
not I_25(n35_0,IN_3_1_l_0);
not I_26(n36_0,n27_0);
nor I_27(n37_0,n36_0,n38_0);
nand I_28(n38_0,N1508_0_r_0,n35_0);
or I_29(n39_0,IN_3_10_l_0,IN_4_10_l_0);
nor I_30(N1371_0_r_5,n28_5,n39_5);
not I_31(N1508_0_r_5,n39_5);
nor I_32(N6147_2_r_5,n28_5,n37_5);
nand I_33(n_429_or_0_5_r_5,n30_5,n32_5);
DFFARX1 I_34(n_431_5_r_5,blif_clk_net_5_r_5,n6_5,G78_5_r_5,);
nand I_35(n_576_5_r_5,n26_5,n27_5);
not I_36(n_102_5_r_5,n28_5);
nand I_37(n_547_5_r_5,n31_5,n32_5);
nor I_38(N1507_6_r_5,n30_5,n32_5);
nor I_39(N1508_6_r_5,n39_5,n41_5);
nand I_40(n_431_5_r_5,n34_5,n35_5);
not I_41(n6_5,blif_reset_net_5_r_5);
nor I_42(n26_5,n29_5,n30_5);
nor I_43(n27_5,n28_5,N1371_0_r_0);
nor I_44(n28_5,n29_5,n44_5);
not I_45(n29_5,n_547_5_r_0);
nand I_46(n30_5,N1508_0_r_5,n43_5);
nor I_47(n31_5,n28_5,n33_5);
nor I_48(n32_5,n40_5,N1508_6_r_0);
nor I_49(n33_5,n29_5,N1371_0_r_0);
or I_50(n34_5,n29_5,N1371_0_r_0);
nand I_51(n35_5,n32_5,n36_5);
not I_52(n36_5,n30_5);
nor I_53(n37_5,N1507_6_r_5,n38_5);
and I_54(n38_5,n39_5,n40_5);
nand I_55(n39_5,n_429_or_0_5_r_0,G78_5_r_0);
nand I_56(n40_5,G78_5_r_0,n_576_5_r_0);
nand I_57(n41_5,n28_5,n42_5);
or I_58(n42_5,n32_5,n36_5);
or I_59(n43_5,N6147_2_r_0,N1507_6_r_0);
nor I_60(n44_5,N1371_0_r_0,N6147_2_r_0);
endmodule


