module test_I11287(I11412,I8854,I1477,I1470,I11327,I11287);
input I11412,I8854,I1477,I1470,I11327;
output I11287;
wire I11576,I8827,I11813,I11895,I11830,I11559,I11310,I11641,I11624;
DFFARX1 I_0(I11895,I1470,I11310,,,I11287,);
nor I_1(I11576,I11559,I11412);
DFFARX1 I_2(I1470,,,I8827,);
DFFARX1 I_3(I8854,I1470,I11310,,,I11813,);
or I_4(I11895,I11830,I11641);
not I_5(I11830,I11813);
DFFARX1 I_6(I1470,I11310,,,I11559,);
not I_7(I11310,I1477);
and I_8(I11641,I11624,I11576);
nand I_9(I11624,I11327,I8827);
endmodule


