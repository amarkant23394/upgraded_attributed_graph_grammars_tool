module test_I4544(I1477,I4544);
input I1477;
output I4544;
wire ;
not I_0(I4544,I1477);
endmodule


