module test_I3798(I1477,I1637,I1504,I1603,I1470,I3798);
input I1477,I1637,I1504,I1603,I1470;
output I3798;
wire I3422,I3781,I1507,I3764,I3747,I3685,I1483,I3388,I3668,I1518,I1668,I1928,I1480,I2038,I1880,I1498,I1976,I2021;
or I_0(I3422,I1483,I1480);
nor I_1(I3781,I3422,I3764);
nor I_2(I1507,I1603,I1637);
not I_3(I3764,I3747);
DFFARX1 I_4(I1504,I1470,I3388,,,I3747,);
and I_5(I3685,I3668,I1498);
DFFARX1 I_6(I1880,I1470,I1518,,,I1483,);
not I_7(I3388,I1477);
DFFARX1 I_8(I1507,I1470,I3388,,,I3668,);
not I_9(I1518,I1477);
not I_10(I1668,I1637);
nor I_11(I1928,I1880,I1668);
DFFARX1 I_12(I1976,I1470,I1518,,,I1480,);
not I_13(I2038,I2021);
DFFARX1 I_14(I1470,I1518,,,I1880,);
nand I_15(I1498,I2038,I1928);
and I_16(I3798,I3685,I3781);
and I_17(I1976,I1637);
DFFARX1 I_18(I1470,I1518,,,I2021,);
endmodule


