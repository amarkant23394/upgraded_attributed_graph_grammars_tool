module test_I2457(I1294,I1492,I1639,I1410,I2070,I1301,I1704,I2457);
input I1294,I1492,I1639,I1410,I2070,I1301,I1704;
output I2457;
wire I2313,I2389,I1322,I2087,I2234,I2440,I1427,I2423,I1331,I1954,I2406,I1937,I1342,I1509,I1304;
DFFARX1 I_0(I1331,I1294,I1937,,,I2313,);
DFFARX1 I_1(I1294,I1937,,,I2389,);
nand I_2(I1322,I1427,I1704);
not I_3(I2087,I2070);
nand I_4(I2234,I1954,I1304);
and I_5(I2440,I2313,I2423);
DFFARX1 I_6(I1294,I1342,,,I1427,);
nor I_7(I2423,I2406,I2087);
nor I_8(I1331,I1639,I1410);
not I_9(I1954,I1322);
not I_10(I2406,I2389);
not I_11(I1937,I1301);
not I_12(I1342,I1301);
or I_13(I2457,I2234,I2440);
DFFARX1 I_14(I1492,I1294,I1342,,,I1509,);
DFFARX1 I_15(I1509,I1294,I1342,,,I1304,);
endmodule


