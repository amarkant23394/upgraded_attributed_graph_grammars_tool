module test_I17481(I13908,I15645,I15730,I13743,I13758,I15928,I13764,I16069,I14162,I17481);
input I13908,I15645,I15730,I13743,I13758,I15928,I13764,I16069,I14162;
output I17481;
wire I15662,I13749,I15832,I15579,I15679,I15597,I16145,I16162,I17430,I15696,I15628,I15976;
nand I_0(I15662,I15645,I13764);
nand I_1(I13749,I14162,I13908);
nand I_2(I15832,I15628,I13749);
nand I_3(I15579,I15662,I15976);
nor I_4(I15679,I15628);
nor I_5(I15597,I15832,I16162);
not I_6(I16145,I16069);
and I_7(I16162,I15696,I16145);
not I_8(I17430,I15579);
nand I_9(I15696,I15679,I13758);
not I_10(I15628,I13743);
nor I_11(I15976,I15928,I15730);
nor I_12(I17481,I17430,I15597);
endmodule


