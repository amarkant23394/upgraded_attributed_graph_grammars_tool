module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_5_r_7,blif_reset_net_5_r_7,N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_5_r_7,blif_reset_net_5_r_7;
output N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,n_102_5_r_7,n_452_7_r_7,n4_7_l_7,n6_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_5_r_7,n6_7,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_5_r_7,n6_7,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
nor I_35(N1371_0_r_7,n53_7,n52_7);
nor I_36(N1508_0_r_7,n51_7,n52_7);
nand I_37(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_38(n_431_5_r_7,blif_clk_net_5_r_7,n6_7,G78_5_r_7,);
nand I_39(n_576_5_r_7,n31_7,n32_7);
nor I_40(n_102_5_r_7,N1508_0_r_0,n_429_or_0_5_r_0);
nand I_41(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_42(n4_7_r_7,blif_clk_net_5_r_7,n6_7,G42_7_r_7,);
nor I_43(n_572_7_r_7,n54_7,n33_7);
nand I_44(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_45(n_549_7_r_7,n53_7,n36_7);
nand I_46(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_47(n_452_7_r_7,n_547_5_r_0,n_569_7_r_0);
nor I_48(n4_7_l_7,n_429_or_0_5_r_0,G78_5_r_0);
not I_49(n6_7,blif_reset_net_5_r_7);
DFFARX1 I_50(n4_7_l_7,blif_clk_net_5_r_7,n6_7,n53_7,);
not I_51(n30_7,n53_7);
and I_52(N3_8_l_7,n50_7,N1371_0_r_0);
DFFARX1 I_53(N3_8_l_7,blif_clk_net_5_r_7,n6_7,n54_7,);
nand I_54(n_431_5_r_7,n40_7,n41_7);
nor I_55(n4_7_r_7,n54_7,n49_7);
and I_56(n31_7,n_102_5_r_7,n39_7);
not I_57(n32_7,n_429_or_0_5_r_0);
nor I_58(n33_7,n34_7,n_573_7_r_0);
and I_59(n34_7,n35_7,G42_7_r_0);
not I_60(n35_7,n_576_5_r_0);
nor I_61(n36_7,n37_7,n_429_or_0_5_r_0);
or I_62(n37_7,n54_7,n_429_or_0_5_r_0);
or I_63(n38_7,n_572_7_r_0,n_549_7_r_0);
nor I_64(n39_7,n_452_7_r_7,N1508_0_r_0);
nand I_65(n40_7,n46_7,n47_7);
nand I_66(n41_7,n42_7,n43_7);
nor I_67(n42_7,n44_7,n45_7);
nor I_68(n43_7,n_572_7_r_0,n_549_7_r_0);
nor I_69(n44_7,n_576_5_r_0,N1371_0_r_0);
nor I_70(n45_7,n_573_7_r_0,N1508_0_r_0);
nand I_71(n46_7,n35_7,G42_7_r_0);
not I_72(n47_7,n_573_7_r_0);
or I_73(n48_7,n_452_7_r_7,N1508_0_r_0);
not I_74(n49_7,n_452_7_r_7);
nand I_75(n50_7,n_549_7_r_0,G78_5_r_0);
and I_76(n51_7,n_452_7_r_7,n45_7);
not I_77(n52_7,n44_7);
endmodule


