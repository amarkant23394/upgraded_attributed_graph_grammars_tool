module test_I2751(I1447,I1431,I1477,I1470,I2751);
input I1447,I1431,I1477,I1470;
output I2751;
wire I3217,I2759,I3200,I3076;
not I_0(I3217,I3200);
not I_1(I2759,I1477);
DFFARX1 I_2(I1431,I1470,I2759,,,I3200,);
DFFARX1 I_3(I1447,I1470,I2759,,,I3076,);
nor I_4(I2751,I3076,I3217);
endmodule


