module test_I3543(I2815,I2668,I2234,I1294,I1301,I3543);
input I2815,I2668,I2234,I1294,I1301;
output I3543;
wire I3263,I2962,I2583,I1902,I2203,I2569,I2566,I2945,I2832;
not I_0(I3263,I2569);
nor I_1(I2962,I2945,I2668);
not I_2(I2583,I1301);
and I_3(I1902,I2234,I2203);
DFFARX1 I_4(I1294,,,I2203,);
nand I_5(I2569,I2832,I2962);
not I_6(I2566,I2945);
DFFARX1 I_7(I1902,I1294,I2583,,,I2945,);
nand I_8(I3543,I3263,I2566);
DFFARX1 I_9(I2815,I1294,I2583,,,I2832,);
endmodule


