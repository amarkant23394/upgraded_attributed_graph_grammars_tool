module test_final(IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_7_r_12,blif_reset_net_7_r_12,N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12);
input IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_7_r_12,blif_reset_net_7_r_12;
output N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12;
wire N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,n_429_or_0_5_r_9,G78_5_r_9,n_576_5_r_9,n_102_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9,n_573_7_r_12,n_452_7_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n8_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12;
nor I_0(N6147_2_r_9,n62_9,n46_9);
not I_1(N1372_4_r_9,n59_9);
nor I_2(N1508_4_r_9,n58_9,n59_9);
nand I_3(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_4(n_431_5_r_9,blif_clk_net_7_r_12,n8_12,G78_5_r_9,);
nand I_5(n_576_5_r_9,n39_9,n40_9);
not I_6(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_7(n_547_5_r_9,IN_3_1_l_9,n43_9);
and I_8(n_42_8_r_9,G18_7_l_9,n44_9);
DFFARX1 I_9(N3_8_r_9,blif_clk_net_7_r_12,n8_12,G199_8_r_9,);
nor I_10(N6147_9_r_9,n41_9,n45_9);
nor I_11(N6134_9_r_9,n45_9,n51_9);
nor I_12(I_BUFF_1_9_r_9,IN_3_1_l_9,n41_9);
nor I_13(n4_7_l_9,G18_7_l_9,IN_1_7_l_9);
DFFARX1 I_14(n4_7_l_9,blif_clk_net_7_r_12,n8_12,n62_9,);
and I_15(N3_8_l_9,IN_6_8_l_9,n57_9);
DFFARX1 I_16(N3_8_l_9,blif_clk_net_7_r_12,n8_12,n63_9,);
not I_17(n38_9,n63_9);
nor I_18(n_431_5_r_9,G15_7_l_9,IN_7_7_l_9);
nor I_19(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_20(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_21(n40_9,n41_9);
nand I_22(n41_9,IN_1_1_l_9,IN_2_1_l_9);
nor I_23(n42_9,IN_9_7_l_9,IN_10_7_l_9);
nor I_24(n43_9,n63_9,n41_9);
nor I_25(n44_9,IN_5_7_l_9,IN_9_7_l_9);
and I_26(n45_9,IN_4_7_l_9,n52_9);
nor I_27(n46_9,n47_9,n48_9);
nor I_28(n47_9,n49_9,n50_9);
not I_29(n48_9,n_429_or_0_5_r_9);
not I_30(n49_9,n42_9);
or I_31(n50_9,n63_9,n51_9);
nor I_32(n51_9,IN_1_8_l_9,IN_3_8_l_9);
nor I_33(n52_9,G15_7_l_9,n49_9);
nor I_34(n53_9,n54_9,n55_9);
nor I_35(n54_9,G15_7_l_9,n56_9);
or I_36(n55_9,IN_10_7_l_9,n44_9);
not I_37(n56_9,IN_4_7_l_9);
nand I_38(n57_9,IN_2_8_l_9,IN_3_8_l_9);
nor I_39(n58_9,n62_9,n60_9);
nand I_40(n59_9,n51_9,n61_9);
nor I_41(n60_9,n38_9,n44_9);
nor I_42(n61_9,G18_7_l_9,IN_5_7_l_9);
nor I_43(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_44(N1508_0_r_12,n30_12,n37_12);
nor I_45(N1507_6_r_12,n25_12,n39_12);
nor I_46(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_47(n1_12,blif_clk_net_7_r_12,n8_12,G42_7_r_12,);
nor I_48(n_572_7_r_12,n23_12,n24_12);
nand I_49(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_50(n_549_7_r_12,n27_12,n28_12);
nand I_51(n_569_7_r_12,n25_12,n26_12);
nand I_52(n_452_7_r_12,G199_8_r_9,N1372_4_r_9);
nand I_53(N6147_9_r_12,n30_12,n31_12);
nor I_54(N6134_9_r_12,n35_12,n36_12);
not I_55(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_56(n1_12,n_573_7_r_12);
not I_57(n8_12,blif_reset_net_7_r_12);
not I_58(n23_12,n36_12);
nor I_59(n24_12,n_452_7_r_12,n_576_5_r_9);
nand I_60(n25_12,n23_12,n40_12);
not I_61(n26_12,n35_12);
not I_62(n27_12,N6134_9_r_12);
nand I_63(n28_12,n26_12,n29_12);
not I_64(n29_12,n24_12);
nand I_65(n30_12,n33_12,n41_12);
nand I_66(n31_12,n32_12,n33_12);
nor I_67(n32_12,n26_12,n34_12);
nor I_68(n33_12,N1508_4_r_9,G78_5_r_9);
nor I_69(n34_12,n42_12,n_547_5_r_9);
nor I_70(n35_12,n38_12,N1372_4_r_9);
nand I_71(n36_12,G78_5_r_9,n_576_5_r_9);
nand I_72(n37_12,n23_12,n35_12);
or I_73(n38_12,N6147_9_r_9,N1508_4_r_9);
not I_74(n39_12,n30_12);
or I_75(n40_12,N6147_2_r_9,N6134_9_r_9);
nor I_76(n41_12,n34_12,n36_12);
nor I_77(n42_12,n_42_8_r_9,N6147_2_r_9);
endmodule


