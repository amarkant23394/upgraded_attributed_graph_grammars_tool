module test_I1543(I1231,I1271,I1255,I1207,I1543);
input I1231,I1271,I1255,I1207;
output I1543;
wire I1492,I1526,I1509;
or I_0(I1543,I1526,I1255);
not I_1(I1492,I1207);
and I_2(I1526,I1509,I1271);
nor I_3(I1509,I1492,I1231);
endmodule


