module test_I17679(I17430,I1477,I15832,I1470,I17611,I17679);
input I17430,I1477,I15832,I1470,I17611;
output I17679;
wire I15582,I17413,I17498,I15597,I17515,I17628,I15600,I15815,I17645,I15573,I17481,I17662,I15928;
not I_0(I15582,I15928);
not I_1(I17413,I1477);
nand I_2(I17498,I17481,I15600);
nor I_3(I15597,I15832);
not I_4(I17515,I17498);
and I_5(I17628,I17611,I15573);
or I_6(I15600,I15832,I15815);
DFFARX1 I_7(I1470,,,I15815,);
or I_8(I17645,I17628,I15582);
nor I_9(I17679,I17662,I17515);
nand I_10(I15573,I15832);
nor I_11(I17481,I17430,I15597);
DFFARX1 I_12(I17645,I1470,I17413,,,I17662,);
DFFARX1 I_13(I1470,,,I15928,);
endmodule


