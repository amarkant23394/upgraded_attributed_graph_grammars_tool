module test_I1424(I1263,I1215,I1424);
input I1263,I1215;
output I1424;
wire I1359;
not I_0(I1359,I1263);
nor I_1(I1424,I1359,I1215);
endmodule


