module test_I4674(I1477,I1470,I1239,I4674);
input I1477,I1470,I1239;
output I4674;
wire I2181,I4544,I2155,I2633;
not I_0(I2181,I1477);
not I_1(I4544,I1477);
DFFARX1 I_2(I2155,I1470,I4544,,,I4674,);
DFFARX1 I_3(I2633,I1470,I2181,,,I2155,);
DFFARX1 I_4(I1239,I1470,I2181,,,I2633,);
endmodule


