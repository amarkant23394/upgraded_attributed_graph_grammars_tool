module test_I2146(I1343,I1231,I1477,I1470,I1375,I1271,I2146);
input I1343,I1231,I1477,I1470,I1375,I1271;
output I2146;
wire I2181,I2232,I2198,I2345,I2393,I2215;
and I_0(I2146,I2232,I2393);
not I_1(I2181,I1477);
DFFARX1 I_2(I2215,I1470,I2181,,,I2232,);
nand I_3(I2198,I1343,I1231);
DFFARX1 I_4(I1375,I1470,I2181,,,I2345,);
DFFARX1 I_5(I2345,I1470,I2181,,,I2393,);
and I_6(I2215,I2198,I1271);
endmodule


