module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_7_r_12,blif_reset_net_7_r_12,N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_7_r_12,blif_reset_net_7_r_12;
output N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,n_573_7_r_12,n_452_7_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n8_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_7_r_12,n8_12,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
nor I_36(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_37(N1508_0_r_12,n30_12,n37_12);
nor I_38(N1507_6_r_12,n25_12,n39_12);
nor I_39(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_40(n1_12,blif_clk_net_7_r_12,n8_12,G42_7_r_12,);
nor I_41(n_572_7_r_12,n23_12,n24_12);
nand I_42(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_43(n_549_7_r_12,n27_12,n28_12);
nand I_44(n_569_7_r_12,n25_12,n26_12);
nand I_45(n_452_7_r_12,n_573_7_r_3,N1507_6_r_3);
nand I_46(N6147_9_r_12,n30_12,n31_12);
nor I_47(N6134_9_r_12,n35_12,n36_12);
not I_48(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_49(n1_12,n_573_7_r_12);
not I_50(n8_12,blif_reset_net_7_r_12);
not I_51(n23_12,n36_12);
nor I_52(n24_12,n_452_7_r_12,G42_7_r_3);
nand I_53(n25_12,n23_12,n40_12);
not I_54(n26_12,n35_12);
not I_55(n27_12,N6134_9_r_12);
nand I_56(n28_12,n26_12,n29_12);
not I_57(n29_12,n24_12);
nand I_58(n30_12,n33_12,n41_12);
nand I_59(n31_12,n32_12,n33_12);
nor I_60(n32_12,n26_12,n34_12);
nor I_61(n33_12,n_549_7_r_3,N1372_1_r_3);
nor I_62(n34_12,n42_12,N1508_6_r_3);
nor I_63(n35_12,n38_12,N1508_1_r_3);
nand I_64(n36_12,N1507_6_r_3,G42_7_r_3);
nand I_65(n37_12,n23_12,n35_12);
or I_66(n38_12,n_452_7_r_3,N1508_6_r_3);
not I_67(n39_12,n30_12);
or I_68(n40_12,N1372_1_r_3,N6134_9_r_3);
nor I_69(n41_12,n34_12,n36_12);
nor I_70(n42_12,n_569_7_r_3,N1508_1_r_3);
endmodule


