module test_I6907_rst(I1477_rst,I6907_rst);
,I6907_rst);
input I1477_rst;
output I6907_rst;
wire ;
not I_0(I6907_rst,I1477_rst);
endmodule


