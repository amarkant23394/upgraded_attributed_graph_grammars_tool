module test_final(G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_17,blif_reset_net_1_r_17,G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17);
input G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_17,blif_reset_net_1_r_17;
output G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17;
wire G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,n_452_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15,n4_1_l_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15,n_431_0_l_17,n6_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17;
DFFARX1 I_0(n_452_1_r_15,blif_clk_net_1_r_17,n6_17,G42_1_r_15,);
and I_1(n_572_1_r_15,n17_15,n19_15);
nand I_2(n_573_1_r_15,n15_15,n18_15);
nor I_3(n_549_1_r_15,n21_15,n22_15);
nand I_4(n_569_1_r_15,n15_15,n20_15);
nor I_5(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_6(G42_1_l_15,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_15,);
nor I_7(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_8(N1_4_r_15,blif_clk_net_1_r_17,n6_17,G199_4_r_15,);
DFFARX1 I_9(n_573_1_l_15,blif_clk_net_1_r_17,n6_17,G214_4_r_15,);
nor I_10(n4_1_l_15,G18_1_l_15,IN_1_1_l_15);
DFFARX1 I_11(n4_1_l_15,blif_clk_net_1_r_17,n6_17,G42_1_l_15,);
not I_12(n15_15,G42_1_l_15);
DFFARX1 I_13(IN_1_3_l_15,blif_clk_net_1_r_17,n6_17,n17_internal_15,);
not I_14(n17_15,n17_internal_15);
DFFARX1 I_15(IN_2_3_l_15,blif_clk_net_1_r_17,n6_17,n30_15,);
nor I_16(n_572_1_l_15,G15_1_l_15,IN_7_1_l_15);
DFFARX1 I_17(n_572_1_l_15,blif_clk_net_1_r_17,n6_17,n14_internal_15,);
not I_18(n14_15,n14_internal_15);
nand I_19(N1_4_r_15,n25_15,n26_15);
or I_20(n_573_1_l_15,IN_5_1_l_15,IN_9_1_l_15);
nor I_21(n18_15,IN_9_1_l_15,IN_10_1_l_15);
nand I_22(n19_15,n27_15,n28_15);
nand I_23(n20_15,IN_4_3_l_15,n30_15);
not I_24(n21_15,n20_15);
and I_25(n22_15,n17_15,n_572_1_l_15);
nor I_26(n23_15,G18_1_l_15,IN_5_1_l_15);
or I_27(n24_15,IN_9_1_l_15,IN_10_1_l_15);
or I_28(n25_15,G18_1_l_15,n_573_1_l_15);
nand I_29(n26_15,n19_15,n23_15);
not I_30(n27_15,IN_10_1_l_15);
nand I_31(n28_15,IN_4_1_l_15,n29_15);
not I_32(n29_15,G15_1_l_15);
DFFARX1 I_33(n4_1_r_17,blif_clk_net_1_r_17,n6_17,G42_1_r_17,);
nor I_34(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_35(n_573_1_r_17,n20_17,n21_17);
nand I_36(n_549_1_r_17,n23_17,n24_17);
nand I_37(n_569_1_r_17,n21_17,n22_17);
not I_38(n_452_1_r_17,n23_17);
DFFARX1 I_39(n19_17,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_17,);
nor I_40(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_41(N1_4_r_17,blif_clk_net_1_r_17,n6_17,G199_4_r_17,);
DFFARX1 I_42(n5_17,blif_clk_net_1_r_17,n6_17,G214_4_r_17,);
or I_43(n_431_0_l_17,n26_17,G199_4_r_15);
not I_44(n6_17,blif_reset_net_1_r_17);
DFFARX1 I_45(n_431_0_l_17,blif_clk_net_1_r_17,n6_17,n20_internal_17,);
not I_46(n20_17,n20_internal_17);
DFFARX1 I_47(n_266_and_0_3_r_15,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_17,);
DFFARX1 I_48(n_549_1_r_15,blif_clk_net_1_r_17,n6_17,n19_internal_17,);
not I_49(n19_17,n19_internal_17);
nor I_50(n4_1_r_17,n5_17,n25_17);
not I_51(n2_17,n29_17);
DFFARX1 I_52(n2_17,blif_clk_net_1_r_17,n6_17,n17_internal_17,);
not I_53(n17_17,n17_internal_17);
nor I_54(N1_4_r_17,n29_17,n31_17);
not I_55(n5_17,G42_1_r_15);
and I_56(n21_17,n32_17,n_572_1_r_15);
not I_57(n22_17,n25_17);
nand I_58(n23_17,n20_17,n22_17);
nand I_59(n24_17,n19_17,n22_17);
nand I_60(n25_17,n30_17,G214_4_r_15);
and I_61(n26_17,n27_17,n_569_1_r_15);
nor I_62(n27_17,n28_17,n_572_1_r_15);
not I_63(n28_17,G42_1_r_15);
nor I_64(n29_17,n28_17,n_573_1_r_15);
and I_65(n30_17,n5_17,n_573_1_r_15);
nor I_66(n31_17,n21_17,G42_1_r_15);
nor I_67(n32_17,G42_1_r_15,ACVQN2_3_r_15);
endmodule


