module test_final(G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_10,blif_reset_net_1_r_10,G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10);
input G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_10,blif_reset_net_1_r_10;
output G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10;
wire G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_452_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14,n4_1_l_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14,n_452_1_r_10,N3_2_l_10,n4_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10;
DFFARX1 I_0(n_452_1_r_14,blif_clk_net_1_r_10,n4_10,G42_1_r_14,);
and I_1(n_572_1_r_14,n18_14,n19_14);
nand I_2(n_573_1_r_14,n16_14,n17_14);
nor I_3(n_549_1_r_14,n20_14,n21_14);
or I_4(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_5(n_452_1_r_14,IN_10_1_l_14,n23_14);
nor I_6(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_7(N3_2_r_14,blif_clk_net_1_r_10,n4_10,G199_2_r_14,);
DFFARX1 I_8(n_572_1_l_14,blif_clk_net_1_r_10,n4_10,ACVQN1_5_r_14,);
not I_9(P6_5_r_14,P6_5_r_internal_14);
nor I_10(n4_1_l_14,G18_1_l_14,IN_1_1_l_14);
DFFARX1 I_11(n4_1_l_14,blif_clk_net_1_r_10,n4_10,n15_internal_14,);
not I_12(n15_14,n15_internal_14);
DFFARX1 I_13(IN_1_3_l_14,blif_clk_net_1_r_10,n4_10,ACVQN2_3_l_14,);
DFFARX1 I_14(IN_2_3_l_14,blif_clk_net_1_r_10,n4_10,ACVQN1_3_l_14,);
and I_15(N3_2_r_14,n26_14,n27_14);
nor I_16(n_572_1_l_14,G15_1_l_14,IN_7_1_l_14);
DFFARX1 I_17(ACVQN2_3_l_14,blif_clk_net_1_r_10,n4_10,P6_5_r_internal_14,);
nor I_18(n16_14,IN_9_1_l_14,IN_10_1_l_14);
not I_19(n17_14,n_572_1_l_14);
nor I_20(n18_14,IN_5_1_l_14,IN_9_1_l_14);
nand I_21(n19_14,IN_4_3_l_14,ACVQN1_3_l_14);
nor I_22(n20_14,G18_1_l_14,IN_5_1_l_14);
nor I_23(n21_14,n15_14,n22_14);
nand I_24(n22_14,n24_14,n25_14);
nand I_25(n23_14,n15_14,n24_14);
not I_26(n24_14,IN_9_1_l_14);
not I_27(n25_14,IN_5_1_l_14);
nor I_28(n26_14,IN_10_1_l_14,n20_14);
nand I_29(n27_14,IN_4_1_l_14,n28_14);
not I_30(n28_14,G15_1_l_14);
DFFARX1 I_31(n4_1_r_10,blif_clk_net_1_r_10,n4_10,G42_1_r_10,);
nor I_32(n_572_1_r_10,n26_10,n3_10);
nand I_33(n_573_1_r_10,n16_10,n18_10);
nand I_34(n_549_1_r_10,n19_10,n20_10);
nor I_35(n_452_1_r_10,n25_10,n21_10);
nor I_36(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_37(N3_2_r_10,blif_clk_net_1_r_10,n4_10,G199_2_r_10,);
DFFARX1 I_38(G199_4_l_10,blif_clk_net_1_r_10,n4_10,ACVQN2_3_r_10,);
nor I_39(n_266_and_0_3_r_10,n17_10,n13_10);
and I_40(N3_2_l_10,n23_10,P6_5_r_14);
not I_41(n4_10,blif_reset_net_1_r_10);
DFFARX1 I_42(N3_2_l_10,blif_clk_net_1_r_10,n4_10,n25_10,);
not I_43(n16_10,n25_10);
DFFARX1 I_44(ACVQN1_5_r_14,blif_clk_net_1_r_10,n4_10,n26_10,);
DFFARX1 I_45(n_42_2_r_14,blif_clk_net_1_r_10,n4_10,ACVQN1_3_l_10,);
and I_46(N1_4_l_10,n24_10,n_549_1_r_14);
DFFARX1 I_47(N1_4_l_10,blif_clk_net_1_r_10,n4_10,G199_4_l_10,);
DFFARX1 I_48(n_569_1_r_14,blif_clk_net_1_r_10,n4_10,n27_10,);
not I_49(n17_10,n27_10);
nor I_50(n4_1_r_10,n27_10,n21_10);
nor I_51(N3_2_r_10,n16_10,n22_10);
not I_52(n3_10,n18_10);
DFFARX1 I_53(n3_10,blif_clk_net_1_r_10,n4_10,n13_internal_10,);
not I_54(n13_10,n13_internal_10);
nand I_55(n18_10,ACVQN1_3_l_10,n_572_1_r_14);
not I_56(n19_10,n_452_1_r_10);
nand I_57(n20_10,n16_10,n26_10);
nor I_58(n21_10,n_573_1_r_14,n_572_1_r_14);
and I_59(n22_10,n26_10,n21_10);
nand I_60(n23_10,G42_1_r_14,n_573_1_r_14);
nand I_61(n24_10,G199_2_r_14,G42_1_r_14);
endmodule


