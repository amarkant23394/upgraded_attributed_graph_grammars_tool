module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_7_r_3,blif_reset_net_7_r_3,N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_7_r_3,blif_reset_net_7_r_3;
output N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,n_572_7_r_3,N6147_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n10_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_7_r_3,n10_3,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
not I_35(N1372_1_r_3,n40_3);
nor I_36(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_37(N1507_6_r_3,n31_3,n42_3);
nor I_38(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_39(n4_7_r_3,blif_clk_net_7_r_3,n10_3,G42_7_r_3,);
nor I_40(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_41(n_573_7_r_3,n30_3,n31_3);
nor I_42(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_43(n_569_7_r_3,n30_3,n32_3);
nor I_44(n_452_7_r_3,n35_3,G42_7_r_4);
not I_45(N6147_9_r_3,n32_3);
nor I_46(N6134_9_r_3,n36_3,n37_3);
not I_47(I_BUFF_1_9_r_3,n45_3);
nor I_48(n4_7_r_3,I_BUFF_1_9_r_3,G42_7_r_4);
not I_49(n10_3,blif_reset_net_7_r_3);
not I_50(n30_3,n39_3);
not I_51(n31_3,n35_3);
nand I_52(n32_3,n41_3,n_549_7_r_4);
nor I_53(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_54(n34_3,n46_3,G42_7_r_4);
nor I_55(n35_3,n43_3,n44_3);
not I_56(n36_3,n34_3);
nor I_57(n37_3,N6147_9_r_3,G42_7_r_4);
or I_58(n38_3,n_572_7_r_3,n34_3);
nor I_59(n39_3,n44_3,N6134_9_r_4);
nand I_60(n40_3,n39_3,G42_7_r_4);
nand I_61(n41_3,n_549_7_r_4,N1508_6_r_4);
nor I_62(n42_3,n34_3,n45_3);
not I_63(n43_3,n_572_7_r_4);
nor I_64(n44_3,N1371_0_r_4,n_572_7_r_4);
nand I_65(n45_3,n49_3,n50_3);
and I_66(n46_3,n47_3,N1507_6_r_4);
nand I_67(n47_3,n41_3,n48_3);
not I_68(n48_3,n_549_7_r_4);
nor I_69(n49_3,N1508_6_r_4,n_452_7_r_4);
or I_70(n50_3,n51_3,N1507_6_r_4);
nor I_71(n51_3,n_569_7_r_4,N1371_0_r_4);
endmodule


