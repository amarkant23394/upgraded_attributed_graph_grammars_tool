module test_I7570(I1477,I7570);
input I1477;
output I7570;
wire ;
not I_0(I7570,I1477);
endmodule


