module test_I16211(I14667,I14856,I1477,I1470,I16211);
input I14667,I14856,I1477,I1470;
output I16211;
wire I16356,I16240,I14356,I16373;
DFFARX1 I_0(I14356,I1470,I16240,,,I16356,);
not I_1(I16240,I1477);
not I_2(I16211,I16373);
nand I_3(I14356,I14667,I14856);
DFFARX1 I_4(I16356,I1470,I16240,,,I16373,);
endmodule


