module test_I8216_rst(I1477_rst,I8216_rst);
,I8216_rst);
input I1477_rst;
output I8216_rst;
wire ;
not I_0(I8216_rst,I1477_rst);
endmodule


