module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_7_r_4,blif_reset_net_7_r_4,N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_7_r_4,blif_reset_net_7_r_4;
output N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,N1508_0_r_4,n_573_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n6_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_7_r_4,n6_4,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_7_r_4,n6_4,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
nor I_35(N1371_0_r_4,n25_4,N1508_0_r_0);
not I_36(N1508_0_r_4,n25_4);
nor I_37(N1507_6_r_4,n32_4,n33_4);
nor I_38(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_39(n4_7_r_4,blif_clk_net_7_r_4,n6_4,G42_7_r_4,);
not I_40(n_572_7_r_4,n_573_7_r_4);
nand I_41(n_573_7_r_4,n21_4,n22_4);
nor I_42(n_549_7_r_4,n24_4,N1508_0_r_0);
nand I_43(n_569_7_r_4,n22_4,n23_4);
nor I_44(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_45(N6147_9_r_4,n28_4);
nor I_46(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_47(I_BUFF_1_9_r_4,n21_4);
nor I_48(n4_7_r_4,N6147_9_r_4,N1508_0_r_0);
not I_49(n6_4,blif_reset_net_7_r_4);
nand I_50(n21_4,n39_4,n40_4);
or I_51(n22_4,n31_4,n_569_7_r_0);
not I_52(n23_4,N1508_0_r_0);
nor I_53(n24_4,n25_4,n26_4);
nand I_54(n25_4,G42_7_r_0,n_429_or_0_5_r_0);
nand I_55(n26_4,n21_4,n27_4);
nand I_56(n27_4,n36_4,n37_4);
nand I_57(n28_4,n38_4,n_572_7_r_0);
nand I_58(n29_4,N1508_0_r_4,n30_4);
nand I_59(n30_4,n34_4,n35_4);
nor I_60(n31_4,N1508_0_r_0,n_549_7_r_0);
not I_61(n32_4,n30_4);
nor I_62(n33_4,n21_4,n28_4);
nand I_63(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_64(n35_4,N1508_0_r_4,n27_4);
not I_65(n36_4,n_573_7_r_0);
nand I_66(n37_4,n_576_5_r_0,n_547_5_r_0);
or I_67(n38_4,N1508_0_r_0,n_549_7_r_0);
nor I_68(n39_4,N1371_0_r_0,G78_5_r_0);
or I_69(n40_4,n41_4,n_429_or_0_5_r_0);
nor I_70(n41_4,G78_5_r_0,N1371_0_r_0);
endmodule


