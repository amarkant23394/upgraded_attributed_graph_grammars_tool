module test_I1393(I1231,I1294,I1301,I1287,I1239,I1393);
input I1231,I1294,I1301,I1287,I1239;
output I1393;
wire I1376,I1342,I1359;
and I_0(I1376,I1359,I1231);
not I_1(I1342,I1301);
nand I_2(I1359,I1287,I1239);
DFFARX1 I_3(I1376,I1294,I1342,,,I1393,);
endmodule


