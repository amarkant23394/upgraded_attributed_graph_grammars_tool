module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_7_r_2,blif_reset_net_7_r_2,N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_7_r_2,blif_reset_net_7_r_2;
output N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,n4_7_l_2,n10_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_7_r_2,n10_2,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
nor I_36(N1371_0_r_2,n32_2,n35_2);
nor I_37(N1508_0_r_2,n32_2,n55_2);
not I_38(N1372_1_r_2,n54_2);
nor I_39(N1508_1_r_2,n59_2,n54_2);
nor I_40(N6147_2_r_2,n42_2,n43_2);
nor I_41(N1507_6_r_2,n40_2,n53_2);
nor I_42(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_43(n4_7_r_2,blif_clk_net_7_r_2,n10_2,G42_7_r_2,);
nor I_44(n_572_7_r_2,n36_2,n37_2);
or I_45(n_573_7_r_2,n34_2,n35_2);
nor I_46(n_549_7_r_2,n40_2,n41_2);
nand I_47(n_569_7_r_2,n38_2,n39_2);
nor I_48(n_452_7_r_2,n59_2,n35_2);
nor I_49(n4_7_l_2,N1372_1_r_3,G42_7_r_3);
not I_50(n10_2,blif_reset_net_7_r_2);
DFFARX1 I_51(n4_7_l_2,blif_clk_net_7_r_2,n10_2,n59_2,);
not I_52(n33_2,n59_2);
and I_53(N3_8_l_2,n49_2,N1372_1_r_3);
DFFARX1 I_54(N3_8_l_2,blif_clk_net_7_r_2,n10_2,n32_internal_2,);
not I_55(n32_2,n32_internal_2);
nor I_56(n4_7_r_2,n59_2,n36_2);
not I_57(n34_2,n39_2);
nor I_58(n35_2,n_452_7_r_3,N1507_6_r_3);
nor I_59(n36_2,N1507_6_r_3,G42_7_r_3);
or I_60(n37_2,N1508_6_r_3,n_549_7_r_3);
not I_61(n38_2,n40_2);
nand I_62(n39_2,n45_2,n57_2);
nor I_63(n40_2,n47_2,N1508_1_r_3);
nor I_64(n41_2,n32_2,n36_2);
not I_65(n42_2,n53_2);
nand I_66(n43_2,n44_2,n45_2);
nand I_67(n44_2,n38_2,n46_2);
not I_68(n45_2,n_549_7_r_3);
nand I_69(n46_2,n47_2,n48_2);
nand I_70(n47_2,G42_7_r_3,N6134_9_r_3);
or I_71(n48_2,N1508_1_r_3,N1508_6_r_3);
nand I_72(n49_2,n_573_7_r_3,N1507_6_r_3);
nand I_73(n50_2,n51_2,n52_2);
not I_74(n51_2,n47_2);
nand I_75(n52_2,n38_2,n53_2);
nor I_76(n53_2,N1507_6_r_3,N1508_6_r_3);
nand I_77(n54_2,n42_2,n56_2);
nor I_78(n55_2,n34_2,n56_2);
nor I_79(n56_2,N1508_1_r_3,N1508_6_r_3);
nand I_80(n57_2,n58_2,n_569_7_r_3);
not I_81(n58_2,N1508_6_r_3);
endmodule


