module test_I17563(I15696,I16145,I15628,I13749,I17563);
input I15696,I16145,I15628,I13749;
output I17563;
wire I15597,I15832,I17532,I16162;
not I_0(I17563,I17532);
nor I_1(I15597,I15832,I16162);
nand I_2(I15832,I15628,I13749);
not I_3(I17532,I15597);
and I_4(I16162,I15696,I16145);
endmodule


