module test_I2344(I1239,I1207,I1294,I1577,I1301,I1223,I2344);
input I1239,I1207,I1294,I1577,I1301,I1223;
output I2344;
wire I2313,I1797,I1749,I1656,I1971,I1334,I1639,I1310,I1410,I1319,I1331,I1780,I1622,I1937,I1342,I1988;
DFFARX1 I_0(I1331,I1294,I1937,,,I2313,);
and I_1(I1797,I1780,I1656);
or I_2(I1749,I1639);
nand I_3(I1656,I1639);
nor I_4(I1971,I1310,I1319);
DFFARX1 I_5(I1797,I1294,I1342,,,I1334,);
and I_6(I1639,I1622,I1207);
DFFARX1 I_7(I1577,I1294,I1342,,,I1310,);
nor I_8(I1410,I1223,I1239);
DFFARX1 I_9(I1749,I1294,I1342,,,I1319,);
nor I_10(I2344,I2313,I1988);
nor I_11(I1331,I1639,I1410);
DFFARX1 I_12(I1294,I1342,,,I1780,);
DFFARX1 I_13(I1294,I1342,,,I1622,);
not I_14(I1937,I1301);
not I_15(I1342,I1301);
nand I_16(I1988,I1971,I1334);
endmodule


