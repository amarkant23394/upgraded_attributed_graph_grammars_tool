module test_I9462(I5737,I8527,I8216,I1470,I9462);
input I5737,I8527,I8216,I1470;
output I9462;
wire I9576,I8202,I8267,I8181,I8360,I8496,I8592,I5719,I8377,I8250,I8462;
not I_0(I9462,I9576);
nor I_1(I9576,I8181,I8202);
nand I_2(I8202,I8267,I8496);
nand I_3(I8267,I8250,I5737);
and I_4(I8181,I8360,I8592);
not I_5(I8360,I5719);
nor I_6(I8496,I8462,I8377);
DFFARX1 I_7(I8527,I1470,I8216,,,I8592,);
DFFARX1 I_8(I1470,,,I5719,);
not I_9(I8377,I8360);
nor I_10(I8250,I5719);
DFFARX1 I_11(I1470,I8216,,,I8462,);
endmodule


