module test_I3396(I1902,I1294,I1301,I3396);
input I1902,I1294,I1301;
output I3396;
wire I3379,I2548,I2583,I2945;
not I_0(I3396,I3379);
not I_1(I3379,I2548);
DFFARX1 I_2(I2945,I1294,I2583,,,I2548,);
not I_3(I2583,I1301);
DFFARX1 I_4(I1902,I1294,I2583,,,I2945,);
endmodule


