module test_I14353(I13231,I1477,I1470,I14353);
input I13231,I1477,I1470;
output I14353;
wire I13361,I13313,I13162,I13197,I14808,I13248,I14370;
DFFARX1 I_0(I13313,I1470,I13197,,,I13361,);
DFFARX1 I_1(I1470,I13197,,,I13313,);
and I_2(I13162,I13248,I13361);
not I_3(I13197,I1477);
not I_4(I14353,I14808);
DFFARX1 I_5(I13162,I1470,I14370,,,I14808,);
DFFARX1 I_6(I13231,I1470,I13197,,,I13248,);
not I_7(I14370,I1477);
endmodule


