module test_final(IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_3_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_4_4_l_2,IN_5_4_l_2,blif_clk_net_5_r_3,blif_reset_net_5_r_3,N1371_0_r_3,N1508_0_r_3,N6147_3_r_3,n_429_or_0_5_r_3,G78_5_r_3,n_576_5_r_3,n_102_5_r_3,n_547_5_r_3,N1508_10_r_3);
input IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_3_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_4_4_l_2,IN_5_4_l_2,blif_clk_net_5_r_3,blif_reset_net_5_r_3;
output N1371_0_r_3,N1508_0_r_3,N6147_3_r_3,n_429_or_0_5_r_3,G78_5_r_3,n_576_5_r_3,n_102_5_r_3,n_547_5_r_3,N1508_10_r_3;
wire N1371_0_r_2,N1508_0_r_2,N6147_3_r_2,n_429_or_0_5_r_2,G78_5_r_2,n_576_5_r_2,n_102_5_r_2,n_547_5_r_2,N1372_10_r_2,N1508_10_r_2,n_431_5_r_2,n21_2,n22_2,n23_2,n24_2,n25_2,n26_2,n27_2,n28_2,n29_2,n30_2,n31_2,n32_2,N1372_10_r_3,N3_8_l_3,n5_3,n39_3,n_431_5_r_3,n22_3,n23_3,n24_3,n25_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3;
nor I_0(N1371_0_r_2,n23_2,n24_2);
not I_1(N1508_0_r_2,n24_2);
nor I_2(N6147_3_r_2,n22_2,n26_2);
nand I_3(n_429_or_0_5_r_2,IN_3_1_l_2,n22_2);
DFFARX1 I_4(n_431_5_r_2,blif_clk_net_5_r_3,n5_3,G78_5_r_2,);
nand I_5(n_576_5_r_2,n21_2,n22_2);
not I_6(n_102_5_r_2,n23_2);
nand I_7(n_547_5_r_2,n22_2,n24_2);
not I_8(N1372_10_r_2,n29_2);
nor I_9(N1508_10_r_2,n28_2,n29_2);
nand I_10(n_431_5_r_2,n_102_5_r_2,n25_2);
nor I_11(n21_2,IN_3_1_l_2,n23_2);
and I_12(n22_2,IN_1_1_l_2,IN_2_1_l_2);
nor I_13(n23_2,n24_2,n31_2);
nand I_14(n24_2,IN_1_4_l_2,IN_2_4_l_2);
nand I_15(n25_2,n26_2,n27_2);
nor I_16(n26_2,IN_1_3_l_2,n30_2);
not I_17(n27_2,n_429_or_0_5_r_2);
nor I_18(n28_2,n22_2,n23_2);
nand I_19(n29_2,N1508_0_r_2,n26_2);
or I_20(n30_2,IN_2_3_l_2,IN_3_3_l_2);
nor I_21(n31_2,IN_5_4_l_2,n32_2);
and I_22(n32_2,IN_3_4_l_2,IN_4_4_l_2);
nor I_23(N1371_0_r_3,n39_3,n37_3);
nor I_24(N1508_0_r_3,n25_3,n37_3);
nor I_25(N6147_3_r_3,N1372_10_r_3,n33_3);
nand I_26(n_429_or_0_5_r_3,N1372_10_r_3,n30_3);
DFFARX1 I_27(n_431_5_r_3,blif_clk_net_5_r_3,n5_3,G78_5_r_3,);
nand I_28(n_576_5_r_3,n22_3,n23_3);
not I_29(n_102_5_r_3,n39_3);
nand I_30(n_547_5_r_3,n26_3,n27_3);
not I_31(N1372_10_r_3,n36_3);
nor I_32(N1508_10_r_3,n35_3,n36_3);
and I_33(N3_8_l_3,n34_3,N1371_0_r_2);
not I_34(n5_3,blif_reset_net_5_r_3);
DFFARX1 I_35(N3_8_l_3,blif_clk_net_5_r_3,n5_3,n39_3,);
nand I_36(n_431_5_r_3,n29_3,n30_3);
nor I_37(n22_3,n24_3,n25_3);
nor I_38(n23_3,n39_3,G78_5_r_2);
not I_39(n24_3,n27_3);
nand I_40(n25_3,N1371_0_r_2,n_547_5_r_2);
nor I_41(n26_3,n39_3,n28_3);
nor I_42(n27_3,N6147_3_r_2,N1508_10_r_2);
not I_43(n28_3,n37_3);
nand I_44(n29_3,N1372_10_r_3,n39_3);
nand I_45(n30_3,n31_3,n32_3);
not I_46(n31_3,n25_3);
not I_47(n32_3,G78_5_r_2);
nand I_48(n33_3,n24_3,n25_3);
nand I_49(n34_3,N6147_3_r_2,G78_5_r_2);
nor I_50(n35_3,n27_3,n31_3);
nand I_51(n36_3,n28_3,n38_3);
nand I_52(n37_3,n_576_5_r_2,n_547_5_r_2);
or I_53(n38_3,N1372_10_r_2,n_576_5_r_2);
endmodule


