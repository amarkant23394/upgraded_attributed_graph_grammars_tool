module test_I11412(I9413,I8879,I6881,I8830,I9049,I1470_clk,I1477_rst,I11412);
input I9413,I8879,I6881,I8830,I9049,I1470_clk,I1477_rst;
output I11412;
wire I11378,I8851,I11327,I9083,I9066,I8848,I11395,I8862_rst;
nor I_0(I11378,I11327,I8848);
or I_1(I8851,I9083,I9066);
not I_2(I11327,I8830);
nand I_3(I9083,I8879,I6881);
DFFARX1 I_4 (I9049,I1470_clk,I8862_rst,I9066);
nor I_5(I8848,I9083,I9413);
nand I_6(I11395,I11378,I8851);
not I_7(I8862_rst,I1477_rst);
not I_8(I11412,I11395);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule