module test_final(G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_17,blif_reset_net_1_r_17,G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17);
input G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_17,blif_reset_net_1_r_17;
output G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17;
wire G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4,n_431_0_l_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n_431_0_l_17,n6_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17;
DFFARX1 I_0(n4_1_r_4,blif_clk_net_1_r_17,n6_17,G42_1_r_4,);
nor I_1(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_2(n_573_1_r_4,G2_0_l_4,n16_4);
nor I_3(n_549_1_r_4,n22_4,n23_4);
nand I_4(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_5(n19_4,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_4,);
nor I_6(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_7(n19_4,blif_clk_net_1_r_17,n6_17,ACVQN1_5_r_4,);
not I_8(P6_5_r_4,P6_5_r_internal_4);
or I_9(n_431_0_l_4,IN_8_0_l_4,n26_4);
DFFARX1 I_10(n_431_0_l_4,blif_clk_net_1_r_17,n6_17,G78_0_l_4,);
DFFARX1 I_11(IN_2_5_l_4,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_4,);
not I_12(n16_4,ACVQN1_5_l_4);
DFFARX1 I_13(IN_1_5_l_4,blif_clk_net_1_r_17,n6_17,n17_internal_4,);
not I_14(n17_4,n17_internal_4);
nor I_15(n4_1_r_4,n30_4,n31_4);
nand I_16(n19_4,G1_0_l_4,n33_4);
DFFARX1 I_17(G78_0_l_4,blif_clk_net_1_r_17,n6_17,n15_internal_4,);
not I_18(n15_4,n15_internal_4);
DFFARX1 I_19(ACVQN1_5_l_4,blif_clk_net_1_r_17,n6_17,P6_5_r_internal_4,);
and I_20(n20_4,IN_11_0_l_4,n16_4);
nor I_21(n21_4,G2_0_l_4,IN_10_0_l_4);
nand I_22(n22_4,G78_0_l_4,n25_4);
nand I_23(n23_4,IN_11_0_l_4,n24_4);
not I_24(n24_4,G2_0_l_4);
not I_25(n25_4,IN_10_0_l_4);
and I_26(n26_4,IN_2_0_l_4,n27_4);
nor I_27(n27_4,IN_4_0_l_4,n28_4);
not I_28(n28_4,G1_0_l_4);
not I_29(n29_4,n30_4);
nand I_30(n30_4,IN_7_0_l_4,n32_4);
nand I_31(n31_4,IN_11_0_l_4,n25_4);
nor I_32(n32_4,G2_0_l_4,n33_4);
not I_33(n33_4,IN_5_0_l_4);
DFFARX1 I_34(n4_1_r_17,blif_clk_net_1_r_17,n6_17,G42_1_r_17,);
nor I_35(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_36(n_573_1_r_17,n20_17,n21_17);
nand I_37(n_549_1_r_17,n23_17,n24_17);
nand I_38(n_569_1_r_17,n21_17,n22_17);
not I_39(n_452_1_r_17,n23_17);
DFFARX1 I_40(n19_17,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_17,);
nor I_41(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_42(N1_4_r_17,blif_clk_net_1_r_17,n6_17,G199_4_r_17,);
DFFARX1 I_43(n5_17,blif_clk_net_1_r_17,n6_17,G214_4_r_17,);
or I_44(n_431_0_l_17,n26_17,G42_1_r_4);
not I_45(n6_17,blif_reset_net_1_r_17);
DFFARX1 I_46(n_431_0_l_17,blif_clk_net_1_r_17,n6_17,n20_internal_17,);
not I_47(n20_17,n20_internal_17);
DFFARX1 I_48(ACVQN1_5_r_4,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_17,);
DFFARX1 I_49(n_572_1_r_4,blif_clk_net_1_r_17,n6_17,n19_internal_17,);
not I_50(n19_17,n19_internal_17);
nor I_51(n4_1_r_17,n5_17,n25_17);
not I_52(n2_17,n29_17);
DFFARX1 I_53(n2_17,blif_clk_net_1_r_17,n6_17,n17_internal_17,);
not I_54(n17_17,n17_internal_17);
nor I_55(N1_4_r_17,n29_17,n31_17);
not I_56(n5_17,n_549_1_r_4);
and I_57(n21_17,n32_17,n_569_1_r_4);
not I_58(n22_17,n25_17);
nand I_59(n23_17,n20_17,n22_17);
nand I_60(n24_17,n19_17,n22_17);
nand I_61(n25_17,n30_17,n_572_1_r_4);
and I_62(n26_17,n27_17,n_266_and_0_3_r_4);
nor I_63(n27_17,n28_17,n_573_1_r_4);
not I_64(n28_17,ACVQN2_3_r_4);
nor I_65(n29_17,n28_17,P6_5_r_4);
and I_66(n30_17,n5_17,P6_5_r_4);
nor I_67(n31_17,n21_17,n_549_1_r_4);
nor I_68(n32_17,G42_1_r_4,n_549_1_r_4);
endmodule


