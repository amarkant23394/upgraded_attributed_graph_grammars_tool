module test_I14341(I1477,I1470,I13508,I13460,I14341);
input I1477,I1470,I13508,I13460;
output I14341;
wire I13177,I13542,I14455,I11302,I11278,I13296,I14370;
nand I_0(I13177,I13296,I13542);
DFFARX1 I_1(I14455,I1470,I14370,,,I14341,);
nor I_2(I13542,I13508,I13460);
DFFARX1 I_3(I13177,I1470,I14370,,,I14455,);
DFFARX1 I_4(I1470,,,I11302,);
DFFARX1 I_5(I1470,,,I11278,);
nor I_6(I13296,I11278,I11302);
not I_7(I14370,I1477);
endmodule


