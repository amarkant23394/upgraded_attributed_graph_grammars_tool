module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_5_r_11,blif_reset_net_5_r_11,N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_5_r_11,blif_reset_net_5_r_11;
output N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,n_102_5_r_11,N1372_10_r_11,n_431_5_r_11,n9_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_5_r_11,n9_11,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
not I_35(N1372_1_r_11,n53_11);
nor I_36(N1508_1_r_11,n39_11,n53_11);
nor I_37(N6147_2_r_11,n48_11,n49_11);
nor I_38(N6147_3_r_11,n44_11,n45_11);
nand I_39(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_40(n_431_5_r_11,blif_clk_net_5_r_11,n9_11,G78_5_r_11,);
nand I_41(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_42(n_102_5_r_11,n39_11);
nand I_43(n_547_5_r_11,n36_11,n37_11);
nor I_44(N1507_6_r_11,n52_11,n57_11);
nor I_45(N1508_6_r_11,n46_11,n51_11);
nor I_46(N1372_10_r_11,n43_11,n47_11);
nor I_47(N1508_10_r_11,n55_11,n56_11);
nand I_48(n_431_5_r_11,n40_11,n41_11);
not I_49(n9_11,blif_reset_net_5_r_11);
nor I_50(n36_11,n38_11,n39_11);
not I_51(n37_11,n40_11);
nor I_52(n38_11,n60_11,N1507_6_r_4);
nor I_53(n39_11,n54_11,N1508_6_r_4);
nand I_54(n40_11,N1507_6_r_4,n_452_7_r_4);
nand I_55(n41_11,n_102_5_r_11,n42_11);
and I_56(n42_11,n58_11,N1371_0_r_4);
not I_57(n43_11,n44_11);
nor I_58(n44_11,n40_11,n_549_7_r_4);
nand I_59(n45_11,n46_11,n47_11);
not I_60(n46_11,n38_11);
nand I_61(n47_11,n59_11,n62_11);
and I_62(n48_11,n37_11,n47_11);
or I_63(n49_11,n44_11,n50_11);
nor I_64(n50_11,n60_11,n61_11);
or I_65(n51_11,n_102_5_r_11,n52_11);
nor I_66(n52_11,n42_11,n57_11);
nand I_67(n53_11,n37_11,n50_11);
or I_68(n54_11,N1508_6_r_4,n_572_7_r_4);
nor I_69(n55_11,n38_11,n42_11);
not I_70(n56_11,N1372_10_r_11);
and I_71(n57_11,n38_11,n50_11);
and I_72(n58_11,n59_11,G42_7_r_4);
or I_73(n59_11,n63_11,n_549_7_r_4);
not I_74(n60_11,N6134_9_r_4);
nor I_75(n61_11,G42_7_r_4,N1371_0_r_4);
nand I_76(n62_11,n_572_7_r_4,n_569_7_r_4);
and I_77(n63_11,n_572_7_r_4,n_569_7_r_4);
endmodule


