module test_I11956(I7550,I1477,I7535,I1470,I11956);
input I7550,I1477,I7535,I1470;
output I11956;
wire I10349,I7538,I10041,I12349,I11973,I10120,I10332;
and I_0(I10349,I10332,I7550);
not I_1(I11956,I12349);
DFFARX1 I_2(I1470,,,I7538,);
nor I_3(I10041,I10349,I10120);
DFFARX1 I_4(I10041,I1470,I11973,,,I12349,);
not I_5(I11973,I1477);
nor I_6(I10120,I7538,I7535);
DFFARX1 I_7(I1470,,,I10332,);
endmodule


