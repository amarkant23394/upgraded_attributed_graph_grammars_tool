module test_I2878(I1351,I2878);
input I1351;
output I2878;
wire I2861;
not I_0(I2878,I2861);
not I_1(I2861,I1351);
endmodule


