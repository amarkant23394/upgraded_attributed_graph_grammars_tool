module test_final(IN_1_1_l,IN_2_1_l,IN_3_1_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,IN_1_6_l,IN_2_6_l,IN_3_6_l,IN_4_6_l,IN_5_6_l,IN_1_8_l,IN_2_8_l,IN_3_8_l,IN_6_8_l,blif_clk_net_5_r,blif_reset_net_5_r,N1371_0_r,N1508_0_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,G42_7_r,n_572_7_r,n_573_7_r,n_549_7_r,n_569_7_r,n_452_7_r);
input IN_1_1_l,IN_2_1_l,IN_3_1_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,IN_1_6_l,IN_2_6_l,IN_3_6_l,IN_4_6_l,IN_5_6_l,IN_1_8_l,IN_2_8_l,IN_3_8_l,IN_6_8_l,blif_clk_net_5_r,blif_reset_net_5_r;
output N1371_0_r,N1508_0_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,G42_7_r,n_572_7_r,n_573_7_r,n_549_7_r,n_569_7_r,n_452_7_r;
wire N1372_1_l,N1508_1_l,n4_1_l,N6147_3_l,n3_3_l,N6138_3_l,N1507_6_l,N1508_6_l,n6_6_l,n7_6_l,n8_6_l,n9_6_l,n_42_8_l,G199_8_l,N3_8_l,n3_8_l,n3_0_r,n4_0_r,n_431_5_r,n2_5_r,n11_5_r,n12_5_r,n13_5_r,n14_5_r,n15_5_r,n16_5_r,n_87_7_r,n4_7_r,n7_7_r;
not I_0(N1372_1_l,n4_1_l);
nor I_1(N1508_1_l,IN_3_1_l,n4_1_l);
nand I_2(n4_1_l,IN_1_1_l,IN_2_1_l);
nor I_3(N6147_3_l,IN_3_3_l,n3_3_l);
not I_4(n3_3_l,N6138_3_l);
nor I_5(N6138_3_l,IN_1_3_l,IN_2_3_l);
nor I_6(N1507_6_l,n8_6_l,n9_6_l);
and I_7(N1508_6_l,IN_2_6_l,n6_6_l);
nor I_8(n6_6_l,n7_6_l,n8_6_l);
not I_9(n7_6_l,IN_1_6_l);
nor I_10(n8_6_l,IN_5_6_l,n9_6_l);
and I_11(n9_6_l,IN_3_6_l,IN_4_6_l);
nor I_12(n_42_8_l,IN_1_8_l,IN_3_8_l);
DFFARX1 I_13(N3_8_l,blif_clk_net_5_r,n2_5_r,G199_8_l,);
and I_14(N3_8_l,IN_6_8_l,n3_8_l);
nand I_15(n3_8_l,IN_2_8_l,IN_3_8_l);
nor I_16(N1371_0_r,n4_0_r,N1507_6_l);
nor I_17(N1508_0_r,n3_0_r,n4_0_r);
nor I_18(n3_0_r,N6147_3_l,G199_8_l);
not I_19(n4_0_r,N1508_1_l);
nand I_20(n_429_or_0_5_r,n12_5_r,N1508_1_l);
DFFARX1 I_21(n_431_5_r,blif_clk_net_5_r,n2_5_r,G78_5_r,);
nand I_22(n_576_5_r,n11_5_r,N6147_3_l);
not I_23(n_102_5_r,N1372_1_l);
nand I_24(n_547_5_r,n13_5_r,N1507_6_l);
or I_25(n_431_5_r,n14_5_r,G199_8_l);
not I_26(n2_5_r,blif_reset_net_5_r);
nor I_27(n11_5_r,n12_5_r,N1372_1_l);
not I_28(n12_5_r,N1508_6_l);
nor I_29(n13_5_r,N1372_1_l,N6147_3_l);
and I_30(n14_5_r,n15_5_r,n_42_8_l);
nor I_31(n15_5_r,n16_5_r,G199_8_l);
not I_32(n16_5_r,N1508_1_l);
DFFARX1 I_33(n4_7_r,blif_clk_net_5_r,n2_5_r,G42_7_r,);
not I_34(n_87_7_r,N1508_6_l);
nor I_35(n_572_7_r,N1372_1_l,N1508_6_l);
or I_36(n_573_7_r,N1507_6_l,n_42_8_l);
nor I_37(n_549_7_r,n7_7_r,N1508_1_l);
or I_38(n_569_7_r,N1508_1_l,N1507_6_l);
nor I_39(n_452_7_r,N1508_6_l,n_42_8_l);
nor I_40(n4_7_r,N1508_6_l,n_42_8_l);
and I_41(n7_7_r,n_87_7_r,N1372_1_l);
endmodule


