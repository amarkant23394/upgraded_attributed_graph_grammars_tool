module test_I10961(I9491,I8216,I8753,I1470,I9525,I8205,I9672,I10961);
input I9491,I8216,I8753,I1470,I9525,I8205,I9672;
output I10961;
wire I8187,I9542,I9720,I10664,I9754,I9771,I9737,I9459,I8178,I9621,I9689,I9471;
DFFARX1 I_0(I1470,I8216,,,I8187,);
DFFARX1 I_1(I9525,I1470,I9491,,,I9542,);
nand I_2(I10961,I10664,I9459);
not I_3(I9720,I9689);
not I_4(I10664,I9471);
DFFARX1 I_5(I8187,I1470,I9491,,,I9754,);
and I_6(I9771,I9754,I8178);
nor I_7(I9737,I9621,I9720);
nand I_8(I9459,I9771,I9737);
DFFARX1 I_9(I8753,I1470,I8216,,,I8178,);
DFFARX1 I_10(I8205,I1470,I9491,,,I9621,);
DFFARX1 I_11(I9672,I1470,I9491,,,I9689,);
nor I_12(I9471,I9689,I9542);
endmodule


