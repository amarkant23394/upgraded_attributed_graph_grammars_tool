module test_I7139(I3470,I1477,I5156,I3380,I3353,I1470,I7139);
input I3470,I1477,I5156,I3380,I3353,I1470;
output I7139;
wire I7122,I5266,I7105,I5085,I5088,I5512,I5249,I3747,I5076,I5079,I5204,I5187,I7088,I5105,I3368;
and I_0(I7122,I7105,I5076);
not I_1(I5266,I5249);
nor I_2(I7105,I7088,I5079);
nand I_3(I5085,I5512,I5266);
DFFARX1 I_4(I1470,I5105,,,I5088,);
DFFARX1 I_5(I3368,I1470,I5105,,,I5512,);
not I_6(I5249,I3380);
DFFARX1 I_7(I1470,,,I3747,);
or I_8(I7139,I7122,I5085);
DFFARX1 I_9(I5204,I1470,I5105,,,I5076,);
DFFARX1 I_10(I5156,I1470,I5105,,,I5079,);
nand I_11(I5204,I5187,I3353);
nor I_12(I5187,I3380);
not I_13(I7088,I5088);
not I_14(I5105,I1477);
nand I_15(I3368,I3747,I3470);
endmodule


