module test_I10052(I1477,I10052);
input I1477;
output I10052;
wire ;
not I_0(I10052,I1477);
endmodule


