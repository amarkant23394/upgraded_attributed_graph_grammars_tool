module test_I10538(I7559,I1477,I7604,I7535,I7731,I1470,I6315,I10538);
input I7559,I1477,I7604,I7535,I7731,I1470,I6315;
output I10538;
wire I7556,I10086,I7621,I7816,I7570,I7850,I7544,I10490,I10052,I10103,I10069;
nand I_0(I7556,I7621,I7850);
and I_1(I10086,I10069,I7544);
nand I_2(I7621,I7604,I6315);
DFFARX1 I_3(I1470,I7570,,,I7816,);
not I_4(I7570,I1477);
nor I_5(I7850,I7816,I7731);
nor I_6(I10538,I10490,I10103);
DFFARX1 I_7(I7621,I1470,I7570,,,I7544,);
DFFARX1 I_8(I7556,I1470,I10052,,,I10490,);
not I_9(I10052,I1477);
DFFARX1 I_10(I10086,I1470,I10052,,,I10103,);
nand I_11(I10069,I7559,I7535);
endmodule


