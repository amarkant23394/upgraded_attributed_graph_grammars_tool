module test_I1560(I1231,I1223,I1294,I1239,I1492,I1301,I1560);
input I1231,I1223,I1294,I1239,I1492,I1301;
output I1560;
wire I1410,I1543,I1376,I1526,I1342,I1509,I1393,I1359;
nor I_0(I1410,I1223,I1239);
and I_1(I1560,I1410,I1543);
nor I_2(I1543,I1393,I1526);
and I_3(I1376,I1359,I1231);
not I_4(I1526,I1509);
not I_5(I1342,I1301);
DFFARX1 I_6(I1492,I1294,I1342,,,I1509,);
DFFARX1 I_7(I1376,I1294,I1342,,,I1393,);
nand I_8(I1359,I1239);
endmodule


