module test_I11302(I8830,I8851,I1477,I1470,I9258,I11302);
input I8830,I8851,I1477,I1470,I9258;
output I11302;
wire I11378,I8827,I11813,I11830,I11847,I11395,I8862,I11327,I11310,I11864,I11624;
nor I_0(I11378,I11327);
DFFARX1 I_1(I9258,I1470,I8862,,,I8827,);
DFFARX1 I_2(I1470,I11310,,,I11813,);
not I_3(I11830,I11813);
DFFARX1 I_4(I11864,I1470,I11310,,,I11302,);
nand I_5(I11847,I11830,I11395);
nand I_6(I11395,I11378,I8851);
not I_7(I8862,I1477);
not I_8(I11327,I8830);
not I_9(I11310,I1477);
and I_10(I11864,I11624,I11847);
nand I_11(I11624,I11327,I8827);
endmodule


