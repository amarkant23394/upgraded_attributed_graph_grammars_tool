module Benchmark_testing85000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2684,I2692,I2700,I2708,I2716,I2724,I2732,I2740,I2748,I2756,I2764,I2772,I2780,I2788,I2796,I2804,I2812,I2820,I2828,I2836,I2844,I2852,I2860,I2868,I2876,I2884,I2892,I2900,I2908,I2916,I2924,I2932,I2940,I2948,I2956,I2964,I2972,I2980,I2988,I2996,I3004,I3012,I3020,I3028,I3036,I3044,I3052,I3060,I3068,I3076,I3084,I3092,I3100,I3108,I3116,I3124,I3132,I3140,I3148,I3156,I3164,I3172,I3180,I3188,I3196,I3204,I3212,I3220,I3228,I3236,I3244,I3252,I3260,I3268,I3276,I3284,I3292,I3300,I3308,I3316,I3324,I3332,I3340,I3348,I3356,I3364,I3372,I3380,I3388,I3396,I3404,I3412,I3420,I3428,I3436,I3444,I3452,I3460,I3468,I3476,I3484,I3492,I3500,I3508,I3516,I3524,I3532,I3540,I3548,I3556,I3563,I3570,I40861,I40852,I40849,I40855,I40843,I40837,I40858,I40846,I40840,I70349,I70361,I70370,I70373,I70358,I70367,I70355,I70364,I70352,I82470,I82482,I82491,I82494,I82479,I82488,I82476,I82485,I82473,I136751,I136763,I136772,I136775,I136760,I136769,I136757,I136766,I136754,I203007,I202983,I202995,I202989,I203004,I202998,I202992,I202986,I203001,I342811,I342835,I342817,I342820,I342808,I342826,I342829,I342814,I342823,I342832,I362837,I362861,I362843,I362846,I362834,I362852,I362855,I362840,I362849,I362858,I399200,I399224,I399206,I399209,I399197,I399215,I399218,I399203,I399212,I399221,I425693,I425672,I425666,I425681,I425669,I425684,I425675,I425678,I425690,I425687,I432221,I432200,I432194,I432209,I432197,I432212,I432203,I432206,I432218,I432215,I529900,I529897,I529882,I529894,I529888,I529876,I529885,I529891,I529879,I530495,I530492,I530477,I530489,I530483,I530471,I530480,I530486,I530474,I538230,I538227,I538212,I538224,I538218,I538206,I538215,I538221,I538209,I748018,I748021,I748003,I748012,I748024,I748015,I748006,I748009,I748027,I752642,I752645,I752627,I752636,I752648,I752639,I752630,I752633,I752651,I861139,I861142,I861133,I861124,I861127,I861136,I861121,I861130,I865882,I865885,I865876,I865867,I865870,I865879,I865864,I865873,I896975,I896978,I896969,I896960,I896963,I896972,I896957,I896966,I898029,I898032,I898023,I898014,I898017,I898026,I898011,I898020,I955594,I955597,I955573,I955585,I955600,I955588,I955582,I955576,I955579,I955591,I965284,I965287,I965263,I965275,I965290,I965278,I965272,I965266,I965269,I965281,I1038282,I1038285,I1038261,I1038273,I1038288,I1038276,I1038270,I1038264,I1038267,I1038279,I1183490,I1183478,I1183499,I1183475,I1183496,I1183487,I1183493,I1183484,I1183481,I1251329,I1251308,I1251311,I1251326,I1251323,I1251320,I1251317,I1251305,I1251314,I1368421,I1368436,I1368418,I1368430,I1368445,I1368442,I1368439,I1368433,I1368427,I1368424);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2684,I2692,I2700,I2708,I2716,I2724,I2732,I2740,I2748,I2756,I2764,I2772,I2780,I2788,I2796,I2804,I2812,I2820,I2828,I2836,I2844,I2852,I2860,I2868,I2876,I2884,I2892,I2900,I2908,I2916,I2924,I2932,I2940,I2948,I2956,I2964,I2972,I2980,I2988,I2996,I3004,I3012,I3020,I3028,I3036,I3044,I3052,I3060,I3068,I3076,I3084,I3092,I3100,I3108,I3116,I3124,I3132,I3140,I3148,I3156,I3164,I3172,I3180,I3188,I3196,I3204,I3212,I3220,I3228,I3236,I3244,I3252,I3260,I3268,I3276,I3284,I3292,I3300,I3308,I3316,I3324,I3332,I3340,I3348,I3356,I3364,I3372,I3380,I3388,I3396,I3404,I3412,I3420,I3428,I3436,I3444,I3452,I3460,I3468,I3476,I3484,I3492,I3500,I3508,I3516,I3524,I3532,I3540,I3548,I3556,I3563,I3570;
output I40861,I40852,I40849,I40855,I40843,I40837,I40858,I40846,I40840,I70349,I70361,I70370,I70373,I70358,I70367,I70355,I70364,I70352,I82470,I82482,I82491,I82494,I82479,I82488,I82476,I82485,I82473,I136751,I136763,I136772,I136775,I136760,I136769,I136757,I136766,I136754,I203007,I202983,I202995,I202989,I203004,I202998,I202992,I202986,I203001,I342811,I342835,I342817,I342820,I342808,I342826,I342829,I342814,I342823,I342832,I362837,I362861,I362843,I362846,I362834,I362852,I362855,I362840,I362849,I362858,I399200,I399224,I399206,I399209,I399197,I399215,I399218,I399203,I399212,I399221,I425693,I425672,I425666,I425681,I425669,I425684,I425675,I425678,I425690,I425687,I432221,I432200,I432194,I432209,I432197,I432212,I432203,I432206,I432218,I432215,I529900,I529897,I529882,I529894,I529888,I529876,I529885,I529891,I529879,I530495,I530492,I530477,I530489,I530483,I530471,I530480,I530486,I530474,I538230,I538227,I538212,I538224,I538218,I538206,I538215,I538221,I538209,I748018,I748021,I748003,I748012,I748024,I748015,I748006,I748009,I748027,I752642,I752645,I752627,I752636,I752648,I752639,I752630,I752633,I752651,I861139,I861142,I861133,I861124,I861127,I861136,I861121,I861130,I865882,I865885,I865876,I865867,I865870,I865879,I865864,I865873,I896975,I896978,I896969,I896960,I896963,I896972,I896957,I896966,I898029,I898032,I898023,I898014,I898017,I898026,I898011,I898020,I955594,I955597,I955573,I955585,I955600,I955588,I955582,I955576,I955579,I955591,I965284,I965287,I965263,I965275,I965290,I965278,I965272,I965266,I965269,I965281,I1038282,I1038285,I1038261,I1038273,I1038288,I1038276,I1038270,I1038264,I1038267,I1038279,I1183490,I1183478,I1183499,I1183475,I1183496,I1183487,I1183493,I1183484,I1183481,I1251329,I1251308,I1251311,I1251326,I1251323,I1251320,I1251317,I1251305,I1251314,I1368421,I1368436,I1368418,I1368430,I1368445,I1368442,I1368439,I1368433,I1368427,I1368424;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2684,I2692,I2700,I2708,I2716,I2724,I2732,I2740,I2748,I2756,I2764,I2772,I2780,I2788,I2796,I2804,I2812,I2820,I2828,I2836,I2844,I2852,I2860,I2868,I2876,I2884,I2892,I2900,I2908,I2916,I2924,I2932,I2940,I2948,I2956,I2964,I2972,I2980,I2988,I2996,I3004,I3012,I3020,I3028,I3036,I3044,I3052,I3060,I3068,I3076,I3084,I3092,I3100,I3108,I3116,I3124,I3132,I3140,I3148,I3156,I3164,I3172,I3180,I3188,I3196,I3204,I3212,I3220,I3228,I3236,I3244,I3252,I3260,I3268,I3276,I3284,I3292,I3300,I3308,I3316,I3324,I3332,I3340,I3348,I3356,I3364,I3372,I3380,I3388,I3396,I3404,I3412,I3420,I3428,I3436,I3444,I3452,I3460,I3468,I3476,I3484,I3492,I3500,I3508,I3516,I3524,I3532,I3540,I3548,I3556,I3563,I3570,I3602,I1238388,I3628,I3636,I3653,I3594,I1238403,I3693,I3701,I3718,I1238400,I3735,I1238409,I3752,I3769,I3573,I3800,I3817,I3834,I1238397,I1238406,I3576,I3865,I3882,I1238394,I3899,I1238385,I3916,I3933,I3950,I3585,I3981,I1238391,I3998,I4015,I3591,I4046,I3588,I4077,I4103,I4111,I4128,I3582,I3579,I4197,I242851,I4223,I4231,I4248,I4189,I242857,I4288,I4296,I4313,I242866,I4330,I242860,I4347,I4364,I4168,I4395,I4412,I4429,I242863,I242869,I4171,I4460,I4477,I242872,I4494,I242848,I4511,I4528,I4545,I4180,I4576,I242854,I4593,I4610,I4186,I4641,I4183,I4672,I4698,I4706,I4723,I4177,I4174,I4792,I1234342,I4818,I4826,I4843,I4784,I1234357,I4883,I4891,I4908,I1234354,I4925,I1234363,I4942,I4959,I4763,I4990,I5007,I5024,I1234351,I1234360,I4766,I5055,I5072,I1234348,I5089,I1234339,I5106,I5123,I5140,I4775,I5171,I1234345,I5188,I5205,I4781,I5236,I4778,I5267,I5293,I5301,I5318,I4772,I4769,I5387,I1056763,I5413,I5421,I1056775,I5438,I5379,I1056760,I5478,I5486,I5503,I5520,I1056757,I5537,I5554,I5358,I5585,I5602,I5619,I1056766,I5361,I5650,I5667,I1056772,I5684,I5701,I5718,I5735,I5370,I5766,I1056769,I5783,I5800,I5376,I5831,I5373,I5862,I1056778,I5888,I5896,I5913,I5367,I5364,I5982,I368646,I6008,I6016,I368637,I6033,I5974,I368640,I6073,I6081,I6098,I368634,I6115,I368643,I6132,I6149,I5953,I6180,I6197,I6214,I368631,I368649,I5956,I6245,I6262,I6279,I368655,I6296,I6313,I6330,I5965,I6361,I368652,I6378,I6395,I5971,I6426,I5968,I6457,I368658,I6483,I6491,I6508,I5962,I5959,I6577,I332810,I6603,I6611,I332801,I6628,I6569,I332804,I6668,I6676,I6693,I332798,I6710,I332807,I6727,I6744,I6548,I6775,I6792,I6809,I332795,I332813,I6551,I6840,I6857,I6874,I332819,I6891,I6908,I6925,I6560,I6956,I332816,I6973,I6990,I6566,I7021,I6563,I7052,I332822,I7078,I7086,I7103,I6557,I6554,I7172,I1193882,I7198,I7206,I7223,I7164,I1193897,I7263,I7271,I7288,I1193894,I7305,I1193903,I7322,I7339,I7143,I7370,I7387,I7404,I1193891,I1193900,I7146,I7435,I7452,I1193888,I7469,I1193879,I7486,I7503,I7520,I7155,I7551,I1193885,I7568,I7585,I7161,I7616,I7158,I7647,I7673,I7681,I7698,I7152,I7149,I7767,I86171,I7793,I7801,I86162,I7818,I7759,I86183,I7858,I7866,I7883,I86159,I7900,I7917,I7934,I7738,I7965,I7982,I7999,I86168,I7741,I8030,I8047,I86180,I8064,I86177,I8081,I8098,I8115,I7750,I8146,I86174,I8163,I8180,I7756,I8211,I7753,I8242,I86165,I8268,I8276,I8293,I7747,I7744,I8362,I39798,I8388,I8396,I39792,I8413,I8354,I39807,I8453,I8461,I8478,I39801,I8495,I39783,I8512,I8529,I8333,I8560,I8577,I8594,I39789,I39795,I8336,I8625,I8642,I39786,I8659,I39804,I8676,I8693,I8710,I8345,I8741,I8758,I8775,I8351,I8806,I8348,I8837,I8863,I8871,I8888,I8342,I8339,I8957,I637030,I8983,I8991,I637048,I9008,I8949,I637042,I9048,I9056,I9073,I637033,I9090,I9107,I9124,I8928,I9155,I9172,I9189,I637039,I637027,I8931,I9220,I9237,I637045,I9254,I637051,I9271,I9288,I9305,I8940,I9336,I9353,I9370,I8946,I9401,I8943,I9432,I637036,I9458,I9466,I9483,I8937,I8934,I9552,I174426,I9578,I9586,I9603,I9544,I174432,I9643,I9651,I9668,I174441,I9685,I174435,I9702,I9719,I9523,I9750,I9767,I9784,I174438,I174444,I9526,I9815,I9832,I174447,I9849,I174423,I9866,I9883,I9900,I9535,I9931,I174429,I9948,I9965,I9541,I9996,I9538,I10027,I10053,I10061,I10078,I9532,I9529,I10147,I916834,I10173,I10181,I916825,I10198,I10139,I916828,I10238,I10246,I10263,I916840,I10280,I916819,I10297,I10314,I10118,I10345,I10362,I10379,I916831,I916837,I10121,I10410,I10427,I916822,I10444,I916813,I10461,I10478,I10495,I10130,I10526,I10543,I10560,I10136,I10591,I10133,I10622,I916816,I10648,I10656,I10673,I10127,I10124,I10742,I708145,I10768,I10776,I708124,I10793,I10734,I708133,I10833,I10841,I10858,I708139,I10875,I708136,I10892,I10909,I10713,I10940,I10957,I10974,I708127,I708121,I10716,I11005,I11022,I708142,I11039,I11056,I11073,I11090,I10725,I11121,I708130,I11138,I11155,I10731,I11186,I10728,I11217,I11243,I11251,I11268,I10722,I10719,I11337,I920710,I11363,I11371,I920701,I11388,I11329,I920704,I11428,I11436,I11453,I920716,I11470,I920695,I11487,I11504,I11308,I11535,I11552,I11569,I920707,I920713,I11311,I11600,I11617,I920698,I11634,I920689,I11651,I11668,I11685,I11320,I11716,I11733,I11750,I11326,I11781,I11323,I11812,I920692,I11838,I11846,I11863,I11317,I11314,I11932,I1226828,I11958,I11966,I11983,I11924,I1226843,I12023,I12031,I12048,I1226840,I12065,I1226849,I12082,I12099,I11903,I12130,I12147,I12164,I1226837,I1226846,I11906,I12195,I12212,I1226834,I12229,I1226825,I12246,I12263,I12280,I11915,I12311,I1226831,I12328,I12345,I11921,I12376,I11918,I12407,I12433,I12441,I12458,I11912,I11909,I12527,I1288912,I12553,I12561,I1288918,I12578,I12519,I1288921,I12618,I12626,I12643,I1288909,I12660,I1288927,I12677,I12694,I12498,I12725,I12742,I12759,I1288924,I1288933,I12501,I12790,I12807,I12824,I1288930,I12841,I12858,I12875,I12510,I12906,I1288915,I12923,I12940,I12516,I12971,I12513,I13002,I13028,I13036,I13053,I12507,I12504,I13122,I1195038,I13148,I13156,I13173,I13114,I1195053,I13213,I13221,I13238,I1195050,I13255,I1195059,I13272,I13289,I13093,I13320,I13337,I13354,I1195047,I1195056,I13096,I13385,I13402,I1195044,I13419,I1195035,I13436,I13453,I13470,I13105,I13501,I1195041,I13518,I13535,I13111,I13566,I13108,I13597,I13623,I13631,I13648,I13102,I13099,I13717,I426231,I13743,I13751,I426213,I13768,I13709,I426225,I13808,I13816,I13833,I426210,I13850,I426219,I13867,I13884,I13688,I13915,I13932,I13949,I426216,I426237,I13691,I13980,I13997,I426228,I14014,I426234,I14031,I14048,I14065,I13700,I14096,I14113,I14130,I13706,I14161,I13703,I14192,I426222,I14218,I14226,I14243,I13697,I13694,I14312,I540586,I14338,I14346,I540607,I14363,I14304,I540604,I14403,I14411,I14428,I14445,I540598,I14462,I14479,I14283,I14510,I14527,I14544,I540601,I540610,I14286,I14575,I14592,I540589,I14609,I540592,I14626,I14643,I14660,I14295,I14691,I14708,I14725,I14301,I14756,I14298,I14787,I540595,I14813,I14821,I14838,I14292,I14289,I14907,I1075837,I14933,I14941,I1075849,I14958,I14899,I1075834,I14998,I15006,I15023,I15040,I1075831,I15057,I15074,I14878,I15105,I15122,I15139,I1075840,I14881,I15170,I15187,I1075846,I15204,I15221,I15238,I15255,I14890,I15286,I1075843,I15303,I15320,I14896,I15351,I14893,I15382,I1075852,I15408,I15416,I15433,I14887,I14884,I15502,I1146486,I15528,I15536,I15553,I15494,I1146501,I15593,I15601,I15618,I1146498,I15635,I1146507,I15652,I15669,I15473,I15700,I15717,I15734,I1146495,I1146504,I15476,I15765,I15782,I1146492,I15799,I1146483,I15816,I15833,I15850,I15485,I15881,I1146489,I15898,I15915,I15491,I15946,I15488,I15977,I16003,I16011,I16028,I15482,I15479,I16100,I1161535,I16126,I16143,I16151,I16168,I1161523,I1161514,I16185,I1161511,I16211,I16092,I16083,I1161517,I16256,I16264,I1161529,I16281,I16080,I1161526,I16321,I16329,I16086,I16074,I16374,I1161520,I16391,I1161532,I16417,I16425,I16068,I16456,I16473,I16490,I16507,I16524,I16089,I16555,I16077,I16071,I16627,I1270345,I16653,I16670,I16678,I16695,I1270363,I1270357,I16712,I1270366,I16738,I16619,I16610,I1270351,I16783,I16791,I1270360,I16808,I16607,I1270348,I16848,I16856,I16613,I16601,I16901,I1270369,I1270354,I16918,I16944,I16952,I16595,I16983,I17000,I17017,I17034,I17051,I16616,I17082,I16604,I16598,I17154,I264274,I17180,I17197,I17205,I17222,I264292,I264277,I17239,I264280,I17265,I17146,I17137,I264268,I17310,I17318,I264271,I17335,I17134,I264283,I17375,I17383,I17140,I17128,I17428,I264289,I264286,I17445,I17471,I17479,I17122,I17510,I17527,I17544,I17561,I17578,I17143,I17609,I17131,I17125,I17681,I604674,I17707,I17724,I17732,I17749,I604659,I604677,I17766,I604671,I17792,I17673,I17664,I604668,I17837,I17845,I17862,I17661,I604662,I17902,I17910,I17667,I17655,I17955,I604683,I604665,I17972,I604680,I17998,I18006,I17649,I18037,I18054,I18071,I18088,I18105,I17670,I18136,I17658,I17652,I18208,I838469,I18234,I18251,I18259,I18276,I838460,I838481,I18293,I838463,I18319,I18200,I18191,I18364,I18372,I838478,I18389,I18188,I838472,I18429,I18437,I18194,I18182,I18482,I838466,I838475,I18499,I18525,I18533,I18176,I18564,I18581,I18598,I18615,I18632,I18197,I18663,I18185,I18179,I18735,I97229,I18761,I18778,I18786,I18803,I97244,I18820,I97247,I18846,I18727,I18718,I97241,I18891,I18899,I97250,I18916,I18715,I97226,I18956,I18964,I18721,I18709,I19009,I97232,I19026,I97235,I19052,I19060,I18703,I19091,I19108,I97238,I19125,I19142,I19159,I18724,I19190,I18712,I18706,I19262,I880629,I19288,I19305,I19313,I19330,I880620,I880641,I19347,I880623,I19373,I19254,I19245,I19418,I19426,I880638,I19443,I19242,I880632,I19483,I19491,I19248,I19236,I19536,I880626,I880635,I19553,I19579,I19587,I19230,I19618,I19635,I19652,I19669,I19686,I19251,I19717,I19239,I19233,I19789,I83000,I19815,I19832,I19840,I19857,I83015,I19874,I83018,I19900,I19781,I19772,I83012,I19945,I19953,I83021,I19970,I19769,I82997,I20010,I20018,I19775,I19763,I20063,I83003,I20080,I83006,I20106,I20114,I19757,I20145,I20162,I83009,I20179,I20196,I20213,I19778,I20244,I19766,I19760,I20316,I479522,I20342,I20359,I20367,I20384,I479525,I20401,I479546,I20427,I20308,I20299,I479534,I20472,I20480,I479537,I20497,I20296,I479543,I20537,I20545,I20302,I20290,I20590,I479540,I479528,I20607,I479531,I20633,I20641,I20284,I20672,I20689,I479549,I20706,I20723,I20740,I20305,I20771,I20293,I20287,I20843,I1330933,I20869,I20886,I20894,I20911,I1330936,I1330942,I20928,I1330951,I20954,I20835,I20826,I1330954,I20999,I21007,I1330945,I21024,I20823,I21064,I21072,I20829,I20817,I21117,I1330960,I1330939,I21134,I1330948,I21160,I21168,I20811,I21199,I21216,I1330957,I21233,I21250,I21267,I20832,I21298,I20820,I20814,I21370,I1200261,I21396,I21413,I21421,I21438,I1200249,I1200240,I21455,I1200237,I21481,I21362,I21353,I1200243,I21526,I21534,I1200255,I21551,I21350,I1200252,I21591,I21599,I21356,I21344,I21644,I1200246,I21661,I1200258,I21687,I21695,I21338,I21726,I21743,I21760,I21777,I21794,I21359,I21825,I21347,I21341,I21897,I870616,I21923,I21940,I21948,I21965,I870607,I870628,I21982,I870610,I22008,I21889,I21880,I22053,I22061,I870625,I22078,I21877,I870619,I22118,I22126,I21883,I21871,I22171,I870613,I870622,I22188,I22214,I22222,I21865,I22253,I22270,I22287,I22304,I22321,I21886,I22352,I21874,I21868,I22424,I750899,I22450,I22467,I22475,I22492,I750914,I750917,I22509,I750896,I22535,I22416,I22407,I750902,I22580,I22588,I750908,I22605,I22404,I22645,I22653,I22410,I22398,I22698,I750911,I750893,I22715,I750905,I22741,I22749,I22392,I22780,I22797,I22814,I22831,I22848,I22413,I22879,I22401,I22395,I22951,I650914,I22977,I22994,I23002,I23019,I650899,I650917,I23036,I650911,I23062,I22943,I22934,I650908,I23107,I23115,I23132,I22931,I650902,I23172,I23180,I22937,I22925,I23225,I650923,I650905,I23242,I650920,I23268,I23276,I22919,I23307,I23324,I23341,I23358,I23375,I22940,I23406,I22928,I22922,I23478,I431106,I23504,I23521,I23529,I23546,I431109,I23563,I431130,I23589,I23470,I23461,I431118,I23634,I23642,I431121,I23659,I23458,I431127,I23699,I23707,I23464,I23452,I23752,I431124,I431112,I23769,I431115,I23795,I23803,I23446,I23834,I23851,I431133,I23868,I23885,I23902,I23467,I23933,I23455,I23449,I24005,I248209,I24031,I24048,I24056,I24073,I248227,I248212,I24090,I248215,I24116,I23997,I23988,I248203,I24161,I24169,I248206,I24186,I23985,I248218,I24226,I24234,I23991,I23979,I24279,I248224,I248221,I24296,I24322,I24330,I23973,I24361,I24378,I24395,I24412,I24429,I23994,I24460,I23982,I23976,I24532,I516514,I24558,I24575,I24583,I24600,I516517,I24617,I516538,I24643,I24524,I24515,I516526,I24688,I24696,I516529,I24713,I24512,I516535,I24753,I24761,I24518,I24506,I24806,I516532,I516520,I24823,I516523,I24849,I24857,I24500,I24888,I24905,I516541,I24922,I24939,I24956,I24521,I24987,I24509,I24503,I25059,I1163847,I25085,I25102,I25110,I25127,I1163835,I1163826,I25144,I1163823,I25170,I25051,I25042,I1163829,I25215,I25223,I1163841,I25240,I25039,I1163838,I25280,I25288,I25045,I25033,I25333,I1163832,I25350,I1163844,I25376,I25384,I25027,I25415,I25432,I25449,I25466,I25483,I25048,I25514,I25036,I25030,I25586,I1320136,I25612,I25629,I25637,I25654,I1320139,I1320133,I25671,I1320142,I25697,I25578,I25569,I1320130,I25742,I25750,I1320145,I25767,I25566,I1320121,I25807,I25815,I25572,I25560,I25860,I1320124,I25877,I25903,I25911,I25554,I25942,I25959,I1320127,I25976,I25993,I26010,I25575,I26041,I25563,I25557,I26113,I138335,I26139,I26156,I26164,I26181,I138350,I26198,I138353,I26224,I26105,I26096,I138347,I26269,I26277,I138356,I26294,I26093,I138332,I26334,I26342,I26099,I26087,I26387,I138338,I26404,I138341,I26430,I26438,I26081,I26469,I26486,I138344,I26503,I26520,I26537,I26102,I26568,I26090,I26084,I26640,I627216,I26666,I26683,I26691,I26708,I627201,I627219,I26725,I627213,I26751,I26632,I26623,I627210,I26796,I26804,I26821,I26620,I627204,I26861,I26869,I26626,I26614,I26914,I627225,I627207,I26931,I627222,I26957,I26965,I26608,I26996,I27013,I27030,I27047,I27064,I26629,I27095,I26617,I26611,I27167,I745119,I27193,I27210,I27218,I27235,I745134,I745137,I27252,I745116,I27278,I27159,I27150,I745122,I27323,I27331,I745128,I27348,I27147,I27388,I27396,I27153,I27141,I27441,I745131,I745113,I27458,I745125,I27484,I27492,I27135,I27523,I27540,I27557,I27574,I27591,I27156,I27622,I27144,I27138,I27694,I58231,I27720,I27737,I27745,I27762,I58246,I27779,I58249,I27805,I27686,I27677,I58243,I27850,I27858,I58252,I27875,I27674,I58228,I27915,I27923,I27680,I27668,I27968,I58234,I27985,I58237,I28011,I28019,I27662,I28050,I28067,I58240,I28084,I28101,I28118,I27683,I28149,I27671,I27665,I28221,I1274153,I28247,I28264,I28272,I28289,I1274171,I1274165,I28306,I1274174,I28332,I28213,I28204,I1274159,I28377,I28385,I1274168,I28402,I28201,I1274156,I28442,I28450,I28207,I28195,I28495,I1274177,I1274162,I28512,I28538,I28546,I28189,I28577,I28594,I28611,I28628,I28645,I28210,I28676,I28198,I28192,I28748,I1165003,I28774,I28791,I28799,I28816,I1164991,I1164982,I28833,I1164979,I28859,I28740,I28731,I1164985,I28904,I28912,I1164997,I28929,I28728,I1164994,I28969,I28977,I28734,I28722,I29022,I1164988,I29039,I1165000,I29065,I29073,I28716,I29104,I29121,I29138,I29155,I29172,I28737,I29203,I28725,I28719,I29275,I903817,I29301,I29318,I29326,I29343,I903808,I903829,I29360,I903811,I29386,I29267,I29258,I29431,I29439,I903826,I29456,I29255,I903820,I29496,I29504,I29261,I29249,I29549,I903814,I903823,I29566,I29592,I29600,I29243,I29631,I29648,I29665,I29682,I29699,I29264,I29730,I29252,I29246,I29802,I302256,I29828,I29845,I29853,I29870,I302253,I302247,I29887,I302241,I29913,I29794,I29785,I302229,I29958,I29966,I302238,I29983,I29782,I302235,I30023,I30031,I29788,I29776,I30076,I302232,I302250,I30093,I30119,I30127,I29770,I30158,I30175,I302244,I30192,I30209,I30226,I29791,I30257,I29779,I29773,I30329,I523586,I30355,I30372,I30380,I30397,I523589,I30414,I523610,I30440,I30321,I30312,I523598,I30485,I30493,I523601,I30510,I30309,I523607,I30550,I30558,I30315,I30303,I30603,I523604,I523592,I30620,I523595,I30646,I30654,I30297,I30685,I30702,I523613,I30719,I30736,I30753,I30318,I30784,I30306,I30300,I30856,I104080,I30882,I30899,I30907,I30924,I104095,I30941,I104098,I30967,I30848,I30839,I104092,I31012,I31020,I104101,I31037,I30836,I104077,I31077,I31085,I30842,I30830,I31130,I104083,I31147,I104086,I31173,I31181,I30824,I31212,I31229,I104089,I31246,I31263,I31280,I30845,I31311,I30833,I30827,I31383,I380252,I31409,I31426,I31434,I31451,I380249,I380243,I31468,I380237,I31494,I31375,I31366,I380225,I31539,I31547,I380234,I31564,I31363,I380231,I31604,I31612,I31369,I31357,I31657,I380228,I380246,I31674,I31700,I31708,I31351,I31739,I31756,I380240,I31773,I31790,I31807,I31372,I31838,I31360,I31354,I31910,I877994,I31936,I31953,I31961,I31978,I877985,I878006,I31995,I877988,I32021,I31902,I31893,I32066,I32074,I878003,I32091,I31890,I877997,I32131,I32139,I31896,I31884,I32184,I877991,I878000,I32201,I32227,I32235,I31878,I32266,I32283,I32300,I32317,I32334,I31899,I32365,I31887,I31881,I32437,I280934,I32463,I32480,I32488,I32505,I280952,I280937,I32522,I280940,I32548,I32429,I32420,I280928,I32593,I32601,I280931,I32618,I32417,I280943,I32658,I32666,I32423,I32411,I32711,I280949,I280946,I32728,I32754,I32762,I32405,I32793,I32810,I32827,I32844,I32861,I32426,I32892,I32414,I32408,I32964,I255349,I32990,I33007,I33015,I33032,I255367,I255352,I33049,I255355,I33075,I32956,I32947,I255343,I33120,I33128,I255346,I33145,I32944,I255358,I33185,I33193,I32950,I32938,I33238,I255364,I255361,I33255,I33281,I33289,I32932,I33320,I33337,I33354,I33371,I33388,I32953,I33419,I32941,I32935,I33491,I942677,I33517,I33534,I33542,I33559,I942653,I942680,I33576,I942665,I33602,I33483,I33474,I942671,I33647,I33655,I942656,I33672,I33471,I942674,I33712,I33720,I33477,I33465,I33765,I942659,I942662,I33782,I33808,I33816,I33459,I33847,I33864,I942668,I33881,I33898,I33915,I33480,I33946,I33468,I33462,I34018,I1317824,I34044,I34061,I34069,I34086,I1317827,I1317821,I34103,I1317830,I34129,I34010,I34001,I1317818,I34174,I34182,I1317833,I34199,I33998,I1317809,I34239,I34247,I34004,I33992,I34292,I1317812,I34309,I34335,I34343,I33986,I34374,I34391,I1317815,I34408,I34425,I34442,I34007,I34473,I33995,I33989,I34545,I519778,I34571,I34588,I34596,I34613,I519781,I34630,I519802,I34656,I34537,I34528,I519790,I34701,I34709,I519793,I34726,I34525,I519799,I34766,I34774,I34531,I34519,I34819,I519796,I519784,I34836,I519787,I34862,I34870,I34513,I34901,I34918,I519805,I34935,I34952,I34969,I34534,I35000,I34522,I34516,I35072,I616812,I35098,I35115,I35123,I35140,I616797,I616815,I35157,I616809,I35183,I35064,I35055,I616806,I35228,I35236,I35253,I35052,I616800,I35293,I35301,I35058,I35046,I35346,I616821,I616803,I35363,I616818,I35389,I35397,I35040,I35428,I35445,I35462,I35479,I35496,I35061,I35527,I35049,I35043,I35599,I1097955,I35625,I35642,I35650,I35667,I1097943,I1097934,I35684,I1097931,I35710,I35591,I35582,I1097937,I35755,I35763,I1097949,I35780,I35579,I1097946,I35820,I35828,I35585,I35573,I35873,I1097940,I35890,I1097952,I35916,I35924,I35567,I35955,I35972,I35989,I36006,I36023,I35588,I36054,I35576,I35570,I36126,I1283945,I36152,I36169,I36177,I36194,I1283963,I1283957,I36211,I1283966,I36237,I36118,I36109,I1283951,I36282,I36290,I1283960,I36307,I36106,I1283948,I36347,I36355,I36112,I36100,I36400,I1283969,I1283954,I36417,I36443,I36451,I36094,I36482,I36499,I36516,I36533,I36550,I36115,I36581,I36103,I36097,I36653,I475714,I36679,I36696,I36704,I36721,I475717,I36738,I475738,I36764,I36645,I36636,I475726,I36809,I36817,I475729,I36834,I36633,I475735,I36874,I36882,I36639,I36627,I36927,I475732,I475720,I36944,I475723,I36970,I36978,I36621,I37009,I37026,I475741,I37043,I37060,I37077,I36642,I37108,I36630,I36624,I37180,I203584,I37206,I37223,I37231,I37248,I203602,I203587,I37265,I203590,I37291,I37172,I37163,I203578,I37336,I37344,I203581,I37361,I37160,I203593,I37401,I37409,I37166,I37154,I37454,I203599,I203596,I37471,I37497,I37505,I37148,I37536,I37553,I37570,I37587,I37604,I37169,I37635,I37157,I37151,I37707,I1351163,I37733,I37750,I37758,I37775,I1351166,I1351172,I37792,I1351181,I37818,I37699,I37690,I1351184,I37863,I37871,I1351175,I37888,I37687,I37928,I37936,I37693,I37681,I37981,I1351190,I1351169,I37998,I1351178,I38024,I38032,I37675,I38063,I38080,I1351187,I38097,I38114,I38131,I37696,I38162,I37684,I37678,I38234,I509986,I38260,I38277,I38285,I38302,I509989,I38319,I510010,I38345,I38226,I38217,I509998,I38390,I38398,I510001,I38415,I38214,I510007,I38455,I38463,I38220,I38208,I38508,I510004,I509992,I38525,I509995,I38551,I38559,I38202,I38590,I38607,I510013,I38624,I38641,I38658,I38223,I38689,I38211,I38205,I38761,I329133,I38787,I38804,I38812,I38829,I329130,I329124,I38846,I329118,I38872,I38753,I38744,I329106,I38917,I38925,I329115,I38942,I38741,I329112,I38982,I38990,I38747,I38735,I39035,I329109,I329127,I39052,I39078,I39086,I38729,I39117,I39134,I329121,I39151,I39168,I39185,I38750,I39216,I38738,I38732,I39288,I876940,I39314,I39331,I39339,I39356,I876931,I876952,I39373,I876934,I39399,I39280,I39271,I39444,I39452,I876949,I39469,I39268,I876943,I39509,I39517,I39274,I39262,I39562,I876937,I876946,I39579,I39605,I39613,I39256,I39644,I39661,I39678,I39695,I39712,I39277,I39743,I39265,I39259,I39815,I1084252,I39841,I39858,I39866,I39883,I1084246,I1084267,I39900,I39926,I1084249,I39971,I39979,I1084258,I39996,I40036,I40044,I40089,I1084264,I40106,I1084255,I40132,I40140,I40171,I40188,I1084261,I40205,I40222,I40239,I40270,I40342,I1162691,I40368,I40385,I40393,I40410,I1162679,I1162670,I40427,I1162667,I40453,I40334,I40325,I1162673,I40498,I40506,I1162685,I40523,I40322,I1162682,I40563,I40571,I40328,I40316,I40616,I1162676,I40633,I1162688,I40659,I40667,I40310,I40698,I40715,I40732,I40749,I40766,I40331,I40797,I40319,I40313,I40869,I1232051,I40895,I40912,I40920,I40937,I1232039,I1232030,I40954,I1232027,I40980,I1232033,I41025,I41033,I1232045,I41050,I1232042,I41090,I41098,I41143,I1232036,I41160,I1232048,I41186,I41194,I41225,I41242,I41259,I41276,I41293,I41324,I41396,I387630,I41422,I41439,I41447,I41464,I387627,I387621,I41481,I387615,I41507,I41388,I41379,I387603,I41552,I41560,I387612,I41577,I41376,I387609,I41617,I41625,I41382,I41370,I41670,I387606,I387624,I41687,I41713,I41721,I41364,I41752,I41769,I387618,I41786,I41803,I41820,I41385,I41851,I41373,I41367,I41923,I949783,I41949,I41966,I41974,I41991,I949759,I949786,I42008,I949771,I42034,I41915,I41906,I949777,I42079,I42087,I949762,I42104,I41903,I949780,I42144,I42152,I41909,I41897,I42197,I949765,I949768,I42214,I42240,I42248,I41891,I42279,I42296,I949774,I42313,I42330,I42347,I41912,I42378,I41900,I41894,I42450,I362334,I42476,I42493,I42501,I42518,I362331,I362325,I42535,I362319,I42561,I42442,I42433,I362307,I42606,I42614,I362316,I42631,I42430,I362313,I42671,I42679,I42436,I42424,I42724,I362310,I362328,I42741,I42767,I42775,I42418,I42806,I42823,I362322,I42840,I42857,I42874,I42439,I42905,I42427,I42421,I42977,I1117029,I43003,I43020,I43028,I43045,I1117017,I1117008,I43062,I1117005,I43088,I42969,I42960,I1117011,I43133,I43141,I1117023,I43158,I42957,I1117020,I43198,I43206,I42963,I42951,I43251,I1117014,I43268,I1117026,I43294,I43302,I42945,I43333,I43350,I43367,I43384,I43401,I42966,I43432,I42954,I42948,I43504,I1192747,I43530,I43547,I43555,I43572,I1192735,I1192726,I43589,I1192723,I43615,I43496,I43487,I1192729,I43660,I43668,I1192741,I43685,I43484,I1192738,I43725,I43733,I43490,I43478,I43778,I1192732,I43795,I1192744,I43821,I43829,I43472,I43860,I43877,I43894,I43911,I43928,I43493,I43959,I43481,I43475,I44031,I495842,I44057,I44074,I44082,I44099,I495845,I44116,I495866,I44142,I44023,I44014,I495854,I44187,I44195,I495857,I44212,I44011,I495863,I44252,I44260,I44017,I44005,I44305,I495860,I495848,I44322,I495851,I44348,I44356,I43999,I44387,I44404,I495869,I44421,I44438,I44455,I44020,I44486,I44008,I44002,I44558,I421858,I44584,I44601,I44609,I44626,I421861,I44643,I421882,I44669,I44550,I44541,I421870,I44714,I44722,I421873,I44739,I44538,I421879,I44779,I44787,I44544,I44532,I44832,I421876,I421864,I44849,I421867,I44875,I44883,I44526,I44914,I44931,I421885,I44948,I44965,I44982,I44547,I45013,I44535,I44529,I45085,I871143,I45111,I45128,I45136,I45153,I871134,I871155,I45170,I871137,I45196,I45077,I45068,I45241,I45249,I871152,I45266,I45065,I871146,I45306,I45314,I45071,I45059,I45359,I871140,I871149,I45376,I45402,I45410,I45053,I45441,I45458,I45475,I45492,I45509,I45074,I45540,I45062,I45056,I45612,I829510,I45638,I45655,I45663,I45680,I829501,I829522,I45697,I829504,I45723,I45604,I45595,I45768,I45776,I829519,I45793,I45592,I829513,I45833,I45841,I45598,I45586,I45886,I829507,I829516,I45903,I45929,I45937,I45580,I45968,I45985,I46002,I46019,I46036,I45601,I46067,I45589,I45583,I46139,I1111249,I46165,I46182,I46190,I46207,I1111237,I1111228,I46224,I1111225,I46250,I46131,I46122,I1111231,I46295,I46303,I1111243,I46320,I46119,I1111240,I46360,I46368,I46125,I46113,I46413,I1111234,I46430,I1111246,I46456,I46464,I46107,I46495,I46512,I46529,I46546,I46563,I46128,I46594,I46116,I46110,I46666,I594848,I46692,I46709,I46717,I46734,I594833,I594851,I46751,I594845,I46777,I46658,I46649,I594842,I46822,I46830,I46847,I46646,I594836,I46887,I46895,I46652,I46640,I46940,I594857,I594839,I46957,I594854,I46983,I46991,I46634,I47022,I47039,I47056,I47073,I47090,I46655,I47121,I46643,I46637,I47193,I901709,I47219,I47236,I47244,I47261,I901700,I901721,I47278,I901703,I47304,I47185,I47176,I47349,I47357,I901718,I47374,I47173,I901712,I47414,I47422,I47179,I47167,I47467,I901706,I901715,I47484,I47510,I47518,I47161,I47549,I47566,I47583,I47600,I47617,I47182,I47648,I47170,I47164,I47720,I962057,I47746,I47763,I47771,I47788,I962033,I962060,I47805,I962045,I47831,I47712,I47703,I962051,I47876,I47884,I962036,I47901,I47700,I962054,I47941,I47949,I47706,I47694,I47994,I962039,I962042,I48011,I48037,I48045,I47688,I48076,I48093,I962048,I48110,I48127,I48144,I47709,I48175,I47697,I47691,I48247,I1309732,I48273,I48290,I48298,I48315,I1309735,I1309729,I48332,I1309738,I48358,I48239,I48230,I1309726,I48403,I48411,I1309741,I48428,I48227,I1309717,I48468,I48476,I48233,I48221,I48521,I1309720,I48538,I48564,I48572,I48215,I48603,I48620,I1309723,I48637,I48654,I48671,I48236,I48702,I48224,I48218,I48774,I831618,I48800,I48817,I48825,I48842,I831609,I831630,I48859,I831612,I48885,I48766,I48757,I48930,I48938,I831627,I48955,I48754,I831621,I48995,I49003,I48760,I48748,I49048,I831615,I831624,I49065,I49091,I49099,I48742,I49130,I49147,I49164,I49181,I49198,I48763,I49229,I48751,I48745,I49301,I1249673,I49327,I49344,I49352,I49369,I1249691,I1249685,I49386,I1249694,I49412,I49293,I49284,I1249679,I49457,I49465,I1249688,I49482,I49281,I1249676,I49522,I49530,I49287,I49275,I49575,I1249697,I1249682,I49592,I49618,I49626,I49269,I49657,I49674,I49691,I49708,I49725,I49290,I49756,I49278,I49272,I49828,I1131479,I49854,I49871,I49879,I49896,I1131467,I1131458,I49913,I1131455,I49939,I49820,I49811,I1131461,I49984,I49992,I1131473,I50009,I49808,I1131470,I50049,I50057,I49814,I49802,I50102,I1131464,I50119,I1131476,I50145,I50153,I49796,I50184,I50201,I50218,I50235,I50252,I49817,I50283,I49805,I49799,I50355,I509442,I50381,I50398,I50406,I50423,I509445,I50440,I509466,I50466,I50347,I50338,I509454,I50511,I50519,I509457,I50536,I50335,I509463,I50576,I50584,I50341,I50329,I50629,I509460,I509448,I50646,I509451,I50672,I50680,I50323,I50711,I50728,I509469,I50745,I50762,I50779,I50344,I50810,I50332,I50326,I50882,I1388053,I50908,I50925,I50933,I50950,I1388056,I1388062,I50967,I1388071,I50993,I50874,I50865,I1388074,I51038,I51046,I1388065,I51063,I50862,I51103,I51111,I50868,I50856,I51156,I1388080,I1388059,I51173,I1388068,I51199,I51207,I50850,I51238,I51255,I1388077,I51272,I51289,I51306,I50871,I51337,I50859,I50853,I51409,I263679,I51435,I51452,I51460,I51477,I263697,I263682,I51494,I263685,I51520,I51401,I51392,I263673,I51565,I51573,I263676,I51590,I51389,I263688,I51630,I51638,I51395,I51383,I51683,I263694,I263691,I51700,I51726,I51734,I51377,I51765,I51782,I51799,I51816,I51833,I51398,I51864,I51386,I51380,I51936,I773441,I51962,I51979,I51987,I52004,I773456,I773459,I52021,I773438,I52047,I51928,I51919,I773444,I52092,I52100,I773450,I52117,I51916,I52157,I52165,I51922,I51910,I52210,I773453,I773435,I52227,I773447,I52253,I52261,I51904,I52292,I52309,I52326,I52343,I52360,I51925,I52391,I51913,I51907,I52463,I794249,I52489,I52506,I52514,I52531,I794264,I794267,I52548,I794246,I52574,I52455,I52446,I794252,I52619,I52627,I794258,I52644,I52443,I52684,I52692,I52449,I52437,I52737,I794261,I794243,I52754,I794255,I52780,I52788,I52431,I52819,I52836,I52853,I52870,I52887,I52452,I52918,I52440,I52434,I52990,I452322,I53016,I53033,I53041,I53058,I452325,I53075,I452346,I53101,I52982,I52973,I452334,I53146,I53154,I452337,I53171,I52970,I452343,I53211,I53219,I52976,I52964,I53264,I452340,I452328,I53281,I452331,I53307,I53315,I52958,I53346,I53363,I452349,I53380,I53397,I53414,I52979,I53445,I52967,I52961,I53517,I1281769,I53543,I53560,I53568,I53585,I1281787,I1281781,I53602,I1281790,I53628,I53509,I53500,I1281775,I53673,I53681,I1281784,I53698,I53497,I1281772,I53738,I53746,I53503,I53491,I53791,I1281793,I1281778,I53808,I53834,I53842,I53485,I53873,I53890,I53907,I53924,I53941,I53506,I53972,I53494,I53488,I54044,I876413,I54070,I54087,I54095,I54112,I876404,I876425,I54129,I876407,I54155,I54036,I54027,I54200,I54208,I876422,I54225,I54024,I876416,I54265,I54273,I54030,I54018,I54318,I876410,I876419,I54335,I54361,I54369,I54012,I54400,I54417,I54434,I54451,I54468,I54033,I54499,I54021,I54015,I54571,I836888,I54597,I54614,I54622,I54639,I836879,I836900,I54656,I836882,I54682,I54563,I54554,I54727,I54735,I836897,I54752,I54551,I836891,I54792,I54800,I54557,I54545,I54845,I836885,I836894,I54862,I54888,I54896,I54539,I54927,I54944,I54961,I54978,I54995,I54560,I55026,I54548,I54542,I55098,I296459,I55124,I55141,I55149,I55166,I296456,I296450,I55183,I296444,I55209,I55090,I55081,I296432,I55254,I55262,I296441,I55279,I55078,I296438,I55319,I55327,I55084,I55072,I55372,I296435,I296453,I55389,I55415,I55423,I55066,I55454,I55471,I296447,I55488,I55505,I55522,I55087,I55553,I55075,I55069,I55625,I634730,I55651,I55668,I55676,I55693,I634715,I634733,I55710,I634727,I55736,I55617,I55608,I634724,I55781,I55789,I55806,I55605,I634718,I55846,I55854,I55611,I55599,I55899,I634739,I634721,I55916,I634736,I55942,I55950,I55593,I55981,I55998,I56015,I56032,I56049,I55614,I56080,I55602,I55596,I56152,I733559,I56178,I56195,I56203,I56220,I733574,I733577,I56237,I733556,I56263,I56144,I56135,I733562,I56308,I56316,I733568,I56333,I56132,I56373,I56381,I56138,I56126,I56426,I733571,I733553,I56443,I733565,I56469,I56477,I56120,I56508,I56525,I56542,I56559,I56576,I56141,I56607,I56129,I56123,I56679,I1185811,I56705,I56722,I56730,I56747,I1185799,I1185790,I56764,I1185787,I56790,I56671,I56662,I1185793,I56835,I56843,I1185805,I56860,I56659,I1185802,I56900,I56908,I56665,I56653,I56953,I1185796,I56970,I1185808,I56996,I57004,I56647,I57035,I57052,I57069,I57086,I57103,I56668,I57134,I56656,I56650,I57206,I1212977,I57232,I57249,I57257,I57274,I1212965,I1212956,I57291,I1212953,I57317,I57198,I57189,I1212959,I57362,I57370,I1212971,I57387,I57186,I1212968,I57427,I57435,I57192,I57180,I57480,I1212962,I57497,I1212974,I57523,I57531,I57174,I57562,I57579,I57596,I57613,I57630,I57195,I57661,I57183,I57177,I57733,I1233207,I57759,I57776,I57784,I57801,I1233195,I1233186,I57818,I1233183,I57844,I57725,I57716,I1233189,I57889,I57897,I1233201,I57914,I57713,I1233198,I57954,I57962,I57719,I57707,I58007,I1233192,I58024,I1233204,I58050,I58058,I57701,I58089,I58106,I58123,I58140,I58157,I57722,I58188,I57710,I57704,I58260,I353902,I58286,I58294,I58311,I353884,I353899,I58328,I353875,I58354,I353878,I58371,I58379,I353893,I58396,I58427,I58444,I353896,I58484,I58506,I353887,I58523,I353881,I58549,I58566,I58588,I58619,I353890,I58636,I58653,I58670,I58701,I58787,I217870,I58813,I58821,I58838,I217864,I217858,I58855,I217879,I58881,I217876,I58898,I58906,I217873,I58923,I58755,I58954,I58971,I58767,I59011,I58776,I59033,I217861,I59050,I217882,I59076,I59093,I58779,I59115,I58764,I59146,I217867,I59163,I59180,I59197,I58773,I59228,I58761,I58770,I58758,I59314,I1380925,I59340,I59348,I59365,I1380919,I1380940,I59382,I1380916,I59408,I1380937,I59425,I59433,I1380934,I59450,I59282,I59481,I59498,I59294,I1380922,I59538,I59303,I59560,I1380931,I1380928,I59577,I1380913,I59603,I59620,I59306,I59642,I59291,I59673,I59690,I59707,I59724,I59300,I59755,I59288,I59297,I59285,I59841,I650330,I59867,I59875,I59892,I650342,I650327,I59909,I650321,I59935,I650336,I59952,I59960,I650324,I59977,I59809,I60008,I60025,I59821,I650333,I60065,I59830,I60087,I650339,I650345,I60104,I60130,I60147,I59833,I60169,I59818,I60200,I60217,I60234,I60251,I59827,I60282,I59815,I59824,I59812,I60368,I771135,I60394,I60402,I60419,I771126,I771144,I60436,I771123,I60462,I60479,I60487,I771129,I60504,I60336,I60535,I60552,I60348,I60592,I60357,I60614,I771141,I771132,I60631,I771147,I60657,I60674,I60360,I60696,I60345,I60727,I771138,I60744,I60761,I60778,I60354,I60809,I60342,I60351,I60339,I60895,I578080,I60921,I60929,I60946,I578092,I578077,I60963,I578071,I60989,I578086,I61006,I61014,I578074,I61031,I60863,I61062,I61079,I60875,I578083,I61119,I60884,I61141,I578089,I578095,I61158,I61184,I61201,I60887,I61223,I60872,I61254,I61271,I61288,I61305,I60881,I61336,I60869,I60878,I60866,I61422,I341781,I61448,I61456,I61473,I341763,I341778,I61490,I341754,I61516,I341757,I61533,I61541,I341772,I61558,I61390,I61589,I61606,I61402,I341775,I61646,I61411,I61668,I341766,I61685,I341760,I61711,I61728,I61414,I61750,I61399,I61781,I341769,I61798,I61815,I61832,I61408,I61863,I61396,I61405,I61393,I61949,I589062,I61975,I61983,I62000,I589074,I589059,I62017,I589053,I62043,I589068,I62060,I62068,I589056,I62085,I61917,I62116,I62133,I61929,I589065,I62173,I61938,I62195,I589071,I589077,I62212,I62238,I62255,I61941,I62277,I61926,I62308,I62325,I62342,I62359,I61935,I62390,I61923,I61932,I61920,I62476,I649752,I62502,I62510,I62527,I649764,I649749,I62544,I649743,I62570,I649758,I62587,I62595,I649746,I62612,I62444,I62643,I62660,I62456,I649755,I62700,I62465,I62722,I649761,I649767,I62739,I62765,I62782,I62468,I62804,I62453,I62835,I62852,I62869,I62886,I62462,I62917,I62450,I62459,I62447,I63003,I407129,I63029,I63037,I63054,I407111,I407126,I63071,I407102,I63097,I407105,I63114,I63122,I407120,I63139,I62971,I63170,I63187,I62983,I407123,I63227,I62992,I63249,I407114,I63266,I407108,I63292,I63309,I62995,I63331,I62980,I63362,I407117,I63379,I63396,I63413,I62989,I63444,I62977,I62986,I62974,I63530,I63556,I63564,I63581,I63598,I63624,I63641,I63649,I63666,I63498,I63697,I63714,I63510,I63754,I63519,I63776,I63793,I63819,I63836,I63522,I63858,I63507,I63889,I63906,I63923,I63940,I63516,I63971,I63504,I63513,I63501,I64057,I1009846,I64083,I64091,I64108,I1009864,I1009858,I64125,I1009837,I64151,I1009855,I64168,I64176,I1009840,I64193,I64025,I64224,I64241,I64037,I1009852,I64281,I64046,I64303,I1009861,I1009849,I64320,I1009843,I64346,I64363,I64049,I64385,I64034,I64416,I64433,I64450,I64467,I64043,I64498,I64031,I64040,I64028,I64584,I361807,I64610,I64618,I64635,I361789,I361804,I64652,I361780,I64678,I361783,I64695,I64703,I361798,I64720,I64552,I64751,I64768,I64564,I361801,I64808,I64573,I64830,I361792,I64847,I361786,I64873,I64890,I64576,I64912,I64561,I64943,I361795,I64960,I64977,I64994,I64570,I65025,I64558,I64567,I64555,I65111,I617384,I65137,I65145,I65162,I617396,I617381,I65179,I617375,I65205,I617390,I65222,I65230,I617378,I65247,I65079,I65278,I65295,I65091,I617387,I65335,I65100,I65357,I617393,I617399,I65374,I65400,I65417,I65103,I65439,I65088,I65470,I65487,I65504,I65521,I65097,I65552,I65085,I65094,I65082,I65638,I437652,I65664,I65672,I65689,I437646,I437637,I65706,I437658,I65732,I437640,I65749,I65757,I437634,I65774,I65606,I65805,I65822,I65618,I65862,I65627,I65884,I437661,I437643,I65901,I437649,I65927,I65944,I65630,I65966,I65615,I65997,I437655,I66014,I66031,I66048,I65624,I66079,I65612,I65621,I65609,I66165,I1286671,I66191,I66199,I66216,I1286665,I1286686,I66233,I1286677,I66259,I1286668,I66276,I66284,I1286680,I66301,I66133,I66332,I66349,I66145,I66389,I66154,I66411,I1286689,I1286674,I66428,I66454,I66471,I66157,I66493,I66142,I66524,I1286683,I66541,I66558,I66575,I66151,I66606,I66139,I66148,I66136,I66692,I226795,I66718,I66726,I66743,I226789,I226783,I66760,I226804,I66786,I226801,I66803,I66811,I226798,I66828,I66660,I66859,I66876,I66672,I66916,I66681,I66938,I226786,I66955,I226807,I66981,I66998,I66684,I67020,I66669,I67051,I226792,I67068,I67085,I67102,I66678,I67133,I66666,I66675,I66663,I67219,I891169,I67245,I67253,I67270,I891166,I891181,I67287,I891163,I67313,I891160,I67330,I67338,I67355,I67187,I67386,I67403,I67199,I67443,I67208,I67465,I891175,I67482,I891178,I67508,I67525,I67211,I67547,I67196,I67578,I891172,I67595,I67612,I67629,I67205,I67660,I67193,I67202,I67190,I67746,I1137241,I67772,I67780,I67797,I1137256,I1137235,I67814,I1137238,I67840,I1137259,I67857,I67865,I67882,I67714,I67913,I67930,I67726,I67970,I67735,I67992,I1137247,I1137244,I68009,I1137250,I68035,I68052,I67738,I68074,I67723,I68105,I1137253,I68122,I68139,I68156,I67732,I68187,I67720,I67729,I67717,I68273,I849009,I68299,I68307,I68324,I849006,I849021,I68341,I849003,I68367,I849000,I68384,I68392,I68409,I68241,I68440,I68457,I68253,I68497,I68262,I68519,I849015,I68536,I849018,I68562,I68579,I68265,I68601,I68250,I68632,I849012,I68649,I68666,I68683,I68259,I68714,I68247,I68256,I68244,I68800,I1258383,I68826,I68834,I68851,I1258377,I1258398,I68868,I1258389,I68894,I1258380,I68911,I68919,I1258392,I68936,I68768,I68967,I68984,I68780,I69024,I68789,I69046,I1258401,I1258386,I69063,I69089,I69106,I68792,I69128,I68777,I69159,I1258395,I69176,I69193,I69210,I68786,I69241,I68774,I68783,I68771,I69327,I1005324,I69353,I69361,I69378,I1005342,I1005336,I69395,I1005315,I69421,I1005333,I69438,I69446,I1005318,I69463,I69295,I69494,I69511,I69307,I1005330,I69551,I69316,I69573,I1005339,I1005327,I69590,I1005321,I69616,I69633,I69319,I69655,I69304,I69686,I69703,I69720,I69737,I69313,I69768,I69301,I69310,I69298,I69854,I1355340,I69880,I69888,I69905,I1355334,I1355355,I69922,I1355331,I69948,I1355352,I69965,I69973,I1355349,I69990,I69822,I70021,I70038,I69834,I1355337,I70078,I69843,I70100,I1355346,I1355343,I70117,I1355328,I70143,I70160,I69846,I70182,I69831,I70213,I70230,I70247,I70264,I69840,I70295,I69828,I69837,I69825,I70381,I1034394,I70407,I70415,I70432,I1034412,I1034406,I70449,I1034385,I70475,I1034403,I70492,I70500,I1034388,I70517,I70548,I70565,I1034400,I70605,I70627,I1034409,I1034397,I70644,I1034391,I70670,I70687,I70709,I70740,I70757,I70774,I70791,I70822,I70908,I1308582,I70934,I70942,I70959,I1308585,I1308579,I70976,I1308576,I71002,I1308561,I71019,I71027,I1308570,I71044,I70876,I71075,I71092,I70888,I71132,I70897,I71154,I1308564,I1308567,I71171,I1308573,I71197,I71214,I70900,I71236,I70885,I71267,I71284,I71301,I71318,I70894,I71349,I70882,I70891,I70879,I71435,I1127415,I71461,I71469,I71486,I1127430,I1127409,I71503,I1127412,I71529,I1127433,I71546,I71554,I71571,I71403,I71602,I71619,I71415,I71659,I71424,I71681,I1127421,I1127418,I71698,I1127424,I71724,I71741,I71427,I71763,I71412,I71794,I1127427,I71811,I71828,I71845,I71421,I71876,I71409,I71418,I71406,I71962,I358645,I71988,I71996,I72013,I358627,I358642,I72030,I358618,I72056,I358621,I72073,I72081,I358636,I72098,I71930,I72129,I72146,I71942,I358639,I72186,I71951,I72208,I358630,I72225,I358624,I72251,I72268,I71954,I72290,I71939,I72321,I358633,I72338,I72355,I72372,I71948,I72403,I71936,I71945,I71933,I72489,I72515,I72523,I72540,I72557,I72583,I72600,I72608,I72625,I72457,I72656,I72673,I72469,I72713,I72478,I72735,I72752,I72778,I72795,I72481,I72817,I72466,I72848,I72865,I72882,I72899,I72475,I72930,I72463,I72472,I72460,I73016,I208350,I73042,I73050,I73067,I208344,I208338,I73084,I208359,I73110,I208356,I73127,I73135,I208353,I73152,I72984,I73183,I73200,I72996,I73240,I73005,I73262,I208341,I73279,I208362,I73305,I73322,I73008,I73344,I72993,I73375,I208347,I73392,I73409,I73426,I73002,I73457,I72990,I72999,I72987,I73543,I887480,I73569,I73577,I73594,I887477,I887492,I73611,I887474,I73637,I887471,I73654,I73662,I73679,I73511,I73710,I73727,I73523,I73767,I73532,I73789,I887486,I73806,I887489,I73832,I73849,I73535,I73871,I73520,I73902,I887483,I73919,I73936,I73953,I73529,I73984,I73517,I73526,I73514,I74070,I526309,I74096,I74104,I74121,I526330,I526324,I74138,I526306,I74164,I74181,I74189,I526318,I74206,I74038,I74237,I74254,I74050,I526315,I74294,I74059,I74316,I526321,I526312,I74333,I74359,I74376,I74062,I74398,I74047,I74429,I526327,I74446,I74463,I74480,I74056,I74511,I74044,I74053,I74041,I74597,I206565,I74623,I74631,I74648,I206559,I206553,I74665,I206574,I74691,I206571,I74708,I74716,I206568,I74733,I74565,I74764,I74781,I74577,I74821,I74586,I74843,I206556,I74860,I206577,I74886,I74903,I74589,I74925,I74574,I74956,I206562,I74973,I74990,I75007,I74583,I75038,I74571,I74580,I74568,I75124,I75150,I75158,I75175,I75192,I75218,I75235,I75243,I75260,I75092,I75291,I75308,I75104,I75348,I75113,I75370,I75387,I75413,I75430,I75116,I75452,I75101,I75483,I75500,I75517,I75534,I75110,I75565,I75098,I75107,I75095,I75651,I471380,I75677,I75685,I75702,I471374,I471365,I75719,I471386,I75745,I471368,I75762,I75770,I471362,I75787,I75619,I75818,I75835,I75631,I75875,I75640,I75897,I471389,I471371,I75914,I471377,I75940,I75957,I75643,I75979,I75628,I76010,I471383,I76027,I76044,I76061,I75637,I76092,I75625,I75634,I75622,I76178,I254760,I76204,I76212,I76229,I254754,I254748,I76246,I254769,I76272,I254766,I76289,I76297,I254763,I76314,I76146,I76345,I76362,I76158,I76402,I76167,I76424,I254751,I76441,I254772,I76467,I76484,I76170,I76506,I76155,I76537,I254757,I76554,I76571,I76588,I76164,I76619,I76152,I76161,I76149,I76705,I379725,I76731,I76739,I76756,I379707,I379722,I76773,I379698,I76799,I379701,I76816,I76824,I379716,I76841,I76673,I76872,I76889,I76685,I379719,I76929,I76694,I76951,I379710,I76968,I379704,I76994,I77011,I76697,I77033,I76682,I77064,I379713,I77081,I77098,I77115,I76691,I77146,I76679,I76688,I76676,I77232,I1174811,I77258,I77266,I77283,I1174826,I1174805,I77300,I1174808,I77326,I1174829,I77343,I77351,I77368,I77200,I77399,I77416,I77212,I77456,I77221,I77478,I1174817,I1174814,I77495,I1174820,I77521,I77538,I77224,I77560,I77209,I77591,I1174823,I77608,I77625,I77642,I77218,I77673,I77206,I77215,I77203,I77759,I555464,I77785,I77793,I77810,I555485,I555479,I77827,I555461,I77853,I77870,I77878,I555473,I77895,I77727,I77926,I77943,I77739,I555470,I77983,I77748,I78005,I555476,I555467,I78022,I78048,I78065,I77751,I78087,I77736,I78118,I555482,I78135,I78152,I78169,I77745,I78200,I77733,I77742,I77730,I78286,I307526,I78312,I78320,I78337,I307508,I307523,I78354,I307499,I78380,I307502,I78397,I78405,I307517,I78422,I78254,I78453,I78470,I78266,I307520,I78510,I78275,I78532,I307511,I78549,I307505,I78575,I78592,I78278,I78614,I78263,I78645,I307514,I78662,I78679,I78696,I78272,I78727,I78260,I78269,I78257,I78813,I573314,I78839,I78847,I78864,I573335,I573329,I78881,I573311,I78907,I78924,I78932,I573323,I78949,I78781,I78980,I78997,I78793,I573320,I79037,I78802,I79059,I573326,I573317,I79076,I79102,I79119,I78805,I79141,I78790,I79172,I573332,I79189,I79206,I79223,I78799,I79254,I78787,I78796,I78784,I79340,I994988,I79366,I79374,I79391,I995006,I995000,I79408,I994979,I79434,I994997,I79451,I79459,I994982,I79476,I79308,I79507,I79524,I79320,I994994,I79564,I79329,I79586,I995003,I994991,I79603,I994985,I79629,I79646,I79332,I79668,I79317,I79699,I79716,I79733,I79750,I79326,I79781,I79314,I79323,I79311,I79867,I336511,I79893,I79901,I79918,I336493,I336508,I79935,I336484,I79961,I336487,I79978,I79986,I336502,I80003,I79835,I80034,I80051,I79847,I336505,I80091,I79856,I80113,I336496,I80130,I336490,I80156,I80173,I79859,I80195,I79844,I80226,I336499,I80243,I80260,I80277,I79853,I80308,I79841,I79850,I79838,I80394,I788475,I80420,I80428,I80445,I788466,I788484,I80462,I788463,I80488,I80505,I80513,I788469,I80530,I80362,I80561,I80578,I80374,I80618,I80383,I80640,I788481,I788472,I80657,I788487,I80683,I80700,I80386,I80722,I80371,I80753,I788478,I80770,I80787,I80804,I80380,I80835,I80368,I80377,I80365,I80921,I176220,I80947,I80955,I80972,I176214,I176208,I80989,I176229,I81015,I176226,I81032,I81040,I176223,I81057,I80889,I81088,I81105,I80901,I81145,I80910,I81167,I176211,I81184,I176232,I81210,I81227,I80913,I81249,I80898,I81280,I176217,I81297,I81314,I81331,I80907,I81362,I80895,I80904,I80892,I81448,I705243,I81474,I81482,I81499,I705234,I705252,I81516,I705231,I81542,I81559,I81567,I705237,I81584,I81416,I81615,I81632,I81428,I81672,I81437,I81694,I705249,I705240,I81711,I705255,I81737,I81754,I81440,I81776,I81425,I81807,I705246,I81824,I81841,I81858,I81434,I81889,I81422,I81431,I81419,I81975,I556059,I82001,I82009,I82026,I556080,I556074,I82043,I556056,I82069,I82086,I82094,I556068,I82111,I81943,I82142,I82159,I81955,I556065,I82199,I81964,I82221,I556071,I556062,I82238,I82264,I82281,I81967,I82303,I81952,I82334,I556077,I82351,I82368,I82385,I81961,I82416,I81949,I81958,I81946,I82502,I342308,I82528,I82536,I82553,I342290,I342305,I82570,I342281,I82596,I342284,I82613,I82621,I342299,I82638,I82669,I82686,I342302,I82726,I82748,I342293,I82765,I342287,I82791,I82808,I82830,I82861,I342296,I82878,I82895,I82912,I82943,I83029,I858495,I83055,I83063,I83080,I858492,I858507,I83097,I858489,I83123,I858486,I83140,I83148,I83165,I83196,I83213,I83253,I83275,I858501,I83292,I858504,I83318,I83335,I83357,I83388,I858498,I83405,I83422,I83439,I83470,I83556,I624898,I83582,I83590,I83607,I624910,I624895,I83624,I624889,I83650,I624904,I83667,I83675,I624892,I83692,I83524,I83723,I83740,I83536,I624901,I83780,I83545,I83802,I624907,I624913,I83819,I83845,I83862,I83548,I83884,I83533,I83915,I83932,I83949,I83966,I83542,I83997,I83530,I83539,I83527,I84083,I1347010,I84109,I84117,I84134,I1347004,I1347025,I84151,I1347001,I84177,I1347022,I84194,I84202,I1347019,I84219,I84051,I84250,I84267,I84063,I1347007,I84307,I84072,I84329,I1347016,I1347013,I84346,I1346998,I84372,I84389,I84075,I84411,I84060,I84442,I84459,I84476,I84493,I84069,I84524,I84057,I84066,I84054,I84610,I205970,I84636,I84644,I84661,I205964,I205958,I84678,I205979,I84704,I205976,I84721,I84729,I205973,I84746,I84578,I84777,I84794,I84590,I84834,I84599,I84856,I205961,I84873,I205982,I84899,I84916,I84602,I84938,I84587,I84969,I205967,I84986,I85003,I85020,I84596,I85051,I84584,I84593,I84581,I85137,I1204867,I85163,I85171,I85188,I1204882,I1204861,I85205,I1204864,I85231,I1204885,I85248,I85256,I85273,I85105,I85304,I85321,I85117,I85361,I85126,I85383,I1204873,I1204870,I85400,I1204876,I85426,I85443,I85129,I85465,I85114,I85496,I1204879,I85513,I85530,I85547,I85123,I85578,I85111,I85120,I85108,I85664,I755529,I85690,I85698,I85715,I755520,I755538,I85732,I755517,I85758,I85775,I85783,I755523,I85800,I85632,I85831,I85848,I85644,I85888,I85653,I85910,I755535,I755526,I85927,I755541,I85953,I85970,I85656,I85992,I85641,I86023,I755532,I86040,I86057,I86074,I85650,I86105,I85638,I85647,I85635,I86191,I1189261,I86217,I86225,I86242,I1189276,I1189255,I86259,I1189258,I86285,I1189279,I86302,I86310,I86327,I86358,I86375,I86415,I86437,I1189267,I1189264,I86454,I1189270,I86480,I86497,I86519,I86550,I1189273,I86567,I86584,I86601,I86632,I86718,I1088176,I86744,I86752,I86769,I1088173,I1088179,I86786,I86812,I86829,I86837,I86854,I86686,I86885,I86902,I86698,I1088182,I86942,I86707,I86964,I1088185,I1088194,I86981,I1088188,I87007,I87024,I86710,I87046,I86695,I87077,I1088191,I87094,I87111,I87128,I86704,I87159,I86692,I86701,I86689,I87245,I446900,I87271,I87279,I87296,I446894,I446885,I87313,I446906,I87339,I446888,I87356,I87364,I446882,I87381,I87213,I87412,I87429,I87225,I87469,I87234,I87491,I446909,I446891,I87508,I446897,I87534,I87551,I87237,I87573,I87222,I87604,I446903,I87621,I87638,I87655,I87231,I87686,I87219,I87228,I87216,I87772,I468660,I87798,I87806,I87823,I468654,I468645,I87840,I468666,I87866,I468648,I87883,I87891,I468642,I87908,I87740,I87939,I87956,I87752,I87996,I87761,I88018,I468669,I468651,I88035,I468657,I88061,I88078,I87764,I88100,I87749,I88131,I468663,I88148,I88165,I88182,I87758,I88213,I87746,I87755,I87743,I88299,I803503,I88325,I88333,I88350,I803494,I803512,I88367,I803491,I88393,I88410,I88418,I803497,I88435,I88267,I88466,I88483,I88279,I88523,I88288,I88545,I803509,I803500,I88562,I803515,I88588,I88605,I88291,I88627,I88276,I88658,I803506,I88675,I88692,I88709,I88285,I88740,I88273,I88282,I88270,I88826,I364442,I88852,I88860,I88877,I364424,I364439,I88894,I364415,I88920,I364418,I88937,I88945,I364433,I88962,I88794,I88993,I89010,I88806,I364436,I89050,I88815,I89072,I364427,I89089,I364421,I89115,I89132,I88818,I89154,I88803,I89185,I364430,I89202,I89219,I89236,I88812,I89267,I88800,I88809,I88797,I89353,I89379,I89387,I89404,I89421,I89447,I89464,I89472,I89489,I89321,I89520,I89537,I89333,I89577,I89342,I89599,I89616,I89642,I89659,I89345,I89681,I89330,I89712,I89729,I89746,I89763,I89339,I89794,I89327,I89336,I89324,I89880,I749171,I89906,I89914,I89931,I749162,I749180,I89948,I749159,I89974,I89991,I89999,I749165,I90016,I89848,I90047,I90064,I89860,I90104,I89869,I90126,I749177,I749168,I90143,I749183,I90169,I90186,I89872,I90208,I89857,I90239,I749174,I90256,I90273,I90290,I89866,I90321,I89854,I89863,I89851,I90407,I257735,I90433,I90441,I90458,I257729,I257723,I90475,I257744,I90501,I257741,I90518,I90526,I257738,I90543,I90375,I90574,I90591,I90387,I90631,I90396,I90653,I257726,I90670,I257747,I90696,I90713,I90399,I90735,I90384,I90766,I257732,I90783,I90800,I90817,I90393,I90848,I90381,I90390,I90378,I90934,I654954,I90960,I90968,I90985,I654966,I654951,I91002,I654945,I91028,I654960,I91045,I91053,I654948,I91070,I90902,I91101,I91118,I90914,I654957,I91158,I90923,I91180,I654963,I654969,I91197,I91223,I91240,I90926,I91262,I90911,I91293,I91310,I91327,I91344,I90920,I91375,I90908,I90917,I90905,I91461,I1271983,I91487,I91495,I91512,I1271977,I1271998,I91529,I1271989,I91555,I1271980,I91572,I91580,I1271992,I91597,I91429,I91628,I91645,I91441,I91685,I91450,I91707,I1272001,I1271986,I91724,I91750,I91767,I91453,I91789,I91438,I91820,I1271995,I91837,I91854,I91871,I91447,I91902,I91435,I91444,I91432,I91988,I92014,I92022,I92039,I92056,I92082,I92099,I92107,I92124,I91956,I92155,I92172,I91968,I92212,I91977,I92234,I92251,I92277,I92294,I91980,I92316,I91965,I92347,I92364,I92381,I92398,I91974,I92429,I91962,I91971,I91959,I92515,I508372,I92541,I92549,I92566,I508366,I508357,I92583,I508378,I92609,I508360,I92626,I92634,I508354,I92651,I92483,I92682,I92699,I92495,I92739,I92504,I92761,I508381,I508363,I92778,I508369,I92804,I92821,I92507,I92843,I92492,I92874,I508375,I92891,I92908,I92925,I92501,I92956,I92489,I92498,I92486,I93042,I219655,I93068,I93076,I93093,I219649,I219643,I93110,I219664,I93136,I219661,I93153,I93161,I219658,I93178,I93010,I93209,I93226,I93022,I93266,I93031,I93288,I219646,I93305,I219667,I93331,I93348,I93034,I93370,I93019,I93401,I219652,I93418,I93435,I93452,I93028,I93483,I93016,I93025,I93013,I93569,I1223363,I93595,I93603,I93620,I1223378,I1223357,I93637,I1223360,I93663,I1223381,I93680,I93688,I93705,I93537,I93736,I93753,I93549,I93793,I93558,I93815,I1223369,I1223366,I93832,I1223372,I93858,I93875,I93561,I93897,I93546,I93928,I1223375,I93945,I93962,I93979,I93555,I94010,I93543,I93552,I93540,I94096,I1007908,I94122,I94130,I94147,I1007926,I1007920,I94164,I1007899,I94190,I1007917,I94207,I94215,I1007902,I94232,I94064,I94263,I94280,I94076,I1007914,I94320,I94085,I94342,I1007923,I1007911,I94359,I1007905,I94385,I94402,I94088,I94424,I94073,I94455,I94472,I94489,I94506,I94082,I94537,I94070,I94079,I94067,I94623,I1273615,I94649,I94657,I94674,I1273609,I1273630,I94691,I1273621,I94717,I1273612,I94734,I94742,I1273624,I94759,I94591,I94790,I94807,I94603,I94847,I94612,I94869,I1273633,I1273618,I94886,I94912,I94929,I94615,I94951,I94600,I94982,I1273627,I94999,I95016,I95033,I94609,I95064,I94597,I94606,I94594,I95150,I1125681,I95176,I95184,I95201,I1125696,I1125675,I95218,I1125678,I95244,I1125699,I95261,I95269,I95286,I95118,I95317,I95334,I95130,I95374,I95139,I95396,I1125687,I1125684,I95413,I1125690,I95439,I95456,I95142,I95478,I95127,I95509,I1125693,I95526,I95543,I95560,I95136,I95591,I95124,I95133,I95121,I95677,I166700,I95703,I95711,I95728,I166694,I166688,I95745,I166709,I95771,I166706,I95788,I95796,I166703,I95813,I95645,I95844,I95861,I95657,I95901,I95666,I95923,I166691,I95940,I166712,I95966,I95983,I95669,I96005,I95654,I96036,I166697,I96053,I96070,I96087,I95663,I96118,I95651,I95660,I95648,I96204,I807549,I96230,I96238,I96255,I807540,I807558,I96272,I807537,I96298,I96315,I96323,I807543,I96340,I96172,I96371,I96388,I96184,I96428,I96193,I96450,I807555,I807546,I96467,I807561,I96493,I96510,I96196,I96532,I96181,I96563,I807552,I96580,I96597,I96614,I96190,I96645,I96178,I96187,I96175,I96731,I601200,I96757,I96765,I96782,I601212,I601197,I96799,I601191,I96825,I601206,I96842,I96850,I601194,I96867,I96699,I96898,I96915,I96711,I601203,I96955,I96720,I96977,I601209,I601215,I96994,I97020,I97037,I96723,I97059,I96708,I97090,I97107,I97124,I97141,I96717,I97172,I96705,I96714,I96702,I97258,I175030,I97284,I97292,I97309,I175024,I175018,I97326,I175039,I97352,I175036,I97369,I97377,I175033,I97394,I97425,I97442,I97482,I97504,I175021,I97521,I175042,I97547,I97564,I97586,I97617,I175027,I97634,I97651,I97668,I97699,I97785,I97811,I97819,I97836,I97853,I97879,I97896,I97904,I97921,I97753,I97952,I97969,I97765,I98009,I97774,I98031,I98048,I98074,I98091,I97777,I98113,I97762,I98144,I98161,I98178,I98195,I97771,I98226,I97759,I97768,I97756,I98312,I832145,I98338,I98346,I98363,I832142,I832157,I98380,I832139,I98406,I832136,I98423,I98431,I98448,I98280,I98479,I98496,I98292,I98536,I98301,I98558,I832151,I98575,I832154,I98601,I98618,I98304,I98640,I98289,I98671,I832148,I98688,I98705,I98722,I98298,I98753,I98286,I98295,I98283,I98839,I285105,I98865,I98873,I98890,I285099,I285093,I98907,I285114,I98933,I285111,I98950,I98958,I285108,I98975,I98807,I99006,I99023,I98819,I99063,I98828,I99085,I285096,I99102,I285117,I99128,I99145,I98831,I99167,I98816,I99198,I285102,I99215,I99232,I99249,I98825,I99280,I98813,I98822,I98810,I99366,I1345820,I99392,I99400,I99417,I1345814,I1345835,I99434,I1345811,I99460,I1345832,I99477,I99485,I1345829,I99502,I99334,I99533,I99550,I99346,I1345817,I99590,I99355,I99612,I1345826,I1345823,I99629,I1345808,I99655,I99672,I99358,I99694,I99343,I99725,I99742,I99759,I99776,I99352,I99807,I99340,I99349,I99337,I99893,I299621,I99919,I99927,I99944,I299603,I299618,I99961,I299594,I99987,I299597,I100004,I100012,I299612,I100029,I99861,I100060,I100077,I99873,I299615,I100117,I99882,I100139,I299606,I100156,I299600,I100182,I100199,I99885,I100221,I99870,I100252,I299609,I100269,I100286,I100303,I99879,I100334,I99867,I99876,I99864,I100420,I1401155,I100446,I100454,I100471,I1401149,I1401170,I100488,I1401146,I100514,I1401167,I100531,I100539,I1401164,I100556,I100388,I100587,I100604,I100400,I1401152,I100644,I100409,I100666,I1401161,I1401158,I100683,I1401143,I100709,I100726,I100412,I100748,I100397,I100779,I100796,I100813,I100830,I100406,I100861,I100394,I100403,I100391,I100947,I692527,I100973,I100981,I100998,I692518,I692536,I101015,I692515,I101041,I101058,I101066,I692521,I101083,I100915,I101114,I101131,I100927,I101171,I100936,I101193,I692533,I692524,I101210,I692539,I101236,I101253,I100939,I101275,I100924,I101306,I692530,I101323,I101340,I101357,I100933,I101388,I100921,I100930,I100918,I101474,I826875,I101500,I101508,I101525,I826872,I826887,I101542,I826869,I101568,I826866,I101585,I101593,I101610,I101442,I101641,I101658,I101454,I101698,I101463,I101720,I826881,I101737,I826884,I101763,I101780,I101466,I101802,I101451,I101833,I826878,I101850,I101867,I101884,I101460,I101915,I101448,I101457,I101445,I102001,I102027,I102035,I102052,I102069,I102095,I102112,I102120,I102137,I101969,I102168,I102185,I101981,I102225,I101990,I102247,I102264,I102290,I102307,I101993,I102329,I101978,I102360,I102377,I102394,I102411,I101987,I102442,I101975,I101984,I101972,I102528,I484980,I102554,I102562,I102579,I484974,I484965,I102596,I484986,I102622,I484968,I102639,I102647,I484962,I102664,I102496,I102695,I102712,I102508,I102752,I102517,I102774,I484989,I484971,I102791,I484977,I102817,I102834,I102520,I102856,I102505,I102887,I484983,I102904,I102921,I102938,I102514,I102969,I102502,I102511,I102499,I103055,I1333325,I103081,I103089,I103106,I1333319,I1333340,I103123,I1333316,I103149,I1333337,I103166,I103174,I1333334,I103191,I103023,I103222,I103239,I103035,I1333322,I103279,I103044,I103301,I1333331,I1333328,I103318,I1333313,I103344,I103361,I103047,I103383,I103032,I103414,I103431,I103448,I103465,I103041,I103496,I103029,I103038,I103026,I103582,I429492,I103608,I103616,I103633,I429486,I429477,I103650,I429498,I103676,I429480,I103693,I103701,I429474,I103718,I103550,I103749,I103766,I103562,I103806,I103571,I103828,I429501,I429483,I103845,I429489,I103871,I103888,I103574,I103910,I103559,I103941,I429495,I103958,I103975,I103992,I103568,I104023,I103556,I103565,I103553,I104109,I996280,I104135,I104143,I104160,I996298,I996292,I104177,I996271,I104203,I996289,I104220,I104228,I996274,I104245,I104276,I104293,I996286,I104333,I104355,I996295,I996283,I104372,I996277,I104398,I104415,I104437,I104468,I104485,I104502,I104519,I104550,I104636,I793677,I104662,I104670,I104687,I793668,I793686,I104704,I793665,I104730,I104747,I104755,I793671,I104772,I104604,I104803,I104820,I104616,I104860,I104625,I104882,I793683,I793674,I104899,I793689,I104925,I104942,I104628,I104964,I104613,I104995,I793680,I105012,I105029,I105046,I104622,I105077,I104610,I104619,I104607,I105163,I211920,I105189,I105197,I105214,I211914,I211908,I105231,I211929,I105257,I211926,I105274,I105282,I211923,I105299,I105131,I105330,I105347,I105143,I105387,I105152,I105409,I211911,I105426,I211932,I105452,I105469,I105155,I105491,I105140,I105522,I211917,I105539,I105556,I105573,I105149,I105604,I105137,I105146,I105134,I105690,I635880,I105716,I105724,I105741,I635892,I635877,I105758,I635871,I105784,I635886,I105801,I105809,I635874,I105826,I105658,I105857,I105874,I105670,I635883,I105914,I105679,I105936,I635889,I635895,I105953,I105979,I105996,I105682,I106018,I105667,I106049,I106066,I106083,I106100,I105676,I106131,I105664,I105673,I105661,I106217,I778071,I106243,I106251,I106268,I778062,I778080,I106285,I778059,I106311,I106328,I106336,I778065,I106353,I106185,I106384,I106401,I106197,I106441,I106206,I106463,I778077,I778068,I106480,I778083,I106506,I106523,I106209,I106545,I106194,I106576,I778074,I106593,I106610,I106627,I106203,I106658,I106191,I106200,I106188,I106744,I669985,I106770,I106778,I106795,I669976,I669994,I106812,I669973,I106838,I106855,I106863,I669979,I106880,I106712,I106911,I106928,I106724,I106968,I106733,I106990,I669991,I669982,I107007,I669997,I107033,I107050,I106736,I107072,I106721,I107103,I669988,I107120,I107137,I107154,I106730,I107185,I106718,I106727,I106715,I107271,I517620,I107297,I107305,I107322,I517614,I517605,I107339,I517626,I107365,I517608,I107382,I107390,I517602,I107407,I107239,I107438,I107455,I107251,I107495,I107260,I107517,I517629,I517611,I107534,I517617,I107560,I107577,I107263,I107599,I107248,I107630,I517623,I107647,I107664,I107681,I107257,I107712,I107245,I107254,I107242,I107798,I333876,I107824,I107832,I107849,I333858,I333873,I107866,I333849,I107892,I333852,I107909,I107917,I333867,I107934,I107766,I107965,I107982,I107778,I333870,I108022,I107787,I108044,I333861,I108061,I333855,I108087,I108104,I107790,I108126,I107775,I108157,I333864,I108174,I108191,I108208,I107784,I108239,I107772,I107781,I107769,I108325,I108351,I108359,I108376,I108393,I108419,I108436,I108444,I108461,I108293,I108492,I108509,I108305,I108549,I108314,I108571,I108588,I108614,I108631,I108317,I108653,I108302,I108684,I108701,I108718,I108735,I108311,I108766,I108299,I108308,I108296,I108852,I1031164,I108878,I108886,I108903,I1031182,I1031176,I108920,I1031155,I108946,I1031173,I108963,I108971,I1031158,I108988,I108820,I109019,I109036,I108832,I1031170,I109076,I108841,I109098,I1031179,I1031167,I109115,I1031161,I109141,I109158,I108844,I109180,I108829,I109211,I109228,I109245,I109262,I108838,I109293,I108826,I108835,I108823,I109379,I1394015,I109405,I109413,I109430,I1394009,I1394030,I109447,I1394006,I109473,I1394027,I109490,I109498,I1394024,I109515,I109347,I109546,I109563,I109359,I1394012,I109603,I109368,I109625,I1394021,I1394018,I109642,I1394003,I109668,I109685,I109371,I109707,I109356,I109738,I109755,I109772,I109789,I109365,I109820,I109353,I109362,I109350,I109906,I638770,I109932,I109940,I109957,I638782,I638767,I109974,I638761,I110000,I638776,I110017,I110025,I638764,I110042,I109874,I110073,I110090,I109886,I638773,I110130,I109895,I110152,I638779,I638785,I110169,I110195,I110212,I109898,I110234,I109883,I110265,I110282,I110299,I110316,I109892,I110347,I109880,I109889,I109877,I110433,I168485,I110459,I110467,I110484,I168479,I168473,I110501,I168494,I110527,I168491,I110544,I110552,I168488,I110569,I110401,I110600,I110617,I110413,I110657,I110422,I110679,I168476,I110696,I168497,I110722,I110739,I110425,I110761,I110410,I110792,I168482,I110809,I110826,I110843,I110419,I110874,I110407,I110416,I110404,I110960,I985944,I110986,I110994,I111011,I985962,I985956,I111028,I985935,I111054,I985953,I111071,I111079,I985938,I111096,I110928,I111127,I111144,I110940,I985950,I111184,I110949,I111206,I985959,I985947,I111223,I985941,I111249,I111266,I110952,I111288,I110937,I111319,I111336,I111353,I111370,I110946,I111401,I110934,I110943,I110931,I111487,I1178857,I111513,I111521,I111538,I1178872,I1178851,I111555,I1178854,I111581,I1178875,I111598,I111606,I111623,I111455,I111654,I111671,I111467,I111711,I111476,I111733,I1178863,I1178860,I111750,I1178866,I111776,I111793,I111479,I111815,I111464,I111846,I1178869,I111863,I111880,I111897,I111473,I111928,I111461,I111470,I111458,I112014,I1240125,I112040,I112048,I112065,I1240140,I1240119,I112082,I1240122,I112108,I1240143,I112125,I112133,I112150,I111982,I112181,I112198,I111994,I112238,I112003,I112260,I1240131,I1240128,I112277,I1240134,I112303,I112320,I112006,I112342,I111991,I112373,I1240137,I112390,I112407,I112424,I112000,I112455,I111988,I111997,I111985,I112541,I787897,I112567,I112575,I112592,I787888,I787906,I112609,I787885,I112635,I112652,I112660,I787891,I112677,I112509,I112708,I112725,I112521,I112765,I112530,I112787,I787903,I787894,I112804,I787909,I112830,I112847,I112533,I112869,I112518,I112900,I787900,I112917,I112934,I112951,I112527,I112982,I112515,I112524,I112512,I113068,I277370,I113094,I113102,I113119,I277364,I277358,I113136,I277379,I113162,I277376,I113179,I113187,I277373,I113204,I113036,I113235,I113252,I113048,I113292,I113057,I113314,I277361,I113331,I277382,I113357,I113374,I113060,I113396,I113045,I113427,I277367,I113444,I113461,I113478,I113054,I113509,I113042,I113051,I113039,I113595,I1329777,I113621,I113629,I113646,I1329783,I1329801,I113663,I1329798,I113689,I1329795,I113706,I113714,I1329789,I113731,I113563,I113762,I113779,I113575,I113819,I113584,I113841,I1329792,I1329780,I113858,I1329804,I113884,I113901,I113587,I113923,I113572,I113954,I1329786,I113971,I113988,I114005,I113581,I114036,I113569,I113578,I113566,I114122,I633568,I114148,I114156,I114173,I633580,I633565,I114190,I633559,I114216,I633574,I114233,I114241,I633562,I114258,I114090,I114289,I114306,I114102,I633571,I114346,I114111,I114368,I633577,I633583,I114385,I114411,I114428,I114114,I114450,I114099,I114481,I114498,I114515,I114532,I114108,I114563,I114096,I114105,I114093,I114649,I908560,I114675,I114683,I114700,I908557,I908572,I114717,I908554,I114743,I908551,I114760,I114768,I114785,I114617,I114816,I114833,I114629,I114873,I114638,I114895,I908566,I114912,I908569,I114938,I114955,I114641,I114977,I114626,I115008,I908563,I115025,I115042,I115059,I114635,I115090,I114623,I114632,I114620,I115176,I365496,I115202,I115210,I115227,I365478,I365493,I115244,I365469,I115270,I365472,I115287,I115295,I365487,I115312,I115144,I115343,I115360,I115156,I365490,I115400,I115165,I115422,I365481,I115439,I365475,I115465,I115482,I115168,I115504,I115153,I115535,I365484,I115552,I115569,I115586,I115162,I115617,I115150,I115159,I115147,I115703,I466484,I115729,I115737,I115754,I466478,I466469,I115771,I466490,I115797,I466472,I115814,I115822,I466466,I115839,I115671,I115870,I115887,I115683,I115927,I115692,I115949,I466493,I466475,I115966,I466481,I115992,I116009,I115695,I116031,I115680,I116062,I466487,I116079,I116096,I116113,I115689,I116144,I115677,I115686,I115674,I116230,I361280,I116256,I116264,I116281,I361262,I361277,I116298,I361253,I116324,I361256,I116341,I116349,I361271,I116366,I116198,I116397,I116414,I116210,I361274,I116454,I116219,I116476,I361265,I116493,I361259,I116519,I116536,I116222,I116558,I116207,I116589,I361268,I116606,I116623,I116640,I116216,I116671,I116204,I116213,I116201,I116757,I1065736,I116783,I116791,I116808,I1065733,I1065739,I116825,I116851,I116868,I116876,I116893,I116725,I116924,I116941,I116737,I1065742,I116981,I116746,I117003,I1065745,I1065754,I117020,I1065748,I117046,I117063,I116749,I117085,I116734,I117116,I1065751,I117133,I117150,I117167,I116743,I117198,I116731,I116740,I116728,I117284,I562604,I117310,I117318,I117335,I562625,I562619,I117352,I562601,I117378,I117395,I117403,I562613,I117420,I117252,I117451,I117468,I117264,I562610,I117508,I117273,I117530,I562616,I562607,I117547,I117573,I117590,I117276,I117612,I117261,I117643,I562622,I117660,I117677,I117694,I117270,I117725,I117258,I117267,I117255,I117811,I322809,I117837,I117845,I117862,I322791,I322806,I117879,I322782,I117905,I322785,I117922,I117930,I322800,I117947,I117779,I117978,I117995,I117791,I322803,I118035,I117800,I118057,I322794,I118074,I322788,I118100,I118117,I117803,I118139,I117788,I118170,I322797,I118187,I118204,I118221,I117797,I118252,I117785,I117794,I117782,I118338,I671141,I118364,I118372,I118389,I671132,I671150,I118406,I671129,I118432,I118449,I118457,I671135,I118474,I118306,I118505,I118522,I118318,I118562,I118327,I118584,I671147,I671138,I118601,I671153,I118627,I118644,I118330,I118666,I118315,I118697,I671144,I118714,I118731,I118748,I118324,I118779,I118312,I118321,I118309,I118865,I1265455,I118891,I118899,I118916,I1265449,I1265470,I118933,I1265461,I118959,I1265452,I118976,I118984,I1265464,I119001,I118833,I119032,I119049,I118845,I119089,I118854,I119111,I1265473,I1265458,I119128,I119154,I119171,I118857,I119193,I118842,I119224,I1265467,I119241,I119258,I119275,I118851,I119306,I118839,I118848,I118836,I119392,I822132,I119418,I119426,I119443,I822129,I822144,I119460,I822126,I119486,I822123,I119503,I119511,I119528,I119360,I119559,I119576,I119372,I119616,I119381,I119638,I822138,I119655,I822141,I119681,I119698,I119384,I119720,I119369,I119751,I822135,I119768,I119785,I119802,I119378,I119833,I119366,I119375,I119363,I119919,I510548,I119945,I119953,I119970,I510542,I510533,I119987,I510554,I120013,I510536,I120030,I120038,I510530,I120055,I119887,I120086,I120103,I119899,I120143,I119908,I120165,I510557,I510539,I120182,I510545,I120208,I120225,I119911,I120247,I119896,I120278,I510551,I120295,I120312,I120329,I119905,I120360,I119893,I119902,I119890,I120446,I377090,I120472,I120480,I120497,I377072,I377087,I120514,I377063,I120540,I377066,I120557,I120565,I377081,I120582,I120414,I120613,I120630,I120426,I377084,I120670,I120435,I120692,I377075,I120709,I377069,I120735,I120752,I120438,I120774,I120423,I120805,I377078,I120822,I120839,I120856,I120432,I120887,I120420,I120429,I120417,I120973,I725473,I120999,I121007,I121024,I725464,I725482,I121041,I725461,I121067,I121084,I121092,I725467,I121109,I120941,I121140,I121157,I120953,I121197,I120962,I121219,I725479,I725470,I121236,I725485,I121262,I121279,I120965,I121301,I120950,I121332,I725476,I121349,I121366,I121383,I120959,I121414,I120947,I120956,I120944,I121500,I783851,I121526,I121534,I121551,I783842,I783860,I121568,I783839,I121594,I121611,I121619,I783845,I121636,I121468,I121667,I121684,I121480,I121724,I121489,I121746,I783857,I783848,I121763,I783863,I121789,I121806,I121492,I121828,I121477,I121859,I783854,I121876,I121893,I121910,I121486,I121941,I121474,I121483,I121471,I122027,I430580,I122053,I122061,I122078,I430574,I430565,I122095,I430586,I122121,I430568,I122138,I122146,I430562,I122163,I121995,I122194,I122211,I122007,I122251,I122016,I122273,I430589,I430571,I122290,I430577,I122316,I122333,I122019,I122355,I122004,I122386,I430583,I122403,I122420,I122437,I122013,I122468,I122001,I122010,I121998,I122554,I957520,I122580,I122588,I122605,I957538,I957532,I122622,I957511,I122648,I957529,I122665,I122673,I957514,I122690,I122522,I122721,I122738,I122534,I957526,I122778,I122543,I122800,I957535,I957523,I122817,I957517,I122843,I122860,I122546,I122882,I122531,I122913,I122930,I122947,I122964,I122540,I122995,I122528,I122537,I122525,I123081,I1243015,I123107,I123115,I123132,I1243030,I1243009,I123149,I1243012,I123175,I1243033,I123192,I123200,I123217,I123049,I123248,I123265,I123061,I123305,I123070,I123327,I1243021,I1243018,I123344,I1243024,I123370,I123387,I123073,I123409,I123058,I123440,I1243027,I123457,I123474,I123491,I123067,I123522,I123055,I123064,I123052,I123608,I615072,I123634,I123642,I123659,I615084,I615069,I123676,I615063,I123702,I615078,I123719,I123727,I615066,I123744,I123576,I123775,I123792,I123588,I615075,I123832,I123597,I123854,I615081,I615087,I123871,I123897,I123914,I123600,I123936,I123585,I123967,I123984,I124001,I124018,I123594,I124049,I123582,I123591,I123579,I124135,I1169609,I124161,I124169,I124186,I1169624,I1169603,I124203,I1169606,I124229,I1169627,I124246,I124254,I124271,I124103,I124302,I124319,I124115,I124359,I124124,I124381,I1169615,I1169612,I124398,I1169618,I124424,I124441,I124127,I124463,I124112,I124494,I1169621,I124511,I124528,I124545,I124121,I124576,I124109,I124118,I124106,I124662,I898547,I124688,I124696,I124713,I898544,I898559,I124730,I898541,I124756,I898538,I124773,I124781,I124798,I124630,I124829,I124846,I124642,I124886,I124651,I124908,I898553,I124925,I898556,I124951,I124968,I124654,I124990,I124639,I125021,I898550,I125038,I125055,I125072,I124648,I125103,I124636,I124645,I124633,I125189,I125215,I125223,I125240,I125257,I125283,I125300,I125308,I125325,I125157,I125356,I125373,I125169,I125413,I125178,I125435,I125452,I125478,I125495,I125181,I125517,I125166,I125548,I125565,I125582,I125599,I125175,I125630,I125163,I125172,I125160,I125716,I639926,I125742,I125750,I125767,I639938,I639923,I125784,I639917,I125810,I639932,I125827,I125835,I639920,I125852,I125684,I125883,I125900,I125696,I639929,I125940,I125705,I125962,I639935,I639941,I125979,I126005,I126022,I125708,I126044,I125693,I126075,I126092,I126109,I126126,I125702,I126157,I125690,I125699,I125687,I126243,I823186,I126269,I126277,I126294,I823183,I823198,I126311,I823180,I126337,I823177,I126354,I126362,I126379,I126211,I126410,I126427,I126223,I126467,I126232,I126489,I823192,I126506,I823195,I126532,I126549,I126235,I126571,I126220,I126602,I823189,I126619,I126636,I126653,I126229,I126684,I126217,I126226,I126214,I126770,I483892,I126796,I126804,I126821,I483886,I483877,I126838,I483898,I126864,I483880,I126881,I126889,I483874,I126906,I126738,I126937,I126954,I126750,I126994,I126759,I127016,I483901,I483883,I127033,I483889,I127059,I127076,I126762,I127098,I126747,I127129,I483895,I127146,I127163,I127180,I126756,I127211,I126744,I126753,I126741,I127297,I1133195,I127323,I127331,I127348,I1133210,I1133189,I127365,I1133192,I127391,I1133213,I127408,I127416,I127433,I127265,I127464,I127481,I127277,I127521,I127286,I127543,I1133201,I1133198,I127560,I1133204,I127586,I127603,I127289,I127625,I127274,I127656,I1133207,I127673,I127690,I127707,I127283,I127738,I127271,I127280,I127268,I127824,I1024704,I127850,I127858,I127875,I1024722,I1024716,I127892,I1024695,I127918,I1024713,I127935,I127943,I1024698,I127960,I127792,I127991,I128008,I127804,I1024710,I128048,I127813,I128070,I1024719,I1024707,I128087,I1024701,I128113,I128130,I127816,I128152,I127801,I128183,I128200,I128217,I128234,I127810,I128265,I127798,I127807,I127795,I128351,I608714,I128377,I128385,I128402,I608726,I608711,I128419,I608705,I128445,I608720,I128462,I128470,I608708,I128487,I128319,I128518,I128535,I128331,I608717,I128575,I128340,I128597,I608723,I608729,I128614,I128640,I128657,I128343,I128679,I128328,I128710,I128727,I128744,I128761,I128337,I128792,I128325,I128334,I128322,I128878,I360753,I128904,I128912,I128929,I360735,I360750,I128946,I360726,I128972,I360729,I128989,I128997,I360744,I129014,I128846,I129045,I129062,I128858,I360747,I129102,I128867,I129124,I360738,I129141,I360732,I129167,I129184,I128870,I129206,I128855,I129237,I360741,I129254,I129271,I129288,I128864,I129319,I128852,I128861,I128849,I129405,I635302,I129431,I129439,I129456,I635314,I635299,I129473,I635293,I129499,I635308,I129516,I129524,I635296,I129541,I129373,I129572,I129589,I129385,I635305,I129629,I129394,I129651,I635311,I635317,I129668,I129694,I129711,I129397,I129733,I129382,I129764,I129781,I129798,I129815,I129391,I129846,I129379,I129388,I129376,I129932,I974316,I129958,I129966,I129983,I974334,I974328,I130000,I974307,I130026,I974325,I130043,I130051,I974310,I130068,I129900,I130099,I130116,I129912,I974322,I130156,I129921,I130178,I974331,I974319,I130195,I974313,I130221,I130238,I129924,I130260,I129909,I130291,I130308,I130325,I130342,I129918,I130373,I129906,I129915,I129903,I130459,I953644,I130485,I130493,I130510,I953662,I953656,I130527,I953635,I130553,I953653,I130570,I130578,I953638,I130595,I130427,I130626,I130643,I130439,I953650,I130683,I130448,I130705,I953659,I953647,I130722,I953641,I130748,I130765,I130451,I130787,I130436,I130818,I130835,I130852,I130869,I130445,I130900,I130433,I130442,I130430,I130986,I131012,I131020,I131037,I131054,I131080,I131097,I131105,I131122,I130954,I131153,I131170,I130966,I131210,I130975,I131232,I131249,I131275,I131292,I130978,I131314,I130963,I131345,I131362,I131379,I131396,I130972,I131427,I130960,I130969,I130957,I131513,I1003386,I131539,I131547,I131564,I1003404,I1003398,I131581,I1003377,I131607,I1003395,I131624,I131632,I1003380,I131649,I131481,I131680,I131697,I131493,I1003392,I131737,I131502,I131759,I1003401,I1003389,I131776,I1003383,I131802,I131819,I131505,I131841,I131490,I131872,I131889,I131906,I131923,I131499,I131954,I131487,I131496,I131484,I132040,I854806,I132066,I132074,I132091,I854803,I854818,I132108,I854800,I132134,I854797,I132151,I132159,I132176,I132008,I132207,I132224,I132020,I132264,I132029,I132286,I854812,I132303,I854815,I132329,I132346,I132032,I132368,I132017,I132399,I854809,I132416,I132433,I132450,I132026,I132481,I132014,I132023,I132011,I132567,I613916,I132593,I132601,I132618,I613928,I613913,I132635,I613907,I132661,I613922,I132678,I132686,I613910,I132703,I132535,I132734,I132751,I132547,I613919,I132791,I132556,I132813,I613925,I613931,I132830,I132856,I132873,I132559,I132895,I132544,I132926,I132943,I132960,I132977,I132553,I133008,I132541,I132550,I132538,I133094,I867981,I133120,I133128,I133145,I867978,I867993,I133162,I867975,I133188,I867972,I133205,I133213,I133230,I133062,I133261,I133278,I133074,I133318,I133083,I133340,I867987,I133357,I867990,I133383,I133400,I133086,I133422,I133071,I133453,I867984,I133470,I133487,I133504,I133080,I133535,I133068,I133077,I133065,I133621,I311742,I133647,I133655,I133672,I311724,I311739,I133689,I311715,I133715,I311718,I133732,I133740,I311733,I133757,I133589,I133788,I133805,I133601,I311736,I133845,I133610,I133867,I311727,I133884,I311721,I133910,I133927,I133613,I133949,I133598,I133980,I311730,I133997,I134014,I134031,I133607,I134062,I133595,I133604,I133592,I134148,I682123,I134174,I134182,I134199,I682114,I682132,I134216,I682111,I134242,I134259,I134267,I682117,I134284,I134116,I134315,I134332,I134128,I134372,I134137,I134394,I682129,I682120,I134411,I682135,I134437,I134454,I134140,I134476,I134125,I134507,I682126,I134524,I134541,I134558,I134134,I134589,I134122,I134131,I134119,I134675,I1395205,I134701,I134709,I134726,I1395199,I1395220,I134743,I1395196,I134769,I1395217,I134786,I134794,I1395214,I134811,I134643,I134842,I134859,I134655,I1395202,I134899,I134664,I134921,I1395211,I1395208,I134938,I1395193,I134964,I134981,I134667,I135003,I134652,I135034,I135051,I135068,I135085,I134661,I135116,I134649,I134658,I134646,I135202,I1129727,I135228,I135236,I135253,I1129742,I1129721,I135270,I1129724,I135296,I1129745,I135313,I135321,I135338,I135170,I135369,I135386,I135182,I135426,I135191,I135448,I1129733,I1129730,I135465,I1129736,I135491,I135508,I135194,I135530,I135179,I135561,I1129739,I135578,I135595,I135612,I135188,I135643,I135176,I135185,I135173,I135729,I308580,I135755,I135763,I135780,I308562,I308577,I135797,I308553,I135823,I308556,I135840,I135848,I308571,I135865,I135697,I135896,I135913,I135709,I308574,I135953,I135718,I135975,I308565,I135992,I308559,I136018,I136035,I135721,I136057,I135706,I136088,I308568,I136105,I136122,I136139,I135715,I136170,I135703,I135712,I135700,I136256,I1233767,I136282,I136290,I136307,I1233782,I1233761,I136324,I1233764,I136350,I1233785,I136367,I136375,I136392,I136224,I136423,I136440,I136236,I136480,I136245,I136502,I1233773,I1233770,I136519,I1233776,I136545,I136562,I136248,I136584,I136233,I136615,I1233779,I136632,I136649,I136666,I136242,I136697,I136230,I136239,I136227,I136783,I136809,I136817,I136834,I136851,I136877,I136894,I136902,I136919,I136950,I136967,I137007,I137029,I137046,I137072,I137089,I137111,I137142,I137159,I137176,I137193,I137224,I137310,I321755,I137336,I137344,I137361,I321737,I321752,I137378,I321728,I137404,I321731,I137421,I137429,I321746,I137446,I137278,I137477,I137494,I137290,I321749,I137534,I137299,I137556,I321740,I137573,I321734,I137599,I137616,I137302,I137638,I137287,I137669,I321743,I137686,I137703,I137720,I137296,I137751,I137284,I137293,I137281,I137837,I137863,I137871,I137888,I137905,I137931,I137948,I137956,I137973,I137805,I138004,I138021,I137817,I138061,I137826,I138083,I138100,I138126,I138143,I137829,I138165,I137814,I138196,I138213,I138230,I138247,I137823,I138278,I137811,I137820,I137808,I138364,I492596,I138390,I138398,I138415,I492590,I492581,I138432,I492602,I138458,I492584,I138475,I138483,I492578,I138500,I138531,I138548,I138588,I138610,I492605,I492587,I138627,I492593,I138653,I138670,I138692,I138723,I492599,I138740,I138757,I138774,I138805,I138891,I292243,I138917,I138925,I138942,I292225,I292240,I138959,I292216,I138985,I292219,I139002,I139010,I292234,I139027,I138859,I139058,I139075,I138871,I292237,I139115,I138880,I139137,I292228,I139154,I292222,I139180,I139197,I138883,I139219,I138868,I139250,I292231,I139267,I139284,I139301,I138877,I139332,I138865,I138874,I138862,I139418,I580392,I139444,I139452,I139469,I580404,I580389,I139486,I580383,I139512,I580398,I139529,I139537,I580386,I139554,I139386,I139585,I139602,I139398,I580395,I139642,I139407,I139664,I580401,I580407,I139681,I139707,I139724,I139410,I139746,I139395,I139777,I139794,I139811,I139828,I139404,I139859,I139392,I139401,I139389,I139945,I668251,I139971,I139979,I139996,I668242,I668260,I140013,I668239,I140039,I140056,I140064,I668245,I140081,I139913,I140112,I140129,I139925,I140169,I139934,I140191,I668257,I668248,I140208,I668263,I140234,I140251,I139937,I140273,I139922,I140304,I668254,I140321,I140338,I140355,I139931,I140386,I139919,I139928,I139916,I140472,I952998,I140498,I140506,I140523,I953016,I953010,I140540,I952989,I140566,I953007,I140583,I140591,I952992,I140608,I140440,I140639,I140656,I140452,I953004,I140696,I140461,I140718,I953013,I953001,I140735,I952995,I140761,I140778,I140464,I140800,I140449,I140831,I140848,I140865,I140882,I140458,I140913,I140446,I140455,I140443,I140999,I685591,I141025,I141033,I141050,I685582,I685600,I141067,I685579,I141093,I141110,I141118,I685585,I141135,I140967,I141166,I141183,I140979,I141223,I140988,I141245,I685597,I685588,I141262,I685603,I141288,I141305,I140991,I141327,I140976,I141358,I685594,I141375,I141392,I141409,I140985,I141440,I140973,I140982,I140970,I141526,I1053955,I141552,I141560,I141577,I1053952,I1053958,I141594,I141620,I141637,I141645,I141662,I141494,I141693,I141710,I141506,I1053961,I141750,I141515,I141772,I1053964,I1053973,I141789,I1053967,I141815,I141832,I141518,I141854,I141503,I141885,I1053970,I141902,I141919,I141936,I141512,I141967,I141500,I141509,I141497,I142053,I1070785,I142079,I142087,I142104,I1070782,I1070788,I142121,I142147,I142164,I142172,I142189,I142021,I142220,I142237,I142033,I1070791,I142277,I142042,I142299,I1070794,I1070803,I142316,I1070797,I142342,I142359,I142045,I142381,I142030,I142412,I1070800,I142429,I142446,I142463,I142039,I142494,I142027,I142036,I142024,I142580,I605824,I142606,I142614,I142631,I605836,I605821,I142648,I605815,I142674,I605830,I142691,I142699,I605818,I142716,I142548,I142747,I142764,I142560,I605827,I142804,I142569,I142826,I605833,I605839,I142843,I142869,I142886,I142572,I142908,I142557,I142939,I142956,I142973,I142990,I142566,I143021,I142554,I142563,I142551,I143107,I1263823,I143133,I143141,I143158,I1263817,I1263838,I143175,I1263829,I143201,I1263820,I143218,I143226,I1263832,I143243,I143075,I143274,I143291,I143087,I143331,I143096,I143353,I1263841,I1263826,I143370,I143396,I143413,I143099,I143435,I143084,I143466,I1263835,I143483,I143500,I143517,I143093,I143548,I143081,I143090,I143078,I143634,I450708,I143660,I143668,I143685,I450702,I450693,I143702,I450714,I143728,I450696,I143745,I143753,I450690,I143770,I143602,I143801,I143818,I143614,I143858,I143623,I143880,I450717,I450699,I143897,I450705,I143923,I143940,I143626,I143962,I143611,I143993,I450711,I144010,I144027,I144044,I143620,I144075,I143608,I143617,I143605,I144161,I383414,I144187,I144195,I144212,I383396,I383411,I144229,I383387,I144255,I383390,I144272,I144280,I383405,I144297,I144129,I144328,I144345,I144141,I383408,I144385,I144150,I144407,I383399,I144424,I383393,I144450,I144467,I144153,I144489,I144138,I144520,I383402,I144537,I144554,I144571,I144147,I144602,I144135,I144144,I144132,I144688,I306999,I144714,I144722,I144739,I306981,I306996,I144756,I306972,I144782,I306975,I144799,I144807,I306990,I144824,I144656,I144855,I144872,I144668,I306993,I144912,I144677,I144934,I306984,I144951,I306978,I144977,I144994,I144680,I145016,I144665,I145047,I306987,I145064,I145081,I145098,I144674,I145129,I144662,I144671,I144659,I145215,I1294710,I145241,I145249,I145266,I1294713,I1294707,I145283,I1294704,I145309,I1294689,I145326,I145334,I1294698,I145351,I145183,I145382,I145399,I145195,I145439,I145204,I145461,I1294692,I1294695,I145478,I1294701,I145504,I145521,I145207,I145543,I145192,I145574,I145591,I145608,I145625,I145201,I145656,I145189,I145198,I145186,I145742,I353375,I145768,I145776,I145793,I353357,I353372,I145810,I353348,I145836,I353351,I145853,I145861,I353366,I145878,I145710,I145909,I145926,I145722,I353369,I145966,I145731,I145988,I353360,I146005,I353354,I146031,I146048,I145734,I146070,I145719,I146101,I353363,I146118,I146135,I146152,I145728,I146183,I145716,I145725,I145713,I146269,I732409,I146295,I146303,I146320,I732400,I732418,I146337,I732397,I146363,I146380,I146388,I732403,I146405,I146237,I146436,I146453,I146249,I146493,I146258,I146515,I732415,I732406,I146532,I732421,I146558,I146575,I146261,I146597,I146246,I146628,I732412,I146645,I146662,I146679,I146255,I146710,I146243,I146252,I146240,I146796,I334930,I146822,I146830,I146847,I334912,I334927,I146864,I334903,I146890,I334906,I146907,I146915,I334921,I146932,I146764,I146963,I146980,I146776,I334924,I147020,I146785,I147042,I334915,I147059,I334909,I147085,I147102,I146788,I147124,I146773,I147155,I334918,I147172,I147189,I147206,I146782,I147237,I146770,I146779,I146767,I147323,I207755,I147349,I147357,I147374,I207749,I207743,I147391,I207764,I147417,I207761,I147434,I147442,I207758,I147459,I147291,I147490,I147507,I147303,I147547,I147312,I147569,I207746,I147586,I207767,I147612,I147629,I147315,I147651,I147300,I147682,I207752,I147699,I147716,I147733,I147309,I147764,I147297,I147306,I147294,I147850,I316485,I147876,I147884,I147901,I316467,I316482,I147918,I316458,I147944,I316461,I147961,I147969,I316476,I147986,I147818,I148017,I148034,I147830,I316479,I148074,I147839,I148096,I316470,I148113,I316464,I148139,I148156,I147842,I148178,I147827,I148209,I316473,I148226,I148243,I148260,I147836,I148291,I147824,I147833,I147821,I148377,I702931,I148403,I148411,I148428,I702922,I702940,I148445,I702919,I148471,I148488,I148496,I702925,I148513,I148345,I148544,I148561,I148357,I148601,I148366,I148623,I702937,I702928,I148640,I702943,I148666,I148683,I148369,I148705,I148354,I148736,I702934,I148753,I148770,I148787,I148363,I148818,I148351,I148360,I148348,I148904,I694261,I148930,I148938,I148955,I694252,I694270,I148972,I694249,I148998,I149015,I149023,I694255,I149040,I148872,I149071,I149088,I148884,I149128,I148893,I149150,I694267,I694258,I149167,I694273,I149193,I149210,I148896,I149232,I148881,I149263,I694264,I149280,I149297,I149314,I148890,I149345,I148878,I148887,I148875,I149431,I1239547,I149457,I149465,I149482,I1239562,I1239541,I149499,I1239544,I149525,I1239565,I149542,I149550,I149567,I149399,I149598,I149615,I149411,I149655,I149420,I149677,I1239553,I1239550,I149694,I1239556,I149720,I149737,I149423,I149759,I149408,I149790,I1239559,I149807,I149824,I149841,I149417,I149872,I149405,I149414,I149402,I149958,I1057882,I149984,I149992,I150009,I1057879,I1057885,I150026,I150052,I150069,I150077,I150094,I149926,I150125,I150142,I149938,I1057888,I150182,I149947,I150204,I1057891,I1057900,I150221,I1057894,I150247,I150264,I149950,I150286,I149935,I150317,I1057897,I150334,I150351,I150368,I149944,I150399,I149932,I149941,I149929,I150485,I843739,I150511,I150519,I150536,I843736,I843751,I150553,I843733,I150579,I843730,I150596,I150604,I150621,I150453,I150652,I150669,I150465,I150709,I150474,I150731,I843745,I150748,I843748,I150774,I150791,I150477,I150813,I150462,I150844,I843742,I150861,I150878,I150895,I150471,I150926,I150459,I150468,I150456,I151012,I381833,I151038,I151046,I151063,I381815,I381830,I151080,I381806,I151106,I381809,I151123,I151131,I381824,I151148,I150980,I151179,I151196,I150992,I381827,I151236,I151001,I151258,I381818,I151275,I381812,I151301,I151318,I151004,I151340,I150989,I151371,I381821,I151388,I151405,I151422,I150998,I151453,I150986,I150995,I150983,I151539,I1052272,I151565,I151573,I151590,I1052269,I1052275,I151607,I151633,I151650,I151658,I151675,I151507,I151706,I151723,I151519,I1052278,I151763,I151528,I151785,I1052281,I1052290,I151802,I1052284,I151828,I151845,I151531,I151867,I151516,I151898,I1052287,I151915,I151932,I151949,I151525,I151980,I151513,I151522,I151510,I152066,I201210,I152092,I152100,I152117,I201204,I201198,I152134,I201219,I152160,I201216,I152177,I152185,I201213,I152202,I152034,I152233,I152250,I152046,I152290,I152055,I152312,I201201,I152329,I201222,I152355,I152372,I152058,I152394,I152043,I152425,I201207,I152442,I152459,I152476,I152052,I152507,I152040,I152049,I152037,I152593,I1206601,I152619,I152627,I152644,I1206616,I1206595,I152661,I1206598,I152687,I1206619,I152704,I152712,I152729,I152561,I152760,I152777,I152573,I152817,I152582,I152839,I1206607,I1206604,I152856,I1206610,I152882,I152899,I152585,I152921,I152570,I152952,I1206613,I152969,I152986,I153003,I152579,I153034,I152567,I152576,I152564,I153120,I711601,I153146,I153154,I153171,I711592,I711610,I153188,I711589,I153214,I153231,I153239,I711595,I153256,I153088,I153287,I153304,I153100,I153344,I153109,I153366,I711607,I711598,I153383,I711613,I153409,I153426,I153112,I153448,I153097,I153479,I711604,I153496,I153513,I153530,I153106,I153561,I153094,I153103,I153091,I153647,I272610,I153673,I153681,I153698,I272604,I272598,I153715,I272619,I153741,I272616,I153758,I153766,I272613,I153783,I153615,I153814,I153831,I153627,I153871,I153636,I153893,I272601,I153910,I272622,I153936,I153953,I153639,I153975,I153624,I154006,I272607,I154023,I154040,I154057,I153633,I154088,I153621,I153630,I153618,I154174,I327552,I154200,I154208,I154225,I327534,I327549,I154242,I327525,I154268,I327528,I154285,I154293,I327543,I154310,I154142,I154341,I154358,I154154,I327546,I154398,I154163,I154420,I327537,I154437,I327531,I154463,I154480,I154166,I154502,I154151,I154533,I327540,I154550,I154567,I154584,I154160,I154615,I154148,I154157,I154145,I154701,I379198,I154727,I154735,I154752,I379180,I379195,I154769,I379171,I154795,I379174,I154812,I154820,I379189,I154837,I154669,I154868,I154885,I154681,I379192,I154925,I154690,I154947,I379183,I154964,I379177,I154990,I155007,I154693,I155029,I154678,I155060,I379186,I155077,I155094,I155111,I154687,I155142,I154675,I154684,I154672,I155228,I1360100,I155254,I155262,I155279,I1360094,I1360115,I155296,I1360091,I155322,I1360112,I155339,I155347,I1360109,I155364,I155196,I155395,I155412,I155208,I1360097,I155452,I155217,I155474,I1360106,I1360103,I155491,I1360088,I155517,I155534,I155220,I155556,I155205,I155587,I155604,I155621,I155638,I155214,I155669,I155202,I155211,I155199,I155755,I1130305,I155781,I155789,I155806,I1130320,I1130299,I155823,I1130302,I155849,I1130323,I155866,I155874,I155891,I155723,I155922,I155939,I155735,I155979,I155744,I156001,I1130311,I1130308,I156018,I1130314,I156044,I156061,I155747,I156083,I155732,I156114,I1130317,I156131,I156148,I156165,I155741,I156196,I155729,I155738,I155726,I156282,I985298,I156308,I156316,I156333,I985316,I985310,I156350,I985289,I156376,I985307,I156393,I156401,I985292,I156418,I156250,I156449,I156466,I156262,I985304,I156506,I156271,I156528,I985313,I985301,I156545,I985295,I156571,I156588,I156274,I156610,I156259,I156641,I156658,I156675,I156692,I156268,I156723,I156256,I156265,I156253,I156809,I1089298,I156835,I156843,I156860,I1089295,I1089301,I156877,I156903,I156920,I156928,I156945,I156777,I156976,I156993,I156789,I1089304,I157033,I156798,I157055,I1089307,I1089316,I157072,I1089310,I157098,I157115,I156801,I157137,I156786,I157168,I1089313,I157185,I157202,I157219,I156795,I157250,I156783,I156792,I156780,I157336,I1293554,I157362,I157370,I157387,I1293557,I1293551,I157404,I1293548,I157430,I1293533,I157447,I157455,I1293542,I157472,I157304,I157503,I157520,I157316,I157560,I157325,I157582,I1293536,I1293539,I157599,I1293545,I157625,I157642,I157328,I157664,I157313,I157695,I157712,I157729,I157746,I157322,I157777,I157310,I157319,I157307,I157863,I228580,I157889,I157897,I157914,I228574,I228568,I157931,I228589,I157957,I228586,I157974,I157982,I228583,I157999,I157831,I158030,I158047,I157843,I158087,I157852,I158109,I228571,I158126,I228592,I158152,I158169,I157855,I158191,I157840,I158222,I228577,I158239,I158256,I158273,I157849,I158304,I157837,I157846,I157834,I158393,I1264364,I158419,I158427,I1264376,I158453,I158461,I1264382,I158478,I1264361,I158495,I158370,I158526,I1264379,I158364,I158557,I158574,I158591,I1264367,I158608,I158625,I158642,I158379,I158376,I158382,I158701,I158718,I158735,I1264385,I1264373,I158761,I158361,I158792,I158800,I1264370,I158385,I158831,I158848,I158865,I158367,I158896,I158913,I158358,I158373,I158988,I159014,I159022,I159048,I159056,I159073,I159090,I158965,I159121,I158959,I159152,I159169,I159186,I159203,I159220,I159237,I158974,I158971,I158977,I159296,I159313,I159330,I159356,I158956,I159387,I159395,I158980,I159426,I159443,I159460,I158962,I159491,I159508,I158953,I158968,I159583,I394990,I159609,I159617,I394987,I159643,I159651,I394984,I159668,I394996,I159685,I159560,I159716,I395005,I159554,I159747,I395002,I159764,I159781,I394981,I159798,I159815,I159832,I159569,I159566,I159572,I159891,I159908,I159925,I394993,I395008,I159951,I159551,I159982,I159990,I394999,I159575,I160021,I160038,I160055,I159557,I160086,I160103,I159548,I159563,I160178,I520890,I160204,I160212,I520884,I160238,I160246,I520881,I160263,I520872,I160280,I160155,I160311,I520875,I160149,I160342,I520878,I160359,I160376,I520866,I520893,I160393,I160410,I160427,I160164,I160161,I160167,I160486,I160503,I160520,I520869,I160546,I160146,I160577,I160585,I520887,I160170,I160616,I160633,I160650,I160152,I160681,I160698,I160143,I160158,I160773,I160799,I160807,I160833,I160841,I160858,I160875,I160750,I160906,I160744,I160937,I160954,I160971,I160988,I161005,I161022,I160759,I160756,I160762,I161081,I161098,I161115,I161141,I160741,I161172,I161180,I160765,I161211,I161228,I161245,I160747,I161276,I161293,I160738,I160753,I161368,I1277964,I161394,I161402,I1277976,I161428,I161436,I1277982,I161453,I1277961,I161470,I161345,I161501,I1277979,I161339,I161532,I161549,I161566,I1277967,I161583,I161600,I161617,I161354,I161351,I161357,I161676,I161693,I161710,I1277985,I1277973,I161736,I161336,I161767,I161775,I1277970,I161360,I161806,I161823,I161840,I161342,I161871,I161888,I161333,I161348,I161963,I350195,I161989,I161997,I350192,I162023,I162031,I350189,I162048,I350201,I162065,I161940,I162096,I350210,I161934,I162127,I350207,I162144,I162161,I350186,I162178,I162195,I162212,I161949,I161946,I161952,I162271,I162288,I162305,I350198,I350213,I162331,I161931,I162362,I162370,I350204,I161955,I162401,I162418,I162435,I161937,I162466,I162483,I161928,I161943,I162558,I411327,I162584,I162592,I411324,I162618,I162626,I411321,I162643,I411333,I162660,I162535,I162691,I411342,I162529,I162722,I411339,I162739,I162756,I411318,I162773,I162790,I162807,I162544,I162541,I162547,I162866,I162883,I162900,I411330,I411345,I162926,I162526,I162957,I162965,I411336,I162550,I162996,I163013,I163030,I162532,I163061,I163078,I162523,I162538,I163153,I776903,I163179,I163187,I776924,I163213,I163221,I163238,I776915,I163255,I163130,I163286,I776912,I163124,I163317,I776921,I163334,I163351,I776906,I163368,I163385,I163402,I163139,I163136,I163142,I163461,I163478,I163495,I776927,I776909,I163521,I163121,I163552,I163560,I776918,I163145,I163591,I163608,I163625,I163127,I163656,I163673,I163118,I163133,I163748,I1130880,I163774,I163782,I1130877,I163808,I163816,I1130886,I163833,I163850,I163725,I163881,I1130889,I163719,I163912,I1130883,I163929,I163946,I1130898,I163963,I163980,I163997,I163734,I163731,I163737,I164056,I164073,I164090,I1130901,I1130895,I164116,I163716,I164147,I164155,I1130892,I163740,I164186,I164203,I164220,I163722,I164251,I164268,I163713,I163728,I164343,I724883,I164369,I164377,I724904,I164403,I164411,I164428,I724895,I164445,I164320,I164476,I724892,I164314,I164507,I724901,I164524,I164541,I724886,I164558,I164575,I164592,I164329,I164326,I164332,I164651,I164668,I164685,I724907,I724889,I164711,I164311,I164742,I164750,I724898,I164335,I164781,I164798,I164815,I164317,I164846,I164863,I164308,I164323,I164938,I1027931,I164964,I164972,I1027952,I164998,I165006,I1027934,I165023,I1027925,I165040,I164915,I165071,I1027937,I164909,I165102,I1027928,I165119,I165136,I1027946,I1027949,I165153,I165170,I165187,I164924,I164921,I164927,I165246,I165263,I165280,I1027940,I1027943,I165306,I164906,I165337,I165345,I164930,I165376,I165393,I165410,I164912,I165441,I165458,I164903,I164918,I165530,I1096775,I165556,I165573,I165522,I165595,I165621,I165629,I165646,I1096778,I165663,I1096790,I165680,I165697,I1096796,I165714,I1096787,I165731,I1096793,I165748,I165498,I165779,I165796,I165813,I165830,I165510,I165504,I165875,I1096784,I165519,I165513,I165920,I165937,I1096781,I165954,I1096799,I165971,I165997,I166005,I165507,I165501,I166059,I166067,I165516,I166125,I1250235,I166151,I166168,I166117,I166190,I1250220,I166216,I166224,I166241,I1250238,I166258,I166275,I166292,I1250241,I166309,I1250232,I166326,I1250229,I166343,I166093,I166374,I166391,I166408,I166425,I166105,I166099,I166470,I1250226,I166114,I166108,I166515,I166532,I1250217,I166549,I1250223,I166566,I166592,I166600,I166102,I166096,I166654,I166662,I166111,I166720,I166746,I166763,I166785,I166811,I166819,I166836,I166853,I166870,I166887,I166904,I166921,I166938,I166969,I166986,I167003,I167020,I167065,I167110,I167127,I167144,I167161,I167187,I167195,I167249,I167257,I167315,I167341,I167358,I167307,I167380,I167406,I167414,I167431,I167448,I167465,I167482,I167499,I167516,I167533,I167283,I167564,I167581,I167598,I167615,I167295,I167289,I167660,I167304,I167298,I167705,I167722,I167739,I167756,I167782,I167790,I167292,I167286,I167844,I167852,I167301,I167910,I167936,I167953,I167902,I167975,I168001,I168009,I168026,I168043,I168060,I168077,I168094,I168111,I168128,I167878,I168159,I168176,I168193,I168210,I167890,I167884,I168255,I167899,I167893,I168300,I168317,I168334,I168351,I168377,I168385,I167887,I167881,I168439,I168447,I167896,I168505,I1082005,I168531,I168548,I168570,I1082014,I168596,I168604,I168621,I1082008,I168638,I1082002,I168655,I168672,I1082017,I168689,I168706,I1082011,I168723,I168754,I168771,I168788,I168805,I168850,I168895,I168912,I1082023,I168929,I1082020,I168946,I168972,I168980,I169034,I169042,I169100,I1056199,I169126,I169143,I169092,I169165,I1056208,I169191,I169199,I169216,I1056202,I169233,I1056196,I169250,I169267,I1056211,I169284,I169301,I1056205,I169318,I169068,I169349,I169366,I169383,I169400,I169080,I169074,I169445,I169089,I169083,I169490,I169507,I1056217,I169524,I1056214,I169541,I169567,I169575,I169077,I169071,I169629,I169637,I169086,I169695,I782695,I169721,I169738,I169687,I169760,I782692,I169786,I169794,I169811,I782698,I169828,I782683,I169845,I169862,I782686,I169879,I782707,I169896,I782704,I169913,I169663,I169944,I169961,I169978,I169995,I169675,I169669,I170040,I169684,I169678,I170085,I170102,I782689,I170119,I782701,I170136,I170162,I170170,I169672,I169666,I170224,I170232,I169681,I170290,I1126831,I170316,I170333,I170282,I170355,I170381,I170389,I170406,I1126834,I170423,I1126846,I170440,I170457,I1126852,I170474,I1126843,I170491,I1126849,I170508,I170258,I170539,I170556,I170573,I170590,I170270,I170264,I170635,I1126840,I170279,I170273,I170680,I170697,I1126837,I170714,I1126855,I170731,I170757,I170765,I170267,I170261,I170819,I170827,I170276,I170885,I170911,I170928,I170877,I170950,I170976,I170984,I171001,I171018,I171035,I171052,I171069,I171086,I171103,I170853,I171134,I171151,I171168,I171185,I170865,I170859,I171230,I170874,I170868,I171275,I171292,I171309,I171326,I171352,I171360,I170862,I170856,I171414,I171422,I170871,I171480,I1250779,I171506,I171523,I171472,I171545,I1250764,I171571,I171579,I171596,I1250782,I171613,I171630,I171647,I1250785,I171664,I1250776,I171681,I1250773,I171698,I171448,I171729,I171746,I171763,I171780,I171460,I171454,I171825,I1250770,I171469,I171463,I171870,I171887,I1250761,I171904,I1250767,I171921,I171947,I171955,I171457,I171451,I172009,I172017,I171466,I172075,I1234917,I172101,I172118,I172067,I172140,I172166,I172174,I172191,I1234920,I172208,I1234932,I172225,I172242,I1234938,I172259,I1234929,I172276,I1234935,I172293,I172043,I172324,I172341,I172358,I172375,I172055,I172049,I172420,I1234926,I172064,I172058,I172465,I172482,I1234923,I172499,I1234941,I172516,I172542,I172550,I172052,I172046,I172604,I172612,I172061,I172670,I1313188,I172696,I172713,I172662,I172735,I1313200,I172761,I172769,I172786,I1313194,I172803,I1313206,I172820,I172837,I1313191,I172854,I1313203,I172871,I1313185,I172888,I172638,I172919,I172936,I172953,I172970,I172650,I172644,I173015,I1313197,I172659,I172653,I173060,I173077,I173094,I173111,I1313209,I173137,I173145,I172647,I172641,I173199,I173207,I172656,I173265,I477914,I173291,I173308,I173257,I173330,I477902,I173356,I173364,I173381,I477911,I173398,I477908,I173415,I173432,I477899,I173449,I477905,I173466,I477890,I173483,I173233,I173514,I173531,I173548,I173565,I173245,I173239,I173610,I173254,I173248,I173655,I173672,I477896,I173689,I477893,I173706,I477917,I173732,I173740,I173242,I173236,I173794,I173802,I173251,I173860,I173886,I173903,I173852,I173925,I173951,I173959,I173976,I173993,I174010,I174027,I174044,I174061,I174078,I173828,I174109,I174126,I174143,I174160,I173840,I173834,I174205,I173849,I173843,I174250,I174267,I174284,I174301,I174327,I174335,I173837,I173831,I174389,I174397,I173846,I174455,I370212,I174481,I174498,I174520,I370227,I174546,I174554,I174571,I370224,I174588,I174605,I174622,I370221,I174639,I370236,I174656,I370233,I174673,I174704,I174721,I174738,I174755,I174800,I370230,I174845,I174862,I370218,I174879,I370239,I174896,I370215,I174922,I174930,I174984,I174992,I175050,I175076,I175093,I175115,I175141,I175149,I175166,I175183,I175200,I175217,I175234,I175251,I175268,I175299,I175316,I175333,I175350,I175395,I175440,I175457,I175474,I175491,I175517,I175525,I175579,I175587,I175645,I951066,I175671,I175688,I175637,I175710,I951075,I175736,I175744,I175761,I951063,I175778,I951054,I175795,I175812,I951060,I175829,I951078,I175846,I951051,I175863,I175613,I175894,I175911,I175928,I175945,I175625,I175619,I175990,I951057,I175634,I175628,I176035,I176052,I951069,I176069,I176086,I951072,I176112,I176120,I175622,I175616,I176174,I176182,I175631,I176240,I661893,I176266,I176283,I176305,I661890,I176331,I176339,I176356,I661896,I176373,I661881,I176390,I176407,I661884,I176424,I661905,I176441,I661902,I176458,I176489,I176506,I176523,I176540,I176585,I176630,I176647,I661887,I176664,I661899,I176681,I176707,I176715,I176769,I176777,I176835,I1066858,I176861,I176878,I176827,I176900,I1066867,I176926,I176934,I176951,I1066861,I176968,I1066855,I176985,I177002,I1066870,I177019,I177036,I1066864,I177053,I176803,I177084,I177101,I177118,I177135,I176815,I176809,I177180,I176824,I176818,I177225,I177242,I1066876,I177259,I1066873,I177276,I177302,I177310,I176812,I176806,I177364,I177372,I176821,I177430,I896436,I177456,I177473,I177422,I177495,I896430,I177521,I177529,I177546,I896448,I177563,I177580,I177597,I177614,I896442,I177631,I896433,I177648,I177398,I177679,I177696,I177713,I177730,I177410,I177404,I177775,I896445,I177419,I177413,I177820,I177837,I896451,I177854,I177871,I896439,I177897,I177905,I177407,I177401,I177959,I177967,I177416,I178025,I1107757,I178051,I178068,I178017,I178090,I178116,I178124,I178141,I1107760,I178158,I1107772,I178175,I178192,I1107778,I178209,I1107769,I178226,I1107775,I178243,I177993,I178274,I178291,I178308,I178325,I178005,I177999,I178370,I1107766,I178014,I178008,I178415,I178432,I1107763,I178449,I1107781,I178466,I178492,I178500,I178002,I177996,I178554,I178562,I178011,I178620,I714491,I178646,I178663,I178612,I178685,I714488,I178711,I178719,I178736,I714494,I178753,I714479,I178770,I178787,I714482,I178804,I714503,I178821,I714500,I178838,I178588,I178869,I178886,I178903,I178920,I178600,I178594,I178965,I178609,I178603,I179010,I179027,I714485,I179044,I714497,I179061,I179087,I179095,I178597,I178591,I179149,I179157,I178606,I179215,I414480,I179241,I179258,I179207,I179280,I414495,I179306,I179314,I179331,I414492,I179348,I179365,I179382,I414489,I179399,I414504,I179416,I414501,I179433,I179183,I179464,I179481,I179498,I179515,I179195,I179189,I179560,I414498,I179204,I179198,I179605,I179622,I414486,I179639,I414507,I179656,I414483,I179682,I179690,I179192,I179186,I179744,I179752,I179201,I179810,I760153,I179836,I179853,I179802,I179875,I760150,I179901,I179909,I179926,I760156,I179943,I760141,I179960,I179977,I760144,I179994,I760165,I180011,I760162,I180028,I179778,I180059,I180076,I180093,I180110,I179790,I179784,I180155,I179799,I179793,I180200,I180217,I760147,I180234,I760159,I180251,I180277,I180285,I179787,I179781,I180339,I180347,I179796,I180405,I180431,I180448,I180397,I180470,I180496,I180504,I180521,I180538,I180555,I180572,I180589,I180606,I180623,I180373,I180654,I180671,I180688,I180705,I180385,I180379,I180750,I180394,I180388,I180795,I180812,I180829,I180846,I180872,I180880,I180382,I180376,I180934,I180942,I180391,I181000,I328579,I181026,I181043,I180992,I181065,I328594,I181091,I181099,I181116,I328591,I181133,I181150,I181167,I328588,I181184,I328603,I181201,I328600,I181218,I180968,I181249,I181266,I181283,I181300,I180980,I180974,I181345,I328597,I180989,I180983,I181390,I181407,I328585,I181424,I328606,I181441,I328582,I181467,I181475,I180977,I180971,I181529,I181537,I180986,I181595,I735877,I181621,I181638,I181587,I181660,I735874,I181686,I181694,I181711,I735880,I181728,I735865,I181745,I181762,I735868,I181779,I735889,I181796,I735886,I181813,I181563,I181844,I181861,I181878,I181895,I181575,I181569,I181940,I181584,I181578,I181985,I182002,I735871,I182019,I735883,I182036,I182062,I182070,I181572,I181566,I182124,I182132,I181581,I182190,I182216,I182233,I182182,I182255,I182281,I182289,I182306,I182323,I182340,I182357,I182374,I182391,I182408,I182158,I182439,I182456,I182473,I182490,I182170,I182164,I182535,I182179,I182173,I182580,I182597,I182614,I182631,I182657,I182665,I182167,I182161,I182719,I182727,I182176,I182785,I1297004,I182811,I182828,I182777,I182850,I1297016,I182876,I182884,I182901,I1297010,I182918,I1297022,I182935,I182952,I1297007,I182969,I1297019,I182986,I1297001,I183003,I182753,I183034,I183051,I183068,I183085,I182765,I182759,I183130,I1297013,I182774,I182768,I183175,I183192,I183209,I183226,I1297025,I183252,I183260,I182762,I182756,I183314,I183322,I182771,I183380,I690215,I183406,I183423,I183372,I183445,I690212,I183471,I183479,I183496,I690218,I183513,I690203,I183530,I183547,I690206,I183564,I690227,I183581,I690224,I183598,I183348,I183629,I183646,I183663,I183680,I183360,I183354,I183725,I183369,I183363,I183770,I183787,I690209,I183804,I690221,I183821,I183847,I183855,I183357,I183351,I183909,I183917,I183366,I183975,I591380,I184001,I184018,I183967,I184040,I591371,I184066,I184074,I184091,I591389,I184108,I591386,I184125,I184142,I591365,I184159,I591368,I184176,I591377,I184193,I183943,I184224,I184241,I184258,I184275,I183955,I183949,I184320,I591383,I183964,I183958,I184365,I184382,I184399,I591374,I184416,I184442,I184450,I183952,I183946,I184504,I184512,I183961,I184570,I614500,I184596,I184613,I184562,I184635,I614491,I184661,I184669,I184686,I614509,I184703,I614506,I184720,I184737,I614485,I184754,I614488,I184771,I614497,I184788,I184538,I184819,I184836,I184853,I184870,I184550,I184544,I184915,I614503,I184559,I184553,I184960,I184977,I184994,I614494,I185011,I185037,I185045,I184547,I184541,I185099,I185107,I184556,I185165,I1257851,I185191,I185208,I185157,I185230,I1257836,I185256,I185264,I185281,I1257854,I185298,I185315,I185332,I1257857,I185349,I1257848,I185366,I1257845,I185383,I185133,I185414,I185431,I185448,I185465,I185145,I185139,I185510,I1257842,I185154,I185148,I185555,I185572,I1257833,I185589,I1257839,I185606,I185632,I185640,I185142,I185136,I185694,I185702,I185151,I185760,I1051150,I185786,I185803,I185752,I185825,I1051159,I185851,I185859,I185876,I1051153,I185893,I1051147,I185910,I185927,I1051162,I185944,I185961,I1051156,I185978,I185728,I186009,I186026,I186043,I186060,I185740,I185734,I186105,I185749,I185743,I186150,I186167,I1051168,I186184,I1051165,I186201,I186227,I186235,I185737,I185731,I186289,I186297,I185746,I186355,I485530,I186381,I186398,I186347,I186420,I485518,I186446,I186454,I186471,I485527,I186488,I485524,I186505,I186522,I485515,I186539,I485521,I186556,I485506,I186573,I186323,I186604,I186621,I186638,I186655,I186335,I186329,I186700,I186344,I186338,I186745,I186762,I485512,I186779,I485509,I186796,I485533,I186822,I186830,I186332,I186326,I186884,I186892,I186341,I186950,I593692,I186976,I186993,I186942,I187015,I593683,I187041,I187049,I187066,I593701,I187083,I593698,I187100,I187117,I593677,I187134,I593680,I187151,I593689,I187168,I186918,I187199,I187216,I187233,I187250,I186930,I186924,I187295,I593695,I186939,I186933,I187340,I187357,I187374,I593686,I187391,I187417,I187425,I186927,I186921,I187479,I187487,I186936,I187545,I578664,I187571,I187588,I187537,I187610,I578655,I187636,I187644,I187661,I578673,I187678,I578670,I187695,I187712,I578649,I187729,I578652,I187746,I578661,I187763,I187513,I187794,I187811,I187828,I187845,I187525,I187519,I187890,I578667,I187534,I187528,I187935,I187952,I187969,I578658,I187986,I188012,I188020,I187522,I187516,I188074,I188082,I187531,I188140,I1046028,I188166,I188183,I188132,I188205,I1046037,I188231,I188239,I188256,I1046025,I188273,I1046016,I188290,I188307,I1046022,I188324,I1046040,I188341,I1046013,I188358,I188108,I188389,I188406,I188423,I188440,I188120,I188114,I188485,I1046019,I188129,I188123,I188530,I188547,I1046031,I188564,I188581,I1046034,I188607,I188615,I188117,I188111,I188669,I188677,I188126,I188735,I767089,I188761,I188778,I188727,I188800,I767086,I188826,I188834,I188851,I767092,I188868,I767077,I188885,I188902,I767080,I188919,I767101,I188936,I767098,I188953,I188703,I188984,I189001,I189018,I189035,I188715,I188709,I189080,I188724,I188718,I189125,I189142,I767083,I189159,I767095,I189176,I189202,I189210,I188712,I188706,I189264,I189272,I188721,I189330,I1048345,I189356,I189373,I189322,I189395,I1048354,I189421,I189429,I189446,I1048348,I189463,I1048342,I189480,I189497,I1048357,I189514,I189531,I1048351,I189548,I189298,I189579,I189596,I189613,I189630,I189310,I189304,I189675,I189319,I189313,I189720,I189737,I1048363,I189754,I1048360,I189771,I189797,I189805,I189307,I189301,I189859,I189867,I189316,I189925,I671719,I189951,I189968,I189917,I189990,I671716,I190016,I190024,I190041,I671722,I190058,I671707,I190075,I190092,I671710,I190109,I671731,I190126,I671728,I190143,I189893,I190174,I190191,I190208,I190225,I189905,I189899,I190270,I189914,I189908,I190315,I190332,I671713,I190349,I671725,I190366,I190392,I190400,I189902,I189896,I190454,I190462,I189911,I190520,I634152,I190546,I190563,I190512,I190585,I634143,I190611,I190619,I190636,I634161,I190653,I634158,I190670,I190687,I634137,I190704,I634140,I190721,I634149,I190738,I190488,I190769,I190786,I190803,I190820,I190500,I190494,I190865,I634155,I190509,I190503,I190910,I190927,I190944,I634146,I190961,I190987,I190995,I190497,I190491,I191049,I191057,I190506,I191115,I1276347,I191141,I191158,I191107,I191180,I1276332,I191206,I191214,I191231,I1276350,I191248,I191265,I191282,I1276353,I191299,I1276344,I191316,I1276341,I191333,I191083,I191364,I191381,I191398,I191415,I191095,I191089,I191460,I1276338,I191104,I191098,I191505,I191522,I1276329,I191539,I1276335,I191556,I191582,I191590,I191092,I191086,I191644,I191652,I191101,I191710,I356510,I191736,I191753,I191702,I191775,I356525,I191801,I191809,I191826,I356522,I191843,I191860,I191877,I356519,I191894,I356534,I191911,I356531,I191928,I191678,I191959,I191976,I191993,I192010,I191690,I191684,I192055,I356528,I191699,I191693,I192100,I192117,I356516,I192134,I356537,I192151,I356513,I192177,I192185,I191687,I191681,I192239,I192247,I191696,I192305,I649180,I192331,I192348,I192297,I192370,I649171,I192396,I192404,I192421,I649189,I192438,I649186,I192455,I192472,I649165,I192489,I649168,I192506,I649177,I192523,I192273,I192554,I192571,I192588,I192605,I192285,I192279,I192650,I649183,I192294,I192288,I192695,I192712,I192729,I649174,I192746,I192772,I192780,I192282,I192276,I192834,I192842,I192291,I192900,I192926,I192943,I192892,I192965,I192991,I192999,I193016,I193033,I193050,I193067,I193084,I193101,I193118,I192868,I193149,I193166,I193183,I193200,I192880,I192874,I193245,I192889,I192883,I193290,I193307,I193324,I193341,I193367,I193375,I192877,I192871,I193429,I193437,I192886,I193495,I193521,I193538,I193487,I193560,I193586,I193594,I193611,I193628,I193645,I193662,I193679,I193696,I193713,I193463,I193744,I193761,I193778,I193795,I193475,I193469,I193840,I193484,I193478,I193885,I193902,I193919,I193936,I193962,I193970,I193472,I193466,I194024,I194032,I193481,I194090,I1122785,I194116,I194133,I194082,I194155,I194181,I194189,I194206,I1122788,I194223,I1122800,I194240,I194257,I1122806,I194274,I1122797,I194291,I1122803,I194308,I194058,I194339,I194356,I194373,I194390,I194070,I194064,I194435,I1122794,I194079,I194073,I194480,I194497,I1122791,I194514,I1122809,I194531,I194557,I194565,I194067,I194061,I194619,I194627,I194076,I194685,I661315,I194711,I194728,I194677,I194750,I661312,I194776,I194784,I194801,I661318,I194818,I661303,I194835,I194852,I661306,I194869,I661327,I194886,I661324,I194903,I194653,I194934,I194951,I194968,I194985,I194665,I194659,I195030,I194674,I194668,I195075,I195092,I661309,I195109,I661321,I195126,I195152,I195160,I194662,I194656,I195214,I195222,I194671,I195280,I675765,I195306,I195323,I195272,I195345,I675762,I195371,I195379,I195396,I675768,I195413,I675753,I195430,I195447,I675756,I195464,I675777,I195481,I675774,I195498,I195248,I195529,I195546,I195563,I195580,I195260,I195254,I195625,I195269,I195263,I195670,I195687,I675759,I195704,I675771,I195721,I195747,I195755,I195257,I195251,I195809,I195817,I195266,I195875,I435482,I195901,I195918,I195867,I195940,I435470,I195966,I195974,I195991,I435479,I196008,I435476,I196025,I196042,I435467,I196059,I435473,I196076,I435458,I196093,I195843,I196124,I196141,I196158,I196175,I195855,I195849,I196220,I195864,I195858,I196265,I196282,I435464,I196299,I435461,I196316,I435485,I196342,I196350,I195852,I195846,I196404,I196412,I195861,I196470,I865343,I196496,I196513,I196462,I196535,I865337,I196561,I196569,I196586,I865355,I196603,I196620,I196637,I196654,I865349,I196671,I865340,I196688,I196438,I196719,I196736,I196753,I196770,I196450,I196444,I196815,I865352,I196459,I196453,I196860,I196877,I865358,I196894,I196911,I865346,I196937,I196945,I196447,I196441,I196999,I197007,I196456,I197065,I1301050,I197091,I197108,I197057,I197130,I1301062,I197156,I197164,I197181,I1301056,I197198,I1301068,I197215,I197232,I1301053,I197249,I1301065,I197266,I1301047,I197283,I197033,I197314,I197331,I197348,I197365,I197045,I197039,I197410,I1301059,I197054,I197048,I197455,I197472,I197489,I197506,I1301071,I197532,I197540,I197042,I197036,I197594,I197602,I197051,I197660,I660159,I197686,I197703,I197652,I197725,I660156,I197751,I197759,I197776,I660162,I197793,I660147,I197810,I197827,I660150,I197844,I660171,I197861,I660168,I197878,I197628,I197909,I197926,I197943,I197960,I197640,I197634,I198005,I197649,I197643,I198050,I198067,I660153,I198084,I660165,I198101,I198127,I198135,I197637,I197631,I198189,I198197,I197646,I198255,I1129143,I198281,I198298,I198247,I198320,I198346,I198354,I198371,I1129146,I198388,I1129158,I198405,I198422,I1129164,I198439,I1129155,I198456,I1129161,I198473,I198223,I198504,I198521,I198538,I198555,I198235,I198229,I198600,I1129152,I198244,I198238,I198645,I198662,I1129149,I198679,I1129167,I198696,I198722,I198730,I198232,I198226,I198784,I198792,I198241,I198850,I1372604,I198876,I198893,I198842,I198915,I1372595,I198941,I198949,I198966,I1372589,I198983,I1372583,I199000,I199017,I1372610,I199034,I199051,I1372607,I199068,I198818,I199099,I199116,I199133,I199150,I198830,I198824,I199195,I1372592,I198839,I198833,I199240,I199257,I1372598,I199274,I1372601,I199291,I1372586,I199317,I199325,I198827,I198821,I199379,I199387,I198836,I199445,I551903,I199471,I199488,I199437,I199510,I551897,I199536,I199544,I199561,I551912,I199578,I551909,I199595,I199612,I551900,I199629,I551891,I199646,I551894,I199663,I199413,I199694,I199711,I199728,I199745,I199425,I199419,I199790,I551915,I199434,I199428,I199835,I199852,I551906,I199869,I199886,I199912,I199920,I199422,I199416,I199974,I199982,I199431,I200040,I200066,I200083,I200032,I200105,I200131,I200139,I200156,I200173,I200190,I200207,I200224,I200241,I200258,I200008,I200289,I200306,I200323,I200340,I200020,I200014,I200385,I200029,I200023,I200430,I200447,I200464,I200481,I200507,I200515,I200017,I200011,I200569,I200577,I200026,I200635,I200661,I200678,I200627,I200700,I200726,I200734,I200751,I200768,I200785,I200802,I200819,I200836,I200853,I200603,I200884,I200901,I200918,I200935,I200615,I200609,I200980,I200624,I200618,I201025,I201042,I201059,I201076,I201102,I201110,I200612,I200606,I201164,I201172,I200621,I201230,I611032,I201256,I201273,I201295,I611023,I201321,I201329,I201346,I611041,I201363,I611038,I201380,I201397,I611017,I201414,I611020,I201431,I611029,I201448,I201479,I201496,I201513,I201530,I201575,I611035,I201620,I201637,I201654,I611026,I201671,I201697,I201705,I201759,I201767,I201825,I1219889,I201851,I201868,I201817,I201890,I201916,I201924,I201941,I1219892,I201958,I1219904,I201975,I201992,I1219910,I202009,I1219901,I202026,I1219907,I202043,I201793,I202074,I202091,I202108,I202125,I201805,I201799,I202170,I1219898,I201814,I201808,I202215,I202232,I1219895,I202249,I1219913,I202266,I202292,I202300,I201802,I201796,I202354,I202362,I201811,I202420,I642822,I202446,I202463,I202412,I202485,I642813,I202511,I202519,I202536,I642831,I202553,I642828,I202570,I202587,I642807,I202604,I642810,I202621,I642819,I202638,I202388,I202669,I202686,I202703,I202720,I202400,I202394,I202765,I642825,I202409,I202403,I202810,I202827,I202844,I642816,I202861,I202887,I202895,I202397,I202391,I202949,I202957,I202406,I203015,I736455,I203041,I203058,I203080,I736452,I203106,I203114,I203131,I736458,I203148,I736443,I203165,I203182,I736446,I203199,I736467,I203216,I736464,I203233,I203264,I203281,I203298,I203315,I203360,I203405,I203422,I736449,I203439,I736461,I203456,I203482,I203490,I203544,I203552,I203610,I1390454,I203636,I203653,I203675,I1390445,I203701,I203709,I203726,I1390439,I203743,I1390433,I203760,I203777,I1390460,I203794,I203811,I1390457,I203828,I203859,I203876,I203893,I203910,I203955,I1390442,I204000,I204017,I1390448,I204034,I1390451,I204051,I1390436,I204077,I204085,I204139,I204147,I204205,I1100243,I204231,I204248,I204197,I204270,I204296,I204304,I204321,I1100246,I204338,I1100258,I204355,I204372,I1100264,I204389,I1100255,I204406,I1100261,I204423,I204173,I204454,I204471,I204488,I204505,I204185,I204179,I204550,I1100252,I204194,I204188,I204595,I204612,I1100249,I204629,I1100267,I204646,I204672,I204680,I204182,I204176,I204734,I204742,I204191,I204800,I204826,I204843,I204792,I204865,I204891,I204899,I204916,I204933,I204950,I204967,I204984,I205001,I205018,I204768,I205049,I205066,I205083,I205100,I204780,I204774,I205145,I204789,I204783,I205190,I205207,I205224,I205241,I205267,I205275,I204777,I204771,I205329,I205337,I204786,I205395,I541193,I205421,I205438,I205387,I205460,I541187,I205486,I205494,I205511,I541202,I205528,I541199,I205545,I205562,I541190,I205579,I541181,I205596,I541184,I205613,I205363,I205644,I205661,I205678,I205695,I205375,I205369,I205740,I541205,I205384,I205378,I205785,I205802,I541196,I205819,I205836,I205862,I205870,I205372,I205366,I205924,I205932,I205381,I205990,I337538,I206016,I206033,I206055,I337553,I206081,I206089,I206106,I337550,I206123,I206140,I206157,I337547,I206174,I337562,I206191,I337559,I206208,I206239,I206256,I206273,I206290,I206335,I337556,I206380,I206397,I337544,I206414,I337565,I206431,I337541,I206457,I206465,I206519,I206527,I206585,I1350589,I206611,I206628,I206650,I1350580,I206676,I206684,I206701,I1350574,I206718,I1350568,I206735,I206752,I1350595,I206769,I206786,I1350592,I206803,I206834,I206851,I206868,I206885,I206930,I1350577,I206975,I206992,I1350583,I207009,I1350586,I207026,I1350571,I207052,I207060,I207114,I207122,I207180,I1005976,I207206,I207223,I207172,I207245,I1005985,I207271,I207279,I207296,I1005973,I207313,I1005964,I207330,I207347,I1005970,I207364,I1005988,I207381,I1005961,I207398,I207148,I207429,I207446,I207463,I207480,I207160,I207154,I207525,I1005967,I207169,I207163,I207570,I207587,I1005979,I207604,I207621,I1005982,I207647,I207655,I207157,I207151,I207709,I207717,I207166,I207775,I889585,I207801,I207818,I207840,I889579,I207866,I207874,I207891,I889597,I207908,I207925,I207942,I207959,I889591,I207976,I889582,I207993,I208024,I208041,I208058,I208075,I208120,I889594,I208165,I208182,I889600,I208199,I208216,I889588,I208242,I208250,I208304,I208312,I208370,I967216,I208396,I208413,I208435,I967225,I208461,I208469,I208486,I967213,I208503,I967204,I208520,I208537,I967210,I208554,I967228,I208571,I967201,I208588,I208619,I208636,I208653,I208670,I208715,I967207,I208760,I208777,I967219,I208794,I208811,I967222,I208837,I208845,I208899,I208907,I208965,I306445,I208991,I209008,I208957,I209030,I306460,I209056,I209064,I209081,I306457,I209098,I209115,I209132,I306454,I209149,I306469,I209166,I306466,I209183,I208933,I209214,I209231,I209248,I209265,I208945,I208939,I209310,I306463,I208954,I208948,I209355,I209372,I306451,I209389,I306472,I209406,I306448,I209432,I209440,I208942,I208936,I209494,I209502,I208951,I209560,I209586,I209603,I209552,I209625,I209651,I209659,I209676,I209693,I209710,I209727,I209744,I209761,I209778,I209528,I209809,I209826,I209843,I209860,I209540,I209534,I209905,I209549,I209543,I209950,I209967,I209984,I210001,I210027,I210035,I209537,I209531,I210089,I210097,I209546,I210155,I210181,I210198,I210147,I210220,I210246,I210254,I210271,I210288,I210305,I210322,I210339,I210356,I210373,I210123,I210404,I210421,I210438,I210455,I210135,I210129,I210500,I210144,I210138,I210545,I210562,I210579,I210596,I210622,I210630,I210132,I210126,I210684,I210692,I210141,I210750,I1271451,I210776,I210793,I210742,I210815,I1271436,I210841,I210849,I210866,I1271454,I210883,I210900,I210917,I1271457,I210934,I1271448,I210951,I1271445,I210968,I210718,I210999,I211016,I211033,I211050,I210730,I210724,I211095,I1271442,I210739,I210733,I211140,I211157,I1271433,I211174,I1271439,I211191,I211217,I211225,I210727,I210721,I211279,I211287,I210736,I211345,I1332144,I211371,I211388,I211337,I211410,I1332135,I211436,I211444,I211461,I1332129,I211478,I1332123,I211495,I211512,I1332150,I211529,I211546,I1332147,I211563,I211313,I211594,I211611,I211628,I211645,I211325,I211319,I211690,I1332132,I211334,I211328,I211735,I211752,I1332138,I211769,I1332141,I211786,I1332126,I211812,I211820,I211322,I211316,I211874,I211882,I211331,I211940,I313823,I211966,I211983,I212005,I313838,I212031,I212039,I212056,I313835,I212073,I212090,I212107,I313832,I212124,I313847,I212141,I313844,I212158,I212189,I212206,I212223,I212240,I212285,I313841,I212330,I212347,I313829,I212364,I313850,I212381,I313826,I212407,I212415,I212469,I212477,I212535,I354929,I212561,I212578,I212527,I212600,I354944,I212626,I212634,I212651,I354941,I212668,I212685,I212702,I354938,I212719,I354953,I212736,I354950,I212753,I212503,I212784,I212801,I212818,I212835,I212515,I212509,I212880,I354947,I212524,I212518,I212925,I212942,I354935,I212959,I354956,I212976,I354932,I213002,I213010,I212512,I212506,I213064,I213072,I212521,I213130,I331741,I213156,I213173,I213122,I213195,I331756,I213221,I213229,I213246,I331753,I213263,I213280,I213297,I331750,I213314,I331765,I213331,I331762,I213348,I213098,I213379,I213396,I213413,I213430,I213110,I213104,I213475,I331759,I213119,I213113,I213520,I213537,I331747,I213554,I331768,I213571,I331744,I213597,I213605,I213107,I213101,I213659,I213667,I213116,I213725,I449082,I213751,I213768,I213717,I213790,I449070,I213816,I213824,I213841,I449079,I213858,I449076,I213875,I213892,I449067,I213909,I449073,I213926,I449058,I213943,I213693,I213974,I213991,I214008,I214025,I213705,I213699,I214070,I213714,I213708,I214115,I214132,I449064,I214149,I449061,I214166,I449085,I214192,I214200,I213702,I213696,I214254,I214262,I213711,I214320,I1051711,I214346,I214363,I214312,I214385,I1051720,I214411,I214419,I214436,I1051714,I214453,I1051708,I214470,I214487,I1051723,I214504,I214521,I1051717,I214538,I214288,I214569,I214586,I214603,I214620,I214300,I214294,I214665,I214309,I214303,I214710,I214727,I1051729,I214744,I1051726,I214761,I214787,I214795,I214297,I214291,I214849,I214857,I214306,I214915,I860073,I214941,I214958,I214907,I214980,I860067,I215006,I215014,I215031,I860085,I215048,I215065,I215082,I215099,I860079,I215116,I860070,I215133,I214883,I215164,I215181,I215198,I215215,I214895,I214889,I215260,I860082,I214904,I214898,I215305,I215322,I860088,I215339,I215356,I860076,I215382,I215390,I214892,I214886,I215444,I215452,I214901,I215510,I357037,I215536,I215553,I215502,I215575,I357052,I215601,I215609,I215626,I357049,I215643,I215660,I215677,I357046,I215694,I357061,I215711,I357058,I215728,I215478,I215759,I215776,I215793,I215810,I215490,I215484,I215855,I357055,I215499,I215493,I215900,I215917,I357043,I215934,I357064,I215951,I357040,I215977,I215985,I215487,I215481,I216039,I216047,I215496,I216105,I216131,I216148,I216097,I216170,I216196,I216204,I216221,I216238,I216255,I216272,I216289,I216306,I216323,I216073,I216354,I216371,I216388,I216405,I216085,I216079,I216450,I216094,I216088,I216495,I216512,I216529,I216546,I216572,I216580,I216082,I216076,I216634,I216642,I216091,I216700,I1262747,I216726,I216743,I216692,I216765,I1262732,I216791,I216799,I216816,I1262750,I216833,I216850,I216867,I1262753,I216884,I1262744,I216901,I1262741,I216918,I216668,I216949,I216966,I216983,I217000,I216680,I216674,I217045,I1262738,I216689,I216683,I217090,I217107,I1262729,I217124,I1262735,I217141,I217167,I217175,I216677,I216671,I217229,I217237,I216686,I217295,I1120473,I217321,I217338,I217287,I217360,I217386,I217394,I217411,I1120476,I217428,I1120488,I217445,I217462,I1120494,I217479,I1120485,I217496,I1120491,I217513,I217263,I217544,I217561,I217578,I217595,I217275,I217269,I217640,I1120482,I217284,I217278,I217685,I217702,I1120479,I217719,I1120497,I217736,I217762,I217770,I217272,I217266,I217824,I217832,I217281,I217890,I734143,I217916,I217933,I217955,I734140,I217981,I217989,I218006,I734146,I218023,I734131,I218040,I218057,I734134,I218074,I734155,I218091,I734152,I218108,I218139,I218156,I218173,I218190,I218235,I218280,I218297,I734137,I218314,I734149,I218331,I218357,I218365,I218419,I218427,I218485,I844790,I218511,I218528,I218477,I218550,I844784,I218576,I218584,I218601,I844802,I218618,I218635,I218652,I218669,I844796,I218686,I844787,I218703,I218453,I218734,I218751,I218768,I218785,I218465,I218459,I218830,I844799,I218474,I218468,I218875,I218892,I844805,I218909,I218926,I844793,I218952,I218960,I218462,I218456,I219014,I219022,I218471,I219080,I686169,I219106,I219123,I219072,I219145,I686166,I219171,I219179,I219196,I686172,I219213,I686157,I219230,I219247,I686160,I219264,I686181,I219281,I686178,I219298,I219048,I219329,I219346,I219363,I219380,I219060,I219054,I219425,I219069,I219063,I219470,I219487,I686163,I219504,I686175,I219521,I219547,I219555,I219057,I219051,I219609,I219617,I219066,I219675,I219701,I219718,I219740,I219766,I219774,I219791,I219808,I219825,I219842,I219859,I219876,I219893,I219924,I219941,I219958,I219975,I220020,I220065,I220082,I220099,I220116,I220142,I220150,I220204,I220212,I220270,I1072468,I220296,I220313,I220262,I220335,I1072477,I220361,I220369,I220386,I1072471,I220403,I1072465,I220420,I220437,I1072480,I220454,I220471,I1072474,I220488,I220238,I220519,I220536,I220553,I220570,I220250,I220244,I220615,I220259,I220253,I220660,I220677,I1072486,I220694,I1072483,I220711,I220737,I220745,I220247,I220241,I220799,I220807,I220256,I220865,I947190,I220891,I220908,I220857,I220930,I947199,I220956,I220964,I220981,I947187,I220998,I947178,I221015,I221032,I947184,I221049,I947202,I221066,I947175,I221083,I220833,I221114,I221131,I221148,I221165,I220845,I220839,I221210,I947181,I220854,I220848,I221255,I221272,I947193,I221289,I221306,I947196,I221332,I221340,I220842,I220836,I221394,I221402,I220851,I221460,I992410,I221486,I221503,I221452,I221525,I992419,I221551,I221559,I221576,I992407,I221593,I992398,I221610,I221627,I992404,I221644,I992422,I221661,I992395,I221678,I221428,I221709,I221726,I221743,I221760,I221440,I221434,I221805,I992401,I221449,I221443,I221850,I221867,I992413,I221884,I221901,I992416,I221927,I221935,I221437,I221431,I221989,I221997,I221446,I222055,I1358919,I222081,I222098,I222047,I222120,I1358910,I222146,I222154,I222171,I1358904,I222188,I1358898,I222205,I222222,I1358925,I222239,I222256,I1358922,I222273,I222023,I222304,I222321,I222338,I222355,I222035,I222029,I222400,I1358907,I222044,I222038,I222445,I222462,I1358913,I222479,I1358916,I222496,I1358901,I222522,I222530,I222032,I222026,I222584,I222592,I222041,I222650,I222676,I222693,I222642,I222715,I222741,I222749,I222766,I222783,I222800,I222817,I222834,I222851,I222868,I222618,I222899,I222916,I222933,I222950,I222630,I222624,I222995,I222639,I222633,I223040,I223057,I223074,I223091,I223117,I223125,I222627,I222621,I223179,I223187,I222636,I223245,I1391049,I223271,I223288,I223237,I223310,I1391040,I223336,I223344,I223361,I1391034,I223378,I1391028,I223395,I223412,I1391055,I223429,I223446,I1391052,I223463,I223213,I223494,I223511,I223528,I223545,I223225,I223219,I223590,I1391037,I223234,I223228,I223635,I223652,I1391043,I223669,I1391046,I223686,I1391031,I223712,I223720,I223222,I223216,I223774,I223782,I223231,I223840,I223866,I223883,I223832,I223905,I223931,I223939,I223956,I223973,I223990,I224007,I224024,I224041,I224058,I223808,I224089,I224106,I224123,I224140,I223820,I223814,I224185,I223829,I223823,I224230,I224247,I224264,I224281,I224307,I224315,I223817,I223811,I224369,I224377,I223826,I224435,I1295848,I224461,I224478,I224427,I224500,I1295860,I224526,I224534,I224551,I1295854,I224568,I1295866,I224585,I224602,I1295851,I224619,I1295863,I224636,I1295845,I224653,I224403,I224684,I224701,I224718,I224735,I224415,I224409,I224780,I1295857,I224424,I224418,I224825,I224842,I224859,I224876,I1295869,I224902,I224910,I224412,I224406,I224964,I224972,I224421,I225030,I395508,I225056,I225073,I225022,I225095,I395523,I225121,I225129,I225146,I395520,I225163,I225180,I225197,I395517,I225214,I395532,I225231,I395529,I225248,I224998,I225279,I225296,I225313,I225330,I225010,I225004,I225375,I395526,I225019,I225013,I225420,I225437,I395514,I225454,I395535,I225471,I395511,I225497,I225505,I225007,I225001,I225559,I225567,I225016,I225625,I326998,I225651,I225668,I225617,I225690,I327013,I225716,I225724,I225741,I327010,I225758,I225775,I225792,I327007,I225809,I327022,I225826,I327019,I225843,I225593,I225874,I225891,I225908,I225925,I225605,I225599,I225970,I327016,I225614,I225608,I226015,I226032,I327004,I226049,I327025,I226066,I327001,I226092,I226100,I225602,I225596,I226154,I226162,I225611,I226220,I798879,I226246,I226263,I226212,I226285,I798876,I226311,I226319,I226336,I798882,I226353,I798867,I226370,I226387,I798870,I226404,I798891,I226421,I798888,I226438,I226188,I226469,I226486,I226503,I226520,I226200,I226194,I226565,I226209,I226203,I226610,I226627,I798873,I226644,I798885,I226661,I226687,I226695,I226197,I226191,I226749,I226757,I226206,I226815,I1372009,I226841,I226858,I226880,I1372000,I226906,I226914,I226931,I1371994,I226948,I1371988,I226965,I226982,I1372015,I226999,I227016,I1372012,I227033,I227064,I227081,I227098,I227115,I227160,I1371997,I227205,I227222,I1372003,I227239,I1372006,I227256,I1371991,I227282,I227290,I227344,I227352,I227410,I934270,I227436,I227453,I227402,I227475,I934279,I227501,I227509,I227526,I934267,I227543,I934258,I227560,I227577,I934264,I227594,I934282,I227611,I934255,I227628,I227378,I227659,I227676,I227693,I227710,I227390,I227384,I227755,I934261,I227399,I227393,I227800,I227817,I934273,I227834,I227851,I934276,I227877,I227885,I227387,I227381,I227939,I227947,I227396,I228005,I228031,I228048,I227997,I228070,I228096,I228104,I228121,I228138,I228155,I228172,I228189,I228206,I228223,I227973,I228254,I228271,I228288,I228305,I227985,I227979,I228350,I227994,I227988,I228395,I228412,I228429,I228446,I228472,I228480,I227982,I227976,I228534,I228542,I227991,I228600,I497498,I228626,I228643,I228665,I497486,I228691,I228699,I228716,I497495,I228733,I497492,I228750,I228767,I497483,I228784,I497489,I228801,I497474,I228818,I228849,I228866,I228883,I228900,I228945,I228990,I229007,I497480,I229024,I497477,I229041,I497501,I229067,I229075,I229129,I229137,I229195,I229221,I229238,I229187,I229260,I229286,I229294,I229311,I229328,I229345,I229362,I229379,I229396,I229413,I229163,I229444,I229461,I229478,I229495,I229175,I229169,I229540,I229184,I229178,I229585,I229602,I229619,I229636,I229662,I229670,I229172,I229166,I229724,I229732,I229181,I229790,I647446,I229816,I229833,I229782,I229855,I647437,I229881,I229889,I229906,I647455,I229923,I647452,I229940,I229957,I647431,I229974,I647434,I229991,I647443,I230008,I229758,I230039,I230056,I230073,I230090,I229770,I229764,I230135,I647449,I229779,I229773,I230180,I230197,I230214,I647440,I230231,I230257,I230265,I229767,I229761,I230319,I230327,I229776,I230385,I758997,I230411,I230428,I230377,I230450,I758994,I230476,I230484,I230501,I759000,I230518,I758985,I230535,I230552,I758988,I230569,I759009,I230586,I759006,I230603,I230353,I230634,I230651,I230668,I230685,I230365,I230359,I230730,I230374,I230368,I230775,I230792,I758991,I230809,I759003,I230826,I230852,I230860,I230362,I230356,I230914,I230922,I230371,I230980,I1294114,I231006,I231023,I230972,I231045,I1294126,I231071,I231079,I231096,I1294120,I231113,I1294132,I231130,I231147,I1294117,I231164,I1294129,I231181,I1294111,I231198,I230948,I231229,I231246,I231263,I231280,I230960,I230954,I231325,I1294123,I230969,I230963,I231370,I231387,I231404,I231421,I1294135,I231447,I231455,I230957,I230951,I231509,I231517,I230966,I231575,I553688,I231601,I231618,I231567,I231640,I553682,I231666,I231674,I231691,I553697,I231708,I553694,I231725,I231742,I553685,I231759,I553676,I231776,I553679,I231793,I231543,I231824,I231841,I231858,I231875,I231555,I231549,I231920,I553700,I231564,I231558,I231965,I231982,I553691,I231999,I232016,I232042,I232050,I231552,I231546,I232104,I232112,I231561,I232170,I232196,I232213,I232162,I232235,I232261,I232269,I232286,I232303,I232320,I232337,I232354,I232371,I232388,I232138,I232419,I232436,I232453,I232470,I232150,I232144,I232515,I232159,I232153,I232560,I232577,I232594,I232611,I232637,I232645,I232147,I232141,I232699,I232707,I232156,I232765,I833196,I232791,I232808,I232757,I232830,I833190,I232856,I232864,I232881,I833208,I232898,I232915,I232932,I232949,I833202,I232966,I833193,I232983,I232733,I233014,I233031,I233048,I233065,I232745,I232739,I233110,I833205,I232754,I232748,I233155,I233172,I833211,I233189,I233206,I833199,I233232,I233240,I232742,I232736,I233294,I233302,I232751,I233360,I233386,I233403,I233352,I233425,I233451,I233459,I233476,I233493,I233510,I233527,I233544,I233561,I233578,I233328,I233609,I233626,I233643,I233660,I233340,I233334,I233705,I233349,I233343,I233750,I233767,I233784,I233801,I233827,I233835,I233337,I233331,I233889,I233897,I233346,I233955,I1101399,I233981,I233998,I233947,I234020,I234046,I234054,I234071,I1101402,I234088,I1101414,I234105,I234122,I1101420,I234139,I1101411,I234156,I1101417,I234173,I233923,I234204,I234221,I234238,I234255,I233935,I233929,I234300,I1101408,I233944,I233938,I234345,I234362,I1101405,I234379,I1101423,I234396,I234422,I234430,I233932,I233926,I234484,I234492,I233941,I234550,I907503,I234576,I234593,I234542,I234615,I907497,I234641,I234649,I234666,I907515,I234683,I234700,I234717,I234734,I907509,I234751,I907500,I234768,I234518,I234799,I234816,I234833,I234850,I234530,I234524,I234895,I907512,I234539,I234533,I234940,I234957,I907518,I234974,I234991,I907506,I235017,I235025,I234527,I234521,I235079,I235087,I234536,I235145,I457786,I235171,I235188,I235137,I235210,I457774,I235236,I235244,I235261,I457783,I235278,I457780,I235295,I235312,I457771,I235329,I457777,I235346,I457762,I235363,I235113,I235394,I235411,I235428,I235445,I235125,I235119,I235490,I235134,I235128,I235535,I235552,I457768,I235569,I457765,I235586,I457789,I235612,I235620,I235122,I235116,I235674,I235682,I235131,I235740,I503482,I235766,I235783,I235732,I235805,I503470,I235831,I235839,I235856,I503479,I235873,I503476,I235890,I235907,I503467,I235924,I503473,I235941,I503458,I235958,I235708,I235989,I236006,I236023,I236040,I235720,I235714,I236085,I235729,I235723,I236130,I236147,I503464,I236164,I503461,I236181,I503485,I236207,I236215,I235717,I235711,I236269,I236277,I235726,I236335,I946544,I236361,I236378,I236327,I236400,I946553,I236426,I236434,I236451,I946541,I236468,I946532,I236485,I236502,I946538,I236519,I946556,I236536,I946529,I236553,I236303,I236584,I236601,I236618,I236635,I236315,I236309,I236680,I946535,I236324,I236318,I236725,I236742,I946547,I236759,I236776,I946550,I236802,I236810,I236312,I236306,I236864,I236872,I236321,I236930,I1102555,I236956,I236973,I236922,I236995,I237021,I237029,I237046,I1102558,I237063,I1102570,I237080,I237097,I1102576,I237114,I1102567,I237131,I1102573,I237148,I236898,I237179,I237196,I237213,I237230,I236910,I236904,I237275,I1102564,I236919,I236913,I237320,I237337,I1102561,I237354,I1102579,I237371,I237397,I237405,I236907,I236901,I237459,I237467,I236916,I237525,I737611,I237551,I237568,I237517,I237590,I737608,I237616,I237624,I237641,I737614,I237658,I737599,I237675,I237692,I737602,I237709,I737623,I237726,I737620,I237743,I237493,I237774,I237791,I237808,I237825,I237505,I237499,I237870,I237514,I237508,I237915,I237932,I737605,I237949,I737617,I237966,I237992,I238000,I237502,I237496,I238054,I238062,I237511,I238120,I1323592,I238146,I238163,I238112,I238185,I1323604,I238211,I238219,I238236,I1323598,I238253,I1323610,I238270,I238287,I1323595,I238304,I1323607,I238321,I1323589,I238338,I238088,I238369,I238386,I238403,I238420,I238100,I238094,I238465,I1323601,I238109,I238103,I238510,I238527,I238544,I238561,I1323613,I238587,I238595,I238097,I238091,I238649,I238657,I238106,I238715,I729519,I238741,I238758,I238707,I238780,I729516,I238806,I238814,I238831,I729522,I238848,I729507,I238865,I238882,I729510,I238899,I729531,I238916,I729528,I238933,I238683,I238964,I238981,I238998,I239015,I238695,I238689,I239060,I238704,I238698,I239105,I239122,I729513,I239139,I729525,I239156,I239182,I239190,I238692,I238686,I239244,I239252,I238701,I239310,I641088,I239336,I239353,I239302,I239375,I641079,I239401,I239409,I239426,I641097,I239443,I641094,I239460,I239477,I641073,I239494,I641076,I239511,I641085,I239528,I239278,I239559,I239576,I239593,I239610,I239290,I239284,I239655,I641091,I239299,I239293,I239700,I239717,I239734,I641082,I239751,I239777,I239785,I239287,I239281,I239839,I239847,I239296,I239905,I535243,I239931,I239948,I239897,I239970,I535237,I239996,I240004,I240021,I535252,I240038,I535249,I240055,I240072,I535240,I240089,I535231,I240106,I535234,I240123,I239873,I240154,I240171,I240188,I240205,I239885,I239879,I240250,I535255,I239894,I239888,I240295,I240312,I535246,I240329,I240346,I240372,I240380,I239882,I239876,I240434,I240442,I239891,I240500,I586178,I240526,I240543,I240492,I240565,I586169,I240591,I240599,I240616,I586187,I240633,I586184,I240650,I240667,I586163,I240684,I586166,I240701,I586175,I240718,I240468,I240749,I240766,I240783,I240800,I240480,I240474,I240845,I586181,I240489,I240483,I240890,I240907,I240924,I586172,I240941,I240967,I240975,I240477,I240471,I241029,I241037,I240486,I241095,I1240697,I241121,I241138,I241087,I241160,I241186,I241194,I241211,I1240700,I241228,I1240712,I241245,I241262,I1240718,I241279,I1240709,I241296,I1240715,I241313,I241063,I241344,I241361,I241378,I241395,I241075,I241069,I241440,I1240706,I241084,I241078,I241485,I241502,I1240703,I241519,I1240721,I241536,I241562,I241570,I241072,I241066,I241624,I241632,I241081,I241690,I419750,I241716,I241733,I241682,I241755,I419765,I241781,I241789,I241806,I419762,I241823,I241840,I241857,I419759,I241874,I419774,I241891,I419771,I241908,I241658,I241939,I241956,I241973,I241990,I241670,I241664,I242035,I419768,I241679,I241673,I242080,I242097,I419756,I242114,I419777,I242131,I419753,I242157,I242165,I241667,I241661,I242219,I242227,I241676,I242285,I242311,I242328,I242277,I242350,I242376,I242384,I242401,I242418,I242435,I242452,I242469,I242486,I242503,I242253,I242534,I242551,I242568,I242585,I242265,I242259,I242630,I242274,I242268,I242675,I242692,I242709,I242726,I242752,I242760,I242262,I242256,I242814,I242822,I242271,I242880,I242906,I242923,I242945,I242971,I242979,I242996,I243013,I243030,I243047,I243064,I243081,I243098,I243129,I243146,I243163,I243180,I243225,I243270,I243287,I243304,I243321,I243347,I243355,I243409,I243417,I243475,I872194,I243501,I243518,I243467,I243540,I872188,I243566,I243574,I243591,I872206,I243608,I243625,I243642,I243659,I872200,I243676,I872191,I243693,I243443,I243724,I243741,I243758,I243775,I243455,I243449,I243820,I872203,I243464,I243458,I243865,I243882,I872209,I243899,I243916,I872197,I243942,I243950,I243452,I243446,I244004,I244012,I243461,I244070,I1061809,I244096,I244113,I244062,I244135,I1061818,I244161,I244169,I244186,I1061812,I244203,I1061806,I244220,I244237,I1061821,I244254,I244271,I1061815,I244288,I244038,I244319,I244336,I244353,I244370,I244050,I244044,I244415,I244059,I244053,I244460,I244477,I1061827,I244494,I1061824,I244511,I244537,I244545,I244047,I244041,I244599,I244607,I244056,I244665,I1316656,I244691,I244708,I244657,I244730,I1316668,I244756,I244764,I244781,I1316662,I244798,I1316674,I244815,I244832,I1316659,I244849,I1316671,I244866,I1316653,I244883,I244633,I244914,I244931,I244948,I244965,I244645,I244639,I245010,I1316665,I244654,I244648,I245055,I245072,I245089,I245106,I1316677,I245132,I245140,I244642,I244636,I245194,I245202,I244651,I245260,I245286,I245303,I245252,I245325,I245351,I245359,I245376,I245393,I245410,I245427,I245444,I245461,I245478,I245228,I245509,I245526,I245543,I245560,I245240,I245234,I245605,I245249,I245243,I245650,I245667,I245684,I245701,I245727,I245735,I245237,I245231,I245789,I245797,I245246,I245855,I294324,I245881,I245898,I245847,I245920,I294339,I245946,I245954,I245971,I294336,I245988,I246005,I246022,I294333,I246039,I294348,I246056,I294345,I246073,I245823,I246104,I246121,I246138,I246155,I245835,I245829,I246200,I294342,I245844,I245838,I246245,I246262,I294330,I246279,I294351,I246296,I294327,I246322,I246330,I245832,I245826,I246384,I246392,I245841,I246450,I482810,I246476,I246493,I246442,I246515,I482798,I246541,I246549,I246566,I482807,I246583,I482804,I246600,I246617,I482795,I246634,I482801,I246651,I482786,I246668,I246418,I246699,I246716,I246733,I246750,I246430,I246424,I246795,I246439,I246433,I246840,I246857,I482792,I246874,I482789,I246891,I482813,I246917,I246925,I246427,I246421,I246979,I246987,I246436,I247045,I965924,I247071,I247088,I247037,I247110,I965933,I247136,I247144,I247161,I965921,I247178,I965912,I247195,I247212,I965918,I247229,I965936,I247246,I965909,I247263,I247013,I247294,I247311,I247328,I247345,I247025,I247019,I247390,I965915,I247034,I247028,I247435,I247452,I965927,I247469,I247486,I965930,I247512,I247520,I247022,I247016,I247574,I247582,I247031,I247640,I1166135,I247666,I247683,I247632,I247705,I247731,I247739,I247756,I1166138,I247773,I1166150,I247790,I247807,I1166156,I247824,I1166147,I247841,I1166153,I247858,I247608,I247889,I247906,I247923,I247940,I247620,I247614,I247985,I1166144,I247629,I247623,I248030,I248047,I1166141,I248064,I1166159,I248081,I248107,I248115,I247617,I247611,I248169,I248177,I247626,I248235,I1181163,I248261,I248278,I248300,I248326,I248334,I248351,I1181166,I248368,I1181178,I248385,I248402,I1181184,I248419,I1181175,I248436,I1181181,I248453,I248484,I248501,I248518,I248535,I248580,I1181172,I248625,I248642,I1181169,I248659,I1181187,I248676,I248702,I248710,I248764,I248772,I248830,I1365464,I248856,I248873,I248822,I248895,I1365455,I248921,I248929,I248946,I1365449,I248963,I1365443,I248980,I248997,I1365470,I249014,I249031,I1365467,I249048,I248798,I249079,I249096,I249113,I249130,I248810,I248804,I249175,I1365452,I248819,I248813,I249220,I249237,I1365458,I249254,I1365461,I249271,I1365446,I249297,I249305,I248807,I248801,I249359,I249367,I248816,I249425,I389711,I249451,I249468,I249417,I249490,I389726,I249516,I249524,I249541,I389723,I249558,I249575,I249592,I389720,I249609,I389735,I249626,I389732,I249643,I249393,I249674,I249691,I249708,I249725,I249405,I249399,I249770,I389729,I249414,I249408,I249815,I249832,I389717,I249849,I389738,I249866,I389714,I249892,I249900,I249402,I249396,I249954,I249962,I249411,I250020,I718537,I250046,I250063,I250012,I250085,I718534,I250111,I250119,I250136,I718540,I250153,I718525,I250170,I250187,I718528,I250204,I718549,I250221,I718546,I250238,I249988,I250269,I250286,I250303,I250320,I250000,I249994,I250365,I250009,I250003,I250410,I250427,I718531,I250444,I718543,I250461,I250487,I250495,I249997,I249991,I250549,I250557,I250006,I250615,I1066297,I250641,I250658,I250607,I250680,I1066306,I250706,I250714,I250731,I1066300,I250748,I1066294,I250765,I250782,I1066309,I250799,I250816,I1066303,I250833,I250583,I250864,I250881,I250898,I250915,I250595,I250589,I250960,I250604,I250598,I251005,I251022,I1066315,I251039,I1066312,I251056,I251082,I251090,I250592,I250586,I251144,I251152,I250601,I251210,I1392239,I251236,I251253,I251202,I251275,I1392230,I251301,I251309,I251326,I1392224,I251343,I1392218,I251360,I251377,I1392245,I251394,I251411,I1392242,I251428,I251178,I251459,I251476,I251493,I251510,I251190,I251184,I251555,I1392227,I251199,I251193,I251600,I251617,I1392233,I251634,I1392236,I251651,I1392221,I251677,I251685,I251187,I251181,I251739,I251747,I251196,I251805,I536433,I251831,I251848,I251797,I251870,I536427,I251896,I251904,I251921,I536442,I251938,I536439,I251955,I251972,I536430,I251989,I536421,I252006,I536424,I252023,I251773,I252054,I252071,I252088,I252105,I251785,I251779,I252150,I536445,I251794,I251788,I252195,I252212,I536436,I252229,I252246,I252272,I252280,I251782,I251776,I252334,I252342,I251791,I252400,I490426,I252426,I252443,I252392,I252465,I490414,I252491,I252499,I252516,I490423,I252533,I490420,I252550,I252567,I490411,I252584,I490417,I252601,I490402,I252618,I252368,I252649,I252666,I252683,I252700,I252380,I252374,I252745,I252389,I252383,I252790,I252807,I490408,I252824,I490405,I252841,I490429,I252867,I252875,I252377,I252371,I252929,I252937,I252386,I252995,I632996,I253021,I253038,I252987,I253060,I632987,I253086,I253094,I253111,I633005,I253128,I633002,I253145,I253162,I632981,I253179,I632984,I253196,I632993,I253213,I252963,I253244,I253261,I253278,I253295,I252975,I252969,I253340,I632999,I252984,I252978,I253385,I253402,I253419,I632990,I253436,I253462,I253470,I252972,I252966,I253524,I253532,I252981,I253590,I253616,I253633,I253582,I253655,I253681,I253689,I253706,I253723,I253740,I253757,I253774,I253791,I253808,I253558,I253839,I253856,I253873,I253890,I253570,I253564,I253935,I253579,I253573,I253980,I253997,I254014,I254031,I254057,I254065,I253567,I253561,I254119,I254127,I253576,I254185,I1191567,I254211,I254228,I254177,I254250,I254276,I254284,I254301,I1191570,I254318,I1191582,I254335,I254352,I1191588,I254369,I1191579,I254386,I1191585,I254403,I254153,I254434,I254451,I254468,I254485,I254165,I254159,I254530,I1191576,I254174,I254168,I254575,I254592,I1191573,I254609,I1191591,I254626,I254652,I254660,I254162,I254156,I254714,I254722,I254171,I254780,I1118161,I254806,I254823,I254845,I254871,I254879,I254896,I1118164,I254913,I1118176,I254930,I254947,I1118182,I254964,I1118173,I254981,I1118179,I254998,I255029,I255046,I255063,I255080,I255125,I1118170,I255170,I255187,I1118167,I255204,I1118185,I255221,I255247,I255255,I255309,I255317,I255375,I255401,I255418,I255440,I255466,I255474,I255491,I255508,I255525,I255542,I255559,I255576,I255593,I255624,I255641,I255658,I255675,I255720,I255765,I255782,I255799,I255816,I255842,I255850,I255904,I255912,I255970,I1238963,I255996,I256013,I255962,I256035,I256061,I256069,I256086,I1238966,I256103,I1238978,I256120,I256137,I1238984,I256154,I1238975,I256171,I1238981,I256188,I255938,I256219,I256236,I256253,I256270,I255950,I255944,I256315,I1238972,I255959,I255953,I256360,I256377,I1238969,I256394,I1238987,I256411,I256437,I256445,I255947,I255941,I256499,I256507,I255956,I256565,I418169,I256591,I256608,I256557,I256630,I418184,I256656,I256664,I256681,I418181,I256698,I256715,I256732,I418178,I256749,I418193,I256766,I418190,I256783,I256533,I256814,I256831,I256848,I256865,I256545,I256539,I256910,I418187,I256554,I256548,I256955,I256972,I418175,I256989,I418196,I257006,I418172,I257032,I257040,I256542,I256536,I257094,I257102,I256551,I257160,I774603,I257186,I257203,I257152,I257225,I774600,I257251,I257259,I257276,I774606,I257293,I774591,I257310,I257327,I774594,I257344,I774615,I257361,I774612,I257378,I257128,I257409,I257426,I257443,I257460,I257140,I257134,I257505,I257149,I257143,I257550,I257567,I774597,I257584,I774609,I257601,I257627,I257635,I257137,I257131,I257689,I257697,I257146,I257755,I257781,I257798,I257820,I257846,I257854,I257871,I257888,I257905,I257922,I257939,I257956,I257973,I258004,I258021,I258038,I258055,I258100,I258145,I258162,I258179,I258196,I258222,I258230,I258284,I258292,I258350,I995640,I258376,I258393,I258342,I258415,I995649,I258441,I258449,I258466,I995637,I258483,I995628,I258500,I258517,I995634,I258534,I995652,I258551,I995625,I258568,I258318,I258599,I258616,I258633,I258650,I258330,I258324,I258695,I995631,I258339,I258333,I258740,I258757,I995643,I258774,I258791,I995646,I258817,I258825,I258327,I258321,I258879,I258887,I258336,I258945,I763043,I258971,I258988,I258937,I259010,I763040,I259036,I259044,I259061,I763046,I259078,I763031,I259095,I259112,I763034,I259129,I763055,I259146,I763052,I259163,I258913,I259194,I259211,I259228,I259245,I258925,I258919,I259290,I258934,I258928,I259335,I259352,I763037,I259369,I763049,I259386,I259412,I259420,I258922,I258916,I259474,I259482,I258931,I259540,I869032,I259566,I259583,I259532,I259605,I869026,I259631,I259639,I259656,I869044,I259673,I259690,I259707,I259724,I869038,I259741,I869029,I259758,I259508,I259789,I259806,I259823,I259840,I259520,I259514,I259885,I869041,I259529,I259523,I259930,I259947,I869047,I259964,I259981,I869035,I260007,I260015,I259517,I259511,I260069,I260077,I259526,I260135,I301702,I260161,I260178,I260127,I260200,I301717,I260226,I260234,I260251,I301714,I260268,I260285,I260302,I301711,I260319,I301726,I260336,I301723,I260353,I260103,I260384,I260401,I260418,I260435,I260115,I260109,I260480,I301720,I260124,I260118,I260525,I260542,I301708,I260559,I301729,I260576,I301705,I260602,I260610,I260112,I260106,I260664,I260672,I260121,I260730,I1243587,I260756,I260773,I260722,I260795,I260821,I260829,I260846,I1243590,I260863,I1243602,I260880,I260897,I1243608,I260914,I1243599,I260931,I1243605,I260948,I260698,I260979,I260996,I261013,I261030,I260710,I260704,I261075,I1243596,I260719,I260713,I261120,I261137,I1243593,I261154,I1243611,I261171,I261197,I261205,I260707,I260701,I261259,I261267,I260716,I261325,I261351,I261368,I261317,I261390,I261416,I261424,I261441,I261458,I261475,I261492,I261509,I261526,I261543,I261293,I261574,I261591,I261608,I261625,I261305,I261299,I261670,I261314,I261308,I261715,I261732,I261749,I261766,I261792,I261800,I261302,I261296,I261854,I261862,I261311,I261920,I956880,I261946,I261963,I261912,I261985,I956889,I262011,I262019,I262036,I956877,I262053,I956868,I262070,I262087,I956874,I262104,I956892,I262121,I956865,I262138,I261888,I262169,I262186,I262203,I262220,I261900,I261894,I262265,I956871,I261909,I261903,I262310,I262327,I956883,I262344,I262361,I956886,I262387,I262395,I261897,I261891,I262449,I262457,I261906,I262515,I1228559,I262541,I262558,I262507,I262580,I262606,I262614,I262631,I1228562,I262648,I1228574,I262665,I262682,I1228580,I262699,I1228571,I262716,I1228577,I262733,I262483,I262764,I262781,I262798,I262815,I262495,I262489,I262860,I1228568,I262504,I262498,I262905,I262922,I1228565,I262939,I1228583,I262956,I262982,I262990,I262492,I262486,I263044,I263052,I262501,I263110,I263136,I263153,I263102,I263175,I263201,I263209,I263226,I263243,I263260,I263277,I263294,I263311,I263328,I263078,I263359,I263376,I263393,I263410,I263090,I263084,I263455,I263099,I263093,I263500,I263517,I263534,I263551,I263577,I263585,I263087,I263081,I263639,I263647,I263096,I263705,I681545,I263731,I263748,I263770,I681542,I263796,I263804,I263821,I681548,I263838,I681533,I263855,I263872,I681536,I263889,I681557,I263906,I681554,I263923,I263954,I263971,I263988,I264005,I264050,I264095,I264112,I681539,I264129,I681551,I264146,I264172,I264180,I264234,I264242,I264300,I417115,I264326,I264343,I264365,I417130,I264391,I264399,I264416,I417127,I264433,I264450,I264467,I417124,I264484,I417139,I264501,I417136,I264518,I264549,I264566,I264583,I264600,I264645,I417133,I264690,I264707,I417121,I264724,I417142,I264741,I417118,I264767,I264775,I264829,I264837,I264895,I931040,I264921,I264938,I264887,I264960,I931049,I264986,I264994,I265011,I931037,I265028,I931028,I265045,I265062,I931034,I265079,I931052,I265096,I931025,I265113,I264863,I265144,I265161,I265178,I265195,I264875,I264869,I265240,I931031,I264884,I264878,I265285,I265302,I931043,I265319,I265336,I931046,I265362,I265370,I264872,I264866,I265424,I265432,I264881,I265490,I1013728,I265516,I265533,I265482,I265555,I1013737,I265581,I265589,I265606,I1013725,I265623,I1013716,I265640,I265657,I1013722,I265674,I1013740,I265691,I1013713,I265708,I265458,I265739,I265756,I265773,I265790,I265470,I265464,I265835,I1013719,I265479,I265473,I265880,I265897,I1013731,I265914,I265931,I1013734,I265957,I265965,I265467,I265461,I266019,I266027,I265476,I266085,I266111,I266128,I266077,I266150,I266176,I266184,I266201,I266218,I266235,I266252,I266269,I266286,I266303,I266053,I266334,I266351,I266368,I266385,I266065,I266059,I266430,I266074,I266068,I266475,I266492,I266509,I266526,I266552,I266560,I266062,I266056,I266614,I266622,I266071,I266680,I1266555,I266706,I266723,I266672,I266745,I1266540,I266771,I266779,I266796,I1266558,I266813,I266830,I266847,I1266561,I266864,I1266552,I266881,I1266549,I266898,I266648,I266929,I266946,I266963,I266980,I266660,I266654,I267025,I1266546,I266669,I266663,I267070,I267087,I1266537,I267104,I1266543,I267121,I267147,I267155,I266657,I266651,I267209,I267217,I266666,I267275,I836358,I267301,I267318,I267267,I267340,I836352,I267366,I267374,I267391,I836370,I267408,I267425,I267442,I267459,I836364,I267476,I836355,I267493,I267243,I267524,I267541,I267558,I267575,I267255,I267249,I267620,I836367,I267264,I267258,I267665,I267682,I836373,I267699,I267716,I836361,I267742,I267750,I267252,I267246,I267804,I267812,I267261,I267870,I1386289,I267896,I267913,I267862,I267935,I1386280,I267961,I267969,I267986,I1386274,I268003,I1386268,I268020,I268037,I1386295,I268054,I268071,I1386292,I268088,I267838,I268119,I268136,I268153,I268170,I267850,I267844,I268215,I1386277,I267859,I267853,I268260,I268277,I1386283,I268294,I1386286,I268311,I1386271,I268337,I268345,I267847,I267841,I268399,I268407,I267856,I268465,I601784,I268491,I268508,I268457,I268530,I601775,I268556,I268564,I268581,I601793,I268598,I601790,I268615,I268632,I601769,I268649,I601772,I268666,I601781,I268683,I268433,I268714,I268731,I268748,I268765,I268445,I268439,I268810,I601787,I268454,I268448,I268855,I268872,I268889,I601778,I268906,I268932,I268940,I268442,I268436,I268994,I269002,I268451,I269060,I673453,I269086,I269103,I269052,I269125,I673450,I269151,I269159,I269176,I673456,I269193,I673441,I269210,I269227,I673444,I269244,I673465,I269261,I673462,I269278,I269028,I269309,I269326,I269343,I269360,I269040,I269034,I269405,I269049,I269043,I269450,I269467,I673447,I269484,I673459,I269501,I269527,I269535,I269037,I269031,I269589,I269597,I269046,I269655,I411845,I269681,I269698,I269647,I269720,I411860,I269746,I269754,I269771,I411857,I269788,I269805,I269822,I411854,I269839,I411869,I269856,I411866,I269873,I269623,I269904,I269921,I269938,I269955,I269635,I269629,I270000,I411863,I269644,I269638,I270045,I270062,I411851,I270079,I411872,I270096,I411848,I270122,I270130,I269632,I269626,I270184,I270192,I269641,I270250,I270276,I270293,I270242,I270315,I270341,I270349,I270366,I270383,I270400,I270417,I270434,I270451,I270468,I270218,I270499,I270516,I270533,I270550,I270230,I270224,I270595,I270239,I270233,I270640,I270657,I270674,I270691,I270717,I270725,I270227,I270221,I270779,I270787,I270236,I270845,I341227,I270871,I270888,I270837,I270910,I341242,I270936,I270944,I270961,I341239,I270978,I270995,I271012,I341236,I271029,I341251,I271046,I341248,I271063,I270813,I271094,I271111,I271128,I271145,I270825,I270819,I271190,I341245,I270834,I270828,I271235,I271252,I341233,I271269,I341254,I271286,I341230,I271312,I271320,I270822,I270816,I271374,I271382,I270831,I271440,I1143015,I271466,I271483,I271432,I271505,I271531,I271539,I271556,I1143018,I271573,I1143030,I271590,I271607,I1143036,I271624,I1143027,I271641,I1143033,I271658,I271408,I271689,I271706,I271723,I271740,I271420,I271414,I271785,I1143024,I271429,I271423,I271830,I271847,I1143021,I271864,I1143039,I271881,I271907,I271915,I271417,I271411,I271969,I271977,I271426,I272035,I741079,I272061,I272078,I272027,I272100,I741076,I272126,I272134,I272151,I741082,I272168,I741067,I272185,I272202,I741070,I272219,I741091,I272236,I741088,I272253,I272003,I272284,I272301,I272318,I272335,I272015,I272009,I272380,I272024,I272018,I272425,I272442,I741073,I272459,I741085,I272476,I272502,I272510,I272012,I272006,I272564,I272572,I272021,I272630,I987242,I272656,I272673,I272695,I987251,I272721,I272729,I272746,I987239,I272763,I987230,I272780,I272797,I987236,I272814,I987254,I272831,I987227,I272848,I272879,I272896,I272913,I272930,I272975,I987233,I273020,I273037,I987245,I273054,I273071,I987248,I273097,I273105,I273159,I273167,I273225,I455066,I273251,I273268,I273217,I273290,I455054,I273316,I273324,I273341,I455063,I273358,I455060,I273375,I273392,I455051,I273409,I455057,I273426,I455042,I273443,I273193,I273474,I273491,I273508,I273525,I273205,I273199,I273570,I273214,I273208,I273615,I273632,I455048,I273649,I455045,I273666,I455069,I273692,I273700,I273202,I273196,I273754,I273762,I273211,I273820,I388657,I273846,I273863,I273812,I273885,I388672,I273911,I273919,I273936,I388669,I273953,I273970,I273987,I388666,I274004,I388681,I274021,I388678,I274038,I273788,I274069,I274086,I274103,I274120,I273800,I273794,I274165,I388675,I273809,I273803,I274210,I274227,I388663,I274244,I388684,I274261,I388660,I274287,I274295,I273797,I273791,I274349,I274357,I273806,I274415,I1175383,I274441,I274458,I274407,I274480,I274506,I274514,I274531,I1175386,I274548,I1175398,I274565,I274582,I1175404,I274599,I1175395,I274616,I1175401,I274633,I274383,I274664,I274681,I274698,I274715,I274395,I274389,I274760,I1175392,I274404,I274398,I274805,I274822,I1175389,I274839,I1175407,I274856,I274882,I274890,I274392,I274386,I274944,I274952,I274401,I275010,I275036,I275053,I275002,I275075,I275101,I275109,I275126,I275143,I275160,I275177,I275194,I275211,I275228,I274978,I275259,I275276,I275293,I275310,I274990,I274984,I275355,I274999,I274993,I275400,I275417,I275434,I275451,I275477,I275485,I274987,I274981,I275539,I275547,I274996,I275605,I275631,I275648,I275597,I275670,I275696,I275704,I275721,I275738,I275755,I275772,I275789,I275806,I275823,I275573,I275854,I275871,I275888,I275905,I275585,I275579,I275950,I275594,I275588,I275995,I276012,I276029,I276046,I276072,I276080,I275582,I275576,I276134,I276142,I275591,I276200,I629528,I276226,I276243,I276192,I276265,I629519,I276291,I276299,I276316,I629537,I276333,I629534,I276350,I276367,I629513,I276384,I629516,I276401,I629525,I276418,I276168,I276449,I276466,I276483,I276500,I276180,I276174,I276545,I629531,I276189,I276183,I276590,I276607,I276624,I629522,I276641,I276667,I276675,I276177,I276171,I276729,I276737,I276186,I276795,I505658,I276821,I276838,I276787,I276860,I505646,I276886,I276894,I276911,I505655,I276928,I505652,I276945,I276962,I505643,I276979,I505649,I276996,I505634,I277013,I276763,I277044,I277061,I277078,I277095,I276775,I276769,I277140,I276784,I276778,I277185,I277202,I505640,I277219,I505637,I277236,I505661,I277262,I277270,I276772,I276766,I277324,I277332,I276781,I277390,I1242431,I277416,I277433,I277455,I277481,I277489,I277506,I1242434,I277523,I1242446,I277540,I277557,I1242452,I277574,I1242443,I277591,I1242449,I277608,I277639,I277656,I277673,I277690,I277735,I1242440,I277780,I277797,I1242437,I277814,I1242455,I277831,I277857,I277865,I277919,I277927,I277985,I587334,I278011,I278028,I277977,I278050,I587325,I278076,I278084,I278101,I587343,I278118,I587340,I278135,I278152,I587319,I278169,I587322,I278186,I587331,I278203,I277953,I278234,I278251,I278268,I278285,I277965,I277959,I278330,I587337,I277974,I277968,I278375,I278392,I278409,I587328,I278426,I278452,I278460,I277962,I277956,I278514,I278522,I277971,I278580,I1275803,I278606,I278623,I278572,I278645,I1275788,I278671,I278679,I278696,I1275806,I278713,I278730,I278747,I1275809,I278764,I1275800,I278781,I1275797,I278798,I278548,I278829,I278846,I278863,I278880,I278560,I278554,I278925,I1275794,I278569,I278563,I278970,I278987,I1275785,I279004,I1275791,I279021,I279047,I279055,I278557,I278551,I279109,I279117,I278566,I279175,I490970,I279201,I279218,I279167,I279240,I490958,I279266,I279274,I279291,I490967,I279308,I490964,I279325,I279342,I490955,I279359,I490961,I279376,I490946,I279393,I279143,I279424,I279441,I279458,I279475,I279155,I279149,I279520,I279164,I279158,I279565,I279582,I490952,I279599,I490949,I279616,I490973,I279642,I279650,I279152,I279146,I279704,I279712,I279161,I279770,I620858,I279796,I279813,I279762,I279835,I620849,I279861,I279869,I279886,I620867,I279903,I620864,I279920,I279937,I620843,I279954,I620846,I279971,I620855,I279988,I279738,I280019,I280036,I280053,I280070,I279750,I279744,I280115,I620861,I279759,I279753,I280160,I280177,I280194,I620852,I280211,I280237,I280245,I279747,I279741,I280299,I280307,I279756,I280365,I478458,I280391,I280408,I280357,I280430,I478446,I280456,I280464,I280481,I478455,I280498,I478452,I280515,I280532,I478443,I280549,I478449,I280566,I478434,I280583,I280333,I280614,I280631,I280648,I280665,I280345,I280339,I280710,I280354,I280348,I280755,I280772,I478440,I280789,I478437,I280806,I478461,I280832,I280840,I280342,I280336,I280894,I280902,I280351,I280960,I513274,I280986,I281003,I281025,I513262,I281051,I281059,I281076,I513271,I281093,I513268,I281110,I281127,I513259,I281144,I513265,I281161,I513250,I281178,I281209,I281226,I281243,I281260,I281305,I281350,I281367,I513256,I281384,I513253,I281401,I513277,I281427,I281435,I281489,I281497,I281555,I756685,I281581,I281598,I281547,I281620,I756682,I281646,I281654,I281671,I756688,I281688,I756673,I281705,I281722,I756676,I281739,I756697,I281756,I756694,I281773,I281523,I281804,I281821,I281838,I281855,I281535,I281529,I281900,I281544,I281538,I281945,I281962,I756679,I281979,I756691,I281996,I282022,I282030,I281532,I281526,I282084,I282092,I281541,I282150,I1046662,I282176,I282193,I282142,I282215,I1046671,I282241,I282249,I282266,I1046665,I282283,I1046659,I282300,I282317,I1046674,I282334,I282351,I1046668,I282368,I282118,I282399,I282416,I282433,I282450,I282130,I282124,I282495,I282139,I282133,I282540,I282557,I1046680,I282574,I1046677,I282591,I282617,I282625,I282127,I282121,I282679,I282687,I282136,I282745,I282771,I282788,I282737,I282810,I282836,I282844,I282861,I282878,I282895,I282912,I282929,I282946,I282963,I282713,I282994,I283011,I283028,I283045,I282725,I282719,I283090,I282734,I282728,I283135,I283152,I283169,I283186,I283212,I283220,I282722,I282716,I283274,I283282,I282731,I283340,I1158043,I283366,I283383,I283332,I283405,I283431,I283439,I283456,I1158046,I283473,I1158058,I283490,I283507,I1158064,I283524,I1158055,I283541,I1158061,I283558,I283308,I283589,I283606,I283623,I283640,I283320,I283314,I283685,I1158052,I283329,I283323,I283730,I283747,I1158049,I283764,I1158067,I283781,I283807,I283815,I283317,I283311,I283869,I283877,I283326,I283935,I928456,I283961,I283978,I283927,I284000,I928465,I284026,I284034,I284051,I928453,I284068,I928444,I284085,I284102,I928450,I284119,I928468,I284136,I928441,I284153,I283903,I284184,I284201,I284218,I284235,I283915,I283909,I284280,I928447,I283924,I283918,I284325,I284342,I928459,I284359,I284376,I928462,I284402,I284410,I283912,I283906,I284464,I284472,I283921,I284530,I921350,I284556,I284573,I284522,I284595,I921359,I284621,I284629,I284646,I921347,I284663,I921338,I284680,I284697,I921344,I284714,I921362,I284731,I921335,I284748,I284498,I284779,I284796,I284813,I284830,I284510,I284504,I284875,I921341,I284519,I284513,I284920,I284937,I921353,I284954,I284971,I921356,I284997,I285005,I284507,I284501,I285059,I285067,I284516,I285125,I688481,I285151,I285168,I285190,I688478,I285216,I285224,I285241,I688484,I285258,I688469,I285275,I285292,I688472,I285309,I688493,I285326,I688490,I285343,I285374,I285391,I285408,I285425,I285470,I285515,I285532,I688475,I285549,I688487,I285566,I285592,I285600,I285654,I285662,I285720,I913827,I285746,I285763,I285712,I285785,I913821,I285811,I285819,I285836,I913839,I285853,I285870,I285887,I285904,I913833,I285921,I913824,I285938,I285688,I285969,I285986,I286003,I286020,I285700,I285694,I286065,I913836,I285709,I285703,I286110,I286127,I913842,I286144,I286161,I913830,I286187,I286195,I285697,I285691,I286249,I286257,I285706,I286315,I286341,I286358,I286307,I286380,I286406,I286414,I286431,I286448,I286465,I286482,I286499,I286516,I286533,I286283,I286564,I286581,I286598,I286615,I286295,I286289,I286660,I286304,I286298,I286705,I286722,I286739,I286756,I286782,I286790,I286292,I286286,I286844,I286852,I286301,I286910,I1004038,I286936,I286953,I286902,I286975,I1004047,I287001,I287009,I287026,I1004035,I287043,I1004026,I287060,I287077,I1004032,I287094,I1004050,I287111,I1004023,I287128,I286878,I287159,I287176,I287193,I287210,I286890,I286884,I287255,I1004029,I286899,I286893,I287300,I287317,I1004041,I287334,I287351,I1004044,I287377,I287385,I286887,I286881,I287439,I287447,I286896,I287508,I541779,I287534,I287542,I541791,I287559,I541776,I287585,I287476,I287607,I541800,I287633,I287641,I541797,I287658,I287684,I287500,I287706,I287482,I541788,I287746,I287763,I287771,I287788,I287485,I287819,I541785,I287836,I541794,I287862,I287870,I287473,I287491,I287915,I541782,I287932,I287494,I287479,I287488,I287497,I288035,I932320,I288061,I288069,I932317,I932335,I288086,I932326,I288112,I288003,I288134,I932341,I288160,I288168,I932323,I288185,I288211,I288027,I288233,I288009,I932329,I288273,I288290,I288298,I288315,I288012,I288346,I932344,I288363,I932332,I288389,I288397,I288000,I288018,I288442,I932338,I288459,I288021,I288006,I288015,I288024,I288562,I1096197,I288588,I288596,I1096212,I288613,I1096215,I288639,I288530,I288661,I1096221,I288687,I288695,I1096203,I288712,I288738,I288554,I288760,I288536,I1096200,I288800,I288817,I288825,I288842,I288539,I288873,I1096206,I288890,I1096218,I288916,I288924,I288527,I288545,I288969,I1096209,I288986,I288548,I288533,I288542,I288551,I289089,I1391644,I289115,I289123,I1391623,I289140,I1391650,I289166,I289057,I289188,I1391638,I289214,I289222,I1391641,I289239,I289265,I289081,I289287,I289063,I1391632,I289327,I289344,I289352,I289369,I289066,I289400,I1391629,I1391626,I289417,I1391647,I289443,I289451,I289054,I289072,I289496,I1391635,I289513,I289075,I289060,I289069,I289078,I289616,I1134923,I289642,I289650,I1134938,I289667,I1134941,I289693,I289584,I289715,I1134947,I289741,I289749,I1134929,I289766,I289792,I289608,I289814,I289590,I1134926,I289854,I289871,I289879,I289896,I289593,I289927,I1134932,I289944,I1134944,I289970,I289978,I289581,I289599,I290023,I1134935,I290040,I289602,I289587,I289596,I289605,I290143,I959452,I290169,I290177,I959449,I959467,I290194,I959458,I290220,I290111,I290242,I959473,I290268,I290276,I959455,I290293,I290319,I290135,I290341,I290117,I959461,I290381,I290398,I290406,I290423,I290120,I290454,I959476,I290471,I959464,I290497,I290505,I290108,I290126,I290550,I959470,I290567,I290129,I290114,I290123,I290132,I290670,I290696,I290704,I290721,I290747,I290638,I290769,I290795,I290803,I290820,I290846,I290662,I290868,I290644,I290908,I290925,I290933,I290950,I290647,I290981,I290998,I291024,I291032,I290635,I290653,I291077,I291094,I290656,I290641,I290650,I290659,I291197,I680389,I291223,I291231,I680380,I680395,I291248,I680401,I291274,I291165,I291296,I680386,I291322,I291330,I291347,I291373,I291189,I291395,I291171,I680383,I291435,I291452,I291460,I291477,I291174,I291508,I680377,I680392,I291525,I291551,I291559,I291162,I291180,I291604,I680398,I291621,I291183,I291168,I291177,I291186,I291724,I646868,I291750,I291758,I646853,I646856,I291775,I646871,I291801,I291692,I291823,I646865,I291849,I291857,I291874,I291900,I291716,I291922,I291698,I646862,I291962,I291979,I291987,I292004,I291701,I292035,I646877,I292052,I646874,I292078,I292086,I291689,I291707,I292131,I646859,I292148,I291710,I291695,I291704,I291713,I292251,I292277,I292285,I292302,I292328,I292350,I292376,I292384,I292401,I292427,I292449,I292489,I292506,I292514,I292531,I292562,I292579,I292605,I292613,I292658,I292675,I292778,I1344044,I292804,I292812,I1344023,I292829,I1344050,I292855,I292746,I292877,I1344038,I292903,I292911,I1344041,I292928,I292954,I292770,I292976,I292752,I1344032,I293016,I293033,I293041,I293058,I292755,I293089,I1344029,I1344026,I293106,I1344047,I293132,I293140,I292743,I292761,I293185,I1344035,I293202,I292764,I292749,I292758,I292767,I293305,I1092151,I293331,I293339,I1092166,I293356,I1092169,I293382,I293273,I293404,I1092175,I293430,I293438,I1092157,I293455,I293481,I293297,I293503,I293279,I1092154,I293543,I293560,I293568,I293585,I293282,I293616,I1092160,I293633,I1092172,I293659,I293667,I293270,I293288,I293712,I1092163,I293729,I293291,I293276,I293285,I293294,I293832,I749749,I293858,I293866,I749740,I749755,I293883,I749761,I293909,I293800,I293931,I749746,I293957,I293965,I293982,I294008,I293824,I294030,I293806,I749743,I294070,I294087,I294095,I294112,I293809,I294143,I749737,I749752,I294160,I294186,I294194,I293797,I293815,I294239,I749758,I294256,I293818,I293803,I293812,I293821,I294359,I1336309,I294385,I294393,I1336288,I294410,I1336315,I294436,I294458,I1336303,I294484,I294492,I1336306,I294509,I294535,I294557,I1336297,I294597,I294614,I294622,I294639,I294670,I1336294,I1336291,I294687,I1336312,I294713,I294721,I294766,I1336300,I294783,I294886,I294912,I294920,I294937,I294963,I294854,I294985,I295011,I295019,I295036,I295062,I294878,I295084,I294860,I295124,I295141,I295149,I295166,I294863,I295197,I295214,I295240,I295248,I294851,I294869,I295293,I295310,I294872,I294857,I294866,I294875,I295413,I1031804,I295439,I295447,I1031801,I1031819,I295464,I1031810,I295490,I295381,I295512,I1031825,I295538,I295546,I1031807,I295563,I295589,I295405,I295611,I295387,I1031813,I295651,I295668,I295676,I295693,I295390,I295724,I1031828,I295741,I1031816,I295767,I295775,I295378,I295396,I295820,I1031822,I295837,I295399,I295384,I295393,I295402,I295940,I1159199,I295966,I295974,I1159214,I295991,I1159217,I296017,I295908,I296039,I1159223,I296065,I296073,I1159205,I296090,I296116,I295932,I296138,I295914,I1159202,I296178,I296195,I296203,I296220,I295917,I296251,I1159208,I296268,I1159220,I296294,I296302,I295905,I295923,I296347,I1159211,I296364,I295926,I295911,I295920,I295929,I296467,I1180007,I296493,I296501,I1180022,I296518,I1180025,I296544,I296566,I1180031,I296592,I296600,I1180013,I296617,I296643,I296665,I1180010,I296705,I296722,I296730,I296747,I296778,I1180016,I296795,I1180028,I296821,I296829,I296874,I1180019,I296891,I296994,I1199081,I297020,I297028,I1199096,I297045,I1199099,I297071,I296962,I297093,I1199105,I297119,I297127,I1199087,I297144,I297170,I296986,I297192,I296968,I1199084,I297232,I297249,I297257,I297274,I296971,I297305,I1199090,I297322,I1199102,I297348,I297356,I296959,I296977,I297401,I1199093,I297418,I296980,I296965,I296974,I296983,I297521,I764199,I297547,I297555,I764190,I764205,I297572,I764211,I297598,I297489,I297620,I764196,I297646,I297654,I297671,I297697,I297513,I297719,I297495,I764193,I297759,I297776,I297784,I297801,I297498,I297832,I764187,I764202,I297849,I297875,I297883,I297486,I297504,I297928,I764208,I297945,I297507,I297492,I297501,I297510,I298048,I1185209,I298074,I298082,I1185224,I298099,I1185227,I298125,I298016,I298147,I1185233,I298173,I298181,I1185215,I298198,I298224,I298040,I298246,I298022,I1185212,I298286,I298303,I298311,I298328,I298025,I298359,I1185218,I298376,I1185230,I298402,I298410,I298013,I298031,I298455,I1185221,I298472,I298034,I298019,I298028,I298037,I298575,I1313778,I298601,I298609,I1313775,I1313766,I298626,I1313763,I298652,I298543,I298674,I1313772,I298700,I298708,I1313781,I298725,I298751,I298567,I298773,I298549,I1313784,I298813,I298830,I298838,I298855,I298552,I298886,I1313769,I298903,I1313787,I298929,I298937,I298540,I298558,I298982,I298999,I298561,I298546,I298555,I298564,I299102,I430030,I299128,I299136,I430042,I430021,I299153,I430045,I299179,I299070,I299201,I430036,I299227,I299235,I430018,I299252,I299278,I299094,I299300,I299076,I430033,I299340,I299357,I299365,I299382,I299079,I299413,I430024,I299430,I430027,I299456,I299464,I299067,I299085,I299509,I430039,I299526,I299088,I299073,I299082,I299091,I299629,I940718,I299655,I299663,I940715,I940733,I299680,I940724,I299706,I299728,I940739,I299754,I299762,I940721,I299779,I299805,I299827,I940727,I299867,I299884,I299892,I299909,I299940,I940742,I299957,I940730,I299983,I299991,I300036,I940736,I300053,I300156,I888001,I300182,I300190,I888004,I887998,I300207,I888010,I300233,I300124,I300255,I888013,I300281,I300289,I300306,I300332,I300148,I300354,I300130,I888016,I300394,I300411,I300419,I300436,I300133,I300467,I888007,I300484,I300510,I300518,I300121,I300139,I300563,I888019,I300580,I300142,I300127,I300136,I300145,I300683,I423502,I300709,I300717,I423514,I423493,I300734,I423517,I300760,I300651,I300782,I423508,I300808,I300816,I423490,I300833,I300859,I300675,I300881,I300657,I423505,I300921,I300938,I300946,I300963,I300660,I300994,I423496,I301011,I423499,I301037,I301045,I300648,I300666,I301090,I423511,I301107,I300669,I300654,I300663,I300672,I301210,I1219311,I301236,I301244,I1219326,I301261,I1219329,I301287,I301178,I301309,I1219335,I301335,I301343,I1219317,I301360,I301386,I301202,I301408,I301184,I1219314,I301448,I301465,I301473,I301490,I301187,I301521,I1219320,I301538,I1219332,I301564,I301572,I301175,I301193,I301617,I1219323,I301634,I301196,I301181,I301190,I301199,I301737,I301763,I301771,I301788,I301814,I301836,I301862,I301870,I301887,I301913,I301935,I301975,I301992,I302000,I302017,I302048,I302065,I302091,I302099,I302144,I302161,I302264,I1152841,I302290,I302298,I1152856,I302315,I1152859,I302341,I302363,I1152865,I302389,I302397,I1152847,I302414,I302440,I302462,I1152844,I302502,I302519,I302527,I302544,I302575,I1152850,I302592,I1152862,I302618,I302626,I302671,I1152853,I302688,I302791,I1278523,I302817,I302825,I1278505,I1278529,I302842,I1278520,I302868,I302759,I302890,I1278526,I302916,I302924,I1278514,I302941,I302967,I302783,I302989,I302765,I303029,I303046,I303054,I303071,I302768,I303102,I1278511,I1278508,I303119,I1278517,I303145,I303153,I302756,I302774,I303198,I303215,I302777,I302762,I302771,I302780,I303318,I938780,I303344,I303352,I938777,I938795,I303369,I938786,I303395,I303286,I303417,I938801,I303443,I303451,I938783,I303468,I303494,I303310,I303516,I303292,I938789,I303556,I303573,I303581,I303598,I303295,I303629,I938804,I303646,I938792,I303672,I303680,I303283,I303301,I303725,I938798,I303742,I303304,I303289,I303298,I303307,I303845,I303871,I303879,I303896,I303922,I303813,I303944,I303970,I303978,I303995,I304021,I303837,I304043,I303819,I304083,I304100,I304108,I304125,I303822,I304156,I304173,I304199,I304207,I303810,I303828,I304252,I304269,I303831,I303816,I303825,I303834,I304372,I498030,I304398,I304406,I498042,I498021,I304423,I498045,I304449,I304340,I304471,I498036,I304497,I304505,I498018,I304522,I304548,I304364,I304570,I304346,I498033,I304610,I304627,I304635,I304652,I304349,I304683,I498024,I304700,I498027,I304726,I304734,I304337,I304355,I304779,I498039,I304796,I304358,I304343,I304352,I304361,I304899,I761309,I304925,I304933,I761300,I761315,I304950,I761321,I304976,I304867,I304998,I761306,I305024,I305032,I305049,I305075,I304891,I305097,I304873,I761303,I305137,I305154,I305162,I305179,I304876,I305210,I761297,I761312,I305227,I305253,I305261,I304864,I304882,I305306,I761318,I305323,I304885,I304870,I304879,I304888,I305426,I305452,I305460,I305477,I305503,I305394,I305525,I305551,I305559,I305576,I305602,I305418,I305624,I305400,I305664,I305681,I305689,I305706,I305403,I305737,I305754,I305780,I305788,I305391,I305409,I305833,I305850,I305412,I305397,I305406,I305415,I305953,I305979,I305987,I306004,I306030,I305921,I306052,I306078,I306086,I306103,I306129,I305945,I306151,I305927,I306191,I306208,I306216,I306233,I305930,I306264,I306281,I306307,I306315,I305918,I305936,I306360,I306377,I305939,I305924,I305933,I305942,I306480,I685013,I306506,I306514,I685004,I685019,I306531,I685025,I306557,I306579,I685010,I306605,I306613,I306630,I306656,I306678,I685007,I306718,I306735,I306743,I306760,I306791,I685001,I685016,I306808,I306834,I306842,I306887,I685022,I306904,I307007,I612766,I307033,I307041,I612751,I612754,I307058,I612769,I307084,I307106,I612763,I307132,I307140,I307157,I307183,I307205,I612760,I307245,I307262,I307270,I307287,I307318,I612775,I307335,I612772,I307361,I307369,I307414,I612757,I307431,I307534,I307560,I307568,I307585,I307611,I307633,I307659,I307667,I307684,I307710,I307732,I307772,I307789,I307797,I307814,I307845,I307862,I307888,I307896,I307941,I307958,I308061,I1122207,I308087,I308095,I1122222,I308112,I1122225,I308138,I308029,I308160,I1122231,I308186,I308194,I1122213,I308211,I308237,I308053,I308259,I308035,I1122210,I308299,I308316,I308324,I308341,I308038,I308372,I1122216,I308389,I1122228,I308415,I308423,I308026,I308044,I308468,I1122219,I308485,I308047,I308032,I308041,I308050,I308588,I527499,I308614,I308622,I527511,I308639,I527496,I308665,I308687,I527520,I308713,I308721,I527517,I308738,I308764,I308786,I527508,I308826,I308843,I308851,I308868,I308899,I527505,I308916,I527514,I308942,I308950,I308995,I527502,I309012,I309115,I309141,I309149,I309166,I309192,I309083,I309214,I309240,I309248,I309265,I309291,I309107,I309313,I309089,I309353,I309370,I309378,I309395,I309092,I309426,I309443,I309469,I309477,I309080,I309098,I309522,I309539,I309101,I309086,I309095,I309104,I309642,I1405924,I309668,I309676,I1405903,I309693,I1405930,I309719,I309610,I309741,I1405918,I309767,I309775,I1405921,I309792,I309818,I309634,I309840,I309616,I1405912,I309880,I309897,I309905,I309922,I309619,I309953,I1405909,I1405906,I309970,I1405927,I309996,I310004,I309607,I309625,I310049,I1405915,I310066,I309628,I309613,I309622,I309631,I310169,I310195,I310203,I310220,I310246,I310137,I310268,I310294,I310302,I310319,I310345,I310161,I310367,I310143,I310407,I310424,I310432,I310449,I310146,I310480,I310497,I310523,I310531,I310134,I310152,I310576,I310593,I310155,I310140,I310149,I310158,I310696,I659581,I310722,I310730,I659572,I659587,I310747,I659593,I310773,I310664,I310795,I659578,I310821,I310829,I310846,I310872,I310688,I310894,I310670,I659575,I310934,I310951,I310959,I310976,I310673,I311007,I659569,I659584,I311024,I311050,I311058,I310661,I310679,I311103,I659590,I311120,I310682,I310667,I310676,I310685,I311223,I879042,I311249,I311257,I879045,I879039,I311274,I879051,I311300,I311191,I311322,I879054,I311348,I311356,I311373,I311399,I311215,I311421,I311197,I879057,I311461,I311478,I311486,I311503,I311200,I311534,I879048,I311551,I311577,I311585,I311188,I311206,I311630,I879060,I311647,I311209,I311194,I311203,I311212,I311750,I1103711,I311776,I311784,I1103726,I311801,I1103729,I311827,I311849,I1103735,I311875,I311883,I1103717,I311900,I311926,I311948,I1103714,I311988,I312005,I312013,I312030,I312061,I1103720,I312078,I1103732,I312104,I312112,I312157,I1103723,I312174,I312277,I312303,I312311,I312328,I312354,I312245,I312376,I312402,I312410,I312427,I312453,I312269,I312475,I312251,I312515,I312532,I312540,I312557,I312254,I312588,I312605,I312631,I312639,I312242,I312260,I312684,I312701,I312263,I312248,I312257,I312266,I312804,I637620,I312830,I312838,I637605,I637608,I312855,I637623,I312881,I312772,I312903,I637617,I312929,I312937,I312954,I312980,I312796,I313002,I312778,I637614,I313042,I313059,I313067,I313084,I312781,I313115,I637629,I313132,I637626,I313158,I313166,I312769,I312787,I313211,I637611,I313228,I312790,I312775,I312784,I312793,I313331,I984646,I313357,I313365,I984643,I984661,I313382,I984652,I313408,I313299,I313430,I984667,I313456,I313464,I984649,I313481,I313507,I313323,I313529,I313305,I984655,I313569,I313586,I313594,I313611,I313308,I313642,I984670,I313659,I984658,I313685,I313693,I313296,I313314,I313738,I984664,I313755,I313317,I313302,I313311,I313320,I313858,I313884,I313892,I313909,I313935,I313957,I313983,I313991,I314008,I314034,I314056,I314096,I314113,I314121,I314138,I314169,I314186,I314212,I314220,I314265,I314282,I314385,I495310,I314411,I314419,I495322,I495301,I314436,I495325,I314462,I314353,I314484,I495316,I314510,I314518,I495298,I314535,I314561,I314377,I314583,I314359,I495313,I314623,I314640,I314648,I314665,I314362,I314696,I495304,I314713,I495307,I314739,I314747,I314350,I314368,I314792,I495319,I314809,I314371,I314356,I314365,I314374,I314912,I1168447,I314938,I314946,I1168462,I314963,I1168465,I314989,I314880,I315011,I1168471,I315037,I315045,I1168453,I315062,I315088,I314904,I315110,I314886,I1168450,I315150,I315167,I315175,I315192,I314889,I315223,I1168456,I315240,I1168468,I315266,I315274,I314877,I314895,I315319,I1168459,I315336,I314898,I314883,I314892,I314901,I315439,I947824,I315465,I315473,I947821,I947839,I315490,I947830,I315516,I315407,I315538,I947845,I315564,I315572,I947827,I315589,I315615,I315431,I315637,I315413,I947833,I315677,I315694,I315702,I315719,I315416,I315750,I947848,I315767,I947836,I315793,I315801,I315404,I315422,I315846,I947842,I315863,I315425,I315410,I315419,I315428,I315966,I847422,I315992,I316000,I847425,I847419,I316017,I847431,I316043,I315934,I316065,I847434,I316091,I316099,I316116,I316142,I315958,I316164,I315940,I847437,I316204,I316221,I316229,I316246,I315943,I316277,I847428,I316294,I316320,I316328,I315931,I315949,I316373,I847440,I316390,I315952,I315937,I315946,I315955,I316493,I954284,I316519,I316527,I954281,I954299,I316544,I954290,I316570,I316592,I954305,I316618,I316626,I954287,I316643,I316669,I316691,I954293,I316731,I316748,I316756,I316773,I316804,I954308,I316821,I954296,I316847,I316855,I316900,I954302,I316917,I317020,I875880,I317046,I317054,I875883,I875877,I317071,I875889,I317097,I316988,I317119,I875892,I317145,I317153,I317170,I317196,I317012,I317218,I316994,I875895,I317258,I317275,I317283,I317300,I316997,I317331,I875886,I317348,I317374,I317382,I316985,I317003,I317427,I875898,I317444,I317006,I316991,I317000,I317009,I317547,I1006610,I317573,I317581,I1006607,I1006625,I317598,I1006616,I317624,I317515,I317646,I1006631,I317672,I317680,I1006613,I317697,I317723,I317539,I317745,I317521,I1006619,I317785,I317802,I317810,I317827,I317524,I317858,I1006634,I317875,I1006622,I317901,I317909,I317512,I317530,I317954,I1006628,I317971,I317533,I317518,I317527,I317536,I318074,I318100,I318108,I318125,I318151,I318042,I318173,I318199,I318207,I318224,I318250,I318066,I318272,I318048,I318312,I318329,I318337,I318354,I318051,I318385,I318402,I318428,I318436,I318039,I318057,I318481,I318498,I318060,I318045,I318054,I318063,I318601,I1366654,I318627,I318635,I1366633,I318652,I1366660,I318678,I318569,I318700,I1366648,I318726,I318734,I1366651,I318751,I318777,I318593,I318799,I318575,I1366642,I318839,I318856,I318864,I318881,I318578,I318912,I1366639,I1366636,I318929,I1366657,I318955,I318963,I318566,I318584,I319008,I1366645,I319025,I318587,I318572,I318581,I318590,I319128,I319154,I319162,I319179,I319205,I319096,I319227,I319253,I319261,I319278,I319304,I319120,I319326,I319102,I319366,I319383,I319391,I319408,I319105,I319439,I319456,I319482,I319490,I319093,I319111,I319535,I319552,I319114,I319099,I319108,I319117,I319655,I932966,I319681,I319689,I932963,I932981,I319706,I932972,I319732,I319623,I319754,I932987,I319780,I319788,I932969,I319805,I319831,I319647,I319853,I319629,I932975,I319893,I319910,I319918,I319935,I319632,I319966,I932990,I319983,I932978,I320009,I320017,I319620,I319638,I320062,I932984,I320079,I319641,I319626,I319635,I319644,I320182,I320208,I320216,I320233,I320259,I320150,I320281,I320307,I320315,I320332,I320358,I320174,I320380,I320156,I320420,I320437,I320445,I320462,I320159,I320493,I320510,I320536,I320544,I320147,I320165,I320589,I320606,I320168,I320153,I320162,I320171,I320709,I616234,I320735,I320743,I616219,I616222,I320760,I616237,I320786,I320677,I320808,I616231,I320834,I320842,I320859,I320885,I320701,I320907,I320683,I616228,I320947,I320964,I320972,I320989,I320686,I321020,I616243,I321037,I616240,I321063,I321071,I320674,I320692,I321116,I616225,I321133,I320695,I320680,I320689,I320698,I321236,I576289,I321262,I321270,I576301,I321287,I576286,I321313,I321204,I321335,I576310,I321361,I321369,I576307,I321386,I321412,I321228,I321434,I321210,I576298,I321474,I321491,I321499,I321516,I321213,I321547,I576295,I321564,I576304,I321590,I321598,I321201,I321219,I321643,I576292,I321660,I321222,I321207,I321216,I321225,I321763,I1241275,I321789,I321797,I1241290,I321814,I1241293,I321840,I321862,I1241299,I321888,I321896,I1241281,I321913,I321939,I321961,I1241278,I322001,I322018,I322026,I322043,I322074,I1241284,I322091,I1241296,I322117,I322125,I322170,I1241287,I322187,I322290,I322316,I322324,I322341,I322367,I322258,I322389,I322415,I322423,I322440,I322466,I322282,I322488,I322264,I322528,I322545,I322553,I322570,I322267,I322601,I322618,I322644,I322652,I322255,I322273,I322697,I322714,I322276,I322261,I322270,I322279,I322817,I1325850,I322843,I322851,I1325877,I1325853,I322868,I1325862,I322894,I322916,I322942,I322950,I1325874,I322967,I322993,I323015,I1325856,I323055,I323072,I323080,I323097,I323128,I1325871,I1325859,I323145,I1325865,I323171,I323179,I323224,I1325868,I323241,I323344,I899595,I323370,I323378,I899598,I899592,I323395,I899604,I323421,I323312,I323443,I899607,I323469,I323477,I323494,I323520,I323336,I323542,I323318,I899610,I323582,I323599,I323607,I323624,I323321,I323655,I899601,I323672,I323698,I323706,I323309,I323327,I323751,I899613,I323768,I323330,I323315,I323324,I323333,I323871,I323897,I323905,I323922,I323948,I323839,I323970,I323996,I324004,I324021,I324047,I323863,I324069,I323845,I324109,I324126,I324134,I324151,I323848,I324182,I324199,I324225,I324233,I323836,I323854,I324278,I324295,I323857,I323842,I323851,I323860,I324398,I324424,I324432,I324449,I324475,I324366,I324497,I324523,I324531,I324548,I324574,I324390,I324596,I324372,I324636,I324653,I324661,I324678,I324375,I324709,I324726,I324752,I324760,I324363,I324381,I324805,I324822,I324384,I324369,I324378,I324387,I324925,I1399974,I324951,I324959,I1399953,I324976,I1399980,I325002,I324893,I325024,I1399968,I325050,I325058,I1399971,I325075,I325101,I324917,I325123,I324899,I1399962,I325163,I325180,I325188,I325205,I324902,I325236,I1399959,I1399956,I325253,I1399977,I325279,I325287,I324890,I324908,I325332,I1399965,I325349,I324911,I324896,I324905,I324914,I325452,I565579,I325478,I325486,I565591,I325503,I565576,I325529,I325420,I325551,I565600,I325577,I325585,I565597,I325602,I325628,I325444,I325650,I325426,I565588,I325690,I325707,I325715,I325732,I325429,I325763,I565585,I325780,I565594,I325806,I325814,I325417,I325435,I325859,I565582,I325876,I325438,I325423,I325432,I325441,I325979,I1112381,I326005,I326013,I1112396,I326030,I1112399,I326056,I325947,I326078,I1112405,I326104,I326112,I1112387,I326129,I326155,I325971,I326177,I325953,I1112384,I326217,I326234,I326242,I326259,I325956,I326290,I1112390,I326307,I1112402,I326333,I326341,I325944,I325962,I326386,I1112393,I326403,I325965,I325950,I325959,I325968,I326506,I488782,I326532,I326540,I488794,I488773,I326557,I488797,I326583,I326474,I326605,I488788,I326631,I326639,I488770,I326656,I326682,I326498,I326704,I326480,I488785,I326744,I326761,I326769,I326786,I326483,I326817,I488776,I326834,I488779,I326860,I326868,I326471,I326489,I326913,I488791,I326930,I326492,I326477,I326486,I326495,I327033,I1196769,I327059,I327067,I1196784,I327084,I1196787,I327110,I327132,I1196793,I327158,I327166,I1196775,I327183,I327209,I327231,I1196772,I327271,I327288,I327296,I327313,I327344,I1196778,I327361,I1196790,I327387,I327395,I327440,I1196781,I327457,I327560,I1180585,I327586,I327594,I1180600,I327611,I1180603,I327637,I327659,I1180609,I327685,I327693,I1180591,I327710,I327736,I327758,I1180588,I327798,I327815,I327823,I327840,I327871,I1180594,I327888,I1180606,I327914,I327922,I327967,I1180597,I327984,I328087,I1170181,I328113,I328121,I1170196,I328138,I1170199,I328164,I328055,I328186,I1170205,I328212,I328220,I1170187,I328237,I328263,I328079,I328285,I328061,I1170184,I328325,I328342,I328350,I328367,I328064,I328398,I1170190,I328415,I1170202,I328441,I328449,I328052,I328070,I328494,I1170193,I328511,I328073,I328058,I328067,I328076,I328614,I473550,I328640,I328648,I473562,I473541,I328665,I473565,I328691,I328713,I473556,I328739,I328747,I473538,I328764,I328790,I328812,I473553,I328852,I328869,I328877,I328894,I328925,I473544,I328942,I473547,I328968,I328976,I329021,I473559,I329038,I329141,I660737,I329167,I329175,I660728,I660743,I329192,I660749,I329218,I329240,I660734,I329266,I329274,I329291,I329317,I329339,I660731,I329379,I329396,I329404,I329421,I329452,I660725,I660740,I329469,I329495,I329503,I329548,I660746,I329565,I329668,I329694,I329702,I329719,I329745,I329636,I329767,I329793,I329801,I329818,I329844,I329660,I329866,I329642,I329906,I329923,I329931,I329948,I329645,I329979,I329996,I330022,I330030,I329633,I329651,I330075,I330092,I329654,I329639,I329648,I329657,I330195,I1150529,I330221,I330229,I1150544,I330246,I1150547,I330272,I330163,I330294,I1150553,I330320,I330328,I1150535,I330345,I330371,I330187,I330393,I330169,I1150532,I330433,I330450,I330458,I330475,I330172,I330506,I1150538,I330523,I1150550,I330549,I330557,I330160,I330178,I330602,I1150541,I330619,I330181,I330166,I330175,I330184,I330722,I330748,I330756,I330773,I330799,I330690,I330821,I330847,I330855,I330872,I330898,I330714,I330920,I330696,I330960,I330977,I330985,I331002,I330699,I331033,I331050,I331076,I331084,I330687,I330705,I331129,I331146,I330708,I330693,I330702,I330711,I331249,I844260,I331275,I331283,I844263,I844257,I331300,I844269,I331326,I331217,I331348,I844272,I331374,I331382,I331399,I331425,I331241,I331447,I331223,I844275,I331487,I331504,I331512,I331529,I331226,I331560,I844266,I331577,I331603,I331611,I331214,I331232,I331656,I844278,I331673,I331235,I331220,I331229,I331238,I331776,I851638,I331802,I331810,I851641,I851635,I331827,I851647,I331853,I331875,I851650,I331901,I331909,I331926,I331952,I331974,I851653,I332014,I332031,I332039,I332056,I332087,I851644,I332104,I332130,I332138,I332183,I851656,I332200,I332303,I332329,I332337,I332354,I332380,I332271,I332402,I332428,I332436,I332453,I332479,I332295,I332501,I332277,I332541,I332558,I332566,I332583,I332280,I332614,I332631,I332657,I332665,I332268,I332286,I332710,I332727,I332289,I332274,I332283,I332292,I332830,I909081,I332856,I332864,I909084,I909078,I332881,I909090,I332907,I332929,I909093,I332955,I332963,I332980,I333006,I333028,I909096,I333068,I333085,I333093,I333110,I333141,I909087,I333158,I333184,I333192,I333237,I909099,I333254,I333357,I1040202,I333383,I333391,I1040199,I1040217,I333408,I1040208,I333434,I333325,I333456,I1040223,I333482,I333490,I1040205,I333507,I333533,I333349,I333555,I333331,I1040211,I333595,I333612,I333620,I333637,I333334,I333668,I1040226,I333685,I1040214,I333711,I333719,I333322,I333340,I333764,I1040220,I333781,I333343,I333328,I333337,I333346,I333884,I333910,I333918,I333935,I333961,I333983,I334009,I334017,I334034,I334060,I334082,I334122,I334139,I334147,I334164,I334195,I334212,I334238,I334246,I334291,I334308,I334411,I450158,I334437,I334445,I450170,I450149,I334462,I450173,I334488,I334379,I334510,I450164,I334536,I334544,I450146,I334561,I334587,I334403,I334609,I334385,I450161,I334649,I334666,I334674,I334691,I334388,I334722,I450152,I334739,I450155,I334765,I334773,I334376,I334394,I334818,I450167,I334835,I334397,I334382,I334391,I334400,I334938,I1402949,I334964,I334972,I1402928,I334989,I1402955,I335015,I335037,I1402943,I335063,I335071,I1402946,I335088,I335114,I335136,I1402937,I335176,I335193,I335201,I335218,I335249,I1402934,I1402931,I335266,I1402952,I335292,I335300,I335345,I1402940,I335362,I335465,I1371414,I335491,I335499,I1371393,I335516,I1371420,I335542,I335433,I335564,I1371408,I335590,I335598,I1371411,I335615,I335641,I335457,I335663,I335439,I1371402,I335703,I335720,I335728,I335745,I335442,I335776,I1371399,I1371396,I335793,I1371417,I335819,I335827,I335430,I335448,I335872,I1371405,I335889,I335451,I335436,I335445,I335454,I335992,I336018,I336026,I336043,I336069,I335960,I336091,I336117,I336125,I336142,I336168,I335984,I336190,I335966,I336230,I336247,I336255,I336272,I335969,I336303,I336320,I336346,I336354,I335957,I335975,I336399,I336416,I335978,I335963,I335972,I335981,I336519,I1071346,I336545,I336553,I1071343,I336570,I1071355,I336596,I336618,I336644,I336652,I1071361,I336669,I336695,I336717,I1071349,I336757,I336774,I336782,I336799,I336830,I1071358,I1071364,I336847,I336873,I336881,I336926,I1071352,I336943,I337046,I806971,I337072,I337080,I806962,I806977,I337097,I806983,I337123,I337014,I337145,I806968,I337171,I337179,I337196,I337222,I337038,I337244,I337020,I806965,I337284,I337301,I337309,I337326,I337023,I337357,I806959,I806974,I337374,I337400,I337408,I337011,I337029,I337453,I806980,I337470,I337032,I337017,I337026,I337035,I337573,I1022760,I337599,I337607,I1022757,I1022775,I337624,I1022766,I337650,I337672,I1022781,I337698,I337706,I1022763,I337723,I337749,I337771,I1022769,I337811,I337828,I337836,I337853,I337884,I1022784,I337901,I1022772,I337927,I337935,I337980,I1022778,I337997,I338100,I624326,I338126,I338134,I624311,I624314,I338151,I624329,I338177,I338068,I338199,I624323,I338225,I338233,I338250,I338276,I338092,I338298,I338074,I624320,I338338,I338355,I338363,I338380,I338077,I338411,I624335,I338428,I624332,I338454,I338462,I338065,I338083,I338507,I624317,I338524,I338086,I338071,I338080,I338089,I338627,I338653,I338661,I338678,I338704,I338595,I338726,I338752,I338760,I338777,I338803,I338619,I338825,I338601,I338865,I338882,I338890,I338907,I338604,I338938,I338955,I338981,I338989,I338592,I338610,I339034,I339051,I338613,I338598,I338607,I338616,I339154,I768245,I339180,I339188,I768236,I768251,I339205,I768257,I339231,I339122,I339253,I768242,I339279,I339287,I339304,I339330,I339146,I339352,I339128,I768239,I339392,I339409,I339417,I339434,I339131,I339465,I768233,I768248,I339482,I339508,I339516,I339119,I339137,I339561,I768254,I339578,I339140,I339125,I339134,I339143,I339681,I1097353,I339707,I339715,I1097368,I339732,I1097371,I339758,I339649,I339780,I1097377,I339806,I339814,I1097359,I339831,I339857,I339673,I339879,I339655,I1097356,I339919,I339936,I339944,I339961,I339658,I339992,I1097362,I340009,I1097374,I340035,I340043,I339646,I339664,I340088,I1097365,I340105,I339667,I339652,I339661,I339670,I340208,I340234,I340242,I340259,I340285,I340176,I340307,I340333,I340341,I340358,I340384,I340200,I340406,I340182,I340446,I340463,I340471,I340488,I340185,I340519,I340536,I340562,I340570,I340173,I340191,I340615,I340632,I340194,I340179,I340188,I340197,I340735,I1229715,I340761,I340769,I1229730,I340786,I1229733,I340812,I340703,I340834,I1229739,I340860,I340868,I1229721,I340885,I340911,I340727,I340933,I340709,I1229718,I340973,I340990,I340998,I341015,I340712,I341046,I1229724,I341063,I1229736,I341089,I341097,I340700,I340718,I341142,I1229727,I341159,I340721,I340706,I340715,I340724,I341262,I1211219,I341288,I341296,I1211234,I341313,I1211237,I341339,I341361,I1211243,I341387,I341395,I1211225,I341412,I341438,I341460,I1211222,I341500,I341517,I341525,I341542,I341573,I1211228,I341590,I1211240,I341616,I341624,I341669,I1211231,I341686,I341789,I802347,I341815,I341823,I802338,I802353,I341840,I802359,I341866,I341888,I802344,I341914,I341922,I341939,I341965,I341987,I802341,I342027,I342044,I342052,I342069,I342100,I802335,I802350,I342117,I342143,I342151,I342196,I802356,I342213,I342316,I342342,I342350,I342367,I342393,I342415,I342441,I342449,I342466,I342492,I342514,I342554,I342571,I342579,I342596,I342627,I342644,I342670,I342678,I342723,I342740,I342843,I342869,I342877,I342894,I342920,I342942,I342968,I342976,I342993,I343019,I343041,I343081,I343098,I343106,I343123,I343154,I343171,I343197,I343205,I343250,I343267,I343370,I582132,I343396,I343404,I582117,I582120,I343421,I582135,I343447,I343338,I343469,I582129,I343495,I343503,I343520,I343546,I343362,I343568,I343344,I582126,I343608,I343625,I343633,I343650,I343347,I343681,I582141,I343698,I582138,I343724,I343732,I343335,I343353,I343777,I582123,I343794,I343356,I343341,I343350,I343359,I343897,I1353564,I343923,I343931,I1353543,I343948,I1353570,I343974,I343865,I343996,I1353558,I344022,I344030,I1353561,I344047,I344073,I343889,I344095,I343871,I1353552,I344135,I344152,I344160,I344177,I343874,I344208,I1353549,I1353546,I344225,I1353567,I344251,I344259,I343862,I343880,I344304,I1353555,I344321,I343883,I343868,I343877,I343886,I344424,I344450,I344458,I344475,I344501,I344392,I344523,I344549,I344557,I344574,I344600,I344416,I344622,I344398,I344662,I344679,I344687,I344704,I344401,I344735,I344752,I344778,I344786,I344389,I344407,I344831,I344848,I344410,I344395,I344404,I344413,I344951,I344977,I344985,I345002,I345028,I344919,I345050,I345076,I345084,I345101,I345127,I344943,I345149,I344925,I345189,I345206,I345214,I345231,I344928,I345262,I345279,I345305,I345313,I344916,I344934,I345358,I345375,I344937,I344922,I344931,I344940,I345478,I1352374,I345504,I345512,I1352353,I345529,I1352380,I345555,I345446,I345577,I1352368,I345603,I345611,I1352371,I345628,I345654,I345470,I345676,I345452,I1352362,I345716,I345733,I345741,I345758,I345455,I345789,I1352359,I1352356,I345806,I1352377,I345832,I345840,I345443,I345461,I345885,I1352365,I345902,I345464,I345449,I345458,I345467,I346005,I874299,I346031,I346039,I874302,I874296,I346056,I874308,I346082,I345973,I346104,I874311,I346130,I346138,I346155,I346181,I345997,I346203,I345979,I874314,I346243,I346260,I346268,I346285,I345982,I346316,I874305,I346333,I346359,I346367,I345970,I345988,I346412,I874317,I346429,I345991,I345976,I345985,I345994,I346532,I980770,I346558,I346566,I980767,I980785,I346583,I980776,I346609,I346500,I346631,I980791,I346657,I346665,I980773,I346682,I346708,I346524,I346730,I346506,I980779,I346770,I346787,I346795,I346812,I346509,I346843,I980794,I346860,I980782,I346886,I346894,I346497,I346515,I346939,I980788,I346956,I346518,I346503,I346512,I346521,I347059,I1172493,I347085,I347093,I1172508,I347110,I1172511,I347136,I347027,I347158,I1172517,I347184,I347192,I1172499,I347209,I347235,I347051,I347257,I347033,I1172496,I347297,I347314,I347322,I347339,I347036,I347370,I1172502,I347387,I1172514,I347413,I347421,I347024,I347042,I347466,I1172505,I347483,I347045,I347030,I347039,I347048,I347586,I347612,I347620,I347637,I347663,I347554,I347685,I347711,I347719,I347736,I347762,I347578,I347784,I347560,I347824,I347841,I347849,I347866,I347563,I347897,I347914,I347940,I347948,I347551,I347569,I347993,I348010,I347572,I347557,I347566,I347575,I348113,I1060687,I348139,I348147,I1060684,I348164,I1060696,I348190,I348081,I348212,I348238,I348246,I1060702,I348263,I348289,I348105,I348311,I348087,I1060690,I348351,I348368,I348376,I348393,I348090,I348424,I1060699,I1060705,I348441,I348467,I348475,I348078,I348096,I348520,I1060693,I348537,I348099,I348084,I348093,I348102,I348640,I1068541,I348666,I348674,I1068538,I348691,I1068550,I348717,I348608,I348739,I348765,I348773,I1068556,I348790,I348816,I348632,I348838,I348614,I1068544,I348878,I348895,I348903,I348920,I348617,I348951,I1068553,I1068559,I348968,I348994,I349002,I348605,I348623,I349047,I1068547,I349064,I348626,I348611,I348620,I348629,I349167,I507278,I349193,I349201,I507290,I507269,I349218,I507293,I349244,I349135,I349266,I507284,I349292,I349300,I507266,I349317,I349343,I349159,I349365,I349141,I507281,I349405,I349422,I349430,I349447,I349144,I349478,I507272,I349495,I507275,I349521,I349529,I349132,I349150,I349574,I507287,I349591,I349153,I349138,I349147,I349156,I349694,I864286,I349720,I349728,I864289,I864283,I349745,I864295,I349771,I349662,I349793,I864298,I349819,I349827,I349844,I349870,I349686,I349892,I349668,I864301,I349932,I349949,I349957,I349974,I349671,I350005,I864292,I350022,I350048,I350056,I349659,I349677,I350101,I864304,I350118,I349680,I349665,I349674,I349683,I350221,I613344,I350247,I350255,I613329,I613332,I350272,I613347,I350298,I350320,I613341,I350346,I350354,I350371,I350397,I350419,I613338,I350459,I350476,I350484,I350501,I350532,I613353,I350549,I613350,I350575,I350583,I350628,I613335,I350645,I350748,I1290080,I350774,I350782,I1290077,I1290068,I350799,I1290065,I350825,I350716,I350847,I1290074,I350873,I350881,I1290083,I350898,I350924,I350740,I350946,I350722,I1290086,I350986,I351003,I351011,I351028,I350725,I351059,I1290071,I351076,I1290089,I351102,I351110,I350713,I350731,I351155,I351172,I350734,I350719,I350728,I350737,I351275,I779227,I351301,I351309,I779218,I779233,I351326,I779239,I351352,I351243,I351374,I779224,I351400,I351408,I351425,I351451,I351267,I351473,I351249,I779221,I351513,I351530,I351538,I351555,I351252,I351586,I779215,I779230,I351603,I351629,I351637,I351240,I351258,I351682,I779236,I351699,I351261,I351246,I351255,I351264,I351802,I618546,I351828,I351836,I618531,I618534,I351853,I618549,I351879,I351770,I351901,I618543,I351927,I351935,I351952,I351978,I351794,I352000,I351776,I618540,I352040,I352057,I352065,I352082,I351779,I352113,I618555,I352130,I618552,I352156,I352164,I351767,I351785,I352209,I618537,I352226,I351788,I351773,I351782,I351791,I352329,I1054516,I352355,I352363,I1054513,I352380,I1054525,I352406,I352297,I352428,I352454,I352462,I1054531,I352479,I352505,I352321,I352527,I352303,I1054519,I352567,I352584,I352592,I352609,I352306,I352640,I1054528,I1054534,I352657,I352683,I352691,I352294,I352312,I352736,I1054522,I352753,I352315,I352300,I352309,I352318,I352856,I1177117,I352882,I352890,I1177132,I352907,I1177135,I352933,I352824,I352955,I1177141,I352981,I352989,I1177123,I353006,I353032,I352848,I353054,I352830,I1177120,I353094,I353111,I353119,I353136,I352833,I353167,I1177126,I353184,I1177138,I353210,I353218,I352821,I352839,I353263,I1177129,I353280,I352842,I352827,I352836,I352845,I353383,I1109491,I353409,I353417,I1109506,I353434,I1109509,I353460,I353482,I1109515,I353508,I353516,I1109497,I353533,I353559,I353581,I1109494,I353621,I353638,I353646,I353663,I353694,I1109500,I353711,I1109512,I353737,I353745,I353790,I1109503,I353807,I353910,I596004,I353936,I353944,I595989,I595992,I353961,I596007,I353987,I354009,I596001,I354035,I354043,I354060,I354086,I354108,I595998,I354148,I354165,I354173,I354190,I354221,I596013,I354238,I596010,I354264,I354272,I354317,I595995,I354334,I354437,I354463,I354471,I354488,I354514,I354405,I354536,I354562,I354570,I354587,I354613,I354429,I354635,I354411,I354675,I354692,I354700,I354717,I354414,I354748,I354765,I354791,I354799,I354402,I354420,I354844,I354861,I354423,I354408,I354417,I354426,I354964,I354990,I354998,I355015,I355041,I355063,I355089,I355097,I355114,I355140,I355162,I355202,I355219,I355227,I355244,I355275,I355292,I355318,I355326,I355371,I355388,I355491,I355517,I355525,I355542,I355568,I355459,I355590,I355616,I355624,I355641,I355667,I355483,I355689,I355465,I355729,I355746,I355754,I355771,I355468,I355802,I355819,I355845,I355853,I355456,I355474,I355898,I355915,I355477,I355462,I355471,I355480,I356018,I774025,I356044,I356052,I774016,I774031,I356069,I774037,I356095,I355986,I356117,I774022,I356143,I356151,I356168,I356194,I356010,I356216,I355992,I774019,I356256,I356273,I356281,I356298,I355995,I356329,I774013,I774028,I356346,I356372,I356380,I355983,I356001,I356425,I774034,I356442,I356004,I355989,I355998,I356007,I356545,I1090995,I356571,I356579,I1091010,I356596,I1091013,I356622,I356644,I1091019,I356670,I356678,I1091001,I356695,I356721,I356743,I1090998,I356783,I356800,I356808,I356825,I356856,I1091004,I356873,I1091016,I356899,I356907,I356952,I1091007,I356969,I357072,I787319,I357098,I357106,I787310,I787325,I357123,I787331,I357149,I357171,I787316,I357197,I357205,I357222,I357248,I357270,I787313,I357310,I357327,I357335,I357352,I357383,I787307,I787322,I357400,I357426,I357434,I357479,I787328,I357496,I357599,I1137813,I357625,I357633,I1137828,I357650,I1137831,I357676,I357567,I357698,I1137837,I357724,I357732,I1137819,I357749,I357775,I357591,I357797,I357573,I1137816,I357837,I357854,I357862,I357879,I357576,I357910,I1137822,I357927,I1137834,I357953,I357961,I357564,I357582,I358006,I1137825,I358023,I357585,I357570,I357579,I357588,I358126,I1135501,I358152,I358160,I1135516,I358177,I1135519,I358203,I358094,I358225,I1135525,I358251,I358259,I1135507,I358276,I358302,I358118,I358324,I358100,I1135504,I358364,I358381,I358389,I358406,I358103,I358437,I1135510,I358454,I1135522,I358480,I358488,I358091,I358109,I358533,I1135513,I358550,I358112,I358097,I358106,I358115,I358653,I358679,I358687,I358704,I358730,I358752,I358778,I358786,I358803,I358829,I358851,I358891,I358908,I358916,I358933,I358964,I358981,I359007,I359015,I359060,I359077,I359180,I543564,I359206,I359214,I543576,I359231,I543561,I359257,I359148,I359279,I543585,I359305,I359313,I543582,I359330,I359356,I359172,I359378,I359154,I543573,I359418,I359435,I359443,I359460,I359157,I359491,I543570,I359508,I543579,I359534,I359542,I359145,I359163,I359587,I543567,I359604,I359166,I359151,I359160,I359169,I359707,I868502,I359733,I359741,I868505,I868499,I359758,I868511,I359784,I359675,I359806,I868514,I359832,I359840,I359857,I359883,I359699,I359905,I359681,I868517,I359945,I359962,I359970,I359987,I359684,I360018,I868508,I360035,I360061,I360069,I359672,I359690,I360114,I868520,I360131,I359693,I359678,I359687,I359696,I360234,I1404139,I360260,I360268,I1404118,I360285,I1404145,I360311,I360202,I360333,I1404133,I360359,I360367,I1404136,I360384,I360410,I360226,I360432,I360208,I1404127,I360472,I360489,I360497,I360514,I360211,I360545,I1404124,I1404121,I360562,I1404142,I360588,I360596,I360199,I360217,I360641,I1404130,I360658,I360220,I360205,I360214,I360223,I360761,I967850,I360787,I360795,I967847,I967865,I360812,I967856,I360838,I360860,I967871,I360886,I360894,I967853,I360911,I360937,I360959,I967859,I360999,I361016,I361024,I361041,I361072,I967874,I361089,I967862,I361115,I361123,I361168,I967868,I361185,I361288,I1080322,I361314,I361322,I1080319,I361339,I1080331,I361365,I361387,I361413,I361421,I1080337,I361438,I361464,I361486,I1080325,I361526,I361543,I361551,I361568,I361599,I1080334,I1080340,I361616,I361642,I361650,I361695,I1080328,I361712,I361815,I956222,I361841,I361849,I956219,I956237,I361866,I956228,I361892,I361914,I956243,I361940,I361948,I956225,I361965,I361991,I362013,I956231,I362053,I362070,I362078,I362095,I362126,I956246,I362143,I956234,I362169,I362177,I362222,I956240,I362239,I362342,I362368,I362376,I362393,I362419,I362441,I362467,I362475,I362492,I362518,I362540,I362580,I362597,I362605,I362622,I362653,I362670,I362696,I362704,I362749,I362766,I362869,I362895,I362903,I362920,I362946,I362968,I362994,I363002,I363019,I363045,I363067,I363107,I363124,I363132,I363149,I363180,I363197,I363223,I363231,I363276,I363293,I363396,I1124519,I363422,I363430,I1124534,I363447,I1124537,I363473,I363364,I363495,I1124543,I363521,I363529,I1124525,I363546,I363572,I363388,I363594,I363370,I1124522,I363634,I363651,I363659,I363676,I363373,I363707,I1124528,I363724,I1124540,I363750,I363758,I363361,I363379,I363803,I1124531,I363820,I363382,I363367,I363376,I363385,I363923,I757841,I363949,I363957,I757832,I757847,I363974,I757853,I364000,I363891,I364022,I757838,I364048,I364056,I364073,I364099,I363915,I364121,I363897,I757835,I364161,I364178,I364186,I364203,I363900,I364234,I757829,I757844,I364251,I364277,I364285,I363888,I363906,I364330,I757850,I364347,I363909,I363894,I363903,I363912,I364450,I981416,I364476,I364484,I981413,I981431,I364501,I981422,I364527,I364549,I981437,I364575,I364583,I981419,I364600,I364626,I364648,I981425,I364688,I364705,I364713,I364730,I364761,I981440,I364778,I981428,I364804,I364812,I364857,I981434,I364874,I364977,I945240,I365003,I365011,I945237,I945255,I365028,I945246,I365054,I364945,I365076,I945261,I365102,I365110,I945243,I365127,I365153,I364969,I365175,I364951,I945249,I365215,I365232,I365240,I365257,I364954,I365288,I945264,I365305,I945252,I365331,I365339,I364942,I364960,I365384,I945258,I365401,I364963,I364948,I364957,I364966,I365504,I365530,I365538,I365555,I365581,I365603,I365629,I365637,I365654,I365680,I365702,I365742,I365759,I365767,I365784,I365815,I365832,I365858,I365866,I365911,I365928,I366031,I1199659,I366057,I366065,I1199674,I366082,I1199677,I366108,I365999,I366130,I1199683,I366156,I366164,I1199665,I366181,I366207,I366023,I366229,I366005,I1199662,I366269,I366286,I366294,I366311,I366008,I366342,I1199668,I366359,I1199680,I366385,I366393,I365996,I366014,I366438,I1199671,I366455,I366017,I366002,I366011,I366020,I366558,I1210641,I366584,I366592,I1210656,I366609,I1210659,I366635,I366526,I366657,I1210665,I366683,I366691,I1210647,I366708,I366734,I366550,I366756,I366532,I1210644,I366796,I366813,I366821,I366838,I366535,I366869,I1210650,I366886,I1210662,I366912,I366920,I366523,I366541,I366965,I1210653,I366982,I366544,I366529,I366538,I366547,I367085,I1282331,I367111,I367119,I1282313,I1282337,I367136,I1282328,I367162,I367053,I367184,I1282334,I367210,I367218,I1282322,I367235,I367261,I367077,I367283,I367059,I367323,I367340,I367348,I367365,I367062,I367396,I1282319,I1282316,I367413,I1282325,I367439,I367447,I367050,I367068,I367492,I367509,I367071,I367056,I367065,I367074,I367612,I679811,I367638,I367646,I679802,I679817,I367663,I679823,I367689,I367580,I367711,I679808,I367737,I367745,I367762,I367788,I367604,I367810,I367586,I679805,I367850,I367867,I367875,I367892,I367589,I367923,I679799,I679814,I367940,I367966,I367974,I367577,I367595,I368019,I679820,I368036,I367598,I367583,I367592,I367601,I368139,I600050,I368165,I368173,I600035,I600038,I368190,I600053,I368216,I368107,I368238,I600047,I368264,I368272,I368289,I368315,I368131,I368337,I368113,I600044,I368377,I368394,I368402,I368419,I368116,I368450,I600059,I368467,I600056,I368493,I368501,I368104,I368122,I368546,I600041,I368563,I368125,I368110,I368119,I368128,I368666,I1170759,I368692,I368700,I1170774,I368717,I1170777,I368743,I368765,I1170783,I368791,I368799,I1170765,I368816,I368842,I368864,I1170762,I368904,I368921,I368929,I368946,I368977,I1170768,I368994,I1170780,I369020,I369028,I369073,I1170771,I369090,I369193,I1218733,I369219,I369227,I1218748,I369244,I1218751,I369270,I369161,I369292,I1218757,I369318,I369326,I1218739,I369343,I369369,I369185,I369391,I369167,I1218736,I369431,I369448,I369456,I369473,I369170,I369504,I1218742,I369521,I1218754,I369547,I369555,I369158,I369176,I369600,I1218745,I369617,I369179,I369164,I369173,I369182,I369720,I713335,I369746,I369754,I713326,I713341,I369771,I713347,I369797,I369688,I369819,I713332,I369845,I369853,I369870,I369896,I369712,I369918,I369694,I713329,I369958,I369975,I369983,I370000,I369697,I370031,I713323,I713338,I370048,I370074,I370082,I369685,I369703,I370127,I713344,I370144,I369706,I369691,I369700,I369709,I370247,I751483,I370273,I370281,I751474,I751489,I370298,I751495,I370324,I370346,I751480,I370372,I370380,I370397,I370423,I370445,I751477,I370485,I370502,I370510,I370527,I370558,I751471,I751486,I370575,I370601,I370609,I370654,I751492,I370671,I370774,I370800,I370808,I370825,I370851,I370742,I370873,I370899,I370907,I370924,I370950,I370766,I370972,I370748,I371012,I371029,I371037,I371054,I370751,I371085,I371102,I371128,I371136,I370739,I370757,I371181,I371198,I370760,I370745,I370754,I370763,I371301,I939426,I371327,I371335,I939423,I939441,I371352,I939432,I371378,I371269,I371400,I939447,I371426,I371434,I939429,I371451,I371477,I371293,I371499,I371275,I939435,I371539,I371556,I371564,I371581,I371278,I371612,I939450,I371629,I939438,I371655,I371663,I371266,I371284,I371708,I939444,I371725,I371287,I371272,I371281,I371290,I371828,I735299,I371854,I371862,I735290,I735305,I371879,I735311,I371905,I371796,I371927,I735296,I371953,I371961,I371978,I372004,I371820,I372026,I371802,I735293,I372066,I372083,I372091,I372108,I371805,I372139,I735287,I735302,I372156,I372182,I372190,I371793,I371811,I372235,I735308,I372252,I371814,I371799,I371808,I371817,I372355,I1123941,I372381,I372389,I1123956,I372406,I1123959,I372432,I372323,I372454,I1123965,I372480,I372488,I1123947,I372505,I372531,I372347,I372553,I372329,I1123944,I372593,I372610,I372618,I372635,I372332,I372666,I1123950,I372683,I1123962,I372709,I372717,I372320,I372338,I372762,I1123953,I372779,I372341,I372326,I372335,I372344,I372882,I372908,I372916,I372933,I372959,I372850,I372981,I373007,I373015,I373032,I373058,I372874,I373080,I372856,I373120,I373137,I373145,I373162,I372859,I373193,I373210,I373236,I373244,I372847,I372865,I373289,I373306,I372868,I372853,I372862,I372871,I373409,I1093307,I373435,I373443,I1093322,I373460,I1093325,I373486,I373377,I373508,I1093331,I373534,I373542,I1093313,I373559,I373585,I373401,I373607,I373383,I1093310,I373647,I373664,I373672,I373689,I373386,I373720,I1093316,I373737,I1093328,I373763,I373771,I373374,I373392,I373816,I1093319,I373833,I373395,I373380,I373389,I373398,I373936,I1373199,I373962,I373970,I1373178,I373987,I1373205,I374013,I373904,I374035,I1373193,I374061,I374069,I1373196,I374086,I374112,I373928,I374134,I373910,I1373187,I374174,I374191,I374199,I374216,I373913,I374247,I1373184,I1373181,I374264,I1373202,I374290,I374298,I373901,I373919,I374343,I1373190,I374360,I373922,I373907,I373916,I373925,I374463,I978832,I374489,I374497,I978829,I978847,I374514,I978838,I374540,I374431,I374562,I978853,I374588,I374596,I978835,I374613,I374639,I374455,I374661,I374437,I978841,I374701,I374718,I374726,I374743,I374440,I374774,I978856,I374791,I978844,I374817,I374825,I374428,I374446,I374870,I978850,I374887,I374449,I374434,I374443,I374452,I374990,I1107179,I375016,I375024,I1107194,I375041,I1107197,I375067,I374958,I375089,I1107203,I375115,I375123,I1107185,I375140,I375166,I374982,I375188,I374964,I1107182,I375228,I375245,I375253,I375270,I374967,I375301,I1107188,I375318,I1107200,I375344,I375352,I374955,I374973,I375397,I1107191,I375414,I374976,I374961,I374970,I374979,I375517,I676343,I375543,I375551,I676334,I676349,I375568,I676355,I375594,I375485,I375616,I676340,I375642,I375650,I375667,I375693,I375509,I375715,I375491,I676337,I375755,I375772,I375780,I375797,I375494,I375828,I676331,I676346,I375845,I375871,I375879,I375482,I375500,I375924,I676352,I375941,I375503,I375488,I375497,I375506,I376044,I678655,I376070,I376078,I678646,I678661,I376095,I678667,I376121,I376012,I376143,I678652,I376169,I376177,I376194,I376220,I376036,I376242,I376018,I678649,I376282,I376299,I376307,I376324,I376021,I376355,I678643,I678658,I376372,I376398,I376406,I376009,I376027,I376451,I678664,I376468,I376030,I376015,I376024,I376033,I376571,I1153997,I376597,I376605,I1154012,I376622,I1154015,I376648,I376539,I376670,I1154021,I376696,I376704,I1154003,I376721,I376747,I376563,I376769,I376545,I1154000,I376809,I376826,I376834,I376851,I376548,I376882,I1154006,I376899,I1154018,I376925,I376933,I376536,I376554,I376978,I1154009,I376995,I376557,I376542,I376551,I376560,I377098,I502926,I377124,I377132,I502938,I502917,I377149,I502941,I377175,I377197,I502932,I377223,I377231,I502914,I377248,I377274,I377296,I502929,I377336,I377353,I377361,I377378,I377409,I502920,I377426,I502923,I377452,I377460,I377505,I502935,I377522,I377625,I825288,I377651,I377659,I825291,I825285,I377676,I825297,I377702,I377593,I377724,I825300,I377750,I377758,I377775,I377801,I377617,I377823,I377599,I825303,I377863,I377880,I377888,I377905,I377602,I377936,I825294,I377953,I377979,I377987,I377590,I377608,I378032,I825306,I378049,I377611,I377596,I377605,I377614,I378152,I945886,I378178,I378186,I945883,I945901,I378203,I945892,I378229,I378120,I378251,I945907,I378277,I378285,I945889,I378302,I378328,I378144,I378350,I378126,I945895,I378390,I378407,I378415,I378432,I378129,I378463,I945910,I378480,I945898,I378506,I378514,I378117,I378135,I378559,I945904,I378576,I378138,I378123,I378132,I378141,I378679,I716803,I378705,I378713,I716794,I716809,I378730,I716815,I378756,I378647,I378778,I716800,I378804,I378812,I378829,I378855,I378671,I378877,I378653,I716797,I378917,I378934,I378942,I378959,I378656,I378990,I716791,I716806,I379007,I379033,I379041,I378644,I378662,I379086,I716812,I379103,I378665,I378650,I378659,I378668,I379206,I461582,I379232,I379240,I461594,I461573,I379257,I461597,I379283,I379305,I461588,I379331,I379339,I461570,I379356,I379382,I379404,I461585,I379444,I379461,I379469,I379486,I379517,I461576,I379534,I461579,I379560,I379568,I379613,I461591,I379630,I379733,I379759,I379767,I379784,I379810,I379832,I379858,I379866,I379883,I379909,I379931,I379971,I379988,I379996,I380013,I380044,I380061,I380087,I380095,I380140,I380157,I380260,I1159777,I380286,I380294,I1159792,I380311,I1159795,I380337,I380359,I1159801,I380385,I380393,I1159783,I380410,I380436,I380458,I1159780,I380498,I380515,I380523,I380540,I380571,I1159786,I380588,I1159798,I380614,I380622,I380667,I1159789,I380684,I380787,I770557,I380813,I380821,I770548,I770563,I380838,I770569,I380864,I380755,I380886,I770554,I380912,I380920,I380937,I380963,I380779,I380985,I380761,I770551,I381025,I381042,I381050,I381067,I380764,I381098,I770545,I770560,I381115,I381141,I381149,I380752,I380770,I381194,I770566,I381211,I380773,I380758,I380767,I380776,I381314,I644556,I381340,I381348,I644541,I644544,I381365,I644559,I381391,I381282,I381413,I644553,I381439,I381447,I381464,I381490,I381306,I381512,I381288,I644550,I381552,I381569,I381577,I381594,I381291,I381625,I644565,I381642,I644562,I381668,I381676,I381279,I381297,I381721,I644547,I381738,I381300,I381285,I381294,I381303,I381841,I381867,I381875,I381892,I381918,I381940,I381966,I381974,I381991,I382017,I382039,I382079,I382096,I382104,I382121,I382152,I382169,I382195,I382203,I382248,I382265,I382368,I493134,I382394,I382402,I493146,I493125,I382419,I493149,I382445,I382336,I382467,I493140,I382493,I382501,I493122,I382518,I382544,I382360,I382566,I382342,I493137,I382606,I382623,I382631,I382648,I382345,I382679,I493128,I382696,I493131,I382722,I382730,I382333,I382351,I382775,I493143,I382792,I382354,I382339,I382348,I382357,I382895,I912243,I382921,I382929,I912246,I912240,I382946,I912252,I382972,I382863,I382994,I912255,I383020,I383028,I383045,I383071,I382887,I383093,I382869,I912258,I383133,I383150,I383158,I383175,I382872,I383206,I912249,I383223,I383249,I383257,I382860,I382878,I383302,I912261,I383319,I382881,I382866,I382875,I382884,I383422,I801769,I383448,I383456,I801760,I801775,I383473,I801781,I383499,I383521,I801766,I383547,I383555,I383572,I383598,I383620,I801763,I383660,I383677,I383685,I383702,I383733,I801757,I801772,I383750,I383776,I383784,I383829,I801778,I383846,I383949,I713913,I383975,I383983,I713904,I713919,I384000,I713925,I384026,I383917,I384048,I713910,I384074,I384082,I384099,I384125,I383941,I384147,I383923,I713907,I384187,I384204,I384212,I384229,I383926,I384260,I713901,I713916,I384277,I384303,I384311,I383914,I383932,I384356,I713922,I384373,I383935,I383920,I383929,I383938,I384476,I695417,I384502,I384510,I695408,I695423,I384527,I695429,I384553,I384444,I384575,I695414,I384601,I384609,I384626,I384652,I384468,I384674,I384450,I695411,I384714,I384731,I384739,I384756,I384453,I384787,I695405,I695420,I384804,I384830,I384838,I384441,I384459,I384883,I695426,I384900,I384462,I384447,I384456,I384465,I385003,I698885,I385029,I385037,I698876,I698891,I385054,I698897,I385080,I384971,I385102,I698882,I385128,I385136,I385153,I385179,I384995,I385201,I384977,I698879,I385241,I385258,I385266,I385283,I384980,I385314,I698873,I698888,I385331,I385357,I385365,I384968,I384986,I385410,I698894,I385427,I384989,I384974,I384983,I384992,I385530,I663627,I385556,I385564,I663618,I663633,I385581,I663639,I385607,I385498,I385629,I663624,I385655,I385663,I385680,I385706,I385522,I385728,I385504,I663621,I385768,I385785,I385793,I385810,I385507,I385841,I663615,I663630,I385858,I385884,I385892,I385495,I385513,I385937,I663636,I385954,I385516,I385501,I385510,I385519,I386057,I386083,I386091,I386108,I386134,I386025,I386156,I386182,I386190,I386207,I386233,I386049,I386255,I386031,I386295,I386312,I386320,I386337,I386034,I386368,I386385,I386411,I386419,I386022,I386040,I386464,I386481,I386043,I386028,I386037,I386046,I386584,I892217,I386610,I386618,I892220,I892214,I386635,I892226,I386661,I386552,I386683,I892229,I386709,I386717,I386734,I386760,I386576,I386782,I386558,I892232,I386822,I386839,I386847,I386864,I386561,I386895,I892223,I386912,I386938,I386946,I386549,I386567,I386991,I892235,I387008,I386570,I386555,I386564,I386573,I387111,I387137,I387145,I387162,I387188,I387079,I387210,I387236,I387244,I387261,I387287,I387103,I387309,I387085,I387349,I387366,I387374,I387391,I387088,I387422,I387439,I387465,I387473,I387076,I387094,I387518,I387535,I387097,I387082,I387091,I387100,I387638,I759575,I387664,I387672,I759566,I759581,I387689,I759587,I387715,I387737,I759572,I387763,I387771,I387788,I387814,I387836,I759569,I387876,I387893,I387901,I387918,I387949,I759563,I759578,I387966,I387992,I388000,I388045,I759584,I388062,I388165,I782117,I388191,I388199,I782108,I782123,I388216,I782129,I388242,I388133,I388264,I782114,I388290,I388298,I388315,I388341,I388157,I388363,I388139,I782111,I388403,I388420,I388428,I388445,I388142,I388476,I782105,I782120,I388493,I388519,I388527,I388130,I388148,I388572,I782126,I388589,I388151,I388136,I388145,I388154,I388692,I1267099,I388718,I388726,I1267081,I1267105,I388743,I1267096,I388769,I388791,I1267102,I388817,I388825,I1267090,I388842,I388868,I388890,I388930,I388947,I388955,I388972,I389003,I1267087,I1267084,I389020,I1267093,I389046,I389054,I389099,I389116,I389219,I852692,I389245,I389253,I852695,I852689,I389270,I852701,I389296,I389187,I389318,I852704,I389344,I389352,I389369,I389395,I389211,I389417,I389193,I852707,I389457,I389474,I389482,I389499,I389196,I389530,I852698,I389547,I389573,I389581,I389184,I389202,I389626,I852710,I389643,I389205,I389190,I389199,I389208,I389746,I389772,I389780,I389797,I389823,I389845,I389871,I389879,I389896,I389922,I389944,I389984,I390001,I390009,I390026,I390057,I390074,I390100,I390108,I390153,I390170,I390273,I767667,I390299,I390307,I767658,I767673,I390324,I767679,I390350,I390241,I390372,I767664,I390398,I390406,I390423,I390449,I390265,I390471,I390247,I767661,I390511,I390528,I390536,I390553,I390250,I390584,I767655,I767670,I390601,I390627,I390635,I390238,I390256,I390680,I767676,I390697,I390259,I390244,I390253,I390262,I390800,I390826,I390834,I390851,I390877,I390768,I390899,I390925,I390933,I390950,I390976,I390792,I390998,I390774,I391038,I391055,I391063,I391080,I390777,I391111,I391128,I391154,I391162,I390765,I390783,I391207,I391224,I390786,I390771,I390780,I390789,I391327,I391353,I391361,I391378,I391404,I391295,I391426,I391452,I391460,I391477,I391503,I391319,I391525,I391301,I391565,I391582,I391590,I391607,I391304,I391638,I391655,I391681,I391689,I391292,I391310,I391734,I391751,I391313,I391298,I391307,I391316,I391854,I1062370,I391880,I391888,I1062367,I391905,I1062379,I391931,I391822,I391953,I391979,I391987,I1062385,I392004,I392030,I391846,I392052,I391828,I1062373,I392092,I392109,I392117,I392134,I391831,I392165,I1062382,I1062388,I392182,I392208,I392216,I391819,I391837,I392261,I1062376,I392278,I391840,I391825,I391834,I391843,I392381,I793099,I392407,I392415,I793090,I793105,I392432,I793111,I392458,I392349,I392480,I793096,I392506,I392514,I392531,I392557,I392373,I392579,I392355,I793093,I392619,I392636,I392644,I392661,I392358,I392692,I793087,I793102,I392709,I392735,I392743,I392346,I392364,I392788,I793108,I392805,I392367,I392352,I392361,I392370,I392908,I1186365,I392934,I392942,I1186380,I392959,I1186383,I392985,I392876,I393007,I1186389,I393033,I393041,I1186371,I393058,I393084,I392900,I393106,I392882,I1186368,I393146,I393163,I393171,I393188,I392885,I393219,I1186374,I393236,I1186386,I393262,I393270,I392873,I392891,I393315,I1186377,I393332,I392894,I392879,I392888,I392897,I393435,I511086,I393461,I393469,I511098,I511077,I393486,I511101,I393512,I393403,I393534,I511092,I393560,I393568,I511074,I393585,I393611,I393427,I393633,I393409,I511089,I393673,I393690,I393698,I393715,I393412,I393746,I511080,I393763,I511083,I393789,I393797,I393400,I393418,I393842,I511095,I393859,I393421,I393406,I393415,I393424,I393962,I853219,I393988,I393996,I853222,I853216,I394013,I853228,I394039,I393930,I394061,I853231,I394087,I394095,I394112,I394138,I393954,I394160,I393936,I853234,I394200,I394217,I394225,I394242,I393939,I394273,I853225,I394290,I394316,I394324,I393927,I393945,I394369,I853237,I394386,I393948,I393933,I393942,I393951,I394489,I1248059,I394515,I394523,I1248041,I1248065,I394540,I1248056,I394566,I394457,I394588,I1248062,I394614,I394622,I1248050,I394639,I394665,I394481,I394687,I394463,I394727,I394744,I394752,I394769,I394466,I394800,I1248047,I1248044,I394817,I1248053,I394843,I394851,I394454,I394472,I394896,I394913,I394475,I394460,I394469,I394478,I395016,I1136079,I395042,I395050,I1136094,I395067,I1136097,I395093,I395115,I1136103,I395141,I395149,I1136085,I395166,I395192,I395214,I1136082,I395254,I395271,I395279,I395296,I395327,I1136088,I395344,I1136100,I395370,I395378,I395423,I1136091,I395440,I395543,I395569,I395577,I395594,I395620,I395642,I395668,I395676,I395693,I395719,I395741,I395781,I395798,I395806,I395823,I395854,I395871,I395897,I395905,I395950,I395967,I396070,I1093885,I396096,I396104,I1093900,I396121,I1093903,I396147,I396038,I396169,I1093909,I396195,I396203,I1093891,I396220,I396246,I396062,I396268,I396044,I1093888,I396308,I396325,I396333,I396350,I396047,I396381,I1093894,I396398,I1093906,I396424,I396432,I396035,I396053,I396477,I1093897,I396494,I396056,I396041,I396050,I396059,I396597,I895906,I396623,I396631,I895909,I895903,I396648,I895915,I396674,I396565,I396696,I895918,I396722,I396730,I396747,I396773,I396589,I396795,I396571,I895921,I396835,I396852,I396860,I396877,I396574,I396908,I895912,I396925,I396951,I396959,I396562,I396580,I397004,I895924,I397021,I396583,I396568,I396577,I396586,I397124,I814221,I397150,I397158,I814224,I814218,I397175,I814230,I397201,I397092,I397223,I814233,I397249,I397257,I397274,I397300,I397116,I397322,I397098,I814236,I397362,I397379,I397387,I397404,I397101,I397435,I814227,I397452,I397478,I397486,I397089,I397107,I397531,I814239,I397548,I397110,I397095,I397104,I397113,I397651,I1023406,I397677,I397685,I1023403,I1023421,I397702,I1023412,I397728,I397619,I397750,I1023427,I397776,I397784,I1023409,I397801,I397827,I397643,I397849,I397625,I1023415,I397889,I397906,I397914,I397931,I397628,I397962,I1023430,I397979,I1023418,I398005,I398013,I397616,I397634,I398058,I1023424,I398075,I397637,I397622,I397631,I397640,I398178,I398204,I398212,I398229,I398255,I398146,I398277,I398303,I398311,I398328,I398354,I398170,I398376,I398152,I398416,I398433,I398441,I398458,I398155,I398489,I398506,I398532,I398540,I398143,I398161,I398585,I398602,I398164,I398149,I398158,I398167,I398705,I1190989,I398731,I398739,I1191004,I398756,I1191007,I398782,I398673,I398804,I1191013,I398830,I398838,I1190995,I398855,I398881,I398697,I398903,I398679,I1190992,I398943,I398960,I398968,I398985,I398682,I399016,I1190998,I399033,I1191010,I399059,I399067,I398670,I398688,I399112,I1191001,I399129,I398691,I398676,I398685,I398694,I399232,I399258,I399266,I399283,I399309,I399331,I399357,I399365,I399382,I399408,I399430,I399470,I399487,I399495,I399512,I399543,I399560,I399586,I399594,I399639,I399656,I399759,I1015008,I399785,I399793,I1015005,I1015023,I399810,I1015014,I399836,I399727,I399858,I1015029,I399884,I399892,I1015011,I399909,I399935,I399751,I399957,I399733,I1015017,I399997,I400014,I400022,I400039,I399736,I400070,I1015032,I400087,I1015020,I400113,I400121,I399724,I399742,I400166,I1015026,I400183,I399745,I399730,I399739,I399748,I400286,I936196,I400312,I400320,I936193,I936211,I400337,I936202,I400363,I400254,I400385,I936217,I400411,I400419,I936199,I400436,I400462,I400278,I400484,I400260,I936205,I400524,I400541,I400549,I400566,I400263,I400597,I936220,I400614,I936208,I400640,I400648,I400251,I400269,I400693,I936214,I400710,I400272,I400257,I400266,I400275,I400813,I1002734,I400839,I400847,I1002731,I1002749,I400864,I1002740,I400890,I400781,I400912,I1002755,I400938,I400946,I1002737,I400963,I400989,I400805,I401011,I400787,I1002743,I401051,I401068,I401076,I401093,I400790,I401124,I1002758,I401141,I1002746,I401167,I401175,I400778,I400796,I401220,I1002752,I401237,I400799,I400784,I400793,I400802,I401340,I401366,I401374,I401391,I401417,I401308,I401439,I401465,I401473,I401490,I401516,I401332,I401538,I401314,I401578,I401595,I401603,I401620,I401317,I401651,I401668,I401694,I401702,I401305,I401323,I401747,I401764,I401326,I401311,I401320,I401329,I401867,I998212,I401893,I401901,I998209,I998227,I401918,I998218,I401944,I401835,I401966,I998233,I401992,I402000,I998215,I402017,I402043,I401859,I402065,I401841,I998221,I402105,I402122,I402130,I402147,I401844,I402178,I998236,I402195,I998224,I402221,I402229,I401832,I401850,I402274,I998230,I402291,I401853,I401838,I401847,I401856,I402394,I402420,I402428,I402445,I402471,I402362,I402493,I402519,I402527,I402544,I402570,I402386,I402592,I402368,I402632,I402649,I402657,I402674,I402371,I402705,I402722,I402748,I402756,I402359,I402377,I402801,I402818,I402380,I402365,I402374,I402383,I402921,I402947,I402955,I402972,I402998,I402889,I403020,I403046,I403054,I403071,I403097,I402913,I403119,I402895,I403159,I403176,I403184,I403201,I402898,I403232,I403249,I403275,I403283,I402886,I402904,I403328,I403345,I402907,I402892,I402901,I402910,I403448,I711023,I403474,I403482,I711014,I711029,I403499,I711035,I403525,I403416,I403547,I711020,I403573,I403581,I403598,I403624,I403440,I403646,I403422,I711017,I403686,I403703,I403711,I403728,I403425,I403759,I711011,I711026,I403776,I403802,I403810,I403413,I403431,I403855,I711032,I403872,I403434,I403419,I403428,I403437,I403975,I927152,I404001,I404009,I927149,I927167,I404026,I927158,I404052,I403943,I404074,I927173,I404100,I404108,I927155,I404125,I404151,I403967,I404173,I403949,I927161,I404213,I404230,I404238,I404255,I403952,I404286,I927176,I404303,I927164,I404329,I404337,I403940,I403958,I404382,I927170,I404399,I403961,I403946,I403955,I403964,I404502,I695995,I404528,I404536,I695986,I696001,I404553,I696007,I404579,I404470,I404601,I695992,I404627,I404635,I404652,I404678,I404494,I404700,I404476,I695989,I404740,I404757,I404765,I404782,I404479,I404813,I695983,I695998,I404830,I404856,I404864,I404467,I404485,I404909,I696004,I404926,I404488,I404473,I404482,I404491,I405029,I1357134,I405055,I405063,I1357113,I405080,I1357140,I405106,I404997,I405128,I1357128,I405154,I405162,I1357131,I405179,I405205,I405021,I405227,I405003,I1357122,I405267,I405284,I405292,I405309,I405006,I405340,I1357119,I1357116,I405357,I1357137,I405383,I405391,I404994,I405012,I405436,I1357125,I405453,I405015,I405000,I405009,I405018,I405556,I1028574,I405582,I405590,I1028571,I1028589,I405607,I1028580,I405633,I405524,I405655,I1028595,I405681,I405689,I1028577,I405706,I405732,I405548,I405754,I405530,I1028583,I405794,I405811,I405819,I405836,I405533,I405867,I1028598,I405884,I1028586,I405910,I405918,I405521,I405539,I405963,I1028592,I405980,I405542,I405527,I405536,I405545,I406083,I824234,I406109,I406117,I824237,I824231,I406134,I824243,I406160,I406051,I406182,I824246,I406208,I406216,I406233,I406259,I406075,I406281,I406057,I824249,I406321,I406338,I406346,I406363,I406060,I406394,I824240,I406411,I406437,I406445,I406048,I406066,I406490,I824252,I406507,I406069,I406054,I406063,I406072,I406610,I406636,I406644,I406661,I406687,I406578,I406709,I406735,I406743,I406760,I406786,I406602,I406808,I406584,I406848,I406865,I406873,I406890,I406587,I406921,I406938,I406964,I406972,I406575,I406593,I407017,I407034,I406596,I406581,I406590,I406599,I407137,I486606,I407163,I407171,I486618,I486597,I407188,I486621,I407214,I407236,I486612,I407262,I407270,I486594,I407287,I407313,I407335,I486609,I407375,I407392,I407400,I407417,I407448,I486600,I407465,I486603,I407491,I407499,I407544,I486615,I407561,I407664,I407690,I407698,I407715,I407741,I407632,I407763,I407789,I407797,I407814,I407840,I407656,I407862,I407638,I407902,I407919,I407927,I407944,I407641,I407975,I407992,I408018,I408026,I407629,I407647,I408071,I408088,I407650,I407635,I407644,I407653,I408191,I625482,I408217,I408225,I625467,I625470,I408242,I625485,I408268,I408159,I408290,I625479,I408316,I408324,I408341,I408367,I408183,I408389,I408165,I625476,I408429,I408446,I408454,I408471,I408168,I408502,I625491,I408519,I625488,I408545,I408553,I408156,I408174,I408598,I625473,I408615,I408177,I408162,I408171,I408180,I408718,I1032450,I408744,I408752,I1032447,I1032465,I408769,I1032456,I408795,I408686,I408817,I1032471,I408843,I408851,I1032453,I408868,I408894,I408710,I408916,I408692,I1032459,I408956,I408973,I408981,I408998,I408695,I409029,I1032474,I409046,I1032462,I409072,I409080,I408683,I408701,I409125,I1032468,I409142,I408704,I408689,I408698,I408707,I409245,I1017592,I409271,I409279,I1017589,I1017607,I409296,I1017598,I409322,I409213,I409344,I1017613,I409370,I409378,I1017595,I409395,I409421,I409237,I409443,I409219,I1017601,I409483,I409500,I409508,I409525,I409222,I409556,I1017616,I409573,I1017604,I409599,I409607,I409210,I409228,I409652,I1017610,I409669,I409231,I409216,I409225,I409234,I409772,I904338,I409798,I409806,I904341,I904335,I409823,I904347,I409849,I409740,I409871,I904350,I409897,I409905,I409922,I409948,I409764,I409970,I409746,I904353,I410010,I410027,I410035,I410052,I409749,I410083,I904344,I410100,I410126,I410134,I409737,I409755,I410179,I904356,I410196,I409758,I409743,I409752,I409761,I410299,I1212375,I410325,I410333,I1212390,I410350,I1212393,I410376,I410267,I410398,I1212399,I410424,I410432,I1212381,I410449,I410475,I410291,I410497,I410273,I1212378,I410537,I410554,I410562,I410579,I410276,I410610,I1212384,I410627,I1212396,I410653,I410661,I410264,I410282,I410706,I1212387,I410723,I410285,I410270,I410279,I410288,I410826,I697729,I410852,I410860,I697720,I697735,I410877,I697741,I410903,I410794,I410925,I697726,I410951,I410959,I410976,I411002,I410818,I411024,I410800,I697723,I411064,I411081,I411089,I411106,I410803,I411137,I697717,I697732,I411154,I411180,I411188,I410791,I410809,I411233,I697738,I411250,I410812,I410797,I410806,I410815,I411353,I411379,I411387,I411404,I411430,I411452,I411478,I411486,I411503,I411529,I411551,I411591,I411608,I411616,I411633,I411664,I411681,I411707,I411715,I411760,I411777,I411880,I1184053,I411906,I411914,I1184068,I411931,I1184071,I411957,I411979,I1184077,I412005,I412013,I1184059,I412030,I412056,I412078,I1184056,I412118,I412135,I412143,I412160,I412191,I1184062,I412208,I1184074,I412234,I412242,I412287,I1184065,I412304,I412407,I451790,I412433,I412441,I451802,I451781,I412458,I451805,I412484,I412375,I412506,I451796,I412532,I412540,I451778,I412557,I412583,I412399,I412605,I412381,I451793,I412645,I412662,I412670,I412687,I412384,I412718,I451784,I412735,I451787,I412761,I412769,I412372,I412390,I412814,I451799,I412831,I412393,I412378,I412387,I412396,I412934,I1379744,I412960,I412968,I1379723,I412985,I1379750,I413011,I412902,I413033,I1379738,I413059,I413067,I1379741,I413084,I413110,I412926,I413132,I412908,I1379732,I413172,I413189,I413197,I413214,I412911,I413245,I1379729,I1379726,I413262,I1379747,I413288,I413296,I412899,I412917,I413341,I1379735,I413358,I412920,I412905,I412914,I412923,I413461,I413487,I413495,I413512,I413538,I413429,I413560,I413586,I413594,I413611,I413637,I413453,I413659,I413435,I413699,I413716,I413724,I413741,I413438,I413772,I413789,I413815,I413823,I413426,I413444,I413868,I413885,I413447,I413432,I413441,I413450,I413988,I414014,I414022,I414039,I414065,I413956,I414087,I414113,I414121,I414138,I414164,I413980,I414186,I413962,I414226,I414243,I414251,I414268,I413965,I414299,I414316,I414342,I414350,I413953,I413971,I414395,I414412,I413974,I413959,I413968,I413977,I414515,I800613,I414541,I414549,I800604,I800619,I414566,I800625,I414592,I414614,I800610,I414640,I414648,I414665,I414691,I414713,I800607,I414753,I414770,I414778,I414795,I414826,I800601,I800616,I414843,I414869,I414877,I414922,I800622,I414939,I415042,I1284507,I415068,I415076,I1284489,I1284513,I415093,I1284504,I415119,I415010,I415141,I1284510,I415167,I415175,I1284498,I415192,I415218,I415034,I415240,I415016,I415280,I415297,I415305,I415322,I415019,I415353,I1284495,I1284492,I415370,I1284501,I415396,I415404,I415007,I415025,I415449,I415466,I415028,I415013,I415022,I415031,I415569,I1190411,I415595,I415603,I1190426,I415620,I1190429,I415646,I415537,I415668,I1190435,I415694,I415702,I1190417,I415719,I415745,I415561,I415767,I415543,I1190414,I415807,I415824,I415832,I415849,I415546,I415880,I1190420,I415897,I1190432,I415923,I415931,I415534,I415552,I415976,I1190423,I415993,I415555,I415540,I415549,I415558,I416096,I905392,I416122,I416130,I905395,I905389,I416147,I905401,I416173,I416064,I416195,I905404,I416221,I416229,I416246,I416272,I416088,I416294,I416070,I905407,I416334,I416351,I416359,I416376,I416073,I416407,I905398,I416424,I416450,I416458,I416061,I416079,I416503,I905410,I416520,I416082,I416067,I416076,I416085,I416623,I416649,I416657,I416674,I416700,I416591,I416722,I416748,I416756,I416773,I416799,I416615,I416821,I416597,I416861,I416878,I416886,I416903,I416600,I416934,I416951,I416977,I416985,I416588,I416606,I417030,I417047,I416609,I416594,I416603,I416612,I417150,I1147639,I417176,I417184,I1147654,I417201,I1147657,I417227,I417249,I1147663,I417275,I417283,I1147645,I417300,I417326,I417348,I1147642,I417388,I417405,I417413,I417430,I417461,I1147648,I417478,I1147660,I417504,I417512,I417557,I1147651,I417574,I417677,I586756,I417703,I417711,I586741,I586744,I417728,I586759,I417754,I417645,I417776,I586753,I417802,I417810,I417827,I417853,I417669,I417875,I417651,I586750,I417915,I417932,I417940,I417957,I417654,I417988,I586765,I418005,I586762,I418031,I418039,I417642,I417660,I418084,I586747,I418101,I417663,I417648,I417657,I417666,I418204,I1357729,I418230,I418238,I1357708,I418255,I1357735,I418281,I418303,I1357723,I418329,I418337,I1357726,I418354,I418380,I418402,I1357717,I418442,I418459,I418467,I418484,I418515,I1357714,I1357711,I418532,I1357732,I418558,I418566,I418611,I1357720,I418628,I418731,I842152,I418757,I418765,I842155,I842149,I418782,I842161,I418808,I418699,I418830,I842164,I418856,I418864,I418881,I418907,I418723,I418929,I418705,I842167,I418969,I418986,I418994,I419011,I418708,I419042,I842158,I419059,I419085,I419093,I418696,I418714,I419138,I842170,I419155,I418717,I418702,I418711,I418720,I419258,I1348804,I419284,I419292,I1348783,I419309,I1348810,I419335,I419226,I419357,I1348798,I419383,I419391,I1348801,I419408,I419434,I419250,I419456,I419232,I1348792,I419496,I419513,I419521,I419538,I419235,I419569,I1348789,I1348786,I419586,I1348807,I419612,I419620,I419223,I419241,I419665,I1348795,I419682,I419244,I419229,I419238,I419247,I419785,I419811,I419819,I419836,I419862,I419884,I419910,I419918,I419935,I419961,I419983,I420023,I420040,I420048,I420065,I420096,I420113,I420139,I420147,I420192,I420209,I420312,I420338,I420346,I420363,I420389,I420280,I420411,I420437,I420445,I420462,I420488,I420304,I420510,I420286,I420550,I420567,I420575,I420592,I420289,I420623,I420640,I420666,I420674,I420277,I420295,I420719,I420736,I420298,I420283,I420292,I420301,I420839,I672297,I420865,I420873,I672288,I672303,I420890,I672309,I420916,I420807,I420938,I672294,I420964,I420972,I420989,I421015,I420831,I421037,I420813,I672291,I421077,I421094,I421102,I421119,I420816,I421150,I672285,I672300,I421167,I421193,I421201,I420804,I420822,I421246,I672306,I421263,I420825,I420810,I420819,I420828,I421366,I421392,I421400,I421417,I421443,I421334,I421465,I421491,I421499,I421516,I421542,I421358,I421564,I421340,I421604,I421621,I421629,I421646,I421343,I421677,I421694,I421720,I421728,I421331,I421349,I421773,I421790,I421352,I421337,I421346,I421355,I421893,I421919,I421936,I421958,I421975,I421992,I422018,I422026,I422052,I422060,I422077,I422117,I422125,I422170,I422187,I422213,I422235,I422252,I422269,I422300,I422317,I422348,I422437,I921987,I422463,I422480,I422429,I422502,I422519,I922002,I921990,I422536,I921981,I422562,I422570,I921993,I422596,I422604,I921984,I422621,I422408,I921999,I422661,I422669,I422402,I422417,I422714,I922008,I921996,I422731,I922005,I422757,I422405,I422779,I422796,I422813,I422420,I422844,I422861,I422411,I422892,I422414,I422426,I422423,I422981,I728932,I423007,I423024,I422973,I423046,I423063,I728953,I728944,I423080,I423106,I423114,I728938,I423140,I423148,I728935,I423165,I422952,I728929,I423205,I423213,I422946,I422961,I423258,I728941,I423275,I728950,I423301,I422949,I423323,I423340,I423357,I422964,I423388,I423405,I728947,I422955,I423436,I422958,I422970,I422967,I423525,I423551,I423568,I423590,I423607,I423624,I423650,I423658,I423684,I423692,I423709,I423749,I423757,I423802,I423819,I423845,I423867,I423884,I423901,I423932,I423949,I423980,I424069,I424095,I424112,I424061,I424134,I424151,I424168,I424194,I424202,I424228,I424236,I424253,I424040,I424293,I424301,I424034,I424049,I424346,I424363,I424389,I424037,I424411,I424428,I424445,I424052,I424476,I424493,I424043,I424524,I424046,I424058,I424055,I424613,I1149376,I424639,I424656,I424605,I424678,I424695,I1149388,I424712,I1149379,I424738,I424746,I1149397,I424772,I424780,I1149373,I424797,I424584,I1149391,I424837,I424845,I424578,I424593,I424890,I1149385,I1149382,I424907,I1149394,I424933,I424581,I424955,I424972,I424989,I424596,I425020,I425037,I424587,I425068,I424590,I424602,I424599,I425157,I885902,I425183,I425200,I425149,I425222,I425239,I885896,I885893,I425256,I885908,I425282,I425290,I425316,I425324,I885890,I425341,I425128,I425381,I425389,I425122,I425137,I425434,I885905,I885899,I425451,I425477,I425125,I425499,I425516,I425533,I425140,I425564,I425581,I885911,I425131,I425612,I425134,I425146,I425143,I425701,I425727,I425744,I425766,I425783,I425800,I425826,I425834,I425860,I425868,I425885,I425925,I425933,I425978,I425995,I426021,I426043,I426060,I426077,I426108,I426125,I426156,I426245,I1382130,I426271,I426288,I426310,I426327,I1382106,I1382127,I426344,I1382124,I426370,I426378,I1382103,I426404,I426412,I1382115,I426429,I1382118,I426469,I426477,I426522,I1382121,I1382109,I426539,I1382112,I426565,I426587,I426604,I426621,I426652,I426669,I426700,I426789,I820027,I426815,I426832,I426781,I426854,I426871,I820021,I820018,I426888,I820033,I426914,I426922,I426948,I426956,I820015,I426973,I426760,I427013,I427021,I426754,I426769,I427066,I820030,I820024,I427083,I427109,I426757,I427131,I427148,I427165,I426772,I427196,I427213,I820036,I426763,I427244,I426766,I426778,I426775,I427333,I752052,I427359,I427376,I427325,I427398,I427415,I752073,I752064,I427432,I427458,I427466,I752058,I427492,I427500,I752055,I427517,I427304,I752049,I427557,I427565,I427298,I427313,I427610,I752061,I427627,I752070,I427653,I427301,I427675,I427692,I427709,I427316,I427740,I427757,I752067,I427307,I427788,I427310,I427322,I427319,I427877,I1095044,I427903,I427920,I427869,I427942,I427959,I1095056,I427976,I1095047,I428002,I428010,I1095065,I428036,I428044,I1095041,I428061,I427848,I1095059,I428101,I428109,I427842,I427857,I428154,I1095053,I1095050,I428171,I1095062,I428197,I427845,I428219,I428236,I428253,I427860,I428284,I428301,I427851,I428332,I427854,I427866,I427863,I428421,I428447,I428464,I428413,I428486,I428503,I428520,I428546,I428554,I428580,I428588,I428605,I428392,I428645,I428653,I428386,I428401,I428698,I428715,I428741,I428389,I428763,I428780,I428797,I428404,I428828,I428845,I428395,I428876,I428398,I428410,I428407,I428965,I428991,I429008,I428957,I429030,I429047,I429064,I429090,I429098,I429124,I429132,I429149,I428936,I429189,I429197,I428930,I428945,I429242,I429259,I429285,I428933,I429307,I429324,I429341,I428948,I429372,I429389,I428939,I429420,I428942,I428954,I428951,I429509,I818973,I429535,I429552,I429574,I429591,I818967,I818964,I429608,I818979,I429634,I429642,I429668,I429676,I818961,I429693,I429733,I429741,I429786,I818976,I818970,I429803,I429829,I429851,I429868,I429885,I429916,I429933,I818982,I429964,I430053,I430079,I430096,I430118,I430135,I430152,I430178,I430186,I430212,I430220,I430237,I430277,I430285,I430330,I430347,I430373,I430395,I430412,I430429,I430460,I430477,I430508,I430597,I1087051,I430623,I430640,I430662,I430679,I1087069,I430696,I1087063,I430722,I430730,I1087057,I430756,I430764,I1087066,I430781,I1087054,I430821,I430829,I430874,I1087072,I430891,I430917,I430939,I430956,I430973,I431004,I431021,I1087060,I431052,I431141,I431167,I431184,I431206,I431223,I431240,I431266,I431274,I431300,I431308,I431325,I431365,I431373,I431418,I431435,I431461,I431483,I431500,I431517,I431548,I431565,I431596,I431685,I431711,I431728,I431677,I431750,I431767,I431784,I431810,I431818,I431844,I431852,I431869,I431656,I431909,I431917,I431650,I431665,I431962,I431979,I432005,I431653,I432027,I432044,I432061,I431668,I432092,I432109,I431659,I432140,I431662,I431674,I431671,I432229,I1059001,I432255,I432272,I432294,I432311,I1059019,I432328,I1059013,I432354,I432362,I1059007,I432388,I432396,I1059016,I432413,I1059004,I432453,I432461,I432506,I1059022,I432523,I432549,I432571,I432588,I432605,I432636,I432653,I1059010,I432684,I432773,I432799,I432816,I432765,I432838,I432855,I432872,I432898,I432906,I432932,I432940,I432957,I432744,I432997,I433005,I432738,I432753,I433050,I433067,I433093,I432741,I433115,I433132,I433149,I432756,I433180,I433197,I432747,I433228,I432750,I432762,I432759,I433317,I756098,I433343,I433360,I433309,I433382,I433399,I756119,I756110,I433416,I433442,I433450,I756104,I433476,I433484,I756101,I433501,I433288,I756095,I433541,I433549,I433282,I433297,I433594,I756107,I433611,I756116,I433637,I433285,I433659,I433676,I433693,I433300,I433724,I433741,I756113,I433291,I433772,I433294,I433306,I433303,I433861,I1194460,I433887,I433904,I433853,I433926,I433943,I1194472,I433960,I1194463,I433986,I433994,I1194481,I434020,I434028,I1194457,I434045,I433832,I1194475,I434085,I434093,I433826,I433841,I434138,I1194469,I1194466,I434155,I1194478,I434181,I433829,I434203,I434220,I434237,I433844,I434268,I434285,I433835,I434316,I433838,I433850,I433847,I434405,I1069660,I434431,I434448,I434397,I434470,I434487,I1069678,I434504,I1069672,I434530,I434538,I1069666,I434564,I434572,I1069675,I434589,I434376,I1069663,I434629,I434637,I434370,I434385,I434682,I1069681,I434699,I434725,I434373,I434747,I434764,I434781,I434388,I434812,I434829,I1069669,I434379,I434860,I434382,I434394,I434391,I434949,I776328,I434975,I434992,I434941,I435014,I435031,I776349,I776340,I435048,I435074,I435082,I776334,I435108,I435116,I776331,I435133,I434920,I776325,I435173,I435181,I434914,I434929,I435226,I776337,I435243,I776346,I435269,I434917,I435291,I435308,I435325,I434932,I435356,I435373,I776343,I434923,I435404,I434926,I434938,I434935,I435493,I435519,I435536,I435558,I435575,I435592,I435618,I435626,I435652,I435660,I435677,I435717,I435725,I435770,I435787,I435813,I435835,I435852,I435869,I435900,I435917,I435948,I436037,I436063,I436080,I436029,I436102,I436119,I436136,I436162,I436170,I436196,I436204,I436221,I436008,I436261,I436269,I436002,I436017,I436314,I436331,I436357,I436005,I436379,I436396,I436413,I436020,I436444,I436461,I436011,I436492,I436014,I436026,I436023,I436581,I1267628,I436607,I436624,I436573,I436646,I436663,I1267640,I1267643,I436680,I1267646,I436706,I436714,I1267631,I436740,I436748,I1267637,I436765,I436552,I1267625,I436805,I436813,I436546,I436561,I436858,I1267649,I436875,I1267634,I436901,I436549,I436923,I436940,I436957,I436564,I436988,I437005,I436555,I437036,I436558,I436570,I436567,I437125,I437151,I437168,I437117,I437190,I437207,I437224,I437250,I437258,I437284,I437292,I437309,I437096,I437349,I437357,I437090,I437105,I437402,I437419,I437445,I437093,I437467,I437484,I437501,I437108,I437532,I437549,I437099,I437580,I437102,I437114,I437111,I437669,I969791,I437695,I437712,I437734,I437751,I969806,I969794,I437768,I969785,I437794,I437802,I969797,I437828,I437836,I969788,I437853,I969803,I437893,I437901,I437946,I969812,I969800,I437963,I969809,I437989,I438011,I438028,I438045,I438076,I438093,I438124,I438213,I1175964,I438239,I438256,I438205,I438278,I438295,I1175976,I438312,I1175967,I438338,I438346,I1175985,I438372,I438380,I1175961,I438397,I438184,I1175979,I438437,I438445,I438178,I438193,I438490,I1175973,I1175970,I438507,I1175982,I438533,I438181,I438555,I438572,I438589,I438196,I438620,I438637,I438187,I438668,I438190,I438202,I438199,I438757,I564984,I438783,I438800,I438749,I438822,I438839,I564987,I565005,I438856,I564993,I438882,I438890,I438916,I438924,I565002,I438941,I438728,I564996,I438981,I438989,I438722,I438737,I439034,I564999,I564981,I439051,I564990,I439077,I438725,I439099,I439116,I439133,I438740,I439164,I439181,I438731,I439212,I438734,I438746,I438743,I439301,I439327,I439344,I439293,I439366,I439383,I439400,I439426,I439434,I439460,I439468,I439485,I439272,I439525,I439533,I439266,I439281,I439578,I439595,I439621,I439269,I439643,I439660,I439677,I439284,I439708,I439725,I439275,I439756,I439278,I439290,I439287,I439845,I439871,I439888,I439837,I439910,I439927,I439944,I439970,I439978,I440004,I440012,I440029,I439816,I440069,I440077,I439810,I439825,I440122,I440139,I440165,I439813,I440187,I440204,I440221,I439828,I440252,I440269,I439819,I440300,I439822,I439834,I439831,I440389,I440415,I440432,I440381,I440454,I440471,I440488,I440514,I440522,I440548,I440556,I440573,I440360,I440613,I440621,I440354,I440369,I440666,I440683,I440709,I440357,I440731,I440748,I440765,I440372,I440796,I440813,I440363,I440844,I440366,I440378,I440375,I440933,I440959,I440976,I440925,I440998,I441015,I441032,I441058,I441066,I441092,I441100,I441117,I440904,I441157,I441165,I440898,I440913,I441210,I441227,I441253,I440901,I441275,I441292,I441309,I440916,I441340,I441357,I440907,I441388,I440910,I440922,I440919,I441477,I1198506,I441503,I441520,I441469,I441542,I441559,I1198518,I441576,I1198509,I441602,I441610,I1198527,I441636,I441644,I1198503,I441661,I441448,I1198521,I441701,I441709,I441442,I441457,I441754,I1198515,I1198512,I441771,I1198524,I441797,I441445,I441819,I441836,I441853,I441460,I441884,I441901,I441451,I441932,I441454,I441466,I441463,I442021,I442047,I442064,I442013,I442086,I442103,I442120,I442146,I442154,I442180,I442188,I442205,I441992,I442245,I442253,I441986,I442001,I442298,I442315,I442341,I441989,I442363,I442380,I442397,I442004,I442428,I442445,I441995,I442476,I441998,I442010,I442007,I442565,I1152266,I442591,I442608,I442557,I442630,I442647,I1152278,I442664,I1152269,I442690,I442698,I1152287,I442724,I442732,I1152263,I442749,I442536,I1152281,I442789,I442797,I442530,I442545,I442842,I1152275,I1152272,I442859,I1152284,I442885,I442533,I442907,I442924,I442941,I442548,I442972,I442989,I442539,I443020,I442542,I442554,I442551,I443109,I748584,I443135,I443152,I443101,I443174,I443191,I748605,I748596,I443208,I443234,I443242,I748590,I443268,I443276,I748587,I443293,I443080,I748581,I443333,I443341,I443074,I443089,I443386,I748593,I443403,I748602,I443429,I443077,I443451,I443468,I443485,I443092,I443516,I443533,I748599,I443083,I443564,I443086,I443098,I443095,I443653,I933615,I443679,I443696,I443645,I443718,I443735,I933630,I933618,I443752,I933609,I443778,I443786,I933621,I443812,I443820,I933612,I443837,I443624,I933627,I443877,I443885,I443618,I443633,I443930,I933636,I933624,I443947,I933633,I443973,I443621,I443995,I444012,I444029,I443636,I444060,I444077,I443627,I444108,I443630,I443642,I443639,I444197,I1306845,I444223,I444240,I444189,I444262,I444279,I1306842,I1306839,I444296,I1306827,I444322,I444330,I1306851,I444356,I444364,I1306836,I444381,I444168,I1306830,I444421,I444429,I444162,I444177,I444474,I1306833,I444491,I1306848,I444517,I444165,I444539,I444556,I444573,I444180,I444604,I444621,I444171,I444652,I444174,I444186,I444183,I444741,I989171,I444767,I444784,I444733,I444806,I444823,I989186,I989174,I444840,I989165,I444866,I444874,I989177,I444900,I444908,I989168,I444925,I444712,I989183,I444965,I444973,I444706,I444721,I445018,I989192,I989180,I445035,I989189,I445061,I444709,I445083,I445100,I445117,I444724,I445148,I445165,I444715,I445196,I444718,I444730,I444727,I445285,I445311,I445328,I445277,I445350,I445367,I445384,I445410,I445418,I445444,I445452,I445469,I445256,I445509,I445517,I445250,I445265,I445562,I445579,I445605,I445253,I445627,I445644,I445661,I445268,I445692,I445709,I445259,I445740,I445262,I445274,I445271,I445829,I445855,I445872,I445821,I445894,I445911,I445928,I445954,I445962,I445988,I445996,I446013,I445800,I446053,I446061,I445794,I445809,I446106,I446123,I446149,I445797,I446171,I446188,I446205,I445812,I446236,I446253,I445803,I446284,I445806,I445818,I445815,I446373,I1171918,I446399,I446416,I446365,I446438,I446455,I1171930,I446472,I1171921,I446498,I446506,I1171939,I446532,I446540,I1171915,I446557,I446344,I1171933,I446597,I446605,I446338,I446353,I446650,I1171927,I1171924,I446667,I1171936,I446693,I446341,I446715,I446732,I446749,I446356,I446780,I446797,I446347,I446828,I446350,I446362,I446359,I446917,I883267,I446943,I446960,I446982,I446999,I883261,I883258,I447016,I883273,I447042,I447050,I447076,I447084,I883255,I447101,I447141,I447149,I447194,I883270,I883264,I447211,I447237,I447259,I447276,I447293,I447324,I447341,I883276,I447372,I447461,I1055635,I447487,I447504,I447453,I447526,I447543,I1055653,I447560,I1055647,I447586,I447594,I1055641,I447620,I447628,I1055650,I447645,I447432,I1055638,I447685,I447693,I447426,I447441,I447738,I1055656,I447755,I447781,I447429,I447803,I447820,I447837,I447444,I447868,I447885,I1055644,I447435,I447916,I447438,I447450,I447447,I448005,I1200818,I448031,I448048,I447997,I448070,I448087,I1200830,I448104,I1200821,I448130,I448138,I1200839,I448164,I448172,I1200815,I448189,I447976,I1200833,I448229,I448237,I447970,I447985,I448282,I1200827,I1200824,I448299,I1200836,I448325,I447973,I448347,I448364,I448381,I447988,I448412,I448429,I447979,I448460,I447982,I447994,I447991,I448549,I1364280,I448575,I448592,I448541,I448614,I448631,I1364256,I1364277,I448648,I1364274,I448674,I448682,I1364253,I448708,I448716,I1364265,I448733,I448520,I1364268,I448773,I448781,I448514,I448529,I448826,I1364271,I1364259,I448843,I1364262,I448869,I448517,I448891,I448908,I448925,I448532,I448956,I448973,I448523,I449004,I448526,I448538,I448535,I449093,I832675,I449119,I449136,I449158,I449175,I832669,I832666,I449192,I832681,I449218,I449226,I449252,I449260,I832663,I449277,I449317,I449325,I449370,I832678,I832672,I449387,I449413,I449435,I449452,I449469,I449500,I449517,I832684,I449548,I449637,I1385105,I449663,I449680,I449629,I449702,I449719,I1385081,I1385102,I449736,I1385099,I449762,I449770,I1385078,I449796,I449804,I1385090,I449821,I449608,I1385093,I449861,I449869,I449602,I449617,I449914,I1385096,I1385084,I449931,I1385087,I449957,I449605,I449979,I449996,I450013,I449620,I450044,I450061,I449611,I450092,I449614,I449626,I449623,I450181,I689050,I450207,I450224,I450246,I450263,I689071,I689062,I450280,I450306,I450314,I689056,I450340,I450348,I689053,I450365,I689047,I450405,I450413,I450458,I689059,I450475,I689068,I450501,I450523,I450540,I450557,I450588,I450605,I689065,I450636,I450725,I1162092,I450751,I450768,I450790,I450807,I1162104,I450824,I1162095,I450850,I450858,I1162113,I450884,I450892,I1162089,I450909,I1162107,I450949,I450957,I451002,I1162101,I1162098,I451019,I1162110,I451045,I451067,I451084,I451101,I451132,I451149,I451180,I451269,I451295,I451312,I451261,I451334,I451351,I451368,I451394,I451402,I451428,I451436,I451453,I451240,I451493,I451501,I451234,I451249,I451546,I451563,I451589,I451237,I451611,I451628,I451645,I451252,I451676,I451693,I451243,I451724,I451246,I451258,I451255,I451813,I906982,I451839,I451856,I451878,I451895,I906976,I906973,I451912,I906988,I451938,I451946,I451972,I451980,I906970,I451997,I452037,I452045,I452090,I906985,I906979,I452107,I452133,I452155,I452172,I452189,I452220,I452237,I906991,I452268,I452357,I811008,I452383,I452400,I452422,I452439,I811029,I811020,I452456,I452482,I452490,I811014,I452516,I452524,I811011,I452541,I811005,I452581,I452589,I452634,I811017,I452651,I811026,I452677,I452699,I452716,I452733,I452764,I452781,I811023,I452812,I452901,I452927,I452944,I452893,I452966,I452983,I453000,I453026,I453034,I453060,I453068,I453085,I452872,I453125,I453133,I452866,I452881,I453178,I453195,I453221,I452869,I453243,I453260,I453277,I452884,I453308,I453325,I452875,I453356,I452878,I452890,I452887,I453445,I539994,I453471,I453488,I453437,I453510,I453527,I539997,I540015,I453544,I540003,I453570,I453578,I453604,I453612,I540012,I453629,I453416,I540006,I453669,I453677,I453410,I453425,I453722,I540009,I539991,I453739,I540000,I453765,I453413,I453787,I453804,I453821,I453428,I453852,I453869,I453419,I453900,I453422,I453434,I453431,I453989,I810430,I454015,I454032,I453981,I454054,I454071,I810451,I810442,I454088,I454114,I454122,I810436,I454148,I454156,I810433,I454173,I453960,I810427,I454213,I454221,I453954,I453969,I454266,I810439,I454283,I810448,I454309,I453957,I454331,I454348,I454365,I453972,I454396,I454413,I810445,I453963,I454444,I453966,I453978,I453975,I454533,I834256,I454559,I454576,I454525,I454598,I454615,I834250,I834247,I454632,I834262,I454658,I454666,I454692,I454700,I834244,I454717,I454504,I454757,I454765,I454498,I454513,I454810,I834259,I834253,I454827,I454853,I454501,I454875,I454892,I454909,I454516,I454940,I454957,I834265,I454507,I454988,I454510,I454522,I454519,I455077,I455103,I455120,I455142,I455159,I455176,I455202,I455210,I455236,I455244,I455261,I455301,I455309,I455354,I455371,I455397,I455419,I455436,I455453,I455484,I455501,I455532,I455621,I1011135,I455647,I455664,I455613,I455686,I455703,I1011150,I1011138,I455720,I1011129,I455746,I455754,I1011141,I455780,I455788,I1011132,I455805,I455592,I1011147,I455845,I455853,I455586,I455601,I455898,I1011156,I1011144,I455915,I1011153,I455941,I455589,I455963,I455980,I455997,I455604,I456028,I456045,I455595,I456076,I455598,I455610,I455607,I456165,I456191,I456208,I456157,I456230,I456247,I456264,I456290,I456298,I456324,I456332,I456349,I456136,I456389,I456397,I456130,I456145,I456442,I456459,I456485,I456133,I456507,I456524,I456541,I456148,I456572,I456589,I456139,I456620,I456142,I456154,I456151,I456709,I969145,I456735,I456752,I456701,I456774,I456791,I969160,I969148,I456808,I969139,I456834,I456842,I969151,I456868,I456876,I969142,I456893,I456680,I969157,I456933,I456941,I456674,I456689,I456986,I969166,I969154,I457003,I969163,I457029,I456677,I457051,I457068,I457085,I456692,I457116,I457133,I456683,I457164,I456686,I456698,I456695,I457253,I982711,I457279,I457296,I457245,I457318,I457335,I982726,I982714,I457352,I982705,I457378,I457386,I982717,I457412,I457420,I982708,I457437,I457224,I982723,I457477,I457485,I457218,I457233,I457530,I982732,I982720,I457547,I982729,I457573,I457221,I457595,I457612,I457629,I457236,I457660,I457677,I457227,I457708,I457230,I457242,I457239,I457797,I1022117,I457823,I457840,I457862,I457879,I1022132,I1022120,I457896,I1022111,I457922,I457930,I1022123,I457956,I457964,I1022114,I457981,I1022129,I458021,I458029,I458074,I1022138,I1022126,I458091,I1022135,I458117,I458139,I458156,I458173,I458204,I458221,I458252,I458341,I1153422,I458367,I458384,I458333,I458406,I458423,I1153434,I458440,I1153425,I458466,I458474,I1153443,I458500,I458508,I1153419,I458525,I458312,I1153437,I458565,I458573,I458306,I458321,I458618,I1153431,I1153428,I458635,I1153440,I458661,I458309,I458683,I458700,I458717,I458324,I458748,I458765,I458315,I458796,I458318,I458330,I458327,I458885,I458911,I458928,I458877,I458950,I458967,I458984,I459010,I459018,I459044,I459052,I459069,I458856,I459109,I459117,I458850,I458865,I459162,I459179,I459205,I458853,I459227,I459244,I459261,I458868,I459292,I459309,I458859,I459340,I458862,I458874,I458871,I459429,I1397005,I459455,I459472,I459421,I459494,I459511,I1396981,I1397002,I459528,I1396999,I459554,I459562,I1396978,I459588,I459596,I1396990,I459613,I459400,I1396993,I459653,I459661,I459394,I459409,I459706,I1396996,I1396984,I459723,I1396987,I459749,I459397,I459771,I459788,I459805,I459412,I459836,I459853,I459403,I459884,I459406,I459418,I459415,I459973,I845323,I459999,I460016,I459965,I460038,I460055,I845317,I845314,I460072,I845329,I460098,I460106,I460132,I460140,I845311,I460157,I459944,I460197,I460205,I459938,I459953,I460250,I845326,I845320,I460267,I460293,I459941,I460315,I460332,I460349,I459956,I460380,I460397,I845332,I459947,I460428,I459950,I459962,I459959,I460517,I1079197,I460543,I460560,I460509,I460582,I460599,I1079215,I460616,I1079209,I460642,I460650,I1079203,I460676,I460684,I1079212,I460701,I460488,I1079200,I460741,I460749,I460482,I460497,I460794,I1079218,I460811,I460837,I460485,I460859,I460876,I460893,I460500,I460924,I460941,I1079206,I460491,I460972,I460494,I460506,I460503,I461061,I819500,I461087,I461104,I461053,I461126,I461143,I819494,I819491,I461160,I819506,I461186,I461194,I461220,I461228,I819488,I461245,I461032,I461285,I461293,I461026,I461041,I461338,I819503,I819497,I461355,I461381,I461029,I461403,I461420,I461437,I461044,I461468,I461485,I819509,I461035,I461516,I461038,I461050,I461047,I461605,I856390,I461631,I461648,I461670,I461687,I856384,I856381,I461704,I856396,I461730,I461738,I461764,I461772,I856378,I461789,I461829,I461837,I461882,I856393,I856387,I461899,I461925,I461947,I461964,I461981,I462012,I462029,I856399,I462060,I462149,I1128568,I462175,I462192,I462141,I462214,I462231,I1128580,I462248,I1128571,I462274,I462282,I1128589,I462308,I462316,I1128565,I462333,I462120,I1128583,I462373,I462381,I462114,I462129,I462426,I1128577,I1128574,I462443,I1128586,I462469,I462117,I462491,I462508,I462525,I462132,I462556,I462573,I462123,I462604,I462126,I462138,I462135,I462693,I1260556,I462719,I462736,I462685,I462758,I462775,I1260568,I1260571,I462792,I1260574,I462818,I462826,I1260559,I462852,I462860,I1260565,I462877,I462664,I1260553,I462917,I462925,I462658,I462673,I462970,I1260577,I462987,I1260562,I463013,I462661,I463035,I463052,I463069,I462676,I463100,I463117,I462667,I463148,I462670,I462682,I462679,I463237,I1377370,I463263,I463280,I463229,I463302,I463319,I1377346,I1377367,I463336,I1377364,I463362,I463370,I1377343,I463396,I463404,I1377355,I463421,I463208,I1377358,I463461,I463469,I463202,I463217,I463514,I1377361,I1377349,I463531,I1377352,I463557,I463205,I463579,I463596,I463613,I463220,I463644,I463661,I463211,I463692,I463214,I463226,I463223,I463781,I1374990,I463807,I463824,I463773,I463846,I463863,I1374966,I1374987,I463880,I1374984,I463906,I463914,I1374963,I463940,I463948,I1374975,I463965,I463752,I1374978,I464005,I464013,I463746,I463761,I464058,I1374981,I1374969,I464075,I1374972,I464101,I463749,I464123,I464140,I464157,I463764,I464188,I464205,I463755,I464236,I463758,I463770,I463767,I464325,I1307423,I464351,I464368,I464317,I464390,I464407,I1307420,I1307417,I464424,I1307405,I464450,I464458,I1307429,I464484,I464492,I1307414,I464509,I464296,I1307408,I464549,I464557,I464290,I464305,I464602,I1307411,I464619,I1307426,I464645,I464293,I464667,I464684,I464701,I464308,I464732,I464749,I464299,I464780,I464302,I464314,I464311,I464869,I464895,I464912,I464861,I464934,I464951,I464968,I464994,I465002,I465028,I465036,I465053,I464840,I465093,I465101,I464834,I464849,I465146,I465163,I465189,I464837,I465211,I465228,I465245,I464852,I465276,I465293,I464843,I465324,I464846,I464858,I464855,I465413,I1036975,I465439,I465456,I465405,I465478,I465495,I1036990,I1036978,I465512,I1036969,I465538,I465546,I1036981,I465572,I465580,I1036972,I465597,I465384,I1036987,I465637,I465645,I465378,I465393,I465690,I1036996,I1036984,I465707,I1036993,I465733,I465381,I465755,I465772,I465789,I465396,I465820,I465837,I465387,I465868,I465390,I465402,I465399,I465957,I962685,I465983,I466000,I465949,I466022,I466039,I962700,I962688,I466056,I962679,I466082,I466090,I962691,I466116,I466124,I962682,I466141,I465928,I962697,I466181,I466189,I465922,I465937,I466234,I962706,I962694,I466251,I962703,I466277,I465925,I466299,I466316,I466333,I465940,I466364,I466381,I465931,I466412,I465934,I465946,I465943,I466501,I643388,I466527,I466544,I466566,I466583,I643385,I643406,I466600,I643409,I466626,I466634,I643394,I466660,I466668,I643397,I466685,I643400,I466725,I466733,I466778,I643391,I466795,I643403,I466821,I466843,I466860,I466877,I466908,I466925,I466956,I467045,I467071,I467088,I467037,I467110,I467127,I467144,I467170,I467178,I467204,I467212,I467229,I467016,I467269,I467277,I467010,I467025,I467322,I467339,I467365,I467013,I467387,I467404,I467421,I467028,I467452,I467469,I467019,I467500,I467022,I467034,I467031,I467589,I467615,I467632,I467581,I467654,I467671,I467688,I467714,I467722,I467748,I467756,I467773,I467560,I467813,I467821,I467554,I467569,I467866,I467883,I467909,I467557,I467931,I467948,I467965,I467572,I467996,I468013,I467563,I468044,I467566,I467578,I467575,I468133,I1311469,I468159,I468176,I468125,I468198,I468215,I1311466,I1311463,I468232,I1311451,I468258,I468266,I1311475,I468292,I468300,I1311460,I468317,I468104,I1311454,I468357,I468365,I468098,I468113,I468410,I1311457,I468427,I1311472,I468453,I468101,I468475,I468492,I468509,I468116,I468540,I468557,I468107,I468588,I468110,I468122,I468119,I468677,I468703,I468720,I468742,I468759,I468776,I468802,I468810,I468836,I468844,I468861,I468901,I468909,I468954,I468971,I468997,I469019,I469036,I469053,I469084,I469101,I469132,I469221,I917465,I469247,I469264,I469213,I469286,I469303,I917480,I917468,I469320,I917459,I469346,I469354,I917471,I469380,I469388,I917462,I469405,I469192,I917477,I469445,I469453,I469186,I469201,I469498,I917486,I917474,I469515,I917483,I469541,I469189,I469563,I469580,I469597,I469204,I469628,I469645,I469195,I469676,I469198,I469210,I469207,I469765,I608130,I469791,I469808,I469757,I469830,I469847,I608127,I608148,I469864,I608151,I469890,I469898,I608136,I469924,I469932,I608139,I469949,I469736,I608142,I469989,I469997,I469730,I469745,I470042,I608133,I470059,I608145,I470085,I469733,I470107,I470124,I470141,I469748,I470172,I470189,I469739,I470220,I469742,I469754,I469751,I470309,I470335,I470352,I470301,I470374,I470391,I470408,I470434,I470442,I470468,I470476,I470493,I470280,I470533,I470541,I470274,I470289,I470586,I470603,I470629,I470277,I470651,I470668,I470685,I470292,I470716,I470733,I470283,I470764,I470286,I470298,I470295,I470853,I470879,I470896,I470845,I470918,I470935,I470952,I470978,I470986,I471012,I471020,I471037,I470824,I471077,I471085,I470818,I470833,I471130,I471147,I471173,I470821,I471195,I471212,I471229,I470836,I471260,I471277,I470827,I471308,I470830,I470842,I470839,I471397,I1363685,I471423,I471440,I471462,I471479,I1363661,I1363682,I471496,I1363679,I471522,I471530,I1363658,I471556,I471564,I1363670,I471581,I1363673,I471621,I471629,I471674,I1363676,I1363664,I471691,I1363667,I471717,I471739,I471756,I471773,I471804,I471821,I471852,I471941,I1323029,I471967,I471984,I471933,I472006,I472023,I1323026,I1323023,I472040,I1323011,I472066,I472074,I1323035,I472100,I472108,I1323020,I472125,I471912,I1323014,I472165,I472173,I471906,I471921,I472218,I1323017,I472235,I1323032,I472261,I471909,I472283,I472300,I472317,I471924,I472348,I472365,I471915,I472396,I471918,I471930,I471927,I472485,I698298,I472511,I472528,I472477,I472550,I472567,I698319,I698310,I472584,I472610,I472618,I698304,I472644,I472652,I698301,I472669,I472456,I698295,I472709,I472717,I472450,I472465,I472762,I698307,I472779,I698316,I472805,I472453,I472827,I472844,I472861,I472468,I472892,I472909,I698313,I472459,I472940,I472462,I472474,I472471,I473029,I1350000,I473055,I473072,I473021,I473094,I473111,I1349976,I1349997,I473128,I1349994,I473154,I473162,I1349973,I473188,I473196,I1349985,I473213,I473000,I1349988,I473253,I473261,I472994,I473009,I473306,I1349991,I1349979,I473323,I1349982,I473349,I472997,I473371,I473388,I473405,I473012,I473436,I473453,I473003,I473484,I473006,I473018,I473015,I473573,I473599,I473616,I473638,I473655,I473672,I473698,I473706,I473732,I473740,I473757,I473797,I473805,I473850,I473867,I473893,I473915,I473932,I473949,I473980,I473997,I474028,I474117,I474143,I474160,I474109,I474182,I474199,I474216,I474242,I474250,I474276,I474284,I474301,I474088,I474341,I474349,I474082,I474097,I474394,I474411,I474437,I474085,I474459,I474476,I474493,I474100,I474524,I474541,I474091,I474572,I474094,I474106,I474103,I474661,I474687,I474704,I474653,I474726,I474743,I474760,I474786,I474794,I474820,I474828,I474845,I474632,I474885,I474893,I474626,I474641,I474938,I474955,I474981,I474629,I475003,I475020,I475037,I474644,I475068,I475085,I474635,I475116,I474638,I474650,I474647,I475205,I994339,I475231,I475248,I475197,I475270,I475287,I994354,I994342,I475304,I994333,I475330,I475338,I994345,I475364,I475372,I994336,I475389,I475176,I994351,I475429,I475437,I475170,I475185,I475482,I994360,I994348,I475499,I994357,I475525,I475173,I475547,I475564,I475581,I475188,I475612,I475629,I475179,I475660,I475182,I475194,I475191,I475749,I1002091,I475775,I475792,I475814,I475831,I1002106,I1002094,I475848,I1002085,I475874,I475882,I1002097,I475908,I475916,I1002088,I475933,I1002103,I475973,I475981,I476026,I1002112,I1002100,I476043,I1002109,I476069,I476091,I476108,I476125,I476156,I476173,I476204,I476293,I883794,I476319,I476336,I476285,I476358,I476375,I883788,I883785,I476392,I883800,I476418,I476426,I476452,I476460,I883782,I476477,I476264,I476517,I476525,I476258,I476273,I476570,I883797,I883791,I476587,I476613,I476261,I476635,I476652,I476669,I476276,I476700,I476717,I883803,I476267,I476748,I476270,I476282,I476279,I476837,I1262188,I476863,I476880,I476829,I476902,I476919,I1262200,I1262203,I476936,I1262206,I476962,I476970,I1262191,I476996,I477004,I1262197,I477021,I476808,I1262185,I477061,I477069,I476802,I476817,I477114,I1262209,I477131,I1262194,I477157,I476805,I477179,I477196,I477213,I476820,I477244,I477261,I476811,I477292,I476814,I476826,I476823,I477381,I477407,I477424,I477373,I477446,I477463,I477480,I477506,I477514,I477540,I477548,I477565,I477352,I477605,I477613,I477346,I477361,I477658,I477675,I477701,I477349,I477723,I477740,I477757,I477364,I477788,I477805,I477355,I477836,I477358,I477370,I477367,I477925,I862187,I477951,I477968,I477990,I478007,I862181,I862178,I478024,I862193,I478050,I478058,I478084,I478092,I862175,I478109,I478149,I478157,I478202,I862190,I862184,I478219,I478245,I478267,I478284,I478301,I478332,I478349,I862196,I478380,I478469,I1248588,I478495,I478512,I478534,I478551,I1248600,I1248603,I478568,I1248606,I478594,I478602,I1248591,I478628,I478636,I1248597,I478653,I1248585,I478693,I478701,I478746,I1248609,I478763,I1248594,I478789,I478811,I478828,I478845,I478876,I478893,I478924,I479013,I1125100,I479039,I479056,I479005,I479078,I479095,I1125112,I479112,I1125103,I479138,I479146,I1125121,I479172,I479180,I1125097,I479197,I478984,I1125115,I479237,I479245,I478978,I478993,I479290,I1125109,I1125106,I479307,I1125118,I479333,I478981,I479355,I479372,I479389,I478996,I479420,I479437,I478987,I479468,I478990,I479002,I478999,I479557,I720262,I479583,I479600,I479622,I479639,I720283,I720274,I479656,I479682,I479690,I720268,I479716,I479724,I720265,I479741,I720259,I479781,I479789,I479834,I720271,I479851,I720280,I479877,I479899,I479916,I479933,I479964,I479981,I720277,I480012,I480101,I1173652,I480127,I480144,I480093,I480166,I480183,I1173664,I480200,I1173655,I480226,I480234,I1173673,I480260,I480268,I1173649,I480285,I480072,I1173667,I480325,I480333,I480066,I480081,I480378,I1173661,I1173658,I480395,I1173670,I480421,I480069,I480443,I480460,I480477,I480084,I480508,I480525,I480075,I480556,I480078,I480090,I480087,I480645,I562009,I480671,I480688,I480637,I480710,I480727,I562012,I562030,I480744,I562018,I480770,I480778,I480804,I480812,I562027,I480829,I480616,I562021,I480869,I480877,I480610,I480625,I480922,I562024,I562006,I480939,I562015,I480965,I480613,I480987,I481004,I481021,I480628,I481052,I481069,I480619,I481100,I480622,I480634,I480631,I481189,I986587,I481215,I481232,I481181,I481254,I481271,I986602,I986590,I481288,I986581,I481314,I481322,I986593,I481348,I481356,I986584,I481373,I481160,I986599,I481413,I481421,I481154,I481169,I481466,I986608,I986596,I481483,I986605,I481509,I481157,I481531,I481548,I481565,I481172,I481596,I481613,I481163,I481644,I481166,I481178,I481175,I481733,I914881,I481759,I481776,I481725,I481798,I481815,I914896,I914884,I481832,I914875,I481858,I481866,I914887,I481892,I481900,I914878,I481917,I481704,I914893,I481957,I481965,I481698,I481713,I482010,I914902,I914890,I482027,I914899,I482053,I481701,I482075,I482092,I482109,I481716,I482140,I482157,I481707,I482188,I481710,I481722,I481719,I482277,I482303,I482320,I482269,I482342,I482359,I482376,I482402,I482410,I482436,I482444,I482461,I482248,I482501,I482509,I482242,I482257,I482554,I482571,I482597,I482245,I482619,I482636,I482653,I482260,I482684,I482701,I482251,I482732,I482254,I482266,I482263,I482821,I1236076,I482847,I482864,I482886,I482903,I1236088,I482920,I1236079,I482946,I482954,I1236097,I482980,I482988,I1236073,I483005,I1236091,I483045,I483053,I483098,I1236085,I1236082,I483115,I1236094,I483141,I483163,I483180,I483197,I483228,I483245,I483276,I483365,I797136,I483391,I483408,I483357,I483430,I483447,I797157,I797148,I483464,I483490,I483498,I797142,I483524,I483532,I797139,I483549,I483336,I797133,I483589,I483597,I483330,I483345,I483642,I797145,I483659,I797154,I483685,I483333,I483707,I483724,I483741,I483348,I483772,I483789,I797151,I483339,I483820,I483342,I483354,I483351,I483909,I1306267,I483935,I483952,I483974,I483991,I1306264,I1306261,I484008,I1306249,I484034,I484042,I1306273,I484068,I484076,I1306258,I484093,I1306252,I484133,I484141,I484186,I1306255,I484203,I1306270,I484229,I484251,I484268,I484285,I484316,I484333,I484364,I484453,I656682,I484479,I484496,I484445,I484518,I484535,I656679,I656700,I484552,I656703,I484578,I484586,I656688,I484612,I484620,I656691,I484637,I484424,I656694,I484677,I484685,I484418,I484433,I484730,I656685,I484747,I656697,I484773,I484421,I484795,I484812,I484829,I484436,I484860,I484877,I484427,I484908,I484430,I484442,I484439,I484997,I653792,I485023,I485040,I485062,I485079,I653789,I653810,I485096,I653813,I485122,I485130,I653798,I485156,I485164,I653801,I485181,I653804,I485221,I485229,I485274,I653795,I485291,I653807,I485317,I485339,I485356,I485373,I485404,I485421,I485452,I485541,I764768,I485567,I485584,I485606,I485623,I764789,I764780,I485640,I485666,I485674,I764774,I485700,I485708,I764771,I485725,I764765,I485765,I485773,I485818,I764777,I485835,I764786,I485861,I485883,I485900,I485917,I485948,I485965,I764783,I485996,I486085,I746850,I486111,I486128,I486077,I486150,I486167,I746871,I746862,I486184,I486210,I486218,I746856,I486244,I486252,I746853,I486269,I486056,I746847,I486309,I486317,I486050,I486065,I486362,I746859,I486379,I746868,I486405,I486053,I486427,I486444,I486461,I486068,I486492,I486509,I746865,I486059,I486540,I486062,I486074,I486071,I486629,I486655,I486672,I486694,I486711,I486728,I486754,I486762,I486788,I486796,I486813,I486853,I486861,I486906,I486923,I486949,I486971,I486988,I487005,I487036,I487053,I487084,I487173,I487199,I487216,I487165,I487238,I487255,I487272,I487298,I487306,I487332,I487340,I487357,I487144,I487397,I487405,I487138,I487153,I487450,I487467,I487493,I487141,I487515,I487532,I487549,I487156,I487580,I487597,I487147,I487628,I487150,I487162,I487159,I487717,I487743,I487760,I487709,I487782,I487799,I487816,I487842,I487850,I487876,I487884,I487901,I487688,I487941,I487949,I487682,I487697,I487994,I488011,I488037,I487685,I488059,I488076,I488093,I487700,I488124,I488141,I487691,I488172,I487694,I487706,I487703,I488261,I547134,I488287,I488304,I488253,I488326,I488343,I547137,I547155,I488360,I547143,I488386,I488394,I488420,I488428,I547152,I488445,I488232,I547146,I488485,I488493,I488226,I488241,I488538,I547149,I547131,I488555,I547140,I488581,I488229,I488603,I488620,I488637,I488244,I488668,I488685,I488235,I488716,I488238,I488250,I488247,I488805,I889064,I488831,I488848,I488870,I488887,I889058,I889055,I488904,I889070,I488930,I488938,I488964,I488972,I889052,I488989,I489029,I489037,I489082,I889067,I889061,I489099,I489125,I489147,I489164,I489181,I489212,I489229,I889073,I489260,I489349,I813176,I489375,I489392,I489341,I489414,I489431,I813170,I813167,I489448,I813182,I489474,I489482,I489508,I489516,I813164,I489533,I489320,I489573,I489581,I489314,I489329,I489626,I813179,I813173,I489643,I489669,I489317,I489691,I489708,I489725,I489332,I489756,I489773,I813185,I489323,I489804,I489326,I489338,I489335,I489893,I684426,I489919,I489936,I489885,I489958,I489975,I684447,I684438,I489992,I490018,I490026,I684432,I490052,I490060,I684429,I490077,I489864,I684423,I490117,I490125,I489858,I489873,I490170,I684435,I490187,I684444,I490213,I489861,I490235,I490252,I490269,I489876,I490300,I490317,I684441,I489867,I490348,I489870,I489882,I489879,I490437,I1091576,I490463,I490480,I490502,I490519,I1091588,I490536,I1091579,I490562,I490570,I1091597,I490596,I490604,I1091573,I490621,I1091591,I490661,I490669,I490714,I1091585,I1091582,I490731,I1091594,I490757,I490779,I490796,I490813,I490844,I490861,I490892,I490981,I491007,I491024,I491046,I491063,I491080,I491106,I491114,I491140,I491148,I491165,I491205,I491213,I491258,I491275,I491301,I491323,I491340,I491357,I491388,I491405,I491436,I491525,I1298175,I491551,I491568,I491517,I491590,I491607,I1298172,I1298169,I491624,I1298157,I491650,I491658,I1298181,I491684,I491692,I1298166,I491709,I491496,I1298160,I491749,I491757,I491490,I491505,I491802,I1298163,I491819,I1298178,I491845,I491493,I491867,I491884,I491901,I491508,I491932,I491949,I491499,I491980,I491502,I491514,I491511,I492069,I1352975,I492095,I492112,I492061,I492134,I492151,I1352951,I1352972,I492168,I1352969,I492194,I492202,I1352948,I492228,I492236,I1352960,I492253,I492040,I1352963,I492293,I492301,I492034,I492049,I492346,I1352966,I1352954,I492363,I1352957,I492389,I492037,I492411,I492428,I492445,I492052,I492476,I492493,I492043,I492524,I492046,I492058,I492055,I492613,I1237810,I492639,I492656,I492678,I492695,I1237822,I492712,I1237813,I492738,I492746,I1237831,I492772,I492780,I1237807,I492797,I1237825,I492837,I492845,I492890,I1237819,I1237816,I492907,I1237828,I492933,I492955,I492972,I492989,I493020,I493037,I493068,I493157,I493183,I493200,I493222,I493239,I493256,I493282,I493290,I493316,I493324,I493341,I493381,I493389,I493434,I493451,I493477,I493499,I493516,I493533,I493564,I493581,I493612,I493701,I704656,I493727,I493744,I493693,I493766,I493783,I704677,I704668,I493800,I493826,I493834,I704662,I493860,I493868,I704659,I493885,I493672,I704653,I493925,I493933,I493666,I493681,I493978,I704665,I493995,I704674,I494021,I493669,I494043,I494060,I494077,I493684,I494108,I494125,I704671,I493675,I494156,I493678,I493690,I493687,I494245,I652636,I494271,I494288,I494237,I494310,I494327,I652633,I652654,I494344,I652657,I494370,I494378,I652642,I494404,I494412,I652645,I494429,I494216,I652648,I494469,I494477,I494210,I494225,I494522,I652639,I494539,I652651,I494565,I494213,I494587,I494604,I494621,I494228,I494652,I494669,I494219,I494700,I494222,I494234,I494231,I494789,I1025347,I494815,I494832,I494781,I494854,I494871,I1025362,I1025350,I494888,I1025341,I494914,I494922,I1025353,I494948,I494956,I1025344,I494973,I494760,I1025359,I495013,I495021,I494754,I494769,I495066,I1025368,I1025356,I495083,I1025365,I495109,I494757,I495131,I495148,I495165,I494772,I495196,I495213,I494763,I495244,I494766,I494778,I494775,I495333,I495359,I495376,I495398,I495415,I495432,I495458,I495466,I495492,I495500,I495517,I495557,I495565,I495610,I495627,I495653,I495675,I495692,I495709,I495740,I495757,I495788,I495877,I495903,I495920,I495942,I495959,I495976,I496002,I496010,I496036,I496044,I496061,I496101,I496109,I496154,I496171,I496197,I496219,I496236,I496253,I496284,I496301,I496332,I496421,I886956,I496447,I496464,I496413,I496486,I496503,I886950,I886947,I496520,I886962,I496546,I496554,I496580,I496588,I886944,I496605,I496392,I496645,I496653,I496386,I496401,I496698,I886959,I886953,I496715,I496741,I496389,I496763,I496780,I496797,I496404,I496828,I496845,I886965,I496395,I496876,I496398,I496410,I496407,I496965,I1078075,I496991,I497008,I496957,I497030,I497047,I1078093,I497064,I1078087,I497090,I497098,I1078081,I497124,I497132,I1078090,I497149,I496936,I1078078,I497189,I497197,I496930,I496945,I497242,I1078096,I497259,I497285,I496933,I497307,I497324,I497341,I496948,I497372,I497389,I1078084,I496939,I497420,I496942,I496954,I496951,I497509,I1333935,I497535,I497552,I497574,I497591,I1333911,I1333932,I497608,I1333929,I497634,I497642,I1333908,I497668,I497676,I1333920,I497693,I1333923,I497733,I497741,I497786,I1333926,I1333914,I497803,I1333917,I497829,I497851,I497868,I497885,I497916,I497933,I497964,I498053,I498079,I498096,I498118,I498135,I498152,I498178,I498186,I498212,I498220,I498237,I498277,I498285,I498330,I498347,I498373,I498395,I498412,I498429,I498460,I498477,I498508,I498597,I498623,I498640,I498589,I498662,I498679,I498696,I498722,I498730,I498756,I498764,I498781,I498568,I498821,I498829,I498562,I498577,I498874,I498891,I498917,I498565,I498939,I498956,I498973,I498580,I499004,I499021,I498571,I499052,I498574,I498586,I498583,I499141,I926509,I499167,I499184,I499133,I499206,I499223,I926524,I926512,I499240,I926503,I499266,I499274,I926515,I499300,I499308,I926506,I499325,I499112,I926521,I499365,I499373,I499106,I499121,I499418,I926530,I926518,I499435,I926527,I499461,I499109,I499483,I499500,I499517,I499124,I499548,I499565,I499115,I499596,I499118,I499130,I499127,I499685,I550109,I499711,I499728,I499677,I499750,I499767,I550112,I550130,I499784,I550118,I499810,I499818,I499844,I499852,I550127,I499869,I499656,I550121,I499909,I499917,I499650,I499665,I499962,I550124,I550106,I499979,I550115,I500005,I499653,I500027,I500044,I500061,I499668,I500092,I500109,I499659,I500140,I499662,I499674,I499671,I500229,I500255,I500272,I500221,I500294,I500311,I500328,I500354,I500362,I500388,I500396,I500413,I500200,I500453,I500461,I500194,I500209,I500506,I500523,I500549,I500197,I500571,I500588,I500605,I500212,I500636,I500653,I500203,I500684,I500206,I500218,I500215,I500773,I500799,I500816,I500765,I500838,I500855,I500872,I500898,I500906,I500932,I500940,I500957,I500744,I500997,I501005,I500738,I500753,I501050,I501067,I501093,I500741,I501115,I501132,I501149,I500756,I501180,I501197,I500747,I501228,I500750,I500762,I500759,I501317,I1158624,I501343,I501360,I501309,I501382,I501399,I1158636,I501416,I1158627,I501442,I501450,I1158645,I501476,I501484,I1158621,I501501,I501288,I1158639,I501541,I501549,I501282,I501297,I501594,I1158633,I1158630,I501611,I1158642,I501637,I501285,I501659,I501676,I501693,I501300,I501724,I501741,I501291,I501772,I501294,I501306,I501303,I501861,I814757,I501887,I501904,I501853,I501926,I501943,I814751,I814748,I501960,I814763,I501986,I501994,I502020,I502028,I814745,I502045,I501832,I502085,I502093,I501826,I501841,I502138,I814760,I814754,I502155,I502181,I501829,I502203,I502220,I502237,I501844,I502268,I502285,I814766,I501835,I502316,I501838,I501850,I501847,I502405,I1289505,I502431,I502448,I502397,I502470,I502487,I1289502,I1289499,I502504,I1289487,I502530,I502538,I1289511,I502564,I502572,I1289496,I502589,I502376,I1289490,I502629,I502637,I502370,I502385,I502682,I1289493,I502699,I1289508,I502725,I502373,I502747,I502764,I502781,I502388,I502812,I502829,I502379,I502860,I502382,I502394,I502391,I502949,I873781,I502975,I502992,I503014,I503031,I873775,I873772,I503048,I873787,I503074,I503082,I503108,I503116,I873769,I503133,I503173,I503181,I503226,I873784,I873778,I503243,I503269,I503291,I503308,I503325,I503356,I503373,I873790,I503404,I503493,I897496,I503519,I503536,I503558,I503575,I897490,I897487,I503592,I897502,I503618,I503626,I503652,I503660,I897484,I503677,I503717,I503725,I503770,I897499,I897493,I503787,I503813,I503835,I503852,I503869,I503900,I503917,I897505,I503948,I504037,I1253484,I504063,I504080,I504029,I504102,I504119,I1253496,I1253499,I504136,I1253502,I504162,I504170,I1253487,I504196,I504204,I1253493,I504221,I504008,I1253481,I504261,I504269,I504002,I504017,I504314,I1253505,I504331,I1253490,I504357,I504005,I504379,I504396,I504413,I504020,I504444,I504461,I504011,I504492,I504014,I504026,I504023,I504581,I1086490,I504607,I504624,I504573,I504646,I504663,I1086508,I504680,I1086502,I504706,I504714,I1086496,I504740,I504748,I1086505,I504765,I504552,I1086493,I504805,I504813,I504546,I504561,I504858,I1086511,I504875,I504901,I504549,I504923,I504940,I504957,I504564,I504988,I505005,I1086499,I504555,I505036,I504558,I504570,I504567,I505125,I570934,I505151,I505168,I505117,I505190,I505207,I570937,I570955,I505224,I570943,I505250,I505258,I505284,I505292,I570952,I505309,I505096,I570946,I505349,I505357,I505090,I505105,I505402,I570949,I570931,I505419,I570940,I505445,I505093,I505467,I505484,I505501,I505108,I505532,I505549,I505099,I505580,I505102,I505114,I505111,I505669,I505695,I505712,I505734,I505751,I505768,I505794,I505802,I505828,I505836,I505853,I505893,I505901,I505946,I505963,I505989,I506011,I506028,I506045,I506076,I506093,I506124,I506213,I506239,I506256,I506205,I506278,I506295,I506312,I506338,I506346,I506372,I506380,I506397,I506184,I506437,I506445,I506178,I506193,I506490,I506507,I506533,I506181,I506555,I506572,I506589,I506196,I506620,I506637,I506187,I506668,I506190,I506202,I506199,I506757,I506783,I506800,I506749,I506822,I506839,I506856,I506882,I506890,I506916,I506924,I506941,I506728,I506981,I506989,I506722,I506737,I507034,I507051,I507077,I506725,I507099,I507116,I507133,I506740,I507164,I507181,I506731,I507212,I506734,I506746,I506743,I507301,I507327,I507344,I507366,I507383,I507400,I507426,I507434,I507460,I507468,I507485,I507525,I507533,I507578,I507595,I507621,I507643,I507660,I507677,I507708,I507725,I507756,I507845,I507871,I507888,I507837,I507910,I507927,I507944,I507970,I507978,I508004,I508012,I508029,I507816,I508069,I508077,I507810,I507825,I508122,I508139,I508165,I507813,I508187,I508204,I508221,I507828,I508252,I508269,I507819,I508300,I507822,I507834,I507831,I508389,I1279052,I508415,I508432,I508454,I508471,I1279064,I1279067,I508488,I1279070,I508514,I508522,I1279055,I508548,I508556,I1279061,I508573,I1279049,I508613,I508621,I508666,I1279073,I508683,I1279058,I508709,I508731,I508748,I508765,I508796,I508813,I508844,I508933,I1339290,I508959,I508976,I508925,I508998,I509015,I1339266,I1339287,I509032,I1339284,I509058,I509066,I1339263,I509092,I509100,I1339275,I509117,I508904,I1339278,I509157,I509165,I508898,I508913,I509210,I1339281,I1339269,I509227,I1339272,I509253,I508901,I509275,I509292,I509309,I508916,I509340,I509357,I508907,I509388,I508910,I508922,I508919,I509477,I509503,I509520,I509542,I509559,I509576,I509602,I509610,I509636,I509644,I509661,I509701,I509709,I509754,I509771,I509797,I509819,I509836,I509853,I509884,I509901,I509932,I510021,I510047,I510064,I510086,I510103,I510120,I510146,I510154,I510180,I510188,I510205,I510245,I510253,I510298,I510315,I510341,I510363,I510380,I510397,I510428,I510445,I510476,I510565,I559034,I510591,I510608,I510630,I510647,I559037,I559055,I510664,I559043,I510690,I510698,I510724,I510732,I559052,I510749,I559046,I510789,I510797,I510842,I559049,I559031,I510859,I559040,I510885,I510907,I510924,I510941,I510972,I510989,I511020,I511109,I952349,I511135,I511152,I511174,I511191,I952364,I952352,I511208,I952343,I511234,I511242,I952355,I511268,I511276,I952346,I511293,I952361,I511333,I511341,I511386,I952370,I952358,I511403,I952367,I511429,I511451,I511468,I511485,I511516,I511533,I511564,I511653,I511679,I511696,I511645,I511718,I511735,I511752,I511778,I511786,I511812,I511820,I511837,I511624,I511877,I511885,I511618,I511633,I511930,I511947,I511973,I511621,I511995,I512012,I512029,I511636,I512060,I512077,I511627,I512108,I511630,I511642,I511639,I512197,I1216424,I512223,I512240,I512189,I512262,I512279,I1216436,I512296,I1216427,I512322,I512330,I1216445,I512356,I512364,I1216421,I512381,I512168,I1216439,I512421,I512429,I512162,I512177,I512474,I1216433,I1216430,I512491,I1216442,I512517,I512165,I512539,I512556,I512573,I512180,I512604,I512621,I512171,I512652,I512174,I512186,I512183,I512741,I512767,I512784,I512733,I512806,I512823,I512840,I512866,I512874,I512900,I512908,I512925,I512712,I512965,I512973,I512706,I512721,I513018,I513035,I513061,I512709,I513083,I513100,I513117,I512724,I513148,I513165,I512715,I513196,I512718,I512730,I512727,I513285,I513311,I513328,I513350,I513367,I513384,I513410,I513418,I513444,I513452,I513469,I513509,I513517,I513562,I513579,I513605,I513627,I513644,I513661,I513692,I513709,I513740,I513829,I1380345,I513855,I513872,I513821,I513894,I513911,I1380321,I1380342,I513928,I1380339,I513954,I513962,I1380318,I513988,I513996,I1380330,I514013,I513800,I1380333,I514053,I514061,I513794,I513809,I514106,I1380336,I1380324,I514123,I1380327,I514149,I513797,I514171,I514188,I514205,I513812,I514236,I514253,I513803,I514284,I513806,I513818,I513815,I514373,I1361305,I514399,I514416,I514365,I514438,I514455,I1361281,I1361302,I514472,I1361299,I514498,I514506,I1361278,I514532,I514540,I1361290,I514557,I514344,I1361293,I514597,I514605,I514338,I514353,I514650,I1361296,I1361284,I514667,I1361287,I514693,I514341,I514715,I514732,I514749,I514356,I514780,I514797,I514347,I514828,I514350,I514362,I514359,I514917,I854282,I514943,I514960,I514909,I514982,I514999,I854276,I854273,I515016,I854288,I515042,I515050,I515076,I515084,I854270,I515101,I514888,I515141,I515149,I514882,I514897,I515194,I854285,I854279,I515211,I515237,I514885,I515259,I515276,I515293,I514900,I515324,I515341,I854291,I514891,I515372,I514894,I514906,I514903,I515461,I1310891,I515487,I515504,I515453,I515526,I515543,I1310888,I1310885,I515560,I1310873,I515586,I515594,I1310897,I515620,I515628,I1310882,I515645,I515432,I1310876,I515685,I515693,I515426,I515441,I515738,I1310879,I515755,I1310894,I515781,I515429,I515803,I515820,I515837,I515444,I515868,I515885,I515435,I515916,I515438,I515450,I515447,I516005,I738180,I516031,I516048,I515997,I516070,I516087,I738201,I738192,I516104,I516130,I516138,I738186,I516164,I516172,I738183,I516189,I515976,I738177,I516229,I516237,I515970,I515985,I516282,I738189,I516299,I738198,I516325,I515973,I516347,I516364,I516381,I515988,I516412,I516429,I738195,I515979,I516460,I515982,I515994,I515991,I516549,I1144752,I516575,I516592,I516614,I516631,I1144764,I516648,I1144755,I516674,I516682,I1144773,I516708,I516716,I1144749,I516733,I1144767,I516773,I516781,I516826,I1144761,I1144758,I516843,I1144770,I516869,I516891,I516908,I516925,I516956,I516973,I517004,I517093,I1007259,I517119,I517136,I517085,I517158,I517175,I1007274,I1007262,I517192,I1007253,I517218,I517226,I1007265,I517252,I517260,I1007256,I517277,I517064,I1007271,I517317,I517325,I517058,I517073,I517370,I1007280,I1007268,I517387,I1007277,I517413,I517061,I517435,I517452,I517469,I517076,I517500,I517517,I517067,I517548,I517070,I517082,I517079,I517637,I542374,I517663,I517680,I517702,I517719,I542377,I542395,I517736,I542383,I517762,I517770,I517796,I517804,I542392,I517821,I542386,I517861,I517869,I517914,I542389,I542371,I517931,I542380,I517957,I517979,I517996,I518013,I518044,I518061,I518092,I518181,I518207,I518224,I518173,I518246,I518263,I518280,I518306,I518314,I518340,I518348,I518365,I518152,I518405,I518413,I518146,I518161,I518458,I518475,I518501,I518149,I518523,I518540,I518557,I518164,I518588,I518605,I518155,I518636,I518158,I518170,I518167,I518725,I937491,I518751,I518768,I518717,I518790,I518807,I937506,I937494,I518824,I937485,I518850,I518858,I937497,I518884,I518892,I937488,I518909,I518696,I937503,I518949,I518957,I518690,I518705,I519002,I937512,I937500,I519019,I937509,I519045,I518693,I519067,I519084,I519101,I518708,I519132,I519149,I518699,I519180,I518702,I518714,I518711,I519269,I519295,I519312,I519261,I519334,I519351,I519368,I519394,I519402,I519428,I519436,I519453,I519240,I519493,I519501,I519234,I519249,I519546,I519563,I519589,I519237,I519611,I519628,I519645,I519252,I519676,I519693,I519243,I519724,I519246,I519258,I519255,I519813,I805806,I519839,I519856,I519878,I519895,I805827,I805818,I519912,I519938,I519946,I805812,I519972,I519980,I805809,I519997,I805803,I520037,I520045,I520090,I805815,I520107,I805824,I520133,I520155,I520172,I520189,I520220,I520237,I805821,I520268,I520357,I778640,I520383,I520400,I520349,I520422,I520439,I778661,I778652,I520456,I520482,I520490,I778646,I520516,I520524,I778643,I520541,I520328,I778637,I520581,I520589,I520322,I520337,I520634,I778649,I520651,I778658,I520677,I520325,I520699,I520716,I520733,I520340,I520764,I520781,I778655,I520331,I520812,I520334,I520346,I520343,I520901,I765346,I520927,I520944,I520966,I520983,I765367,I765358,I521000,I521026,I521034,I765352,I521060,I521068,I765349,I521085,I765343,I521125,I521133,I521178,I765355,I521195,I765364,I521221,I521243,I521260,I521277,I521308,I521325,I765361,I521356,I521445,I521471,I521488,I521437,I521510,I521527,I521544,I521570,I521578,I521604,I521612,I521629,I521416,I521669,I521677,I521410,I521425,I521722,I521739,I521765,I521413,I521787,I521804,I521821,I521428,I521852,I521869,I521419,I521900,I521422,I521434,I521431,I521989,I1316093,I522015,I522032,I521981,I522054,I522071,I1316090,I1316087,I522088,I1316075,I522114,I522122,I1316099,I522148,I522156,I1316084,I522173,I521960,I1316078,I522213,I522221,I521954,I521969,I522266,I1316081,I522283,I1316096,I522309,I521957,I522331,I522348,I522365,I521972,I522396,I522413,I521963,I522444,I521966,I521978,I521975,I522533,I522559,I522576,I522525,I522598,I522615,I522632,I522658,I522666,I522692,I522700,I522717,I522504,I522757,I522765,I522498,I522513,I522810,I522827,I522853,I522501,I522875,I522892,I522909,I522516,I522940,I522957,I522507,I522988,I522510,I522522,I522519,I523077,I971729,I523103,I523120,I523069,I523142,I523159,I971744,I971732,I523176,I971723,I523202,I523210,I971735,I523236,I523244,I971726,I523261,I523048,I971741,I523301,I523309,I523042,I523057,I523354,I971750,I971738,I523371,I971747,I523397,I523045,I523419,I523436,I523453,I523060,I523484,I523501,I523051,I523532,I523054,I523066,I523063,I523621,I789622,I523647,I523664,I523686,I523703,I789643,I789634,I523720,I523746,I523754,I789628,I523780,I523788,I789625,I523805,I789619,I523845,I523853,I523898,I789631,I523915,I789640,I523941,I523963,I523980,I523997,I524028,I524045,I789637,I524076,I524165,I1013073,I524191,I524208,I524157,I524230,I524247,I1013088,I1013076,I524264,I1013067,I524290,I524298,I1013079,I524324,I524332,I1013070,I524349,I524136,I1013085,I524389,I524397,I524130,I524145,I524442,I1013094,I1013082,I524459,I1013091,I524485,I524133,I524507,I524524,I524541,I524148,I524572,I524589,I524139,I524620,I524142,I524154,I524151,I524709,I524735,I524752,I524701,I524774,I524791,I524808,I524834,I524842,I524868,I524876,I524893,I524680,I524933,I524941,I524674,I524689,I524986,I525003,I525029,I524677,I525051,I525068,I525085,I524692,I525116,I525133,I524683,I525164,I524686,I524698,I524695,I525253,I837945,I525279,I525296,I525245,I525318,I525335,I837939,I837936,I525352,I837951,I525378,I525386,I525412,I525420,I837933,I525437,I525224,I525477,I525485,I525218,I525233,I525530,I837948,I837942,I525547,I525573,I525221,I525595,I525612,I525629,I525236,I525660,I525677,I837954,I525227,I525708,I525230,I525242,I525239,I525797,I881686,I525823,I525840,I525789,I525862,I525879,I881680,I881677,I525896,I881692,I525922,I525930,I525956,I525964,I881674,I525981,I525768,I526021,I526029,I525762,I525777,I526074,I881689,I881683,I526091,I526117,I525765,I526139,I526156,I526173,I525780,I526204,I526221,I881695,I525771,I526252,I525774,I525786,I525783,I526338,I862711,I526364,I526381,I862708,I526412,I526420,I526437,I526454,I862705,I526471,I862720,I526488,I526505,I526522,I526553,I862714,I526570,I862702,I526587,I526632,I526649,I526680,I862723,I526697,I526728,I526745,I862717,I526762,I526788,I526796,I526827,I526844,I526875,I526933,I837415,I526959,I526976,I526925,I837412,I527007,I527015,I527032,I527049,I837409,I527066,I837424,I527083,I527100,I527117,I526922,I527148,I837418,I527165,I837406,I527182,I526907,I526919,I527227,I527244,I526913,I527275,I837427,I527292,I526901,I527323,I527340,I837421,I527357,I527383,I527391,I526910,I527422,I527439,I526916,I527470,I526904,I527528,I679230,I527554,I527571,I679224,I527602,I527610,I679221,I527627,I527644,I679233,I527661,I679236,I527678,I527695,I527712,I527743,I679245,I527760,I679239,I527777,I527822,I527839,I527870,I679227,I527887,I527918,I679242,I527935,I527952,I527978,I527986,I528017,I528034,I528065,I528123,I528149,I528166,I528115,I528197,I528205,I528222,I528239,I528256,I528273,I528290,I528307,I528112,I528338,I528355,I528372,I528097,I528109,I528417,I528434,I528103,I528465,I528482,I528091,I528513,I528530,I528547,I528573,I528581,I528100,I528612,I528629,I528106,I528660,I528094,I528718,I835834,I528744,I528761,I528710,I835831,I528792,I528800,I528817,I528834,I835828,I528851,I835843,I528868,I528885,I528902,I528707,I528933,I835837,I528950,I835825,I528967,I528692,I528704,I529012,I529029,I528698,I529060,I835846,I529077,I528686,I529108,I529125,I835840,I529142,I529168,I529176,I528695,I529207,I529224,I528701,I529255,I528689,I529313,I529339,I529356,I529305,I529387,I529395,I529412,I529429,I529446,I529463,I529480,I529497,I529302,I529528,I529545,I529562,I529287,I529299,I529607,I529624,I529293,I529655,I529672,I529281,I529703,I529720,I529737,I529763,I529771,I529290,I529802,I529819,I529296,I529850,I529284,I529908,I1387458,I529934,I529951,I1387464,I529982,I529990,I1387479,I530007,I530024,I1387470,I530041,I1387467,I530058,I530075,I530092,I530123,I530140,I1387482,I530157,I530202,I530219,I530250,I1387476,I530267,I530298,I1387461,I530315,I1387473,I530332,I1387485,I530358,I530366,I530397,I530414,I530445,I530503,I599460,I530529,I530546,I599472,I530577,I530585,I599457,I530602,I530619,I599475,I530636,I599466,I530653,I530670,I530687,I530718,I599478,I530735,I599481,I530752,I530797,I530814,I530845,I530862,I530893,I599469,I530910,I599463,I530927,I530953,I530961,I530992,I531009,I531040,I531098,I531124,I531141,I531090,I531172,I531180,I531197,I531214,I531231,I531248,I531265,I531282,I531087,I531313,I531330,I531347,I531072,I531084,I531392,I531409,I531078,I531440,I531457,I531066,I531488,I531505,I531522,I531548,I531556,I531075,I531587,I531604,I531081,I531635,I531069,I531693,I531719,I531736,I531685,I531767,I531775,I531792,I531809,I531826,I531843,I531860,I531877,I531682,I531908,I531925,I531942,I531667,I531679,I531987,I532004,I531673,I532035,I532052,I531661,I532083,I532100,I532117,I532143,I532151,I531670,I532182,I532199,I531676,I532230,I531664,I532288,I1136675,I532314,I532331,I532280,I1136657,I532362,I532370,I1136663,I532387,I532404,I1136678,I532421,I1136669,I532438,I532455,I532472,I532277,I532503,I1136681,I532520,I1136660,I532537,I532262,I532274,I532582,I532599,I532268,I532630,I1136666,I532647,I532256,I532678,I1136672,I532695,I532712,I532738,I532746,I532265,I532777,I532794,I532271,I532825,I532259,I532883,I532909,I532926,I532875,I532957,I532965,I532982,I532999,I533016,I533033,I533050,I533067,I532872,I533098,I533115,I533132,I532857,I532869,I533177,I533194,I532863,I533225,I533242,I532851,I533273,I533290,I533307,I533333,I533341,I532860,I533372,I533389,I532866,I533420,I532854,I533478,I900655,I533504,I533521,I533470,I900652,I533552,I533560,I533577,I533594,I900649,I533611,I900664,I533628,I533645,I533662,I533467,I533693,I900658,I533710,I900646,I533727,I533452,I533464,I533772,I533789,I533458,I533820,I900667,I533837,I533446,I533868,I533885,I900661,I533902,I533928,I533936,I533455,I533967,I533984,I533461,I534015,I533449,I534073,I1103151,I534099,I534116,I534065,I1103133,I534147,I534155,I1103139,I534172,I534189,I1103154,I534206,I1103145,I534223,I534240,I534257,I534062,I534288,I1103157,I534305,I1103136,I534322,I534047,I534059,I534367,I534384,I534053,I534415,I1103142,I534432,I534041,I534463,I1103148,I534480,I534497,I534523,I534531,I534050,I534562,I534579,I534056,I534610,I534044,I534668,I534694,I534711,I534660,I534742,I534750,I534767,I534784,I534801,I534818,I534835,I534852,I534657,I534883,I534900,I534917,I534642,I534654,I534962,I534979,I534648,I535010,I535027,I534636,I535058,I535075,I535092,I535118,I535126,I534645,I535157,I535174,I534651,I535205,I534639,I535263,I535289,I535306,I535337,I535345,I535362,I535379,I535396,I535413,I535430,I535447,I535478,I535495,I535512,I535557,I535574,I535605,I535622,I535653,I535670,I535687,I535713,I535721,I535752,I535769,I535800,I535858,I535884,I535901,I535850,I535932,I535940,I535957,I535974,I535991,I536008,I536025,I536042,I535847,I536073,I536090,I536107,I535832,I535844,I536152,I536169,I535838,I536200,I536217,I535826,I536248,I536265,I536282,I536308,I536316,I535835,I536347,I536364,I535841,I536395,I535829,I536453,I597148,I536479,I536496,I597160,I536527,I536535,I597145,I536552,I536569,I597163,I536586,I597154,I536603,I536620,I536637,I536668,I597166,I536685,I597169,I536702,I536747,I536764,I536795,I536812,I536843,I597157,I536860,I597151,I536877,I536903,I536911,I536942,I536959,I536990,I537048,I537074,I537091,I537040,I537122,I537130,I537147,I537164,I537181,I537198,I537215,I537232,I537037,I537263,I537280,I537297,I537022,I537034,I537342,I537359,I537028,I537390,I537407,I537016,I537438,I537455,I537472,I537498,I537506,I537025,I537537,I537554,I537031,I537585,I537019,I537643,I537669,I537686,I537635,I537717,I537725,I537742,I537759,I537776,I537793,I537810,I537827,I537632,I537858,I537875,I537892,I537617,I537629,I537937,I537954,I537623,I537985,I538002,I537611,I538033,I538050,I538067,I538093,I538101,I537620,I538132,I538149,I537626,I538180,I537614,I538238,I866400,I538264,I538281,I866397,I538312,I538320,I538337,I538354,I866394,I538371,I866409,I538388,I538405,I538422,I538453,I866403,I538470,I866391,I538487,I538532,I538549,I538580,I866412,I538597,I538628,I538645,I866406,I538662,I538688,I538696,I538727,I538744,I538775,I538833,I538859,I538876,I538825,I538907,I538915,I538932,I538949,I538966,I538983,I539000,I539017,I538822,I539048,I539065,I539082,I538807,I538819,I539127,I539144,I538813,I539175,I539192,I538801,I539223,I539240,I539257,I539283,I539291,I538810,I539322,I539339,I538816,I539370,I538804,I539428,I1126271,I539454,I539471,I539420,I1126253,I539502,I539510,I1126259,I539527,I539544,I1126274,I539561,I1126265,I539578,I539595,I539612,I539417,I539643,I1126277,I539660,I1126256,I539677,I539402,I539414,I539722,I539739,I539408,I539770,I1126262,I539787,I539396,I539818,I1126268,I539835,I539852,I539878,I539886,I539405,I539917,I539934,I539411,I539965,I539399,I540023,I540049,I540066,I540097,I540105,I540122,I540139,I540156,I540173,I540190,I540207,I540238,I540255,I540272,I540317,I540334,I540365,I540382,I540413,I540430,I540447,I540473,I540481,I540512,I540529,I540560,I540618,I779802,I540644,I540661,I779796,I540692,I540700,I779793,I540717,I540734,I779805,I540751,I779808,I540768,I540785,I540802,I540833,I779817,I540850,I779811,I540867,I540912,I540929,I540960,I779799,I540977,I541008,I779814,I541025,I541042,I541068,I541076,I541107,I541124,I541155,I541213,I1319552,I541239,I541256,I1319558,I541287,I541295,I1319546,I541312,I541329,I1319549,I541346,I1319555,I541363,I541380,I541397,I541428,I541445,I1319564,I541462,I541507,I541524,I541555,I1319543,I541572,I541603,I1319567,I541620,I541637,I1319561,I541663,I541671,I541702,I541719,I541750,I541808,I541834,I541851,I541882,I541890,I541907,I541924,I541941,I541958,I541975,I541992,I542023,I542040,I542057,I542102,I542119,I542150,I542167,I542198,I542215,I542232,I542258,I542266,I542297,I542314,I542345,I542403,I691946,I542429,I542446,I691940,I542477,I542485,I691937,I542502,I542519,I691949,I542536,I691952,I542553,I542570,I542587,I542618,I691961,I542635,I691955,I542652,I542697,I542714,I542745,I691943,I542762,I542793,I691958,I542810,I542827,I542853,I542861,I542892,I542909,I542940,I542998,I543024,I543041,I542990,I543072,I543080,I543097,I543114,I543131,I543148,I543165,I543182,I542987,I543213,I543230,I543247,I542972,I542984,I543292,I543309,I542978,I543340,I543357,I542966,I543388,I543405,I543422,I543448,I543456,I542975,I543487,I543504,I542981,I543535,I542969,I543593,I655526,I543619,I543636,I655538,I543667,I543675,I655523,I543692,I543709,I655541,I543726,I655532,I543743,I543760,I543777,I543808,I655544,I543825,I655547,I543842,I543887,I543904,I543935,I543952,I543983,I655535,I544000,I655529,I544017,I544043,I544051,I544082,I544099,I544130,I544188,I1355923,I544214,I544231,I544180,I1355929,I544262,I544270,I1355944,I544287,I544304,I1355935,I544321,I1355932,I544338,I544355,I544372,I544177,I544403,I544420,I1355947,I544437,I544162,I544174,I544482,I544499,I544168,I544530,I1355941,I544547,I544156,I544578,I1355926,I544595,I1355938,I544612,I1355950,I544638,I544646,I544165,I544677,I544694,I544171,I544725,I544159,I544783,I1119913,I544809,I544826,I544775,I1119895,I544857,I544865,I1119901,I544882,I544899,I1119916,I544916,I1119907,I544933,I544950,I544967,I544772,I544998,I1119919,I545015,I1119898,I545032,I544757,I544769,I545077,I545094,I544763,I545125,I1119904,I545142,I544751,I545173,I1119910,I545190,I545207,I545233,I545241,I544760,I545272,I545289,I544766,I545320,I544754,I545378,I645122,I545404,I545421,I545370,I645134,I545452,I545460,I645119,I545477,I545494,I645137,I545511,I645128,I545528,I545545,I545562,I545367,I545593,I645140,I545610,I645143,I545627,I545352,I545364,I545672,I545689,I545358,I545720,I545737,I545346,I545768,I645131,I545785,I645125,I545802,I545828,I545836,I545355,I545867,I545884,I545361,I545915,I545349,I545973,I545999,I546016,I545965,I546047,I546055,I546072,I546089,I546106,I546123,I546140,I546157,I545962,I546188,I546205,I546222,I545947,I545959,I546267,I546284,I545953,I546315,I546332,I545941,I546363,I546380,I546397,I546423,I546431,I545950,I546462,I546479,I545956,I546510,I545944,I546568,I1000808,I546594,I546611,I546560,I1000796,I546642,I546650,I1000793,I546667,I546684,I1000805,I546701,I1000802,I546718,I546735,I546752,I546557,I546783,I1000811,I546800,I1000814,I546817,I546542,I546554,I546862,I546879,I546548,I546910,I1000817,I546927,I546536,I546958,I1000820,I546975,I1000799,I546992,I547018,I547026,I546545,I547057,I547074,I546551,I547105,I546539,I547163,I547189,I547206,I547237,I547245,I547262,I547279,I547296,I547313,I547330,I547347,I547378,I547395,I547412,I547457,I547474,I547505,I547522,I547553,I547570,I547587,I547613,I547621,I547652,I547669,I547700,I547758,I547784,I547801,I547750,I547832,I547840,I547857,I547874,I547891,I547908,I547925,I547942,I547747,I547973,I547990,I548007,I547732,I547744,I548052,I548069,I547738,I548100,I548117,I547726,I548148,I548165,I548182,I548208,I548216,I547735,I548247,I548264,I547741,I548295,I547729,I548353,I548379,I548396,I548345,I548427,I548435,I548452,I548469,I548486,I548503,I548520,I548537,I548342,I548568,I548585,I548602,I548327,I548339,I548647,I548664,I548333,I548695,I548712,I548321,I548743,I548760,I548777,I548803,I548811,I548330,I548842,I548859,I548336,I548890,I548324,I548948,I940084,I548974,I548991,I548940,I940072,I549022,I549030,I940069,I549047,I549064,I940081,I549081,I940078,I549098,I549115,I549132,I548937,I549163,I940087,I549180,I940090,I549197,I548922,I548934,I549242,I549259,I548928,I549290,I940093,I549307,I548916,I549338,I940096,I549355,I940075,I549372,I549398,I549406,I548925,I549437,I549454,I548931,I549485,I548919,I549543,I944606,I549569,I549586,I549535,I944594,I549617,I549625,I944591,I549642,I549659,I944603,I549676,I944600,I549693,I549710,I549727,I549532,I549758,I944609,I549775,I944612,I549792,I549517,I549529,I549837,I549854,I549523,I549885,I944615,I549902,I549511,I549933,I944618,I549950,I944597,I549967,I549993,I550001,I549520,I550032,I550049,I549526,I550080,I549514,I550138,I894858,I550164,I550181,I894855,I550212,I550220,I550237,I550254,I894852,I550271,I894867,I550288,I550305,I550322,I550353,I894861,I550370,I894849,I550387,I550432,I550449,I550480,I894870,I550497,I550528,I550545,I894864,I550562,I550588,I550596,I550627,I550644,I550675,I550733,I690790,I550759,I550776,I550725,I690784,I550807,I550815,I690781,I550832,I550849,I690793,I550866,I690796,I550883,I550900,I550917,I550722,I550948,I690805,I550965,I690799,I550982,I550707,I550719,I551027,I551044,I550713,I551075,I690787,I551092,I550701,I551123,I690802,I551140,I551157,I551183,I551191,I550710,I551222,I551239,I550716,I551270,I550704,I551328,I659000,I551354,I551371,I551320,I658994,I551402,I551410,I658991,I551427,I551444,I659003,I551461,I659006,I551478,I551495,I551512,I551317,I551543,I659015,I551560,I659009,I551577,I551302,I551314,I551622,I551639,I551308,I551670,I658997,I551687,I551296,I551718,I659012,I551735,I551752,I551778,I551786,I551305,I551817,I551834,I551311,I551865,I551299,I551923,I740498,I551949,I551966,I740492,I551997,I552005,I740489,I552022,I552039,I740501,I552056,I740504,I552073,I552090,I552107,I552138,I740513,I552155,I740507,I552172,I552217,I552234,I552265,I740495,I552282,I552313,I740510,I552330,I552347,I552373,I552381,I552412,I552429,I552460,I552518,I697148,I552544,I552561,I552510,I697142,I552592,I552600,I697139,I552617,I552634,I697151,I552651,I697154,I552668,I552685,I552702,I552507,I552733,I697163,I552750,I697157,I552767,I552492,I552504,I552812,I552829,I552498,I552860,I697145,I552877,I552486,I552908,I697160,I552925,I552942,I552968,I552976,I552495,I553007,I553024,I552501,I553055,I552489,I553113,I857441,I553139,I553156,I553105,I857438,I553187,I553195,I553212,I553229,I857435,I553246,I857450,I553263,I553280,I553297,I553102,I553328,I857444,I553345,I857432,I553362,I553087,I553099,I553407,I553424,I553093,I553455,I857453,I553472,I553081,I553503,I553520,I857447,I553537,I553563,I553571,I553090,I553602,I553619,I553096,I553650,I553084,I553708,I553734,I553751,I553782,I553790,I553807,I553824,I553841,I553858,I553875,I553892,I553923,I553940,I553957,I554002,I554019,I554050,I554067,I554098,I554115,I554132,I554158,I554166,I554197,I554214,I554245,I554303,I1044090,I554329,I554346,I554295,I1044078,I554377,I554385,I1044075,I554402,I554419,I1044087,I554436,I1044084,I554453,I554470,I554487,I554292,I554518,I1044093,I554535,I1044096,I554552,I554277,I554289,I554597,I554614,I554283,I554645,I1044099,I554662,I554271,I554693,I1044102,I554710,I1044081,I554727,I554753,I554761,I554280,I554792,I554809,I554286,I554840,I554274,I554898,I1149969,I554924,I554941,I554890,I1149951,I554972,I554980,I1149957,I554997,I555014,I1149972,I555031,I1149963,I555048,I555065,I555082,I554887,I555113,I1149975,I555130,I1149954,I555147,I554872,I554884,I555192,I555209,I554878,I555240,I1149960,I555257,I554866,I555288,I1149966,I555305,I555322,I555348,I555356,I554875,I555387,I555404,I554881,I555435,I554869,I555493,I555519,I555536,I555567,I555575,I555592,I555609,I555626,I555643,I555660,I555677,I555708,I555725,I555742,I555787,I555804,I555835,I555852,I555883,I555900,I555917,I555943,I555951,I555982,I555999,I556030,I556088,I1213549,I556114,I556131,I1213531,I556162,I556170,I1213537,I556187,I556204,I1213552,I556221,I1213543,I556238,I556255,I556272,I556303,I1213555,I556320,I1213534,I556337,I556382,I556399,I556430,I1213540,I556447,I556478,I1213546,I556495,I556512,I556538,I556546,I556577,I556594,I556625,I556683,I712754,I556709,I556726,I556675,I712748,I556757,I556765,I712745,I556782,I556799,I712757,I556816,I712760,I556833,I556850,I556867,I556672,I556898,I712769,I556915,I712763,I556932,I556657,I556669,I556977,I556994,I556663,I557025,I712751,I557042,I556651,I557073,I712766,I557090,I557107,I557133,I557141,I556660,I557172,I557189,I556666,I557220,I556654,I557278,I715644,I557304,I557321,I557270,I715638,I557352,I557360,I715635,I557377,I557394,I715647,I557411,I715650,I557428,I557445,I557462,I557267,I557493,I715659,I557510,I715653,I557527,I557252,I557264,I557572,I557589,I557258,I557620,I715641,I557637,I557246,I557668,I715656,I557685,I557702,I557728,I557736,I557255,I557767,I557784,I557261,I557815,I557249,I557873,I557899,I557916,I557865,I557947,I557955,I557972,I557989,I558006,I558023,I558040,I558057,I557862,I558088,I558105,I558122,I557847,I557859,I558167,I558184,I557853,I558215,I558232,I557841,I558263,I558280,I558297,I558323,I558331,I557850,I558362,I558379,I557856,I558410,I557844,I558468,I558494,I558511,I558460,I558542,I558550,I558567,I558584,I558601,I558618,I558635,I558652,I558457,I558683,I558700,I558717,I558442,I558454,I558762,I558779,I558448,I558810,I558827,I558436,I558858,I558875,I558892,I558918,I558926,I558445,I558957,I558974,I558451,I559005,I558439,I559063,I1084807,I559089,I559106,I1084810,I559137,I559145,I1084813,I559162,I559179,I1084825,I559196,I1084816,I559213,I559230,I559247,I559278,I1084822,I559295,I559312,I559357,I559374,I559405,I559422,I559453,I1084819,I559470,I559487,I1084828,I559513,I559521,I559552,I559569,I559600,I559658,I559684,I559701,I559650,I559732,I559740,I559757,I559774,I559791,I559808,I559825,I559842,I559647,I559873,I559890,I559907,I559632,I559644,I559952,I559969,I559638,I560000,I560017,I559626,I560048,I560065,I560082,I560108,I560116,I559635,I560147,I560164,I559641,I560195,I559629,I560253,I560279,I560296,I560245,I560327,I560335,I560352,I560369,I560386,I560403,I560420,I560437,I560242,I560468,I560485,I560502,I560227,I560239,I560547,I560564,I560233,I560595,I560612,I560221,I560643,I560660,I560677,I560703,I560711,I560230,I560742,I560759,I560236,I560790,I560224,I560848,I880102,I560874,I560891,I560840,I880099,I560922,I560930,I560947,I560964,I880096,I560981,I880111,I560998,I561015,I561032,I560837,I561063,I880105,I561080,I880093,I561097,I560822,I560834,I561142,I561159,I560828,I561190,I880114,I561207,I560816,I561238,I561255,I880108,I561272,I561298,I561306,I560825,I561337,I561354,I560831,I561385,I560819,I561443,I561469,I561486,I561435,I561517,I561525,I561542,I561559,I561576,I561593,I561610,I561627,I561432,I561658,I561675,I561692,I561417,I561429,I561737,I561754,I561423,I561785,I561802,I561411,I561833,I561850,I561867,I561893,I561901,I561420,I561932,I561949,I561426,I561980,I561414,I562038,I1232623,I562064,I562081,I1232605,I562112,I562120,I1232611,I562137,I562154,I1232626,I562171,I1232617,I562188,I562205,I562222,I562253,I1232629,I562270,I1232608,I562287,I562332,I562349,I562380,I1232614,I562397,I562428,I1232620,I562445,I562462,I562488,I562496,I562527,I562544,I562575,I562633,I609864,I562659,I562676,I609876,I562707,I562715,I609861,I562732,I562749,I609879,I562766,I609870,I562783,I562800,I562817,I562848,I609882,I562865,I609885,I562882,I562927,I562944,I562975,I562992,I563023,I609873,I563040,I609867,I563057,I563083,I563091,I563122,I563139,I563170,I563228,I563254,I563271,I563220,I563302,I563310,I563327,I563344,I563361,I563378,I563395,I563412,I563217,I563443,I563460,I563477,I563202,I563214,I563522,I563539,I563208,I563570,I563587,I563196,I563618,I563635,I563652,I563678,I563686,I563205,I563717,I563734,I563211,I563765,I563199,I563823,I705818,I563849,I563866,I563815,I705812,I563897,I563905,I705809,I563922,I563939,I705821,I563956,I705824,I563973,I563990,I564007,I563812,I564038,I705833,I564055,I705827,I564072,I563797,I563809,I564117,I564134,I563803,I564165,I705815,I564182,I563791,I564213,I705830,I564230,I564247,I564273,I564281,I563800,I564312,I564329,I563806,I564360,I563794,I564418,I1310304,I564444,I564461,I564410,I1310310,I564492,I564500,I1310298,I564517,I564534,I1310301,I564551,I1310307,I564568,I564585,I564602,I564407,I564633,I564650,I1310316,I564667,I564392,I564404,I564712,I564729,I564398,I564760,I1310295,I564777,I564386,I564808,I1310319,I564825,I564842,I1310313,I564868,I564876,I564395,I564907,I564924,I564401,I564955,I564389,I565013,I565039,I565056,I565087,I565095,I565112,I565129,I565146,I565163,I565180,I565197,I565228,I565245,I565262,I565307,I565324,I565355,I565372,I565403,I565420,I565437,I565463,I565471,I565502,I565519,I565550,I565608,I964632,I565634,I565651,I964620,I565682,I565690,I964617,I565707,I565724,I964629,I565741,I964626,I565758,I565775,I565792,I565823,I964635,I565840,I964638,I565857,I565902,I565919,I565950,I964641,I565967,I565998,I964644,I566015,I964623,I566032,I566058,I566066,I566097,I566114,I566145,I566203,I566229,I566246,I566195,I566277,I566285,I566302,I566319,I566336,I566353,I566370,I566387,I566192,I566418,I566435,I566452,I566177,I566189,I566497,I566514,I566183,I566545,I566562,I566171,I566593,I566610,I566627,I566653,I566661,I566180,I566692,I566709,I566186,I566740,I566174,I566798,I667670,I566824,I566841,I566790,I667664,I566872,I566880,I667661,I566897,I566914,I667673,I566931,I667676,I566948,I566965,I566982,I566787,I567013,I667685,I567030,I667679,I567047,I566772,I566784,I567092,I567109,I566778,I567140,I667667,I567157,I566766,I567188,I667682,I567205,I567222,I567248,I567256,I566775,I567287,I567304,I566781,I567335,I566769,I567393,I567419,I567436,I567385,I567467,I567475,I567492,I567509,I567526,I567543,I567560,I567577,I567382,I567608,I567625,I567642,I567367,I567379,I567687,I567704,I567373,I567735,I567752,I567361,I567783,I567800,I567817,I567843,I567851,I567370,I567882,I567899,I567376,I567930,I567364,I567988,I960110,I568014,I568031,I567980,I960098,I568062,I568070,I960095,I568087,I568104,I960107,I568121,I960104,I568138,I568155,I568172,I567977,I568203,I960113,I568220,I960116,I568237,I567962,I567974,I568282,I568299,I567968,I568330,I960119,I568347,I567956,I568378,I960122,I568395,I960101,I568412,I568438,I568446,I567965,I568477,I568494,I567971,I568525,I567959,I568583,I761884,I568609,I568626,I568575,I761878,I568657,I568665,I761875,I568682,I568699,I761887,I568716,I761890,I568733,I568750,I568767,I568572,I568798,I761899,I568815,I761893,I568832,I568557,I568569,I568877,I568894,I568563,I568925,I761881,I568942,I568551,I568973,I761896,I568990,I569007,I569033,I569041,I568560,I569072,I569089,I568566,I569120,I568554,I569178,I1244183,I569204,I569221,I569170,I1244165,I569252,I569260,I1244171,I569277,I569294,I1244186,I569311,I1244177,I569328,I569345,I569362,I569167,I569393,I1244189,I569410,I1244168,I569427,I569152,I569164,I569472,I569489,I569158,I569520,I1244174,I569537,I569146,I569568,I1244180,I569585,I569602,I569628,I569636,I569155,I569667,I569684,I569161,I569715,I569149,I569773,I1020188,I569799,I569816,I569765,I1020176,I569847,I569855,I1020173,I569872,I569889,I1020185,I569906,I1020182,I569923,I569940,I569957,I569762,I569988,I1020191,I570005,I1020194,I570022,I569747,I569759,I570067,I570084,I569753,I570115,I1020197,I570132,I569741,I570163,I1020200,I570180,I1020179,I570197,I570223,I570231,I569750,I570262,I570279,I569756,I570310,I569744,I570368,I570394,I570411,I570360,I570442,I570450,I570467,I570484,I570501,I570518,I570535,I570552,I570357,I570583,I570600,I570617,I570342,I570354,I570662,I570679,I570348,I570710,I570727,I570336,I570758,I570775,I570792,I570818,I570826,I570345,I570857,I570874,I570351,I570905,I570339,I570963,I809280,I570989,I571006,I809274,I571037,I571045,I809271,I571062,I571079,I809283,I571096,I809286,I571113,I571130,I571147,I571178,I809295,I571195,I809289,I571212,I571257,I571274,I571305,I809277,I571322,I571353,I809292,I571370,I571387,I571413,I571421,I571452,I571469,I571500,I571558,I1042798,I571584,I571601,I571550,I1042786,I571632,I571640,I1042783,I571657,I571674,I1042795,I571691,I1042792,I571708,I571725,I571742,I571547,I571773,I1042801,I571790,I1042804,I571807,I571532,I571544,I571852,I571869,I571538,I571900,I1042807,I571917,I571526,I571948,I1042810,I571965,I1042789,I571982,I572008,I572016,I571535,I572047,I572064,I571541,I572095,I571529,I572153,I572179,I572196,I572145,I572227,I572235,I572252,I572269,I572286,I572303,I572320,I572337,I572142,I572368,I572385,I572402,I572127,I572139,I572447,I572464,I572133,I572495,I572512,I572121,I572543,I572560,I572577,I572603,I572611,I572130,I572642,I572659,I572136,I572690,I572124,I572748,I1261097,I572774,I572791,I572740,I1261112,I572822,I572830,I1261121,I572847,I572864,I1261100,I572881,I1261106,I572898,I572915,I572932,I572737,I572963,I1261118,I572980,I1261115,I572997,I572722,I572734,I573042,I573059,I572728,I573090,I573107,I572716,I573138,I1261109,I573155,I1261103,I573172,I573198,I573206,I572725,I573237,I573254,I572731,I573285,I572719,I573343,I573369,I573386,I573417,I573425,I573442,I573459,I573476,I573493,I573510,I573527,I573558,I573575,I573592,I573637,I573654,I573685,I573702,I573733,I573750,I573767,I573793,I573801,I573832,I573849,I573880,I573938,I573964,I573981,I573930,I574012,I574020,I574037,I574054,I574071,I574088,I574105,I574122,I573927,I574153,I574170,I574187,I573912,I573924,I574232,I574249,I573918,I574280,I574297,I573906,I574328,I574345,I574362,I574388,I574396,I573915,I574427,I574444,I573921,I574475,I573909,I574533,I931686,I574559,I574576,I574525,I931674,I574607,I574615,I931671,I574632,I574649,I931683,I574666,I931680,I574683,I574700,I574717,I574522,I574748,I931689,I574765,I931692,I574782,I574507,I574519,I574827,I574844,I574513,I574875,I931695,I574892,I574501,I574923,I931698,I574940,I931677,I574957,I574983,I574991,I574510,I575022,I575039,I574516,I575070,I574504,I575128,I1203723,I575154,I575171,I575120,I1203705,I575202,I575210,I1203711,I575227,I575244,I1203726,I575261,I1203717,I575278,I575295,I575312,I575117,I575343,I1203729,I575360,I1203708,I575377,I575102,I575114,I575422,I575439,I575108,I575470,I1203714,I575487,I575096,I575518,I1203720,I575535,I575552,I575578,I575586,I575105,I575617,I575634,I575111,I575665,I575099,I575723,I575749,I575766,I575715,I575797,I575805,I575822,I575839,I575856,I575873,I575890,I575907,I575712,I575938,I575955,I575972,I575697,I575709,I576017,I576034,I575703,I576065,I576082,I575691,I576113,I576130,I576147,I576173,I576181,I575700,I576212,I576229,I575706,I576260,I575694,I576318,I1329231,I576344,I576361,I1329237,I576392,I576400,I1329240,I576417,I576434,I1329243,I576451,I1329228,I576468,I576485,I576502,I576533,I1329234,I576550,I1329216,I576567,I576612,I576629,I576660,I576677,I576708,I1329225,I576725,I1329222,I576742,I1329219,I576768,I576776,I576807,I576824,I576855,I576913,I834780,I576939,I576956,I576905,I834777,I576987,I576995,I577012,I577029,I834774,I577046,I834789,I577063,I577080,I577097,I576902,I577128,I834783,I577145,I834771,I577162,I576887,I576899,I577207,I577224,I576893,I577255,I834792,I577272,I576881,I577303,I577320,I834786,I577337,I577363,I577371,I576890,I577402,I577419,I576896,I577450,I576884,I577508,I1076392,I577534,I577551,I577500,I1076395,I577582,I577590,I1076398,I577607,I577624,I1076410,I577641,I1076401,I577658,I577675,I577692,I577497,I577723,I1076407,I577740,I577757,I577482,I577494,I577802,I577819,I577488,I577850,I577867,I577476,I577898,I1076404,I577915,I577932,I1076413,I577958,I577966,I577485,I577997,I578014,I577491,I578045,I577479,I578103,I578129,I578137,I578163,I578171,I578188,I578205,I578222,I578239,I578270,I578287,I578304,I578321,I578366,I578411,I578428,I578445,I578476,I578493,I578510,I578536,I578544,I578589,I578606,I578623,I578681,I578707,I578715,I578741,I578749,I578766,I578783,I578800,I578817,I578848,I578865,I578882,I578899,I578944,I578989,I579006,I579023,I579054,I579071,I579088,I579114,I579122,I579167,I579184,I579201,I579259,I915527,I579285,I579293,I915524,I579319,I579327,I915521,I579344,I915548,I579361,I579378,I915536,I579395,I579245,I579426,I579443,I579460,I915542,I579477,I915533,I579242,I579233,I579522,I579236,I579230,I579567,I915530,I579584,I579601,I579239,I579632,I915545,I579649,I915539,I579666,I579692,I579700,I579227,I579251,I579745,I579762,I579779,I579248,I579837,I1315509,I579863,I579871,I1315521,I579897,I579905,I1315512,I579922,I1315500,I579939,I579956,I1315497,I579973,I579823,I580004,I580021,I580038,I1315503,I580055,I579820,I579811,I580100,I579814,I579808,I580145,I1315518,I580162,I580179,I579817,I580210,I1315506,I580227,I580244,I1315515,I580270,I580278,I579805,I579829,I580323,I580340,I580357,I579826,I580415,I1298747,I580441,I580449,I1298759,I580475,I580483,I1298750,I580500,I1298738,I580517,I580534,I1298735,I580551,I580582,I580599,I580616,I1298741,I580633,I580678,I580723,I1298756,I580740,I580757,I580788,I1298744,I580805,I580822,I1298753,I580848,I580856,I580901,I580918,I580935,I580993,I726617,I581019,I581027,I726629,I581053,I581061,I726620,I581078,I726623,I581095,I581112,I726626,I581129,I580979,I581160,I581177,I581194,I581211,I726632,I580976,I580967,I581256,I580970,I580964,I581301,I726638,I581318,I581335,I580973,I581366,I581383,I726635,I581400,I726641,I581426,I581434,I580961,I580985,I581479,I581496,I581513,I580982,I581571,I1235495,I581597,I581605,I1235501,I581631,I581639,I581656,I1235498,I581673,I581690,I1235516,I581707,I581557,I581738,I581755,I581772,I1235519,I581789,I581554,I581545,I581834,I581548,I581542,I581879,I1235504,I581896,I581913,I581551,I581944,I1235510,I581961,I1235507,I581978,I1235513,I582004,I582012,I581539,I581563,I582057,I582074,I582091,I581560,I582149,I582175,I582183,I582209,I582217,I582234,I582251,I582268,I582285,I582316,I582333,I582350,I582367,I582412,I582457,I582474,I582491,I582522,I582539,I582556,I582582,I582590,I582635,I582652,I582669,I582727,I582753,I582761,I582787,I582795,I582812,I582829,I582846,I582863,I582713,I582894,I582911,I582928,I582945,I582710,I582701,I582990,I582704,I582698,I583035,I583052,I583069,I582707,I583100,I583117,I583134,I583160,I583168,I582695,I582719,I583213,I583230,I583247,I582716,I583305,I1064071,I583331,I583339,I1064062,I583365,I583373,I1064056,I583390,I1064068,I583407,I583424,I1064059,I583441,I583291,I583472,I583489,I583506,I1064065,I583523,I1064050,I583288,I583279,I583568,I583282,I583276,I583613,I583630,I583647,I583285,I583678,I1064053,I583695,I583712,I583738,I583746,I583273,I583297,I583791,I583808,I583825,I583294,I583883,I583909,I583917,I583943,I583951,I583968,I583985,I584002,I584019,I583869,I584050,I584067,I584084,I584101,I583866,I583857,I584146,I583860,I583854,I584191,I584208,I584225,I583863,I584256,I584273,I584290,I584316,I584324,I583851,I583875,I584369,I584386,I584403,I583872,I584461,I584487,I584495,I584521,I584529,I584546,I584563,I584580,I584597,I584447,I584628,I584645,I584662,I584679,I584444,I584435,I584724,I584438,I584432,I584769,I584786,I584803,I584441,I584834,I584851,I584868,I584894,I584902,I584429,I584453,I584947,I584964,I584981,I584450,I585039,I585065,I585073,I585099,I585107,I585124,I585141,I585158,I585175,I585025,I585206,I585223,I585240,I585257,I585022,I585013,I585302,I585016,I585010,I585347,I585364,I585381,I585019,I585412,I585429,I585446,I585472,I585480,I585007,I585031,I585525,I585542,I585559,I585028,I585617,I743379,I585643,I585651,I743391,I585677,I585685,I743382,I585702,I743385,I585719,I585736,I743388,I585753,I585603,I585784,I585801,I585818,I585835,I743394,I585600,I585591,I585880,I585594,I585588,I585925,I743400,I585942,I585959,I585597,I585990,I586007,I743397,I586024,I743403,I586050,I586058,I585585,I585609,I586103,I586120,I586137,I585606,I586195,I586221,I586229,I586255,I586263,I586280,I586297,I586314,I586331,I586362,I586379,I586396,I586413,I586458,I586503,I586520,I586537,I586568,I586585,I586602,I586628,I586636,I586681,I586698,I586715,I586773,I586799,I586807,I586833,I586841,I586858,I586875,I586892,I586909,I586940,I586957,I586974,I586991,I587036,I587081,I587098,I587115,I587146,I587163,I587180,I587206,I587214,I587259,I587276,I587293,I587351,I587377,I587385,I587411,I587419,I587436,I587453,I587470,I587487,I587518,I587535,I587552,I587569,I587614,I587659,I587676,I587693,I587724,I587741,I587758,I587784,I587792,I587837,I587854,I587871,I587929,I587955,I587963,I587989,I587997,I588014,I588031,I588048,I588065,I587915,I588096,I588113,I588130,I588147,I587912,I587903,I588192,I587906,I587900,I588237,I588254,I588271,I587909,I588302,I588319,I588336,I588362,I588370,I587897,I587921,I588415,I588432,I588449,I587918,I588507,I588533,I588541,I588567,I588575,I588592,I588609,I588626,I588643,I588493,I588674,I588691,I588708,I588725,I588490,I588481,I588770,I588484,I588478,I588815,I588832,I588849,I588487,I588880,I588897,I588914,I588940,I588948,I588475,I588499,I588993,I589010,I589027,I588496,I589085,I664771,I589111,I589119,I664783,I589145,I589153,I664774,I589170,I664777,I589187,I589204,I664780,I589221,I589252,I589269,I589286,I589303,I664786,I589348,I589393,I664792,I589410,I589427,I589458,I589475,I664789,I589492,I664795,I589518,I589526,I589571,I589588,I589605,I589663,I589689,I589697,I589723,I589731,I589748,I589765,I589782,I589799,I589649,I589830,I589847,I589864,I589881,I589646,I589637,I589926,I589640,I589634,I589971,I589988,I590005,I589643,I590036,I590053,I590070,I590096,I590104,I589631,I589655,I590149,I590166,I590183,I589652,I590241,I1106023,I590267,I590275,I1106029,I590301,I590309,I590326,I1106026,I590343,I590360,I1106044,I590377,I590227,I590408,I590425,I590442,I1106047,I590459,I590224,I590215,I590504,I590218,I590212,I590549,I1106032,I590566,I590583,I590221,I590614,I1106038,I590631,I1106035,I590648,I1106041,I590674,I590682,I590209,I590233,I590727,I590744,I590761,I590230,I590819,I1358303,I590845,I590853,I590879,I590887,I1358327,I590904,I1358309,I590921,I590938,I1358324,I590955,I590805,I590986,I591003,I591020,I1358306,I591037,I1358315,I590802,I590793,I591082,I590796,I590790,I591127,I1358312,I591144,I591161,I590799,I591192,I1358321,I591209,I1358330,I591226,I1358318,I591252,I591260,I590787,I590811,I591305,I591322,I591339,I590808,I591397,I1160355,I591423,I591431,I1160361,I591457,I591465,I591482,I1160358,I591499,I591516,I1160376,I591533,I591564,I591581,I591598,I1160379,I591615,I591660,I591705,I1160364,I591722,I591739,I591770,I1160370,I591787,I1160367,I591804,I1160373,I591830,I591838,I591883,I591900,I591917,I591975,I592001,I592009,I592035,I592043,I592060,I592077,I592094,I592111,I591961,I592142,I592159,I592176,I592193,I591958,I591949,I592238,I591952,I591946,I592283,I592300,I592317,I591955,I592348,I592365,I592382,I592408,I592416,I591943,I591967,I592461,I592478,I592495,I591964,I592553,I1263291,I592579,I592587,I1263285,I592613,I592621,I1263294,I592638,I1263273,I592655,I592672,I1263282,I592689,I592539,I592720,I592737,I592754,I1263297,I592771,I1263276,I592536,I592527,I592816,I592530,I592524,I592861,I1263279,I592878,I592895,I592533,I592926,I1263288,I592943,I592960,I592986,I592994,I592521,I592545,I593039,I593056,I593073,I592542,I593131,I593157,I593165,I593191,I593199,I593216,I593233,I593250,I593267,I593117,I593298,I593315,I593332,I593349,I593114,I593105,I593394,I593108,I593102,I593439,I593456,I593473,I593111,I593504,I593521,I593538,I593564,I593572,I593099,I593123,I593617,I593634,I593651,I593120,I593709,I786151,I593735,I593743,I786163,I593769,I593777,I786154,I593794,I786157,I593811,I593828,I786160,I593845,I593876,I593893,I593910,I593927,I786166,I593972,I594017,I786172,I594034,I594051,I594082,I594099,I786169,I594116,I786175,I594142,I594150,I594195,I594212,I594229,I594287,I594313,I594321,I594347,I594355,I594372,I594389,I594406,I594423,I594273,I594454,I594471,I594488,I594505,I594270,I594261,I594550,I594264,I594258,I594595,I594612,I594629,I594267,I594660,I594677,I594694,I594720,I594728,I594255,I594279,I594773,I594790,I594807,I594276,I594865,I594891,I594899,I594925,I594933,I594950,I594967,I594984,I595001,I595032,I595049,I595066,I595083,I595128,I595173,I595190,I595207,I595238,I595255,I595272,I595298,I595306,I595351,I595368,I595385,I595443,I595469,I595477,I595503,I595511,I595528,I595545,I595562,I595579,I595429,I595610,I595627,I595644,I595661,I595426,I595417,I595706,I595420,I595414,I595751,I595768,I595785,I595423,I595816,I595833,I595850,I595876,I595884,I595411,I595435,I595929,I595946,I595963,I595432,I596021,I1201971,I596047,I596055,I1201977,I596081,I596089,I596106,I1201974,I596123,I596140,I1201992,I596157,I596188,I596205,I596222,I1201995,I596239,I596284,I596329,I1201980,I596346,I596363,I596394,I1201986,I596411,I1201983,I596428,I1201989,I596454,I596462,I596507,I596524,I596541,I596599,I700607,I596625,I596633,I700619,I596659,I596667,I700610,I596684,I700613,I596701,I596718,I700616,I596735,I596585,I596766,I596783,I596800,I596817,I700622,I596582,I596573,I596862,I596576,I596570,I596907,I700628,I596924,I596941,I596579,I596972,I596989,I700625,I597006,I700631,I597032,I597040,I596567,I596591,I597085,I597102,I597119,I596588,I597177,I597203,I597211,I597237,I597245,I597262,I597279,I597296,I597313,I597344,I597361,I597378,I597395,I597440,I597485,I597502,I597519,I597550,I597567,I597584,I597610,I597618,I597663,I597680,I597697,I597755,I597781,I597789,I597815,I597823,I597840,I597857,I597874,I597891,I597741,I597922,I597939,I597956,I597973,I597738,I597729,I598018,I597732,I597726,I598063,I598080,I598097,I597735,I598128,I598145,I598162,I598188,I598196,I597723,I597747,I598241,I598258,I598275,I597744,I598333,I780371,I598359,I598367,I780383,I598393,I598401,I780374,I598418,I780377,I598435,I598452,I780380,I598469,I598319,I598500,I598517,I598534,I598551,I780386,I598316,I598307,I598596,I598310,I598304,I598641,I780392,I598658,I598675,I598313,I598706,I598723,I780389,I598740,I780395,I598766,I598774,I598301,I598325,I598819,I598836,I598853,I598322,I598911,I598937,I598945,I598971,I598979,I598996,I599013,I599030,I599047,I598897,I599078,I599095,I599112,I599129,I598894,I598885,I599174,I598888,I598882,I599219,I599236,I599253,I598891,I599284,I599301,I599318,I599344,I599352,I598879,I598903,I599397,I599414,I599431,I598900,I599489,I599515,I599523,I599549,I599557,I599574,I599591,I599608,I599625,I599656,I599673,I599690,I599707,I599752,I599797,I599814,I599831,I599862,I599879,I599896,I599922,I599930,I599975,I599992,I600009,I600067,I1132033,I600093,I600101,I1132039,I600127,I600135,I600152,I1132036,I600169,I600186,I1132054,I600203,I600234,I600251,I600268,I1132057,I600285,I600330,I600375,I1132042,I600392,I600409,I600440,I1132048,I600457,I1132045,I600474,I1132051,I600500,I600508,I600553,I600570,I600587,I600645,I1370798,I600671,I600679,I600705,I600713,I1370822,I600730,I1370804,I600747,I600764,I1370819,I600781,I600631,I600812,I600829,I600846,I1370801,I600863,I1370810,I600628,I600619,I600908,I600622,I600616,I600953,I1370807,I600970,I600987,I600625,I601018,I1370816,I601035,I1370825,I601052,I1370813,I601078,I601086,I600613,I600637,I601131,I601148,I601165,I600634,I601223,I601249,I601257,I601283,I601291,I601308,I601325,I601342,I601359,I601390,I601407,I601424,I601441,I601486,I601531,I601548,I601565,I601596,I601613,I601630,I601656,I601664,I601709,I601726,I601743,I601801,I601827,I601835,I601861,I601869,I601886,I601903,I601920,I601937,I601968,I601985,I602002,I602019,I602064,I602109,I602126,I602143,I602174,I602191,I602208,I602234,I602242,I602287,I602304,I602321,I602379,I602405,I602413,I602439,I602447,I602464,I602481,I602498,I602515,I602365,I602546,I602563,I602580,I602597,I602362,I602353,I602642,I602356,I602350,I602687,I602704,I602721,I602359,I602752,I602769,I602786,I602812,I602820,I602347,I602371,I602865,I602882,I602899,I602368,I602957,I602983,I602991,I603017,I603025,I603042,I603059,I603076,I603093,I602943,I603124,I603141,I603158,I603175,I602940,I602931,I603220,I602934,I602928,I603265,I603282,I603299,I602937,I603330,I603347,I603364,I603390,I603398,I602925,I602949,I603443,I603460,I603477,I602946,I603535,I1140703,I603561,I603569,I1140709,I603595,I603603,I603620,I1140706,I603637,I603654,I1140724,I603671,I603521,I603702,I603719,I603736,I1140727,I603753,I603518,I603509,I603798,I603512,I603506,I603843,I1140712,I603860,I603877,I603515,I603908,I1140718,I603925,I1140715,I603942,I1140721,I603968,I603976,I603503,I603527,I604021,I604038,I604055,I603524,I604113,I604139,I604147,I604173,I604181,I604198,I604215,I604232,I604249,I604099,I604280,I604297,I604314,I604331,I604096,I604087,I604376,I604090,I604084,I604421,I604438,I604455,I604093,I604486,I604503,I604520,I604546,I604554,I604081,I604105,I604599,I604616,I604633,I604102,I604691,I785573,I604717,I604725,I785585,I604751,I604759,I785576,I604776,I785579,I604793,I604810,I785582,I604827,I604858,I604875,I604892,I604909,I785588,I604954,I604999,I785594,I605016,I605033,I605064,I605081,I785591,I605098,I785597,I605124,I605132,I605177,I605194,I605211,I605269,I1087633,I605295,I605303,I1087624,I605329,I605337,I1087618,I605354,I1087630,I605371,I605388,I1087621,I605405,I605255,I605436,I605453,I605470,I1087627,I605487,I1087612,I605252,I605243,I605532,I605246,I605240,I605577,I605594,I605611,I605249,I605642,I1087615,I605659,I605676,I605702,I605710,I605237,I605261,I605755,I605772,I605789,I605258,I605847,I605873,I605881,I605907,I605915,I605932,I605949,I605966,I605983,I606014,I606031,I606048,I606065,I606110,I606155,I606172,I606189,I606220,I606237,I606254,I606280,I606288,I606333,I606350,I606367,I606425,I833723,I606451,I606459,I606485,I606493,I833720,I606510,I833735,I606527,I606544,I833729,I606561,I606411,I606592,I606609,I606626,I833726,I606643,I833717,I606408,I606399,I606688,I606402,I606396,I606733,I833738,I606750,I606767,I606405,I606798,I606815,I606832,I833732,I606858,I606866,I606393,I606417,I606911,I606928,I606945,I606414,I607003,I607029,I607037,I607063,I607071,I607088,I607105,I607122,I607139,I606989,I607170,I607187,I607204,I607221,I606986,I606977,I607266,I606980,I606974,I607311,I607328,I607345,I606983,I607376,I607393,I607410,I607436,I607444,I606971,I606995,I607489,I607506,I607523,I606992,I607581,I607607,I607615,I607641,I607649,I607666,I607683,I607700,I607717,I607567,I607748,I607765,I607782,I607799,I607564,I607555,I607844,I607558,I607552,I607889,I607906,I607923,I607561,I607954,I607971,I607988,I608014,I608022,I607549,I607573,I608067,I608084,I608101,I607570,I608159,I608185,I608193,I608219,I608227,I608244,I608261,I608278,I608295,I608326,I608343,I608360,I608377,I608422,I608467,I608484,I608501,I608532,I608549,I608566,I608592,I608600,I608645,I608662,I608679,I608737,I608763,I608771,I608797,I608805,I608822,I608839,I608856,I608873,I608904,I608921,I608938,I608955,I609000,I609045,I609062,I609079,I609110,I609127,I609144,I609170,I609178,I609223,I609240,I609257,I609315,I609341,I609349,I609375,I609383,I609400,I609417,I609434,I609451,I609301,I609482,I609499,I609516,I609533,I609298,I609289,I609578,I609292,I609286,I609623,I609640,I609657,I609295,I609688,I609705,I609722,I609748,I609756,I609283,I609307,I609801,I609818,I609835,I609304,I609893,I609919,I609927,I609953,I609961,I609978,I609995,I610012,I610029,I610060,I610077,I610094,I610111,I610156,I610201,I610218,I610235,I610266,I610283,I610300,I610326,I610334,I610379,I610396,I610413,I610471,I948473,I610497,I610505,I948470,I610531,I610539,I948467,I610556,I948494,I610573,I610590,I948482,I610607,I610457,I610638,I610655,I610672,I948488,I610689,I948479,I610454,I610445,I610734,I610448,I610442,I610779,I948476,I610796,I610813,I610451,I610844,I948491,I610861,I948485,I610878,I610904,I610912,I610439,I610463,I610957,I610974,I610991,I610460,I611049,I1207751,I611075,I611083,I1207757,I611109,I611117,I611134,I1207754,I611151,I611168,I1207772,I611185,I611216,I611233,I611250,I1207775,I611267,I611312,I611357,I1207760,I611374,I611391,I611422,I1207766,I611439,I1207763,I611456,I1207769,I611482,I611490,I611535,I611552,I611569,I611627,I611653,I611661,I611687,I611695,I611712,I611729,I611746,I611763,I611613,I611794,I611811,I611828,I611845,I611610,I611601,I611890,I611604,I611598,I611935,I611952,I611969,I611607,I612000,I612017,I612034,I612060,I612068,I611595,I611619,I612113,I612130,I612147,I611616,I612205,I612231,I612239,I612265,I612273,I612290,I612307,I612324,I612341,I612191,I612372,I612389,I612406,I612423,I612188,I612179,I612468,I612182,I612176,I612513,I612530,I612547,I612185,I612578,I612595,I612612,I612638,I612646,I612173,I612197,I612691,I612708,I612725,I612194,I612783,I1354733,I612809,I612817,I612843,I612851,I1354757,I612868,I1354739,I612885,I612902,I1354754,I612919,I612950,I612967,I612984,I1354736,I613001,I1354745,I613046,I613091,I1354742,I613108,I613125,I613156,I1354751,I613173,I1354760,I613190,I1354748,I613216,I613224,I613269,I613286,I613303,I613361,I820548,I613387,I613395,I613421,I613429,I820545,I613446,I820560,I613463,I613480,I820554,I613497,I613528,I613545,I613562,I820551,I613579,I820542,I613624,I613669,I820563,I613686,I613703,I613734,I613751,I613768,I820557,I613794,I613802,I613847,I613864,I613881,I613939,I747425,I613965,I613973,I747437,I613999,I614007,I747428,I614024,I747431,I614041,I614058,I747434,I614075,I614106,I614123,I614140,I614157,I747440,I614202,I614247,I747446,I614264,I614281,I614312,I614329,I747443,I614346,I747449,I614372,I614380,I614425,I614442,I614459,I614517,I1182319,I614543,I614551,I1182325,I614577,I614585,I614602,I1182322,I614619,I614636,I1182340,I614653,I614684,I614701,I614718,I1182343,I614735,I614780,I614825,I1182328,I614842,I614859,I614890,I1182334,I614907,I1182331,I614924,I1182337,I614950,I614958,I615003,I615020,I615037,I615095,I1132611,I615121,I615129,I1132617,I615155,I615163,I615180,I1132614,I615197,I615214,I1132632,I615231,I615262,I615279,I615296,I1132635,I615313,I615358,I615403,I1132620,I615420,I615437,I615468,I1132626,I615485,I1132623,I615502,I1132629,I615528,I615536,I615581,I615598,I615615,I615673,I1164401,I615699,I615707,I1164407,I615733,I615741,I615758,I1164404,I615775,I615792,I1164422,I615809,I615659,I615840,I615857,I615874,I1164425,I615891,I615656,I615647,I615936,I615650,I615644,I615981,I1164410,I615998,I616015,I615653,I616046,I1164416,I616063,I1164413,I616080,I1164419,I616106,I616114,I615641,I615665,I616159,I616176,I616193,I615662,I616251,I616277,I616285,I616311,I616319,I616336,I616353,I616370,I616387,I616418,I616435,I616452,I616469,I616514,I616559,I616576,I616593,I616624,I616641,I616658,I616684,I616692,I616737,I616754,I616771,I616829,I817386,I616855,I616863,I616889,I616897,I817383,I616914,I817398,I616931,I616948,I817392,I616965,I616996,I617013,I617030,I817389,I617047,I817380,I617092,I617137,I817401,I617154,I617171,I617202,I617219,I617236,I817395,I617262,I617270,I617315,I617332,I617349,I617407,I841101,I617433,I617441,I617467,I617475,I841098,I617492,I841113,I617509,I617526,I841107,I617543,I617574,I617591,I617608,I841104,I617625,I841095,I617670,I617715,I841116,I617732,I617749,I617780,I617797,I617814,I841110,I617840,I617848,I617893,I617910,I617927,I617985,I1151685,I618011,I618019,I1151691,I618045,I618053,I618070,I1151688,I618087,I618104,I1151706,I618121,I617971,I618152,I618169,I618186,I1151709,I618203,I617968,I617959,I618248,I617962,I617956,I618293,I1151694,I618310,I618327,I617965,I618358,I1151700,I618375,I1151697,I618392,I1151703,I618418,I618426,I617953,I617977,I618471,I618488,I618505,I617974,I618563,I618589,I618597,I618623,I618631,I618648,I618665,I618682,I618699,I618730,I618747,I618764,I618781,I618826,I618871,I618888,I618905,I618936,I618953,I618970,I618996,I619004,I619049,I619066,I619083,I619141,I975605,I619167,I619175,I975602,I619201,I619209,I975599,I619226,I975626,I619243,I619260,I975614,I619277,I619127,I619308,I619325,I619342,I975620,I619359,I975611,I619124,I619115,I619404,I619118,I619112,I619449,I975608,I619466,I619483,I619121,I619514,I975623,I619531,I975617,I619548,I619574,I619582,I619109,I619133,I619627,I619644,I619661,I619130,I619719,I619745,I619753,I619779,I619787,I619804,I619821,I619838,I619855,I619705,I619886,I619903,I619920,I619937,I619702,I619693,I619982,I619696,I619690,I620027,I620044,I620061,I619699,I620092,I620109,I620126,I620152,I620160,I619687,I619711,I620205,I620222,I620239,I619708,I620297,I620323,I620331,I620357,I620365,I620382,I620399,I620416,I620433,I620283,I620464,I620481,I620498,I620515,I620280,I620271,I620560,I620274,I620268,I620605,I620622,I620639,I620277,I620670,I620687,I620704,I620730,I620738,I620265,I620289,I620783,I620800,I620817,I620286,I620875,I620901,I620909,I620935,I620943,I620960,I620977,I620994,I621011,I621042,I621059,I621076,I621093,I621138,I621183,I621200,I621217,I621248,I621265,I621282,I621308,I621316,I621361,I621378,I621395,I621453,I621479,I621487,I621513,I621521,I621538,I621555,I621572,I621589,I621439,I621620,I621637,I621654,I621671,I621436,I621427,I621716,I621430,I621424,I621761,I621778,I621795,I621433,I621826,I621843,I621860,I621886,I621894,I621421,I621445,I621939,I621956,I621973,I621442,I622031,I1088755,I622057,I622065,I1088746,I622091,I622099,I1088740,I622116,I1088752,I622133,I622150,I1088743,I622167,I622017,I622198,I622215,I622232,I1088749,I622249,I1088734,I622014,I622005,I622294,I622008,I622002,I622339,I622356,I622373,I622011,I622404,I1088737,I622421,I622438,I622464,I622472,I621999,I622023,I622517,I622534,I622551,I622020,I622609,I1397573,I622635,I622643,I622669,I622677,I1397597,I622694,I1397579,I622711,I622728,I1397594,I622745,I622595,I622776,I622793,I622810,I1397576,I622827,I1397585,I622592,I622583,I622872,I622586,I622580,I622917,I1397582,I622934,I622951,I622589,I622982,I1397591,I622999,I1397600,I623016,I1397588,I623042,I623050,I622577,I622601,I623095,I623112,I623129,I622598,I623187,I623213,I623221,I623247,I623255,I623272,I623289,I623306,I623323,I623173,I623354,I623371,I623388,I623405,I623170,I623161,I623450,I623164,I623158,I623495,I623512,I623529,I623167,I623560,I623577,I623594,I623620,I623628,I623155,I623179,I623673,I623690,I623707,I623176,I623765,I623791,I623799,I623825,I623833,I623850,I623867,I623884,I623901,I623751,I623932,I623949,I623966,I623983,I623748,I623739,I624028,I623742,I623736,I624073,I624090,I624107,I623745,I624138,I624155,I624172,I624198,I624206,I623733,I623757,I624251,I624268,I624285,I623754,I624343,I1047241,I624369,I624377,I1047232,I624403,I624411,I1047226,I624428,I1047238,I624445,I624462,I1047229,I624479,I624510,I624527,I624544,I1047235,I624561,I1047220,I624606,I624651,I624668,I624685,I624716,I1047223,I624733,I624750,I624776,I624784,I624829,I624846,I624863,I624921,I1297591,I624947,I624955,I1297603,I624981,I624989,I1297594,I625006,I1297582,I625023,I625040,I1297579,I625057,I625088,I625105,I625122,I1297585,I625139,I625184,I625229,I1297600,I625246,I625263,I625294,I1297588,I625311,I625328,I1297597,I625354,I625362,I625407,I625424,I625441,I625499,I1299903,I625525,I625533,I1299915,I625559,I625567,I1299906,I625584,I1299894,I625601,I625618,I1299891,I625635,I625666,I625683,I625700,I1299897,I625717,I625762,I625807,I1299912,I625824,I625841,I625872,I1299900,I625889,I625906,I1299909,I625932,I625940,I625985,I626002,I626019,I626077,I626103,I626111,I626137,I626145,I626162,I626179,I626196,I626213,I626063,I626244,I626261,I626278,I626295,I626060,I626051,I626340,I626054,I626048,I626385,I626402,I626419,I626057,I626450,I626467,I626484,I626510,I626518,I626045,I626069,I626563,I626580,I626597,I626066,I626655,I1000153,I626681,I626689,I1000150,I626715,I626723,I1000147,I626740,I1000174,I626757,I626774,I1000162,I626791,I626641,I626822,I626839,I626856,I1000168,I626873,I1000159,I626638,I626629,I626918,I626632,I626626,I626963,I1000156,I626980,I626997,I626635,I627028,I1000171,I627045,I1000165,I627062,I627088,I627096,I626623,I626647,I627141,I627158,I627175,I626644,I627233,I627259,I627267,I627293,I627301,I627318,I627335,I627352,I627369,I627400,I627417,I627434,I627451,I627496,I627541,I627558,I627575,I627606,I627623,I627640,I627666,I627674,I627719,I627736,I627753,I627811,I1274715,I627837,I627845,I1274709,I627871,I627879,I1274718,I627896,I1274697,I627913,I627930,I1274706,I627947,I627797,I627978,I627995,I628012,I1274721,I628029,I1274700,I627794,I627785,I628074,I627788,I627782,I628119,I1274703,I628136,I628153,I627791,I628184,I1274712,I628201,I628218,I628244,I628252,I627779,I627803,I628297,I628314,I628331,I627800,I628389,I628415,I628423,I628449,I628457,I628474,I628491,I628508,I628525,I628375,I628556,I628573,I628590,I628607,I628372,I628363,I628652,I628366,I628360,I628697,I628714,I628731,I628369,I628762,I628779,I628796,I628822,I628830,I628357,I628381,I628875,I628892,I628909,I628378,I628967,I628993,I629001,I629027,I629035,I629052,I629069,I629086,I629103,I628953,I629134,I629151,I629168,I629185,I628950,I628941,I629230,I628944,I628938,I629275,I629292,I629309,I628947,I629340,I629357,I629374,I629400,I629408,I628935,I628959,I629453,I629470,I629487,I628956,I629545,I1273083,I629571,I629579,I1273077,I629605,I629613,I1273086,I629630,I1273065,I629647,I629664,I1273074,I629681,I629712,I629729,I629746,I1273089,I629763,I1273068,I629808,I629853,I1273071,I629870,I629887,I629918,I1273080,I629935,I629952,I629978,I629986,I630031,I630048,I630065,I630123,I1349378,I630149,I630157,I630183,I630191,I1349402,I630208,I1349384,I630225,I630242,I1349399,I630259,I630109,I630290,I630307,I630324,I1349381,I630341,I1349390,I630106,I630097,I630386,I630100,I630094,I630431,I1349387,I630448,I630465,I630103,I630496,I1349396,I630513,I1349405,I630530,I1349393,I630556,I630564,I630091,I630115,I630609,I630626,I630643,I630112,I630701,I1346403,I630727,I630735,I630761,I630769,I1346427,I630786,I1346409,I630803,I630820,I1346424,I630837,I630687,I630868,I630885,I630902,I1346406,I630919,I1346415,I630684,I630675,I630964,I630678,I630672,I631009,I1346412,I631026,I631043,I630681,I631074,I1346421,I631091,I1346430,I631108,I1346418,I631134,I631142,I630669,I630693,I631187,I631204,I631221,I630690,I631279,I631305,I631313,I631339,I631347,I631364,I631381,I631398,I631415,I631265,I631446,I631463,I631480,I631497,I631262,I631253,I631542,I631256,I631250,I631587,I631604,I631621,I631259,I631652,I631669,I631686,I631712,I631720,I631247,I631271,I631765,I631782,I631799,I631268,I631857,I1389838,I631883,I631891,I631917,I631925,I1389862,I631942,I1389844,I631959,I631976,I1389859,I631993,I631843,I632024,I632041,I632058,I1389841,I632075,I1389850,I631840,I631831,I632120,I631834,I631828,I632165,I1389847,I632182,I632199,I631837,I632230,I1389856,I632247,I1389865,I632264,I1389853,I632290,I632298,I631825,I631849,I632343,I632360,I632377,I631846,I632435,I632461,I632469,I632495,I632503,I632520,I632537,I632554,I632571,I632421,I632602,I632619,I632636,I632653,I632418,I632409,I632698,I632412,I632406,I632743,I632760,I632777,I632415,I632808,I632825,I632842,I632868,I632876,I632403,I632427,I632921,I632938,I632955,I632424,I633013,I1101977,I633039,I633047,I1101983,I633073,I633081,I633098,I1101980,I633115,I633132,I1101998,I633149,I633180,I633197,I633214,I1102001,I633231,I633276,I633321,I1101986,I633338,I633355,I633386,I1101992,I633403,I1101989,I633420,I1101995,I633446,I633454,I633499,I633516,I633533,I633591,I633617,I633625,I633651,I633659,I633676,I633693,I633710,I633727,I633758,I633775,I633792,I633809,I633854,I633899,I633916,I633933,I633964,I633981,I633998,I634024,I634032,I634077,I634094,I634111,I634169,I918757,I634195,I634203,I918754,I634229,I634237,I918751,I634254,I918778,I634271,I634288,I918766,I634305,I634336,I634353,I634370,I918772,I634387,I918763,I634432,I634477,I918760,I634494,I634511,I634542,I918775,I634559,I918769,I634576,I634602,I634610,I634655,I634672,I634689,I634747,I634773,I634781,I634807,I634815,I634832,I634849,I634866,I634883,I634914,I634931,I634948,I634965,I635010,I635055,I635072,I635089,I635120,I635137,I635154,I635180,I635188,I635233,I635250,I635267,I635325,I635351,I635359,I635385,I635393,I635410,I635427,I635444,I635461,I635492,I635509,I635526,I635543,I635588,I635633,I635650,I635667,I635698,I635715,I635732,I635758,I635766,I635811,I635828,I635845,I635903,I732975,I635929,I635937,I732987,I635963,I635971,I732978,I635988,I732981,I636005,I636022,I732984,I636039,I636070,I636087,I636104,I636121,I732990,I636166,I636211,I732996,I636228,I636245,I636276,I636293,I732993,I636310,I732999,I636336,I636344,I636389,I636406,I636423,I636481,I636507,I636515,I636541,I636549,I636566,I636583,I636600,I636617,I636467,I636648,I636665,I636682,I636699,I636464,I636455,I636744,I636458,I636452,I636789,I636806,I636823,I636461,I636854,I636871,I636888,I636914,I636922,I636449,I636473,I636967,I636984,I637001,I636470,I637059,I1035037,I637085,I637093,I1035034,I637119,I637127,I1035031,I637144,I1035058,I637161,I637178,I1035046,I637195,I637226,I637243,I637260,I1035052,I637277,I1035043,I637322,I637367,I1035040,I637384,I637401,I637432,I1035055,I637449,I1035049,I637466,I637492,I637500,I637545,I637562,I637579,I637637,I637663,I637671,I637697,I637705,I637722,I637739,I637756,I637773,I637804,I637821,I637838,I637855,I637900,I637945,I637962,I637979,I638010,I638027,I638044,I638070,I638078,I638123,I638140,I638157,I638215,I979481,I638241,I638249,I979478,I638275,I638283,I979475,I638300,I979502,I638317,I638334,I979490,I638351,I638201,I638382,I638399,I638416,I979496,I638433,I979487,I638198,I638189,I638478,I638192,I638186,I638523,I979484,I638540,I638557,I638195,I638588,I979499,I638605,I979493,I638622,I638648,I638656,I638183,I638207,I638701,I638718,I638735,I638204,I638793,I723149,I638819,I638827,I723161,I638853,I638861,I723152,I638878,I723155,I638895,I638912,I723158,I638929,I638960,I638977,I638994,I639011,I723164,I639056,I639101,I723170,I639118,I639135,I639166,I639183,I723167,I639200,I723173,I639226,I639234,I639279,I639296,I639313,I639371,I1245339,I639397,I639405,I1245333,I639431,I639439,I1245342,I639456,I1245321,I639473,I639490,I1245330,I639507,I639357,I639538,I639555,I639572,I1245345,I639589,I1245324,I639354,I639345,I639634,I639348,I639342,I639679,I1245327,I639696,I639713,I639351,I639744,I1245336,I639761,I639778,I639804,I639812,I639339,I639363,I639857,I639874,I639891,I639360,I639949,I727195,I639975,I639983,I727207,I640009,I640017,I727198,I640034,I727201,I640051,I640068,I727204,I640085,I640116,I640133,I640150,I640167,I727210,I640212,I640257,I727216,I640274,I640291,I640322,I640339,I727213,I640356,I727219,I640382,I640390,I640435,I640452,I640469,I640527,I640553,I640561,I640587,I640595,I640612,I640629,I640646,I640663,I640513,I640694,I640711,I640728,I640745,I640510,I640501,I640790,I640504,I640498,I640835,I640852,I640869,I640507,I640900,I640917,I640934,I640960,I640968,I640495,I640519,I641013,I641030,I641047,I640516,I641105,I806381,I641131,I641139,I806393,I641165,I641173,I806384,I641190,I806387,I641207,I641224,I806390,I641241,I641272,I641289,I641306,I641323,I806396,I641368,I641413,I806402,I641430,I641447,I641478,I641495,I806399,I641512,I806405,I641538,I641546,I641591,I641608,I641625,I641683,I641709,I641717,I641743,I641751,I641768,I641785,I641802,I641819,I641669,I641850,I641867,I641884,I641901,I641666,I641657,I641946,I641660,I641654,I641991,I642008,I642025,I641663,I642056,I642073,I642090,I642116,I642124,I641651,I641675,I642169,I642186,I642203,I641672,I642261,I1295279,I642287,I642295,I1295291,I642321,I642329,I1295282,I642346,I1295270,I642363,I642380,I1295267,I642397,I642247,I642428,I642445,I642462,I1295273,I642479,I642244,I642235,I642524,I642238,I642232,I642569,I1295288,I642586,I642603,I642241,I642634,I1295276,I642651,I642668,I1295285,I642694,I642702,I642229,I642253,I642747,I642764,I642781,I642250,I642839,I662459,I642865,I642873,I662471,I642899,I642907,I662462,I642924,I662465,I642941,I642958,I662468,I642975,I643006,I643023,I643040,I643057,I662474,I643102,I643147,I662480,I643164,I643181,I643212,I643229,I662477,I643246,I662483,I643272,I643280,I643325,I643342,I643359,I643417,I643443,I643451,I643477,I643485,I643502,I643519,I643536,I643553,I643584,I643601,I643618,I643635,I643680,I643725,I643742,I643759,I643790,I643807,I643824,I643850,I643858,I643903,I643920,I643937,I643995,I741645,I644021,I644029,I741657,I644055,I644063,I741648,I644080,I741651,I644097,I644114,I741654,I644131,I643981,I644162,I644179,I644196,I644213,I741660,I643978,I643969,I644258,I643972,I643966,I644303,I741666,I644320,I644337,I643975,I644368,I644385,I741663,I644402,I741669,I644428,I644436,I643963,I643987,I644481,I644498,I644515,I643984,I644573,I1145905,I644599,I644607,I1145911,I644633,I644641,I644658,I1145908,I644675,I644692,I1145926,I644709,I644740,I644757,I644774,I1145929,I644791,I644836,I644881,I1145914,I644898,I644915,I644946,I1145920,I644963,I1145917,I644980,I1145923,I645006,I645014,I645059,I645076,I645093,I645151,I645177,I645185,I645211,I645219,I645236,I645253,I645270,I645287,I645318,I645335,I645352,I645369,I645414,I645459,I645476,I645493,I645524,I645541,I645558,I645584,I645592,I645637,I645654,I645671,I645729,I645755,I645763,I645789,I645797,I645814,I645831,I645848,I645865,I645715,I645896,I645913,I645930,I645947,I645712,I645703,I645992,I645706,I645700,I646037,I646054,I646071,I645709,I646102,I646119,I646136,I646162,I646170,I645697,I645721,I646215,I646232,I646249,I645718,I646307,I646333,I646341,I646367,I646375,I646392,I646409,I646426,I646443,I646293,I646474,I646491,I646508,I646525,I646290,I646281,I646570,I646284,I646278,I646615,I646632,I646649,I646287,I646680,I646697,I646714,I646740,I646748,I646275,I646299,I646793,I646810,I646827,I646296,I646885,I1400548,I646911,I646919,I646945,I646953,I1400572,I646970,I1400554,I646987,I647004,I1400569,I647021,I647052,I647069,I647086,I1400551,I647103,I1400560,I647148,I647193,I1400557,I647210,I647227,I647258,I1400566,I647275,I1400575,I647292,I1400563,I647318,I647326,I647371,I647388,I647405,I647463,I977543,I647489,I647497,I977540,I647523,I647531,I977537,I647548,I977564,I647565,I647582,I977552,I647599,I647630,I647647,I647664,I977558,I647681,I977549,I647726,I647771,I977546,I647788,I647805,I647836,I977561,I647853,I977555,I647870,I647896,I647904,I647949,I647966,I647983,I648041,I648067,I648075,I648101,I648109,I648126,I648143,I648160,I648177,I648027,I648208,I648225,I648242,I648259,I648024,I648015,I648304,I648018,I648012,I648349,I648366,I648383,I648021,I648414,I648431,I648448,I648474,I648482,I648009,I648033,I648527,I648544,I648561,I648030,I648619,I648645,I648653,I648679,I648687,I648704,I648721,I648738,I648755,I648605,I648786,I648803,I648820,I648837,I648602,I648593,I648882,I648596,I648590,I648927,I648944,I648961,I648599,I648992,I649009,I649026,I649052,I649060,I648587,I648611,I649105,I649122,I649139,I648608,I649197,I649223,I649231,I649257,I649265,I649282,I649299,I649316,I649333,I649364,I649381,I649398,I649415,I649460,I649505,I649522,I649539,I649570,I649587,I649604,I649630,I649638,I649683,I649700,I649717,I649775,I886423,I649801,I649809,I649835,I649843,I886420,I649860,I886435,I649877,I649894,I886429,I649911,I649942,I649959,I649976,I886426,I649993,I886417,I650038,I650083,I886438,I650100,I650117,I650148,I650165,I650182,I886432,I650208,I650216,I650261,I650278,I650295,I650353,I650379,I650387,I650413,I650421,I650438,I650455,I650472,I650489,I650520,I650537,I650554,I650571,I650616,I650661,I650678,I650695,I650726,I650743,I650760,I650786,I650794,I650839,I650856,I650873,I650931,I650957,I650965,I650991,I650999,I651016,I651033,I651050,I651067,I651098,I651115,I651132,I651149,I651194,I651239,I651256,I651273,I651304,I651321,I651338,I651364,I651372,I651417,I651434,I651451,I651509,I651535,I651543,I651569,I651577,I651594,I651611,I651628,I651645,I651495,I651676,I651693,I651710,I651727,I651492,I651483,I651772,I651486,I651480,I651817,I651834,I651851,I651489,I651882,I651899,I651916,I651942,I651950,I651477,I651501,I651995,I652012,I652029,I651498,I652087,I652113,I652121,I652147,I652155,I652172,I652189,I652206,I652223,I652073,I652254,I652271,I652288,I652305,I652070,I652061,I652350,I652064,I652058,I652395,I652412,I652429,I652067,I652460,I652477,I652494,I652520,I652528,I652055,I652079,I652573,I652590,I652607,I652076,I652665,I652691,I652699,I652725,I652733,I652750,I652767,I652784,I652801,I652832,I652849,I652866,I652883,I652928,I652973,I652990,I653007,I653038,I653055,I653072,I653098,I653106,I653151,I653168,I653185,I653243,I722571,I653269,I653277,I722583,I653303,I653311,I722574,I653328,I722577,I653345,I653362,I722580,I653379,I653229,I653410,I653427,I653444,I653461,I722586,I653226,I653217,I653506,I653220,I653214,I653551,I722592,I653568,I653585,I653223,I653616,I653633,I722589,I653650,I722595,I653676,I653684,I653211,I653235,I653729,I653746,I653763,I653232,I653821,I653847,I653855,I653881,I653889,I653906,I653923,I653940,I653957,I653988,I654005,I654022,I654039,I654084,I654129,I654146,I654163,I654194,I654211,I654228,I654254,I654262,I654307,I654324,I654341,I654399,I654425,I654433,I654459,I654467,I654484,I654501,I654518,I654535,I654385,I654566,I654583,I654600,I654617,I654382,I654373,I654662,I654376,I654370,I654707,I654724,I654741,I654379,I654772,I654789,I654806,I654832,I654840,I654367,I654391,I654885,I654902,I654919,I654388,I654977,I856911,I655003,I655011,I655037,I655045,I856908,I655062,I856923,I655079,I655096,I856917,I655113,I655144,I655161,I655178,I856914,I655195,I856905,I655240,I655285,I856926,I655302,I655319,I655350,I655367,I655384,I856920,I655410,I655418,I655463,I655480,I655497,I655555,I655581,I655589,I655615,I655623,I655640,I655657,I655674,I655691,I655722,I655739,I655756,I655773,I655818,I655863,I655880,I655897,I655928,I655945,I655962,I655988,I655996,I656041,I656058,I656075,I656133,I656159,I656167,I656193,I656201,I656218,I656235,I656252,I656269,I656119,I656300,I656317,I656334,I656351,I656116,I656107,I656396,I656110,I656104,I656441,I656458,I656475,I656113,I656506,I656523,I656540,I656566,I656574,I656101,I656125,I656619,I656636,I656653,I656122,I656711,I656737,I656745,I656771,I656779,I656796,I656813,I656830,I656847,I656878,I656895,I656912,I656929,I656974,I657019,I657036,I657053,I657084,I657101,I657118,I657144,I657152,I657197,I657214,I657231,I657289,I745691,I657315,I657323,I745703,I657349,I657357,I745694,I657374,I745697,I657391,I657408,I745700,I657425,I657275,I657456,I657473,I657490,I657507,I745706,I657272,I657263,I657552,I657266,I657260,I657597,I745712,I657614,I657631,I657269,I657662,I657679,I745709,I657696,I745715,I657722,I657730,I657257,I657281,I657775,I657792,I657809,I657278,I657867,I657893,I657901,I657927,I657935,I657952,I657969,I657986,I658003,I657853,I658034,I658051,I658068,I658085,I657850,I657841,I658130,I657844,I657838,I658175,I658192,I658209,I657847,I658240,I658257,I658274,I658300,I658308,I657835,I657859,I658353,I658370,I658387,I657856,I658445,I1247497,I658471,I658479,I658496,I1247500,I1247509,I658513,I1247512,I658539,I658547,I1247521,I1247503,I658573,I658581,I658598,I658615,I658632,I658428,I658672,I658680,I658697,I658714,I658731,I658431,I658762,I1247518,I658779,I1247515,I658805,I658813,I658413,I658844,I658422,I658875,I658892,I658434,I658923,I1247506,I658425,I658416,I658419,I658437,I659023,I659049,I659057,I659074,I659091,I659117,I659125,I659151,I659159,I659176,I659193,I659210,I659250,I659258,I659275,I659292,I659309,I659340,I659357,I659383,I659391,I659422,I659453,I659470,I659501,I659601,I831097,I659627,I659635,I659652,I831085,I831103,I659669,I831100,I659695,I659703,I831091,I831088,I659729,I659737,I659754,I659771,I659788,I831082,I659828,I659836,I659853,I659870,I659887,I659918,I659935,I659961,I659969,I660000,I660031,I660048,I660079,I831094,I660179,I660205,I660213,I660230,I660247,I660273,I660281,I660307,I660315,I660332,I660349,I660366,I660406,I660414,I660431,I660448,I660465,I660496,I660513,I660539,I660547,I660578,I660609,I660626,I660657,I660757,I1098527,I660783,I660791,I660808,I1098509,I1098521,I660825,I1098524,I660851,I660859,I1098518,I1098515,I660885,I660893,I660910,I660927,I660944,I1098533,I660984,I660992,I661009,I661026,I661043,I661074,I1098512,I661091,I661117,I661125,I661156,I661187,I661204,I661235,I1098530,I661335,I1119335,I661361,I661369,I661386,I1119317,I1119329,I661403,I1119332,I661429,I661437,I1119326,I1119323,I661463,I661471,I661488,I661505,I661522,I1119341,I661562,I661570,I661587,I661604,I661621,I661652,I1119320,I661669,I661695,I661703,I661734,I661765,I661782,I661813,I1119338,I661913,I1090435,I661939,I661947,I661964,I1090417,I1090429,I661981,I1090432,I662007,I662015,I1090426,I1090423,I662041,I662049,I662066,I662083,I662100,I1090441,I662140,I662148,I662165,I662182,I662199,I662230,I1090420,I662247,I662273,I662281,I662312,I662343,I662360,I662391,I1090438,I662491,I1081447,I662517,I662525,I662542,I1081444,I1081462,I662559,I1081459,I662585,I662593,I1081441,I662619,I662627,I662644,I662661,I662678,I1081453,I662718,I662726,I662743,I662760,I662777,I662808,I1081456,I662825,I662851,I662859,I662890,I662921,I662938,I662969,I1081450,I663069,I1074715,I663095,I663103,I663120,I1074712,I1074730,I663137,I1074727,I663163,I663171,I1074709,I663197,I663205,I663222,I663239,I663256,I663052,I1074721,I663296,I663304,I663321,I663338,I663355,I663055,I663386,I1074724,I663403,I663429,I663437,I663037,I663468,I663046,I663499,I663516,I663058,I663547,I1074718,I663049,I663040,I663043,I663061,I663647,I859555,I663673,I663681,I663698,I859543,I859561,I663715,I859558,I663741,I663749,I859549,I859546,I663775,I663783,I663800,I663817,I663834,I859540,I663874,I663882,I663899,I663916,I663933,I663964,I663981,I664007,I664015,I664046,I664077,I664094,I664125,I859552,I664225,I1042161,I664251,I664259,I664276,I1042137,I1042152,I664293,I1042164,I664319,I664327,I1042149,I1042140,I664353,I664361,I664378,I664395,I664412,I664208,I664452,I664460,I664477,I664494,I664511,I664211,I664542,I1042155,I1042146,I664559,I1042158,I664585,I664593,I664193,I664624,I664202,I664655,I664672,I664214,I664703,I1042143,I664205,I664196,I664199,I664217,I664803,I908039,I664829,I664837,I664854,I908027,I908045,I664871,I908042,I664897,I664905,I908033,I908030,I664931,I664939,I664956,I664973,I664990,I908024,I665030,I665038,I665055,I665072,I665089,I665120,I665137,I665163,I665171,I665202,I665233,I665250,I665281,I908036,I665381,I665407,I665415,I665432,I665449,I665475,I665483,I665509,I665517,I665534,I665551,I665568,I665364,I665608,I665616,I665633,I665650,I665667,I665367,I665698,I665715,I665741,I665749,I665349,I665780,I665358,I665811,I665828,I665370,I665859,I665361,I665352,I665355,I665373,I665959,I1157483,I665985,I665993,I666010,I1157465,I1157477,I666027,I1157480,I666053,I666061,I1157474,I1157471,I666087,I666095,I666112,I666129,I666146,I665942,I1157489,I666186,I666194,I666211,I666228,I666245,I665945,I666276,I1157468,I666293,I666319,I666327,I665927,I666358,I665936,I666389,I666406,I665948,I666437,I1157486,I665939,I665930,I665933,I665951,I666537,I666563,I666571,I666588,I666605,I666631,I666639,I666665,I666673,I666690,I666707,I666724,I666520,I666764,I666772,I666789,I666806,I666823,I666523,I666854,I666871,I666897,I666905,I666505,I666936,I666514,I666967,I666984,I666526,I667015,I666517,I666508,I666511,I666529,I667115,I1166731,I667141,I667149,I667166,I1166713,I1166725,I667183,I1166728,I667209,I667217,I1166722,I1166719,I667243,I667251,I667268,I667285,I667302,I667098,I1166737,I667342,I667350,I667367,I667384,I667401,I667101,I667432,I1166716,I667449,I667475,I667483,I667083,I667514,I667092,I667545,I667562,I667104,I667593,I1166734,I667095,I667086,I667089,I667107,I667693,I667719,I667727,I667744,I667761,I667787,I667795,I667821,I667829,I667846,I667863,I667880,I667920,I667928,I667945,I667962,I667979,I668010,I668027,I668053,I668061,I668092,I668123,I668140,I668171,I668271,I1223953,I668297,I668305,I668322,I1223935,I1223947,I668339,I1223950,I668365,I668373,I1223944,I1223941,I668399,I668407,I668424,I668441,I668458,I1223959,I668498,I668506,I668523,I668540,I668557,I668588,I1223938,I668605,I668631,I668639,I668670,I668701,I668718,I668749,I1223956,I668849,I1178291,I668875,I668883,I668900,I1178273,I1178285,I668917,I1178288,I668943,I668951,I1178282,I1178279,I668977,I668985,I669002,I669019,I669036,I668832,I1178297,I669076,I669084,I669101,I669118,I669135,I668835,I669166,I1178276,I669183,I669209,I669217,I668817,I669248,I668826,I669279,I669296,I668838,I669327,I1178294,I668829,I668820,I668823,I668841,I669427,I1029887,I669453,I669461,I669478,I1029863,I1029878,I669495,I1029890,I669521,I669529,I1029875,I1029866,I669555,I669563,I669580,I669597,I669614,I669410,I669654,I669662,I669679,I669696,I669713,I669413,I669744,I1029881,I1029872,I669761,I1029884,I669787,I669795,I669395,I669826,I669404,I669857,I669874,I669416,I669905,I1029869,I669407,I669398,I669401,I669419,I670005,I670031,I670039,I670056,I670073,I670099,I670107,I670133,I670141,I670158,I670175,I670192,I670232,I670240,I670257,I670274,I670291,I670322,I670339,I670365,I670373,I670404,I670435,I670452,I670483,I670583,I1252937,I670609,I670617,I670634,I1252940,I1252949,I670651,I1252952,I670677,I670685,I1252961,I1252943,I670711,I670719,I670736,I670753,I670770,I670566,I670810,I670818,I670835,I670852,I670869,I670569,I670900,I1252958,I670917,I1252955,I670943,I670951,I670551,I670982,I670560,I671013,I671030,I670572,I671061,I1252946,I670563,I670554,I670557,I670575,I671161,I1169043,I671187,I671195,I671212,I1169025,I1169037,I671229,I1169040,I671255,I671263,I1169034,I1169031,I671289,I671297,I671314,I671331,I671348,I1169049,I671388,I671396,I671413,I671430,I671447,I671478,I1169028,I671495,I671521,I671529,I671560,I671591,I671608,I671639,I1169046,I671739,I1364875,I671765,I671773,I671790,I1364860,I1364848,I671807,I1364863,I671833,I671841,I1364866,I671867,I671875,I671892,I671909,I671926,I1364854,I671966,I671974,I671991,I672008,I672025,I672056,I1364851,I1364857,I672073,I1364872,I672099,I672107,I672138,I672169,I672186,I672217,I1364869,I672317,I672343,I672351,I672368,I672385,I672411,I672419,I672445,I672453,I672470,I672487,I672504,I672544,I672552,I672569,I672586,I672603,I672634,I672651,I672677,I672685,I672716,I672747,I672764,I672795,I672895,I930403,I672921,I672929,I672946,I930379,I930394,I672963,I930406,I672989,I672997,I930391,I930382,I673023,I673031,I673048,I673065,I673082,I672878,I673122,I673130,I673147,I673164,I673181,I672881,I673212,I930397,I930388,I673229,I930400,I673255,I673263,I672863,I673294,I672872,I673325,I673342,I672884,I673373,I930385,I672875,I672866,I672869,I672887,I673473,I1141877,I673499,I673507,I673524,I1141859,I1141871,I673541,I1141874,I673567,I673575,I1141868,I1141865,I673601,I673609,I673626,I673643,I673660,I1141883,I673700,I673708,I673725,I673742,I673759,I673790,I1141862,I673807,I673833,I673841,I673872,I673903,I673920,I673951,I1141880,I674051,I674077,I674085,I674102,I674119,I674145,I674153,I674179,I674187,I674204,I674221,I674238,I674034,I674278,I674286,I674303,I674320,I674337,I674037,I674368,I674385,I674411,I674419,I674019,I674450,I674028,I674481,I674498,I674040,I674529,I674031,I674022,I674025,I674043,I674629,I863771,I674655,I674663,I674680,I863759,I863777,I674697,I863774,I674723,I674731,I863765,I863762,I674757,I674765,I674782,I674799,I674816,I674612,I863756,I674856,I674864,I674881,I674898,I674915,I674615,I674946,I674963,I674989,I674997,I674597,I675028,I674606,I675059,I675076,I674618,I675107,I863768,I674609,I674600,I674603,I674621,I675207,I675233,I675241,I675258,I675275,I675301,I675309,I675335,I675343,I675360,I675377,I675394,I675190,I675434,I675442,I675459,I675476,I675493,I675193,I675524,I675541,I675567,I675575,I675175,I675606,I675184,I675637,I675654,I675196,I675685,I675187,I675178,I675181,I675199,I675785,I1291221,I675811,I675819,I675836,I1291245,I1291227,I675853,I1291233,I675879,I675887,I1291239,I1291224,I675913,I675921,I675938,I675955,I675972,I1291236,I676012,I676020,I676037,I676054,I676071,I676102,I1291242,I1291230,I676119,I676145,I676153,I676184,I676215,I676232,I676263,I676363,I821611,I676389,I676397,I676414,I821599,I821617,I676431,I821614,I676457,I676465,I821605,I821602,I676491,I676499,I676516,I676533,I676550,I821596,I676590,I676598,I676615,I676632,I676649,I676680,I676697,I676723,I676731,I676762,I676793,I676810,I676841,I821608,I676941,I825827,I676967,I676975,I676992,I825815,I825833,I677009,I825830,I677035,I677043,I825821,I825818,I677069,I677077,I677094,I677111,I677128,I676924,I825812,I677168,I677176,I677193,I677210,I677227,I676927,I677258,I677275,I677301,I677309,I676909,I677340,I676918,I677371,I677388,I676930,I677419,I825824,I676921,I676912,I676915,I676933,I677519,I677545,I677553,I677570,I677587,I677613,I677621,I677647,I677655,I677672,I677689,I677706,I677502,I677746,I677754,I677771,I677788,I677805,I677505,I677836,I677853,I677879,I677887,I677487,I677918,I677496,I677949,I677966,I677508,I677997,I677499,I677490,I677493,I677511,I678097,I678123,I678131,I678148,I678165,I678191,I678199,I678225,I678233,I678250,I678267,I678284,I678080,I678324,I678332,I678349,I678366,I678383,I678083,I678414,I678431,I678457,I678465,I678065,I678496,I678074,I678527,I678544,I678086,I678575,I678077,I678068,I678071,I678089,I678675,I678701,I678709,I678726,I678743,I678769,I678777,I678803,I678811,I678828,I678845,I678862,I678902,I678910,I678927,I678944,I678961,I678992,I679009,I679035,I679043,I679074,I679105,I679122,I679153,I679253,I679279,I679287,I679304,I679321,I679347,I679355,I679381,I679389,I679406,I679423,I679440,I679480,I679488,I679505,I679522,I679539,I679570,I679587,I679613,I679621,I679652,I679683,I679700,I679731,I679831,I1251849,I679857,I679865,I679882,I1251852,I1251861,I679899,I1251864,I679925,I679933,I1251873,I1251855,I679959,I679967,I679984,I680001,I680018,I680058,I680066,I680083,I680100,I680117,I680148,I1251870,I680165,I1251867,I680191,I680199,I680230,I680261,I680278,I680309,I1251858,I680409,I680435,I680443,I680460,I680477,I680503,I680511,I680537,I680545,I680562,I680579,I680596,I680636,I680644,I680661,I680678,I680695,I680726,I680743,I680769,I680777,I680808,I680839,I680856,I680887,I680987,I958827,I681013,I681021,I681038,I958803,I958818,I681055,I958830,I681081,I681089,I958815,I958806,I681115,I681123,I681140,I681157,I681174,I680970,I681214,I681222,I681239,I681256,I681273,I680973,I681304,I958821,I958812,I681321,I958824,I681347,I681355,I680955,I681386,I680964,I681417,I681434,I680976,I681465,I958809,I680967,I680958,I680961,I680979,I681565,I1344645,I681591,I681599,I681616,I1344630,I1344618,I681633,I1344633,I681659,I681667,I1344636,I681693,I681701,I681718,I681735,I681752,I1344624,I681792,I681800,I681817,I681834,I681851,I681882,I1344621,I1344627,I681899,I1344642,I681925,I681933,I681964,I681995,I682012,I682043,I1344639,I682143,I682169,I682177,I682194,I682211,I682237,I682245,I682271,I682279,I682296,I682313,I682330,I682370,I682378,I682395,I682412,I682429,I682460,I682477,I682503,I682511,I682542,I682573,I682590,I682621,I682721,I682747,I682755,I682772,I682789,I682815,I682823,I682849,I682857,I682874,I682891,I682908,I682704,I682948,I682956,I682973,I682990,I683007,I682707,I683038,I683055,I683081,I683089,I682689,I683120,I682698,I683151,I683168,I682710,I683199,I682701,I682692,I682695,I682713,I683299,I683325,I683333,I683350,I683367,I683393,I683401,I683427,I683435,I683452,I683469,I683486,I683282,I683526,I683534,I683551,I683568,I683585,I683285,I683616,I683633,I683659,I683667,I683267,I683698,I683276,I683729,I683746,I683288,I683777,I683279,I683270,I683273,I683291,I683877,I1275241,I683903,I683911,I683928,I1275244,I1275253,I683945,I1275256,I683971,I683979,I1275265,I1275247,I684005,I684013,I684030,I684047,I684064,I683860,I684104,I684112,I684129,I684146,I684163,I683863,I684194,I1275262,I684211,I1275259,I684237,I684245,I683845,I684276,I683854,I684307,I684324,I683866,I684355,I1275250,I683857,I683848,I683851,I683869,I684455,I1128005,I684481,I684489,I684506,I1127987,I1127999,I684523,I1128002,I684549,I684557,I1127996,I1127993,I684583,I684591,I684608,I684625,I684642,I1128011,I684682,I684690,I684707,I684724,I684741,I684772,I1127990,I684789,I684815,I684823,I684854,I684885,I684902,I684933,I1128008,I685033,I685059,I685067,I685084,I685101,I685127,I685135,I685161,I685169,I685186,I685203,I685220,I685260,I685268,I685285,I685302,I685319,I685350,I685367,I685393,I685401,I685432,I685463,I685480,I685511,I685611,I1334530,I685637,I685645,I685662,I1334515,I1334503,I685679,I1334518,I685705,I685713,I1334521,I685739,I685747,I685764,I685781,I685798,I1334509,I685838,I685846,I685863,I685880,I685897,I685928,I1334506,I1334512,I685945,I1334527,I685971,I685979,I686010,I686041,I686058,I686089,I1334524,I686189,I847961,I686215,I686223,I686240,I847949,I847967,I686257,I847964,I686283,I686291,I847955,I847952,I686317,I686325,I686342,I686359,I686376,I847946,I686416,I686424,I686441,I686458,I686475,I686506,I686523,I686549,I686557,I686588,I686619,I686636,I686667,I847958,I686767,I872730,I686793,I686801,I686818,I872718,I872736,I686835,I872733,I686861,I686869,I872724,I872721,I686895,I686903,I686920,I686937,I686954,I686750,I872715,I686994,I687002,I687019,I687036,I687053,I686753,I687084,I687101,I687127,I687135,I686735,I687166,I686744,I687197,I687214,I686756,I687245,I872727,I686747,I686738,I686741,I686759,I687345,I1268169,I687371,I687379,I687396,I1268172,I1268181,I687413,I1268184,I687439,I687447,I1268193,I1268175,I687473,I687481,I687498,I687515,I687532,I687328,I687572,I687580,I687597,I687614,I687631,I687331,I687662,I1268190,I687679,I1268187,I687705,I687713,I687313,I687744,I687322,I687775,I687792,I687334,I687823,I1268178,I687325,I687316,I687319,I687337,I687923,I1011799,I687949,I687957,I687974,I1011775,I1011790,I687991,I1011802,I688017,I688025,I1011787,I1011778,I688051,I688059,I688076,I688093,I688110,I687906,I688150,I688158,I688175,I688192,I688209,I687909,I688240,I1011793,I1011784,I688257,I1011796,I688283,I688291,I687891,I688322,I687900,I688353,I688370,I687912,I688401,I1011781,I687903,I687894,I687897,I687915,I688501,I688527,I688535,I688552,I688569,I688595,I688603,I688629,I688637,I688654,I688671,I688688,I688728,I688736,I688753,I688770,I688787,I688818,I688835,I688861,I688869,I688900,I688931,I688948,I688979,I689079,I982083,I689105,I689113,I689130,I982059,I982074,I689147,I982086,I689173,I689181,I982071,I982062,I689207,I689215,I689232,I689249,I689266,I689306,I689314,I689331,I689348,I689365,I689396,I982077,I982068,I689413,I982080,I689439,I689447,I689478,I689509,I689526,I689557,I982065,I689657,I1043453,I689683,I689691,I689708,I1043429,I1043444,I689725,I1043456,I689751,I689759,I1043441,I1043432,I689785,I689793,I689810,I689827,I689844,I689640,I689884,I689892,I689909,I689926,I689943,I689643,I689974,I1043447,I1043438,I689991,I1043450,I690017,I690025,I689625,I690056,I689634,I690087,I690104,I689646,I690135,I1043435,I689637,I689628,I689631,I689649,I690235,I925235,I690261,I690269,I690286,I925211,I925226,I690303,I925238,I690329,I690337,I925223,I925214,I690363,I690371,I690388,I690405,I690422,I690462,I690470,I690487,I690504,I690521,I690552,I925229,I925220,I690569,I925232,I690595,I690603,I690634,I690665,I690682,I690713,I925217,I690813,I690839,I690847,I690864,I690881,I690907,I690915,I690941,I690949,I690966,I690983,I691000,I691040,I691048,I691065,I691082,I691099,I691130,I691147,I691173,I691181,I691212,I691243,I691260,I691291,I691391,I691417,I691425,I691442,I691459,I691485,I691493,I691519,I691527,I691544,I691561,I691578,I691374,I691618,I691626,I691643,I691660,I691677,I691377,I691708,I691725,I691751,I691759,I691359,I691790,I691368,I691821,I691838,I691380,I691869,I691371,I691362,I691365,I691383,I691969,I691995,I692003,I692020,I692037,I692063,I692071,I692097,I692105,I692122,I692139,I692156,I692196,I692204,I692221,I692238,I692255,I692286,I692303,I692329,I692337,I692368,I692399,I692416,I692447,I692547,I1270889,I692573,I692581,I692598,I1270892,I1270901,I692615,I1270904,I692641,I692649,I1270913,I1270895,I692675,I692683,I692700,I692717,I692734,I692774,I692782,I692799,I692816,I692833,I692864,I1270910,I692881,I1270907,I692907,I692915,I692946,I692977,I692994,I693025,I1270898,I693125,I918129,I693151,I693159,I693176,I918105,I918120,I693193,I918132,I693219,I693227,I918117,I918108,I693253,I693261,I693278,I693295,I693312,I693108,I693352,I693360,I693377,I693394,I693411,I693111,I693442,I918123,I918114,I693459,I918126,I693485,I693493,I693093,I693524,I693102,I693555,I693572,I693114,I693603,I918111,I693105,I693096,I693099,I693117,I693703,I812125,I693729,I693737,I693754,I812113,I812131,I693771,I812128,I693797,I693805,I812119,I812116,I693831,I693839,I693856,I693873,I693890,I693686,I812110,I693930,I693938,I693955,I693972,I693989,I693689,I694020,I694037,I694063,I694071,I693671,I694102,I693680,I694133,I694150,I693692,I694181,I812122,I693683,I693674,I693677,I693695,I694281,I694307,I694315,I694332,I694349,I694375,I694383,I694409,I694417,I694434,I694451,I694468,I694508,I694516,I694533,I694550,I694567,I694598,I694615,I694641,I694649,I694680,I694711,I694728,I694759,I694859,I913309,I694885,I694893,I694910,I913297,I913315,I694927,I913312,I694953,I694961,I913303,I913300,I694987,I694995,I695012,I695029,I695046,I694842,I913294,I695086,I695094,I695111,I695128,I695145,I694845,I695176,I695193,I695219,I695227,I694827,I695258,I694836,I695289,I695306,I694848,I695337,I913306,I694839,I694830,I694833,I694851,I695437,I1065178,I695463,I695471,I695488,I1065175,I1065193,I695505,I1065190,I695531,I695539,I1065172,I695565,I695573,I695590,I695607,I695624,I1065184,I695664,I695672,I695689,I695706,I695723,I695754,I1065187,I695771,I695797,I695805,I695836,I695867,I695884,I695915,I1065181,I696015,I696041,I696049,I696066,I696083,I696109,I696117,I696143,I696151,I696168,I696185,I696202,I696242,I696250,I696267,I696284,I696301,I696332,I696349,I696375,I696383,I696414,I696445,I696462,I696493,I696593,I1049470,I696619,I696627,I696644,I1049467,I1049485,I696661,I1049482,I696687,I696695,I1049464,I696721,I696729,I696746,I696763,I696780,I696576,I1049476,I696820,I696828,I696845,I696862,I696879,I696579,I696910,I1049479,I696927,I696953,I696961,I696561,I696992,I696570,I697023,I697040,I696582,I697071,I1049473,I696573,I696564,I696567,I696585,I697171,I697197,I697205,I697222,I697239,I697265,I697273,I697299,I697307,I697324,I697341,I697358,I697398,I697406,I697423,I697440,I697457,I697488,I697505,I697531,I697539,I697570,I697601,I697618,I697649,I697749,I697775,I697783,I697800,I697817,I697843,I697851,I697877,I697885,I697902,I697919,I697936,I697976,I697984,I698001,I698018,I698035,I698066,I698083,I698109,I698117,I698148,I698179,I698196,I698227,I698327,I1144189,I698353,I698361,I698378,I1144171,I1144183,I698395,I1144186,I698421,I698429,I1144180,I1144177,I698455,I698463,I698480,I698497,I698514,I1144195,I698554,I698562,I698579,I698596,I698613,I698644,I1144174,I698661,I698687,I698695,I698726,I698757,I698774,I698805,I1144192,I698905,I1173089,I698931,I698939,I698956,I1173071,I1173083,I698973,I1173086,I698999,I699007,I1173080,I1173077,I699033,I699041,I699058,I699075,I699092,I1173095,I699132,I699140,I699157,I699174,I699191,I699222,I1173074,I699239,I699265,I699273,I699304,I699335,I699352,I699383,I1173092,I699483,I699509,I699517,I699534,I699551,I699577,I699585,I699611,I699619,I699636,I699653,I699670,I699466,I699710,I699718,I699735,I699752,I699769,I699469,I699800,I699817,I699843,I699851,I699451,I699882,I699460,I699913,I699930,I699472,I699961,I699463,I699454,I699457,I699475,I700061,I700087,I700095,I700112,I700129,I700155,I700163,I700189,I700197,I700214,I700231,I700248,I700044,I700288,I700296,I700313,I700330,I700347,I700047,I700378,I700395,I700421,I700429,I700029,I700460,I700038,I700491,I700508,I700050,I700539,I700041,I700032,I700035,I700053,I700639,I700665,I700673,I700690,I700707,I700733,I700741,I700767,I700775,I700792,I700809,I700826,I700866,I700874,I700891,I700908,I700925,I700956,I700973,I700999,I701007,I701038,I701069,I701086,I701117,I701217,I701243,I701251,I701268,I701285,I701311,I701319,I701345,I701353,I701370,I701387,I701404,I701200,I701444,I701452,I701469,I701486,I701503,I701203,I701534,I701551,I701577,I701585,I701185,I701616,I701194,I701647,I701664,I701206,I701695,I701197,I701188,I701191,I701209,I701795,I701821,I701829,I701846,I701863,I701889,I701897,I701923,I701931,I701948,I701965,I701982,I701778,I702022,I702030,I702047,I702064,I702081,I701781,I702112,I702129,I702155,I702163,I701763,I702194,I701772,I702225,I702242,I701784,I702273,I701775,I701766,I701769,I701787,I702373,I1012445,I702399,I702407,I702424,I1012421,I1012436,I702441,I1012448,I702467,I702475,I1012433,I1012424,I702501,I702509,I702526,I702543,I702560,I702356,I702600,I702608,I702625,I702642,I702659,I702359,I702690,I1012439,I1012430,I702707,I1012442,I702733,I702741,I702341,I702772,I702350,I702803,I702820,I702362,I702851,I1012427,I702353,I702344,I702347,I702365,I702951,I811598,I702977,I702985,I703002,I811586,I811604,I703019,I811601,I703045,I703053,I811592,I811589,I703079,I703087,I703104,I703121,I703138,I811583,I703178,I703186,I703203,I703220,I703237,I703268,I703285,I703311,I703319,I703350,I703381,I703398,I703429,I811595,I703529,I991773,I703555,I703563,I703580,I991749,I991764,I703597,I991776,I703623,I703631,I991761,I991752,I703657,I703665,I703682,I703699,I703716,I703512,I703756,I703764,I703781,I703798,I703815,I703515,I703846,I991767,I991758,I703863,I991770,I703889,I703897,I703497,I703928,I703506,I703959,I703976,I703518,I704007,I991755,I703509,I703500,I703503,I703521,I704107,I1141299,I704133,I704141,I704158,I1141281,I1141293,I704175,I1141296,I704201,I704209,I1141290,I1141287,I704235,I704243,I704260,I704277,I704294,I704090,I1141305,I704334,I704342,I704359,I704376,I704393,I704093,I704424,I1141284,I704441,I704467,I704475,I704075,I704506,I704084,I704537,I704554,I704096,I704585,I1141302,I704087,I704078,I704081,I704099,I704685,I1290643,I704711,I704719,I704736,I1290667,I1290649,I704753,I1290655,I704779,I704787,I1290661,I1290646,I704813,I704821,I704838,I704855,I704872,I1290658,I704912,I704920,I704937,I704954,I704971,I705002,I1290664,I1290652,I705019,I705045,I705053,I705084,I705115,I705132,I705163,I705263,I827408,I705289,I705297,I705314,I827396,I827414,I705331,I827411,I705357,I705365,I827402,I827399,I705391,I705399,I705416,I705433,I705450,I827393,I705490,I705498,I705515,I705532,I705549,I705580,I705597,I705623,I705631,I705662,I705693,I705710,I705741,I827405,I705841,I705867,I705875,I705892,I705909,I705935,I705943,I705969,I705977,I705994,I706011,I706028,I706068,I706076,I706093,I706110,I706127,I706158,I706175,I706201,I706209,I706240,I706271,I706288,I706319,I706419,I1207191,I706445,I706453,I706470,I1207173,I1207185,I706487,I1207188,I706513,I706521,I1207182,I1207179,I706547,I706555,I706572,I706589,I706606,I706402,I1207197,I706646,I706654,I706671,I706688,I706705,I706405,I706736,I1207176,I706753,I706779,I706787,I706387,I706818,I706396,I706849,I706866,I706408,I706897,I1207194,I706399,I706390,I706393,I706411,I706997,I707023,I707031,I707048,I707065,I707091,I707099,I707125,I707133,I707150,I707167,I707184,I706980,I707224,I707232,I707249,I707266,I707283,I706983,I707314,I707331,I707357,I707365,I706965,I707396,I706974,I707427,I707444,I706986,I707475,I706977,I706968,I706971,I706989,I707575,I1378560,I707601,I707609,I707626,I1378545,I1378533,I707643,I1378548,I707669,I707677,I1378551,I707703,I707711,I707728,I707745,I707762,I707558,I1378539,I707802,I707810,I707827,I707844,I707861,I707561,I707892,I1378536,I1378542,I707909,I1378557,I707935,I707943,I707543,I707974,I707552,I708005,I708022,I707564,I708053,I1378554,I707555,I707546,I707549,I707567,I708153,I973685,I708179,I708187,I708204,I973661,I973676,I708221,I973688,I708247,I708255,I973673,I973664,I708281,I708289,I708306,I708323,I708340,I708380,I708388,I708405,I708422,I708439,I708470,I973679,I973670,I708487,I973682,I708513,I708521,I708552,I708583,I708600,I708631,I973667,I708731,I708757,I708765,I708782,I708799,I708825,I708833,I708859,I708867,I708884,I708901,I708918,I708714,I708958,I708966,I708983,I709000,I709017,I708717,I709048,I709065,I709091,I709099,I708699,I709130,I708708,I709161,I709178,I708720,I709209,I708711,I708702,I708705,I708723,I709309,I816868,I709335,I709343,I709360,I816856,I816874,I709377,I816871,I709403,I709411,I816862,I816859,I709437,I709445,I709462,I709479,I709496,I709292,I816853,I709536,I709544,I709561,I709578,I709595,I709295,I709626,I709643,I709669,I709677,I709277,I709708,I709286,I709739,I709756,I709298,I709787,I816865,I709289,I709280,I709283,I709301,I709887,I1374395,I709913,I709921,I709938,I1374380,I1374368,I709955,I1374383,I709981,I709989,I1374386,I710015,I710023,I710040,I710057,I710074,I709870,I1374374,I710114,I710122,I710139,I710156,I710173,I709873,I710204,I1374371,I1374377,I710221,I1374392,I710247,I710255,I709855,I710286,I709864,I710317,I710334,I709876,I710365,I1374389,I709867,I709858,I709861,I709879,I710465,I1026011,I710491,I710499,I710516,I1025987,I1026002,I710533,I1026014,I710559,I710567,I1025999,I1025990,I710593,I710601,I710618,I710635,I710652,I710448,I710692,I710700,I710717,I710734,I710751,I710451,I710782,I1026005,I1025996,I710799,I1026008,I710825,I710833,I710433,I710864,I710442,I710895,I710912,I710454,I710943,I1025993,I710445,I710436,I710439,I710457,I711043,I711069,I711077,I711094,I711111,I711137,I711145,I711171,I711179,I711196,I711213,I711230,I711270,I711278,I711295,I711312,I711329,I711360,I711377,I711403,I711411,I711442,I711473,I711490,I711521,I711621,I958181,I711647,I711655,I711672,I958157,I958172,I711689,I958184,I711715,I711723,I958169,I958160,I711749,I711757,I711774,I711791,I711808,I711848,I711856,I711873,I711890,I711907,I711938,I958175,I958166,I711955,I958178,I711981,I711989,I712020,I712051,I712068,I712099,I958163,I712199,I712225,I712233,I712250,I712267,I712293,I712301,I712327,I712335,I712352,I712369,I712386,I712182,I712426,I712434,I712451,I712468,I712485,I712185,I712516,I712533,I712559,I712567,I712167,I712598,I712176,I712629,I712646,I712188,I712677,I712179,I712170,I712173,I712191,I712777,I1058446,I712803,I712811,I712828,I1058443,I1058461,I712845,I1058458,I712871,I712879,I1058440,I712905,I712913,I712930,I712947,I712964,I1058452,I713004,I713012,I713029,I713046,I713063,I713094,I1058455,I713111,I713137,I713145,I713176,I713207,I713224,I713255,I1058449,I713355,I1074154,I713381,I713389,I713406,I1074151,I1074169,I713423,I1074166,I713449,I713457,I1074148,I713483,I713491,I713508,I713525,I713542,I1074160,I713582,I713590,I713607,I713624,I713641,I713672,I1074163,I713689,I713715,I713723,I713754,I713785,I713802,I713833,I1074157,I713933,I1182915,I713959,I713967,I713984,I1182897,I1182909,I714001,I1182912,I714027,I714035,I1182906,I1182903,I714061,I714069,I714086,I714103,I714120,I1182921,I714160,I714168,I714185,I714202,I714219,I714250,I1182900,I714267,I714293,I714301,I714332,I714363,I714380,I714411,I1182918,I714511,I714537,I714545,I714562,I714579,I714605,I714613,I714639,I714647,I714664,I714681,I714698,I714738,I714746,I714763,I714780,I714797,I714828,I714845,I714871,I714879,I714910,I714941,I714958,I714989,I715089,I715115,I715123,I715140,I715157,I715183,I715191,I715217,I715225,I715242,I715259,I715276,I715072,I715316,I715324,I715341,I715358,I715375,I715075,I715406,I715423,I715449,I715457,I715057,I715488,I715066,I715519,I715536,I715078,I715567,I715069,I715060,I715063,I715081,I715667,I715693,I715701,I715718,I715735,I715761,I715769,I715795,I715803,I715820,I715837,I715854,I715894,I715902,I715919,I715936,I715953,I715984,I716001,I716027,I716035,I716066,I716097,I716114,I716145,I716245,I716271,I716279,I716296,I716313,I716339,I716347,I716373,I716381,I716398,I716415,I716432,I716228,I716472,I716480,I716497,I716514,I716531,I716231,I716562,I716579,I716605,I716613,I716213,I716644,I716222,I716675,I716692,I716234,I716723,I716225,I716216,I716219,I716237,I716823,I840056,I716849,I716857,I716874,I840044,I840062,I716891,I840059,I716917,I716925,I840050,I840047,I716951,I716959,I716976,I716993,I717010,I840041,I717050,I717058,I717075,I717092,I717109,I717140,I717157,I717183,I717191,I717222,I717253,I717270,I717301,I840053,I717401,I1001463,I717427,I717435,I717452,I1001439,I1001454,I717469,I1001466,I717495,I717503,I1001451,I1001442,I717529,I717537,I717554,I717571,I717588,I717384,I717628,I717636,I717653,I717670,I717687,I717387,I717718,I1001457,I1001448,I717735,I1001460,I717761,I717769,I717369,I717800,I717378,I717831,I717848,I717390,I717879,I1001445,I717381,I717372,I717375,I717393,I717979,I718005,I718013,I718030,I718047,I718073,I718081,I718107,I718115,I718132,I718149,I718166,I717962,I718206,I718214,I718231,I718248,I718265,I717965,I718296,I718313,I718339,I718347,I717947,I718378,I717956,I718409,I718426,I717968,I718457,I717959,I717950,I717953,I717971,I718557,I718583,I718591,I718608,I718625,I718651,I718659,I718685,I718693,I718710,I718727,I718744,I718784,I718792,I718809,I718826,I718843,I718874,I718891,I718917,I718925,I718956,I718987,I719004,I719035,I719135,I719161,I719169,I719186,I719203,I719229,I719237,I719263,I719271,I719288,I719305,I719322,I719118,I719362,I719370,I719387,I719404,I719421,I719121,I719452,I719469,I719495,I719503,I719103,I719534,I719112,I719565,I719582,I719124,I719613,I719115,I719106,I719109,I719127,I719713,I719739,I719747,I719764,I719781,I719807,I719815,I719841,I719849,I719866,I719883,I719900,I719696,I719940,I719948,I719965,I719982,I719999,I719699,I720030,I720047,I720073,I720081,I719681,I720112,I719690,I720143,I720160,I719702,I720191,I719693,I719684,I719687,I719705,I720291,I720317,I720325,I720342,I720359,I720385,I720393,I720419,I720427,I720444,I720461,I720478,I720518,I720526,I720543,I720560,I720577,I720608,I720625,I720651,I720659,I720690,I720721,I720738,I720769,I720869,I1261641,I720895,I720903,I720920,I1261644,I1261653,I720937,I1261656,I720963,I720971,I1261665,I1261647,I720997,I721005,I721022,I721039,I721056,I720852,I721096,I721104,I721121,I721138,I721155,I720855,I721186,I1261662,I721203,I1261659,I721229,I721237,I720837,I721268,I720846,I721299,I721316,I720858,I721347,I1261650,I720849,I720840,I720843,I720861,I721447,I906458,I721473,I721481,I721498,I906446,I906464,I721515,I906461,I721541,I721549,I906452,I906449,I721575,I721583,I721600,I721617,I721634,I721430,I906443,I721674,I721682,I721699,I721716,I721733,I721433,I721764,I721781,I721807,I721815,I721415,I721846,I721424,I721877,I721894,I721436,I721925,I906455,I721427,I721418,I721421,I721439,I722025,I722051,I722059,I722076,I722093,I722119,I722127,I722153,I722161,I722178,I722195,I722212,I722008,I722252,I722260,I722277,I722294,I722311,I722011,I722342,I722359,I722385,I722393,I721993,I722424,I722002,I722455,I722472,I722014,I722503,I722005,I721996,I721999,I722017,I722603,I722629,I722637,I722654,I722671,I722697,I722705,I722731,I722739,I722756,I722773,I722790,I722830,I722838,I722855,I722872,I722889,I722920,I722937,I722963,I722971,I723002,I723033,I723050,I723081,I723181,I723207,I723215,I723232,I723249,I723275,I723283,I723309,I723317,I723334,I723351,I723368,I723408,I723416,I723433,I723450,I723467,I723498,I723515,I723541,I723549,I723580,I723611,I723628,I723659,I723759,I723785,I723793,I723810,I723827,I723853,I723861,I723887,I723895,I723912,I723929,I723946,I723742,I723986,I723994,I724011,I724028,I724045,I723745,I724076,I724093,I724119,I724127,I723727,I724158,I723736,I724189,I724206,I723748,I724237,I723739,I723730,I723733,I723751,I724337,I1249129,I724363,I724371,I724388,I1249132,I1249141,I724405,I1249144,I724431,I724439,I1249153,I1249135,I724465,I724473,I724490,I724507,I724524,I724320,I724564,I724572,I724589,I724606,I724623,I724323,I724654,I1249150,I724671,I1249147,I724697,I724705,I724305,I724736,I724314,I724767,I724784,I724326,I724815,I1249138,I724317,I724308,I724311,I724329,I724915,I863244,I724941,I724949,I724966,I863232,I863250,I724983,I863247,I725009,I725017,I863238,I863235,I725043,I725051,I725068,I725085,I725102,I863229,I725142,I725150,I725167,I725184,I725201,I725232,I725249,I725275,I725283,I725314,I725345,I725362,I725393,I863241,I725493,I884324,I725519,I725527,I725544,I884312,I884330,I725561,I884327,I725587,I725595,I884318,I884315,I725621,I725629,I725646,I725663,I725680,I884309,I725720,I725728,I725745,I725762,I725779,I725810,I725827,I725853,I725861,I725892,I725923,I725940,I725971,I884321,I726071,I726097,I726105,I726122,I726139,I726165,I726173,I726199,I726207,I726224,I726241,I726258,I726054,I726298,I726306,I726323,I726340,I726357,I726057,I726388,I726405,I726431,I726439,I726039,I726470,I726048,I726501,I726518,I726060,I726549,I726051,I726042,I726045,I726063,I726649,I726675,I726683,I726700,I726717,I726743,I726751,I726777,I726785,I726802,I726819,I726836,I726876,I726884,I726901,I726918,I726935,I726966,I726983,I727009,I727017,I727048,I727079,I727096,I727127,I727227,I727253,I727261,I727278,I727295,I727321,I727329,I727355,I727363,I727380,I727397,I727414,I727454,I727462,I727479,I727496,I727513,I727544,I727561,I727587,I727595,I727626,I727657,I727674,I727705,I727805,I835313,I727831,I727839,I727856,I835301,I835319,I727873,I835316,I727899,I727907,I835307,I835304,I727933,I727941,I727958,I727975,I727992,I727788,I835298,I728032,I728040,I728057,I728074,I728091,I727791,I728122,I728139,I728165,I728173,I727773,I728204,I727782,I728235,I728252,I727794,I728283,I835310,I727785,I727776,I727779,I727797,I728383,I728409,I728417,I728434,I728451,I728477,I728485,I728511,I728519,I728536,I728553,I728570,I728366,I728610,I728618,I728635,I728652,I728669,I728369,I728700,I728717,I728743,I728751,I728351,I728782,I728360,I728813,I728830,I728372,I728861,I728363,I728354,I728357,I728375,I728961,I1389270,I728987,I728995,I729012,I1389255,I1389243,I729029,I1389258,I729055,I729063,I1389261,I729089,I729097,I729114,I729131,I729148,I1389249,I729188,I729196,I729213,I729230,I729247,I729278,I1389246,I1389252,I729295,I1389267,I729321,I729329,I729360,I729391,I729408,I729439,I1389264,I729539,I1138409,I729565,I729573,I729590,I1138391,I1138403,I729607,I1138406,I729633,I729641,I1138400,I1138397,I729667,I729675,I729692,I729709,I729726,I1138415,I729766,I729774,I729791,I729808,I729825,I729856,I1138394,I729873,I729899,I729907,I729938,I729969,I729986,I730017,I1138412,I730117,I730143,I730151,I730168,I730185,I730211,I730219,I730245,I730253,I730270,I730287,I730304,I730100,I730344,I730352,I730369,I730386,I730403,I730103,I730434,I730451,I730477,I730485,I730085,I730516,I730094,I730547,I730564,I730106,I730595,I730097,I730088,I730091,I730109,I730695,I882216,I730721,I730729,I730746,I882204,I882222,I730763,I882219,I730789,I730797,I882210,I882207,I730823,I730831,I730848,I730865,I730882,I730678,I882201,I730922,I730930,I730947,I730964,I730981,I730681,I731012,I731029,I731055,I731063,I730663,I731094,I730672,I731125,I731142,I730684,I731173,I882213,I730675,I730666,I730669,I730687,I731273,I1301625,I731299,I731307,I731324,I1301649,I1301631,I731341,I1301637,I731367,I731375,I1301643,I1301628,I731401,I731409,I731426,I731443,I731460,I731256,I1301640,I731500,I731508,I731525,I731542,I731559,I731259,I731590,I1301646,I1301634,I731607,I731633,I731641,I731241,I731672,I731250,I731703,I731720,I731262,I731751,I731253,I731244,I731247,I731265,I731851,I1204301,I731877,I731885,I731902,I1204283,I1204295,I731919,I1204298,I731945,I731953,I1204292,I1204289,I731979,I731987,I732004,I732021,I732038,I731834,I1204307,I732078,I732086,I732103,I732120,I732137,I731837,I732168,I1204286,I732185,I732211,I732219,I731819,I732250,I731828,I732281,I732298,I731840,I732329,I1204304,I731831,I731822,I731825,I731843,I732429,I732455,I732463,I732480,I732497,I732523,I732531,I732557,I732565,I732582,I732599,I732616,I732656,I732664,I732681,I732698,I732715,I732746,I732763,I732789,I732797,I732828,I732859,I732876,I732907,I733007,I733033,I733041,I733058,I733075,I733101,I733109,I733135,I733143,I733160,I733177,I733194,I733234,I733242,I733259,I733276,I733293,I733324,I733341,I733367,I733375,I733406,I733437,I733454,I733485,I733585,I1050592,I733611,I733619,I733636,I1050589,I1050607,I733653,I1050604,I733679,I733687,I1050586,I733713,I733721,I733738,I733755,I733772,I1050598,I733812,I733820,I733837,I733854,I733871,I733902,I1050601,I733919,I733945,I733953,I733984,I734015,I734032,I734063,I1050595,I734163,I734189,I734197,I734214,I734231,I734257,I734265,I734291,I734299,I734316,I734333,I734350,I734390,I734398,I734415,I734432,I734449,I734480,I734497,I734523,I734531,I734562,I734593,I734610,I734641,I734741,I734767,I734775,I734792,I734809,I734835,I734843,I734869,I734877,I734894,I734911,I734928,I734724,I734968,I734976,I734993,I735010,I735027,I734727,I735058,I735075,I735101,I735109,I734709,I735140,I734718,I735171,I735188,I734730,I735219,I734721,I734712,I734715,I734733,I735319,I735345,I735353,I735370,I735387,I735413,I735421,I735447,I735455,I735472,I735489,I735506,I735546,I735554,I735571,I735588,I735605,I735636,I735653,I735679,I735687,I735718,I735749,I735766,I735797,I735897,I1145345,I735923,I735931,I735948,I1145327,I1145339,I735965,I1145342,I735991,I735999,I1145336,I1145333,I736025,I736033,I736050,I736067,I736084,I1145351,I736124,I736132,I736149,I736166,I736183,I736214,I1145330,I736231,I736257,I736265,I736296,I736327,I736344,I736375,I1145348,I736475,I920067,I736501,I736509,I736526,I920043,I920058,I736543,I920070,I736569,I736577,I920055,I920046,I736603,I736611,I736628,I736645,I736662,I736702,I736710,I736727,I736744,I736761,I736792,I920061,I920052,I736809,I920064,I736835,I736843,I736874,I736905,I736922,I736953,I920049,I737053,I1201411,I737079,I737087,I737104,I1201393,I1201405,I737121,I1201408,I737147,I737155,I1201402,I1201399,I737181,I737189,I737206,I737223,I737240,I737036,I1201417,I737280,I737288,I737305,I737322,I737339,I737039,I737370,I1201396,I737387,I737413,I737421,I737021,I737452,I737030,I737483,I737500,I737042,I737531,I1201414,I737033,I737024,I737027,I737045,I737631,I737657,I737665,I737682,I737699,I737725,I737733,I737759,I737767,I737784,I737801,I737818,I737858,I737866,I737883,I737900,I737917,I737948,I737965,I737991,I737999,I738030,I738061,I738078,I738109,I738209,I738235,I738243,I738260,I738277,I738303,I738311,I738337,I738345,I738362,I738379,I738396,I738436,I738444,I738461,I738478,I738495,I738526,I738543,I738569,I738577,I738608,I738639,I738656,I738687,I738787,I1370230,I738813,I738821,I738838,I1370215,I1370203,I738855,I1370218,I738881,I738889,I1370221,I738915,I738923,I738940,I738957,I738974,I738770,I1370209,I739014,I739022,I739039,I739056,I739073,I738773,I739104,I1370206,I1370212,I739121,I1370227,I739147,I739155,I738755,I739186,I738764,I739217,I739234,I738776,I739265,I1370224,I738767,I738758,I738761,I738779,I739365,I1188117,I739391,I739399,I739416,I1188099,I1188111,I739433,I1188114,I739459,I739467,I1188108,I1188105,I739493,I739501,I739518,I739535,I739552,I739348,I1188123,I739592,I739600,I739617,I739634,I739651,I739351,I739682,I1188102,I739699,I739725,I739733,I739333,I739764,I739342,I739795,I739812,I739354,I739843,I1188120,I739345,I739336,I739339,I739357,I739943,I739969,I739977,I739994,I740011,I740037,I740045,I740071,I740079,I740096,I740113,I740130,I739926,I740170,I740178,I740195,I740212,I740229,I739929,I740260,I740277,I740303,I740311,I739911,I740342,I739920,I740373,I740390,I739932,I740421,I739923,I739914,I739917,I739935,I740521,I740547,I740555,I740572,I740589,I740615,I740623,I740649,I740657,I740674,I740691,I740708,I740748,I740756,I740773,I740790,I740807,I740838,I740855,I740881,I740889,I740920,I740951,I740968,I740999,I741099,I741125,I741133,I741150,I741167,I741193,I741201,I741227,I741235,I741252,I741269,I741286,I741326,I741334,I741351,I741368,I741385,I741416,I741433,I741459,I741467,I741498,I741529,I741546,I741577,I741677,I993065,I741703,I741711,I741728,I993041,I993056,I741745,I993068,I741771,I741779,I993053,I993044,I741805,I741813,I741830,I741847,I741864,I741904,I741912,I741929,I741946,I741963,I741994,I993059,I993050,I742011,I993062,I742037,I742045,I742076,I742107,I742124,I742155,I993047,I742255,I1070227,I742281,I742289,I742306,I1070224,I1070242,I742323,I1070239,I742349,I742357,I1070221,I742383,I742391,I742408,I742425,I742442,I742238,I1070233,I742482,I742490,I742507,I742524,I742541,I742241,I742572,I1070236,I742589,I742615,I742623,I742223,I742654,I742232,I742685,I742702,I742244,I742733,I1070230,I742235,I742226,I742229,I742247,I742833,I742859,I742867,I742884,I742901,I742927,I742935,I742961,I742969,I742986,I743003,I743020,I742816,I743060,I743068,I743085,I743102,I743119,I742819,I743150,I743167,I743193,I743201,I742801,I743232,I742810,I743263,I743280,I742822,I743311,I742813,I742804,I742807,I742825,I743411,I743437,I743445,I743462,I743479,I743505,I743513,I743539,I743547,I743564,I743581,I743598,I743638,I743646,I743663,I743680,I743697,I743728,I743745,I743771,I743779,I743810,I743841,I743858,I743889,I743989,I744015,I744023,I744040,I744057,I744083,I744091,I744117,I744125,I744142,I744159,I744176,I743972,I744216,I744224,I744241,I744258,I744275,I743975,I744306,I744323,I744349,I744357,I743957,I744388,I743966,I744419,I744436,I743978,I744467,I743969,I743960,I743963,I743981,I744567,I744593,I744601,I744618,I744635,I744661,I744669,I744695,I744703,I744720,I744737,I744754,I744550,I744794,I744802,I744819,I744836,I744853,I744553,I744884,I744901,I744927,I744935,I744535,I744966,I744544,I744997,I745014,I744556,I745045,I744547,I744538,I744541,I744559,I745145,I745171,I745179,I745196,I745213,I745239,I745247,I745273,I745281,I745298,I745315,I745332,I745372,I745380,I745397,I745414,I745431,I745462,I745479,I745505,I745513,I745544,I745575,I745592,I745623,I745723,I745749,I745757,I745774,I745791,I745817,I745825,I745851,I745859,I745876,I745893,I745910,I745950,I745958,I745975,I745992,I746009,I746040,I746057,I746083,I746091,I746122,I746153,I746170,I746201,I746301,I1314341,I746327,I746335,I746352,I1314365,I1314347,I746369,I1314353,I746395,I746403,I1314359,I1314344,I746429,I746437,I746454,I746471,I746488,I746284,I1314356,I746528,I746536,I746553,I746570,I746587,I746287,I746618,I1314362,I1314350,I746635,I746661,I746669,I746269,I746700,I746278,I746731,I746748,I746290,I746779,I746281,I746272,I746275,I746293,I746879,I1376180,I746905,I746913,I746930,I1376165,I1376153,I746947,I1376168,I746973,I746981,I1376171,I747007,I747015,I747032,I747049,I747066,I1376159,I747106,I747114,I747131,I747148,I747165,I747196,I1376156,I1376162,I747213,I1376177,I747239,I747247,I747278,I747309,I747326,I747357,I1376174,I747457,I747483,I747491,I747508,I747525,I747551,I747559,I747585,I747593,I747610,I747627,I747644,I747684,I747692,I747709,I747726,I747743,I747774,I747791,I747817,I747825,I747856,I747887,I747904,I747935,I748035,I1338100,I748061,I748069,I748086,I1338085,I1338073,I748103,I1338088,I748129,I748137,I1338091,I748163,I748171,I748188,I748205,I748222,I1338079,I748262,I748270,I748287,I748304,I748321,I748352,I1338076,I1338082,I748369,I1338097,I748395,I748403,I748434,I748465,I748482,I748513,I1338094,I748613,I1236669,I748639,I748647,I748664,I1236651,I1236663,I748681,I1236666,I748707,I748715,I1236660,I1236657,I748741,I748749,I748766,I748783,I748800,I1236675,I748840,I748848,I748865,I748882,I748899,I748930,I1236654,I748947,I748973,I748981,I749012,I749043,I749060,I749091,I1236672,I749191,I1279593,I749217,I749225,I749242,I1279596,I1279605,I749259,I1279608,I749285,I749293,I1279617,I1279599,I749319,I749327,I749344,I749361,I749378,I749418,I749426,I749443,I749460,I749477,I749508,I1279614,I749525,I1279611,I749551,I749559,I749590,I749621,I749638,I749669,I1279602,I749769,I1292955,I749795,I749803,I749820,I1292979,I1292961,I749837,I1292967,I749863,I749871,I1292973,I1292958,I749897,I749905,I749922,I749939,I749956,I1292970,I749996,I750004,I750021,I750038,I750055,I750086,I1292976,I1292964,I750103,I750129,I750137,I750168,I750199,I750216,I750247,I750347,I750373,I750381,I750398,I750415,I750441,I750449,I750475,I750483,I750500,I750517,I750534,I750330,I750574,I750582,I750599,I750616,I750633,I750333,I750664,I750681,I750707,I750715,I750315,I750746,I750324,I750777,I750794,I750336,I750825,I750327,I750318,I750321,I750339,I750925,I826354,I750951,I750959,I750976,I826342,I826360,I750993,I826357,I751019,I751027,I826348,I826345,I751053,I751061,I751078,I751095,I751112,I826339,I751152,I751160,I751177,I751194,I751211,I751242,I751259,I751285,I751293,I751324,I751355,I751372,I751403,I826351,I751503,I751529,I751537,I751554,I751571,I751597,I751605,I751631,I751639,I751656,I751673,I751690,I751730,I751738,I751755,I751772,I751789,I751820,I751837,I751863,I751871,I751902,I751933,I751950,I751981,I752081,I1241871,I752107,I752115,I752132,I1241853,I1241865,I752149,I1241868,I752175,I752183,I1241862,I1241859,I752209,I752217,I752234,I752251,I752268,I1241877,I752308,I752316,I752333,I752350,I752367,I752398,I1241856,I752415,I752441,I752449,I752480,I752511,I752528,I752559,I1241874,I752659,I1259465,I752685,I752693,I752710,I1259468,I1259477,I752727,I1259480,I752753,I752761,I1259489,I1259471,I752787,I752795,I752812,I752829,I752846,I752886,I752894,I752911,I752928,I752945,I752976,I1259486,I752993,I1259483,I753019,I753027,I753058,I753089,I753106,I753137,I1259474,I753237,I960765,I753263,I753271,I753288,I960741,I960756,I753305,I960768,I753331,I753339,I960753,I960744,I753365,I753373,I753390,I753407,I753424,I753220,I753464,I753472,I753489,I753506,I753523,I753223,I753554,I960759,I960750,I753571,I960762,I753597,I753605,I753205,I753636,I753214,I753667,I753684,I753226,I753715,I960747,I753217,I753208,I753211,I753229,I753815,I753841,I753849,I753866,I753883,I753909,I753917,I753943,I753951,I753968,I753985,I754002,I753798,I754042,I754050,I754067,I754084,I754101,I753801,I754132,I754149,I754175,I754183,I753783,I754214,I753792,I754245,I754262,I753804,I754293,I753795,I753786,I753789,I753807,I754393,I754419,I754427,I754444,I754461,I754487,I754495,I754521,I754529,I754546,I754563,I754580,I754376,I754620,I754628,I754645,I754662,I754679,I754379,I754710,I754727,I754753,I754761,I754361,I754792,I754370,I754823,I754840,I754382,I754871,I754373,I754364,I754367,I754385,I754971,I754997,I755005,I755022,I755039,I755065,I755073,I755099,I755107,I755124,I755141,I755158,I754954,I755198,I755206,I755223,I755240,I755257,I754957,I755288,I755305,I755331,I755339,I754939,I755370,I754948,I755401,I755418,I754960,I755449,I754951,I754942,I754945,I754963,I755549,I755575,I755583,I755600,I755617,I755643,I755651,I755677,I755685,I755702,I755719,I755736,I755776,I755784,I755801,I755818,I755835,I755866,I755883,I755909,I755917,I755948,I755979,I755996,I756027,I756127,I756153,I756161,I756178,I756195,I756221,I756229,I756255,I756263,I756280,I756297,I756314,I756354,I756362,I756379,I756396,I756413,I756444,I756461,I756487,I756495,I756526,I756557,I756574,I756605,I756705,I1123381,I756731,I756739,I756756,I1123363,I1123375,I756773,I1123378,I756799,I756807,I1123372,I1123369,I756833,I756841,I756858,I756875,I756892,I1123387,I756932,I756940,I756957,I756974,I756991,I757022,I1123366,I757039,I757065,I757073,I757104,I757135,I757152,I757183,I1123384,I757283,I757309,I757317,I757334,I757351,I757377,I757385,I757411,I757419,I757436,I757453,I757470,I757266,I757510,I757518,I757535,I757552,I757569,I757269,I757600,I757617,I757643,I757651,I757251,I757682,I757260,I757713,I757730,I757272,I757761,I757263,I757254,I757257,I757275,I757861,I757887,I757895,I757912,I757929,I757955,I757963,I757989,I757997,I758014,I758031,I758048,I758088,I758096,I758113,I758130,I758147,I758178,I758195,I758221,I758229,I758260,I758291,I758308,I758339,I758439,I758465,I758473,I758490,I758507,I758533,I758541,I758567,I758575,I758592,I758609,I758626,I758422,I758666,I758674,I758691,I758708,I758725,I758425,I758756,I758773,I758799,I758807,I758407,I758838,I758416,I758869,I758886,I758428,I758917,I758419,I758410,I758413,I758431,I759017,I1394625,I759043,I759051,I759068,I1394610,I1394598,I759085,I1394613,I759111,I759119,I1394616,I759145,I759153,I759170,I759187,I759204,I1394604,I759244,I759252,I759269,I759286,I759303,I759334,I1394601,I1394607,I759351,I1394622,I759377,I759385,I759416,I759447,I759464,I759495,I1394619,I759595,I1342265,I759621,I759629,I759646,I1342250,I1342238,I759663,I1342253,I759689,I759697,I1342256,I759723,I759731,I759748,I759765,I759782,I1342244,I759822,I759830,I759847,I759864,I759881,I759912,I1342241,I1342247,I759929,I1342262,I759955,I759963,I759994,I760025,I760042,I760073,I1342259,I760173,I760199,I760207,I760224,I760241,I760267,I760275,I760301,I760309,I760326,I760343,I760360,I760400,I760408,I760425,I760442,I760459,I760490,I760507,I760533,I760541,I760572,I760603,I760620,I760651,I760751,I760777,I760785,I760802,I760819,I760845,I760853,I760879,I760887,I760904,I760921,I760938,I760734,I760978,I760986,I761003,I761020,I761037,I760737,I761068,I761085,I761111,I761119,I760719,I761150,I760728,I761181,I761198,I760740,I761229,I760731,I760722,I760725,I760743,I761329,I761355,I761363,I761380,I761397,I761423,I761431,I761457,I761465,I761482,I761499,I761516,I761556,I761564,I761581,I761598,I761615,I761646,I761663,I761689,I761697,I761728,I761759,I761776,I761807,I761907,I1176557,I761933,I761941,I761958,I1176539,I1176551,I761975,I1176554,I762001,I762009,I1176548,I1176545,I762035,I762043,I762060,I762077,I762094,I1176563,I762134,I762142,I762159,I762176,I762193,I762224,I1176542,I762241,I762267,I762275,I762306,I762337,I762354,I762385,I1176560,I762485,I762511,I762519,I762536,I762553,I762579,I762587,I762613,I762621,I762638,I762655,I762672,I762468,I762712,I762720,I762737,I762754,I762771,I762471,I762802,I762819,I762845,I762853,I762453,I762884,I762462,I762915,I762932,I762474,I762963,I762465,I762456,I762459,I762477,I763063,I763089,I763097,I763114,I763131,I763157,I763165,I763191,I763199,I763216,I763233,I763250,I763290,I763298,I763315,I763332,I763349,I763380,I763397,I763423,I763431,I763462,I763493,I763510,I763541,I763641,I1155749,I763667,I763675,I763692,I1155731,I1155743,I763709,I1155746,I763735,I763743,I1155740,I1155737,I763769,I763777,I763794,I763811,I763828,I763624,I1155755,I763868,I763876,I763893,I763910,I763927,I763627,I763958,I1155734,I763975,I764001,I764009,I763609,I764040,I763618,I764071,I764088,I763630,I764119,I1155752,I763621,I763612,I763615,I763633,I764219,I1304515,I764245,I764253,I764270,I1304539,I1304521,I764287,I1304527,I764313,I764321,I1304533,I1304518,I764347,I764355,I764372,I764389,I764406,I1304530,I764446,I764454,I764471,I764488,I764505,I764536,I1304536,I1304524,I764553,I764579,I764587,I764618,I764649,I764666,I764697,I764797,I764823,I764831,I764848,I764865,I764891,I764899,I764925,I764933,I764950,I764967,I764984,I765024,I765032,I765049,I765066,I765083,I765114,I765131,I765157,I765165,I765196,I765227,I765244,I765275,I765375,I765401,I765409,I765426,I765443,I765469,I765477,I765503,I765511,I765528,I765545,I765562,I765602,I765610,I765627,I765644,I765661,I765692,I765709,I765735,I765743,I765774,I765805,I765822,I765853,I765953,I1106619,I765979,I765987,I766004,I1106601,I1106613,I766021,I1106616,I766047,I766055,I1106610,I1106607,I766081,I766089,I766106,I766123,I766140,I765936,I1106625,I766180,I766188,I766205,I766222,I766239,I765939,I766270,I1106604,I766287,I766313,I766321,I765921,I766352,I765930,I766383,I766400,I765942,I766431,I1106622,I765933,I765924,I765927,I765945,I766531,I766557,I766565,I766582,I766599,I766625,I766633,I766659,I766667,I766684,I766701,I766718,I766514,I766758,I766766,I766783,I766800,I766817,I766517,I766848,I766865,I766891,I766899,I766499,I766930,I766508,I766961,I766978,I766520,I767009,I766511,I766502,I766505,I766523,I767109,I767135,I767143,I767160,I767177,I767203,I767211,I767237,I767245,I767262,I767279,I767296,I767336,I767344,I767361,I767378,I767395,I767426,I767443,I767469,I767477,I767508,I767539,I767556,I767587,I767687,I1312607,I767713,I767721,I767738,I1312631,I1312613,I767755,I1312619,I767781,I767789,I1312625,I1312610,I767815,I767823,I767840,I767857,I767874,I1312622,I767914,I767922,I767939,I767956,I767973,I768004,I1312628,I1312616,I768021,I768047,I768055,I768086,I768117,I768134,I768165,I768265,I768291,I768299,I768316,I768333,I768359,I768367,I768393,I768401,I768418,I768435,I768452,I768492,I768500,I768517,I768534,I768551,I768582,I768599,I768625,I768633,I768664,I768695,I768712,I768743,I768843,I768869,I768877,I768894,I768911,I768937,I768945,I768971,I768979,I768996,I769013,I769030,I768826,I769070,I769078,I769095,I769112,I769129,I768829,I769160,I769177,I769203,I769211,I768811,I769242,I768820,I769273,I769290,I768832,I769321,I768823,I768814,I768817,I768835,I769421,I1379155,I769447,I769455,I769472,I1379140,I1379128,I769489,I1379143,I769515,I769523,I1379146,I769549,I769557,I769574,I769591,I769608,I769404,I1379134,I769648,I769656,I769673,I769690,I769707,I769407,I769738,I1379131,I1379137,I769755,I1379152,I769781,I769789,I769389,I769820,I769398,I769851,I769868,I769410,I769899,I1379149,I769401,I769392,I769395,I769413,I769999,I1392840,I770025,I770033,I770050,I1392825,I1392813,I770067,I1392828,I770093,I770101,I1392831,I770127,I770135,I770152,I770169,I770186,I769982,I1392819,I770226,I770234,I770251,I770268,I770285,I769985,I770316,I1392816,I1392822,I770333,I1392837,I770359,I770367,I769967,I770398,I769976,I770429,I770446,I769988,I770477,I1392834,I769979,I769970,I769973,I769991,I770577,I1280137,I770603,I770611,I770628,I1280140,I1280149,I770645,I1280152,I770671,I770679,I1280161,I1280143,I770705,I770713,I770730,I770747,I770764,I770804,I770812,I770829,I770846,I770863,I770894,I1280158,I770911,I1280155,I770937,I770945,I770976,I771007,I771024,I771055,I1280146,I771155,I771181,I771189,I771206,I771223,I771249,I771257,I771283,I771291,I771308,I771325,I771342,I771382,I771390,I771407,I771424,I771441,I771472,I771489,I771515,I771523,I771554,I771585,I771602,I771633,I771733,I1288331,I771759,I771767,I771784,I1288355,I1288337,I771801,I1288343,I771827,I771835,I1288349,I1288334,I771861,I771869,I771886,I771903,I771920,I771716,I1288346,I771960,I771968,I771985,I772002,I772019,I771719,I772050,I1288352,I1288340,I772067,I772093,I772101,I771701,I772132,I771710,I772163,I772180,I771722,I772211,I771713,I771704,I771707,I771725,I772311,I772337,I772345,I772362,I772379,I772405,I772413,I772439,I772447,I772464,I772481,I772498,I772294,I772538,I772546,I772563,I772580,I772597,I772297,I772628,I772645,I772671,I772679,I772279,I772710,I772288,I772741,I772758,I772300,I772789,I772291,I772282,I772285,I772303,I772889,I1080886,I772915,I772923,I772940,I1080883,I1080901,I772957,I1080898,I772983,I772991,I1080880,I773017,I773025,I773042,I773059,I773076,I772872,I1080892,I773116,I773124,I773141,I773158,I773175,I772875,I773206,I1080895,I773223,I773249,I773257,I772857,I773288,I772866,I773319,I773336,I772878,I773367,I1080889,I772869,I772860,I772863,I772881,I773467,I1309139,I773493,I773501,I773518,I1309163,I1309145,I773535,I1309151,I773561,I773569,I1309157,I1309142,I773595,I773603,I773620,I773637,I773654,I1309154,I773694,I773702,I773719,I773736,I773753,I773784,I1309160,I1309148,I773801,I773827,I773835,I773866,I773897,I773914,I773945,I774045,I774071,I774079,I774096,I774113,I774139,I774147,I774173,I774181,I774198,I774215,I774232,I774272,I774280,I774297,I774314,I774331,I774362,I774379,I774405,I774413,I774444,I774475,I774492,I774523,I774623,I912782,I774649,I774657,I774674,I912770,I912788,I774691,I912785,I774717,I774725,I912776,I912773,I774751,I774759,I774776,I774793,I774810,I912767,I774850,I774858,I774875,I774892,I774909,I774940,I774957,I774983,I774991,I775022,I775053,I775070,I775101,I912779,I775201,I775227,I775235,I775252,I775269,I775295,I775303,I775329,I775337,I775354,I775371,I775388,I775184,I775428,I775436,I775453,I775470,I775487,I775187,I775518,I775535,I775561,I775569,I775169,I775600,I775178,I775631,I775648,I775190,I775679,I775181,I775172,I775175,I775193,I775779,I775805,I775813,I775830,I775847,I775873,I775881,I775907,I775915,I775932,I775949,I775966,I775762,I776006,I776014,I776031,I776048,I776065,I775765,I776096,I776113,I776139,I776147,I775747,I776178,I775756,I776209,I776226,I775768,I776257,I775759,I775750,I775753,I775771,I776357,I1179447,I776383,I776391,I776408,I1179429,I1179441,I776425,I1179444,I776451,I776459,I1179438,I1179435,I776485,I776493,I776510,I776527,I776544,I1179453,I776584,I776592,I776609,I776626,I776643,I776674,I1179432,I776691,I776717,I776725,I776756,I776787,I776804,I776835,I1179450,I776935,I776961,I776969,I776986,I777003,I777029,I777037,I777063,I777071,I777088,I777105,I777122,I777162,I777170,I777187,I777204,I777221,I777252,I777269,I777295,I777303,I777334,I777365,I777382,I777413,I777513,I1375585,I777539,I777547,I777564,I1375570,I1375558,I777581,I1375573,I777607,I777615,I1375576,I777641,I777649,I777666,I777683,I777700,I777496,I1375564,I777740,I777748,I777765,I777782,I777799,I777499,I777830,I1375561,I1375567,I777847,I1375582,I777873,I777881,I777481,I777912,I777490,I777943,I777960,I777502,I777991,I1375579,I777493,I777484,I777487,I777505,I778091,I778117,I778125,I778142,I778159,I778185,I778193,I778219,I778227,I778244,I778261,I778278,I778318,I778326,I778343,I778360,I778377,I778408,I778425,I778451,I778459,I778490,I778521,I778538,I778569,I778669,I1326987,I778695,I778703,I778720,I1326975,I1326993,I778737,I1326984,I778763,I778771,I1326999,I1326996,I778797,I778805,I778822,I778839,I778856,I1326978,I778896,I778904,I778921,I778938,I778955,I778986,I1326972,I779003,I1326981,I779029,I779037,I779068,I779099,I779116,I779147,I1326990,I779247,I779273,I779281,I779298,I779315,I779341,I779349,I779375,I779383,I779400,I779417,I779434,I779474,I779482,I779499,I779516,I779533,I779564,I779581,I779607,I779615,I779646,I779677,I779694,I779725,I779825,I866933,I779851,I779859,I779876,I866921,I866939,I779893,I866936,I779919,I779927,I866927,I866924,I779953,I779961,I779978,I779995,I780012,I866918,I780052,I780060,I780077,I780094,I780111,I780142,I780159,I780185,I780193,I780224,I780255,I780272,I780303,I866930,I780403,I1302203,I780429,I780437,I780454,I1302227,I1302209,I780471,I1302215,I780497,I780505,I1302221,I1302206,I780531,I780539,I780556,I780573,I780590,I1302218,I780630,I780638,I780655,I780672,I780689,I780720,I1302224,I1302212,I780737,I780763,I780771,I780802,I780833,I780850,I780881,I780981,I1285577,I781007,I781015,I781032,I1285580,I1285589,I781049,I1285592,I781075,I781083,I1285601,I1285583,I781109,I781117,I781134,I781151,I781168,I780964,I781208,I781216,I781233,I781250,I781267,I780967,I781298,I1285598,I781315,I1285595,I781341,I781349,I780949,I781380,I780958,I781411,I781428,I780970,I781459,I1285586,I780961,I780952,I780955,I780973,I781559,I846380,I781585,I781593,I781610,I846368,I846386,I781627,I846383,I781653,I781661,I846374,I846371,I781687,I781695,I781712,I781729,I781746,I781542,I846365,I781786,I781794,I781811,I781828,I781845,I781545,I781876,I781893,I781919,I781927,I781527,I781958,I781536,I781989,I782006,I781548,I782037,I846377,I781539,I781530,I781533,I781551,I782137,I782163,I782171,I782188,I782205,I782231,I782239,I782265,I782273,I782290,I782307,I782324,I782364,I782372,I782389,I782406,I782423,I782454,I782471,I782497,I782505,I782536,I782567,I782584,I782615,I782715,I782741,I782749,I782766,I782783,I782809,I782817,I782843,I782851,I782868,I782885,I782902,I782942,I782950,I782967,I782984,I783001,I783032,I783049,I783075,I783083,I783114,I783145,I783162,I783193,I783293,I783319,I783327,I783344,I783361,I783387,I783395,I783421,I783429,I783446,I783463,I783480,I783276,I783520,I783528,I783545,I783562,I783579,I783279,I783610,I783627,I783653,I783661,I783261,I783692,I783270,I783723,I783740,I783282,I783771,I783273,I783264,I783267,I783285,I783871,I1282857,I783897,I783905,I783922,I1282860,I1282869,I783939,I1282872,I783965,I783973,I1282881,I1282863,I783999,I784007,I784024,I784041,I784058,I784098,I784106,I784123,I784140,I784157,I784188,I1282878,I784205,I1282875,I784231,I784239,I784270,I784301,I784318,I784349,I1282866,I784449,I1064617,I784475,I784483,I784500,I1064614,I1064632,I784517,I1064629,I784543,I784551,I1064611,I784577,I784585,I784602,I784619,I784636,I784432,I1064623,I784676,I784684,I784701,I784718,I784735,I784435,I784766,I1064626,I784783,I784809,I784817,I784417,I784848,I784426,I784879,I784896,I784438,I784927,I1064620,I784429,I784420,I784423,I784441,I785027,I785053,I785061,I785078,I785095,I785121,I785129,I785155,I785163,I785180,I785197,I785214,I785010,I785254,I785262,I785279,I785296,I785313,I785013,I785344,I785361,I785387,I785395,I784995,I785426,I785004,I785457,I785474,I785016,I785505,I785007,I784998,I785001,I785019,I785605,I785631,I785639,I785656,I785673,I785699,I785707,I785733,I785741,I785758,I785775,I785792,I785832,I785840,I785857,I785874,I785891,I785922,I785939,I785965,I785973,I786004,I786035,I786052,I786083,I786183,I1073593,I786209,I786217,I786234,I1073590,I1073608,I786251,I1073605,I786277,I786285,I1073587,I786311,I786319,I786336,I786353,I786370,I1073599,I786410,I786418,I786435,I786452,I786469,I786500,I1073602,I786517,I786543,I786551,I786582,I786613,I786630,I786661,I1073596,I786761,I786787,I786795,I786812,I786829,I786855,I786863,I786889,I786897,I786914,I786931,I786948,I786744,I786988,I786996,I787013,I787030,I787047,I786747,I787078,I787095,I787121,I787129,I786729,I787160,I786738,I787191,I787208,I786750,I787239,I786741,I786732,I786735,I786753,I787339,I1230311,I787365,I787373,I787390,I1230293,I1230305,I787407,I1230308,I787433,I787441,I1230302,I1230299,I787467,I787475,I787492,I787509,I787526,I1230317,I787566,I787574,I787591,I787608,I787625,I787656,I1230296,I787673,I787699,I787707,I787738,I787769,I787786,I787817,I1230314,I787917,I1351785,I787943,I787951,I787968,I1351770,I1351758,I787985,I1351773,I788011,I788019,I1351776,I788045,I788053,I788070,I788087,I788104,I1351764,I788144,I788152,I788169,I788186,I788203,I788234,I1351761,I1351767,I788251,I1351782,I788277,I788285,I788316,I788347,I788364,I788395,I1351779,I788495,I788521,I788529,I788546,I788563,I788589,I788597,I788623,I788631,I788648,I788665,I788682,I788722,I788730,I788747,I788764,I788781,I788812,I788829,I788855,I788863,I788894,I788925,I788942,I788973,I789073,I789099,I789107,I789124,I789141,I789167,I789175,I789201,I789209,I789226,I789243,I789260,I789056,I789300,I789308,I789325,I789342,I789359,I789059,I789390,I789407,I789433,I789441,I789041,I789472,I789050,I789503,I789520,I789062,I789551,I789053,I789044,I789047,I789065,I789651,I789677,I789685,I789702,I789719,I789745,I789753,I789779,I789787,I789804,I789821,I789838,I789878,I789886,I789903,I789920,I789937,I789968,I789985,I790011,I790019,I790050,I790081,I790098,I790129,I790229,I790255,I790263,I790280,I790297,I790323,I790331,I790357,I790365,I790382,I790399,I790416,I790212,I790456,I790464,I790481,I790498,I790515,I790215,I790546,I790563,I790589,I790597,I790197,I790628,I790206,I790659,I790676,I790218,I790707,I790209,I790200,I790203,I790221,I790807,I790833,I790841,I790858,I790875,I790901,I790909,I790935,I790943,I790960,I790977,I790994,I790790,I791034,I791042,I791059,I791076,I791093,I790793,I791124,I791141,I791167,I791175,I790775,I791206,I790784,I791237,I791254,I790796,I791285,I790787,I790778,I790781,I790799,I791385,I791411,I791419,I791436,I791453,I791479,I791487,I791513,I791521,I791538,I791555,I791572,I791368,I791612,I791620,I791637,I791654,I791671,I791371,I791702,I791719,I791745,I791753,I791353,I791784,I791362,I791815,I791832,I791374,I791863,I791365,I791356,I791359,I791377,I791963,I791989,I791997,I792014,I792031,I792057,I792065,I792091,I792099,I792116,I792133,I792150,I791946,I792190,I792198,I792215,I792232,I792249,I791949,I792280,I792297,I792323,I792331,I791931,I792362,I791940,I792393,I792410,I791952,I792441,I791943,I791934,I791937,I791955,I792541,I1143611,I792567,I792575,I792592,I1143593,I1143605,I792609,I1143608,I792635,I792643,I1143602,I1143599,I792669,I792677,I792694,I792711,I792728,I792524,I1143617,I792768,I792776,I792793,I792810,I792827,I792527,I792858,I1143596,I792875,I792901,I792909,I792509,I792940,I792518,I792971,I792988,I792530,I793019,I1143614,I792521,I792512,I792515,I792533,I793119,I793145,I793153,I793170,I793187,I793213,I793221,I793247,I793255,I793272,I793289,I793306,I793346,I793354,I793371,I793388,I793405,I793436,I793453,I793479,I793487,I793518,I793549,I793566,I793597,I793697,I1189851,I793723,I793731,I793748,I1189833,I1189845,I793765,I1189848,I793791,I793799,I1189842,I1189839,I793825,I793833,I793850,I793867,I793884,I1189857,I793924,I793932,I793949,I793966,I793983,I794014,I1189836,I794031,I794057,I794065,I794096,I794127,I794144,I794175,I1189854,I794275,I1300469,I794301,I794309,I794326,I1300493,I1300475,I794343,I1300481,I794369,I794377,I1300487,I1300472,I794403,I794411,I794428,I794445,I794462,I1300484,I794502,I794510,I794527,I794544,I794561,I794592,I1300490,I1300478,I794609,I794635,I794643,I794674,I794705,I794722,I794753,I794853,I794879,I794887,I794904,I794921,I794947,I794955,I794981,I794989,I795006,I795023,I795040,I794836,I795080,I795088,I795105,I795122,I795139,I794839,I795170,I795187,I795213,I795221,I794821,I795252,I794830,I795283,I795300,I794842,I795331,I794833,I794824,I794827,I794845,I795431,I795457,I795465,I795482,I795499,I795525,I795533,I795559,I795567,I795584,I795601,I795618,I795414,I795658,I795666,I795683,I795700,I795717,I795417,I795748,I795765,I795791,I795799,I795399,I795830,I795408,I795861,I795878,I795420,I795909,I795411,I795402,I795405,I795423,I796009,I796035,I796043,I796060,I796077,I796103,I796111,I796137,I796145,I796162,I796179,I796196,I795992,I796236,I796244,I796261,I796278,I796295,I795995,I796326,I796343,I796369,I796377,I795977,I796408,I795986,I796439,I796456,I795998,I796487,I795989,I795980,I795983,I796001,I796587,I1174245,I796613,I796621,I796638,I1174227,I1174239,I796655,I1174242,I796681,I796689,I1174236,I1174233,I796715,I796723,I796740,I796757,I796774,I796570,I1174251,I796814,I796822,I796839,I796856,I796873,I796573,I796904,I1174230,I796921,I796947,I796955,I796555,I796986,I796564,I797017,I797034,I796576,I797065,I1174248,I796567,I796558,I796561,I796579,I797165,I797191,I797199,I797216,I797233,I797259,I797267,I797293,I797301,I797318,I797335,I797352,I797392,I797400,I797417,I797434,I797451,I797482,I797499,I797525,I797533,I797564,I797595,I797612,I797643,I797743,I1382725,I797769,I797777,I797794,I1382710,I1382698,I797811,I1382713,I797837,I797845,I1382716,I797871,I797879,I797896,I797913,I797930,I797726,I1382704,I797970,I797978,I797995,I798012,I798029,I797729,I798060,I1382701,I1382707,I798077,I1382722,I798103,I798111,I797711,I798142,I797720,I798173,I798190,I797732,I798221,I1382719,I797723,I797714,I797717,I797735,I798321,I798347,I798355,I798372,I798389,I798415,I798423,I798449,I798457,I798474,I798491,I798508,I798304,I798548,I798556,I798573,I798590,I798607,I798307,I798638,I798655,I798681,I798689,I798289,I798720,I798298,I798751,I798768,I798310,I798799,I798301,I798292,I798295,I798313,I798899,I861663,I798925,I798933,I798950,I861651,I861669,I798967,I861666,I798993,I799001,I861657,I861654,I799027,I799035,I799052,I799069,I799086,I861648,I799126,I799134,I799151,I799168,I799185,I799216,I799233,I799259,I799267,I799298,I799329,I799346,I799377,I861660,I799477,I799503,I799511,I799528,I799545,I799571,I799579,I799605,I799613,I799630,I799647,I799664,I799460,I799704,I799712,I799729,I799746,I799763,I799463,I799794,I799811,I799837,I799845,I799445,I799876,I799454,I799907,I799924,I799466,I799955,I799457,I799448,I799451,I799469,I800055,I800081,I800089,I800106,I800123,I800149,I800157,I800183,I800191,I800208,I800225,I800242,I800038,I800282,I800290,I800307,I800324,I800341,I800041,I800372,I800389,I800415,I800423,I800023,I800454,I800032,I800485,I800502,I800044,I800533,I800035,I800026,I800029,I800047,I800633,I923297,I800659,I800667,I800684,I923273,I923288,I800701,I923300,I800727,I800735,I923285,I923276,I800761,I800769,I800786,I800803,I800820,I800860,I800868,I800885,I800902,I800919,I800950,I923291,I923282,I800967,I923294,I800993,I801001,I801032,I801063,I801080,I801111,I923279,I801211,I801237,I801245,I801262,I801279,I801305,I801313,I801339,I801347,I801364,I801381,I801398,I801194,I801438,I801446,I801463,I801480,I801497,I801197,I801528,I801545,I801571,I801579,I801179,I801610,I801188,I801641,I801658,I801200,I801689,I801191,I801182,I801185,I801203,I801789,I801815,I801823,I801840,I801857,I801883,I801891,I801917,I801925,I801942,I801959,I801976,I802016,I802024,I802041,I802058,I802075,I802106,I802123,I802149,I802157,I802188,I802219,I802236,I802267,I802367,I802393,I802401,I802418,I802435,I802461,I802469,I802495,I802503,I802520,I802537,I802554,I802594,I802602,I802619,I802636,I802653,I802684,I802701,I802727,I802735,I802766,I802797,I802814,I802845,I802945,I950429,I802971,I802979,I802996,I950405,I950420,I803013,I950432,I803039,I803047,I950417,I950408,I803073,I803081,I803098,I803115,I803132,I802928,I803172,I803180,I803197,I803214,I803231,I802931,I803262,I950423,I950414,I803279,I950426,I803305,I803313,I802913,I803344,I802922,I803375,I803392,I802934,I803423,I950411,I802925,I802916,I802919,I802937,I803523,I970455,I803549,I803557,I803574,I970431,I970446,I803591,I970458,I803617,I803625,I970443,I970434,I803651,I803659,I803676,I803693,I803710,I803750,I803758,I803775,I803792,I803809,I803840,I970449,I970440,I803857,I970452,I803883,I803891,I803922,I803953,I803970,I804001,I970437,I804101,I804127,I804135,I804152,I804169,I804195,I804203,I804229,I804237,I804254,I804271,I804288,I804084,I804328,I804336,I804353,I804370,I804387,I804087,I804418,I804435,I804461,I804469,I804069,I804500,I804078,I804531,I804548,I804090,I804579,I804081,I804072,I804075,I804093,I804679,I804705,I804713,I804730,I804747,I804773,I804781,I804807,I804815,I804832,I804849,I804866,I804662,I804906,I804914,I804931,I804948,I804965,I804665,I804996,I805013,I805039,I805047,I804647,I805078,I804656,I805109,I805126,I804668,I805157,I804659,I804650,I804653,I804671,I805257,I805283,I805291,I805308,I805325,I805351,I805359,I805385,I805393,I805410,I805427,I805444,I805240,I805484,I805492,I805509,I805526,I805543,I805243,I805574,I805591,I805617,I805625,I805225,I805656,I805234,I805687,I805704,I805246,I805735,I805237,I805228,I805231,I805249,I805835,I993711,I805861,I805869,I805886,I993687,I993702,I805903,I993714,I805929,I805937,I993699,I993690,I805963,I805971,I805988,I806005,I806022,I806062,I806070,I806087,I806104,I806121,I806152,I993705,I993696,I806169,I993708,I806195,I806203,I806234,I806265,I806282,I806313,I993693,I806413,I935571,I806439,I806447,I806464,I935547,I935562,I806481,I935574,I806507,I806515,I935559,I935550,I806541,I806549,I806566,I806583,I806600,I806640,I806648,I806665,I806682,I806699,I806730,I935565,I935556,I806747,I935568,I806773,I806781,I806812,I806843,I806860,I806891,I935553,I806991,I807017,I807025,I807042,I807059,I807085,I807093,I807119,I807127,I807144,I807161,I807178,I807218,I807226,I807243,I807260,I807277,I807308,I807325,I807351,I807359,I807390,I807421,I807438,I807469,I807569,I807595,I807603,I807620,I807637,I807663,I807671,I807697,I807705,I807722,I807739,I807756,I807796,I807804,I807821,I807838,I807855,I807886,I807903,I807929,I807937,I807968,I807999,I808016,I808047,I808147,I808173,I808181,I808198,I808215,I808241,I808249,I808275,I808283,I808300,I808317,I808334,I808130,I808374,I808382,I808399,I808416,I808433,I808133,I808464,I808481,I808507,I808515,I808115,I808546,I808124,I808577,I808594,I808136,I808625,I808127,I808118,I808121,I808139,I808725,I1401765,I808751,I808759,I808776,I1401750,I1401738,I808793,I1401753,I808819,I808827,I1401756,I808853,I808861,I808878,I808895,I808912,I808708,I1401744,I808952,I808960,I808977,I808994,I809011,I808711,I809042,I1401741,I1401747,I809059,I1401762,I809085,I809093,I808693,I809124,I808702,I809155,I809172,I808714,I809203,I1401759,I808705,I808696,I808699,I808717,I809303,I1287753,I809329,I809337,I809354,I1287777,I1287759,I809371,I1287765,I809397,I809405,I1287771,I1287756,I809431,I809439,I809456,I809473,I809490,I1287768,I809530,I809538,I809555,I809572,I809589,I809620,I1287774,I1287762,I809637,I809663,I809671,I809702,I809733,I809750,I809781,I809881,I949137,I809907,I809915,I809932,I949113,I949128,I809949,I949140,I809975,I809983,I949125,I949116,I810009,I810017,I810034,I810051,I810068,I809864,I810108,I810116,I810133,I810150,I810167,I809867,I810198,I949131,I949122,I810215,I949134,I810241,I810249,I809849,I810280,I809858,I810311,I810328,I809870,I810359,I949119,I809861,I809852,I809855,I809873,I810459,I902242,I810485,I810493,I810510,I902230,I902248,I810527,I902245,I810553,I810561,I902236,I902233,I810587,I810595,I810612,I810629,I810646,I902227,I810686,I810694,I810711,I810728,I810745,I810776,I810793,I810819,I810827,I810858,I810889,I810906,I810937,I902239,I811037,I811063,I811071,I811088,I811105,I811131,I811139,I811165,I811173,I811190,I811207,I811224,I811264,I811272,I811289,I811306,I811323,I811354,I811371,I811397,I811405,I811436,I811467,I811484,I811515,I811612,I811638,I811646,I811663,I811680,I811706,I811737,I811745,I811762,I811788,I811796,I811836,I811872,I811889,I811915,I811923,I811940,I811971,I811988,I812005,I812036,I812067,I812084,I812139,I812165,I812173,I812190,I812207,I812233,I812264,I812272,I812289,I812315,I812323,I812363,I812399,I812416,I812442,I812450,I812467,I812498,I812515,I812532,I812563,I812594,I812611,I812666,I1083133,I812692,I812700,I812717,I1083142,I1083130,I812734,I1083127,I812760,I812655,I812791,I812799,I1083124,I812816,I812842,I812850,I812658,I812890,I812649,I812640,I812926,I1083145,I1083136,I812943,I1083139,I812969,I812977,I812994,I812643,I813025,I813042,I813059,I812652,I813090,I812637,I813121,I813138,I812646,I813193,I813219,I813227,I813244,I813261,I813287,I813318,I813326,I813343,I813369,I813377,I813417,I813453,I813470,I813496,I813504,I813521,I813552,I813569,I813586,I813617,I813648,I813665,I813720,I1134363,I813746,I813754,I813771,I1134345,I813788,I1134351,I813814,I813709,I1134348,I813845,I813853,I1134357,I813870,I813896,I813904,I813712,I1134369,I813944,I813703,I813694,I813980,I1134360,I1134354,I813997,I814023,I814031,I814048,I813697,I814079,I1134366,I814096,I814113,I813706,I814144,I813691,I814175,I814192,I813700,I814247,I814273,I814281,I814298,I814315,I814341,I814372,I814380,I814397,I814423,I814431,I814471,I814507,I814524,I814550,I814558,I814575,I814606,I814623,I814640,I814671,I814702,I814719,I814774,I814800,I814808,I814825,I814842,I814868,I814899,I814907,I814924,I814950,I814958,I814998,I815034,I815051,I815077,I815085,I815102,I815133,I815150,I815167,I815198,I815229,I815246,I815301,I815327,I815335,I815352,I815369,I815395,I815290,I815426,I815434,I815451,I815477,I815485,I815293,I815525,I815284,I815275,I815561,I815578,I815604,I815612,I815629,I815278,I815660,I815677,I815694,I815287,I815725,I815272,I815756,I815773,I815281,I815828,I1045370,I815854,I815862,I815879,I1045385,I1045367,I815896,I815922,I815817,I1045376,I815953,I815961,I1045394,I815978,I816004,I816012,I815820,I1045391,I816052,I815811,I815802,I816088,I1045388,I1045379,I816105,I1045373,I816131,I816139,I816156,I815805,I816187,I1045382,I816204,I816221,I815814,I816252,I815799,I816283,I816300,I815808,I816355,I816381,I816389,I816406,I816423,I816449,I816344,I816480,I816488,I816505,I816531,I816539,I816347,I816579,I816338,I816329,I816615,I816632,I816658,I816666,I816683,I816332,I816714,I816731,I816748,I816341,I816779,I816326,I816810,I816827,I816335,I816882,I816908,I816916,I816933,I816950,I816976,I817007,I817015,I817032,I817058,I817066,I817106,I817142,I817159,I817185,I817193,I817210,I817241,I817258,I817275,I817306,I817337,I817354,I817409,I1209503,I817435,I817443,I817460,I1209485,I817477,I1209491,I817503,I1209488,I817534,I817542,I1209497,I817559,I817585,I817593,I1209509,I817633,I817669,I1209500,I1209494,I817686,I817712,I817720,I817737,I817768,I1209506,I817785,I817802,I817833,I817864,I817881,I817936,I817962,I817970,I817987,I818004,I818030,I817925,I818061,I818069,I818086,I818112,I818120,I817928,I818160,I817919,I817910,I818196,I818213,I818239,I818247,I818264,I817913,I818295,I818312,I818329,I817922,I818360,I817907,I818391,I818408,I817916,I818463,I980124,I818489,I818497,I818514,I980139,I980121,I818531,I818557,I818452,I980130,I818588,I818596,I980148,I818613,I818639,I818647,I818455,I980145,I818687,I818446,I818437,I818723,I980142,I980133,I818740,I980127,I818766,I818774,I818791,I818440,I818822,I980136,I818839,I818856,I818449,I818887,I818434,I818918,I818935,I818443,I818990,I819016,I819024,I819041,I819058,I819084,I819115,I819123,I819140,I819166,I819174,I819214,I819250,I819267,I819293,I819301,I819318,I819349,I819366,I819383,I819414,I819445,I819462,I819517,I819543,I819551,I819568,I819585,I819611,I819642,I819650,I819667,I819693,I819701,I819741,I819777,I819794,I819820,I819828,I819845,I819876,I819893,I819910,I819941,I819972,I819989,I820044,I820070,I820078,I820095,I820112,I820138,I820169,I820177,I820194,I820220,I820228,I820268,I820304,I820321,I820347,I820355,I820372,I820403,I820420,I820437,I820468,I820499,I820516,I820571,I820597,I820605,I820622,I820639,I820665,I820696,I820704,I820721,I820747,I820755,I820795,I820831,I820848,I820874,I820882,I820899,I820930,I820947,I820964,I820995,I821026,I821043,I821098,I1264917,I821124,I821132,I821149,I1264923,I1264905,I821166,I1264914,I821192,I821087,I1264920,I821223,I821231,I1264908,I821248,I821274,I821282,I821090,I1264926,I821322,I821081,I821072,I821358,I1264911,I821375,I1264929,I821401,I821409,I821426,I821075,I821457,I821474,I821491,I821084,I821522,I821069,I821553,I821570,I821078,I821625,I821651,I821659,I821676,I821693,I821719,I821750,I821758,I821775,I821801,I821809,I821849,I821885,I821902,I821928,I821936,I821953,I821984,I822001,I822018,I822049,I822080,I822097,I822152,I1138987,I822178,I822186,I822203,I1138969,I822220,I1138975,I822246,I1138972,I822277,I822285,I1138981,I822302,I822328,I822336,I1138993,I822376,I822412,I1138984,I1138978,I822429,I822455,I822463,I822480,I822511,I1138990,I822528,I822545,I822576,I822607,I822624,I822679,I822705,I822713,I822730,I822747,I822773,I822668,I822804,I822812,I822829,I822855,I822863,I822671,I822903,I822662,I822653,I822939,I822956,I822982,I822990,I823007,I822656,I823038,I823055,I823072,I822665,I823103,I822650,I823134,I823151,I822659,I823206,I1094481,I823232,I823240,I823257,I1094463,I823274,I1094469,I823300,I1094466,I823331,I823339,I1094475,I823356,I823382,I823390,I1094487,I823430,I823466,I1094478,I1094472,I823483,I823509,I823517,I823534,I823565,I1094484,I823582,I823599,I823630,I823661,I823678,I823733,I823759,I823767,I823784,I823801,I823827,I823722,I823858,I823866,I823883,I823909,I823917,I823725,I823957,I823716,I823707,I823993,I824010,I824036,I824044,I824061,I823710,I824092,I824109,I824126,I823719,I824157,I823704,I824188,I824205,I823713,I824260,I824286,I824294,I824311,I824328,I824354,I824385,I824393,I824410,I824436,I824444,I824484,I824520,I824537,I824563,I824571,I824588,I824619,I824636,I824653,I824684,I824715,I824732,I824787,I824813,I824821,I824838,I824855,I824881,I824776,I824912,I824920,I824937,I824963,I824971,I824779,I825011,I824770,I824761,I825047,I825064,I825090,I825098,I825115,I824764,I825146,I825163,I825180,I824773,I825211,I824758,I825242,I825259,I824767,I825314,I825340,I825348,I825365,I825382,I825408,I825439,I825447,I825464,I825490,I825498,I825538,I825574,I825591,I825617,I825625,I825642,I825673,I825690,I825707,I825738,I825769,I825786,I825841,I825867,I825875,I825892,I825909,I825935,I825966,I825974,I825991,I826017,I826025,I826065,I826101,I826118,I826144,I826152,I826169,I826200,I826217,I826234,I826265,I826296,I826313,I826368,I826394,I826402,I826419,I826436,I826462,I826493,I826501,I826518,I826544,I826552,I826592,I826628,I826645,I826671,I826679,I826696,I826727,I826744,I826761,I826792,I826823,I826840,I826895,I963328,I826921,I826929,I826946,I963343,I963325,I826963,I826989,I963334,I827020,I827028,I963352,I827045,I827071,I827079,I963349,I827119,I827155,I963346,I963337,I827172,I963331,I827198,I827206,I827223,I827254,I963340,I827271,I827288,I827319,I827350,I827367,I827422,I1405323,I827448,I827456,I827473,I1405320,I1405329,I827490,I1405308,I827516,I1405311,I827547,I827555,I1405326,I827572,I827598,I827606,I1405332,I827646,I827682,I1405314,I1405335,I827699,I1405317,I827725,I827733,I827750,I827781,I827798,I827815,I827846,I827877,I827894,I827949,I1211815,I827975,I827983,I828000,I1211797,I828017,I1211803,I828043,I827938,I1211800,I828074,I828082,I1211809,I828099,I828125,I828133,I827941,I1211821,I828173,I827932,I827923,I828209,I1211812,I1211806,I828226,I828252,I828260,I828277,I827926,I828308,I1211818,I828325,I828342,I827935,I828373,I827920,I828404,I828421,I827929,I828476,I828502,I828510,I828527,I828544,I828570,I828465,I828601,I828609,I828626,I828652,I828660,I828468,I828700,I828459,I828450,I828736,I828753,I828779,I828787,I828804,I828453,I828835,I828852,I828869,I828462,I828900,I828447,I828931,I828948,I828456,I829003,I1305111,I829029,I829037,I829054,I1305093,I1305096,I829071,I1305108,I829097,I828992,I1305117,I829128,I829136,I1305102,I829153,I829179,I829187,I828995,I1305114,I829227,I828986,I828977,I829263,I1305105,I1305099,I829280,I829306,I829314,I829331,I828980,I829362,I829379,I829396,I828989,I829427,I828974,I829458,I829475,I828983,I829530,I829556,I829564,I829581,I829598,I829624,I829655,I829663,I829680,I829706,I829714,I829754,I829790,I829807,I829833,I829841,I829858,I829889,I829906,I829923,I829954,I829985,I830002,I830057,I830083,I830091,I830108,I830125,I830151,I830046,I830182,I830190,I830207,I830233,I830241,I830049,I830281,I830040,I830031,I830317,I830334,I830360,I830368,I830385,I830034,I830416,I830433,I830450,I830043,I830481,I830028,I830512,I830529,I830037,I830584,I830610,I830618,I830635,I830652,I830678,I830573,I830709,I830717,I830734,I830760,I830768,I830576,I830808,I830567,I830558,I830844,I830861,I830887,I830895,I830912,I830561,I830943,I830960,I830977,I830570,I831008,I830555,I831039,I831056,I830564,I831111,I1104307,I831137,I831145,I831162,I1104289,I831179,I1104295,I831205,I1104292,I831236,I831244,I1104301,I831261,I831287,I831295,I1104313,I831335,I831371,I1104304,I1104298,I831388,I831414,I831422,I831439,I831470,I1104310,I831487,I831504,I831535,I831566,I831583,I831638,I943948,I831664,I831672,I831689,I943963,I943945,I831706,I831732,I943954,I831763,I831771,I943972,I831788,I831814,I831822,I943969,I831862,I831898,I943966,I943957,I831915,I943951,I831941,I831949,I831966,I831997,I943960,I832014,I832031,I832062,I832093,I832110,I832165,I832191,I832199,I832216,I832233,I832259,I832290,I832298,I832315,I832341,I832349,I832389,I832425,I832442,I832468,I832476,I832493,I832524,I832541,I832558,I832589,I832620,I832637,I832692,I832718,I832726,I832743,I832760,I832786,I832817,I832825,I832842,I832868,I832876,I832916,I832952,I832969,I832995,I833003,I833020,I833051,I833068,I833085,I833116,I833147,I833164,I833219,I1167309,I833245,I833253,I833270,I1167291,I833287,I1167297,I833313,I1167294,I833344,I833352,I1167303,I833369,I833395,I833403,I1167315,I833443,I833479,I1167306,I1167300,I833496,I833522,I833530,I833547,I833578,I1167312,I833595,I833612,I833643,I833674,I833691,I833746,I833772,I833780,I833797,I833814,I833840,I833871,I833879,I833896,I833922,I833930,I833970,I834006,I834023,I834049,I834057,I834074,I834105,I834122,I834139,I834170,I834201,I834218,I834273,I1269813,I834299,I834307,I834324,I1269819,I1269801,I834341,I1269810,I834367,I1269816,I834398,I834406,I1269804,I834423,I834449,I834457,I1269822,I834497,I834533,I1269807,I834550,I1269825,I834576,I834584,I834601,I834632,I834649,I834666,I834697,I834728,I834745,I834800,I1009194,I834826,I834834,I834851,I1009209,I1009191,I834868,I834894,I1009200,I834925,I834933,I1009218,I834950,I834976,I834984,I1009215,I835024,I835060,I1009212,I1009203,I835077,I1009197,I835103,I835111,I835128,I835159,I1009206,I835176,I835193,I835224,I835255,I835272,I835327,I1019530,I835353,I835361,I835378,I1019545,I1019527,I835395,I835421,I1019536,I835452,I835460,I1019554,I835477,I835503,I835511,I1019551,I835551,I835587,I1019548,I1019539,I835604,I1019533,I835630,I835638,I835655,I835686,I1019542,I835703,I835720,I835751,I835782,I835799,I835854,I835880,I835888,I835905,I835922,I835948,I835979,I835987,I836004,I836030,I836038,I836078,I836114,I836131,I836157,I836165,I836182,I836213,I836230,I836247,I836278,I836309,I836326,I836381,I836407,I836415,I836432,I836449,I836475,I836506,I836514,I836531,I836557,I836565,I836605,I836641,I836658,I836684,I836692,I836709,I836740,I836757,I836774,I836805,I836836,I836853,I836908,I836934,I836942,I836959,I836976,I837002,I837033,I837041,I837058,I837084,I837092,I837132,I837168,I837185,I837211,I837219,I837236,I837267,I837284,I837301,I837332,I837363,I837380,I837435,I1171355,I837461,I837469,I837486,I1171337,I837503,I1171343,I837529,I1171340,I837560,I837568,I1171349,I837585,I837611,I837619,I1171361,I837659,I837695,I1171352,I1171346,I837712,I837738,I837746,I837763,I837794,I1171358,I837811,I837828,I837859,I837890,I837907,I837962,I1396398,I837988,I837996,I838013,I1396395,I1396404,I838030,I1396383,I838056,I1396386,I838087,I838095,I1396401,I838112,I838138,I838146,I1396407,I838186,I838222,I1396389,I1396410,I838239,I1396392,I838265,I838273,I838290,I838321,I838338,I838355,I838386,I838417,I838434,I838489,I838515,I838523,I838540,I838557,I838583,I838614,I838622,I838639,I838665,I838673,I838713,I838749,I838766,I838792,I838800,I838817,I838848,I838865,I838882,I838913,I838944,I838961,I839016,I839042,I839050,I839067,I839084,I839110,I839005,I839141,I839149,I839166,I839192,I839200,I839008,I839240,I838999,I838990,I839276,I839293,I839319,I839327,I839344,I838993,I839375,I839392,I839409,I839002,I839440,I838987,I839471,I839488,I838996,I839543,I839569,I839577,I839594,I839611,I839637,I839532,I839668,I839676,I839693,I839719,I839727,I839535,I839767,I839526,I839517,I839803,I839820,I839846,I839854,I839871,I839520,I839902,I839919,I839936,I839529,I839967,I839514,I839998,I840015,I839523,I840070,I840096,I840104,I840121,I840138,I840164,I840195,I840203,I840220,I840246,I840254,I840294,I840330,I840347,I840373,I840381,I840398,I840429,I840446,I840463,I840494,I840525,I840542,I840597,I1048912,I840623,I840631,I840648,I1048921,I1048909,I840665,I1048906,I840691,I840586,I840722,I840730,I1048903,I840747,I840773,I840781,I840589,I840821,I840580,I840571,I840857,I1048924,I1048915,I840874,I1048918,I840900,I840908,I840925,I840574,I840956,I840973,I840990,I840583,I841021,I840568,I841052,I841069,I840577,I841124,I841150,I841158,I841175,I841192,I841218,I841249,I841257,I841274,I841300,I841308,I841348,I841384,I841401,I841427,I841435,I841452,I841483,I841500,I841517,I841548,I841579,I841596,I841651,I1318983,I841677,I841685,I841702,I1318965,I1318968,I841719,I1318980,I841745,I841640,I1318989,I841776,I841784,I1318974,I841801,I841827,I841835,I841643,I1318986,I841875,I841634,I841625,I841911,I1318977,I1318971,I841928,I841954,I841962,I841979,I841628,I842010,I842027,I842044,I841637,I842075,I841622,I842106,I842123,I841631,I842178,I922630,I842204,I842212,I842229,I922645,I922627,I842246,I842272,I922636,I842303,I842311,I922654,I842328,I842354,I842362,I922651,I842402,I842438,I922648,I922639,I842455,I922633,I842481,I842489,I842506,I842537,I922642,I842554,I842571,I842602,I842633,I842650,I842705,I842731,I842739,I842756,I842773,I842799,I842694,I842830,I842838,I842855,I842881,I842889,I842697,I842929,I842688,I842679,I842965,I842982,I843008,I843016,I843033,I842682,I843064,I843081,I843098,I842691,I843129,I842676,I843160,I843177,I842685,I843232,I1076962,I843258,I843266,I843283,I1076971,I1076959,I843300,I1076956,I843326,I843221,I843357,I843365,I1076953,I843382,I843408,I843416,I843224,I843456,I843215,I843206,I843492,I1076974,I1076965,I843509,I1076968,I843535,I843543,I843560,I843209,I843591,I843608,I843625,I843218,I843656,I843203,I843687,I843704,I843212,I843759,I843785,I843793,I843810,I843827,I843853,I843884,I843892,I843909,I843935,I843943,I843983,I844019,I844036,I844062,I844070,I844087,I844118,I844135,I844152,I844183,I844214,I844231,I844286,I844312,I844320,I844337,I844354,I844380,I844411,I844419,I844436,I844462,I844470,I844510,I844546,I844563,I844589,I844597,I844614,I844645,I844662,I844679,I844710,I844741,I844758,I844813,I844839,I844847,I844864,I844881,I844907,I844938,I844946,I844963,I844989,I844997,I845037,I845073,I845090,I845116,I845124,I845141,I845172,I845189,I845206,I845237,I845268,I845285,I845340,I845366,I845374,I845391,I845408,I845434,I845465,I845473,I845490,I845516,I845524,I845564,I845600,I845617,I845643,I845651,I845668,I845699,I845716,I845733,I845764,I845795,I845812,I845867,I845893,I845901,I845918,I845935,I845961,I845856,I845992,I846000,I846017,I846043,I846051,I845859,I846091,I845850,I845841,I846127,I846144,I846170,I846178,I846195,I845844,I846226,I846243,I846260,I845853,I846291,I845838,I846322,I846339,I845847,I846394,I846420,I846428,I846445,I846462,I846488,I846519,I846527,I846544,I846570,I846578,I846618,I846654,I846671,I846697,I846705,I846722,I846753,I846770,I846787,I846818,I846849,I846866,I846921,I1217017,I846947,I846955,I846972,I1216999,I846989,I1217005,I847015,I846910,I1217002,I847046,I847054,I1217011,I847071,I847097,I847105,I846913,I1217023,I847145,I846904,I846895,I847181,I1217014,I1217008,I847198,I847224,I847232,I847249,I846898,I847280,I1217020,I847297,I847314,I846907,I847345,I846892,I847376,I847393,I846901,I847448,I847474,I847482,I847499,I847516,I847542,I847573,I847581,I847598,I847624,I847632,I847672,I847708,I847725,I847751,I847759,I847776,I847807,I847824,I847841,I847872,I847903,I847920,I847975,I848001,I848009,I848026,I848043,I848069,I848100,I848108,I848125,I848151,I848159,I848199,I848235,I848252,I848278,I848286,I848303,I848334,I848351,I848368,I848399,I848430,I848447,I848502,I976248,I848528,I848536,I848553,I976263,I976245,I848570,I848596,I848491,I976254,I848627,I848635,I976272,I848652,I848678,I848686,I848494,I976269,I848726,I848485,I848476,I848762,I976266,I976257,I848779,I976251,I848805,I848813,I848830,I848479,I848861,I976260,I848878,I848895,I848488,I848926,I848473,I848957,I848974,I848482,I849029,I849055,I849063,I849080,I849097,I849123,I849154,I849162,I849179,I849205,I849213,I849253,I849289,I849306,I849332,I849340,I849357,I849388,I849405,I849422,I849453,I849484,I849501,I849556,I849582,I849590,I849607,I849624,I849650,I849545,I849681,I849689,I849706,I849732,I849740,I849548,I849780,I849539,I849530,I849816,I849833,I849859,I849867,I849884,I849533,I849915,I849932,I849949,I849542,I849980,I849527,I850011,I850028,I849536,I850083,I1303377,I850109,I850117,I850134,I1303359,I1303362,I850151,I1303374,I850177,I850072,I1303383,I850208,I850216,I1303368,I850233,I850259,I850267,I850075,I1303380,I850307,I850066,I850057,I850343,I1303371,I1303365,I850360,I850386,I850394,I850411,I850060,I850442,I850459,I850476,I850069,I850507,I850054,I850538,I850555,I850063,I850610,I1314937,I850636,I850644,I850661,I1314919,I1314922,I850678,I1314934,I850704,I850599,I1314943,I850735,I850743,I1314928,I850760,I850786,I850794,I850602,I1314940,I850834,I850593,I850584,I850870,I1314931,I1314925,I850887,I850913,I850921,I850938,I850587,I850969,I850986,I851003,I850596,I851034,I850581,I851065,I851082,I850590,I851137,I851163,I851171,I851188,I851205,I851231,I851126,I851262,I851270,I851287,I851313,I851321,I851129,I851361,I851120,I851111,I851397,I851414,I851440,I851448,I851465,I851114,I851496,I851513,I851530,I851123,I851561,I851108,I851592,I851609,I851117,I851664,I1222797,I851690,I851698,I851715,I1222779,I851732,I1222785,I851758,I1222782,I851789,I851797,I1222791,I851814,I851840,I851848,I1222803,I851888,I851924,I1222794,I1222788,I851941,I851967,I851975,I851992,I852023,I1222800,I852040,I852057,I852088,I852119,I852136,I852191,I852217,I852225,I852242,I852259,I852285,I852180,I852316,I852324,I852341,I852367,I852375,I852183,I852415,I852174,I852165,I852451,I852468,I852494,I852502,I852519,I852168,I852550,I852567,I852584,I852177,I852615,I852162,I852646,I852663,I852171,I852718,I1148235,I852744,I852752,I852769,I1148217,I852786,I1148223,I852812,I1148220,I852843,I852851,I1148229,I852868,I852894,I852902,I1148241,I852942,I852978,I1148232,I1148226,I852995,I853021,I853029,I853046,I853077,I1148238,I853094,I853111,I853142,I853173,I853190,I853245,I853271,I853279,I853296,I853313,I853339,I853370,I853378,I853395,I853421,I853429,I853469,I853505,I853522,I853548,I853556,I853573,I853604,I853621,I853638,I853669,I853700,I853717,I853772,I853798,I853806,I853823,I853840,I853866,I853761,I853897,I853905,I853922,I853948,I853956,I853764,I853996,I853755,I853746,I854032,I854049,I854075,I854083,I854100,I853749,I854131,I854148,I854165,I853758,I854196,I853743,I854227,I854244,I853752,I854299,I1399373,I854325,I854333,I854350,I1399370,I1399379,I854367,I1399358,I854393,I1399361,I854424,I854432,I1399376,I854449,I854475,I854483,I1399382,I854523,I854559,I1399364,I1399385,I854576,I1399367,I854602,I854610,I854627,I854658,I854675,I854692,I854723,I854754,I854771,I854826,I854852,I854860,I854877,I854894,I854920,I854951,I854959,I854976,I855002,I855010,I855050,I855086,I855103,I855129,I855137,I855154,I855185,I855202,I855219,I855250,I855281,I855298,I855353,I1024052,I855379,I855387,I855404,I1024067,I1024049,I855421,I855447,I855342,I1024058,I855478,I855486,I1024076,I855503,I855529,I855537,I855345,I1024073,I855577,I855336,I855327,I855613,I1024070,I1024061,I855630,I1024055,I855656,I855664,I855681,I855330,I855712,I1024064,I855729,I855746,I855339,I855777,I855324,I855808,I855825,I855333,I855880,I855906,I855914,I855931,I855948,I855974,I855869,I856005,I856013,I856030,I856056,I856064,I855872,I856104,I855863,I855854,I856140,I856157,I856183,I856191,I856208,I855857,I856239,I856256,I856273,I855866,I856304,I855851,I856335,I856352,I855860,I856407,I856433,I856441,I856458,I856475,I856501,I856532,I856540,I856557,I856583,I856591,I856631,I856667,I856684,I856710,I856718,I856735,I856766,I856783,I856800,I856831,I856862,I856879,I856934,I856960,I856968,I856985,I857002,I857028,I857059,I857067,I857084,I857110,I857118,I857158,I857194,I857211,I857237,I857245,I857262,I857293,I857310,I857327,I857358,I857389,I857406,I857461,I1085938,I857487,I857495,I857512,I1085947,I1085935,I857529,I1085932,I857555,I857586,I857594,I1085929,I857611,I857637,I857645,I857685,I857721,I1085950,I1085941,I857738,I1085944,I857764,I857772,I857789,I857820,I857837,I857854,I857885,I857916,I857933,I857988,I858014,I858022,I858039,I858056,I858082,I857977,I858113,I858121,I858138,I858164,I858172,I857980,I858212,I857971,I857962,I858248,I858265,I858291,I858299,I858316,I857965,I858347,I858364,I858381,I857974,I858412,I857959,I858443,I858460,I857968,I858515,I858541,I858549,I858566,I858583,I858609,I858640,I858648,I858665,I858691,I858699,I858739,I858775,I858792,I858818,I858826,I858843,I858874,I858891,I858908,I858939,I858970,I858987,I859042,I919400,I859068,I859076,I859093,I919415,I919397,I859110,I859136,I859031,I919406,I859167,I859175,I919424,I859192,I859218,I859226,I859034,I919421,I859266,I859025,I859016,I859302,I919418,I919409,I859319,I919403,I859345,I859353,I859370,I859019,I859401,I919412,I859418,I859435,I859028,I859466,I859013,I859497,I859514,I859022,I859569,I1104885,I859595,I859603,I859620,I1104867,I859637,I1104873,I859663,I1104870,I859694,I859702,I1104879,I859719,I859745,I859753,I1104891,I859793,I859829,I1104882,I1104876,I859846,I859872,I859880,I859897,I859928,I1104888,I859945,I859962,I859993,I860024,I860041,I860096,I860122,I860130,I860147,I860164,I860190,I860221,I860229,I860246,I860272,I860280,I860320,I860356,I860373,I860399,I860407,I860424,I860455,I860472,I860489,I860520,I860551,I860568,I860623,I860649,I860657,I860674,I860691,I860717,I860612,I860748,I860756,I860773,I860799,I860807,I860615,I860847,I860606,I860597,I860883,I860900,I860926,I860934,I860951,I860600,I860982,I860999,I861016,I860609,I861047,I860594,I861078,I861095,I860603,I861150,I861176,I861184,I861201,I861218,I861244,I861275,I861283,I861300,I861326,I861334,I861374,I861410,I861427,I861453,I861461,I861478,I861509,I861526,I861543,I861574,I861605,I861622,I861677,I976894,I861703,I861711,I861728,I976909,I976891,I861745,I861771,I976900,I861802,I861810,I976918,I861827,I861853,I861861,I976915,I861901,I861937,I976912,I976903,I861954,I976897,I861980,I861988,I862005,I862036,I976906,I862053,I862070,I862101,I862132,I862149,I862204,I862230,I862238,I862255,I862272,I862298,I862329,I862337,I862354,I862380,I862388,I862428,I862464,I862481,I862507,I862515,I862532,I862563,I862580,I862597,I862628,I862659,I862676,I862731,I1165575,I862757,I862765,I862782,I1165557,I862799,I1165563,I862825,I1165560,I862856,I862864,I1165569,I862881,I862907,I862915,I1165581,I862955,I862991,I1165572,I1165566,I863008,I863034,I863042,I863059,I863090,I1165578,I863107,I863124,I863155,I863186,I863203,I863258,I1197943,I863284,I863292,I863309,I1197925,I863326,I1197931,I863352,I1197928,I863383,I863391,I1197937,I863408,I863434,I863442,I1197949,I863482,I863518,I1197940,I1197934,I863535,I863561,I863569,I863586,I863617,I1197946,I863634,I863651,I863682,I863713,I863730,I863785,I863811,I863819,I863836,I863853,I863879,I863910,I863918,I863935,I863961,I863969,I864009,I864045,I864062,I864088,I864096,I864113,I864144,I864161,I864178,I864209,I864240,I864257,I864312,I1067425,I864338,I864346,I864363,I1067434,I1067422,I864380,I1067419,I864406,I864437,I864445,I1067416,I864462,I864488,I864496,I864536,I864572,I1067437,I1067428,I864589,I1067431,I864615,I864623,I864640,I864671,I864688,I864705,I864736,I864767,I864784,I864839,I864865,I864873,I864890,I864907,I864933,I864828,I864964,I864972,I864989,I865015,I865023,I864831,I865063,I864822,I864813,I865099,I865116,I865142,I865150,I865167,I864816,I865198,I865215,I865232,I864825,I865263,I864810,I865294,I865311,I864819,I865366,I1095637,I865392,I865400,I865417,I1095619,I865434,I1095625,I865460,I1095622,I865491,I865499,I1095631,I865516,I865542,I865550,I1095643,I865590,I865626,I1095634,I1095628,I865643,I865669,I865677,I865694,I865725,I1095640,I865742,I865759,I865790,I865821,I865838,I865893,I1004672,I865919,I865927,I865944,I1004687,I1004669,I865961,I865987,I1004678,I866018,I866026,I1004696,I866043,I866069,I866077,I1004693,I866117,I866153,I1004690,I1004681,I866170,I1004675,I866196,I866204,I866221,I866252,I1004684,I866269,I866286,I866317,I866348,I866365,I866420,I943302,I866446,I866454,I866471,I943317,I943299,I866488,I866514,I943308,I866545,I866553,I943326,I866570,I866596,I866604,I943323,I866644,I866680,I943320,I943311,I866697,I943305,I866723,I866731,I866748,I866779,I943314,I866796,I866813,I866844,I866875,I866892,I866947,I866973,I866981,I866998,I867015,I867041,I867072,I867080,I867097,I867123,I867131,I867171,I867207,I867224,I867250,I867258,I867275,I867306,I867323,I867340,I867371,I867402,I867419,I867474,I1339873,I867500,I867508,I867525,I1339870,I1339879,I867542,I1339858,I867568,I867463,I1339861,I867599,I867607,I1339876,I867624,I867650,I867658,I867466,I1339882,I867698,I867457,I867448,I867734,I1339864,I1339885,I867751,I1339867,I867777,I867785,I867802,I867451,I867833,I867850,I867867,I867460,I867898,I867445,I867929,I867946,I867454,I868001,I1331543,I868027,I868035,I868052,I1331540,I1331549,I868069,I1331528,I868095,I1331531,I868126,I868134,I1331546,I868151,I868177,I868185,I1331552,I868225,I868261,I1331534,I1331555,I868278,I1331537,I868304,I868312,I868329,I868360,I868377,I868394,I868425,I868456,I868473,I868528,I1203145,I868554,I868562,I868579,I1203127,I868596,I1203133,I868622,I1203130,I868653,I868661,I1203139,I868678,I868704,I868712,I1203151,I868752,I868788,I1203142,I1203136,I868805,I868831,I868839,I868856,I868887,I1203148,I868904,I868921,I868952,I868983,I869000,I869055,I869081,I869089,I869106,I869123,I869149,I869180,I869188,I869205,I869231,I869239,I869279,I869315,I869332,I869358,I869366,I869383,I869414,I869431,I869448,I869479,I869510,I869527,I869582,I869608,I869616,I869633,I869650,I869676,I869571,I869707,I869715,I869732,I869758,I869766,I869574,I869806,I869565,I869556,I869842,I869859,I869885,I869893,I869910,I869559,I869941,I869958,I869975,I869568,I870006,I869553,I870037,I870054,I869562,I870109,I870135,I870143,I870160,I870177,I870203,I870098,I870234,I870242,I870259,I870285,I870293,I870101,I870333,I870092,I870083,I870369,I870386,I870412,I870420,I870437,I870086,I870468,I870485,I870502,I870095,I870533,I870080,I870564,I870581,I870089,I870636,I1205457,I870662,I870670,I870687,I1205439,I870704,I1205445,I870730,I1205442,I870761,I870769,I1205451,I870786,I870812,I870820,I1205463,I870860,I870896,I1205454,I1205448,I870913,I870939,I870947,I870964,I870995,I1205460,I871012,I871029,I871060,I871091,I871108,I871163,I871189,I871197,I871214,I871231,I871257,I871288,I871296,I871313,I871339,I871347,I871387,I871423,I871440,I871466,I871474,I871491,I871522,I871539,I871556,I871587,I871618,I871635,I871690,I871716,I871724,I871741,I871758,I871784,I871679,I871815,I871823,I871840,I871866,I871874,I871682,I871914,I871673,I871664,I871950,I871967,I871993,I872001,I872018,I871667,I872049,I872066,I872083,I871676,I872114,I871661,I872145,I872162,I871670,I872217,I1221063,I872243,I872251,I872268,I1221045,I872285,I1221051,I872311,I1221048,I872342,I872350,I1221057,I872367,I872393,I872401,I1221069,I872441,I872477,I1221060,I1221054,I872494,I872520,I872528,I872545,I872576,I1221066,I872593,I872610,I872641,I872672,I872689,I872744,I872770,I872778,I872795,I872812,I872838,I872869,I872877,I872894,I872920,I872928,I872968,I873004,I873021,I873047,I873055,I873072,I873103,I873120,I873137,I873168,I873199,I873216,I873271,I873297,I873305,I873322,I873339,I873365,I873260,I873396,I873404,I873421,I873447,I873455,I873263,I873495,I873254,I873245,I873531,I873548,I873574,I873582,I873599,I873248,I873630,I873647,I873664,I873257,I873695,I873242,I873726,I873743,I873251,I873798,I873824,I873832,I873849,I873866,I873892,I873923,I873931,I873948,I873974,I873982,I874022,I874058,I874075,I874101,I874109,I874126,I874157,I874174,I874191,I874222,I874253,I874270,I874325,I874351,I874359,I874376,I874393,I874419,I874450,I874458,I874475,I874501,I874509,I874549,I874585,I874602,I874628,I874636,I874653,I874684,I874701,I874718,I874749,I874780,I874797,I874852,I874878,I874886,I874903,I874920,I874946,I874841,I874977,I874985,I875002,I875028,I875036,I874844,I875076,I874835,I874826,I875112,I875129,I875155,I875163,I875180,I874829,I875211,I875228,I875245,I874838,I875276,I874823,I875307,I875324,I874832,I875379,I925860,I875405,I875413,I875430,I925875,I925857,I875447,I875473,I875368,I925866,I875504,I875512,I925884,I875529,I875555,I875563,I875371,I925881,I875603,I875362,I875353,I875639,I925878,I925869,I875656,I925863,I875682,I875690,I875707,I875356,I875738,I925872,I875755,I875772,I875365,I875803,I875350,I875834,I875851,I875359,I875906,I875932,I875940,I875957,I875974,I876000,I876031,I876039,I876056,I876082,I876090,I876130,I876166,I876183,I876209,I876217,I876234,I876265,I876282,I876299,I876330,I876361,I876378,I876433,I1167887,I876459,I876467,I876484,I1167869,I876501,I1167875,I876527,I1167872,I876558,I876566,I1167881,I876583,I876609,I876617,I1167893,I876657,I876693,I1167884,I1167878,I876710,I876736,I876744,I876761,I876792,I1167890,I876809,I876826,I876857,I876888,I876905,I876960,I876986,I876994,I877011,I877028,I877054,I877085,I877093,I877110,I877136,I877144,I877184,I877220,I877237,I877263,I877271,I877288,I877319,I877336,I877353,I877384,I877415,I877432,I877487,I877513,I877521,I877538,I877555,I877581,I877476,I877612,I877620,I877637,I877663,I877671,I877479,I877711,I877470,I877461,I877747,I877764,I877790,I877798,I877815,I877464,I877846,I877863,I877880,I877473,I877911,I877458,I877942,I877959,I877467,I878014,I1118757,I878040,I878048,I878065,I1118739,I878082,I1118745,I878108,I1118742,I878139,I878147,I1118751,I878164,I878190,I878198,I1118763,I878238,I878274,I1118754,I1118748,I878291,I878317,I878325,I878342,I878373,I1118760,I878390,I878407,I878438,I878469,I878486,I878541,I878567,I878575,I878592,I878609,I878635,I878530,I878666,I878674,I878691,I878717,I878725,I878533,I878765,I878524,I878515,I878801,I878818,I878844,I878852,I878869,I878518,I878900,I878917,I878934,I878527,I878965,I878512,I878996,I879013,I878521,I879068,I879094,I879102,I879119,I879136,I879162,I879193,I879201,I879218,I879244,I879252,I879292,I879328,I879345,I879371,I879379,I879396,I879427,I879444,I879461,I879492,I879523,I879540,I879595,I879621,I879629,I879646,I879663,I879689,I879584,I879720,I879728,I879745,I879771,I879779,I879587,I879819,I879578,I879569,I879855,I879872,I879898,I879906,I879923,I879572,I879954,I879971,I879988,I879581,I880019,I879566,I880050,I880067,I879575,I880122,I1115289,I880148,I880156,I880173,I1115271,I880190,I1115277,I880216,I1115274,I880247,I880255,I1115283,I880272,I880298,I880306,I1115295,I880346,I880382,I1115286,I1115280,I880399,I880425,I880433,I880450,I880481,I1115292,I880498,I880515,I880546,I880577,I880594,I880649,I880675,I880683,I880700,I880717,I880743,I880774,I880782,I880799,I880825,I880833,I880873,I880909,I880926,I880952,I880960,I880977,I881008,I881025,I881042,I881073,I881104,I881121,I881176,I881202,I881210,I881227,I881244,I881270,I881165,I881301,I881309,I881326,I881352,I881360,I881168,I881400,I881159,I881150,I881436,I881453,I881479,I881487,I881504,I881153,I881535,I881552,I881569,I881162,I881600,I881147,I881631,I881648,I881156,I881703,I881729,I881737,I881754,I881771,I881797,I881828,I881836,I881853,I881879,I881887,I881927,I881963,I881980,I882006,I882014,I882031,I882062,I882079,I882096,I882127,I882158,I882175,I882230,I882256,I882264,I882281,I882298,I882324,I882355,I882363,I882380,I882406,I882414,I882454,I882490,I882507,I882533,I882541,I882558,I882589,I882606,I882623,I882654,I882685,I882702,I882757,I882783,I882791,I882808,I882825,I882851,I882746,I882882,I882890,I882907,I882933,I882941,I882749,I882981,I882740,I882731,I883017,I883034,I883060,I883068,I883085,I882734,I883116,I883133,I883150,I882743,I883181,I882728,I883212,I883229,I882737,I883284,I1299331,I883310,I883318,I883335,I1299313,I1299316,I883352,I1299328,I883378,I1299337,I883409,I883417,I1299322,I883434,I883460,I883468,I1299334,I883508,I883544,I1299325,I1299319,I883561,I883587,I883595,I883612,I883643,I883660,I883677,I883708,I883739,I883756,I883811,I883837,I883845,I883862,I883879,I883905,I883936,I883944,I883961,I883987,I883995,I884035,I884071,I884088,I884114,I884122,I884139,I884170,I884187,I884204,I884235,I884266,I884283,I884338,I884364,I884372,I884389,I884406,I884432,I884463,I884471,I884488,I884514,I884522,I884562,I884598,I884615,I884641,I884649,I884666,I884697,I884714,I884731,I884762,I884793,I884810,I884865,I884891,I884899,I884916,I884933,I884959,I884854,I884990,I884998,I885015,I885041,I885049,I884857,I885089,I884848,I884839,I885125,I885142,I885168,I885176,I885193,I884842,I885224,I885241,I885258,I884851,I885289,I884836,I885320,I885337,I884845,I885392,I885418,I885426,I885443,I885460,I885486,I885381,I885517,I885525,I885542,I885568,I885576,I885384,I885616,I885375,I885366,I885652,I885669,I885695,I885703,I885720,I885369,I885751,I885768,I885785,I885378,I885816,I885363,I885847,I885864,I885372,I885919,I885945,I885953,I885970,I885987,I886013,I886044,I886052,I886069,I886095,I886103,I886143,I886179,I886196,I886222,I886230,I886247,I886278,I886295,I886312,I886343,I886374,I886391,I886446,I886472,I886480,I886497,I886514,I886540,I886571,I886579,I886596,I886622,I886630,I886670,I886706,I886723,I886749,I886757,I886774,I886805,I886822,I886839,I886870,I886901,I886918,I886973,I886999,I887007,I887024,I887041,I887067,I887098,I887106,I887123,I887149,I887157,I887197,I887233,I887250,I887276,I887284,I887301,I887332,I887349,I887366,I887397,I887428,I887445,I887500,I887526,I887534,I887551,I887568,I887594,I887625,I887633,I887650,I887676,I887684,I887724,I887760,I887777,I887803,I887811,I887828,I887859,I887876,I887893,I887924,I887955,I887972,I888027,I888053,I888061,I888078,I888095,I888121,I888152,I888160,I888177,I888203,I888211,I888251,I888287,I888304,I888330,I888338,I888355,I888386,I888403,I888420,I888451,I888482,I888499,I888554,I888580,I888588,I888605,I888622,I888648,I888543,I888679,I888687,I888704,I888730,I888738,I888546,I888778,I888537,I888528,I888814,I888831,I888857,I888865,I888882,I888531,I888913,I888930,I888947,I888540,I888978,I888525,I889009,I889026,I888534,I889081,I889107,I889115,I889132,I889149,I889175,I889206,I889214,I889231,I889257,I889265,I889305,I889341,I889358,I889384,I889392,I889409,I889440,I889457,I889474,I889505,I889536,I889553,I889608,I889634,I889642,I889659,I889676,I889702,I889733,I889741,I889758,I889784,I889792,I889832,I889868,I889885,I889911,I889919,I889936,I889967,I889984,I890001,I890032,I890063,I890080,I890135,I890161,I890169,I890186,I890203,I890229,I890124,I890260,I890268,I890285,I890311,I890319,I890127,I890359,I890118,I890109,I890395,I890412,I890438,I890446,I890463,I890112,I890494,I890511,I890528,I890121,I890559,I890106,I890590,I890607,I890115,I890662,I890688,I890696,I890713,I890730,I890756,I890651,I890787,I890795,I890812,I890838,I890846,I890654,I890886,I890645,I890636,I890922,I890939,I890965,I890973,I890990,I890639,I891021,I891038,I891055,I890648,I891086,I890633,I891117,I891134,I890642,I891189,I891215,I891223,I891240,I891257,I891283,I891314,I891322,I891339,I891365,I891373,I891413,I891449,I891466,I891492,I891500,I891517,I891548,I891565,I891582,I891613,I891644,I891661,I891716,I1035680,I891742,I891750,I891767,I1035695,I1035677,I891784,I891810,I891705,I1035686,I891841,I891849,I1035704,I891866,I891892,I891900,I891708,I1035701,I891940,I891699,I891690,I891976,I1035698,I1035689,I891993,I1035683,I892019,I892027,I892044,I891693,I892075,I1035692,I892092,I892109,I891702,I892140,I891687,I892171,I892188,I891696,I892243,I892269,I892277,I892294,I892311,I892337,I892368,I892376,I892393,I892419,I892427,I892467,I892503,I892520,I892546,I892554,I892571,I892602,I892619,I892636,I892667,I892698,I892715,I892770,I892796,I892804,I892821,I892838,I892864,I892759,I892895,I892903,I892920,I892946,I892954,I892762,I892994,I892753,I892744,I893030,I893047,I893073,I893081,I893098,I892747,I893129,I893146,I893163,I892756,I893194,I892741,I893225,I893242,I892750,I893297,I1140143,I893323,I893331,I893348,I1140125,I893365,I1140131,I893391,I893286,I1140128,I893422,I893430,I1140137,I893447,I893473,I893481,I893289,I1140149,I893521,I893280,I893271,I893557,I1140140,I1140134,I893574,I893600,I893608,I893625,I893274,I893656,I1140146,I893673,I893690,I893283,I893721,I893268,I893752,I893769,I893277,I893824,I1227999,I893850,I893858,I893875,I1227981,I893892,I1227987,I893918,I893813,I1227984,I893949,I893957,I1227993,I893974,I894000,I894008,I893816,I1228005,I894048,I893807,I893798,I894084,I1227996,I1227990,I894101,I894127,I894135,I894152,I893801,I894183,I1228002,I894200,I894217,I893810,I894248,I893795,I894279,I894296,I893804,I894351,I894377,I894385,I894402,I894419,I894445,I894340,I894476,I894484,I894501,I894527,I894535,I894343,I894575,I894334,I894325,I894611,I894628,I894654,I894662,I894679,I894328,I894710,I894727,I894744,I894337,I894775,I894322,I894806,I894823,I894331,I894878,I894904,I894912,I894929,I894946,I894972,I895003,I895011,I895028,I895054,I895062,I895102,I895138,I895155,I895181,I895189,I895206,I895237,I895254,I895271,I895302,I895333,I895350,I895405,I895431,I895439,I895456,I895473,I895499,I895394,I895530,I895538,I895555,I895581,I895589,I895397,I895629,I895388,I895379,I895665,I895682,I895708,I895716,I895733,I895382,I895764,I895781,I895798,I895391,I895829,I895376,I895860,I895877,I895385,I895932,I895958,I895966,I895983,I896000,I896026,I896057,I896065,I896082,I896108,I896116,I896156,I896192,I896209,I896235,I896243,I896260,I896291,I896308,I896325,I896356,I896387,I896404,I896459,I990460,I896485,I896493,I896510,I990475,I990457,I896527,I896553,I990466,I896584,I896592,I990484,I896609,I896635,I896643,I990481,I896683,I896719,I990478,I990469,I896736,I990463,I896762,I896770,I896787,I896818,I990472,I896835,I896852,I896883,I896914,I896931,I896986,I1280693,I897012,I897020,I897037,I1280699,I1280681,I897054,I1280690,I897080,I1280696,I897111,I897119,I1280684,I897136,I897162,I897170,I1280702,I897210,I897246,I1280687,I897263,I1280705,I897289,I897297,I897314,I897345,I897362,I897379,I897410,I897441,I897458,I897513,I1038910,I897539,I897547,I897564,I1038925,I1038907,I897581,I897607,I1038916,I897638,I897646,I1038934,I897663,I897689,I897697,I1038931,I897737,I897773,I1038928,I1038919,I897790,I1038913,I897816,I897824,I897841,I897872,I1038922,I897889,I897906,I897937,I897968,I897985,I898040,I898066,I898074,I898091,I898108,I898134,I898165,I898173,I898190,I898216,I898224,I898264,I898300,I898317,I898343,I898351,I898368,I898399,I898416,I898433,I898464,I898495,I898512,I898567,I1053400,I898593,I898601,I898618,I1053409,I1053397,I898635,I1053394,I898661,I898692,I898700,I1053391,I898717,I898743,I898751,I898791,I898827,I1053412,I1053403,I898844,I1053406,I898870,I898878,I898895,I898926,I898943,I898960,I898991,I899022,I899039,I899094,I899120,I899128,I899145,I899162,I899188,I899083,I899219,I899227,I899244,I899270,I899278,I899086,I899318,I899077,I899068,I899354,I899371,I899397,I899405,I899422,I899071,I899453,I899470,I899487,I899080,I899518,I899065,I899549,I899566,I899074,I899621,I899647,I899655,I899672,I899689,I899715,I899746,I899754,I899771,I899797,I899805,I899845,I899881,I899898,I899924,I899932,I899949,I899980,I899997,I900014,I900045,I900076,I900093,I900148,I900174,I900182,I900199,I900216,I900242,I900137,I900273,I900281,I900298,I900324,I900332,I900140,I900372,I900131,I900122,I900408,I900425,I900451,I900459,I900476,I900125,I900507,I900524,I900541,I900134,I900572,I900119,I900603,I900620,I900128,I900675,I900701,I900709,I900726,I900743,I900769,I900800,I900808,I900825,I900851,I900859,I900899,I900935,I900952,I900978,I900986,I901003,I901034,I901051,I901068,I901099,I901130,I901147,I901202,I901228,I901236,I901253,I901270,I901296,I901191,I901327,I901335,I901352,I901378,I901386,I901194,I901426,I901185,I901176,I901462,I901479,I901505,I901513,I901530,I901179,I901561,I901578,I901595,I901188,I901626,I901173,I901657,I901674,I901182,I901729,I901755,I901763,I901780,I901797,I901823,I901854,I901862,I901879,I901905,I901913,I901953,I901989,I902006,I902032,I902040,I902057,I902088,I902105,I902122,I902153,I902184,I902201,I902256,I1057327,I902282,I902290,I902307,I1057336,I1057324,I902324,I1057321,I902350,I902381,I902389,I1057318,I902406,I902432,I902440,I902480,I902516,I1057339,I1057330,I902533,I1057333,I902559,I902567,I902584,I902615,I902632,I902649,I902680,I902711,I902728,I902783,I902809,I902817,I902834,I902851,I902877,I902772,I902908,I902916,I902933,I902959,I902967,I902775,I903007,I902766,I902757,I903043,I903060,I903086,I903094,I903111,I902760,I903142,I903159,I903176,I902769,I903207,I902754,I903238,I903255,I902763,I903310,I903336,I903344,I903361,I903378,I903404,I903299,I903435,I903443,I903460,I903486,I903494,I903302,I903534,I903293,I903284,I903570,I903587,I903613,I903621,I903638,I903287,I903669,I903686,I903703,I903296,I903734,I903281,I903765,I903782,I903290,I903837,I903863,I903871,I903888,I903905,I903931,I903962,I903970,I903987,I904013,I904021,I904061,I904097,I904114,I904140,I904148,I904165,I904196,I904213,I904230,I904261,I904292,I904309,I904364,I904390,I904398,I904415,I904432,I904458,I904489,I904497,I904514,I904540,I904548,I904588,I904624,I904641,I904667,I904675,I904692,I904723,I904740,I904757,I904788,I904819,I904836,I904891,I904917,I904925,I904942,I904959,I904985,I904880,I905016,I905024,I905041,I905067,I905075,I904883,I905115,I904874,I904865,I905151,I905168,I905194,I905202,I905219,I904868,I905250,I905267,I905284,I904877,I905315,I904862,I905346,I905363,I904871,I905418,I905444,I905452,I905469,I905486,I905512,I905543,I905551,I905568,I905594,I905602,I905642,I905678,I905695,I905721,I905729,I905746,I905777,I905794,I905811,I905842,I905873,I905890,I905945,I905971,I905979,I905996,I906013,I906039,I905934,I906070,I906078,I906095,I906121,I906129,I905937,I906169,I905928,I905919,I906205,I906222,I906248,I906256,I906273,I905922,I906304,I906321,I906338,I905931,I906369,I905916,I906400,I906417,I905925,I906472,I906498,I906506,I906523,I906540,I906566,I906597,I906605,I906622,I906648,I906656,I906696,I906732,I906749,I906775,I906783,I906800,I906831,I906848,I906865,I906896,I906927,I906944,I906999,I907025,I907033,I907050,I907067,I907093,I907124,I907132,I907149,I907175,I907183,I907223,I907259,I907276,I907302,I907310,I907327,I907358,I907375,I907392,I907423,I907454,I907471,I907526,I983354,I907552,I907560,I907577,I983369,I983351,I907594,I907620,I983360,I907651,I907659,I983378,I907676,I907702,I907710,I983375,I907750,I907786,I983372,I983363,I907803,I983357,I907829,I907837,I907854,I907885,I983366,I907902,I907919,I907950,I907981,I907998,I908053,I908079,I908087,I908104,I908121,I908147,I908178,I908186,I908203,I908229,I908237,I908277,I908313,I908330,I908356,I908364,I908381,I908412,I908429,I908446,I908477,I908508,I908525,I908580,I908606,I908614,I908631,I908648,I908674,I908705,I908713,I908730,I908756,I908764,I908804,I908840,I908857,I908883,I908891,I908908,I908939,I908956,I908973,I909004,I909035,I909052,I909107,I909133,I909141,I909158,I909175,I909201,I909232,I909240,I909257,I909283,I909291,I909331,I909367,I909384,I909410,I909418,I909435,I909466,I909483,I909500,I909531,I909562,I909579,I909634,I909660,I909668,I909685,I909702,I909728,I909623,I909759,I909767,I909784,I909810,I909818,I909626,I909858,I909617,I909608,I909894,I909911,I909937,I909945,I909962,I909611,I909993,I910010,I910027,I909620,I910058,I909605,I910089,I910106,I909614,I910161,I989814,I910187,I910195,I910212,I989829,I989811,I910229,I910255,I910150,I989820,I910286,I910294,I989838,I910311,I910337,I910345,I910153,I989835,I910385,I910144,I910135,I910421,I989832,I989823,I910438,I989817,I910464,I910472,I910489,I910138,I910520,I989826,I910537,I910554,I910147,I910585,I910132,I910616,I910633,I910141,I910688,I1067986,I910714,I910722,I910739,I1067995,I1067983,I910756,I1067980,I910782,I910677,I910813,I910821,I1067977,I910838,I910864,I910872,I910680,I910912,I910671,I910662,I910948,I1067998,I1067989,I910965,I1067992,I910991,I910999,I911016,I910665,I911047,I911064,I911081,I910674,I911112,I910659,I911143,I911160,I910668,I911215,I911241,I911249,I911266,I911283,I911309,I911204,I911340,I911348,I911365,I911391,I911399,I911207,I911439,I911198,I911189,I911475,I911492,I911518,I911526,I911543,I911192,I911574,I911591,I911608,I911201,I911639,I911186,I911670,I911687,I911195,I911742,I911768,I911776,I911793,I911810,I911836,I911731,I911867,I911875,I911892,I911918,I911926,I911734,I911966,I911725,I911716,I912002,I912019,I912045,I912053,I912070,I911719,I912101,I912118,I912135,I911728,I912166,I911713,I912197,I912214,I911722,I912269,I1014362,I912295,I912303,I912320,I1014377,I1014359,I912337,I912363,I1014368,I912394,I912402,I1014386,I912419,I912445,I912453,I1014383,I912493,I912529,I1014380,I1014371,I912546,I1014365,I912572,I912580,I912597,I912628,I1014374,I912645,I912662,I912693,I912724,I912741,I912796,I912822,I912830,I912847,I912864,I912890,I912921,I912929,I912946,I912972,I912980,I913020,I913056,I913073,I913099,I913107,I913124,I913155,I913172,I913189,I913220,I913251,I913268,I913323,I913349,I913357,I913374,I913391,I913417,I913448,I913456,I913473,I913499,I913507,I913547,I913583,I913600,I913626,I913634,I913651,I913682,I913699,I913716,I913747,I913778,I913795,I913850,I1192163,I913876,I913884,I913901,I1192145,I913918,I1192151,I913944,I1192148,I913975,I913983,I1192157,I914000,I914026,I914034,I1192169,I914074,I914110,I1192160,I1192154,I914127,I914153,I914161,I914178,I914209,I1192166,I914226,I914243,I914274,I914305,I914322,I914377,I914403,I914411,I914428,I914445,I914471,I914366,I914502,I914510,I914527,I914553,I914561,I914369,I914601,I914360,I914351,I914637,I914654,I914680,I914688,I914705,I914354,I914736,I914753,I914770,I914363,I914801,I914348,I914832,I914849,I914357,I914910,I1321286,I914936,I1321280,I914953,I914961,I914978,I1321289,I914995,I1321301,I915012,I1321283,I915029,I915046,I915077,I915094,I915125,I915142,I1321277,I915159,I915190,I915230,I915238,I915255,I915272,I1321298,I915289,I915320,I1321292,I915337,I915354,I1321295,I915380,I915402,I915419,I915450,I915495,I915556,I915582,I915599,I915607,I915624,I915641,I915658,I915675,I915692,I915723,I915740,I915771,I915788,I915805,I915836,I915876,I915884,I915901,I915918,I915935,I915966,I915983,I916000,I916026,I916048,I916065,I916096,I916141,I916202,I916228,I916245,I916253,I916270,I916287,I916304,I916321,I916338,I916188,I916369,I916386,I916191,I916417,I916434,I916451,I916167,I916482,I916179,I916522,I916530,I916547,I916564,I916581,I916194,I916612,I916629,I916646,I916672,I916182,I916694,I916711,I916176,I916742,I916170,I916173,I916787,I916185,I916848,I916874,I916891,I916899,I916916,I916933,I916950,I916967,I916984,I917015,I917032,I917063,I917080,I917097,I917128,I917168,I917176,I917193,I917210,I917227,I917258,I917275,I917292,I917318,I917340,I917357,I917388,I917433,I917494,I917520,I917537,I917545,I917562,I917579,I917596,I917613,I917630,I917661,I917678,I917709,I917726,I917743,I917774,I917814,I917822,I917839,I917856,I917873,I917904,I917921,I917938,I917964,I917986,I918003,I918034,I918079,I918140,I1407688,I918166,I1407712,I918183,I918191,I918208,I1407694,I918225,I1407703,I918242,I918259,I1407709,I918276,I918307,I918324,I918355,I918372,I1407706,I918389,I918420,I918460,I918468,I918485,I918502,I1407700,I918519,I918550,I1407691,I918567,I1407715,I918584,I1407697,I918610,I918632,I918649,I918680,I918725,I918786,I1330338,I918812,I1330362,I918829,I918837,I918854,I1330344,I918871,I1330353,I918888,I918905,I1330359,I918922,I918953,I918970,I919001,I919018,I1330356,I919035,I919066,I919106,I919114,I919131,I919148,I1330350,I919165,I919196,I1330341,I919213,I1330365,I919230,I1330347,I919256,I919278,I919295,I919326,I919371,I919432,I919458,I919475,I919483,I919500,I919517,I919534,I919551,I919568,I919599,I919616,I919647,I919664,I919681,I919712,I919752,I919760,I919777,I919794,I919811,I919842,I919859,I919876,I919902,I919924,I919941,I919972,I920017,I920078,I920104,I920121,I920129,I920146,I920163,I920180,I920197,I920214,I920245,I920262,I920293,I920310,I920327,I920358,I920398,I920406,I920423,I920440,I920457,I920488,I920505,I920522,I920548,I920570,I920587,I920618,I920663,I920724,I920750,I920767,I920775,I920792,I920809,I920826,I920843,I920860,I920891,I920908,I920939,I920956,I920973,I921004,I921044,I921052,I921069,I921086,I921103,I921134,I921151,I921168,I921194,I921216,I921233,I921264,I921309,I921370,I921396,I921413,I921421,I921438,I921455,I921472,I921489,I921506,I921537,I921554,I921585,I921602,I921619,I921650,I921690,I921698,I921715,I921732,I921749,I921780,I921797,I921814,I921840,I921862,I921879,I921910,I921955,I922016,I1254587,I922042,I1254593,I922059,I922067,I922084,I1254590,I922101,I1254569,I922118,I1254572,I922135,I1254578,I922152,I922183,I922200,I922231,I922248,I922265,I922296,I922336,I922344,I922361,I922378,I1254581,I922395,I922426,I922443,I1254575,I922460,I1254584,I922486,I922508,I922525,I922556,I922601,I922662,I922688,I922705,I922713,I922730,I922747,I922764,I922781,I922798,I922829,I922846,I922877,I922894,I922911,I922942,I922982,I922990,I923007,I923024,I923041,I923072,I923089,I923106,I923132,I923154,I923171,I923202,I923247,I923308,I923334,I923351,I923359,I923376,I923393,I923410,I923427,I923444,I923475,I923492,I923523,I923540,I923557,I923588,I923628,I923636,I923653,I923670,I923687,I923718,I923735,I923752,I923778,I923800,I923817,I923848,I923893,I923954,I1099105,I923980,I1099087,I923997,I924005,I924022,I1099096,I924039,I1099108,I924056,I1099090,I924073,I1099099,I924090,I923940,I924121,I924138,I923943,I924169,I924186,I1099111,I924203,I923919,I924234,I923931,I924274,I924282,I924299,I924316,I924333,I923946,I924364,I1099093,I924381,I1099102,I924398,I924424,I923934,I924446,I924463,I923928,I924494,I923922,I923925,I924539,I923937,I924600,I924626,I924643,I924651,I924668,I924685,I924702,I924719,I924736,I924586,I924767,I924784,I924589,I924815,I924832,I924849,I924565,I924880,I924577,I924920,I924928,I924945,I924962,I924979,I924592,I925010,I925027,I925044,I925070,I924580,I925092,I925109,I924574,I925140,I924568,I924571,I925185,I924583,I925246,I925272,I925289,I925297,I925314,I925331,I925348,I925365,I925382,I925413,I925430,I925461,I925478,I925495,I925526,I925566,I925574,I925591,I925608,I925625,I925656,I925673,I925690,I925716,I925738,I925755,I925786,I925831,I925892,I925918,I925935,I925943,I925960,I925977,I925994,I926011,I926028,I926059,I926076,I926107,I926124,I926141,I926172,I926212,I926220,I926237,I926254,I926271,I926302,I926319,I926336,I926362,I926384,I926401,I926432,I926477,I926538,I926564,I926581,I926589,I926606,I926623,I926640,I926657,I926674,I926705,I926722,I926753,I926770,I926787,I926818,I926858,I926866,I926883,I926900,I926917,I926948,I926965,I926982,I927008,I927030,I927047,I927078,I927123,I927184,I927210,I927227,I927235,I927252,I927269,I927286,I927303,I927320,I927351,I927368,I927399,I927416,I927433,I927464,I927504,I927512,I927529,I927546,I927563,I927594,I927611,I927628,I927654,I927676,I927693,I927724,I927769,I927830,I927856,I927873,I927881,I927898,I927915,I927932,I927949,I927966,I927816,I927997,I928014,I927819,I928045,I928062,I928079,I927795,I928110,I927807,I928150,I928158,I928175,I928192,I928209,I927822,I928240,I928257,I928274,I928300,I927810,I928322,I928339,I927804,I928370,I927798,I927801,I928415,I927813,I928476,I928502,I928519,I928527,I928544,I928561,I928578,I928595,I928612,I928643,I928660,I928691,I928708,I928725,I928756,I928796,I928804,I928821,I928838,I928855,I928886,I928903,I928920,I928946,I928968,I928985,I929016,I929061,I929122,I929148,I929165,I929173,I929190,I929207,I929224,I929241,I929258,I929108,I929289,I929306,I929111,I929337,I929354,I929371,I929087,I929402,I929099,I929442,I929450,I929467,I929484,I929501,I929114,I929532,I929549,I929566,I929592,I929102,I929614,I929631,I929096,I929662,I929090,I929093,I929707,I929105,I929768,I1230889,I929794,I1230871,I929811,I929819,I929836,I1230880,I929853,I1230892,I929870,I1230874,I929887,I1230883,I929904,I929754,I929935,I929952,I929757,I929983,I930000,I1230895,I930017,I929733,I930048,I929745,I930088,I930096,I930113,I930130,I930147,I929760,I930178,I1230877,I930195,I1230886,I930212,I930238,I929748,I930260,I930277,I929742,I930308,I929736,I929739,I930353,I929751,I930414,I930440,I930457,I930465,I930482,I930499,I930516,I930533,I930550,I930581,I930598,I930629,I930646,I930663,I930694,I930734,I930742,I930759,I930776,I930793,I930824,I930841,I930858,I930884,I930906,I930923,I930954,I930999,I931060,I1156327,I931086,I1156309,I931103,I931111,I931128,I1156318,I931145,I1156330,I931162,I1156312,I931179,I1156321,I931196,I931227,I931244,I931275,I931292,I1156333,I931309,I931340,I931380,I931388,I931405,I931422,I931439,I931470,I1156315,I931487,I1156324,I931504,I931530,I931552,I931569,I931600,I931645,I931706,I931732,I931749,I931757,I931774,I931791,I931808,I931825,I931842,I931873,I931890,I931921,I931938,I931955,I931986,I932026,I932034,I932051,I932068,I932085,I932116,I932133,I932150,I932176,I932198,I932215,I932246,I932291,I932352,I1110087,I932378,I1110069,I932395,I932403,I932420,I1110078,I932437,I1110090,I932454,I1110072,I932471,I1110081,I932488,I932519,I932536,I932567,I932584,I1110093,I932601,I932632,I932672,I932680,I932697,I932714,I932731,I932762,I1110075,I932779,I1110084,I932796,I932822,I932844,I932861,I932892,I932937,I932998,I933024,I933041,I933049,I933066,I933083,I933100,I933117,I933134,I933165,I933182,I933213,I933230,I933247,I933278,I933318,I933326,I933343,I933360,I933377,I933408,I933425,I933442,I933468,I933490,I933507,I933538,I933583,I933644,I933670,I933687,I933695,I933712,I933729,I933746,I933763,I933780,I933811,I933828,I933859,I933876,I933893,I933924,I933964,I933972,I933989,I934006,I934023,I934054,I934071,I934088,I934114,I934136,I934153,I934184,I934229,I934290,I934316,I934333,I934341,I934358,I934375,I934392,I934409,I934426,I934457,I934474,I934505,I934522,I934539,I934570,I934610,I934618,I934635,I934652,I934669,I934700,I934717,I934734,I934760,I934782,I934799,I934830,I934875,I934936,I934962,I934979,I934987,I935004,I935021,I935038,I935055,I935072,I934922,I935103,I935120,I934925,I935151,I935168,I935185,I934901,I935216,I934913,I935256,I935264,I935281,I935298,I935315,I934928,I935346,I935363,I935380,I935406,I934916,I935428,I935445,I934910,I935476,I934904,I934907,I935521,I934919,I935582,I935608,I935625,I935633,I935650,I935667,I935684,I935701,I935718,I935749,I935766,I935797,I935814,I935831,I935862,I935902,I935910,I935927,I935944,I935961,I935992,I936009,I936026,I936052,I936074,I936091,I936122,I936167,I936228,I936254,I936271,I936279,I936296,I936313,I936330,I936347,I936364,I936395,I936412,I936443,I936460,I936477,I936508,I936548,I936556,I936573,I936590,I936607,I936638,I936655,I936672,I936698,I936720,I936737,I936768,I936813,I936874,I936900,I936917,I936925,I936942,I936959,I936976,I936993,I937010,I936860,I937041,I937058,I936863,I937089,I937106,I937123,I936839,I937154,I936851,I937194,I937202,I937219,I937236,I937253,I936866,I937284,I937301,I937318,I937344,I936854,I937366,I937383,I936848,I937414,I936842,I936845,I937459,I936857,I937520,I937546,I937563,I937571,I937588,I937605,I937622,I937639,I937656,I937687,I937704,I937735,I937752,I937769,I937800,I937840,I937848,I937865,I937882,I937899,I937930,I937947,I937964,I937990,I938012,I938029,I938060,I938105,I938166,I1208347,I938192,I1208329,I938209,I938217,I938234,I1208338,I938251,I1208350,I938268,I1208332,I938285,I1208341,I938302,I938152,I938333,I938350,I938155,I938381,I938398,I1208353,I938415,I938131,I938446,I938143,I938486,I938494,I938511,I938528,I938545,I938158,I938576,I1208335,I938593,I1208344,I938610,I938636,I938146,I938658,I938675,I938140,I938706,I938134,I938137,I938751,I938149,I938812,I938838,I938855,I938863,I938880,I938897,I938914,I938931,I938948,I938979,I938996,I939027,I939044,I939061,I939092,I939132,I939140,I939157,I939174,I939191,I939222,I939239,I939256,I939282,I939304,I939321,I939352,I939397,I939458,I1335693,I939484,I1335717,I939501,I939509,I939526,I1335699,I939543,I1335708,I939560,I939577,I1335714,I939594,I939625,I939642,I939673,I939690,I1335711,I939707,I939738,I939778,I939786,I939803,I939820,I1335705,I939837,I939868,I1335696,I939885,I1335720,I939902,I1335702,I939928,I939950,I939967,I939998,I940043,I940104,I940130,I940147,I940155,I940172,I940189,I940206,I940223,I940240,I940271,I940288,I940319,I940336,I940353,I940384,I940424,I940432,I940449,I940466,I940483,I940514,I940531,I940548,I940574,I940596,I940613,I940644,I940689,I940750,I940776,I940793,I940801,I940818,I940835,I940852,I940869,I940886,I940917,I940934,I940965,I940982,I940999,I941030,I941070,I941078,I941095,I941112,I941129,I941160,I941177,I941194,I941220,I941242,I941259,I941290,I941335,I941396,I1341643,I941422,I1341667,I941439,I941447,I941464,I1341649,I941481,I1341658,I941498,I941515,I1341664,I941532,I941382,I941563,I941580,I941385,I941611,I941628,I1341661,I941645,I941361,I941676,I941373,I941716,I941724,I941741,I941758,I1341655,I941775,I941388,I941806,I1341646,I941823,I1341670,I941840,I1341652,I941866,I941376,I941888,I941905,I941370,I941936,I941364,I941367,I941981,I941379,I942042,I942068,I942085,I942093,I942110,I942127,I942144,I942161,I942178,I942028,I942209,I942226,I942031,I942257,I942274,I942291,I942007,I942322,I942019,I942362,I942370,I942387,I942404,I942421,I942034,I942452,I942469,I942486,I942512,I942022,I942534,I942551,I942016,I942582,I942010,I942013,I942627,I942025,I942688,I942714,I942731,I942739,I942756,I942773,I942790,I942807,I942824,I942855,I942872,I942903,I942920,I942937,I942968,I943008,I943016,I943033,I943050,I943067,I943098,I943115,I943132,I943158,I943180,I943197,I943228,I943273,I943334,I1071904,I943360,I1071907,I943377,I943385,I943402,I943419,I1071916,I943436,I1071925,I943453,I1071913,I943470,I943501,I943518,I943549,I943566,I1071919,I943583,I943614,I943654,I943662,I943679,I943696,I1071910,I943713,I943744,I1071922,I943761,I943778,I943804,I943826,I943843,I943874,I943919,I943980,I944006,I944023,I944031,I944048,I944065,I944082,I944099,I944116,I944147,I944164,I944195,I944212,I944229,I944260,I944300,I944308,I944325,I944342,I944359,I944390,I944407,I944424,I944450,I944472,I944489,I944520,I944565,I944626,I944652,I944669,I944677,I944694,I944711,I944728,I944745,I944762,I944793,I944810,I944841,I944858,I944875,I944906,I944946,I944954,I944971,I944988,I945005,I945036,I945053,I945070,I945096,I945118,I945135,I945166,I945211,I945272,I945298,I945315,I945323,I945340,I945357,I945374,I945391,I945408,I945439,I945456,I945487,I945504,I945521,I945552,I945592,I945600,I945617,I945634,I945651,I945682,I945699,I945716,I945742,I945764,I945781,I945812,I945857,I945918,I945944,I945961,I945969,I945986,I946003,I946020,I946037,I946054,I946085,I946102,I946133,I946150,I946167,I946198,I946238,I946246,I946263,I946280,I946297,I946328,I946345,I946362,I946388,I946410,I946427,I946458,I946503,I946564,I1148813,I946590,I1148795,I946607,I946615,I946632,I1148804,I946649,I1148816,I946666,I1148798,I946683,I1148807,I946700,I946731,I946748,I946779,I946796,I1148819,I946813,I946844,I946884,I946892,I946909,I946926,I946943,I946974,I1148801,I946991,I1148810,I947008,I947034,I947056,I947073,I947104,I947149,I947210,I947236,I947253,I947261,I947278,I947295,I947312,I947329,I947346,I947377,I947394,I947425,I947442,I947459,I947490,I947530,I947538,I947555,I947572,I947589,I947620,I947637,I947654,I947680,I947702,I947719,I947750,I947795,I947856,I947882,I947899,I947907,I947924,I947941,I947958,I947975,I947992,I948023,I948040,I948071,I948088,I948105,I948136,I948176,I948184,I948201,I948218,I948235,I948266,I948283,I948300,I948326,I948348,I948365,I948396,I948441,I948502,I948528,I948545,I948553,I948570,I948587,I948604,I948621,I948638,I948669,I948686,I948717,I948734,I948751,I948782,I948822,I948830,I948847,I948864,I948881,I948912,I948929,I948946,I948972,I948994,I949011,I949042,I949087,I949148,I1369013,I949174,I1369037,I949191,I949199,I949216,I1369019,I949233,I1369028,I949250,I949267,I1369034,I949284,I949315,I949332,I949363,I949380,I1369031,I949397,I949428,I949468,I949476,I949493,I949510,I1369025,I949527,I949558,I1369016,I949575,I1369040,I949592,I1369022,I949618,I949640,I949657,I949688,I949733,I949794,I949820,I949837,I949845,I949862,I949879,I949896,I949913,I949930,I949961,I949978,I950009,I950026,I950043,I950074,I950114,I950122,I950139,I950156,I950173,I950204,I950221,I950238,I950264,I950286,I950303,I950334,I950379,I950440,I950466,I950483,I950491,I950508,I950525,I950542,I950559,I950576,I950607,I950624,I950655,I950672,I950689,I950720,I950760,I950768,I950785,I950802,I950819,I950850,I950867,I950884,I950910,I950932,I950949,I950980,I951025,I951086,I1255131,I951112,I1255137,I951129,I951137,I951154,I1255134,I951171,I1255113,I951188,I1255116,I951205,I1255122,I951222,I951253,I951270,I951301,I951318,I951335,I951366,I951406,I951414,I951431,I951448,I1255125,I951465,I951496,I951513,I1255119,I951530,I1255128,I951556,I951578,I951595,I951626,I951671,I951732,I951758,I951775,I951783,I951800,I951817,I951834,I951851,I951868,I951718,I951899,I951916,I951721,I951947,I951964,I951981,I951697,I952012,I951709,I952052,I952060,I952077,I952094,I952111,I951724,I952142,I952159,I952176,I952202,I951712,I952224,I952241,I951706,I952272,I951700,I951703,I952317,I951715,I952378,I952404,I952421,I952429,I952446,I952463,I952480,I952497,I952514,I952545,I952562,I952593,I952610,I952627,I952658,I952698,I952706,I952723,I952740,I952757,I952788,I952805,I952822,I952848,I952870,I952887,I952918,I952963,I953024,I953050,I953067,I953075,I953092,I953109,I953126,I953143,I953160,I953191,I953208,I953239,I953256,I953273,I953304,I953344,I953352,I953369,I953386,I953403,I953434,I953451,I953468,I953494,I953516,I953533,I953564,I953609,I953670,I953696,I953713,I953721,I953738,I953755,I953772,I953789,I953806,I953837,I953854,I953885,I953902,I953919,I953950,I953990,I953998,I954015,I954032,I954049,I954080,I954097,I954114,I954140,I954162,I954179,I954210,I954255,I954316,I954342,I954359,I954367,I954384,I954401,I954418,I954435,I954452,I954483,I954500,I954531,I954548,I954565,I954596,I954636,I954644,I954661,I954678,I954695,I954726,I954743,I954760,I954786,I954808,I954825,I954856,I954901,I954962,I954988,I955005,I955013,I955030,I955047,I955064,I955081,I955098,I954948,I955129,I955146,I954951,I955177,I955194,I955211,I954927,I955242,I954939,I955282,I955290,I955307,I955324,I955341,I954954,I955372,I955389,I955406,I955432,I954942,I955454,I955471,I954936,I955502,I954930,I954933,I955547,I954945,I955608,I1341048,I955634,I1341072,I955651,I955659,I955676,I1341054,I955693,I1341063,I955710,I955727,I1341069,I955744,I955775,I955792,I955823,I955840,I1341066,I955857,I955888,I955928,I955936,I955953,I955970,I1341060,I955987,I956018,I1341051,I956035,I1341075,I956052,I1341057,I956078,I956100,I956117,I956148,I956193,I956254,I956280,I956297,I956305,I956322,I956339,I956356,I956373,I956390,I956421,I956438,I956469,I956486,I956503,I956534,I956574,I956582,I956599,I956616,I956633,I956664,I956681,I956698,I956724,I956746,I956763,I956794,I956839,I956900,I956926,I956943,I956951,I956968,I956985,I957002,I957019,I957036,I957067,I957084,I957115,I957132,I957149,I957180,I957220,I957228,I957245,I957262,I957279,I957310,I957327,I957344,I957370,I957392,I957409,I957440,I957485,I957546,I957572,I957589,I957597,I957614,I957631,I957648,I957665,I957682,I957713,I957730,I957761,I957778,I957795,I957826,I957866,I957874,I957891,I957908,I957925,I957956,I957973,I957990,I958016,I958038,I958055,I958086,I958131,I958192,I1112977,I958218,I1112959,I958235,I958243,I958260,I1112968,I958277,I1112980,I958294,I1112962,I958311,I1112971,I958328,I958359,I958376,I958407,I958424,I1112983,I958441,I958472,I958512,I958520,I958537,I958554,I958571,I958602,I1112965,I958619,I1112974,I958636,I958662,I958684,I958701,I958732,I958777,I958838,I958864,I958881,I958889,I958906,I958923,I958940,I958957,I958974,I959005,I959022,I959053,I959070,I959087,I959118,I959158,I959166,I959183,I959200,I959217,I959248,I959265,I959282,I959308,I959330,I959347,I959378,I959423,I959484,I959510,I959527,I959535,I959552,I959569,I959586,I959603,I959620,I959651,I959668,I959699,I959716,I959733,I959764,I959804,I959812,I959829,I959846,I959863,I959894,I959911,I959928,I959954,I959976,I959993,I960024,I960069,I960130,I960156,I960173,I960181,I960198,I960215,I960232,I960249,I960266,I960297,I960314,I960345,I960362,I960379,I960410,I960450,I960458,I960475,I960492,I960509,I960540,I960557,I960574,I960600,I960622,I960639,I960670,I960715,I960776,I960802,I960819,I960827,I960844,I960861,I960878,I960895,I960912,I960943,I960960,I960991,I961008,I961025,I961056,I961096,I961104,I961121,I961138,I961155,I961186,I961203,I961220,I961246,I961268,I961285,I961316,I961361,I961422,I1258939,I961448,I1258945,I961465,I961473,I961490,I1258942,I961507,I1258921,I961524,I1258924,I961541,I1258930,I961558,I961408,I961589,I961606,I961411,I961637,I961654,I961671,I961387,I961702,I961399,I961742,I961750,I961767,I961784,I1258933,I961801,I961414,I961832,I961849,I1258927,I961866,I1258936,I961892,I961402,I961914,I961931,I961396,I961962,I961390,I961393,I962007,I961405,I962068,I962094,I962111,I962119,I962136,I962153,I962170,I962187,I962204,I962235,I962252,I962283,I962300,I962317,I962348,I962388,I962396,I962413,I962430,I962447,I962478,I962495,I962512,I962538,I962560,I962577,I962608,I962653,I962714,I962740,I962757,I962765,I962782,I962799,I962816,I962833,I962850,I962881,I962898,I962929,I962946,I962963,I962994,I963034,I963042,I963059,I963076,I963093,I963124,I963141,I963158,I963184,I963206,I963223,I963254,I963299,I963360,I1383888,I963386,I1383912,I963403,I963411,I963428,I1383894,I963445,I1383903,I963462,I963479,I1383909,I963496,I963527,I963544,I963575,I963592,I1383906,I963609,I963640,I963680,I963688,I963705,I963722,I1383900,I963739,I963770,I1383891,I963787,I1383915,I963804,I1383897,I963830,I963852,I963869,I963900,I963945,I964006,I964032,I964049,I964057,I964074,I964091,I964108,I964125,I964142,I963992,I964173,I964190,I963995,I964221,I964238,I964255,I963971,I964286,I963983,I964326,I964334,I964351,I964368,I964385,I963998,I964416,I964433,I964450,I964476,I963986,I964498,I964515,I963980,I964546,I963974,I963977,I964591,I963989,I964652,I964678,I964695,I964703,I964720,I964737,I964754,I964771,I964788,I964819,I964836,I964867,I964884,I964901,I964932,I964972,I964980,I964997,I965014,I965031,I965062,I965079,I965096,I965122,I965144,I965161,I965192,I965237,I965298,I1218173,I965324,I1218155,I965341,I965349,I965366,I1218164,I965383,I1218176,I965400,I1218158,I965417,I1218167,I965434,I965465,I965482,I965513,I965530,I1218179,I965547,I965578,I965618,I965626,I965643,I965660,I965677,I965708,I1218161,I965725,I1218170,I965742,I965768,I965790,I965807,I965838,I965883,I965944,I1226265,I965970,I1226247,I965987,I965995,I966012,I1226256,I966029,I1226268,I966046,I1226250,I966063,I1226259,I966080,I966111,I966128,I966159,I966176,I1226271,I966193,I966224,I966264,I966272,I966289,I966306,I966323,I966354,I1226253,I966371,I1226262,I966388,I966414,I966436,I966453,I966484,I966529,I966590,I966616,I966633,I966641,I966658,I966675,I966692,I966709,I966726,I966576,I966757,I966774,I966579,I966805,I966822,I966839,I966555,I966870,I966567,I966910,I966918,I966935,I966952,I966969,I966582,I967000,I967017,I967034,I967060,I966570,I967082,I967099,I966564,I967130,I966558,I966561,I967175,I966573,I967236,I1321864,I967262,I1321858,I967279,I967287,I967304,I1321867,I967321,I1321879,I967338,I1321861,I967355,I967372,I967403,I967420,I967451,I967468,I1321855,I967485,I967516,I967556,I967564,I967581,I967598,I1321876,I967615,I967646,I1321870,I967663,I967680,I1321873,I967706,I967728,I967745,I967776,I967821,I967882,I967908,I967925,I967933,I967950,I967967,I967984,I968001,I968018,I968049,I968066,I968097,I968114,I968131,I968162,I968202,I968210,I968227,I968244,I968261,I968292,I968309,I968326,I968352,I968374,I968391,I968422,I968467,I968528,I968554,I968571,I968579,I968596,I968613,I968630,I968647,I968664,I968514,I968695,I968712,I968517,I968743,I968760,I968777,I968493,I968808,I968505,I968848,I968856,I968873,I968890,I968907,I968520,I968938,I968955,I968972,I968998,I968508,I969020,I969037,I968502,I969068,I968496,I968499,I969113,I968511,I969174,I969200,I969217,I969225,I969242,I969259,I969276,I969293,I969310,I969341,I969358,I969389,I969406,I969423,I969454,I969494,I969502,I969519,I969536,I969553,I969584,I969601,I969618,I969644,I969666,I969683,I969714,I969759,I969820,I969846,I969863,I969871,I969888,I969905,I969922,I969939,I969956,I969987,I970004,I970035,I970052,I970069,I970100,I970140,I970148,I970165,I970182,I970199,I970230,I970247,I970264,I970290,I970312,I970329,I970360,I970405,I970466,I970492,I970509,I970517,I970534,I970551,I970568,I970585,I970602,I970633,I970650,I970681,I970698,I970715,I970746,I970786,I970794,I970811,I970828,I970845,I970876,I970893,I970910,I970936,I970958,I970975,I971006,I971051,I971112,I971138,I971155,I971163,I971180,I971197,I971214,I971231,I971248,I971098,I971279,I971296,I971101,I971327,I971344,I971361,I971077,I971392,I971089,I971432,I971440,I971457,I971474,I971491,I971104,I971522,I971539,I971556,I971582,I971092,I971604,I971621,I971086,I971652,I971080,I971083,I971697,I971095,I971758,I971784,I971801,I971809,I971826,I971843,I971860,I971877,I971894,I971925,I971942,I971973,I971990,I972007,I972038,I972078,I972086,I972103,I972120,I972137,I972168,I972185,I972202,I972228,I972250,I972267,I972298,I972343,I972404,I972430,I972447,I972455,I972472,I972489,I972506,I972523,I972540,I972390,I972571,I972588,I972393,I972619,I972636,I972653,I972369,I972684,I972381,I972724,I972732,I972749,I972766,I972783,I972396,I972814,I972831,I972848,I972874,I972384,I972896,I972913,I972378,I972944,I972372,I972375,I972989,I972387,I973050,I973076,I973093,I973101,I973118,I973135,I973152,I973169,I973186,I973036,I973217,I973234,I973039,I973265,I973282,I973299,I973015,I973330,I973027,I973370,I973378,I973395,I973412,I973429,I973042,I973460,I973477,I973494,I973520,I973030,I973542,I973559,I973024,I973590,I973018,I973021,I973635,I973033,I973696,I973722,I973739,I973747,I973764,I973781,I973798,I973815,I973832,I973863,I973880,I973911,I973928,I973945,I973976,I974016,I974024,I974041,I974058,I974075,I974106,I974123,I974140,I974166,I974188,I974205,I974236,I974281,I974342,I974368,I974385,I974393,I974410,I974427,I974444,I974461,I974478,I974509,I974526,I974557,I974574,I974591,I974622,I974662,I974670,I974687,I974704,I974721,I974752,I974769,I974786,I974812,I974834,I974851,I974882,I974927,I974988,I975014,I975031,I975039,I975056,I975073,I975090,I975107,I975124,I974974,I975155,I975172,I974977,I975203,I975220,I975237,I974953,I975268,I974965,I975308,I975316,I975333,I975350,I975367,I974980,I975398,I975415,I975432,I975458,I974968,I975480,I975497,I974962,I975528,I974956,I974959,I975573,I974971,I975634,I975660,I975677,I975685,I975702,I975719,I975736,I975753,I975770,I975801,I975818,I975849,I975866,I975883,I975914,I975954,I975962,I975979,I975996,I976013,I976044,I976061,I976078,I976104,I976126,I976143,I976174,I976219,I976280,I976306,I976323,I976331,I976348,I976365,I976382,I976399,I976416,I976447,I976464,I976495,I976512,I976529,I976560,I976600,I976608,I976625,I976642,I976659,I976690,I976707,I976724,I976750,I976772,I976789,I976820,I976865,I976926,I976952,I976969,I976977,I976994,I977011,I977028,I977045,I977062,I977093,I977110,I977141,I977158,I977175,I977206,I977246,I977254,I977271,I977288,I977305,I977336,I977353,I977370,I977396,I977418,I977435,I977466,I977511,I977572,I977598,I977615,I977623,I977640,I977657,I977674,I977691,I977708,I977739,I977756,I977787,I977804,I977821,I977852,I977892,I977900,I977917,I977934,I977951,I977982,I977999,I978016,I978042,I978064,I978081,I978112,I978157,I978218,I1225109,I978244,I1225091,I978261,I978269,I978286,I1225100,I978303,I1225112,I978320,I1225094,I978337,I1225103,I978354,I978204,I978385,I978402,I978207,I978433,I978450,I1225115,I978467,I978183,I978498,I978195,I978538,I978546,I978563,I978580,I978597,I978210,I978628,I1225097,I978645,I1225106,I978662,I978688,I978198,I978710,I978727,I978192,I978758,I978186,I978189,I978803,I978201,I978864,I978890,I978907,I978915,I978932,I978949,I978966,I978983,I979000,I979031,I979048,I979079,I979096,I979113,I979144,I979184,I979192,I979209,I979226,I979243,I979274,I979291,I979308,I979334,I979356,I979373,I979404,I979449,I979510,I979536,I979553,I979561,I979578,I979595,I979612,I979629,I979646,I979677,I979694,I979725,I979742,I979759,I979790,I979830,I979838,I979855,I979872,I979889,I979920,I979937,I979954,I979980,I980002,I980019,I980050,I980095,I980156,I980182,I980199,I980207,I980224,I980241,I980258,I980275,I980292,I980323,I980340,I980371,I980388,I980405,I980436,I980476,I980484,I980501,I980518,I980535,I980566,I980583,I980600,I980626,I980648,I980665,I980696,I980741,I980802,I980828,I980845,I980853,I980870,I980887,I980904,I980921,I980938,I980969,I980986,I981017,I981034,I981051,I981082,I981122,I981130,I981147,I981164,I981181,I981212,I981229,I981246,I981272,I981294,I981311,I981342,I981387,I981448,I1100839,I981474,I1100821,I981491,I981499,I981516,I1100830,I981533,I1100842,I981550,I1100824,I981567,I1100833,I981584,I981615,I981632,I981663,I981680,I1100845,I981697,I981728,I981768,I981776,I981793,I981810,I981827,I981858,I1100827,I981875,I1100836,I981892,I981918,I981940,I981957,I981988,I982033,I982094,I982120,I982137,I982145,I982162,I982179,I982196,I982213,I982230,I982261,I982278,I982309,I982326,I982343,I982374,I982414,I982422,I982439,I982456,I982473,I982504,I982521,I982538,I982564,I982586,I982603,I982634,I982679,I982740,I982766,I982783,I982791,I982808,I982825,I982842,I982859,I982876,I982907,I982924,I982955,I982972,I982989,I983020,I983060,I983068,I983085,I983102,I983119,I983150,I983167,I983184,I983210,I983232,I983249,I983280,I983325,I983386,I983412,I983429,I983437,I983454,I983471,I983488,I983505,I983522,I983553,I983570,I983601,I983618,I983635,I983666,I983706,I983714,I983731,I983748,I983765,I983796,I983813,I983830,I983856,I983878,I983895,I983926,I983971,I984032,I984058,I984075,I984083,I984100,I984117,I984134,I984151,I984168,I984018,I984199,I984216,I984021,I984247,I984264,I984281,I983997,I984312,I984009,I984352,I984360,I984377,I984394,I984411,I984024,I984442,I984459,I984476,I984502,I984012,I984524,I984541,I984006,I984572,I984000,I984003,I984617,I984015,I984678,I1244761,I984704,I1244743,I984721,I984729,I984746,I1244752,I984763,I1244764,I984780,I1244746,I984797,I1244755,I984814,I984845,I984862,I984893,I984910,I1244767,I984927,I984958,I984998,I985006,I985023,I985040,I985057,I985088,I1244749,I985105,I1244758,I985122,I985148,I985170,I985187,I985218,I985263,I985324,I1385673,I985350,I1385697,I985367,I985375,I985392,I1385679,I985409,I1385688,I985426,I985443,I1385694,I985460,I985491,I985508,I985539,I985556,I1385691,I985573,I985604,I985644,I985652,I985669,I985686,I1385685,I985703,I985734,I1385676,I985751,I1385700,I985768,I1385682,I985794,I985816,I985833,I985864,I985909,I985970,I1398763,I985996,I1398787,I986013,I986021,I986038,I1398769,I986055,I1398778,I986072,I986089,I1398784,I986106,I986137,I986154,I986185,I986202,I1398781,I986219,I986250,I986290,I986298,I986315,I986332,I1398775,I986349,I986380,I1398766,I986397,I1398790,I986414,I1398772,I986440,I986462,I986479,I986510,I986555,I986616,I986642,I986659,I986667,I986684,I986701,I986718,I986735,I986752,I986783,I986800,I986831,I986848,I986865,I986896,I986936,I986944,I986961,I986978,I986995,I987026,I987043,I987060,I987086,I987108,I987125,I987156,I987201,I987262,I1403523,I987288,I1403547,I987305,I987313,I987330,I1403529,I987347,I1403538,I987364,I987381,I1403544,I987398,I987429,I987446,I987477,I987494,I1403541,I987511,I987542,I987582,I987590,I987607,I987624,I1403535,I987641,I987672,I1403526,I987689,I1403550,I987706,I1403532,I987732,I987754,I987771,I987802,I987847,I987908,I987934,I987951,I987959,I987976,I987993,I988010,I988027,I988044,I987894,I988075,I988092,I987897,I988123,I988140,I988157,I987873,I988188,I987885,I988228,I988236,I988253,I988270,I988287,I987900,I988318,I988335,I988352,I988378,I987888,I988400,I988417,I987882,I988448,I987876,I987879,I988493,I987891,I988554,I1083685,I988580,I1083688,I988597,I988605,I988622,I988639,I1083697,I988656,I1083706,I988673,I1083694,I988690,I988540,I988721,I988738,I988543,I988769,I988786,I1083700,I988803,I988519,I988834,I988531,I988874,I988882,I988899,I988916,I1083691,I988933,I988546,I988964,I1083703,I988981,I988998,I989024,I988534,I989046,I989063,I988528,I989094,I988522,I988525,I989139,I988537,I989200,I989226,I989243,I989251,I989268,I989285,I989302,I989319,I989336,I989367,I989384,I989415,I989432,I989449,I989480,I989520,I989528,I989545,I989562,I989579,I989610,I989627,I989644,I989670,I989692,I989709,I989740,I989785,I989846,I989872,I989889,I989897,I989914,I989931,I989948,I989965,I989982,I990013,I990030,I990061,I990078,I990095,I990126,I990166,I990174,I990191,I990208,I990225,I990256,I990273,I990290,I990316,I990338,I990355,I990386,I990431,I990492,I990518,I990535,I990543,I990560,I990577,I990594,I990611,I990628,I990659,I990676,I990707,I990724,I990741,I990772,I990812,I990820,I990837,I990854,I990871,I990902,I990919,I990936,I990962,I990984,I991001,I991032,I991077,I991138,I1115867,I991164,I1115849,I991181,I991189,I991206,I1115858,I991223,I1115870,I991240,I1115852,I991257,I1115861,I991274,I991124,I991305,I991322,I991127,I991353,I991370,I1115873,I991387,I991103,I991418,I991115,I991458,I991466,I991483,I991500,I991517,I991130,I991548,I1115855,I991565,I1115864,I991582,I991608,I991118,I991630,I991647,I991112,I991678,I991106,I991109,I991723,I991121,I991784,I991810,I991827,I991835,I991852,I991869,I991886,I991903,I991920,I991951,I991968,I991999,I992016,I992033,I992064,I992104,I992112,I992129,I992146,I992163,I992194,I992211,I992228,I992254,I992276,I992293,I992324,I992369,I992430,I992456,I992473,I992481,I992498,I992515,I992532,I992549,I992566,I992597,I992614,I992645,I992662,I992679,I992710,I992750,I992758,I992775,I992792,I992809,I992840,I992857,I992874,I992900,I992922,I992939,I992970,I993015,I993076,I993102,I993119,I993127,I993144,I993161,I993178,I993195,I993212,I993243,I993260,I993291,I993308,I993325,I993356,I993396,I993404,I993421,I993438,I993455,I993486,I993503,I993520,I993546,I993568,I993585,I993616,I993661,I993722,I993748,I993765,I993773,I993790,I993807,I993824,I993841,I993858,I993889,I993906,I993937,I993954,I993971,I994002,I994042,I994050,I994067,I994084,I994101,I994132,I994149,I994166,I994192,I994214,I994231,I994262,I994307,I994368,I1114711,I994394,I1114693,I994411,I994419,I994436,I1114702,I994453,I1114714,I994470,I1114696,I994487,I1114705,I994504,I994535,I994552,I994583,I994600,I1114717,I994617,I994648,I994688,I994696,I994713,I994730,I994747,I994778,I1114699,I994795,I1114708,I994812,I994838,I994860,I994877,I994908,I994953,I995014,I995040,I995057,I995065,I995082,I995099,I995116,I995133,I995150,I995181,I995198,I995229,I995246,I995263,I995294,I995334,I995342,I995359,I995376,I995393,I995424,I995441,I995458,I995484,I995506,I995523,I995554,I995599,I995660,I995686,I995703,I995711,I995728,I995745,I995762,I995779,I995796,I995827,I995844,I995875,I995892,I995909,I995940,I995980,I995988,I996005,I996022,I996039,I996070,I996087,I996104,I996130,I996152,I996169,I996200,I996245,I996306,I996332,I996349,I996357,I996374,I996391,I996408,I996425,I996442,I996473,I996490,I996521,I996538,I996555,I996586,I996626,I996634,I996651,I996668,I996685,I996716,I996733,I996750,I996776,I996798,I996815,I996846,I996891,I996952,I996978,I996995,I997003,I997020,I997037,I997054,I997071,I997088,I996938,I997119,I997136,I996941,I997167,I997184,I997201,I996917,I997232,I996929,I997272,I997280,I997297,I997314,I997331,I996944,I997362,I997379,I997396,I997422,I996932,I997444,I997461,I996926,I997492,I996920,I996923,I997537,I996935,I997598,I997624,I997641,I997649,I997666,I997683,I997700,I997717,I997734,I997584,I997765,I997782,I997587,I997813,I997830,I997847,I997563,I997878,I997575,I997918,I997926,I997943,I997960,I997977,I997590,I998008,I998025,I998042,I998068,I997578,I998090,I998107,I997572,I998138,I997566,I997569,I998183,I997581,I998244,I998270,I998287,I998295,I998312,I998329,I998346,I998363,I998380,I998411,I998428,I998459,I998476,I998493,I998524,I998564,I998572,I998589,I998606,I998623,I998654,I998671,I998688,I998714,I998736,I998753,I998784,I998829,I998890,I998916,I998933,I998941,I998958,I998975,I998992,I999009,I999026,I998876,I999057,I999074,I998879,I999105,I999122,I999139,I998855,I999170,I998867,I999210,I999218,I999235,I999252,I999269,I998882,I999300,I999317,I999334,I999360,I998870,I999382,I999399,I998864,I999430,I998858,I998861,I999475,I998873,I999536,I999562,I999579,I999587,I999604,I999621,I999638,I999655,I999672,I999522,I999703,I999720,I999525,I999751,I999768,I999785,I999501,I999816,I999513,I999856,I999864,I999881,I999898,I999915,I999528,I999946,I999963,I999980,I1000006,I999516,I1000028,I1000045,I999510,I1000076,I999504,I999507,I1000121,I999519,I1000182,I1000208,I1000225,I1000233,I1000250,I1000267,I1000284,I1000301,I1000318,I1000349,I1000366,I1000397,I1000414,I1000431,I1000462,I1000502,I1000510,I1000527,I1000544,I1000561,I1000592,I1000609,I1000626,I1000652,I1000674,I1000691,I1000722,I1000767,I1000828,I1000854,I1000871,I1000879,I1000896,I1000913,I1000930,I1000947,I1000964,I1000995,I1001012,I1001043,I1001060,I1001077,I1001108,I1001148,I1001156,I1001173,I1001190,I1001207,I1001238,I1001255,I1001272,I1001298,I1001320,I1001337,I1001368,I1001413,I1001474,I1001500,I1001517,I1001525,I1001542,I1001559,I1001576,I1001593,I1001610,I1001641,I1001658,I1001689,I1001706,I1001723,I1001754,I1001794,I1001802,I1001819,I1001836,I1001853,I1001884,I1001901,I1001918,I1001944,I1001966,I1001983,I1002014,I1002059,I1002120,I1002146,I1002163,I1002171,I1002188,I1002205,I1002222,I1002239,I1002256,I1002287,I1002304,I1002335,I1002352,I1002369,I1002400,I1002440,I1002448,I1002465,I1002482,I1002499,I1002530,I1002547,I1002564,I1002590,I1002612,I1002629,I1002660,I1002705,I1002766,I1002792,I1002809,I1002817,I1002834,I1002851,I1002868,I1002885,I1002902,I1002933,I1002950,I1002981,I1002998,I1003015,I1003046,I1003086,I1003094,I1003111,I1003128,I1003145,I1003176,I1003193,I1003210,I1003236,I1003258,I1003275,I1003306,I1003351,I1003412,I1003438,I1003455,I1003463,I1003480,I1003497,I1003514,I1003531,I1003548,I1003579,I1003596,I1003627,I1003644,I1003661,I1003692,I1003732,I1003740,I1003757,I1003774,I1003791,I1003822,I1003839,I1003856,I1003882,I1003904,I1003921,I1003952,I1003997,I1004058,I1004084,I1004101,I1004109,I1004126,I1004143,I1004160,I1004177,I1004194,I1004225,I1004242,I1004273,I1004290,I1004307,I1004338,I1004378,I1004386,I1004403,I1004420,I1004437,I1004468,I1004485,I1004502,I1004528,I1004550,I1004567,I1004598,I1004643,I1004704,I1307992,I1004730,I1307986,I1004747,I1004755,I1004772,I1307995,I1004789,I1308007,I1004806,I1307989,I1004823,I1004840,I1004871,I1004888,I1004919,I1004936,I1307983,I1004953,I1004984,I1005024,I1005032,I1005049,I1005066,I1308004,I1005083,I1005114,I1307998,I1005131,I1005148,I1308001,I1005174,I1005196,I1005213,I1005244,I1005289,I1005350,I1202567,I1005376,I1202549,I1005393,I1005401,I1005418,I1202558,I1005435,I1202570,I1005452,I1202552,I1005469,I1202561,I1005486,I1005517,I1005534,I1005565,I1005582,I1202573,I1005599,I1005630,I1005670,I1005678,I1005695,I1005712,I1005729,I1005760,I1202555,I1005777,I1202564,I1005794,I1005820,I1005842,I1005859,I1005890,I1005935,I1005996,I1006022,I1006039,I1006047,I1006064,I1006081,I1006098,I1006115,I1006132,I1006163,I1006180,I1006211,I1006228,I1006245,I1006276,I1006316,I1006324,I1006341,I1006358,I1006375,I1006406,I1006423,I1006440,I1006466,I1006488,I1006505,I1006536,I1006581,I1006642,I1006668,I1006685,I1006693,I1006710,I1006727,I1006744,I1006761,I1006778,I1006809,I1006826,I1006857,I1006874,I1006891,I1006922,I1006962,I1006970,I1006987,I1007004,I1007021,I1007052,I1007069,I1007086,I1007112,I1007134,I1007151,I1007182,I1007227,I1007288,I1007314,I1007331,I1007339,I1007356,I1007373,I1007390,I1007407,I1007424,I1007455,I1007472,I1007503,I1007520,I1007537,I1007568,I1007608,I1007616,I1007633,I1007650,I1007667,I1007698,I1007715,I1007732,I1007758,I1007780,I1007797,I1007828,I1007873,I1007934,I1007960,I1007977,I1007985,I1008002,I1008019,I1008036,I1008053,I1008070,I1008101,I1008118,I1008149,I1008166,I1008183,I1008214,I1008254,I1008262,I1008279,I1008296,I1008313,I1008344,I1008361,I1008378,I1008404,I1008426,I1008443,I1008474,I1008519,I1008580,I1008606,I1008623,I1008631,I1008648,I1008665,I1008682,I1008699,I1008716,I1008566,I1008747,I1008764,I1008569,I1008795,I1008812,I1008829,I1008545,I1008860,I1008557,I1008900,I1008908,I1008925,I1008942,I1008959,I1008572,I1008990,I1009007,I1009024,I1009050,I1008560,I1009072,I1009089,I1008554,I1009120,I1008548,I1008551,I1009165,I1008563,I1009226,I1078636,I1009252,I1078639,I1009269,I1009277,I1009294,I1009311,I1078648,I1009328,I1078657,I1009345,I1078645,I1009362,I1009393,I1009410,I1009441,I1009458,I1078651,I1009475,I1009506,I1009546,I1009554,I1009571,I1009588,I1078642,I1009605,I1009636,I1078654,I1009653,I1009670,I1009696,I1009718,I1009735,I1009766,I1009811,I1009872,I1009898,I1009915,I1009923,I1009940,I1009957,I1009974,I1009991,I1010008,I1010039,I1010056,I1010087,I1010104,I1010121,I1010152,I1010192,I1010200,I1010217,I1010234,I1010251,I1010282,I1010299,I1010316,I1010342,I1010364,I1010381,I1010412,I1010457,I1010518,I1085368,I1010544,I1085371,I1010561,I1010569,I1010586,I1010603,I1085380,I1010620,I1085389,I1010637,I1085377,I1010654,I1010504,I1010685,I1010702,I1010507,I1010733,I1010750,I1085383,I1010767,I1010483,I1010798,I1010495,I1010838,I1010846,I1010863,I1010880,I1085374,I1010897,I1010510,I1010928,I1085386,I1010945,I1010962,I1010988,I1010498,I1011010,I1011027,I1010492,I1011058,I1010486,I1010489,I1011103,I1010501,I1011164,I1011190,I1011207,I1011215,I1011232,I1011249,I1011266,I1011283,I1011300,I1011331,I1011348,I1011379,I1011396,I1011413,I1011444,I1011484,I1011492,I1011509,I1011526,I1011543,I1011574,I1011591,I1011608,I1011634,I1011656,I1011673,I1011704,I1011749,I1011810,I1011836,I1011853,I1011861,I1011878,I1011895,I1011912,I1011929,I1011946,I1011977,I1011994,I1012025,I1012042,I1012059,I1012090,I1012130,I1012138,I1012155,I1012172,I1012189,I1012220,I1012237,I1012254,I1012280,I1012302,I1012319,I1012350,I1012395,I1012456,I1108931,I1012482,I1108913,I1012499,I1012507,I1012524,I1108922,I1012541,I1108934,I1012558,I1108916,I1012575,I1108925,I1012592,I1012623,I1012640,I1012671,I1012688,I1108937,I1012705,I1012736,I1012776,I1012784,I1012801,I1012818,I1012835,I1012866,I1108919,I1012883,I1108928,I1012900,I1012926,I1012948,I1012965,I1012996,I1013041,I1013102,I1013128,I1013145,I1013153,I1013170,I1013187,I1013204,I1013221,I1013238,I1013269,I1013286,I1013317,I1013334,I1013351,I1013382,I1013422,I1013430,I1013447,I1013464,I1013481,I1013512,I1013529,I1013546,I1013572,I1013594,I1013611,I1013642,I1013687,I1013748,I1013774,I1013791,I1013799,I1013816,I1013833,I1013850,I1013867,I1013884,I1013915,I1013932,I1013963,I1013980,I1013997,I1014028,I1014068,I1014076,I1014093,I1014110,I1014127,I1014158,I1014175,I1014192,I1014218,I1014240,I1014257,I1014288,I1014333,I1014394,I1014420,I1014437,I1014445,I1014462,I1014479,I1014496,I1014513,I1014530,I1014561,I1014578,I1014609,I1014626,I1014643,I1014674,I1014714,I1014722,I1014739,I1014756,I1014773,I1014804,I1014821,I1014838,I1014864,I1014886,I1014903,I1014934,I1014979,I1015040,I1229155,I1015066,I1229137,I1015083,I1015091,I1015108,I1229146,I1015125,I1229158,I1015142,I1229140,I1015159,I1229149,I1015176,I1015207,I1015224,I1015255,I1015272,I1229161,I1015289,I1015320,I1015360,I1015368,I1015385,I1015402,I1015419,I1015450,I1229143,I1015467,I1229152,I1015484,I1015510,I1015532,I1015549,I1015580,I1015625,I1015686,I1015712,I1015729,I1015737,I1015754,I1015771,I1015788,I1015805,I1015822,I1015672,I1015853,I1015870,I1015675,I1015901,I1015918,I1015935,I1015651,I1015966,I1015663,I1016006,I1016014,I1016031,I1016048,I1016065,I1015678,I1016096,I1016113,I1016130,I1016156,I1015666,I1016178,I1016195,I1015660,I1016226,I1015654,I1015657,I1016271,I1015669,I1016332,I1016358,I1016375,I1016383,I1016400,I1016417,I1016434,I1016451,I1016468,I1016318,I1016499,I1016516,I1016321,I1016547,I1016564,I1016581,I1016297,I1016612,I1016309,I1016652,I1016660,I1016677,I1016694,I1016711,I1016324,I1016742,I1016759,I1016776,I1016802,I1016312,I1016824,I1016841,I1016306,I1016872,I1016300,I1016303,I1016917,I1016315,I1016978,I1017004,I1017021,I1017029,I1017046,I1017063,I1017080,I1017097,I1017114,I1016964,I1017145,I1017162,I1016967,I1017193,I1017210,I1017227,I1016943,I1017258,I1016955,I1017298,I1017306,I1017323,I1017340,I1017357,I1016970,I1017388,I1017405,I1017422,I1017448,I1016958,I1017470,I1017487,I1016952,I1017518,I1016946,I1016949,I1017563,I1016961,I1017624,I1147079,I1017650,I1147061,I1017667,I1017675,I1017692,I1147070,I1017709,I1147082,I1017726,I1147064,I1017743,I1147073,I1017760,I1017791,I1017808,I1017839,I1017856,I1147085,I1017873,I1017904,I1017944,I1017952,I1017969,I1017986,I1018003,I1018034,I1147067,I1018051,I1147076,I1018068,I1018094,I1018116,I1018133,I1018164,I1018209,I1018270,I1018296,I1018313,I1018321,I1018338,I1018355,I1018372,I1018389,I1018406,I1018256,I1018437,I1018454,I1018259,I1018485,I1018502,I1018519,I1018235,I1018550,I1018247,I1018590,I1018598,I1018615,I1018632,I1018649,I1018262,I1018680,I1018697,I1018714,I1018740,I1018250,I1018762,I1018779,I1018244,I1018810,I1018238,I1018241,I1018855,I1018253,I1018916,I1018942,I1018959,I1018967,I1018984,I1019001,I1019018,I1019035,I1019052,I1018902,I1019083,I1019100,I1018905,I1019131,I1019148,I1019165,I1018881,I1019196,I1018893,I1019236,I1019244,I1019261,I1019278,I1019295,I1018908,I1019326,I1019343,I1019360,I1019386,I1018896,I1019408,I1019425,I1018890,I1019456,I1018884,I1018887,I1019501,I1018899,I1019562,I1019588,I1019605,I1019613,I1019630,I1019647,I1019664,I1019681,I1019698,I1019729,I1019746,I1019777,I1019794,I1019811,I1019842,I1019882,I1019890,I1019907,I1019924,I1019941,I1019972,I1019989,I1020006,I1020032,I1020054,I1020071,I1020102,I1020147,I1020208,I1217595,I1020234,I1217577,I1020251,I1020259,I1020276,I1217586,I1020293,I1217598,I1020310,I1217580,I1020327,I1217589,I1020344,I1020375,I1020392,I1020423,I1020440,I1217601,I1020457,I1020488,I1020528,I1020536,I1020553,I1020570,I1020587,I1020618,I1217583,I1020635,I1217592,I1020652,I1020678,I1020700,I1020717,I1020748,I1020793,I1020854,I1020880,I1020897,I1020905,I1020922,I1020939,I1020956,I1020973,I1020990,I1020840,I1021021,I1021038,I1020843,I1021069,I1021086,I1021103,I1020819,I1021134,I1020831,I1021174,I1021182,I1021199,I1021216,I1021233,I1020846,I1021264,I1021281,I1021298,I1021324,I1020834,I1021346,I1021363,I1020828,I1021394,I1020822,I1020825,I1021439,I1020837,I1021500,I1061245,I1021526,I1061248,I1021543,I1021551,I1021568,I1021585,I1061257,I1021602,I1061266,I1021619,I1061254,I1021636,I1021486,I1021667,I1021684,I1021489,I1021715,I1021732,I1061260,I1021749,I1021465,I1021780,I1021477,I1021820,I1021828,I1021845,I1021862,I1061251,I1021879,I1021492,I1021910,I1061263,I1021927,I1021944,I1021970,I1021480,I1021992,I1022009,I1021474,I1022040,I1021468,I1021471,I1022085,I1021483,I1022146,I1114133,I1022172,I1114115,I1022189,I1022197,I1022214,I1114124,I1022231,I1114136,I1022248,I1114118,I1022265,I1114127,I1022282,I1022313,I1022330,I1022361,I1022378,I1114139,I1022395,I1022426,I1022466,I1022474,I1022491,I1022508,I1022525,I1022556,I1114121,I1022573,I1114130,I1022590,I1022616,I1022638,I1022655,I1022686,I1022731,I1022792,I1022818,I1022835,I1022843,I1022860,I1022877,I1022894,I1022911,I1022928,I1022959,I1022976,I1023007,I1023024,I1023041,I1023072,I1023112,I1023120,I1023137,I1023154,I1023171,I1023202,I1023219,I1023236,I1023262,I1023284,I1023301,I1023332,I1023377,I1023438,I1023464,I1023481,I1023489,I1023506,I1023523,I1023540,I1023557,I1023574,I1023605,I1023622,I1023653,I1023670,I1023687,I1023718,I1023758,I1023766,I1023783,I1023800,I1023817,I1023848,I1023865,I1023882,I1023908,I1023930,I1023947,I1023978,I1024023,I1024084,I1024110,I1024127,I1024135,I1024152,I1024169,I1024186,I1024203,I1024220,I1024251,I1024268,I1024299,I1024316,I1024333,I1024364,I1024404,I1024412,I1024429,I1024446,I1024463,I1024494,I1024511,I1024528,I1024554,I1024576,I1024593,I1024624,I1024669,I1024730,I1024756,I1024773,I1024781,I1024798,I1024815,I1024832,I1024849,I1024866,I1024897,I1024914,I1024945,I1024962,I1024979,I1025010,I1025050,I1025058,I1025075,I1025092,I1025109,I1025140,I1025157,I1025174,I1025200,I1025222,I1025239,I1025270,I1025315,I1025376,I1025402,I1025419,I1025427,I1025444,I1025461,I1025478,I1025495,I1025512,I1025543,I1025560,I1025591,I1025608,I1025625,I1025656,I1025696,I1025704,I1025721,I1025738,I1025755,I1025786,I1025803,I1025820,I1025846,I1025868,I1025885,I1025916,I1025961,I1026022,I1026048,I1026065,I1026073,I1026090,I1026107,I1026124,I1026141,I1026158,I1026189,I1026206,I1026237,I1026254,I1026271,I1026302,I1026342,I1026350,I1026367,I1026384,I1026401,I1026432,I1026449,I1026466,I1026492,I1026514,I1026531,I1026562,I1026607,I1026668,I1026694,I1026711,I1026719,I1026736,I1026753,I1026770,I1026787,I1026804,I1026654,I1026835,I1026852,I1026657,I1026883,I1026900,I1026917,I1026633,I1026948,I1026645,I1026988,I1026996,I1027013,I1027030,I1027047,I1026660,I1027078,I1027095,I1027112,I1027138,I1026648,I1027160,I1027177,I1026642,I1027208,I1026636,I1026639,I1027253,I1026651,I1027314,I1027340,I1027357,I1027365,I1027382,I1027399,I1027416,I1027433,I1027450,I1027300,I1027481,I1027498,I1027303,I1027529,I1027546,I1027563,I1027279,I1027594,I1027291,I1027634,I1027642,I1027659,I1027676,I1027693,I1027306,I1027724,I1027741,I1027758,I1027784,I1027294,I1027806,I1027823,I1027288,I1027854,I1027282,I1027285,I1027899,I1027297,I1027960,I1362468,I1027986,I1362492,I1028003,I1028011,I1028028,I1362474,I1028045,I1362483,I1028062,I1028079,I1362489,I1028096,I1028127,I1028144,I1028175,I1028192,I1362486,I1028209,I1028240,I1028280,I1028288,I1028305,I1028322,I1362480,I1028339,I1028370,I1362471,I1028387,I1362495,I1028404,I1362477,I1028430,I1028452,I1028469,I1028500,I1028545,I1028606,I1177713,I1028632,I1177695,I1028649,I1028657,I1028674,I1177704,I1028691,I1177716,I1028708,I1177698,I1028725,I1177707,I1028742,I1028773,I1028790,I1028821,I1028838,I1177719,I1028855,I1028886,I1028926,I1028934,I1028951,I1028968,I1028985,I1029016,I1177701,I1029033,I1177710,I1029050,I1029076,I1029098,I1029115,I1029146,I1029191,I1029252,I1029278,I1029295,I1029303,I1029320,I1029337,I1029354,I1029371,I1029388,I1029238,I1029419,I1029436,I1029241,I1029467,I1029484,I1029501,I1029217,I1029532,I1029229,I1029572,I1029580,I1029597,I1029614,I1029631,I1029244,I1029662,I1029679,I1029696,I1029722,I1029232,I1029744,I1029761,I1029226,I1029792,I1029220,I1029223,I1029837,I1029235,I1029898,I1029924,I1029941,I1029949,I1029966,I1029983,I1030000,I1030017,I1030034,I1030065,I1030082,I1030113,I1030130,I1030147,I1030178,I1030218,I1030226,I1030243,I1030260,I1030277,I1030308,I1030325,I1030342,I1030368,I1030390,I1030407,I1030438,I1030483,I1030544,I1030570,I1030587,I1030595,I1030612,I1030629,I1030646,I1030663,I1030680,I1030530,I1030711,I1030728,I1030533,I1030759,I1030776,I1030793,I1030509,I1030824,I1030521,I1030864,I1030872,I1030889,I1030906,I1030923,I1030536,I1030954,I1030971,I1030988,I1031014,I1030524,I1031036,I1031053,I1030518,I1031084,I1030512,I1030515,I1031129,I1030527,I1031190,I1395788,I1031216,I1395812,I1031233,I1031241,I1031258,I1395794,I1031275,I1395803,I1031292,I1031309,I1395809,I1031326,I1031357,I1031374,I1031405,I1031422,I1395806,I1031439,I1031470,I1031510,I1031518,I1031535,I1031552,I1395800,I1031569,I1031600,I1395791,I1031617,I1395815,I1031634,I1395797,I1031660,I1031682,I1031699,I1031730,I1031775,I1031836,I1031862,I1031879,I1031887,I1031904,I1031921,I1031938,I1031955,I1031972,I1032003,I1032020,I1032051,I1032068,I1032085,I1032116,I1032156,I1032164,I1032181,I1032198,I1032215,I1032246,I1032263,I1032280,I1032306,I1032328,I1032345,I1032376,I1032421,I1032482,I1032508,I1032525,I1032533,I1032550,I1032567,I1032584,I1032601,I1032618,I1032649,I1032666,I1032697,I1032714,I1032731,I1032762,I1032802,I1032810,I1032827,I1032844,I1032861,I1032892,I1032909,I1032926,I1032952,I1032974,I1032991,I1033022,I1033067,I1033128,I1033154,I1033171,I1033179,I1033196,I1033213,I1033230,I1033247,I1033264,I1033114,I1033295,I1033312,I1033117,I1033343,I1033360,I1033377,I1033093,I1033408,I1033105,I1033448,I1033456,I1033473,I1033490,I1033507,I1033120,I1033538,I1033555,I1033572,I1033598,I1033108,I1033620,I1033637,I1033102,I1033668,I1033096,I1033099,I1033713,I1033111,I1033774,I1033800,I1033817,I1033825,I1033842,I1033859,I1033876,I1033893,I1033910,I1033760,I1033941,I1033958,I1033763,I1033989,I1034006,I1034023,I1033739,I1034054,I1033751,I1034094,I1034102,I1034119,I1034136,I1034153,I1033766,I1034184,I1034201,I1034218,I1034244,I1033754,I1034266,I1034283,I1033748,I1034314,I1033742,I1033745,I1034359,I1033757,I1034420,I1034446,I1034463,I1034471,I1034488,I1034505,I1034522,I1034539,I1034556,I1034587,I1034604,I1034635,I1034652,I1034669,I1034700,I1034740,I1034748,I1034765,I1034782,I1034799,I1034830,I1034847,I1034864,I1034890,I1034912,I1034929,I1034960,I1035005,I1035066,I1035092,I1035109,I1035117,I1035134,I1035151,I1035168,I1035185,I1035202,I1035233,I1035250,I1035281,I1035298,I1035315,I1035346,I1035386,I1035394,I1035411,I1035428,I1035445,I1035476,I1035493,I1035510,I1035536,I1035558,I1035575,I1035606,I1035651,I1035712,I1035738,I1035755,I1035763,I1035780,I1035797,I1035814,I1035831,I1035848,I1035879,I1035896,I1035927,I1035944,I1035961,I1035992,I1036032,I1036040,I1036057,I1036074,I1036091,I1036122,I1036139,I1036156,I1036182,I1036204,I1036221,I1036252,I1036297,I1036358,I1036384,I1036401,I1036409,I1036426,I1036443,I1036460,I1036477,I1036494,I1036344,I1036525,I1036542,I1036347,I1036573,I1036590,I1036607,I1036323,I1036638,I1036335,I1036678,I1036686,I1036703,I1036720,I1036737,I1036350,I1036768,I1036785,I1036802,I1036828,I1036338,I1036850,I1036867,I1036332,I1036898,I1036326,I1036329,I1036943,I1036341,I1037004,I1037030,I1037047,I1037055,I1037072,I1037089,I1037106,I1037123,I1037140,I1037171,I1037188,I1037219,I1037236,I1037253,I1037284,I1037324,I1037332,I1037349,I1037366,I1037383,I1037414,I1037431,I1037448,I1037474,I1037496,I1037513,I1037544,I1037589,I1037650,I1214127,I1037676,I1214109,I1037693,I1037701,I1037718,I1214118,I1037735,I1214130,I1037752,I1214112,I1037769,I1214121,I1037786,I1037636,I1037817,I1037834,I1037639,I1037865,I1037882,I1214133,I1037899,I1037615,I1037930,I1037627,I1037970,I1037978,I1037995,I1038012,I1038029,I1037642,I1038060,I1214115,I1038077,I1214124,I1038094,I1038120,I1037630,I1038142,I1038159,I1037624,I1038190,I1037618,I1037621,I1038235,I1037633,I1038296,I1038322,I1038339,I1038347,I1038364,I1038381,I1038398,I1038415,I1038432,I1038463,I1038480,I1038511,I1038528,I1038545,I1038576,I1038616,I1038624,I1038641,I1038658,I1038675,I1038706,I1038723,I1038740,I1038766,I1038788,I1038805,I1038836,I1038881,I1038942,I1038968,I1038985,I1038993,I1039010,I1039027,I1039044,I1039061,I1039078,I1039109,I1039126,I1039157,I1039174,I1039191,I1039222,I1039262,I1039270,I1039287,I1039304,I1039321,I1039352,I1039369,I1039386,I1039412,I1039434,I1039451,I1039482,I1039527,I1039588,I1039614,I1039631,I1039639,I1039656,I1039673,I1039690,I1039707,I1039724,I1039574,I1039755,I1039772,I1039577,I1039803,I1039820,I1039837,I1039553,I1039868,I1039565,I1039908,I1039916,I1039933,I1039950,I1039967,I1039580,I1039998,I1040015,I1040032,I1040058,I1039568,I1040080,I1040097,I1039562,I1040128,I1039556,I1039559,I1040173,I1039571,I1040234,I1040260,I1040277,I1040285,I1040302,I1040319,I1040336,I1040353,I1040370,I1040401,I1040418,I1040449,I1040466,I1040483,I1040514,I1040554,I1040562,I1040579,I1040596,I1040613,I1040644,I1040661,I1040678,I1040704,I1040726,I1040743,I1040774,I1040819,I1040880,I1040906,I1040923,I1040931,I1040948,I1040965,I1040982,I1040999,I1041016,I1040866,I1041047,I1041064,I1040869,I1041095,I1041112,I1041129,I1040845,I1041160,I1040857,I1041200,I1041208,I1041225,I1041242,I1041259,I1040872,I1041290,I1041307,I1041324,I1041350,I1040860,I1041372,I1041389,I1040854,I1041420,I1040848,I1040851,I1041465,I1040863,I1041526,I1041552,I1041569,I1041577,I1041594,I1041611,I1041628,I1041645,I1041662,I1041512,I1041693,I1041710,I1041515,I1041741,I1041758,I1041775,I1041491,I1041806,I1041503,I1041846,I1041854,I1041871,I1041888,I1041905,I1041518,I1041936,I1041953,I1041970,I1041996,I1041506,I1042018,I1042035,I1041500,I1042066,I1041494,I1041497,I1042111,I1041509,I1042172,I1042198,I1042215,I1042223,I1042240,I1042257,I1042274,I1042291,I1042308,I1042339,I1042356,I1042387,I1042404,I1042421,I1042452,I1042492,I1042500,I1042517,I1042534,I1042551,I1042582,I1042599,I1042616,I1042642,I1042664,I1042681,I1042712,I1042757,I1042818,I1042844,I1042861,I1042869,I1042886,I1042903,I1042920,I1042937,I1042954,I1042985,I1043002,I1043033,I1043050,I1043067,I1043098,I1043138,I1043146,I1043163,I1043180,I1043197,I1043228,I1043245,I1043262,I1043288,I1043310,I1043327,I1043358,I1043403,I1043464,I1043490,I1043507,I1043515,I1043532,I1043549,I1043566,I1043583,I1043600,I1043631,I1043648,I1043679,I1043696,I1043713,I1043744,I1043784,I1043792,I1043809,I1043826,I1043843,I1043874,I1043891,I1043908,I1043934,I1043956,I1043973,I1044004,I1044049,I1044110,I1044136,I1044153,I1044161,I1044178,I1044195,I1044212,I1044229,I1044246,I1044277,I1044294,I1044325,I1044342,I1044359,I1044390,I1044430,I1044438,I1044455,I1044472,I1044489,I1044520,I1044537,I1044554,I1044580,I1044602,I1044619,I1044650,I1044695,I1044756,I1044782,I1044799,I1044807,I1044824,I1044841,I1044858,I1044875,I1044892,I1044742,I1044923,I1044940,I1044745,I1044971,I1044988,I1045005,I1044721,I1045036,I1044733,I1045076,I1045084,I1045101,I1045118,I1045135,I1044748,I1045166,I1045183,I1045200,I1045226,I1044736,I1045248,I1045265,I1044730,I1045296,I1044724,I1044727,I1045341,I1044739,I1045402,I1116445,I1045428,I1116427,I1045445,I1045453,I1045470,I1116436,I1045487,I1116448,I1045504,I1116430,I1045521,I1116439,I1045538,I1045569,I1045586,I1045617,I1045634,I1116451,I1045651,I1045682,I1045722,I1045730,I1045747,I1045764,I1045781,I1045812,I1116433,I1045829,I1116442,I1045846,I1045872,I1045894,I1045911,I1045942,I1045987,I1046048,I1046074,I1046091,I1046099,I1046116,I1046133,I1046150,I1046167,I1046184,I1046215,I1046232,I1046263,I1046280,I1046297,I1046328,I1046368,I1046376,I1046393,I1046410,I1046427,I1046458,I1046475,I1046492,I1046518,I1046540,I1046557,I1046588,I1046633,I1046688,I1046714,I1046731,I1046753,I1046779,I1046787,I1046804,I1046821,I1046838,I1046855,I1046872,I1046889,I1046920,I1046951,I1046968,I1046985,I1047002,I1047033,I1047078,I1047095,I1047112,I1047138,I1047146,I1047177,I1047194,I1047249,I1047275,I1047292,I1047314,I1047340,I1047348,I1047365,I1047382,I1047399,I1047416,I1047433,I1047450,I1047481,I1047512,I1047529,I1047546,I1047563,I1047594,I1047639,I1047656,I1047673,I1047699,I1047707,I1047738,I1047755,I1047810,I1404728,I1047836,I1047853,I1047802,I1047875,I1404722,I1047901,I1047909,I1404713,I1047926,I1047943,I1404740,I1047960,I1404725,I1404734,I1047977,I1047994,I1404719,I1048011,I1047784,I1048042,I1047787,I1048073,I1404737,I1048090,I1048107,I1048124,I1047796,I1048155,I1047799,I1047793,I1048200,I1404731,I1048217,I1048234,I1404716,I1048260,I1048268,I1047781,I1048299,I1048316,I1047790,I1048371,I1048397,I1048414,I1048436,I1048462,I1048470,I1048487,I1048504,I1048521,I1048538,I1048555,I1048572,I1048603,I1048634,I1048651,I1048668,I1048685,I1048716,I1048761,I1048778,I1048795,I1048821,I1048829,I1048860,I1048877,I1048932,I1048958,I1048975,I1048997,I1049023,I1049031,I1049048,I1049065,I1049082,I1049099,I1049116,I1049133,I1049164,I1049195,I1049212,I1049229,I1049246,I1049277,I1049322,I1049339,I1049356,I1049382,I1049390,I1049421,I1049438,I1049493,I1049519,I1049536,I1049558,I1049584,I1049592,I1049609,I1049626,I1049643,I1049660,I1049677,I1049694,I1049725,I1049756,I1049773,I1049790,I1049807,I1049838,I1049883,I1049900,I1049917,I1049943,I1049951,I1049982,I1049999,I1050054,I1050080,I1050097,I1050046,I1050119,I1050145,I1050153,I1050170,I1050187,I1050204,I1050221,I1050238,I1050255,I1050028,I1050286,I1050031,I1050317,I1050334,I1050351,I1050368,I1050040,I1050399,I1050043,I1050037,I1050444,I1050461,I1050478,I1050504,I1050512,I1050025,I1050543,I1050560,I1050034,I1050615,I1260015,I1050641,I1050658,I1050680,I1260021,I1050706,I1050714,I1260030,I1050731,I1050748,I1260009,I1050765,I1260012,I1050782,I1050799,I1260024,I1050816,I1050847,I1050878,I1260018,I1050895,I1050912,I1050929,I1050960,I1051005,I1260033,I1051022,I1051039,I1260027,I1051065,I1051073,I1051104,I1051121,I1051176,I1051202,I1051219,I1051241,I1051267,I1051275,I1051292,I1051309,I1051326,I1051343,I1051360,I1051377,I1051408,I1051439,I1051456,I1051473,I1051490,I1051521,I1051566,I1051583,I1051600,I1051626,I1051634,I1051665,I1051682,I1051737,I1051763,I1051780,I1051802,I1051828,I1051836,I1051853,I1051870,I1051887,I1051904,I1051921,I1051938,I1051969,I1052000,I1052017,I1052034,I1052051,I1052082,I1052127,I1052144,I1052161,I1052187,I1052195,I1052226,I1052243,I1052298,I1286127,I1052324,I1052341,I1052363,I1286133,I1052389,I1052397,I1286142,I1052414,I1052431,I1286121,I1052448,I1286124,I1052465,I1052482,I1286136,I1052499,I1052530,I1052561,I1286130,I1052578,I1052595,I1052612,I1052643,I1052688,I1286145,I1052705,I1052722,I1286139,I1052748,I1052756,I1052787,I1052804,I1052859,I1181756,I1052885,I1052902,I1052851,I1052924,I1181747,I1052950,I1052958,I1181744,I1052975,I1052992,I1181753,I1053009,I1181762,I1053026,I1053043,I1181741,I1053060,I1052833,I1053091,I1052836,I1053122,I1181750,I1053139,I1053156,I1053173,I1052845,I1053204,I1052848,I1052842,I1053249,I1181765,I1053266,I1053283,I1181759,I1053309,I1053317,I1052830,I1053348,I1053365,I1052839,I1053420,I1111818,I1053446,I1053463,I1053485,I1111809,I1053511,I1053519,I1111806,I1053536,I1053553,I1111815,I1053570,I1111824,I1053587,I1053604,I1111803,I1053621,I1053652,I1053683,I1111812,I1053700,I1053717,I1053734,I1053765,I1053810,I1111827,I1053827,I1053844,I1111821,I1053870,I1053878,I1053909,I1053926,I1053981,I1054007,I1054024,I1054046,I1054072,I1054080,I1054097,I1054114,I1054131,I1054148,I1054165,I1054182,I1054213,I1054244,I1054261,I1054278,I1054295,I1054326,I1054371,I1054388,I1054405,I1054431,I1054439,I1054470,I1054487,I1054542,I1054568,I1054585,I1054607,I1054633,I1054641,I1054658,I1054675,I1054692,I1054709,I1054726,I1054743,I1054774,I1054805,I1054822,I1054839,I1054856,I1054887,I1054932,I1054949,I1054966,I1054992,I1055000,I1055031,I1055048,I1055103,I1055129,I1055146,I1055095,I1055168,I1055194,I1055202,I1055219,I1055236,I1055253,I1055270,I1055287,I1055304,I1055077,I1055335,I1055080,I1055366,I1055383,I1055400,I1055417,I1055089,I1055448,I1055092,I1055086,I1055493,I1055510,I1055527,I1055553,I1055561,I1055074,I1055592,I1055609,I1055083,I1055664,I1055690,I1055707,I1055729,I1055755,I1055763,I1055780,I1055797,I1055814,I1055831,I1055848,I1055865,I1055896,I1055927,I1055944,I1055961,I1055978,I1056009,I1056054,I1056071,I1056088,I1056114,I1056122,I1056153,I1056170,I1056225,I1056251,I1056268,I1056290,I1056316,I1056324,I1056341,I1056358,I1056375,I1056392,I1056409,I1056426,I1056457,I1056488,I1056505,I1056522,I1056539,I1056570,I1056615,I1056632,I1056649,I1056675,I1056683,I1056714,I1056731,I1056786,I1056812,I1056829,I1056851,I1056877,I1056885,I1056902,I1056919,I1056936,I1056953,I1056970,I1056987,I1057018,I1057049,I1057066,I1057083,I1057100,I1057131,I1057176,I1057193,I1057210,I1057236,I1057244,I1057275,I1057292,I1057347,I1057373,I1057390,I1057412,I1057438,I1057446,I1057463,I1057480,I1057497,I1057514,I1057531,I1057548,I1057579,I1057610,I1057627,I1057644,I1057661,I1057692,I1057737,I1057754,I1057771,I1057797,I1057805,I1057836,I1057853,I1057908,I1057934,I1057951,I1057973,I1057999,I1058007,I1058024,I1058041,I1058058,I1058075,I1058092,I1058109,I1058140,I1058171,I1058188,I1058205,I1058222,I1058253,I1058298,I1058315,I1058332,I1058358,I1058366,I1058397,I1058414,I1058469,I1058495,I1058512,I1058534,I1058560,I1058568,I1058585,I1058602,I1058619,I1058636,I1058653,I1058670,I1058701,I1058732,I1058749,I1058766,I1058783,I1058814,I1058859,I1058876,I1058893,I1058919,I1058927,I1058958,I1058975,I1059030,I1059056,I1059073,I1059095,I1059121,I1059129,I1059146,I1059163,I1059180,I1059197,I1059214,I1059231,I1059262,I1059293,I1059310,I1059327,I1059344,I1059375,I1059420,I1059437,I1059454,I1059480,I1059488,I1059519,I1059536,I1059591,I1332733,I1059617,I1059634,I1059583,I1059656,I1332727,I1059682,I1059690,I1332718,I1059707,I1059724,I1332745,I1059741,I1332730,I1332739,I1059758,I1059775,I1332724,I1059792,I1059565,I1059823,I1059568,I1059854,I1332742,I1059871,I1059888,I1059905,I1059577,I1059936,I1059580,I1059574,I1059981,I1332736,I1059998,I1060015,I1332721,I1060041,I1060049,I1059562,I1060080,I1060097,I1059571,I1060152,I1342848,I1060178,I1060195,I1060144,I1060217,I1342842,I1060243,I1060251,I1342833,I1060268,I1060285,I1342860,I1060302,I1342845,I1342854,I1060319,I1060336,I1342839,I1060353,I1060126,I1060384,I1060129,I1060415,I1342857,I1060432,I1060449,I1060466,I1060138,I1060497,I1060141,I1060135,I1060542,I1342851,I1060559,I1060576,I1342836,I1060602,I1060610,I1060123,I1060641,I1060658,I1060132,I1060713,I1060739,I1060756,I1060778,I1060804,I1060812,I1060829,I1060846,I1060863,I1060880,I1060897,I1060914,I1060945,I1060976,I1060993,I1061010,I1061027,I1061058,I1061103,I1061120,I1061137,I1061163,I1061171,I1061202,I1061219,I1061274,I1061300,I1061317,I1061339,I1061365,I1061373,I1061390,I1061407,I1061424,I1061441,I1061458,I1061475,I1061506,I1061537,I1061554,I1061571,I1061588,I1061619,I1061664,I1061681,I1061698,I1061724,I1061732,I1061763,I1061780,I1061835,I1061861,I1061878,I1061900,I1061926,I1061934,I1061951,I1061968,I1061985,I1062002,I1062019,I1062036,I1062067,I1062098,I1062115,I1062132,I1062149,I1062180,I1062225,I1062242,I1062259,I1062285,I1062293,I1062324,I1062341,I1062396,I1062422,I1062439,I1062461,I1062487,I1062495,I1062512,I1062529,I1062546,I1062563,I1062580,I1062597,I1062628,I1062659,I1062676,I1062693,I1062710,I1062741,I1062786,I1062803,I1062820,I1062846,I1062854,I1062885,I1062902,I1062957,I1062983,I1063000,I1062949,I1063022,I1063048,I1063056,I1063073,I1063090,I1063107,I1063124,I1063141,I1063158,I1062931,I1063189,I1062934,I1063220,I1063237,I1063254,I1063271,I1062943,I1063302,I1062946,I1062940,I1063347,I1063364,I1063381,I1063407,I1063415,I1062928,I1063446,I1063463,I1062937,I1063518,I1063544,I1063561,I1063510,I1063583,I1063609,I1063617,I1063634,I1063651,I1063668,I1063685,I1063702,I1063719,I1063492,I1063750,I1063495,I1063781,I1063798,I1063815,I1063832,I1063504,I1063863,I1063507,I1063501,I1063908,I1063925,I1063942,I1063968,I1063976,I1063489,I1064007,I1064024,I1063498,I1064079,I1064105,I1064122,I1064144,I1064170,I1064178,I1064195,I1064212,I1064229,I1064246,I1064263,I1064280,I1064311,I1064342,I1064359,I1064376,I1064393,I1064424,I1064469,I1064486,I1064503,I1064529,I1064537,I1064568,I1064585,I1064640,I1064666,I1064683,I1064705,I1064731,I1064739,I1064756,I1064773,I1064790,I1064807,I1064824,I1064841,I1064872,I1064903,I1064920,I1064937,I1064954,I1064985,I1065030,I1065047,I1065064,I1065090,I1065098,I1065129,I1065146,I1065201,I1065227,I1065244,I1065266,I1065292,I1065300,I1065317,I1065334,I1065351,I1065368,I1065385,I1065402,I1065433,I1065464,I1065481,I1065498,I1065515,I1065546,I1065591,I1065608,I1065625,I1065651,I1065659,I1065690,I1065707,I1065762,I1065788,I1065805,I1065827,I1065853,I1065861,I1065878,I1065895,I1065912,I1065929,I1065946,I1065963,I1065994,I1066025,I1066042,I1066059,I1066076,I1066107,I1066152,I1066169,I1066186,I1066212,I1066220,I1066251,I1066268,I1066323,I1066349,I1066366,I1066388,I1066414,I1066422,I1066439,I1066456,I1066473,I1066490,I1066507,I1066524,I1066555,I1066586,I1066603,I1066620,I1066637,I1066668,I1066713,I1066730,I1066747,I1066773,I1066781,I1066812,I1066829,I1066884,I1066910,I1066927,I1066949,I1066975,I1066983,I1067000,I1067017,I1067034,I1067051,I1067068,I1067085,I1067116,I1067147,I1067164,I1067181,I1067198,I1067229,I1067274,I1067291,I1067308,I1067334,I1067342,I1067373,I1067390,I1067445,I1067471,I1067488,I1067510,I1067536,I1067544,I1067561,I1067578,I1067595,I1067612,I1067629,I1067646,I1067677,I1067708,I1067725,I1067742,I1067759,I1067790,I1067835,I1067852,I1067869,I1067895,I1067903,I1067934,I1067951,I1068006,I1068032,I1068049,I1068071,I1068097,I1068105,I1068122,I1068139,I1068156,I1068173,I1068190,I1068207,I1068238,I1068269,I1068286,I1068303,I1068320,I1068351,I1068396,I1068413,I1068430,I1068456,I1068464,I1068495,I1068512,I1068567,I1068593,I1068610,I1068632,I1068658,I1068666,I1068683,I1068700,I1068717,I1068734,I1068751,I1068768,I1068799,I1068830,I1068847,I1068864,I1068881,I1068912,I1068957,I1068974,I1068991,I1069017,I1069025,I1069056,I1069073,I1069128,I1069154,I1069171,I1069120,I1069193,I1069219,I1069227,I1069244,I1069261,I1069278,I1069295,I1069312,I1069329,I1069102,I1069360,I1069105,I1069391,I1069408,I1069425,I1069442,I1069114,I1069473,I1069117,I1069111,I1069518,I1069535,I1069552,I1069578,I1069586,I1069099,I1069617,I1069634,I1069108,I1069689,I1221638,I1069715,I1069732,I1069754,I1221629,I1069780,I1069788,I1221626,I1069805,I1069822,I1221635,I1069839,I1221644,I1069856,I1069873,I1221623,I1069890,I1069921,I1069952,I1221632,I1069969,I1069986,I1070003,I1070034,I1070079,I1221647,I1070096,I1070113,I1221641,I1070139,I1070147,I1070178,I1070195,I1070250,I1070276,I1070293,I1070315,I1070341,I1070349,I1070366,I1070383,I1070400,I1070417,I1070434,I1070451,I1070482,I1070513,I1070530,I1070547,I1070564,I1070595,I1070640,I1070657,I1070674,I1070700,I1070708,I1070739,I1070756,I1070811,I1070837,I1070854,I1070876,I1070902,I1070910,I1070927,I1070944,I1070961,I1070978,I1070995,I1071012,I1071043,I1071074,I1071091,I1071108,I1071125,I1071156,I1071201,I1071218,I1071235,I1071261,I1071269,I1071300,I1071317,I1071372,I1237244,I1071398,I1071415,I1071437,I1237235,I1071463,I1071471,I1237232,I1071488,I1071505,I1237241,I1071522,I1237250,I1071539,I1071556,I1237229,I1071573,I1071604,I1071635,I1237238,I1071652,I1071669,I1071686,I1071717,I1071762,I1237253,I1071779,I1071796,I1237247,I1071822,I1071830,I1071861,I1071878,I1071933,I1071959,I1071976,I1071998,I1072024,I1072032,I1072049,I1072066,I1072083,I1072100,I1072117,I1072134,I1072165,I1072196,I1072213,I1072230,I1072247,I1072278,I1072323,I1072340,I1072357,I1072383,I1072391,I1072422,I1072439,I1072494,I1072520,I1072537,I1072559,I1072585,I1072593,I1072610,I1072627,I1072644,I1072661,I1072678,I1072695,I1072726,I1072757,I1072774,I1072791,I1072808,I1072839,I1072884,I1072901,I1072918,I1072944,I1072952,I1072983,I1073000,I1073055,I1073081,I1073098,I1073047,I1073120,I1073146,I1073154,I1073171,I1073188,I1073205,I1073222,I1073239,I1073256,I1073029,I1073287,I1073032,I1073318,I1073335,I1073352,I1073369,I1073041,I1073400,I1073044,I1073038,I1073445,I1073462,I1073479,I1073505,I1073513,I1073026,I1073544,I1073561,I1073035,I1073616,I1073642,I1073659,I1073681,I1073707,I1073715,I1073732,I1073749,I1073766,I1073783,I1073800,I1073817,I1073848,I1073879,I1073896,I1073913,I1073930,I1073961,I1074006,I1074023,I1074040,I1074066,I1074074,I1074105,I1074122,I1074177,I1360698,I1074203,I1074220,I1074242,I1360692,I1074268,I1074276,I1360683,I1074293,I1074310,I1360710,I1074327,I1360695,I1360704,I1074344,I1074361,I1360689,I1074378,I1074409,I1074440,I1360707,I1074457,I1074474,I1074491,I1074522,I1074567,I1360701,I1074584,I1074601,I1360686,I1074627,I1074635,I1074666,I1074683,I1074738,I1074764,I1074781,I1074803,I1074829,I1074837,I1074854,I1074871,I1074888,I1074905,I1074922,I1074939,I1074970,I1075001,I1075018,I1075035,I1075052,I1075083,I1075128,I1075145,I1075162,I1075188,I1075196,I1075227,I1075244,I1075299,I1075325,I1075342,I1075291,I1075364,I1075390,I1075398,I1075415,I1075432,I1075449,I1075466,I1075483,I1075500,I1075273,I1075531,I1075276,I1075562,I1075579,I1075596,I1075613,I1075285,I1075644,I1075288,I1075282,I1075689,I1075706,I1075723,I1075749,I1075757,I1075270,I1075788,I1075805,I1075279,I1075860,I1075886,I1075903,I1075925,I1075951,I1075959,I1075976,I1075993,I1076010,I1076027,I1076044,I1076061,I1076092,I1076123,I1076140,I1076157,I1076174,I1076205,I1076250,I1076267,I1076284,I1076310,I1076318,I1076349,I1076366,I1076421,I1076447,I1076464,I1076486,I1076512,I1076520,I1076537,I1076554,I1076571,I1076588,I1076605,I1076622,I1076653,I1076684,I1076701,I1076718,I1076735,I1076766,I1076811,I1076828,I1076845,I1076871,I1076879,I1076910,I1076927,I1076982,I1077008,I1077025,I1077047,I1077073,I1077081,I1077098,I1077115,I1077132,I1077149,I1077166,I1077183,I1077214,I1077245,I1077262,I1077279,I1077296,I1077327,I1077372,I1077389,I1077406,I1077432,I1077440,I1077471,I1077488,I1077543,I1077569,I1077586,I1077535,I1077608,I1077634,I1077642,I1077659,I1077676,I1077693,I1077710,I1077727,I1077744,I1077517,I1077775,I1077520,I1077806,I1077823,I1077840,I1077857,I1077529,I1077888,I1077532,I1077526,I1077933,I1077950,I1077967,I1077993,I1078001,I1077514,I1078032,I1078049,I1077523,I1078104,I1078130,I1078147,I1078169,I1078195,I1078203,I1078220,I1078237,I1078254,I1078271,I1078288,I1078305,I1078336,I1078367,I1078384,I1078401,I1078418,I1078449,I1078494,I1078511,I1078528,I1078554,I1078562,I1078593,I1078610,I1078665,I1078691,I1078708,I1078730,I1078756,I1078764,I1078781,I1078798,I1078815,I1078832,I1078849,I1078866,I1078897,I1078928,I1078945,I1078962,I1078979,I1079010,I1079055,I1079072,I1079089,I1079115,I1079123,I1079154,I1079171,I1079226,I1277423,I1079252,I1079269,I1079291,I1277429,I1079317,I1079325,I1277438,I1079342,I1079359,I1277417,I1079376,I1277420,I1079393,I1079410,I1277432,I1079427,I1079458,I1079489,I1277426,I1079506,I1079523,I1079540,I1079571,I1079616,I1277441,I1079633,I1079650,I1277435,I1079676,I1079684,I1079715,I1079732,I1079787,I1092744,I1079813,I1079830,I1079779,I1079852,I1092735,I1079878,I1079886,I1092732,I1079903,I1079920,I1092741,I1079937,I1092750,I1079954,I1079971,I1092729,I1079988,I1079761,I1080019,I1079764,I1080050,I1092738,I1080067,I1080084,I1080101,I1079773,I1080132,I1079776,I1079770,I1080177,I1092753,I1080194,I1080211,I1092747,I1080237,I1080245,I1079758,I1080276,I1080293,I1079767,I1080348,I1080374,I1080391,I1080413,I1080439,I1080447,I1080464,I1080481,I1080498,I1080515,I1080532,I1080549,I1080580,I1080611,I1080628,I1080645,I1080662,I1080693,I1080738,I1080755,I1080772,I1080798,I1080806,I1080837,I1080854,I1080909,I1080935,I1080952,I1080974,I1081000,I1081008,I1081025,I1081042,I1081059,I1081076,I1081093,I1081110,I1081141,I1081172,I1081189,I1081206,I1081223,I1081254,I1081299,I1081316,I1081333,I1081359,I1081367,I1081398,I1081415,I1081470,I1081496,I1081513,I1081535,I1081561,I1081569,I1081586,I1081603,I1081620,I1081637,I1081654,I1081671,I1081702,I1081733,I1081750,I1081767,I1081784,I1081815,I1081860,I1081877,I1081894,I1081920,I1081928,I1081959,I1081976,I1082031,I1328115,I1082057,I1082074,I1082096,I1328100,I1082122,I1082130,I1328109,I1082147,I1082164,I1328103,I1082181,I1328121,I1328118,I1082198,I1082215,I1328094,I1082232,I1082263,I1082294,I1328097,I1082311,I1082328,I1082345,I1082376,I1082421,I1082438,I1328112,I1082455,I1328106,I1082481,I1082489,I1082520,I1082537,I1082592,I1082618,I1082635,I1082584,I1082657,I1082683,I1082691,I1082708,I1082725,I1082742,I1082759,I1082776,I1082793,I1082566,I1082824,I1082569,I1082855,I1082872,I1082889,I1082906,I1082578,I1082937,I1082581,I1082575,I1082982,I1082999,I1083016,I1083042,I1083050,I1082563,I1083081,I1083098,I1082572,I1083153,I1083179,I1083196,I1083218,I1083244,I1083252,I1083269,I1083286,I1083303,I1083320,I1083337,I1083354,I1083385,I1083416,I1083433,I1083450,I1083467,I1083498,I1083543,I1083560,I1083577,I1083603,I1083611,I1083642,I1083659,I1083714,I1083740,I1083757,I1083779,I1083805,I1083813,I1083830,I1083847,I1083864,I1083881,I1083898,I1083915,I1083946,I1083977,I1083994,I1084011,I1084028,I1084059,I1084104,I1084121,I1084138,I1084164,I1084172,I1084203,I1084220,I1084275,I1084301,I1084318,I1084340,I1084366,I1084374,I1084391,I1084408,I1084425,I1084442,I1084459,I1084476,I1084507,I1084538,I1084555,I1084572,I1084589,I1084620,I1084665,I1084682,I1084699,I1084725,I1084733,I1084764,I1084781,I1084836,I1084862,I1084879,I1084901,I1084927,I1084935,I1084952,I1084969,I1084986,I1085003,I1085020,I1085037,I1085068,I1085099,I1085116,I1085133,I1085150,I1085181,I1085226,I1085243,I1085260,I1085286,I1085294,I1085325,I1085342,I1085397,I1085423,I1085440,I1085462,I1085488,I1085496,I1085513,I1085530,I1085547,I1085564,I1085581,I1085598,I1085629,I1085660,I1085677,I1085694,I1085711,I1085742,I1085787,I1085804,I1085821,I1085847,I1085855,I1085886,I1085903,I1085958,I1117598,I1085984,I1086001,I1086023,I1117589,I1086049,I1086057,I1117586,I1086074,I1086091,I1117595,I1086108,I1117604,I1086125,I1086142,I1117583,I1086159,I1086190,I1086221,I1117592,I1086238,I1086255,I1086272,I1086303,I1086348,I1117607,I1086365,I1086382,I1117601,I1086408,I1086416,I1086447,I1086464,I1086519,I1086545,I1086562,I1086584,I1086610,I1086618,I1086635,I1086652,I1086669,I1086686,I1086703,I1086720,I1086751,I1086782,I1086799,I1086816,I1086833,I1086864,I1086909,I1086926,I1086943,I1086969,I1086977,I1087008,I1087025,I1087080,I1215280,I1087106,I1087123,I1087145,I1215271,I1087171,I1087179,I1215268,I1087196,I1087213,I1215277,I1087230,I1215286,I1087247,I1087264,I1215265,I1087281,I1087312,I1087343,I1215274,I1087360,I1087377,I1087394,I1087425,I1087470,I1215289,I1087487,I1087504,I1215283,I1087530,I1087538,I1087569,I1087586,I1087641,I1087667,I1087684,I1087706,I1087732,I1087740,I1087757,I1087774,I1087791,I1087808,I1087825,I1087842,I1087873,I1087904,I1087921,I1087938,I1087955,I1087986,I1088031,I1088048,I1088065,I1088091,I1088099,I1088130,I1088147,I1088202,I1088228,I1088245,I1088267,I1088293,I1088301,I1088318,I1088335,I1088352,I1088369,I1088386,I1088403,I1088434,I1088465,I1088482,I1088499,I1088516,I1088547,I1088592,I1088609,I1088626,I1088652,I1088660,I1088691,I1088708,I1088763,I1088789,I1088806,I1088828,I1088854,I1088862,I1088879,I1088896,I1088913,I1088930,I1088947,I1088964,I1088995,I1089026,I1089043,I1089060,I1089077,I1089108,I1089153,I1089170,I1089187,I1089213,I1089221,I1089252,I1089269,I1089324,I1089350,I1089367,I1089389,I1089415,I1089423,I1089440,I1089457,I1089474,I1089491,I1089508,I1089525,I1089556,I1089587,I1089604,I1089621,I1089638,I1089669,I1089714,I1089731,I1089748,I1089774,I1089782,I1089813,I1089830,I1089885,I1089911,I1089928,I1089877,I1089950,I1089976,I1089984,I1090001,I1090018,I1090035,I1090052,I1090069,I1090086,I1089859,I1090117,I1089862,I1090148,I1090165,I1090182,I1090199,I1089871,I1090230,I1089874,I1089868,I1090275,I1090292,I1090309,I1090335,I1090343,I1089856,I1090374,I1090391,I1089865,I1090449,I1090475,I1090483,I1090523,I1090531,I1090548,I1090565,I1090605,I1090627,I1090644,I1090670,I1090678,I1090695,I1090712,I1090729,I1090746,I1090791,I1090822,I1090839,I1090865,I1090873,I1090904,I1090921,I1090938,I1090955,I1091027,I1091053,I1091061,I1091101,I1091109,I1091126,I1091143,I1091183,I1091205,I1091222,I1091248,I1091256,I1091273,I1091290,I1091307,I1091324,I1091369,I1091400,I1091417,I1091443,I1091451,I1091482,I1091499,I1091516,I1091533,I1091605,I1091631,I1091639,I1091679,I1091687,I1091704,I1091721,I1091761,I1091783,I1091800,I1091826,I1091834,I1091851,I1091868,I1091885,I1091902,I1091947,I1091978,I1091995,I1092021,I1092029,I1092060,I1092077,I1092094,I1092111,I1092183,I1092209,I1092217,I1092257,I1092265,I1092282,I1092299,I1092339,I1092361,I1092378,I1092404,I1092412,I1092429,I1092446,I1092463,I1092480,I1092525,I1092556,I1092573,I1092599,I1092607,I1092638,I1092655,I1092672,I1092689,I1092761,I1092787,I1092795,I1092835,I1092843,I1092860,I1092877,I1092917,I1092939,I1092956,I1092982,I1092990,I1093007,I1093024,I1093041,I1093058,I1093103,I1093134,I1093151,I1093177,I1093185,I1093216,I1093233,I1093250,I1093267,I1093339,I1093365,I1093373,I1093413,I1093421,I1093438,I1093455,I1093495,I1093517,I1093534,I1093560,I1093568,I1093585,I1093602,I1093619,I1093636,I1093681,I1093712,I1093729,I1093755,I1093763,I1093794,I1093811,I1093828,I1093845,I1093917,I1093943,I1093951,I1093991,I1093999,I1094016,I1094033,I1094073,I1094095,I1094112,I1094138,I1094146,I1094163,I1094180,I1094197,I1094214,I1094259,I1094290,I1094307,I1094333,I1094341,I1094372,I1094389,I1094406,I1094423,I1094495,I1094521,I1094529,I1094569,I1094577,I1094594,I1094611,I1094651,I1094673,I1094690,I1094716,I1094724,I1094741,I1094758,I1094775,I1094792,I1094837,I1094868,I1094885,I1094911,I1094919,I1094950,I1094967,I1094984,I1095001,I1095073,I1328655,I1095099,I1095107,I1328682,I1328664,I1095147,I1095155,I1328673,I1095172,I1328676,I1095189,I1095229,I1095251,I1328670,I1095268,I1095294,I1095302,I1095319,I1328658,I1095336,I1328661,I1095353,I1095370,I1095415,I1328679,I1095446,I1095463,I1328667,I1095489,I1095497,I1095528,I1095545,I1095562,I1095579,I1095651,I1095677,I1095685,I1095725,I1095733,I1095750,I1095767,I1095807,I1095829,I1095846,I1095872,I1095880,I1095897,I1095914,I1095931,I1095948,I1095993,I1096024,I1096041,I1096067,I1096075,I1096106,I1096123,I1096140,I1096157,I1096229,I1324167,I1096255,I1096263,I1324194,I1324176,I1096303,I1096311,I1324185,I1096328,I1324188,I1096345,I1096385,I1096407,I1324182,I1096424,I1096450,I1096458,I1096475,I1324170,I1096492,I1324173,I1096509,I1096526,I1096571,I1324191,I1096602,I1096619,I1324179,I1096645,I1096653,I1096684,I1096701,I1096718,I1096735,I1096807,I1096833,I1096841,I1096881,I1096889,I1096906,I1096923,I1096963,I1096985,I1097002,I1097028,I1097036,I1097053,I1097070,I1097087,I1097104,I1097149,I1097180,I1097197,I1097223,I1097231,I1097262,I1097279,I1097296,I1097313,I1097385,I1269278,I1097411,I1097419,I1269272,I1269257,I1097459,I1097467,I1269263,I1097484,I1269275,I1097501,I1097541,I1097563,I1097580,I1097606,I1097614,I1097631,I1269281,I1097648,I1269269,I1097665,I1097682,I1097727,I1269260,I1097758,I1097775,I1269266,I1097801,I1097809,I1097840,I1097857,I1097874,I1097891,I1097963,I1097989,I1097997,I1098037,I1098045,I1098062,I1098079,I1098119,I1098141,I1098158,I1098184,I1098192,I1098209,I1098226,I1098243,I1098260,I1098305,I1098336,I1098353,I1098379,I1098387,I1098418,I1098435,I1098452,I1098469,I1098541,I1098567,I1098575,I1098615,I1098623,I1098640,I1098657,I1098697,I1098719,I1098736,I1098762,I1098770,I1098787,I1098804,I1098821,I1098838,I1098883,I1098914,I1098931,I1098957,I1098965,I1098996,I1099013,I1099030,I1099047,I1099119,I1099145,I1099153,I1099193,I1099201,I1099218,I1099235,I1099275,I1099297,I1099314,I1099340,I1099348,I1099365,I1099382,I1099399,I1099416,I1099461,I1099492,I1099509,I1099535,I1099543,I1099574,I1099591,I1099608,I1099625,I1099697,I1099723,I1099731,I1099680,I1099771,I1099779,I1099796,I1099813,I1099668,I1099853,I1099689,I1099875,I1099892,I1099918,I1099926,I1099943,I1099960,I1099977,I1099994,I1099665,I1099686,I1100039,I1099677,I1100070,I1100087,I1100113,I1100121,I1099683,I1100152,I1100169,I1100186,I1100203,I1099674,I1099671,I1100275,I1100301,I1100309,I1100349,I1100357,I1100374,I1100391,I1100431,I1100453,I1100470,I1100496,I1100504,I1100521,I1100538,I1100555,I1100572,I1100617,I1100648,I1100665,I1100691,I1100699,I1100730,I1100747,I1100764,I1100781,I1100853,I1100879,I1100887,I1100927,I1100935,I1100952,I1100969,I1101009,I1101031,I1101048,I1101074,I1101082,I1101099,I1101116,I1101133,I1101150,I1101195,I1101226,I1101243,I1101269,I1101277,I1101308,I1101325,I1101342,I1101359,I1101431,I1101457,I1101465,I1101505,I1101513,I1101530,I1101547,I1101587,I1101609,I1101626,I1101652,I1101660,I1101677,I1101694,I1101711,I1101728,I1101773,I1101804,I1101821,I1101847,I1101855,I1101886,I1101903,I1101920,I1101937,I1102009,I1102035,I1102043,I1102083,I1102091,I1102108,I1102125,I1102165,I1102187,I1102204,I1102230,I1102238,I1102255,I1102272,I1102289,I1102306,I1102351,I1102382,I1102399,I1102425,I1102433,I1102464,I1102481,I1102498,I1102515,I1102587,I1102613,I1102621,I1102661,I1102669,I1102686,I1102703,I1102743,I1102765,I1102782,I1102808,I1102816,I1102833,I1102850,I1102867,I1102884,I1102929,I1102960,I1102977,I1103003,I1103011,I1103042,I1103059,I1103076,I1103093,I1103165,I1103191,I1103199,I1103239,I1103247,I1103264,I1103281,I1103321,I1103343,I1103360,I1103386,I1103394,I1103411,I1103428,I1103445,I1103462,I1103507,I1103538,I1103555,I1103581,I1103589,I1103620,I1103637,I1103654,I1103671,I1103743,I1103769,I1103777,I1103817,I1103825,I1103842,I1103859,I1103899,I1103921,I1103938,I1103964,I1103972,I1103989,I1104006,I1104023,I1104040,I1104085,I1104116,I1104133,I1104159,I1104167,I1104198,I1104215,I1104232,I1104249,I1104321,I1104347,I1104355,I1104395,I1104403,I1104420,I1104437,I1104477,I1104499,I1104516,I1104542,I1104550,I1104567,I1104584,I1104601,I1104618,I1104663,I1104694,I1104711,I1104737,I1104745,I1104776,I1104793,I1104810,I1104827,I1104899,I1104925,I1104933,I1104973,I1104981,I1104998,I1105015,I1105055,I1105077,I1105094,I1105120,I1105128,I1105145,I1105162,I1105179,I1105196,I1105241,I1105272,I1105289,I1105315,I1105323,I1105354,I1105371,I1105388,I1105405,I1105477,I1105503,I1105511,I1105460,I1105551,I1105559,I1105576,I1105593,I1105448,I1105633,I1105469,I1105655,I1105672,I1105698,I1105706,I1105723,I1105740,I1105757,I1105774,I1105445,I1105466,I1105819,I1105457,I1105850,I1105867,I1105893,I1105901,I1105463,I1105932,I1105949,I1105966,I1105983,I1105454,I1105451,I1106055,I1335125,I1106081,I1106089,I1335107,I1335098,I1106129,I1106137,I1335113,I1106154,I1335101,I1106171,I1106211,I1106233,I1335110,I1106250,I1106276,I1106284,I1106301,I1335119,I1106318,I1106335,I1106352,I1106397,I1335122,I1106428,I1106445,I1335116,I1335104,I1106471,I1106479,I1106510,I1106527,I1106544,I1106561,I1106633,I1106659,I1106667,I1106707,I1106715,I1106732,I1106749,I1106789,I1106811,I1106828,I1106854,I1106862,I1106879,I1106896,I1106913,I1106930,I1106975,I1107006,I1107023,I1107049,I1107057,I1107088,I1107105,I1107122,I1107139,I1107211,I1107237,I1107245,I1107285,I1107293,I1107310,I1107327,I1107367,I1107389,I1107406,I1107432,I1107440,I1107457,I1107474,I1107491,I1107508,I1107553,I1107584,I1107601,I1107627,I1107635,I1107666,I1107683,I1107700,I1107717,I1107789,I1393435,I1107815,I1107823,I1393417,I1393408,I1107863,I1107871,I1393423,I1107888,I1393411,I1107905,I1107945,I1107967,I1393420,I1107984,I1108010,I1108018,I1108035,I1393429,I1108052,I1108069,I1108086,I1108131,I1393432,I1108162,I1108179,I1393426,I1393414,I1108205,I1108213,I1108244,I1108261,I1108278,I1108295,I1108367,I1108393,I1108401,I1108350,I1108441,I1108449,I1108466,I1108483,I1108338,I1108523,I1108359,I1108545,I1108562,I1108588,I1108596,I1108613,I1108630,I1108647,I1108664,I1108335,I1108356,I1108709,I1108347,I1108740,I1108757,I1108783,I1108791,I1108353,I1108822,I1108839,I1108856,I1108873,I1108344,I1108341,I1108945,I1108971,I1108979,I1109019,I1109027,I1109044,I1109061,I1109101,I1109123,I1109140,I1109166,I1109174,I1109191,I1109208,I1109225,I1109242,I1109287,I1109318,I1109335,I1109361,I1109369,I1109400,I1109417,I1109434,I1109451,I1109523,I1109549,I1109557,I1109597,I1109605,I1109622,I1109639,I1109679,I1109701,I1109718,I1109744,I1109752,I1109769,I1109786,I1109803,I1109820,I1109865,I1109896,I1109913,I1109939,I1109947,I1109978,I1109995,I1110012,I1110029,I1110101,I1110127,I1110135,I1110175,I1110183,I1110200,I1110217,I1110257,I1110279,I1110296,I1110322,I1110330,I1110347,I1110364,I1110381,I1110398,I1110443,I1110474,I1110491,I1110517,I1110525,I1110556,I1110573,I1110590,I1110607,I1110679,I1110705,I1110713,I1110662,I1110753,I1110761,I1110778,I1110795,I1110650,I1110835,I1110671,I1110857,I1110874,I1110900,I1110908,I1110925,I1110942,I1110959,I1110976,I1110647,I1110668,I1111021,I1110659,I1111052,I1111069,I1111095,I1111103,I1110665,I1111134,I1111151,I1111168,I1111185,I1110656,I1110653,I1111257,I1111283,I1111291,I1111331,I1111339,I1111356,I1111373,I1111413,I1111435,I1111452,I1111478,I1111486,I1111503,I1111520,I1111537,I1111554,I1111599,I1111630,I1111647,I1111673,I1111681,I1111712,I1111729,I1111746,I1111763,I1111835,I1111861,I1111869,I1111909,I1111917,I1111934,I1111951,I1111991,I1112013,I1112030,I1112056,I1112064,I1112081,I1112098,I1112115,I1112132,I1112177,I1112208,I1112225,I1112251,I1112259,I1112290,I1112307,I1112324,I1112341,I1112413,I1347620,I1112439,I1112447,I1347602,I1347593,I1112487,I1112495,I1347608,I1112512,I1347596,I1112529,I1112569,I1112591,I1347605,I1112608,I1112634,I1112642,I1112659,I1347614,I1112676,I1112693,I1112710,I1112755,I1347617,I1112786,I1112803,I1347611,I1347599,I1112829,I1112837,I1112868,I1112885,I1112902,I1112919,I1112991,I1113017,I1113025,I1113065,I1113073,I1113090,I1113107,I1113147,I1113169,I1113186,I1113212,I1113220,I1113237,I1113254,I1113271,I1113288,I1113333,I1113364,I1113381,I1113407,I1113415,I1113446,I1113463,I1113480,I1113497,I1113569,I1113595,I1113603,I1113552,I1113643,I1113651,I1113668,I1113685,I1113540,I1113725,I1113561,I1113747,I1113764,I1113790,I1113798,I1113815,I1113832,I1113849,I1113866,I1113537,I1113558,I1113911,I1113549,I1113942,I1113959,I1113985,I1113993,I1113555,I1114024,I1114041,I1114058,I1114075,I1113546,I1113543,I1114147,I1114173,I1114181,I1114221,I1114229,I1114246,I1114263,I1114303,I1114325,I1114342,I1114368,I1114376,I1114393,I1114410,I1114427,I1114444,I1114489,I1114520,I1114537,I1114563,I1114571,I1114602,I1114619,I1114636,I1114653,I1114725,I1114751,I1114759,I1114799,I1114807,I1114824,I1114841,I1114881,I1114903,I1114920,I1114946,I1114954,I1114971,I1114988,I1115005,I1115022,I1115067,I1115098,I1115115,I1115141,I1115149,I1115180,I1115197,I1115214,I1115231,I1115303,I1115329,I1115337,I1115377,I1115385,I1115402,I1115419,I1115459,I1115481,I1115498,I1115524,I1115532,I1115549,I1115566,I1115583,I1115600,I1115645,I1115676,I1115693,I1115719,I1115727,I1115758,I1115775,I1115792,I1115809,I1115881,I1115907,I1115915,I1115955,I1115963,I1115980,I1115997,I1116037,I1116059,I1116076,I1116102,I1116110,I1116127,I1116144,I1116161,I1116178,I1116223,I1116254,I1116271,I1116297,I1116305,I1116336,I1116353,I1116370,I1116387,I1116459,I1116485,I1116493,I1116533,I1116541,I1116558,I1116575,I1116615,I1116637,I1116654,I1116680,I1116688,I1116705,I1116722,I1116739,I1116756,I1116801,I1116832,I1116849,I1116875,I1116883,I1116914,I1116931,I1116948,I1116965,I1117037,I1117063,I1117071,I1117111,I1117119,I1117136,I1117153,I1117193,I1117215,I1117232,I1117258,I1117266,I1117283,I1117300,I1117317,I1117334,I1117379,I1117410,I1117427,I1117453,I1117461,I1117492,I1117509,I1117526,I1117543,I1117615,I1345240,I1117641,I1117649,I1345222,I1345213,I1117689,I1117697,I1345228,I1117714,I1345216,I1117731,I1117771,I1117793,I1345225,I1117810,I1117836,I1117844,I1117861,I1345234,I1117878,I1117895,I1117912,I1117957,I1345237,I1117988,I1118005,I1345231,I1345219,I1118031,I1118039,I1118070,I1118087,I1118104,I1118121,I1118193,I1118219,I1118227,I1118267,I1118275,I1118292,I1118309,I1118349,I1118371,I1118388,I1118414,I1118422,I1118439,I1118456,I1118473,I1118490,I1118535,I1118566,I1118583,I1118609,I1118617,I1118648,I1118665,I1118682,I1118699,I1118771,I1118797,I1118805,I1118845,I1118853,I1118870,I1118887,I1118927,I1118949,I1118966,I1118992,I1119000,I1119017,I1119034,I1119051,I1119068,I1119113,I1119144,I1119161,I1119187,I1119195,I1119226,I1119243,I1119260,I1119277,I1119349,I1119375,I1119383,I1119423,I1119431,I1119448,I1119465,I1119505,I1119527,I1119544,I1119570,I1119578,I1119595,I1119612,I1119629,I1119646,I1119691,I1119722,I1119739,I1119765,I1119773,I1119804,I1119821,I1119838,I1119855,I1119927,I1256766,I1119953,I1119961,I1256760,I1256745,I1120001,I1120009,I1256751,I1120026,I1256763,I1120043,I1120083,I1120105,I1120122,I1120148,I1120156,I1120173,I1256769,I1120190,I1256757,I1120207,I1120224,I1120269,I1256748,I1120300,I1120317,I1256754,I1120343,I1120351,I1120382,I1120399,I1120416,I1120433,I1120505,I1348215,I1120531,I1120539,I1348197,I1348188,I1120579,I1120587,I1348203,I1120604,I1348191,I1120621,I1120661,I1120683,I1348200,I1120700,I1120726,I1120734,I1120751,I1348209,I1120768,I1120785,I1120802,I1120847,I1348212,I1120878,I1120895,I1348206,I1348194,I1120921,I1120929,I1120960,I1120977,I1120994,I1121011,I1121083,I1121109,I1121117,I1121066,I1121157,I1121165,I1121182,I1121199,I1121054,I1121239,I1121075,I1121261,I1121278,I1121304,I1121312,I1121329,I1121346,I1121363,I1121380,I1121051,I1121072,I1121425,I1121063,I1121456,I1121473,I1121499,I1121507,I1121069,I1121538,I1121555,I1121572,I1121589,I1121060,I1121057,I1121661,I1121687,I1121695,I1121644,I1121735,I1121743,I1121760,I1121777,I1121632,I1121817,I1121653,I1121839,I1121856,I1121882,I1121890,I1121907,I1121924,I1121941,I1121958,I1121629,I1121650,I1122003,I1121641,I1122034,I1122051,I1122077,I1122085,I1121647,I1122116,I1122133,I1122150,I1122167,I1121638,I1121635,I1122239,I1122265,I1122273,I1122313,I1122321,I1122338,I1122355,I1122395,I1122417,I1122434,I1122460,I1122468,I1122485,I1122502,I1122519,I1122536,I1122581,I1122612,I1122629,I1122655,I1122663,I1122694,I1122711,I1122728,I1122745,I1122817,I1377965,I1122843,I1122851,I1377947,I1377938,I1122891,I1122899,I1377953,I1122916,I1377941,I1122933,I1122973,I1122995,I1377950,I1123012,I1123038,I1123046,I1123063,I1377959,I1123080,I1123097,I1123114,I1123159,I1377962,I1123190,I1123207,I1377956,I1377944,I1123233,I1123241,I1123272,I1123289,I1123306,I1123323,I1123395,I1123421,I1123429,I1123469,I1123477,I1123494,I1123511,I1123551,I1123573,I1123590,I1123616,I1123624,I1123641,I1123658,I1123675,I1123692,I1123737,I1123768,I1123785,I1123811,I1123819,I1123850,I1123867,I1123884,I1123901,I1123973,I1123999,I1124007,I1124047,I1124055,I1124072,I1124089,I1124129,I1124151,I1124168,I1124194,I1124202,I1124219,I1124236,I1124253,I1124270,I1124315,I1124346,I1124363,I1124389,I1124397,I1124428,I1124445,I1124462,I1124479,I1124551,I1124577,I1124585,I1124625,I1124633,I1124650,I1124667,I1124707,I1124729,I1124746,I1124772,I1124780,I1124797,I1124814,I1124831,I1124848,I1124893,I1124924,I1124941,I1124967,I1124975,I1125006,I1125023,I1125040,I1125057,I1125129,I1125155,I1125163,I1125203,I1125211,I1125228,I1125245,I1125285,I1125307,I1125324,I1125350,I1125358,I1125375,I1125392,I1125409,I1125426,I1125471,I1125502,I1125519,I1125545,I1125553,I1125584,I1125601,I1125618,I1125635,I1125707,I1292401,I1125733,I1125741,I1292383,I1292392,I1125781,I1125789,I1292377,I1125806,I1292389,I1125823,I1125863,I1125885,I1292380,I1125902,I1125928,I1125936,I1125953,I1125970,I1125987,I1126004,I1126049,I1292398,I1126080,I1126097,I1292386,I1292395,I1126123,I1126131,I1126162,I1126179,I1126196,I1126213,I1126285,I1126311,I1126319,I1126359,I1126367,I1126384,I1126401,I1126441,I1126463,I1126480,I1126506,I1126514,I1126531,I1126548,I1126565,I1126582,I1126627,I1126658,I1126675,I1126701,I1126709,I1126740,I1126757,I1126774,I1126791,I1126863,I1126889,I1126897,I1126937,I1126945,I1126962,I1126979,I1127019,I1127041,I1127058,I1127084,I1127092,I1127109,I1127126,I1127143,I1127160,I1127205,I1127236,I1127253,I1127279,I1127287,I1127318,I1127335,I1127352,I1127369,I1127441,I1127467,I1127475,I1127515,I1127523,I1127540,I1127557,I1127597,I1127619,I1127636,I1127662,I1127670,I1127687,I1127704,I1127721,I1127738,I1127783,I1127814,I1127831,I1127857,I1127865,I1127896,I1127913,I1127930,I1127947,I1128019,I1128045,I1128053,I1128093,I1128101,I1128118,I1128135,I1128175,I1128197,I1128214,I1128240,I1128248,I1128265,I1128282,I1128299,I1128316,I1128361,I1128392,I1128409,I1128435,I1128443,I1128474,I1128491,I1128508,I1128525,I1128597,I1128623,I1128631,I1128671,I1128679,I1128696,I1128713,I1128753,I1128775,I1128792,I1128818,I1128826,I1128843,I1128860,I1128877,I1128894,I1128939,I1128970,I1128987,I1129013,I1129021,I1129052,I1129069,I1129086,I1129103,I1129175,I1129201,I1129209,I1129249,I1129257,I1129274,I1129291,I1129331,I1129353,I1129370,I1129396,I1129404,I1129421,I1129438,I1129455,I1129472,I1129517,I1129548,I1129565,I1129591,I1129599,I1129630,I1129647,I1129664,I1129681,I1129753,I1129779,I1129787,I1129827,I1129835,I1129852,I1129869,I1129909,I1129931,I1129948,I1129974,I1129982,I1129999,I1130016,I1130033,I1130050,I1130095,I1130126,I1130143,I1130169,I1130177,I1130208,I1130225,I1130242,I1130259,I1130331,I1130357,I1130365,I1130405,I1130413,I1130430,I1130447,I1130487,I1130509,I1130526,I1130552,I1130560,I1130577,I1130594,I1130611,I1130628,I1130673,I1130704,I1130721,I1130747,I1130755,I1130786,I1130803,I1130820,I1130837,I1130909,I1130935,I1130943,I1130983,I1130991,I1131008,I1131025,I1131065,I1131087,I1131104,I1131130,I1131138,I1131155,I1131172,I1131189,I1131206,I1131251,I1131282,I1131299,I1131325,I1131333,I1131364,I1131381,I1131398,I1131415,I1131487,I1131513,I1131521,I1131561,I1131569,I1131586,I1131603,I1131643,I1131665,I1131682,I1131708,I1131716,I1131733,I1131750,I1131767,I1131784,I1131829,I1131860,I1131877,I1131903,I1131911,I1131942,I1131959,I1131976,I1131993,I1132065,I1132091,I1132099,I1132139,I1132147,I1132164,I1132181,I1132221,I1132243,I1132260,I1132286,I1132294,I1132311,I1132328,I1132345,I1132362,I1132407,I1132438,I1132455,I1132481,I1132489,I1132520,I1132537,I1132554,I1132571,I1132643,I1132669,I1132677,I1132717,I1132725,I1132742,I1132759,I1132799,I1132821,I1132838,I1132864,I1132872,I1132889,I1132906,I1132923,I1132940,I1132985,I1133016,I1133033,I1133059,I1133067,I1133098,I1133115,I1133132,I1133149,I1133221,I1133247,I1133255,I1133295,I1133303,I1133320,I1133337,I1133377,I1133399,I1133416,I1133442,I1133450,I1133467,I1133484,I1133501,I1133518,I1133563,I1133594,I1133611,I1133637,I1133645,I1133676,I1133693,I1133710,I1133727,I1133799,I1133825,I1133833,I1133782,I1133873,I1133881,I1133898,I1133915,I1133770,I1133955,I1133791,I1133977,I1133994,I1134020,I1134028,I1134045,I1134062,I1134079,I1134096,I1133767,I1133788,I1134141,I1133779,I1134172,I1134189,I1134215,I1134223,I1133785,I1134254,I1134271,I1134288,I1134305,I1133776,I1133773,I1134377,I1134403,I1134411,I1134451,I1134459,I1134476,I1134493,I1134533,I1134555,I1134572,I1134598,I1134606,I1134623,I1134640,I1134657,I1134674,I1134719,I1134750,I1134767,I1134793,I1134801,I1134832,I1134849,I1134866,I1134883,I1134955,I1134981,I1134989,I1135029,I1135037,I1135054,I1135071,I1135111,I1135133,I1135150,I1135176,I1135184,I1135201,I1135218,I1135235,I1135252,I1135297,I1135328,I1135345,I1135371,I1135379,I1135410,I1135427,I1135444,I1135461,I1135533,I1135559,I1135567,I1135607,I1135615,I1135632,I1135649,I1135689,I1135711,I1135728,I1135754,I1135762,I1135779,I1135796,I1135813,I1135830,I1135875,I1135906,I1135923,I1135949,I1135957,I1135988,I1136005,I1136022,I1136039,I1136111,I1136137,I1136145,I1136185,I1136193,I1136210,I1136227,I1136267,I1136289,I1136306,I1136332,I1136340,I1136357,I1136374,I1136391,I1136408,I1136453,I1136484,I1136501,I1136527,I1136535,I1136566,I1136583,I1136600,I1136617,I1136689,I1136715,I1136723,I1136763,I1136771,I1136788,I1136805,I1136845,I1136867,I1136884,I1136910,I1136918,I1136935,I1136952,I1136969,I1136986,I1137031,I1137062,I1137079,I1137105,I1137113,I1137144,I1137161,I1137178,I1137195,I1137267,I1137293,I1137301,I1137341,I1137349,I1137366,I1137383,I1137423,I1137445,I1137462,I1137488,I1137496,I1137513,I1137530,I1137547,I1137564,I1137609,I1137640,I1137657,I1137683,I1137691,I1137722,I1137739,I1137756,I1137773,I1137845,I1137871,I1137879,I1137919,I1137927,I1137944,I1137961,I1138001,I1138023,I1138040,I1138066,I1138074,I1138091,I1138108,I1138125,I1138142,I1138187,I1138218,I1138235,I1138261,I1138269,I1138300,I1138317,I1138334,I1138351,I1138423,I1138449,I1138457,I1138497,I1138505,I1138522,I1138539,I1138579,I1138601,I1138618,I1138644,I1138652,I1138669,I1138686,I1138703,I1138720,I1138765,I1138796,I1138813,I1138839,I1138847,I1138878,I1138895,I1138912,I1138929,I1139001,I1139027,I1139035,I1139075,I1139083,I1139100,I1139117,I1139157,I1139179,I1139196,I1139222,I1139230,I1139247,I1139264,I1139281,I1139298,I1139343,I1139374,I1139391,I1139417,I1139425,I1139456,I1139473,I1139490,I1139507,I1139579,I1407120,I1139605,I1139613,I1407102,I1139562,I1407093,I1139653,I1139661,I1407108,I1139678,I1407096,I1139695,I1139550,I1139735,I1139571,I1139757,I1407105,I1139774,I1139800,I1139808,I1139825,I1407114,I1139842,I1139859,I1139876,I1139547,I1139568,I1139921,I1407117,I1139559,I1139952,I1139969,I1407111,I1407099,I1139995,I1140003,I1139565,I1140034,I1140051,I1140068,I1140085,I1139556,I1139553,I1140157,I1140183,I1140191,I1140231,I1140239,I1140256,I1140273,I1140313,I1140335,I1140352,I1140378,I1140386,I1140403,I1140420,I1140437,I1140454,I1140499,I1140530,I1140547,I1140573,I1140581,I1140612,I1140629,I1140646,I1140663,I1140735,I1140761,I1140769,I1140809,I1140817,I1140834,I1140851,I1140891,I1140913,I1140930,I1140956,I1140964,I1140981,I1140998,I1141015,I1141032,I1141077,I1141108,I1141125,I1141151,I1141159,I1141190,I1141207,I1141224,I1141241,I1141313,I1141339,I1141347,I1141387,I1141395,I1141412,I1141429,I1141469,I1141491,I1141508,I1141534,I1141542,I1141559,I1141576,I1141593,I1141610,I1141655,I1141686,I1141703,I1141729,I1141737,I1141768,I1141785,I1141802,I1141819,I1141891,I1141917,I1141925,I1141965,I1141973,I1141990,I1142007,I1142047,I1142069,I1142086,I1142112,I1142120,I1142137,I1142154,I1142171,I1142188,I1142233,I1142264,I1142281,I1142307,I1142315,I1142346,I1142363,I1142380,I1142397,I1142469,I1142495,I1142503,I1142452,I1142543,I1142551,I1142568,I1142585,I1142440,I1142625,I1142461,I1142647,I1142664,I1142690,I1142698,I1142715,I1142732,I1142749,I1142766,I1142437,I1142458,I1142811,I1142449,I1142842,I1142859,I1142885,I1142893,I1142455,I1142924,I1142941,I1142958,I1142975,I1142446,I1142443,I1143047,I1143073,I1143081,I1143121,I1143129,I1143146,I1143163,I1143203,I1143225,I1143242,I1143268,I1143276,I1143293,I1143310,I1143327,I1143344,I1143389,I1143420,I1143437,I1143463,I1143471,I1143502,I1143519,I1143536,I1143553,I1143625,I1143651,I1143659,I1143699,I1143707,I1143724,I1143741,I1143781,I1143803,I1143820,I1143846,I1143854,I1143871,I1143888,I1143905,I1143922,I1143967,I1143998,I1144015,I1144041,I1144049,I1144080,I1144097,I1144114,I1144131,I1144203,I1144229,I1144237,I1144277,I1144285,I1144302,I1144319,I1144359,I1144381,I1144398,I1144424,I1144432,I1144449,I1144466,I1144483,I1144500,I1144545,I1144576,I1144593,I1144619,I1144627,I1144658,I1144675,I1144692,I1144709,I1144781,I1144807,I1144815,I1144855,I1144863,I1144880,I1144897,I1144937,I1144959,I1144976,I1145002,I1145010,I1145027,I1145044,I1145061,I1145078,I1145123,I1145154,I1145171,I1145197,I1145205,I1145236,I1145253,I1145270,I1145287,I1145359,I1145385,I1145393,I1145433,I1145441,I1145458,I1145475,I1145515,I1145537,I1145554,I1145580,I1145588,I1145605,I1145622,I1145639,I1145656,I1145701,I1145732,I1145749,I1145775,I1145783,I1145814,I1145831,I1145848,I1145865,I1145937,I1369635,I1145963,I1145971,I1369617,I1369608,I1146011,I1146019,I1369623,I1146036,I1369611,I1146053,I1146093,I1146115,I1369620,I1146132,I1146158,I1146166,I1146183,I1369629,I1146200,I1146217,I1146234,I1146279,I1369632,I1146310,I1146327,I1369626,I1369614,I1146353,I1146361,I1146392,I1146409,I1146426,I1146443,I1146515,I1146541,I1146549,I1146589,I1146597,I1146614,I1146631,I1146671,I1146693,I1146710,I1146736,I1146744,I1146761,I1146778,I1146795,I1146812,I1146857,I1146888,I1146905,I1146931,I1146939,I1146970,I1146987,I1147004,I1147021,I1147093,I1147119,I1147127,I1147167,I1147175,I1147192,I1147209,I1147249,I1147271,I1147288,I1147314,I1147322,I1147339,I1147356,I1147373,I1147390,I1147435,I1147466,I1147483,I1147509,I1147517,I1147548,I1147565,I1147582,I1147599,I1147671,I1147697,I1147705,I1147745,I1147753,I1147770,I1147787,I1147827,I1147849,I1147866,I1147892,I1147900,I1147917,I1147934,I1147951,I1147968,I1148013,I1148044,I1148061,I1148087,I1148095,I1148126,I1148143,I1148160,I1148177,I1148249,I1148275,I1148283,I1148323,I1148331,I1148348,I1148365,I1148405,I1148427,I1148444,I1148470,I1148478,I1148495,I1148512,I1148529,I1148546,I1148591,I1148622,I1148639,I1148665,I1148673,I1148704,I1148721,I1148738,I1148755,I1148827,I1148853,I1148861,I1148901,I1148909,I1148926,I1148943,I1148983,I1149005,I1149022,I1149048,I1149056,I1149073,I1149090,I1149107,I1149124,I1149169,I1149200,I1149217,I1149243,I1149251,I1149282,I1149299,I1149316,I1149333,I1149405,I1381535,I1149431,I1149439,I1381517,I1381508,I1149479,I1149487,I1381523,I1149504,I1381511,I1149521,I1149561,I1149583,I1381520,I1149600,I1149626,I1149634,I1149651,I1381529,I1149668,I1149685,I1149702,I1149747,I1381532,I1149778,I1149795,I1381526,I1381514,I1149821,I1149829,I1149860,I1149877,I1149894,I1149911,I1149983,I1363090,I1150009,I1150017,I1363072,I1363063,I1150057,I1150065,I1363078,I1150082,I1363066,I1150099,I1150139,I1150161,I1363075,I1150178,I1150204,I1150212,I1150229,I1363084,I1150246,I1150263,I1150280,I1150325,I1363087,I1150356,I1150373,I1363081,I1363069,I1150399,I1150407,I1150438,I1150455,I1150472,I1150489,I1150561,I1150587,I1150595,I1150635,I1150643,I1150660,I1150677,I1150717,I1150739,I1150756,I1150782,I1150790,I1150807,I1150824,I1150841,I1150858,I1150903,I1150934,I1150951,I1150977,I1150985,I1151016,I1151033,I1151050,I1151067,I1151139,I1151165,I1151173,I1151122,I1151213,I1151221,I1151238,I1151255,I1151110,I1151295,I1151131,I1151317,I1151334,I1151360,I1151368,I1151385,I1151402,I1151419,I1151436,I1151107,I1151128,I1151481,I1151119,I1151512,I1151529,I1151555,I1151563,I1151125,I1151594,I1151611,I1151628,I1151645,I1151116,I1151113,I1151717,I1151743,I1151751,I1151791,I1151799,I1151816,I1151833,I1151873,I1151895,I1151912,I1151938,I1151946,I1151963,I1151980,I1151997,I1152014,I1152059,I1152090,I1152107,I1152133,I1152141,I1152172,I1152189,I1152206,I1152223,I1152295,I1266014,I1152321,I1152329,I1266008,I1265993,I1152369,I1152377,I1265999,I1152394,I1266011,I1152411,I1152451,I1152473,I1152490,I1152516,I1152524,I1152541,I1266017,I1152558,I1266005,I1152575,I1152592,I1152637,I1265996,I1152668,I1152685,I1266002,I1152711,I1152719,I1152750,I1152767,I1152784,I1152801,I1152873,I1152899,I1152907,I1152947,I1152955,I1152972,I1152989,I1153029,I1153051,I1153068,I1153094,I1153102,I1153119,I1153136,I1153153,I1153170,I1153215,I1153246,I1153263,I1153289,I1153297,I1153328,I1153345,I1153362,I1153379,I1153451,I1153477,I1153485,I1153525,I1153533,I1153550,I1153567,I1153607,I1153629,I1153646,I1153672,I1153680,I1153697,I1153714,I1153731,I1153748,I1153793,I1153824,I1153841,I1153867,I1153875,I1153906,I1153923,I1153940,I1153957,I1154029,I1154055,I1154063,I1154103,I1154111,I1154128,I1154145,I1154185,I1154207,I1154224,I1154250,I1154258,I1154275,I1154292,I1154309,I1154326,I1154371,I1154402,I1154419,I1154445,I1154453,I1154484,I1154501,I1154518,I1154535,I1154607,I1154633,I1154641,I1154590,I1154681,I1154689,I1154706,I1154723,I1154578,I1154763,I1154599,I1154785,I1154802,I1154828,I1154836,I1154853,I1154870,I1154887,I1154904,I1154575,I1154596,I1154949,I1154587,I1154980,I1154997,I1155023,I1155031,I1154593,I1155062,I1155079,I1155096,I1155113,I1154584,I1154581,I1155185,I1155211,I1155219,I1155168,I1155259,I1155267,I1155284,I1155301,I1155156,I1155341,I1155177,I1155363,I1155380,I1155406,I1155414,I1155431,I1155448,I1155465,I1155482,I1155153,I1155174,I1155527,I1155165,I1155558,I1155575,I1155601,I1155609,I1155171,I1155640,I1155657,I1155674,I1155691,I1155162,I1155159,I1155763,I1343455,I1155789,I1155797,I1343437,I1343428,I1155837,I1155845,I1343443,I1155862,I1343431,I1155879,I1155919,I1155941,I1343440,I1155958,I1155984,I1155992,I1156009,I1343449,I1156026,I1156043,I1156060,I1156105,I1343452,I1156136,I1156153,I1343446,I1343434,I1156179,I1156187,I1156218,I1156235,I1156252,I1156269,I1156341,I1156367,I1156375,I1156415,I1156423,I1156440,I1156457,I1156497,I1156519,I1156536,I1156562,I1156570,I1156587,I1156604,I1156621,I1156638,I1156683,I1156714,I1156731,I1156757,I1156765,I1156796,I1156813,I1156830,I1156847,I1156919,I1156945,I1156953,I1156902,I1156993,I1157001,I1157018,I1157035,I1156890,I1157075,I1156911,I1157097,I1157114,I1157140,I1157148,I1157165,I1157182,I1157199,I1157216,I1156887,I1156908,I1157261,I1156899,I1157292,I1157309,I1157335,I1157343,I1156905,I1157374,I1157391,I1157408,I1157425,I1156896,I1156893,I1157497,I1157523,I1157531,I1157571,I1157579,I1157596,I1157613,I1157653,I1157675,I1157692,I1157718,I1157726,I1157743,I1157760,I1157777,I1157794,I1157839,I1157870,I1157887,I1157913,I1157921,I1157952,I1157969,I1157986,I1158003,I1158075,I1158101,I1158109,I1158149,I1158157,I1158174,I1158191,I1158231,I1158253,I1158270,I1158296,I1158304,I1158321,I1158338,I1158355,I1158372,I1158417,I1158448,I1158465,I1158491,I1158499,I1158530,I1158547,I1158564,I1158581,I1158653,I1158679,I1158687,I1158727,I1158735,I1158752,I1158769,I1158809,I1158831,I1158848,I1158874,I1158882,I1158899,I1158916,I1158933,I1158950,I1158995,I1159026,I1159043,I1159069,I1159077,I1159108,I1159125,I1159142,I1159159,I1159231,I1159257,I1159265,I1159305,I1159313,I1159330,I1159347,I1159387,I1159409,I1159426,I1159452,I1159460,I1159477,I1159494,I1159511,I1159528,I1159573,I1159604,I1159621,I1159647,I1159655,I1159686,I1159703,I1159720,I1159737,I1159809,I1159835,I1159843,I1159883,I1159891,I1159908,I1159925,I1159965,I1159987,I1160004,I1160030,I1160038,I1160055,I1160072,I1160089,I1160106,I1160151,I1160182,I1160199,I1160225,I1160233,I1160264,I1160281,I1160298,I1160315,I1160387,I1160413,I1160421,I1160461,I1160469,I1160486,I1160503,I1160543,I1160565,I1160582,I1160608,I1160616,I1160633,I1160650,I1160667,I1160684,I1160729,I1160760,I1160777,I1160803,I1160811,I1160842,I1160859,I1160876,I1160893,I1160965,I1276894,I1160991,I1160999,I1276888,I1160948,I1276873,I1161039,I1161047,I1276879,I1161064,I1276891,I1161081,I1160936,I1161121,I1160957,I1161143,I1161160,I1161186,I1161194,I1161211,I1276897,I1161228,I1276885,I1161245,I1161262,I1160933,I1160954,I1161307,I1276876,I1160945,I1161338,I1161355,I1276882,I1161381,I1161389,I1160951,I1161420,I1161437,I1161454,I1161471,I1160942,I1160939,I1161543,I1161569,I1161577,I1161617,I1161625,I1161642,I1161659,I1161699,I1161721,I1161738,I1161764,I1161772,I1161789,I1161806,I1161823,I1161840,I1161885,I1161916,I1161933,I1161959,I1161967,I1161998,I1162015,I1162032,I1162049,I1162121,I1162147,I1162155,I1162195,I1162203,I1162220,I1162237,I1162277,I1162299,I1162316,I1162342,I1162350,I1162367,I1162384,I1162401,I1162418,I1162463,I1162494,I1162511,I1162537,I1162545,I1162576,I1162593,I1162610,I1162627,I1162699,I1162725,I1162733,I1162773,I1162781,I1162798,I1162815,I1162855,I1162877,I1162894,I1162920,I1162928,I1162945,I1162962,I1162979,I1162996,I1163041,I1163072,I1163089,I1163115,I1163123,I1163154,I1163171,I1163188,I1163205,I1163277,I1163303,I1163311,I1163260,I1163351,I1163359,I1163376,I1163393,I1163248,I1163433,I1163269,I1163455,I1163472,I1163498,I1163506,I1163523,I1163540,I1163557,I1163574,I1163245,I1163266,I1163619,I1163257,I1163650,I1163667,I1163693,I1163701,I1163263,I1163732,I1163749,I1163766,I1163783,I1163254,I1163251,I1163855,I1388675,I1163881,I1163889,I1388657,I1388648,I1163929,I1163937,I1388663,I1163954,I1388651,I1163971,I1164011,I1164033,I1388660,I1164050,I1164076,I1164084,I1164101,I1388669,I1164118,I1164135,I1164152,I1164197,I1388672,I1164228,I1164245,I1388666,I1388654,I1164271,I1164279,I1164310,I1164327,I1164344,I1164361,I1164433,I1255678,I1164459,I1164467,I1255672,I1255657,I1164507,I1164515,I1255663,I1164532,I1255675,I1164549,I1164589,I1164611,I1164628,I1164654,I1164662,I1164679,I1255681,I1164696,I1255669,I1164713,I1164730,I1164775,I1255660,I1164806,I1164823,I1255666,I1164849,I1164857,I1164888,I1164905,I1164922,I1164939,I1165011,I1165037,I1165045,I1165085,I1165093,I1165110,I1165127,I1165167,I1165189,I1165206,I1165232,I1165240,I1165257,I1165274,I1165291,I1165308,I1165353,I1165384,I1165401,I1165427,I1165435,I1165466,I1165483,I1165500,I1165517,I1165589,I1165615,I1165623,I1165663,I1165671,I1165688,I1165705,I1165745,I1165767,I1165784,I1165810,I1165818,I1165835,I1165852,I1165869,I1165886,I1165931,I1165962,I1165979,I1166005,I1166013,I1166044,I1166061,I1166078,I1166095,I1166167,I1166193,I1166201,I1166241,I1166249,I1166266,I1166283,I1166323,I1166345,I1166362,I1166388,I1166396,I1166413,I1166430,I1166447,I1166464,I1166509,I1166540,I1166557,I1166583,I1166591,I1166622,I1166639,I1166656,I1166673,I1166745,I1166771,I1166779,I1166819,I1166827,I1166844,I1166861,I1166901,I1166923,I1166940,I1166966,I1166974,I1166991,I1167008,I1167025,I1167042,I1167087,I1167118,I1167135,I1167161,I1167169,I1167200,I1167217,I1167234,I1167251,I1167323,I1167349,I1167357,I1167397,I1167405,I1167422,I1167439,I1167479,I1167501,I1167518,I1167544,I1167552,I1167569,I1167586,I1167603,I1167620,I1167665,I1167696,I1167713,I1167739,I1167747,I1167778,I1167795,I1167812,I1167829,I1167901,I1167927,I1167935,I1167975,I1167983,I1168000,I1168017,I1168057,I1168079,I1168096,I1168122,I1168130,I1168147,I1168164,I1168181,I1168198,I1168243,I1168274,I1168291,I1168317,I1168325,I1168356,I1168373,I1168390,I1168407,I1168479,I1168505,I1168513,I1168553,I1168561,I1168578,I1168595,I1168635,I1168657,I1168674,I1168700,I1168708,I1168725,I1168742,I1168759,I1168776,I1168821,I1168852,I1168869,I1168895,I1168903,I1168934,I1168951,I1168968,I1168985,I1169057,I1169083,I1169091,I1169131,I1169139,I1169156,I1169173,I1169213,I1169235,I1169252,I1169278,I1169286,I1169303,I1169320,I1169337,I1169354,I1169399,I1169430,I1169447,I1169473,I1169481,I1169512,I1169529,I1169546,I1169563,I1169635,I1245886,I1169661,I1169669,I1245880,I1245865,I1169709,I1169717,I1245871,I1169734,I1245883,I1169751,I1169791,I1169813,I1169830,I1169856,I1169864,I1169881,I1245889,I1169898,I1245877,I1169915,I1169932,I1169977,I1245868,I1170008,I1170025,I1245874,I1170051,I1170059,I1170090,I1170107,I1170124,I1170141,I1170213,I1170239,I1170247,I1170287,I1170295,I1170312,I1170329,I1170369,I1170391,I1170408,I1170434,I1170442,I1170459,I1170476,I1170493,I1170510,I1170555,I1170586,I1170603,I1170629,I1170637,I1170668,I1170685,I1170702,I1170719,I1170791,I1170817,I1170825,I1170865,I1170873,I1170890,I1170907,I1170947,I1170969,I1170986,I1171012,I1171020,I1171037,I1171054,I1171071,I1171088,I1171133,I1171164,I1171181,I1171207,I1171215,I1171246,I1171263,I1171280,I1171297,I1171369,I1171395,I1171403,I1171443,I1171451,I1171468,I1171485,I1171525,I1171547,I1171564,I1171590,I1171598,I1171615,I1171632,I1171649,I1171666,I1171711,I1171742,I1171759,I1171785,I1171793,I1171824,I1171841,I1171858,I1171875,I1171947,I1171973,I1171981,I1172021,I1172029,I1172046,I1172063,I1172103,I1172125,I1172142,I1172168,I1172176,I1172193,I1172210,I1172227,I1172244,I1172289,I1172320,I1172337,I1172363,I1172371,I1172402,I1172419,I1172436,I1172453,I1172525,I1172551,I1172559,I1172599,I1172607,I1172624,I1172641,I1172681,I1172703,I1172720,I1172746,I1172754,I1172771,I1172788,I1172805,I1172822,I1172867,I1172898,I1172915,I1172941,I1172949,I1172980,I1172997,I1173014,I1173031,I1173103,I1173129,I1173137,I1173177,I1173185,I1173202,I1173219,I1173259,I1173281,I1173298,I1173324,I1173332,I1173349,I1173366,I1173383,I1173400,I1173445,I1173476,I1173493,I1173519,I1173527,I1173558,I1173575,I1173592,I1173609,I1173681,I1173707,I1173715,I1173755,I1173763,I1173780,I1173797,I1173837,I1173859,I1173876,I1173902,I1173910,I1173927,I1173944,I1173961,I1173978,I1174023,I1174054,I1174071,I1174097,I1174105,I1174136,I1174153,I1174170,I1174187,I1174259,I1174285,I1174293,I1174333,I1174341,I1174358,I1174375,I1174415,I1174437,I1174454,I1174480,I1174488,I1174505,I1174522,I1174539,I1174556,I1174601,I1174632,I1174649,I1174675,I1174683,I1174714,I1174731,I1174748,I1174765,I1174837,I1174863,I1174871,I1174911,I1174919,I1174936,I1174953,I1174993,I1175015,I1175032,I1175058,I1175066,I1175083,I1175100,I1175117,I1175134,I1175179,I1175210,I1175227,I1175253,I1175261,I1175292,I1175309,I1175326,I1175343,I1175415,I1175441,I1175449,I1175489,I1175497,I1175514,I1175531,I1175571,I1175593,I1175610,I1175636,I1175644,I1175661,I1175678,I1175695,I1175712,I1175757,I1175788,I1175805,I1175831,I1175839,I1175870,I1175887,I1175904,I1175921,I1175993,I1176019,I1176027,I1176067,I1176075,I1176092,I1176109,I1176149,I1176171,I1176188,I1176214,I1176222,I1176239,I1176256,I1176273,I1176290,I1176335,I1176366,I1176383,I1176409,I1176417,I1176448,I1176465,I1176482,I1176499,I1176571,I1176597,I1176605,I1176645,I1176653,I1176670,I1176687,I1176727,I1176749,I1176766,I1176792,I1176800,I1176817,I1176834,I1176851,I1176868,I1176913,I1176944,I1176961,I1176987,I1176995,I1177026,I1177043,I1177060,I1177077,I1177149,I1177175,I1177183,I1177223,I1177231,I1177248,I1177265,I1177305,I1177327,I1177344,I1177370,I1177378,I1177395,I1177412,I1177429,I1177446,I1177491,I1177522,I1177539,I1177565,I1177573,I1177604,I1177621,I1177638,I1177655,I1177727,I1177753,I1177761,I1177801,I1177809,I1177826,I1177843,I1177883,I1177905,I1177922,I1177948,I1177956,I1177973,I1177990,I1178007,I1178024,I1178069,I1178100,I1178117,I1178143,I1178151,I1178182,I1178199,I1178216,I1178233,I1178305,I1178331,I1178339,I1178379,I1178387,I1178404,I1178421,I1178461,I1178483,I1178500,I1178526,I1178534,I1178551,I1178568,I1178585,I1178602,I1178647,I1178678,I1178695,I1178721,I1178729,I1178760,I1178777,I1178794,I1178811,I1178883,I1178909,I1178917,I1178957,I1178965,I1178982,I1178999,I1179039,I1179061,I1179078,I1179104,I1179112,I1179129,I1179146,I1179163,I1179180,I1179225,I1179256,I1179273,I1179299,I1179307,I1179338,I1179355,I1179372,I1179389,I1179461,I1179487,I1179495,I1179535,I1179543,I1179560,I1179577,I1179617,I1179639,I1179656,I1179682,I1179690,I1179707,I1179724,I1179741,I1179758,I1179803,I1179834,I1179851,I1179877,I1179885,I1179916,I1179933,I1179950,I1179967,I1180039,I1376775,I1180065,I1180073,I1376757,I1376748,I1180113,I1180121,I1376763,I1180138,I1376751,I1180155,I1180195,I1180217,I1376760,I1180234,I1180260,I1180268,I1180285,I1376769,I1180302,I1180319,I1180336,I1180381,I1376772,I1180412,I1180429,I1376766,I1376754,I1180455,I1180463,I1180494,I1180511,I1180528,I1180545,I1180617,I1180643,I1180651,I1180691,I1180699,I1180716,I1180733,I1180773,I1180795,I1180812,I1180838,I1180846,I1180863,I1180880,I1180897,I1180914,I1180959,I1180990,I1181007,I1181033,I1181041,I1181072,I1181089,I1181106,I1181123,I1181195,I1318411,I1181221,I1181229,I1318393,I1318402,I1181269,I1181277,I1318387,I1181294,I1318399,I1181311,I1181351,I1181373,I1318390,I1181390,I1181416,I1181424,I1181441,I1181458,I1181475,I1181492,I1181537,I1318408,I1181568,I1181585,I1318396,I1318405,I1181611,I1181619,I1181650,I1181667,I1181684,I1181701,I1181773,I1181799,I1181807,I1181847,I1181855,I1181872,I1181889,I1181929,I1181951,I1181968,I1181994,I1182002,I1182019,I1182036,I1182053,I1182070,I1182115,I1182146,I1182163,I1182189,I1182197,I1182228,I1182245,I1182262,I1182279,I1182351,I1285054,I1182377,I1182385,I1285048,I1285033,I1182425,I1182433,I1285039,I1182450,I1285051,I1182467,I1182507,I1182529,I1182546,I1182572,I1182580,I1182597,I1285057,I1182614,I1285045,I1182631,I1182648,I1182693,I1285036,I1182724,I1182741,I1285042,I1182767,I1182775,I1182806,I1182823,I1182840,I1182857,I1182929,I1182955,I1182963,I1183003,I1183011,I1183028,I1183045,I1183085,I1183107,I1183124,I1183150,I1183158,I1183175,I1183192,I1183209,I1183226,I1183271,I1183302,I1183319,I1183345,I1183353,I1183384,I1183401,I1183418,I1183435,I1183507,I1183533,I1183541,I1183581,I1183589,I1183606,I1183623,I1183663,I1183685,I1183702,I1183728,I1183736,I1183753,I1183770,I1183787,I1183804,I1183849,I1183880,I1183897,I1183923,I1183931,I1183962,I1183979,I1183996,I1184013,I1184085,I1184111,I1184119,I1184159,I1184167,I1184184,I1184201,I1184241,I1184263,I1184280,I1184306,I1184314,I1184331,I1184348,I1184365,I1184382,I1184427,I1184458,I1184475,I1184501,I1184509,I1184540,I1184557,I1184574,I1184591,I1184663,I1184689,I1184697,I1184646,I1184737,I1184745,I1184762,I1184779,I1184634,I1184819,I1184655,I1184841,I1184858,I1184884,I1184892,I1184909,I1184926,I1184943,I1184960,I1184631,I1184652,I1185005,I1184643,I1185036,I1185053,I1185079,I1185087,I1184649,I1185118,I1185135,I1185152,I1185169,I1184640,I1184637,I1185241,I1185267,I1185275,I1185315,I1185323,I1185340,I1185357,I1185397,I1185419,I1185436,I1185462,I1185470,I1185487,I1185504,I1185521,I1185538,I1185583,I1185614,I1185631,I1185657,I1185665,I1185696,I1185713,I1185730,I1185747,I1185819,I1402360,I1185845,I1185853,I1402342,I1402333,I1185893,I1185901,I1402348,I1185918,I1402336,I1185935,I1185975,I1185997,I1402345,I1186014,I1186040,I1186048,I1186065,I1402354,I1186082,I1186099,I1186116,I1186161,I1402357,I1186192,I1186209,I1402351,I1402339,I1186235,I1186243,I1186274,I1186291,I1186308,I1186325,I1186397,I1186423,I1186431,I1186471,I1186479,I1186496,I1186513,I1186553,I1186575,I1186592,I1186618,I1186626,I1186643,I1186660,I1186677,I1186694,I1186739,I1186770,I1186787,I1186813,I1186821,I1186852,I1186869,I1186886,I1186903,I1186975,I1187001,I1187009,I1186958,I1187049,I1187057,I1187074,I1187091,I1186946,I1187131,I1186967,I1187153,I1187170,I1187196,I1187204,I1187221,I1187238,I1187255,I1187272,I1186943,I1186964,I1187317,I1186955,I1187348,I1187365,I1187391,I1187399,I1186961,I1187430,I1187447,I1187464,I1187481,I1186952,I1186949,I1187553,I1187579,I1187587,I1187536,I1187627,I1187635,I1187652,I1187669,I1187524,I1187709,I1187545,I1187731,I1187748,I1187774,I1187782,I1187799,I1187816,I1187833,I1187850,I1187521,I1187542,I1187895,I1187533,I1187926,I1187943,I1187969,I1187977,I1187539,I1188008,I1188025,I1188042,I1188059,I1187530,I1187527,I1188131,I1188157,I1188165,I1188205,I1188213,I1188230,I1188247,I1188287,I1188309,I1188326,I1188352,I1188360,I1188377,I1188394,I1188411,I1188428,I1188473,I1188504,I1188521,I1188547,I1188555,I1188586,I1188603,I1188620,I1188637,I1188709,I1188735,I1188743,I1188692,I1188783,I1188791,I1188808,I1188825,I1188680,I1188865,I1188701,I1188887,I1188904,I1188930,I1188938,I1188955,I1188972,I1188989,I1189006,I1188677,I1188698,I1189051,I1188689,I1189082,I1189099,I1189125,I1189133,I1188695,I1189164,I1189181,I1189198,I1189215,I1188686,I1188683,I1189287,I1189313,I1189321,I1189361,I1189369,I1189386,I1189403,I1189443,I1189465,I1189482,I1189508,I1189516,I1189533,I1189550,I1189567,I1189584,I1189629,I1189660,I1189677,I1189703,I1189711,I1189742,I1189759,I1189776,I1189793,I1189865,I1367850,I1189891,I1189899,I1367832,I1367823,I1189939,I1189947,I1367838,I1189964,I1367826,I1189981,I1190021,I1190043,I1367835,I1190060,I1190086,I1190094,I1190111,I1367844,I1190128,I1190145,I1190162,I1190207,I1367847,I1190238,I1190255,I1367841,I1367829,I1190281,I1190289,I1190320,I1190337,I1190354,I1190371,I1190443,I1190469,I1190477,I1190517,I1190525,I1190542,I1190559,I1190599,I1190621,I1190638,I1190664,I1190672,I1190689,I1190706,I1190723,I1190740,I1190785,I1190816,I1190833,I1190859,I1190867,I1190898,I1190915,I1190932,I1190949,I1191021,I1191047,I1191055,I1191095,I1191103,I1191120,I1191137,I1191177,I1191199,I1191216,I1191242,I1191250,I1191267,I1191284,I1191301,I1191318,I1191363,I1191394,I1191411,I1191437,I1191445,I1191476,I1191493,I1191510,I1191527,I1191599,I1191625,I1191633,I1191673,I1191681,I1191698,I1191715,I1191755,I1191777,I1191794,I1191820,I1191828,I1191845,I1191862,I1191879,I1191896,I1191941,I1191972,I1191989,I1192015,I1192023,I1192054,I1192071,I1192088,I1192105,I1192177,I1192203,I1192211,I1192251,I1192259,I1192276,I1192293,I1192333,I1192355,I1192372,I1192398,I1192406,I1192423,I1192440,I1192457,I1192474,I1192519,I1192550,I1192567,I1192593,I1192601,I1192632,I1192649,I1192666,I1192683,I1192755,I1192781,I1192789,I1192829,I1192837,I1192854,I1192871,I1192911,I1192933,I1192950,I1192976,I1192984,I1193001,I1193018,I1193035,I1193052,I1193097,I1193128,I1193145,I1193171,I1193179,I1193210,I1193227,I1193244,I1193261,I1193333,I1193359,I1193367,I1193316,I1193407,I1193415,I1193432,I1193449,I1193304,I1193489,I1193325,I1193511,I1193528,I1193554,I1193562,I1193579,I1193596,I1193613,I1193630,I1193301,I1193322,I1193675,I1193313,I1193706,I1193723,I1193749,I1193757,I1193319,I1193788,I1193805,I1193822,I1193839,I1193310,I1193307,I1193911,I1383320,I1193937,I1193945,I1383302,I1383293,I1193985,I1193993,I1383308,I1194010,I1383296,I1194027,I1194067,I1194089,I1383305,I1194106,I1194132,I1194140,I1194157,I1383314,I1194174,I1194191,I1194208,I1194253,I1383317,I1194284,I1194301,I1383311,I1383299,I1194327,I1194335,I1194366,I1194383,I1194400,I1194417,I1194489,I1194515,I1194523,I1194563,I1194571,I1194588,I1194605,I1194645,I1194667,I1194684,I1194710,I1194718,I1194735,I1194752,I1194769,I1194786,I1194831,I1194862,I1194879,I1194905,I1194913,I1194944,I1194961,I1194978,I1194995,I1195067,I1195093,I1195101,I1195141,I1195149,I1195166,I1195183,I1195223,I1195245,I1195262,I1195288,I1195296,I1195313,I1195330,I1195347,I1195364,I1195409,I1195440,I1195457,I1195483,I1195491,I1195522,I1195539,I1195556,I1195573,I1195645,I1195671,I1195679,I1195628,I1195719,I1195727,I1195744,I1195761,I1195616,I1195801,I1195637,I1195823,I1195840,I1195866,I1195874,I1195891,I1195908,I1195925,I1195942,I1195613,I1195634,I1195987,I1195625,I1196018,I1196035,I1196061,I1196069,I1195631,I1196100,I1196117,I1196134,I1196151,I1195622,I1195619,I1196223,I1196249,I1196257,I1196206,I1196297,I1196305,I1196322,I1196339,I1196194,I1196379,I1196215,I1196401,I1196418,I1196444,I1196452,I1196469,I1196486,I1196503,I1196520,I1196191,I1196212,I1196565,I1196203,I1196596,I1196613,I1196639,I1196647,I1196209,I1196678,I1196695,I1196712,I1196729,I1196200,I1196197,I1196801,I1196827,I1196835,I1196875,I1196883,I1196900,I1196917,I1196957,I1196979,I1196996,I1197022,I1197030,I1197047,I1197064,I1197081,I1197098,I1197143,I1197174,I1197191,I1197217,I1197225,I1197256,I1197273,I1197290,I1197307,I1197379,I1197405,I1197413,I1197362,I1197453,I1197461,I1197478,I1197495,I1197350,I1197535,I1197371,I1197557,I1197574,I1197600,I1197608,I1197625,I1197642,I1197659,I1197676,I1197347,I1197368,I1197721,I1197359,I1197752,I1197769,I1197795,I1197803,I1197365,I1197834,I1197851,I1197868,I1197885,I1197356,I1197353,I1197957,I1197983,I1197991,I1198031,I1198039,I1198056,I1198073,I1198113,I1198135,I1198152,I1198178,I1198186,I1198203,I1198220,I1198237,I1198254,I1198299,I1198330,I1198347,I1198373,I1198381,I1198412,I1198429,I1198446,I1198463,I1198535,I1198561,I1198569,I1198609,I1198617,I1198634,I1198651,I1198691,I1198713,I1198730,I1198756,I1198764,I1198781,I1198798,I1198815,I1198832,I1198877,I1198908,I1198925,I1198951,I1198959,I1198990,I1199007,I1199024,I1199041,I1199113,I1199139,I1199147,I1199187,I1199195,I1199212,I1199229,I1199269,I1199291,I1199308,I1199334,I1199342,I1199359,I1199376,I1199393,I1199410,I1199455,I1199486,I1199503,I1199529,I1199537,I1199568,I1199585,I1199602,I1199619,I1199691,I1199717,I1199725,I1199765,I1199773,I1199790,I1199807,I1199847,I1199869,I1199886,I1199912,I1199920,I1199937,I1199954,I1199971,I1199988,I1200033,I1200064,I1200081,I1200107,I1200115,I1200146,I1200163,I1200180,I1200197,I1200269,I1200295,I1200303,I1200343,I1200351,I1200368,I1200385,I1200425,I1200447,I1200464,I1200490,I1200498,I1200515,I1200532,I1200549,I1200566,I1200611,I1200642,I1200659,I1200685,I1200693,I1200724,I1200741,I1200758,I1200775,I1200847,I1336910,I1200873,I1200881,I1336892,I1336883,I1200921,I1200929,I1336898,I1200946,I1336886,I1200963,I1201003,I1201025,I1336895,I1201042,I1201068,I1201076,I1201093,I1336904,I1201110,I1201127,I1201144,I1201189,I1336907,I1201220,I1201237,I1336901,I1336889,I1201263,I1201271,I1201302,I1201319,I1201336,I1201353,I1201425,I1201451,I1201459,I1201499,I1201507,I1201524,I1201541,I1201581,I1201603,I1201620,I1201646,I1201654,I1201671,I1201688,I1201705,I1201722,I1201767,I1201798,I1201815,I1201841,I1201849,I1201880,I1201897,I1201914,I1201931,I1202003,I1202029,I1202037,I1202077,I1202085,I1202102,I1202119,I1202159,I1202181,I1202198,I1202224,I1202232,I1202249,I1202266,I1202283,I1202300,I1202345,I1202376,I1202393,I1202419,I1202427,I1202458,I1202475,I1202492,I1202509,I1202581,I1202607,I1202615,I1202655,I1202663,I1202680,I1202697,I1202737,I1202759,I1202776,I1202802,I1202810,I1202827,I1202844,I1202861,I1202878,I1202923,I1202954,I1202971,I1202997,I1203005,I1203036,I1203053,I1203070,I1203087,I1203159,I1203185,I1203193,I1203233,I1203241,I1203258,I1203275,I1203315,I1203337,I1203354,I1203380,I1203388,I1203405,I1203422,I1203439,I1203456,I1203501,I1203532,I1203549,I1203575,I1203583,I1203614,I1203631,I1203648,I1203665,I1203737,I1203763,I1203771,I1203811,I1203819,I1203836,I1203853,I1203893,I1203915,I1203932,I1203958,I1203966,I1203983,I1204000,I1204017,I1204034,I1204079,I1204110,I1204127,I1204153,I1204161,I1204192,I1204209,I1204226,I1204243,I1204315,I1204341,I1204349,I1204389,I1204397,I1204414,I1204431,I1204471,I1204493,I1204510,I1204536,I1204544,I1204561,I1204578,I1204595,I1204612,I1204657,I1204688,I1204705,I1204731,I1204739,I1204770,I1204787,I1204804,I1204821,I1204893,I1204919,I1204927,I1204967,I1204975,I1204992,I1205009,I1205049,I1205071,I1205088,I1205114,I1205122,I1205139,I1205156,I1205173,I1205190,I1205235,I1205266,I1205283,I1205309,I1205317,I1205348,I1205365,I1205382,I1205399,I1205471,I1361900,I1205497,I1205505,I1361882,I1361873,I1205545,I1205553,I1361888,I1205570,I1361876,I1205587,I1205627,I1205649,I1361885,I1205666,I1205692,I1205700,I1205717,I1361894,I1205734,I1205751,I1205768,I1205813,I1361897,I1205844,I1205861,I1361891,I1361879,I1205887,I1205895,I1205926,I1205943,I1205960,I1205977,I1206049,I1206075,I1206083,I1206032,I1206123,I1206131,I1206148,I1206165,I1206020,I1206205,I1206041,I1206227,I1206244,I1206270,I1206278,I1206295,I1206312,I1206329,I1206346,I1206017,I1206038,I1206391,I1206029,I1206422,I1206439,I1206465,I1206473,I1206035,I1206504,I1206521,I1206538,I1206555,I1206026,I1206023,I1206627,I1206653,I1206661,I1206701,I1206709,I1206726,I1206743,I1206783,I1206805,I1206822,I1206848,I1206856,I1206873,I1206890,I1206907,I1206924,I1206969,I1207000,I1207017,I1207043,I1207051,I1207082,I1207099,I1207116,I1207133,I1207205,I1207231,I1207239,I1207279,I1207287,I1207304,I1207321,I1207361,I1207383,I1207400,I1207426,I1207434,I1207451,I1207468,I1207485,I1207502,I1207547,I1207578,I1207595,I1207621,I1207629,I1207660,I1207677,I1207694,I1207711,I1207783,I1207809,I1207817,I1207857,I1207865,I1207882,I1207899,I1207939,I1207961,I1207978,I1208004,I1208012,I1208029,I1208046,I1208063,I1208080,I1208125,I1208156,I1208173,I1208199,I1208207,I1208238,I1208255,I1208272,I1208289,I1208361,I1208387,I1208395,I1208435,I1208443,I1208460,I1208477,I1208517,I1208539,I1208556,I1208582,I1208590,I1208607,I1208624,I1208641,I1208658,I1208703,I1208734,I1208751,I1208777,I1208785,I1208816,I1208833,I1208850,I1208867,I1208939,I1208965,I1208973,I1208922,I1209013,I1209021,I1209038,I1209055,I1208910,I1209095,I1208931,I1209117,I1209134,I1209160,I1209168,I1209185,I1209202,I1209219,I1209236,I1208907,I1208928,I1209281,I1208919,I1209312,I1209329,I1209355,I1209363,I1208925,I1209394,I1209411,I1209428,I1209445,I1208916,I1208913,I1209517,I1209543,I1209551,I1209591,I1209599,I1209616,I1209633,I1209673,I1209695,I1209712,I1209738,I1209746,I1209763,I1209780,I1209797,I1209814,I1209859,I1209890,I1209907,I1209933,I1209941,I1209972,I1209989,I1210006,I1210023,I1210095,I1340480,I1210121,I1210129,I1340462,I1210078,I1340453,I1210169,I1210177,I1340468,I1210194,I1340456,I1210211,I1210066,I1210251,I1210087,I1210273,I1340465,I1210290,I1210316,I1210324,I1210341,I1340474,I1210358,I1210375,I1210392,I1210063,I1210084,I1210437,I1340477,I1210075,I1210468,I1210485,I1340471,I1340459,I1210511,I1210519,I1210081,I1210550,I1210567,I1210584,I1210601,I1210072,I1210069,I1210673,I1210699,I1210707,I1210747,I1210755,I1210772,I1210789,I1210829,I1210851,I1210868,I1210894,I1210902,I1210919,I1210936,I1210953,I1210970,I1211015,I1211046,I1211063,I1211089,I1211097,I1211128,I1211145,I1211162,I1211179,I1211251,I1211277,I1211285,I1211325,I1211333,I1211350,I1211367,I1211407,I1211429,I1211446,I1211472,I1211480,I1211497,I1211514,I1211531,I1211548,I1211593,I1211624,I1211641,I1211667,I1211675,I1211706,I1211723,I1211740,I1211757,I1211829,I1359520,I1211855,I1211863,I1359502,I1359493,I1211903,I1211911,I1359508,I1211928,I1359496,I1211945,I1211985,I1212007,I1359505,I1212024,I1212050,I1212058,I1212075,I1359514,I1212092,I1212109,I1212126,I1212171,I1359517,I1212202,I1212219,I1359511,I1359499,I1212245,I1212253,I1212284,I1212301,I1212318,I1212335,I1212407,I1212433,I1212441,I1212481,I1212489,I1212506,I1212523,I1212563,I1212585,I1212602,I1212628,I1212636,I1212653,I1212670,I1212687,I1212704,I1212749,I1212780,I1212797,I1212823,I1212831,I1212862,I1212879,I1212896,I1212913,I1212985,I1213011,I1213019,I1213059,I1213067,I1213084,I1213101,I1213141,I1213163,I1213180,I1213206,I1213214,I1213231,I1213248,I1213265,I1213282,I1213327,I1213358,I1213375,I1213401,I1213409,I1213440,I1213457,I1213474,I1213491,I1213563,I1213589,I1213597,I1213637,I1213645,I1213662,I1213679,I1213719,I1213741,I1213758,I1213784,I1213792,I1213809,I1213826,I1213843,I1213860,I1213905,I1213936,I1213953,I1213979,I1213987,I1214018,I1214035,I1214052,I1214069,I1214141,I1214167,I1214175,I1214215,I1214223,I1214240,I1214257,I1214297,I1214319,I1214336,I1214362,I1214370,I1214387,I1214404,I1214421,I1214438,I1214483,I1214514,I1214531,I1214557,I1214565,I1214596,I1214613,I1214630,I1214647,I1214719,I1214745,I1214753,I1214702,I1214793,I1214801,I1214818,I1214835,I1214690,I1214875,I1214711,I1214897,I1214914,I1214940,I1214948,I1214965,I1214982,I1214999,I1215016,I1214687,I1214708,I1215061,I1214699,I1215092,I1215109,I1215135,I1215143,I1214705,I1215174,I1215191,I1215208,I1215225,I1214696,I1214693,I1215297,I1246430,I1215323,I1215331,I1246424,I1246409,I1215371,I1215379,I1246415,I1215396,I1246427,I1215413,I1215453,I1215475,I1215492,I1215518,I1215526,I1215543,I1246433,I1215560,I1246421,I1215577,I1215594,I1215639,I1246412,I1215670,I1215687,I1246418,I1215713,I1215721,I1215752,I1215769,I1215786,I1215803,I1215875,I1337505,I1215901,I1215909,I1337487,I1215858,I1337478,I1215949,I1215957,I1337493,I1215974,I1337481,I1215991,I1215846,I1216031,I1215867,I1216053,I1337490,I1216070,I1216096,I1216104,I1216121,I1337499,I1216138,I1216155,I1216172,I1215843,I1215864,I1216217,I1337502,I1215855,I1216248,I1216265,I1337496,I1337484,I1216291,I1216299,I1215861,I1216330,I1216347,I1216364,I1216381,I1215852,I1215849,I1216453,I1356545,I1216479,I1216487,I1356527,I1356518,I1216527,I1216535,I1356533,I1216552,I1356521,I1216569,I1216609,I1216631,I1356530,I1216648,I1216674,I1216682,I1216699,I1356539,I1216716,I1216733,I1216750,I1216795,I1356542,I1216826,I1216843,I1356536,I1356524,I1216869,I1216877,I1216908,I1216925,I1216942,I1216959,I1217031,I1217057,I1217065,I1217105,I1217113,I1217130,I1217147,I1217187,I1217209,I1217226,I1217252,I1217260,I1217277,I1217294,I1217311,I1217328,I1217373,I1217404,I1217421,I1217447,I1217455,I1217486,I1217503,I1217520,I1217537,I1217609,I1217635,I1217643,I1217683,I1217691,I1217708,I1217725,I1217765,I1217787,I1217804,I1217830,I1217838,I1217855,I1217872,I1217889,I1217906,I1217951,I1217982,I1217999,I1218025,I1218033,I1218064,I1218081,I1218098,I1218115,I1218187,I1218213,I1218221,I1218261,I1218269,I1218286,I1218303,I1218343,I1218365,I1218382,I1218408,I1218416,I1218433,I1218450,I1218467,I1218484,I1218529,I1218560,I1218577,I1218603,I1218611,I1218642,I1218659,I1218676,I1218693,I1218765,I1218791,I1218799,I1218839,I1218847,I1218864,I1218881,I1218921,I1218943,I1218960,I1218986,I1218994,I1219011,I1219028,I1219045,I1219062,I1219107,I1219138,I1219155,I1219181,I1219189,I1219220,I1219237,I1219254,I1219271,I1219343,I1219369,I1219377,I1219417,I1219425,I1219442,I1219459,I1219499,I1219521,I1219538,I1219564,I1219572,I1219589,I1219606,I1219623,I1219640,I1219685,I1219716,I1219733,I1219759,I1219767,I1219798,I1219815,I1219832,I1219849,I1219921,I1219947,I1219955,I1219995,I1220003,I1220020,I1220037,I1220077,I1220099,I1220116,I1220142,I1220150,I1220167,I1220184,I1220201,I1220218,I1220263,I1220294,I1220311,I1220337,I1220345,I1220376,I1220393,I1220410,I1220427,I1220499,I1366065,I1220525,I1220533,I1366047,I1220482,I1366038,I1220573,I1220581,I1366053,I1220598,I1366041,I1220615,I1220470,I1220655,I1220491,I1220677,I1366050,I1220694,I1220720,I1220728,I1220745,I1366059,I1220762,I1220779,I1220796,I1220467,I1220488,I1220841,I1366062,I1220479,I1220872,I1220889,I1366056,I1366044,I1220915,I1220923,I1220485,I1220954,I1220971,I1220988,I1221005,I1220476,I1220473,I1221077,I1221103,I1221111,I1221151,I1221159,I1221176,I1221193,I1221233,I1221255,I1221272,I1221298,I1221306,I1221323,I1221340,I1221357,I1221374,I1221419,I1221450,I1221467,I1221493,I1221501,I1221532,I1221549,I1221566,I1221583,I1221655,I1303961,I1221681,I1221689,I1303943,I1303952,I1221729,I1221737,I1303937,I1221754,I1303949,I1221771,I1221811,I1221833,I1303940,I1221850,I1221876,I1221884,I1221901,I1221918,I1221935,I1221952,I1221997,I1303958,I1222028,I1222045,I1303946,I1303955,I1222071,I1222079,I1222110,I1222127,I1222144,I1222161,I1222233,I1222259,I1222267,I1222216,I1222307,I1222315,I1222332,I1222349,I1222204,I1222389,I1222225,I1222411,I1222428,I1222454,I1222462,I1222479,I1222496,I1222513,I1222530,I1222201,I1222222,I1222575,I1222213,I1222606,I1222623,I1222649,I1222657,I1222219,I1222688,I1222705,I1222722,I1222739,I1222210,I1222207,I1222811,I1222837,I1222845,I1222885,I1222893,I1222910,I1222927,I1222967,I1222989,I1223006,I1223032,I1223040,I1223057,I1223074,I1223091,I1223108,I1223153,I1223184,I1223201,I1223227,I1223235,I1223266,I1223283,I1223300,I1223317,I1223389,I1223415,I1223423,I1223463,I1223471,I1223488,I1223505,I1223545,I1223567,I1223584,I1223610,I1223618,I1223635,I1223652,I1223669,I1223686,I1223731,I1223762,I1223779,I1223805,I1223813,I1223844,I1223861,I1223878,I1223895,I1223967,I1223993,I1224001,I1224041,I1224049,I1224066,I1224083,I1224123,I1224145,I1224162,I1224188,I1224196,I1224213,I1224230,I1224247,I1224264,I1224309,I1224340,I1224357,I1224383,I1224391,I1224422,I1224439,I1224456,I1224473,I1224545,I1224571,I1224579,I1224528,I1224619,I1224627,I1224644,I1224661,I1224516,I1224701,I1224537,I1224723,I1224740,I1224766,I1224774,I1224791,I1224808,I1224825,I1224842,I1224513,I1224534,I1224887,I1224525,I1224918,I1224935,I1224961,I1224969,I1224531,I1225000,I1225017,I1225034,I1225051,I1224522,I1224519,I1225123,I1367255,I1225149,I1225157,I1367237,I1367228,I1225197,I1225205,I1367243,I1225222,I1367231,I1225239,I1225279,I1225301,I1367240,I1225318,I1225344,I1225352,I1225369,I1367249,I1225386,I1225403,I1225420,I1225465,I1367252,I1225496,I1225513,I1367246,I1367234,I1225539,I1225547,I1225578,I1225595,I1225612,I1225629,I1225701,I1225727,I1225735,I1225684,I1225775,I1225783,I1225800,I1225817,I1225672,I1225857,I1225693,I1225879,I1225896,I1225922,I1225930,I1225947,I1225964,I1225981,I1225998,I1225669,I1225690,I1226043,I1225681,I1226074,I1226091,I1226117,I1226125,I1225687,I1226156,I1226173,I1226190,I1226207,I1225678,I1225675,I1226279,I1246974,I1226305,I1226313,I1246968,I1246953,I1226353,I1226361,I1246959,I1226378,I1246971,I1226395,I1226435,I1226457,I1226474,I1226500,I1226508,I1226525,I1246977,I1226542,I1246965,I1226559,I1226576,I1226621,I1246956,I1226652,I1226669,I1246962,I1226695,I1226703,I1226734,I1226751,I1226768,I1226785,I1226857,I1226883,I1226891,I1226931,I1226939,I1226956,I1226973,I1227013,I1227035,I1227052,I1227078,I1227086,I1227103,I1227120,I1227137,I1227154,I1227199,I1227230,I1227247,I1227273,I1227281,I1227312,I1227329,I1227346,I1227363,I1227435,I1227461,I1227469,I1227418,I1227509,I1227517,I1227534,I1227551,I1227406,I1227591,I1227427,I1227613,I1227630,I1227656,I1227664,I1227681,I1227698,I1227715,I1227732,I1227403,I1227424,I1227777,I1227415,I1227808,I1227825,I1227851,I1227859,I1227421,I1227890,I1227907,I1227924,I1227941,I1227412,I1227409,I1228013,I1228039,I1228047,I1228087,I1228095,I1228112,I1228129,I1228169,I1228191,I1228208,I1228234,I1228242,I1228259,I1228276,I1228293,I1228310,I1228355,I1228386,I1228403,I1228429,I1228437,I1228468,I1228485,I1228502,I1228519,I1228591,I1256222,I1228617,I1228625,I1256216,I1256201,I1228665,I1228673,I1256207,I1228690,I1256219,I1228707,I1228747,I1228769,I1228786,I1228812,I1228820,I1228837,I1256225,I1228854,I1256213,I1228871,I1228888,I1228933,I1256204,I1228964,I1228981,I1256210,I1229007,I1229015,I1229046,I1229063,I1229080,I1229097,I1229169,I1229195,I1229203,I1229243,I1229251,I1229268,I1229285,I1229325,I1229347,I1229364,I1229390,I1229398,I1229415,I1229432,I1229449,I1229466,I1229511,I1229542,I1229559,I1229585,I1229593,I1229624,I1229641,I1229658,I1229675,I1229747,I1229773,I1229781,I1229821,I1229829,I1229846,I1229863,I1229903,I1229925,I1229942,I1229968,I1229976,I1229993,I1230010,I1230027,I1230044,I1230089,I1230120,I1230137,I1230163,I1230171,I1230202,I1230219,I1230236,I1230253,I1230325,I1287230,I1230351,I1230359,I1287224,I1287209,I1230399,I1230407,I1287215,I1230424,I1287227,I1230441,I1230481,I1230503,I1230520,I1230546,I1230554,I1230571,I1287233,I1230588,I1287221,I1230605,I1230622,I1230667,I1287212,I1230698,I1230715,I1287218,I1230741,I1230749,I1230780,I1230797,I1230814,I1230831,I1230903,I1230929,I1230937,I1230977,I1230985,I1231002,I1231019,I1231059,I1231081,I1231098,I1231124,I1231132,I1231149,I1231166,I1231183,I1231200,I1231245,I1231276,I1231293,I1231319,I1231327,I1231358,I1231375,I1231392,I1231409,I1231481,I1231507,I1231515,I1231464,I1231555,I1231563,I1231580,I1231597,I1231452,I1231637,I1231473,I1231659,I1231676,I1231702,I1231710,I1231727,I1231744,I1231761,I1231778,I1231449,I1231470,I1231823,I1231461,I1231854,I1231871,I1231897,I1231905,I1231467,I1231936,I1231953,I1231970,I1231987,I1231458,I1231455,I1232059,I1232085,I1232093,I1232133,I1232141,I1232158,I1232175,I1232215,I1232237,I1232254,I1232280,I1232288,I1232305,I1232322,I1232339,I1232356,I1232401,I1232432,I1232449,I1232475,I1232483,I1232514,I1232531,I1232548,I1232565,I1232637,I1232663,I1232671,I1232711,I1232719,I1232736,I1232753,I1232793,I1232815,I1232832,I1232858,I1232866,I1232883,I1232900,I1232917,I1232934,I1232979,I1233010,I1233027,I1233053,I1233061,I1233092,I1233109,I1233126,I1233143,I1233215,I1233241,I1233249,I1233289,I1233297,I1233314,I1233331,I1233371,I1233393,I1233410,I1233436,I1233444,I1233461,I1233478,I1233495,I1233512,I1233557,I1233588,I1233605,I1233631,I1233639,I1233670,I1233687,I1233704,I1233721,I1233793,I1233819,I1233827,I1233867,I1233875,I1233892,I1233909,I1233949,I1233971,I1233988,I1234014,I1234022,I1234039,I1234056,I1234073,I1234090,I1234135,I1234166,I1234183,I1234209,I1234217,I1234248,I1234265,I1234282,I1234299,I1234371,I1234397,I1234405,I1234445,I1234453,I1234470,I1234487,I1234527,I1234549,I1234566,I1234592,I1234600,I1234617,I1234634,I1234651,I1234668,I1234713,I1234744,I1234761,I1234787,I1234795,I1234826,I1234843,I1234860,I1234877,I1234949,I1234975,I1234983,I1235023,I1235031,I1235048,I1235065,I1235105,I1235127,I1235144,I1235170,I1235178,I1235195,I1235212,I1235229,I1235246,I1235291,I1235322,I1235339,I1235365,I1235373,I1235404,I1235421,I1235438,I1235455,I1235527,I1235553,I1235561,I1235601,I1235609,I1235626,I1235643,I1235683,I1235705,I1235722,I1235748,I1235756,I1235773,I1235790,I1235807,I1235824,I1235869,I1235900,I1235917,I1235943,I1235951,I1235982,I1235999,I1236016,I1236033,I1236105,I1236131,I1236139,I1236179,I1236187,I1236204,I1236221,I1236261,I1236283,I1236300,I1236326,I1236334,I1236351,I1236368,I1236385,I1236402,I1236447,I1236478,I1236495,I1236521,I1236529,I1236560,I1236577,I1236594,I1236611,I1236683,I1327533,I1236709,I1236717,I1327560,I1327542,I1236757,I1236765,I1327551,I1236782,I1327554,I1236799,I1236839,I1236861,I1327548,I1236878,I1236904,I1236912,I1236929,I1327536,I1236946,I1327539,I1236963,I1236980,I1237025,I1327557,I1237056,I1237073,I1327545,I1237099,I1237107,I1237138,I1237155,I1237172,I1237189,I1237261,I1237287,I1237295,I1237335,I1237343,I1237360,I1237377,I1237417,I1237439,I1237456,I1237482,I1237490,I1237507,I1237524,I1237541,I1237558,I1237603,I1237634,I1237651,I1237677,I1237685,I1237716,I1237733,I1237750,I1237767,I1237839,I1237865,I1237873,I1237913,I1237921,I1237938,I1237955,I1237995,I1238017,I1238034,I1238060,I1238068,I1238085,I1238102,I1238119,I1238136,I1238181,I1238212,I1238229,I1238255,I1238263,I1238294,I1238311,I1238328,I1238345,I1238417,I1238443,I1238451,I1238491,I1238499,I1238516,I1238533,I1238573,I1238595,I1238612,I1238638,I1238646,I1238663,I1238680,I1238697,I1238714,I1238759,I1238790,I1238807,I1238833,I1238841,I1238872,I1238889,I1238906,I1238923,I1238995,I1239021,I1239029,I1239069,I1239077,I1239094,I1239111,I1239151,I1239173,I1239190,I1239216,I1239224,I1239241,I1239258,I1239275,I1239292,I1239337,I1239368,I1239385,I1239411,I1239419,I1239450,I1239467,I1239484,I1239501,I1239573,I1239599,I1239607,I1239647,I1239655,I1239672,I1239689,I1239729,I1239751,I1239768,I1239794,I1239802,I1239819,I1239836,I1239853,I1239870,I1239915,I1239946,I1239963,I1239989,I1239997,I1240028,I1240045,I1240062,I1240079,I1240151,I1240177,I1240185,I1240225,I1240233,I1240250,I1240267,I1240307,I1240329,I1240346,I1240372,I1240380,I1240397,I1240414,I1240431,I1240448,I1240493,I1240524,I1240541,I1240567,I1240575,I1240606,I1240623,I1240640,I1240657,I1240729,I1240755,I1240763,I1240803,I1240811,I1240828,I1240845,I1240885,I1240907,I1240924,I1240950,I1240958,I1240975,I1240992,I1241009,I1241026,I1241071,I1241102,I1241119,I1241145,I1241153,I1241184,I1241201,I1241218,I1241235,I1241307,I1241333,I1241341,I1241381,I1241389,I1241406,I1241423,I1241463,I1241485,I1241502,I1241528,I1241536,I1241553,I1241570,I1241587,I1241604,I1241649,I1241680,I1241697,I1241723,I1241731,I1241762,I1241779,I1241796,I1241813,I1241885,I1241911,I1241919,I1241959,I1241967,I1241984,I1242001,I1242041,I1242063,I1242080,I1242106,I1242114,I1242131,I1242148,I1242165,I1242182,I1242227,I1242258,I1242275,I1242301,I1242309,I1242340,I1242357,I1242374,I1242391,I1242463,I1242489,I1242497,I1242537,I1242545,I1242562,I1242579,I1242619,I1242641,I1242658,I1242684,I1242692,I1242709,I1242726,I1242743,I1242760,I1242805,I1242836,I1242853,I1242879,I1242887,I1242918,I1242935,I1242952,I1242969,I1243041,I1243067,I1243075,I1243115,I1243123,I1243140,I1243157,I1243197,I1243219,I1243236,I1243262,I1243270,I1243287,I1243304,I1243321,I1243338,I1243383,I1243414,I1243431,I1243457,I1243465,I1243496,I1243513,I1243530,I1243547,I1243619,I1243645,I1243653,I1243693,I1243701,I1243718,I1243735,I1243775,I1243797,I1243814,I1243840,I1243848,I1243865,I1243882,I1243899,I1243916,I1243961,I1243992,I1244009,I1244035,I1244043,I1244074,I1244091,I1244108,I1244125,I1244197,I1317255,I1244223,I1244231,I1317237,I1317246,I1244271,I1244279,I1317231,I1244296,I1317243,I1244313,I1244353,I1244375,I1317234,I1244392,I1244418,I1244426,I1244443,I1244460,I1244477,I1244494,I1244539,I1317252,I1244570,I1244587,I1317240,I1317249,I1244613,I1244621,I1244652,I1244669,I1244686,I1244703,I1244775,I1244801,I1244809,I1244849,I1244857,I1244874,I1244891,I1244931,I1244953,I1244970,I1244996,I1245004,I1245021,I1245038,I1245055,I1245072,I1245117,I1245148,I1245165,I1245191,I1245199,I1245230,I1245247,I1245264,I1245281,I1245353,I1324755,I1245379,I1245387,I1324740,I1324752,I1245413,I1245430,I1245452,I1324746,I1245469,I1324737,I1245486,I1324731,I1245503,I1245520,I1245551,I1324743,I1245568,I1324728,I1245585,I1324749,I1245602,I1245647,I1324734,I1245664,I1245681,I1245740,I1245766,I1245774,I1245791,I1245808,I1245839,I1245897,I1245923,I1245931,I1245957,I1245974,I1245996,I1246013,I1246030,I1246047,I1246064,I1246095,I1246112,I1246129,I1246146,I1246191,I1246208,I1246225,I1246284,I1246310,I1246318,I1246335,I1246352,I1246383,I1246441,I1246467,I1246475,I1246501,I1246518,I1246540,I1246557,I1246574,I1246591,I1246608,I1246639,I1246656,I1246673,I1246690,I1246735,I1246752,I1246769,I1246828,I1246854,I1246862,I1246879,I1246896,I1246927,I1246985,I1247011,I1247019,I1247045,I1247062,I1247084,I1247101,I1247118,I1247135,I1247152,I1247183,I1247200,I1247217,I1247234,I1247279,I1247296,I1247313,I1247372,I1247398,I1247406,I1247423,I1247440,I1247471,I1247529,I1247555,I1247563,I1247589,I1247606,I1247628,I1247645,I1247662,I1247679,I1247696,I1247727,I1247744,I1247761,I1247778,I1247823,I1247840,I1247857,I1247916,I1247942,I1247950,I1247967,I1247984,I1248015,I1248073,I1248099,I1248107,I1248133,I1248150,I1248172,I1248189,I1248206,I1248223,I1248240,I1248271,I1248288,I1248305,I1248322,I1248367,I1248384,I1248401,I1248460,I1248486,I1248494,I1248511,I1248528,I1248559,I1248617,I1248643,I1248651,I1248677,I1248694,I1248716,I1248733,I1248750,I1248767,I1248784,I1248815,I1248832,I1248849,I1248866,I1248911,I1248928,I1248945,I1249004,I1249030,I1249038,I1249055,I1249072,I1249103,I1249161,I1249187,I1249195,I1249221,I1249238,I1249260,I1249277,I1249294,I1249311,I1249328,I1249359,I1249376,I1249393,I1249410,I1249455,I1249472,I1249489,I1249548,I1249574,I1249582,I1249599,I1249616,I1249647,I1249705,I1249731,I1249739,I1249765,I1249782,I1249804,I1249821,I1249838,I1249855,I1249872,I1249903,I1249920,I1249937,I1249954,I1249999,I1250016,I1250033,I1250092,I1250118,I1250126,I1250143,I1250160,I1250191,I1250249,I1250275,I1250283,I1250309,I1250326,I1250348,I1250365,I1250382,I1250399,I1250416,I1250447,I1250464,I1250481,I1250498,I1250543,I1250560,I1250577,I1250636,I1250662,I1250670,I1250687,I1250704,I1250735,I1250793,I1250819,I1250827,I1250853,I1250870,I1250892,I1250909,I1250926,I1250943,I1250960,I1250991,I1251008,I1251025,I1251042,I1251087,I1251104,I1251121,I1251180,I1251206,I1251214,I1251231,I1251248,I1251279,I1251337,I1251363,I1251371,I1251397,I1251414,I1251436,I1251453,I1251470,I1251487,I1251504,I1251535,I1251552,I1251569,I1251586,I1251631,I1251648,I1251665,I1251724,I1251750,I1251758,I1251775,I1251792,I1251823,I1251881,I1251907,I1251915,I1251941,I1251958,I1251980,I1251997,I1252014,I1252031,I1252048,I1252079,I1252096,I1252113,I1252130,I1252175,I1252192,I1252209,I1252268,I1252294,I1252302,I1252319,I1252336,I1252367,I1252425,I1252451,I1252459,I1252485,I1252502,I1252417,I1252524,I1252541,I1252558,I1252575,I1252592,I1252396,I1252623,I1252640,I1252657,I1252674,I1252399,I1252414,I1252719,I1252736,I1252753,I1252411,I1252408,I1252405,I1252812,I1252838,I1252846,I1252863,I1252880,I1252393,I1252911,I1252402,I1252969,I1252995,I1253003,I1253029,I1253046,I1253068,I1253085,I1253102,I1253119,I1253136,I1253167,I1253184,I1253201,I1253218,I1253263,I1253280,I1253297,I1253356,I1253382,I1253390,I1253407,I1253424,I1253455,I1253513,I1253539,I1253547,I1253573,I1253590,I1253612,I1253629,I1253646,I1253663,I1253680,I1253711,I1253728,I1253745,I1253762,I1253807,I1253824,I1253841,I1253900,I1253926,I1253934,I1253951,I1253968,I1253999,I1254057,I1254083,I1254091,I1254117,I1254134,I1254049,I1254156,I1254173,I1254190,I1254207,I1254224,I1254028,I1254255,I1254272,I1254289,I1254306,I1254031,I1254046,I1254351,I1254368,I1254385,I1254043,I1254040,I1254037,I1254444,I1254470,I1254478,I1254495,I1254512,I1254025,I1254543,I1254034,I1254601,I1254627,I1254635,I1254661,I1254678,I1254700,I1254717,I1254734,I1254751,I1254768,I1254799,I1254816,I1254833,I1254850,I1254895,I1254912,I1254929,I1254988,I1255014,I1255022,I1255039,I1255056,I1255087,I1255145,I1255171,I1255179,I1255205,I1255222,I1255244,I1255261,I1255278,I1255295,I1255312,I1255343,I1255360,I1255377,I1255394,I1255439,I1255456,I1255473,I1255532,I1255558,I1255566,I1255583,I1255600,I1255631,I1255689,I1255715,I1255723,I1255749,I1255766,I1255788,I1255805,I1255822,I1255839,I1255856,I1255887,I1255904,I1255921,I1255938,I1255983,I1256000,I1256017,I1256076,I1256102,I1256110,I1256127,I1256144,I1256175,I1256233,I1256259,I1256267,I1256293,I1256310,I1256332,I1256349,I1256366,I1256383,I1256400,I1256431,I1256448,I1256465,I1256482,I1256527,I1256544,I1256561,I1256620,I1256646,I1256654,I1256671,I1256688,I1256719,I1256777,I1256803,I1256811,I1256837,I1256854,I1256876,I1256893,I1256910,I1256927,I1256944,I1256975,I1256992,I1257009,I1257026,I1257071,I1257088,I1257105,I1257164,I1257190,I1257198,I1257215,I1257232,I1257263,I1257321,I1373800,I1257347,I1257355,I1373785,I1373779,I1257381,I1257398,I1257313,I1257420,I1373773,I1257437,I1373794,I1257454,I1373782,I1257471,I1257488,I1257292,I1257519,I1373791,I1257536,I1373797,I1257553,I1373788,I1257570,I1257295,I1257310,I1257615,I1373776,I1257632,I1257649,I1257307,I1257304,I1257301,I1257708,I1257734,I1257742,I1257759,I1257776,I1257289,I1257807,I1257298,I1257865,I1257891,I1257899,I1257925,I1257942,I1257964,I1257981,I1257998,I1258015,I1258032,I1258063,I1258080,I1258097,I1258114,I1258159,I1258176,I1258193,I1258252,I1258278,I1258286,I1258303,I1258320,I1258351,I1258409,I1258435,I1258443,I1258469,I1258486,I1258508,I1258525,I1258542,I1258559,I1258576,I1258607,I1258624,I1258641,I1258658,I1258703,I1258720,I1258737,I1258796,I1258822,I1258830,I1258847,I1258864,I1258895,I1258953,I1258979,I1258987,I1259013,I1259030,I1259052,I1259069,I1259086,I1259103,I1259120,I1259151,I1259168,I1259185,I1259202,I1259247,I1259264,I1259281,I1259340,I1259366,I1259374,I1259391,I1259408,I1259439,I1259497,I1259523,I1259531,I1259557,I1259574,I1259596,I1259613,I1259630,I1259647,I1259664,I1259695,I1259712,I1259729,I1259746,I1259791,I1259808,I1259825,I1259884,I1259910,I1259918,I1259935,I1259952,I1259983,I1260041,I1260067,I1260075,I1260101,I1260118,I1260140,I1260157,I1260174,I1260191,I1260208,I1260239,I1260256,I1260273,I1260290,I1260335,I1260352,I1260369,I1260428,I1260454,I1260462,I1260479,I1260496,I1260527,I1260585,I1260611,I1260619,I1260645,I1260662,I1260684,I1260701,I1260718,I1260735,I1260752,I1260783,I1260800,I1260817,I1260834,I1260879,I1260896,I1260913,I1260972,I1260998,I1261006,I1261023,I1261040,I1261071,I1261129,I1261155,I1261163,I1261189,I1261206,I1261228,I1261245,I1261262,I1261279,I1261296,I1261327,I1261344,I1261361,I1261378,I1261423,I1261440,I1261457,I1261516,I1261542,I1261550,I1261567,I1261584,I1261615,I1261673,I1261699,I1261707,I1261733,I1261750,I1261772,I1261789,I1261806,I1261823,I1261840,I1261871,I1261888,I1261905,I1261922,I1261967,I1261984,I1262001,I1262060,I1262086,I1262094,I1262111,I1262128,I1262159,I1262217,I1262243,I1262251,I1262277,I1262294,I1262316,I1262333,I1262350,I1262367,I1262384,I1262415,I1262432,I1262449,I1262466,I1262511,I1262528,I1262545,I1262604,I1262630,I1262638,I1262655,I1262672,I1262703,I1262761,I1262787,I1262795,I1262821,I1262838,I1262860,I1262877,I1262894,I1262911,I1262928,I1262959,I1262976,I1262993,I1263010,I1263055,I1263072,I1263089,I1263148,I1263174,I1263182,I1263199,I1263216,I1263247,I1263305,I1263331,I1263339,I1263365,I1263382,I1263404,I1263421,I1263438,I1263455,I1263472,I1263503,I1263520,I1263537,I1263554,I1263599,I1263616,I1263633,I1263692,I1263718,I1263726,I1263743,I1263760,I1263791,I1263849,I1263875,I1263883,I1263909,I1263926,I1263948,I1263965,I1263982,I1263999,I1264016,I1264047,I1264064,I1264081,I1264098,I1264143,I1264160,I1264177,I1264236,I1264262,I1264270,I1264287,I1264304,I1264335,I1264393,I1264419,I1264427,I1264453,I1264470,I1264492,I1264509,I1264526,I1264543,I1264560,I1264591,I1264608,I1264625,I1264642,I1264687,I1264704,I1264721,I1264780,I1264806,I1264814,I1264831,I1264848,I1264879,I1264937,I1264963,I1264971,I1264997,I1265014,I1265036,I1265053,I1265070,I1265087,I1265104,I1265135,I1265152,I1265169,I1265186,I1265231,I1265248,I1265265,I1265324,I1265350,I1265358,I1265375,I1265392,I1265423,I1265481,I1265507,I1265515,I1265541,I1265558,I1265580,I1265597,I1265614,I1265631,I1265648,I1265679,I1265696,I1265713,I1265730,I1265775,I1265792,I1265809,I1265868,I1265894,I1265902,I1265919,I1265936,I1265967,I1266025,I1266051,I1266059,I1266085,I1266102,I1266124,I1266141,I1266158,I1266175,I1266192,I1266223,I1266240,I1266257,I1266274,I1266319,I1266336,I1266353,I1266412,I1266438,I1266446,I1266463,I1266480,I1266511,I1266569,I1266595,I1266603,I1266629,I1266646,I1266668,I1266685,I1266702,I1266719,I1266736,I1266767,I1266784,I1266801,I1266818,I1266863,I1266880,I1266897,I1266956,I1266982,I1266990,I1267007,I1267024,I1267055,I1267113,I1267139,I1267147,I1267173,I1267190,I1267212,I1267229,I1267246,I1267263,I1267280,I1267311,I1267328,I1267345,I1267362,I1267407,I1267424,I1267441,I1267500,I1267526,I1267534,I1267551,I1267568,I1267599,I1267657,I1267683,I1267691,I1267717,I1267734,I1267756,I1267773,I1267790,I1267807,I1267824,I1267855,I1267872,I1267889,I1267906,I1267951,I1267968,I1267985,I1268044,I1268070,I1268078,I1268095,I1268112,I1268143,I1268201,I1268227,I1268235,I1268261,I1268278,I1268300,I1268317,I1268334,I1268351,I1268368,I1268399,I1268416,I1268433,I1268450,I1268495,I1268512,I1268529,I1268588,I1268614,I1268622,I1268639,I1268656,I1268687,I1268745,I1268771,I1268779,I1268805,I1268822,I1268737,I1268844,I1268861,I1268878,I1268895,I1268912,I1268716,I1268943,I1268960,I1268977,I1268994,I1268719,I1268734,I1269039,I1269056,I1269073,I1268731,I1268728,I1268725,I1269132,I1269158,I1269166,I1269183,I1269200,I1268713,I1269231,I1268722,I1269289,I1269315,I1269323,I1269349,I1269366,I1269388,I1269405,I1269422,I1269439,I1269456,I1269487,I1269504,I1269521,I1269538,I1269583,I1269600,I1269617,I1269676,I1269702,I1269710,I1269727,I1269744,I1269775,I1269833,I1269859,I1269867,I1269893,I1269910,I1269932,I1269949,I1269966,I1269983,I1270000,I1270031,I1270048,I1270065,I1270082,I1270127,I1270144,I1270161,I1270220,I1270246,I1270254,I1270271,I1270288,I1270319,I1270377,I1270403,I1270411,I1270437,I1270454,I1270476,I1270493,I1270510,I1270527,I1270544,I1270575,I1270592,I1270609,I1270626,I1270671,I1270688,I1270705,I1270764,I1270790,I1270798,I1270815,I1270832,I1270863,I1270921,I1270947,I1270955,I1270981,I1270998,I1271020,I1271037,I1271054,I1271071,I1271088,I1271119,I1271136,I1271153,I1271170,I1271215,I1271232,I1271249,I1271308,I1271334,I1271342,I1271359,I1271376,I1271407,I1271465,I1271491,I1271499,I1271525,I1271542,I1271564,I1271581,I1271598,I1271615,I1271632,I1271663,I1271680,I1271697,I1271714,I1271759,I1271776,I1271793,I1271852,I1271878,I1271886,I1271903,I1271920,I1271951,I1272009,I1272035,I1272043,I1272069,I1272086,I1272108,I1272125,I1272142,I1272159,I1272176,I1272207,I1272224,I1272241,I1272258,I1272303,I1272320,I1272337,I1272396,I1272422,I1272430,I1272447,I1272464,I1272495,I1272553,I1406525,I1272579,I1272587,I1406510,I1406504,I1272613,I1272630,I1272545,I1272652,I1406498,I1272669,I1406519,I1272686,I1406507,I1272703,I1272720,I1272524,I1272751,I1406516,I1272768,I1406522,I1272785,I1406513,I1272802,I1272527,I1272542,I1272847,I1406501,I1272864,I1272881,I1272539,I1272536,I1272533,I1272940,I1272966,I1272974,I1272991,I1273008,I1272521,I1273039,I1272530,I1273097,I1273123,I1273131,I1273157,I1273174,I1273196,I1273213,I1273230,I1273247,I1273264,I1273295,I1273312,I1273329,I1273346,I1273391,I1273408,I1273425,I1273484,I1273510,I1273518,I1273535,I1273552,I1273583,I1273641,I1273667,I1273675,I1273701,I1273718,I1273740,I1273757,I1273774,I1273791,I1273808,I1273839,I1273856,I1273873,I1273890,I1273935,I1273952,I1273969,I1274028,I1274054,I1274062,I1274079,I1274096,I1274127,I1274185,I1274211,I1274219,I1274245,I1274262,I1274284,I1274301,I1274318,I1274335,I1274352,I1274383,I1274400,I1274417,I1274434,I1274479,I1274496,I1274513,I1274572,I1274598,I1274606,I1274623,I1274640,I1274671,I1274729,I1274755,I1274763,I1274789,I1274806,I1274828,I1274845,I1274862,I1274879,I1274896,I1274927,I1274944,I1274961,I1274978,I1275023,I1275040,I1275057,I1275116,I1275142,I1275150,I1275167,I1275184,I1275215,I1275273,I1275299,I1275307,I1275333,I1275350,I1275372,I1275389,I1275406,I1275423,I1275440,I1275471,I1275488,I1275505,I1275522,I1275567,I1275584,I1275601,I1275660,I1275686,I1275694,I1275711,I1275728,I1275759,I1275817,I1275843,I1275851,I1275877,I1275894,I1275916,I1275933,I1275950,I1275967,I1275984,I1276015,I1276032,I1276049,I1276066,I1276111,I1276128,I1276145,I1276204,I1276230,I1276238,I1276255,I1276272,I1276303,I1276361,I1276387,I1276395,I1276421,I1276438,I1276460,I1276477,I1276494,I1276511,I1276528,I1276559,I1276576,I1276593,I1276610,I1276655,I1276672,I1276689,I1276748,I1276774,I1276782,I1276799,I1276816,I1276847,I1276905,I1276931,I1276939,I1276965,I1276982,I1277004,I1277021,I1277038,I1277055,I1277072,I1277103,I1277120,I1277137,I1277154,I1277199,I1277216,I1277233,I1277292,I1277318,I1277326,I1277343,I1277360,I1277391,I1277449,I1277475,I1277483,I1277509,I1277526,I1277548,I1277565,I1277582,I1277599,I1277616,I1277647,I1277664,I1277681,I1277698,I1277743,I1277760,I1277777,I1277836,I1277862,I1277870,I1277887,I1277904,I1277935,I1277993,I1278019,I1278027,I1278053,I1278070,I1278092,I1278109,I1278126,I1278143,I1278160,I1278191,I1278208,I1278225,I1278242,I1278287,I1278304,I1278321,I1278380,I1278406,I1278414,I1278431,I1278448,I1278479,I1278537,I1278563,I1278571,I1278597,I1278614,I1278636,I1278653,I1278670,I1278687,I1278704,I1278735,I1278752,I1278769,I1278786,I1278831,I1278848,I1278865,I1278924,I1278950,I1278958,I1278975,I1278992,I1279023,I1279081,I1279107,I1279115,I1279141,I1279158,I1279180,I1279197,I1279214,I1279231,I1279248,I1279279,I1279296,I1279313,I1279330,I1279375,I1279392,I1279409,I1279468,I1279494,I1279502,I1279519,I1279536,I1279567,I1279625,I1279651,I1279659,I1279685,I1279702,I1279724,I1279741,I1279758,I1279775,I1279792,I1279823,I1279840,I1279857,I1279874,I1279919,I1279936,I1279953,I1280012,I1280038,I1280046,I1280063,I1280080,I1280111,I1280169,I1326438,I1280195,I1280203,I1326423,I1326435,I1280229,I1280246,I1280268,I1326429,I1280285,I1326420,I1280302,I1326414,I1280319,I1280336,I1280367,I1326426,I1280384,I1326411,I1280401,I1326432,I1280418,I1280463,I1326417,I1280480,I1280497,I1280556,I1280582,I1280590,I1280607,I1280624,I1280655,I1280713,I1280739,I1280747,I1280773,I1280790,I1280812,I1280829,I1280846,I1280863,I1280880,I1280911,I1280928,I1280945,I1280962,I1281007,I1281024,I1281041,I1281100,I1281126,I1281134,I1281151,I1281168,I1281199,I1281257,I1281283,I1281291,I1281317,I1281334,I1281249,I1281356,I1281373,I1281390,I1281407,I1281424,I1281228,I1281455,I1281472,I1281489,I1281506,I1281231,I1281246,I1281551,I1281568,I1281585,I1281243,I1281240,I1281237,I1281644,I1281670,I1281678,I1281695,I1281712,I1281225,I1281743,I1281234,I1281801,I1281827,I1281835,I1281861,I1281878,I1281900,I1281917,I1281934,I1281951,I1281968,I1281999,I1282016,I1282033,I1282050,I1282095,I1282112,I1282129,I1282188,I1282214,I1282222,I1282239,I1282256,I1282287,I1282345,I1282371,I1282379,I1282405,I1282422,I1282444,I1282461,I1282478,I1282495,I1282512,I1282543,I1282560,I1282577,I1282594,I1282639,I1282656,I1282673,I1282732,I1282758,I1282766,I1282783,I1282800,I1282831,I1282889,I1282915,I1282923,I1282949,I1282966,I1282988,I1283005,I1283022,I1283039,I1283056,I1283087,I1283104,I1283121,I1283138,I1283183,I1283200,I1283217,I1283276,I1283302,I1283310,I1283327,I1283344,I1283375,I1283433,I1398195,I1283459,I1283467,I1398180,I1398174,I1283493,I1283510,I1283425,I1283532,I1398168,I1283549,I1398189,I1283566,I1398177,I1283583,I1283600,I1283404,I1283631,I1398186,I1283648,I1398192,I1283665,I1398183,I1283682,I1283407,I1283422,I1283727,I1398171,I1283744,I1283761,I1283419,I1283416,I1283413,I1283820,I1283846,I1283854,I1283871,I1283888,I1283401,I1283919,I1283410,I1283977,I1284003,I1284011,I1284037,I1284054,I1284076,I1284093,I1284110,I1284127,I1284144,I1284175,I1284192,I1284209,I1284226,I1284271,I1284288,I1284305,I1284364,I1284390,I1284398,I1284415,I1284432,I1284463,I1284521,I1284547,I1284555,I1284581,I1284598,I1284620,I1284637,I1284654,I1284671,I1284688,I1284719,I1284736,I1284753,I1284770,I1284815,I1284832,I1284849,I1284908,I1284934,I1284942,I1284959,I1284976,I1285007,I1285065,I1285091,I1285099,I1285125,I1285142,I1285164,I1285181,I1285198,I1285215,I1285232,I1285263,I1285280,I1285297,I1285314,I1285359,I1285376,I1285393,I1285452,I1285478,I1285486,I1285503,I1285520,I1285551,I1285609,I1285635,I1285643,I1285669,I1285686,I1285708,I1285725,I1285742,I1285759,I1285776,I1285807,I1285824,I1285841,I1285858,I1285903,I1285920,I1285937,I1285996,I1286022,I1286030,I1286047,I1286064,I1286095,I1286153,I1286179,I1286187,I1286213,I1286230,I1286252,I1286269,I1286286,I1286303,I1286320,I1286351,I1286368,I1286385,I1286402,I1286447,I1286464,I1286481,I1286540,I1286566,I1286574,I1286591,I1286608,I1286639,I1286697,I1286723,I1286731,I1286757,I1286774,I1286796,I1286813,I1286830,I1286847,I1286864,I1286895,I1286912,I1286929,I1286946,I1286991,I1287008,I1287025,I1287084,I1287110,I1287118,I1287135,I1287152,I1287183,I1287241,I1287267,I1287275,I1287301,I1287318,I1287340,I1287357,I1287374,I1287391,I1287408,I1287439,I1287456,I1287473,I1287490,I1287535,I1287552,I1287569,I1287628,I1287654,I1287662,I1287679,I1287696,I1287727,I1287785,I1287811,I1287819,I1287836,I1287862,I1287870,I1287887,I1287904,I1287921,I1287938,I1287969,I1287986,I1288003,I1288034,I1288051,I1288091,I1288099,I1288130,I1288147,I1288164,I1288181,I1288212,I1288243,I1288269,I1288291,I1288363,I1288389,I1288397,I1288414,I1288440,I1288448,I1288465,I1288482,I1288499,I1288516,I1288547,I1288564,I1288581,I1288612,I1288629,I1288669,I1288677,I1288708,I1288725,I1288742,I1288759,I1288790,I1288821,I1288847,I1288869,I1288941,I1288967,I1288975,I1288992,I1289018,I1289026,I1289043,I1289060,I1289077,I1289094,I1289125,I1289142,I1289159,I1289190,I1289207,I1289247,I1289255,I1289286,I1289303,I1289320,I1289337,I1289368,I1289399,I1289425,I1289447,I1289519,I1289545,I1289553,I1289570,I1289596,I1289604,I1289621,I1289638,I1289655,I1289672,I1289703,I1289720,I1289737,I1289768,I1289785,I1289825,I1289833,I1289864,I1289881,I1289898,I1289915,I1289946,I1289977,I1290003,I1290025,I1290097,I1290123,I1290131,I1290148,I1290174,I1290182,I1290199,I1290216,I1290233,I1290250,I1290281,I1290298,I1290315,I1290346,I1290363,I1290403,I1290411,I1290442,I1290459,I1290476,I1290493,I1290524,I1290555,I1290581,I1290603,I1290675,I1290701,I1290709,I1290726,I1290752,I1290760,I1290777,I1290794,I1290811,I1290828,I1290859,I1290876,I1290893,I1290924,I1290941,I1290981,I1290989,I1291020,I1291037,I1291054,I1291071,I1291102,I1291133,I1291159,I1291181,I1291253,I1291279,I1291287,I1291304,I1291330,I1291338,I1291355,I1291372,I1291389,I1291406,I1291437,I1291454,I1291471,I1291502,I1291519,I1291559,I1291567,I1291598,I1291615,I1291632,I1291649,I1291680,I1291711,I1291737,I1291759,I1291831,I1384507,I1291857,I1291865,I1384498,I1291882,I1384483,I1291908,I1291916,I1291933,I1384486,I1291950,I1384495,I1291967,I1291984,I1384492,I1291823,I1292015,I1384504,I1292032,I1292049,I1291802,I1292080,I1384489,I1292097,I1291808,I1292137,I1292145,I1291817,I1292176,I1384510,I1292193,I1292210,I1292227,I1291820,I1292258,I1291799,I1292289,I1384501,I1292315,I1291814,I1292337,I1291811,I1291805,I1292409,I1292435,I1292443,I1292460,I1292486,I1292494,I1292511,I1292528,I1292545,I1292562,I1292593,I1292610,I1292627,I1292658,I1292675,I1292715,I1292723,I1292754,I1292771,I1292788,I1292805,I1292836,I1292867,I1292893,I1292915,I1292987,I1293013,I1293021,I1293038,I1293064,I1293072,I1293089,I1293106,I1293123,I1293140,I1293171,I1293188,I1293205,I1293236,I1293253,I1293293,I1293301,I1293332,I1293349,I1293366,I1293383,I1293414,I1293445,I1293471,I1293493,I1293565,I1293591,I1293599,I1293616,I1293642,I1293650,I1293667,I1293684,I1293701,I1293718,I1293749,I1293766,I1293783,I1293814,I1293831,I1293871,I1293879,I1293910,I1293927,I1293944,I1293961,I1293992,I1294023,I1294049,I1294071,I1294143,I1294169,I1294177,I1294194,I1294220,I1294228,I1294245,I1294262,I1294279,I1294296,I1294327,I1294344,I1294361,I1294392,I1294409,I1294449,I1294457,I1294488,I1294505,I1294522,I1294539,I1294570,I1294601,I1294627,I1294649,I1294721,I1294747,I1294755,I1294772,I1294798,I1294806,I1294823,I1294840,I1294857,I1294874,I1294905,I1294922,I1294939,I1294970,I1294987,I1295027,I1295035,I1295066,I1295083,I1295100,I1295117,I1295148,I1295179,I1295205,I1295227,I1295299,I1295325,I1295333,I1295350,I1295376,I1295384,I1295401,I1295418,I1295435,I1295452,I1295483,I1295500,I1295517,I1295548,I1295565,I1295605,I1295613,I1295644,I1295661,I1295678,I1295695,I1295726,I1295757,I1295783,I1295805,I1295877,I1295903,I1295911,I1295928,I1295954,I1295962,I1295979,I1295996,I1296013,I1296030,I1296061,I1296078,I1296095,I1296126,I1296143,I1296183,I1296191,I1296222,I1296239,I1296256,I1296273,I1296304,I1296335,I1296361,I1296383,I1296455,I1296481,I1296489,I1296506,I1296532,I1296540,I1296557,I1296574,I1296591,I1296608,I1296447,I1296639,I1296656,I1296673,I1296426,I1296704,I1296721,I1296432,I1296761,I1296769,I1296441,I1296800,I1296817,I1296834,I1296851,I1296444,I1296882,I1296423,I1296913,I1296939,I1296438,I1296961,I1296435,I1296429,I1297033,I1297059,I1297067,I1297084,I1297110,I1297118,I1297135,I1297152,I1297169,I1297186,I1297217,I1297234,I1297251,I1297282,I1297299,I1297339,I1297347,I1297378,I1297395,I1297412,I1297429,I1297460,I1297491,I1297517,I1297539,I1297611,I1297637,I1297645,I1297662,I1297688,I1297696,I1297713,I1297730,I1297747,I1297764,I1297795,I1297812,I1297829,I1297860,I1297877,I1297917,I1297925,I1297956,I1297973,I1297990,I1298007,I1298038,I1298069,I1298095,I1298117,I1298189,I1298215,I1298223,I1298240,I1298266,I1298274,I1298291,I1298308,I1298325,I1298342,I1298373,I1298390,I1298407,I1298438,I1298455,I1298495,I1298503,I1298534,I1298551,I1298568,I1298585,I1298616,I1298647,I1298673,I1298695,I1298767,I1298793,I1298801,I1298818,I1298844,I1298852,I1298869,I1298886,I1298903,I1298920,I1298951,I1298968,I1298985,I1299016,I1299033,I1299073,I1299081,I1299112,I1299129,I1299146,I1299163,I1299194,I1299225,I1299251,I1299273,I1299345,I1299371,I1299379,I1299396,I1299422,I1299430,I1299447,I1299464,I1299481,I1299498,I1299529,I1299546,I1299563,I1299594,I1299611,I1299651,I1299659,I1299690,I1299707,I1299724,I1299741,I1299772,I1299803,I1299829,I1299851,I1299923,I1299949,I1299957,I1299974,I1300000,I1300008,I1300025,I1300042,I1300059,I1300076,I1300107,I1300124,I1300141,I1300172,I1300189,I1300229,I1300237,I1300268,I1300285,I1300302,I1300319,I1300350,I1300381,I1300407,I1300429,I1300501,I1300527,I1300535,I1300552,I1300578,I1300586,I1300603,I1300620,I1300637,I1300654,I1300685,I1300702,I1300719,I1300750,I1300767,I1300807,I1300815,I1300846,I1300863,I1300880,I1300897,I1300928,I1300959,I1300985,I1301007,I1301079,I1301105,I1301113,I1301130,I1301156,I1301164,I1301181,I1301198,I1301215,I1301232,I1301263,I1301280,I1301297,I1301328,I1301345,I1301385,I1301393,I1301424,I1301441,I1301458,I1301475,I1301506,I1301537,I1301563,I1301585,I1301657,I1301683,I1301691,I1301708,I1301734,I1301742,I1301759,I1301776,I1301793,I1301810,I1301841,I1301858,I1301875,I1301906,I1301923,I1301963,I1301971,I1302002,I1302019,I1302036,I1302053,I1302084,I1302115,I1302141,I1302163,I1302235,I1302261,I1302269,I1302286,I1302312,I1302320,I1302337,I1302354,I1302371,I1302388,I1302419,I1302436,I1302453,I1302484,I1302501,I1302541,I1302549,I1302580,I1302597,I1302614,I1302631,I1302662,I1302693,I1302719,I1302741,I1302813,I1302839,I1302847,I1302864,I1302890,I1302898,I1302915,I1302932,I1302949,I1302966,I1302805,I1302997,I1303014,I1303031,I1302784,I1303062,I1303079,I1302790,I1303119,I1303127,I1302799,I1303158,I1303175,I1303192,I1303209,I1302802,I1303240,I1302781,I1303271,I1303297,I1302796,I1303319,I1302793,I1302787,I1303391,I1303417,I1303425,I1303442,I1303468,I1303476,I1303493,I1303510,I1303527,I1303544,I1303575,I1303592,I1303609,I1303640,I1303657,I1303697,I1303705,I1303736,I1303753,I1303770,I1303787,I1303818,I1303849,I1303875,I1303897,I1303969,I1303995,I1304003,I1304020,I1304046,I1304054,I1304071,I1304088,I1304105,I1304122,I1304153,I1304170,I1304187,I1304218,I1304235,I1304275,I1304283,I1304314,I1304331,I1304348,I1304365,I1304396,I1304427,I1304453,I1304475,I1304547,I1304573,I1304581,I1304598,I1304624,I1304632,I1304649,I1304666,I1304683,I1304700,I1304731,I1304748,I1304765,I1304796,I1304813,I1304853,I1304861,I1304892,I1304909,I1304926,I1304943,I1304974,I1305005,I1305031,I1305053,I1305125,I1305151,I1305159,I1305176,I1305202,I1305210,I1305227,I1305244,I1305261,I1305278,I1305309,I1305326,I1305343,I1305374,I1305391,I1305431,I1305439,I1305470,I1305487,I1305504,I1305521,I1305552,I1305583,I1305609,I1305631,I1305703,I1305729,I1305737,I1305754,I1305780,I1305788,I1305805,I1305822,I1305839,I1305856,I1305695,I1305887,I1305904,I1305921,I1305674,I1305952,I1305969,I1305680,I1306009,I1306017,I1305689,I1306048,I1306065,I1306082,I1306099,I1305692,I1306130,I1305671,I1306161,I1306187,I1305686,I1306209,I1305683,I1305677,I1306281,I1306307,I1306315,I1306332,I1306358,I1306366,I1306383,I1306400,I1306417,I1306434,I1306465,I1306482,I1306499,I1306530,I1306547,I1306587,I1306595,I1306626,I1306643,I1306660,I1306677,I1306708,I1306739,I1306765,I1306787,I1306859,I1306885,I1306893,I1306910,I1306936,I1306944,I1306961,I1306978,I1306995,I1307012,I1307043,I1307060,I1307077,I1307108,I1307125,I1307165,I1307173,I1307204,I1307221,I1307238,I1307255,I1307286,I1307317,I1307343,I1307365,I1307437,I1307463,I1307471,I1307488,I1307514,I1307522,I1307539,I1307556,I1307573,I1307590,I1307621,I1307638,I1307655,I1307686,I1307703,I1307743,I1307751,I1307782,I1307799,I1307816,I1307833,I1307864,I1307895,I1307921,I1307943,I1308015,I1308041,I1308049,I1308066,I1308092,I1308100,I1308117,I1308134,I1308151,I1308168,I1308199,I1308216,I1308233,I1308264,I1308281,I1308321,I1308329,I1308360,I1308377,I1308394,I1308411,I1308442,I1308473,I1308499,I1308521,I1308593,I1308619,I1308627,I1308644,I1308670,I1308678,I1308695,I1308712,I1308729,I1308746,I1308777,I1308794,I1308811,I1308842,I1308859,I1308899,I1308907,I1308938,I1308955,I1308972,I1308989,I1309020,I1309051,I1309077,I1309099,I1309171,I1386887,I1309197,I1309205,I1386878,I1309222,I1386863,I1309248,I1309256,I1309273,I1386866,I1309290,I1386875,I1309307,I1309324,I1386872,I1309355,I1386884,I1309372,I1309389,I1309420,I1386869,I1309437,I1309477,I1309485,I1309516,I1386890,I1309533,I1309550,I1309567,I1309598,I1309629,I1386881,I1309655,I1309677,I1309749,I1309775,I1309783,I1309800,I1309826,I1309834,I1309851,I1309868,I1309885,I1309902,I1309933,I1309950,I1309967,I1309998,I1310015,I1310055,I1310063,I1310094,I1310111,I1310128,I1310145,I1310176,I1310207,I1310233,I1310255,I1310327,I1310353,I1310361,I1310378,I1310404,I1310412,I1310429,I1310446,I1310463,I1310480,I1310511,I1310528,I1310545,I1310576,I1310593,I1310633,I1310641,I1310672,I1310689,I1310706,I1310723,I1310754,I1310785,I1310811,I1310833,I1310905,I1310931,I1310939,I1310956,I1310982,I1310990,I1311007,I1311024,I1311041,I1311058,I1311089,I1311106,I1311123,I1311154,I1311171,I1311211,I1311219,I1311250,I1311267,I1311284,I1311301,I1311332,I1311363,I1311389,I1311411,I1311483,I1311509,I1311517,I1311534,I1311560,I1311568,I1311585,I1311602,I1311619,I1311636,I1311667,I1311684,I1311701,I1311732,I1311749,I1311789,I1311797,I1311828,I1311845,I1311862,I1311879,I1311910,I1311941,I1311967,I1311989,I1312061,I1312087,I1312095,I1312112,I1312138,I1312146,I1312163,I1312180,I1312197,I1312214,I1312053,I1312245,I1312262,I1312279,I1312032,I1312310,I1312327,I1312038,I1312367,I1312375,I1312047,I1312406,I1312423,I1312440,I1312457,I1312050,I1312488,I1312029,I1312519,I1312545,I1312044,I1312567,I1312041,I1312035,I1312639,I1312665,I1312673,I1312690,I1312716,I1312724,I1312741,I1312758,I1312775,I1312792,I1312823,I1312840,I1312857,I1312888,I1312905,I1312945,I1312953,I1312984,I1313001,I1313018,I1313035,I1313066,I1313097,I1313123,I1313145,I1313217,I1313243,I1313251,I1313268,I1313294,I1313302,I1313319,I1313336,I1313353,I1313370,I1313401,I1313418,I1313435,I1313466,I1313483,I1313523,I1313531,I1313562,I1313579,I1313596,I1313613,I1313644,I1313675,I1313701,I1313723,I1313795,I1313821,I1313829,I1313846,I1313872,I1313880,I1313897,I1313914,I1313931,I1313948,I1313979,I1313996,I1314013,I1314044,I1314061,I1314101,I1314109,I1314140,I1314157,I1314174,I1314191,I1314222,I1314253,I1314279,I1314301,I1314373,I1354162,I1314399,I1314407,I1354153,I1314424,I1354138,I1314450,I1314458,I1314475,I1354141,I1314492,I1354150,I1314509,I1314526,I1354147,I1314557,I1354159,I1314574,I1314591,I1314622,I1354144,I1314639,I1314679,I1314687,I1314718,I1354165,I1314735,I1314752,I1314769,I1314800,I1314831,I1354156,I1314857,I1314879,I1314951,I1314977,I1314985,I1315002,I1315028,I1315036,I1315053,I1315070,I1315087,I1315104,I1315135,I1315152,I1315169,I1315200,I1315217,I1315257,I1315265,I1315296,I1315313,I1315330,I1315347,I1315378,I1315409,I1315435,I1315457,I1315529,I1315555,I1315563,I1315580,I1315606,I1315614,I1315631,I1315648,I1315665,I1315682,I1315713,I1315730,I1315747,I1315778,I1315795,I1315835,I1315843,I1315874,I1315891,I1315908,I1315925,I1315956,I1315987,I1316013,I1316035,I1316107,I1316133,I1316141,I1316158,I1316184,I1316192,I1316209,I1316226,I1316243,I1316260,I1316291,I1316308,I1316325,I1316356,I1316373,I1316413,I1316421,I1316452,I1316469,I1316486,I1316503,I1316534,I1316565,I1316591,I1316613,I1316685,I1316711,I1316719,I1316736,I1316762,I1316770,I1316787,I1316804,I1316821,I1316838,I1316869,I1316886,I1316903,I1316934,I1316951,I1316991,I1316999,I1317030,I1317047,I1317064,I1317081,I1317112,I1317143,I1317169,I1317191,I1317263,I1317289,I1317297,I1317314,I1317340,I1317348,I1317365,I1317382,I1317399,I1317416,I1317447,I1317464,I1317481,I1317512,I1317529,I1317569,I1317577,I1317608,I1317625,I1317642,I1317659,I1317690,I1317721,I1317747,I1317769,I1317841,I1317867,I1317875,I1317892,I1317918,I1317926,I1317943,I1317960,I1317977,I1317994,I1318025,I1318042,I1318059,I1318090,I1318107,I1318147,I1318155,I1318186,I1318203,I1318220,I1318237,I1318268,I1318299,I1318325,I1318347,I1318419,I1318445,I1318453,I1318470,I1318496,I1318504,I1318521,I1318538,I1318555,I1318572,I1318603,I1318620,I1318637,I1318668,I1318685,I1318725,I1318733,I1318764,I1318781,I1318798,I1318815,I1318846,I1318877,I1318903,I1318925,I1318997,I1338692,I1319023,I1319031,I1338683,I1319048,I1338668,I1319074,I1319082,I1319099,I1338671,I1319116,I1338680,I1319133,I1319150,I1338677,I1319181,I1338689,I1319198,I1319215,I1319246,I1338674,I1319263,I1319303,I1319311,I1319342,I1338695,I1319359,I1319376,I1319393,I1319424,I1319455,I1338686,I1319481,I1319503,I1319575,I1319601,I1319609,I1319626,I1319652,I1319660,I1319677,I1319694,I1319711,I1319728,I1319759,I1319776,I1319793,I1319824,I1319841,I1319881,I1319889,I1319920,I1319937,I1319954,I1319971,I1320002,I1320033,I1320059,I1320081,I1320153,I1320179,I1320187,I1320204,I1320230,I1320238,I1320255,I1320272,I1320289,I1320306,I1320337,I1320354,I1320371,I1320402,I1320419,I1320459,I1320467,I1320498,I1320515,I1320532,I1320549,I1320580,I1320611,I1320637,I1320659,I1320731,I1320757,I1320765,I1320782,I1320808,I1320816,I1320833,I1320850,I1320867,I1320884,I1320723,I1320915,I1320932,I1320949,I1320702,I1320980,I1320997,I1320708,I1321037,I1321045,I1320717,I1321076,I1321093,I1321110,I1321127,I1320720,I1321158,I1320699,I1321189,I1321215,I1320714,I1321237,I1320711,I1320705,I1321309,I1321335,I1321343,I1321360,I1321386,I1321394,I1321411,I1321428,I1321445,I1321462,I1321493,I1321510,I1321527,I1321558,I1321575,I1321615,I1321623,I1321654,I1321671,I1321688,I1321705,I1321736,I1321767,I1321793,I1321815,I1321887,I1321913,I1321921,I1321938,I1321964,I1321972,I1321989,I1322006,I1322023,I1322040,I1322071,I1322088,I1322105,I1322136,I1322153,I1322193,I1322201,I1322232,I1322249,I1322266,I1322283,I1322314,I1322345,I1322371,I1322393,I1322465,I1322491,I1322499,I1322516,I1322542,I1322550,I1322567,I1322584,I1322601,I1322618,I1322457,I1322649,I1322666,I1322683,I1322436,I1322714,I1322731,I1322442,I1322771,I1322779,I1322451,I1322810,I1322827,I1322844,I1322861,I1322454,I1322892,I1322433,I1322923,I1322949,I1322448,I1322971,I1322445,I1322439,I1323043,I1323069,I1323077,I1323094,I1323120,I1323128,I1323145,I1323162,I1323179,I1323196,I1323227,I1323244,I1323261,I1323292,I1323309,I1323349,I1323357,I1323388,I1323405,I1323422,I1323439,I1323470,I1323501,I1323527,I1323549,I1323621,I1323647,I1323655,I1323672,I1323698,I1323706,I1323723,I1323740,I1323757,I1323774,I1323805,I1323822,I1323839,I1323870,I1323887,I1323927,I1323935,I1323966,I1323983,I1324000,I1324017,I1324048,I1324079,I1324105,I1324127,I1324202,I1324228,I1324236,I1324253,I1324279,I1324287,I1324304,I1324321,I1324352,I1324383,I1324400,I1324417,I1324434,I1324451,I1324482,I1324541,I1324558,I1324584,I1324606,I1324632,I1324640,I1324657,I1324688,I1324763,I1324789,I1324797,I1324814,I1324840,I1324848,I1324865,I1324882,I1324913,I1324944,I1324961,I1324978,I1324995,I1325012,I1325043,I1325102,I1325119,I1325145,I1325167,I1325193,I1325201,I1325218,I1325249,I1325324,I1325350,I1325358,I1325375,I1325401,I1325409,I1325426,I1325443,I1325310,I1325474,I1325313,I1325505,I1325522,I1325539,I1325556,I1325573,I1325298,I1325604,I1325301,I1325295,I1325292,I1325663,I1325680,I1325706,I1325316,I1325728,I1325754,I1325762,I1325779,I1325307,I1325810,I1325289,I1325304,I1325885,I1325911,I1325919,I1325936,I1325962,I1325970,I1325987,I1326004,I1326035,I1326066,I1326083,I1326100,I1326117,I1326134,I1326165,I1326224,I1326241,I1326267,I1326289,I1326315,I1326323,I1326340,I1326371,I1326446,I1326472,I1326480,I1326497,I1326523,I1326531,I1326548,I1326565,I1326596,I1326627,I1326644,I1326661,I1326678,I1326695,I1326726,I1326785,I1326802,I1326828,I1326850,I1326876,I1326884,I1326901,I1326932,I1327007,I1327033,I1327041,I1327058,I1327084,I1327092,I1327109,I1327126,I1327157,I1327188,I1327205,I1327222,I1327239,I1327256,I1327287,I1327346,I1327363,I1327389,I1327411,I1327437,I1327445,I1327462,I1327493,I1327568,I1327594,I1327602,I1327619,I1327645,I1327653,I1327670,I1327687,I1327718,I1327749,I1327766,I1327783,I1327800,I1327817,I1327848,I1327907,I1327924,I1327950,I1327972,I1327998,I1328006,I1328023,I1328054,I1328129,I1328155,I1328163,I1328180,I1328206,I1328214,I1328231,I1328248,I1328279,I1328310,I1328327,I1328344,I1328361,I1328378,I1328409,I1328468,I1328485,I1328511,I1328533,I1328559,I1328567,I1328584,I1328615,I1328690,I1328716,I1328724,I1328741,I1328767,I1328775,I1328792,I1328809,I1328840,I1328871,I1328888,I1328905,I1328922,I1328939,I1328970,I1329029,I1329046,I1329072,I1329094,I1329120,I1329128,I1329145,I1329176,I1329251,I1329277,I1329285,I1329302,I1329328,I1329336,I1329353,I1329370,I1329401,I1329432,I1329449,I1329466,I1329483,I1329500,I1329531,I1329590,I1329607,I1329633,I1329655,I1329681,I1329689,I1329706,I1329737,I1329812,I1329838,I1329846,I1329863,I1329889,I1329897,I1329914,I1329931,I1329962,I1329993,I1330010,I1330027,I1330044,I1330061,I1330092,I1330151,I1330168,I1330194,I1330216,I1330242,I1330250,I1330267,I1330298,I1330373,I1330399,I1330416,I1330424,I1330469,I1330486,I1330503,I1330520,I1330537,I1330554,I1330571,I1330602,I1330619,I1330664,I1330681,I1330698,I1330729,I1330755,I1330763,I1330794,I1330811,I1330828,I1330854,I1330862,I1330879,I1330968,I1330994,I1331011,I1331019,I1331064,I1331081,I1331098,I1331115,I1331132,I1331149,I1331166,I1331197,I1331214,I1331259,I1331276,I1331293,I1331324,I1331350,I1331358,I1331389,I1331406,I1331423,I1331449,I1331457,I1331474,I1331563,I1331589,I1331606,I1331614,I1331659,I1331676,I1331693,I1331710,I1331727,I1331744,I1331761,I1331792,I1331809,I1331854,I1331871,I1331888,I1331919,I1331945,I1331953,I1331984,I1332001,I1332018,I1332044,I1332052,I1332069,I1332158,I1332184,I1332201,I1332209,I1332254,I1332271,I1332288,I1332305,I1332322,I1332339,I1332356,I1332387,I1332404,I1332449,I1332466,I1332483,I1332514,I1332540,I1332548,I1332579,I1332596,I1332613,I1332639,I1332647,I1332664,I1332753,I1332779,I1332796,I1332804,I1332849,I1332866,I1332883,I1332900,I1332917,I1332934,I1332951,I1332982,I1332999,I1333044,I1333061,I1333078,I1333109,I1333135,I1333143,I1333174,I1333191,I1333208,I1333234,I1333242,I1333259,I1333348,I1333374,I1333391,I1333399,I1333444,I1333461,I1333478,I1333495,I1333512,I1333529,I1333546,I1333577,I1333594,I1333639,I1333656,I1333673,I1333704,I1333730,I1333738,I1333769,I1333786,I1333803,I1333829,I1333837,I1333854,I1333943,I1333969,I1333986,I1333994,I1334039,I1334056,I1334073,I1334090,I1334107,I1334124,I1334141,I1334172,I1334189,I1334234,I1334251,I1334268,I1334299,I1334325,I1334333,I1334364,I1334381,I1334398,I1334424,I1334432,I1334449,I1334538,I1334564,I1334581,I1334589,I1334634,I1334651,I1334668,I1334685,I1334702,I1334719,I1334736,I1334767,I1334784,I1334829,I1334846,I1334863,I1334894,I1334920,I1334928,I1334959,I1334976,I1334993,I1335019,I1335027,I1335044,I1335133,I1335159,I1335176,I1335184,I1335229,I1335246,I1335263,I1335280,I1335297,I1335314,I1335331,I1335362,I1335379,I1335424,I1335441,I1335458,I1335489,I1335515,I1335523,I1335554,I1335571,I1335588,I1335614,I1335622,I1335639,I1335728,I1335754,I1335771,I1335779,I1335824,I1335841,I1335858,I1335875,I1335892,I1335909,I1335926,I1335957,I1335974,I1336019,I1336036,I1336053,I1336084,I1336110,I1336118,I1336149,I1336166,I1336183,I1336209,I1336217,I1336234,I1336323,I1336349,I1336366,I1336374,I1336419,I1336436,I1336453,I1336470,I1336487,I1336504,I1336521,I1336552,I1336569,I1336614,I1336631,I1336648,I1336679,I1336705,I1336713,I1336744,I1336761,I1336778,I1336804,I1336812,I1336829,I1336918,I1336944,I1336961,I1336969,I1337014,I1337031,I1337048,I1337065,I1337082,I1337099,I1337116,I1337147,I1337164,I1337209,I1337226,I1337243,I1337274,I1337300,I1337308,I1337339,I1337356,I1337373,I1337399,I1337407,I1337424,I1337513,I1337539,I1337556,I1337564,I1337609,I1337626,I1337643,I1337660,I1337677,I1337694,I1337711,I1337742,I1337759,I1337804,I1337821,I1337838,I1337869,I1337895,I1337903,I1337934,I1337951,I1337968,I1337994,I1338002,I1338019,I1338108,I1338134,I1338151,I1338159,I1338204,I1338221,I1338238,I1338255,I1338272,I1338289,I1338306,I1338337,I1338354,I1338399,I1338416,I1338433,I1338464,I1338490,I1338498,I1338529,I1338546,I1338563,I1338589,I1338597,I1338614,I1338703,I1338729,I1338746,I1338754,I1338799,I1338816,I1338833,I1338850,I1338867,I1338884,I1338901,I1338932,I1338949,I1338994,I1339011,I1339028,I1339059,I1339085,I1339093,I1339124,I1339141,I1339158,I1339184,I1339192,I1339209,I1339298,I1339324,I1339341,I1339349,I1339394,I1339411,I1339428,I1339445,I1339462,I1339479,I1339496,I1339527,I1339544,I1339589,I1339606,I1339623,I1339654,I1339680,I1339688,I1339719,I1339736,I1339753,I1339779,I1339787,I1339804,I1339893,I1339919,I1339936,I1339944,I1339989,I1340006,I1340023,I1340040,I1340057,I1340074,I1340091,I1340122,I1340139,I1340184,I1340201,I1340218,I1340249,I1340275,I1340283,I1340314,I1340331,I1340348,I1340374,I1340382,I1340399,I1340488,I1340514,I1340531,I1340539,I1340584,I1340601,I1340618,I1340635,I1340652,I1340669,I1340686,I1340717,I1340734,I1340779,I1340796,I1340813,I1340844,I1340870,I1340878,I1340909,I1340926,I1340943,I1340969,I1340977,I1340994,I1341083,I1341109,I1341126,I1341134,I1341179,I1341196,I1341213,I1341230,I1341247,I1341264,I1341281,I1341312,I1341329,I1341374,I1341391,I1341408,I1341439,I1341465,I1341473,I1341504,I1341521,I1341538,I1341564,I1341572,I1341589,I1341678,I1341704,I1341721,I1341729,I1341774,I1341791,I1341808,I1341825,I1341842,I1341859,I1341876,I1341907,I1341924,I1341969,I1341986,I1342003,I1342034,I1342060,I1342068,I1342099,I1342116,I1342133,I1342159,I1342167,I1342184,I1342273,I1342299,I1342316,I1342324,I1342369,I1342386,I1342403,I1342420,I1342437,I1342454,I1342471,I1342502,I1342519,I1342564,I1342581,I1342598,I1342629,I1342655,I1342663,I1342694,I1342711,I1342728,I1342754,I1342762,I1342779,I1342868,I1342894,I1342911,I1342919,I1342964,I1342981,I1342998,I1343015,I1343032,I1343049,I1343066,I1343097,I1343114,I1343159,I1343176,I1343193,I1343224,I1343250,I1343258,I1343289,I1343306,I1343323,I1343349,I1343357,I1343374,I1343463,I1343489,I1343506,I1343514,I1343559,I1343576,I1343593,I1343610,I1343627,I1343644,I1343661,I1343692,I1343709,I1343754,I1343771,I1343788,I1343819,I1343845,I1343853,I1343884,I1343901,I1343918,I1343944,I1343952,I1343969,I1344058,I1344084,I1344101,I1344109,I1344154,I1344171,I1344188,I1344205,I1344222,I1344239,I1344256,I1344287,I1344304,I1344349,I1344366,I1344383,I1344414,I1344440,I1344448,I1344479,I1344496,I1344513,I1344539,I1344547,I1344564,I1344653,I1344679,I1344696,I1344704,I1344749,I1344766,I1344783,I1344800,I1344817,I1344834,I1344851,I1344882,I1344899,I1344944,I1344961,I1344978,I1345009,I1345035,I1345043,I1345074,I1345091,I1345108,I1345134,I1345142,I1345159,I1345248,I1345274,I1345291,I1345299,I1345344,I1345361,I1345378,I1345395,I1345412,I1345429,I1345446,I1345477,I1345494,I1345539,I1345556,I1345573,I1345604,I1345630,I1345638,I1345669,I1345686,I1345703,I1345729,I1345737,I1345754,I1345843,I1345869,I1345886,I1345894,I1345939,I1345956,I1345973,I1345990,I1346007,I1346024,I1346041,I1346072,I1346089,I1346134,I1346151,I1346168,I1346199,I1346225,I1346233,I1346264,I1346281,I1346298,I1346324,I1346332,I1346349,I1346438,I1346464,I1346481,I1346489,I1346534,I1346551,I1346568,I1346585,I1346602,I1346619,I1346636,I1346667,I1346684,I1346729,I1346746,I1346763,I1346794,I1346820,I1346828,I1346859,I1346876,I1346893,I1346919,I1346927,I1346944,I1347033,I1347059,I1347076,I1347084,I1347129,I1347146,I1347163,I1347180,I1347197,I1347214,I1347231,I1347262,I1347279,I1347324,I1347341,I1347358,I1347389,I1347415,I1347423,I1347454,I1347471,I1347488,I1347514,I1347522,I1347539,I1347628,I1347654,I1347671,I1347679,I1347724,I1347741,I1347758,I1347775,I1347792,I1347809,I1347826,I1347857,I1347874,I1347919,I1347936,I1347953,I1347984,I1348010,I1348018,I1348049,I1348066,I1348083,I1348109,I1348117,I1348134,I1348223,I1348249,I1348266,I1348274,I1348319,I1348336,I1348353,I1348370,I1348387,I1348404,I1348421,I1348452,I1348469,I1348514,I1348531,I1348548,I1348579,I1348605,I1348613,I1348644,I1348661,I1348678,I1348704,I1348712,I1348729,I1348818,I1348844,I1348861,I1348869,I1348914,I1348931,I1348948,I1348965,I1348982,I1348999,I1349016,I1349047,I1349064,I1349109,I1349126,I1349143,I1349174,I1349200,I1349208,I1349239,I1349256,I1349273,I1349299,I1349307,I1349324,I1349413,I1349439,I1349456,I1349464,I1349509,I1349526,I1349543,I1349560,I1349577,I1349594,I1349611,I1349642,I1349659,I1349704,I1349721,I1349738,I1349769,I1349795,I1349803,I1349834,I1349851,I1349868,I1349894,I1349902,I1349919,I1350008,I1350034,I1350051,I1350059,I1350104,I1350121,I1350138,I1350155,I1350172,I1350189,I1350206,I1350237,I1350254,I1350299,I1350316,I1350333,I1350364,I1350390,I1350398,I1350429,I1350446,I1350463,I1350489,I1350497,I1350514,I1350603,I1350629,I1350646,I1350654,I1350699,I1350716,I1350733,I1350750,I1350767,I1350784,I1350801,I1350832,I1350849,I1350894,I1350911,I1350928,I1350959,I1350985,I1350993,I1351024,I1351041,I1351058,I1351084,I1351092,I1351109,I1351198,I1351224,I1351241,I1351249,I1351294,I1351311,I1351328,I1351345,I1351362,I1351379,I1351396,I1351427,I1351444,I1351489,I1351506,I1351523,I1351554,I1351580,I1351588,I1351619,I1351636,I1351653,I1351679,I1351687,I1351704,I1351793,I1351819,I1351836,I1351844,I1351889,I1351906,I1351923,I1351940,I1351957,I1351974,I1351991,I1352022,I1352039,I1352084,I1352101,I1352118,I1352149,I1352175,I1352183,I1352214,I1352231,I1352248,I1352274,I1352282,I1352299,I1352388,I1352414,I1352431,I1352439,I1352484,I1352501,I1352518,I1352535,I1352552,I1352569,I1352586,I1352617,I1352634,I1352679,I1352696,I1352713,I1352744,I1352770,I1352778,I1352809,I1352826,I1352843,I1352869,I1352877,I1352894,I1352983,I1353009,I1353026,I1353034,I1353079,I1353096,I1353113,I1353130,I1353147,I1353164,I1353181,I1353212,I1353229,I1353274,I1353291,I1353308,I1353339,I1353365,I1353373,I1353404,I1353421,I1353438,I1353464,I1353472,I1353489,I1353578,I1353604,I1353621,I1353629,I1353674,I1353691,I1353708,I1353725,I1353742,I1353759,I1353776,I1353807,I1353824,I1353869,I1353886,I1353903,I1353934,I1353960,I1353968,I1353999,I1354016,I1354033,I1354059,I1354067,I1354084,I1354173,I1354199,I1354216,I1354224,I1354269,I1354286,I1354303,I1354320,I1354337,I1354354,I1354371,I1354402,I1354419,I1354464,I1354481,I1354498,I1354529,I1354555,I1354563,I1354594,I1354611,I1354628,I1354654,I1354662,I1354679,I1354768,I1354794,I1354811,I1354819,I1354864,I1354881,I1354898,I1354915,I1354932,I1354949,I1354966,I1354997,I1355014,I1355059,I1355076,I1355093,I1355124,I1355150,I1355158,I1355189,I1355206,I1355223,I1355249,I1355257,I1355274,I1355363,I1355389,I1355406,I1355414,I1355459,I1355476,I1355493,I1355510,I1355527,I1355544,I1355561,I1355592,I1355609,I1355654,I1355671,I1355688,I1355719,I1355745,I1355753,I1355784,I1355801,I1355818,I1355844,I1355852,I1355869,I1355958,I1355984,I1356001,I1356009,I1356054,I1356071,I1356088,I1356105,I1356122,I1356139,I1356156,I1356187,I1356204,I1356249,I1356266,I1356283,I1356314,I1356340,I1356348,I1356379,I1356396,I1356413,I1356439,I1356447,I1356464,I1356553,I1356579,I1356596,I1356604,I1356649,I1356666,I1356683,I1356700,I1356717,I1356734,I1356751,I1356782,I1356799,I1356844,I1356861,I1356878,I1356909,I1356935,I1356943,I1356974,I1356991,I1357008,I1357034,I1357042,I1357059,I1357148,I1357174,I1357191,I1357199,I1357244,I1357261,I1357278,I1357295,I1357312,I1357329,I1357346,I1357377,I1357394,I1357439,I1357456,I1357473,I1357504,I1357530,I1357538,I1357569,I1357586,I1357603,I1357629,I1357637,I1357654,I1357743,I1357769,I1357786,I1357794,I1357839,I1357856,I1357873,I1357890,I1357907,I1357924,I1357941,I1357972,I1357989,I1358034,I1358051,I1358068,I1358099,I1358125,I1358133,I1358164,I1358181,I1358198,I1358224,I1358232,I1358249,I1358338,I1358364,I1358381,I1358389,I1358434,I1358451,I1358468,I1358485,I1358502,I1358519,I1358536,I1358567,I1358584,I1358629,I1358646,I1358663,I1358694,I1358720,I1358728,I1358759,I1358776,I1358793,I1358819,I1358827,I1358844,I1358933,I1358959,I1358976,I1358984,I1359029,I1359046,I1359063,I1359080,I1359097,I1359114,I1359131,I1359162,I1359179,I1359224,I1359241,I1359258,I1359289,I1359315,I1359323,I1359354,I1359371,I1359388,I1359414,I1359422,I1359439,I1359528,I1359554,I1359571,I1359579,I1359624,I1359641,I1359658,I1359675,I1359692,I1359709,I1359726,I1359757,I1359774,I1359819,I1359836,I1359853,I1359884,I1359910,I1359918,I1359949,I1359966,I1359983,I1360009,I1360017,I1360034,I1360123,I1360149,I1360166,I1360174,I1360219,I1360236,I1360253,I1360270,I1360287,I1360304,I1360321,I1360352,I1360369,I1360414,I1360431,I1360448,I1360479,I1360505,I1360513,I1360544,I1360561,I1360578,I1360604,I1360612,I1360629,I1360718,I1360744,I1360761,I1360769,I1360814,I1360831,I1360848,I1360865,I1360882,I1360899,I1360916,I1360947,I1360964,I1361009,I1361026,I1361043,I1361074,I1361100,I1361108,I1361139,I1361156,I1361173,I1361199,I1361207,I1361224,I1361313,I1361339,I1361356,I1361364,I1361409,I1361426,I1361443,I1361460,I1361477,I1361494,I1361511,I1361542,I1361559,I1361604,I1361621,I1361638,I1361669,I1361695,I1361703,I1361734,I1361751,I1361768,I1361794,I1361802,I1361819,I1361908,I1361934,I1361951,I1361959,I1362004,I1362021,I1362038,I1362055,I1362072,I1362089,I1362106,I1362137,I1362154,I1362199,I1362216,I1362233,I1362264,I1362290,I1362298,I1362329,I1362346,I1362363,I1362389,I1362397,I1362414,I1362503,I1362529,I1362546,I1362554,I1362599,I1362616,I1362633,I1362650,I1362667,I1362684,I1362701,I1362732,I1362749,I1362794,I1362811,I1362828,I1362859,I1362885,I1362893,I1362924,I1362941,I1362958,I1362984,I1362992,I1363009,I1363098,I1363124,I1363141,I1363149,I1363194,I1363211,I1363228,I1363245,I1363262,I1363279,I1363296,I1363327,I1363344,I1363389,I1363406,I1363423,I1363454,I1363480,I1363488,I1363519,I1363536,I1363553,I1363579,I1363587,I1363604,I1363693,I1363719,I1363736,I1363744,I1363789,I1363806,I1363823,I1363840,I1363857,I1363874,I1363891,I1363922,I1363939,I1363984,I1364001,I1364018,I1364049,I1364075,I1364083,I1364114,I1364131,I1364148,I1364174,I1364182,I1364199,I1364288,I1364314,I1364331,I1364339,I1364384,I1364401,I1364418,I1364435,I1364452,I1364469,I1364486,I1364517,I1364534,I1364579,I1364596,I1364613,I1364644,I1364670,I1364678,I1364709,I1364726,I1364743,I1364769,I1364777,I1364794,I1364883,I1364909,I1364926,I1364934,I1364979,I1364996,I1365013,I1365030,I1365047,I1365064,I1365081,I1365112,I1365129,I1365174,I1365191,I1365208,I1365239,I1365265,I1365273,I1365304,I1365321,I1365338,I1365364,I1365372,I1365389,I1365478,I1365504,I1365521,I1365529,I1365574,I1365591,I1365608,I1365625,I1365642,I1365659,I1365676,I1365707,I1365724,I1365769,I1365786,I1365803,I1365834,I1365860,I1365868,I1365899,I1365916,I1365933,I1365959,I1365967,I1365984,I1366073,I1366099,I1366116,I1366124,I1366169,I1366186,I1366203,I1366220,I1366237,I1366254,I1366271,I1366302,I1366319,I1366364,I1366381,I1366398,I1366429,I1366455,I1366463,I1366494,I1366511,I1366528,I1366554,I1366562,I1366579,I1366668,I1366694,I1366711,I1366719,I1366764,I1366781,I1366798,I1366815,I1366832,I1366849,I1366866,I1366897,I1366914,I1366959,I1366976,I1366993,I1367024,I1367050,I1367058,I1367089,I1367106,I1367123,I1367149,I1367157,I1367174,I1367263,I1367289,I1367306,I1367314,I1367359,I1367376,I1367393,I1367410,I1367427,I1367444,I1367461,I1367492,I1367509,I1367554,I1367571,I1367588,I1367619,I1367645,I1367653,I1367684,I1367701,I1367718,I1367744,I1367752,I1367769,I1367858,I1367884,I1367901,I1367909,I1367954,I1367971,I1367988,I1368005,I1368022,I1368039,I1368056,I1368087,I1368104,I1368149,I1368166,I1368183,I1368214,I1368240,I1368248,I1368279,I1368296,I1368313,I1368339,I1368347,I1368364,I1368453,I1368479,I1368496,I1368504,I1368549,I1368566,I1368583,I1368600,I1368617,I1368634,I1368651,I1368682,I1368699,I1368744,I1368761,I1368778,I1368809,I1368835,I1368843,I1368874,I1368891,I1368908,I1368934,I1368942,I1368959,I1369048,I1369074,I1369091,I1369099,I1369144,I1369161,I1369178,I1369195,I1369212,I1369229,I1369246,I1369277,I1369294,I1369339,I1369356,I1369373,I1369404,I1369430,I1369438,I1369469,I1369486,I1369503,I1369529,I1369537,I1369554,I1369643,I1369669,I1369686,I1369694,I1369739,I1369756,I1369773,I1369790,I1369807,I1369824,I1369841,I1369872,I1369889,I1369934,I1369951,I1369968,I1369999,I1370025,I1370033,I1370064,I1370081,I1370098,I1370124,I1370132,I1370149,I1370238,I1370264,I1370281,I1370289,I1370334,I1370351,I1370368,I1370385,I1370402,I1370419,I1370436,I1370467,I1370484,I1370529,I1370546,I1370563,I1370594,I1370620,I1370628,I1370659,I1370676,I1370693,I1370719,I1370727,I1370744,I1370833,I1370859,I1370876,I1370884,I1370929,I1370946,I1370963,I1370980,I1370997,I1371014,I1371031,I1371062,I1371079,I1371124,I1371141,I1371158,I1371189,I1371215,I1371223,I1371254,I1371271,I1371288,I1371314,I1371322,I1371339,I1371428,I1371454,I1371471,I1371479,I1371524,I1371541,I1371558,I1371575,I1371592,I1371609,I1371626,I1371657,I1371674,I1371719,I1371736,I1371753,I1371784,I1371810,I1371818,I1371849,I1371866,I1371883,I1371909,I1371917,I1371934,I1372023,I1372049,I1372066,I1372074,I1372119,I1372136,I1372153,I1372170,I1372187,I1372204,I1372221,I1372252,I1372269,I1372314,I1372331,I1372348,I1372379,I1372405,I1372413,I1372444,I1372461,I1372478,I1372504,I1372512,I1372529,I1372618,I1372644,I1372661,I1372669,I1372714,I1372731,I1372748,I1372765,I1372782,I1372799,I1372816,I1372847,I1372864,I1372909,I1372926,I1372943,I1372974,I1373000,I1373008,I1373039,I1373056,I1373073,I1373099,I1373107,I1373124,I1373213,I1373239,I1373256,I1373264,I1373309,I1373326,I1373343,I1373360,I1373377,I1373394,I1373411,I1373442,I1373459,I1373504,I1373521,I1373538,I1373569,I1373595,I1373603,I1373634,I1373651,I1373668,I1373694,I1373702,I1373719,I1373808,I1373834,I1373851,I1373859,I1373904,I1373921,I1373938,I1373955,I1373972,I1373989,I1374006,I1374037,I1374054,I1374099,I1374116,I1374133,I1374164,I1374190,I1374198,I1374229,I1374246,I1374263,I1374289,I1374297,I1374314,I1374403,I1374429,I1374446,I1374454,I1374499,I1374516,I1374533,I1374550,I1374567,I1374584,I1374601,I1374632,I1374649,I1374694,I1374711,I1374728,I1374759,I1374785,I1374793,I1374824,I1374841,I1374858,I1374884,I1374892,I1374909,I1374998,I1375024,I1375041,I1375049,I1375094,I1375111,I1375128,I1375145,I1375162,I1375179,I1375196,I1375227,I1375244,I1375289,I1375306,I1375323,I1375354,I1375380,I1375388,I1375419,I1375436,I1375453,I1375479,I1375487,I1375504,I1375593,I1375619,I1375636,I1375644,I1375689,I1375706,I1375723,I1375740,I1375757,I1375774,I1375791,I1375822,I1375839,I1375884,I1375901,I1375918,I1375949,I1375975,I1375983,I1376014,I1376031,I1376048,I1376074,I1376082,I1376099,I1376188,I1376214,I1376231,I1376239,I1376284,I1376301,I1376318,I1376335,I1376352,I1376369,I1376386,I1376417,I1376434,I1376479,I1376496,I1376513,I1376544,I1376570,I1376578,I1376609,I1376626,I1376643,I1376669,I1376677,I1376694,I1376783,I1376809,I1376826,I1376834,I1376879,I1376896,I1376913,I1376930,I1376947,I1376964,I1376981,I1377012,I1377029,I1377074,I1377091,I1377108,I1377139,I1377165,I1377173,I1377204,I1377221,I1377238,I1377264,I1377272,I1377289,I1377378,I1377404,I1377421,I1377429,I1377474,I1377491,I1377508,I1377525,I1377542,I1377559,I1377576,I1377607,I1377624,I1377669,I1377686,I1377703,I1377734,I1377760,I1377768,I1377799,I1377816,I1377833,I1377859,I1377867,I1377884,I1377973,I1377999,I1378016,I1378024,I1378069,I1378086,I1378103,I1378120,I1378137,I1378154,I1378171,I1378202,I1378219,I1378264,I1378281,I1378298,I1378329,I1378355,I1378363,I1378394,I1378411,I1378428,I1378454,I1378462,I1378479,I1378568,I1378594,I1378611,I1378619,I1378664,I1378681,I1378698,I1378715,I1378732,I1378749,I1378766,I1378797,I1378814,I1378859,I1378876,I1378893,I1378924,I1378950,I1378958,I1378989,I1379006,I1379023,I1379049,I1379057,I1379074,I1379163,I1379189,I1379206,I1379214,I1379259,I1379276,I1379293,I1379310,I1379327,I1379344,I1379361,I1379392,I1379409,I1379454,I1379471,I1379488,I1379519,I1379545,I1379553,I1379584,I1379601,I1379618,I1379644,I1379652,I1379669,I1379758,I1379784,I1379801,I1379809,I1379854,I1379871,I1379888,I1379905,I1379922,I1379939,I1379956,I1379987,I1380004,I1380049,I1380066,I1380083,I1380114,I1380140,I1380148,I1380179,I1380196,I1380213,I1380239,I1380247,I1380264,I1380353,I1380379,I1380396,I1380404,I1380449,I1380466,I1380483,I1380500,I1380517,I1380534,I1380551,I1380582,I1380599,I1380644,I1380661,I1380678,I1380709,I1380735,I1380743,I1380774,I1380791,I1380808,I1380834,I1380842,I1380859,I1380948,I1380974,I1380991,I1380999,I1381044,I1381061,I1381078,I1381095,I1381112,I1381129,I1381146,I1381177,I1381194,I1381239,I1381256,I1381273,I1381304,I1381330,I1381338,I1381369,I1381386,I1381403,I1381429,I1381437,I1381454,I1381543,I1381569,I1381586,I1381594,I1381639,I1381656,I1381673,I1381690,I1381707,I1381724,I1381741,I1381772,I1381789,I1381834,I1381851,I1381868,I1381899,I1381925,I1381933,I1381964,I1381981,I1381998,I1382024,I1382032,I1382049,I1382138,I1382164,I1382181,I1382189,I1382234,I1382251,I1382268,I1382285,I1382302,I1382319,I1382336,I1382367,I1382384,I1382429,I1382446,I1382463,I1382494,I1382520,I1382528,I1382559,I1382576,I1382593,I1382619,I1382627,I1382644,I1382733,I1382759,I1382776,I1382784,I1382829,I1382846,I1382863,I1382880,I1382897,I1382914,I1382931,I1382962,I1382979,I1383024,I1383041,I1383058,I1383089,I1383115,I1383123,I1383154,I1383171,I1383188,I1383214,I1383222,I1383239,I1383328,I1383354,I1383371,I1383379,I1383424,I1383441,I1383458,I1383475,I1383492,I1383509,I1383526,I1383557,I1383574,I1383619,I1383636,I1383653,I1383684,I1383710,I1383718,I1383749,I1383766,I1383783,I1383809,I1383817,I1383834,I1383923,I1383949,I1383966,I1383974,I1384019,I1384036,I1384053,I1384070,I1384087,I1384104,I1384121,I1384152,I1384169,I1384214,I1384231,I1384248,I1384279,I1384305,I1384313,I1384344,I1384361,I1384378,I1384404,I1384412,I1384429,I1384518,I1384544,I1384561,I1384569,I1384614,I1384631,I1384648,I1384665,I1384682,I1384699,I1384716,I1384747,I1384764,I1384809,I1384826,I1384843,I1384874,I1384900,I1384908,I1384939,I1384956,I1384973,I1384999,I1385007,I1385024,I1385113,I1385139,I1385156,I1385164,I1385209,I1385226,I1385243,I1385260,I1385277,I1385294,I1385311,I1385342,I1385359,I1385404,I1385421,I1385438,I1385469,I1385495,I1385503,I1385534,I1385551,I1385568,I1385594,I1385602,I1385619,I1385708,I1385734,I1385751,I1385759,I1385804,I1385821,I1385838,I1385855,I1385872,I1385889,I1385906,I1385937,I1385954,I1385999,I1386016,I1386033,I1386064,I1386090,I1386098,I1386129,I1386146,I1386163,I1386189,I1386197,I1386214,I1386303,I1386329,I1386346,I1386354,I1386399,I1386416,I1386433,I1386450,I1386467,I1386484,I1386501,I1386532,I1386549,I1386594,I1386611,I1386628,I1386659,I1386685,I1386693,I1386724,I1386741,I1386758,I1386784,I1386792,I1386809,I1386898,I1386924,I1386941,I1386949,I1386994,I1387011,I1387028,I1387045,I1387062,I1387079,I1387096,I1387127,I1387144,I1387189,I1387206,I1387223,I1387254,I1387280,I1387288,I1387319,I1387336,I1387353,I1387379,I1387387,I1387404,I1387493,I1387519,I1387536,I1387544,I1387589,I1387606,I1387623,I1387640,I1387657,I1387674,I1387691,I1387722,I1387739,I1387784,I1387801,I1387818,I1387849,I1387875,I1387883,I1387914,I1387931,I1387948,I1387974,I1387982,I1387999,I1388088,I1388114,I1388131,I1388139,I1388184,I1388201,I1388218,I1388235,I1388252,I1388269,I1388286,I1388317,I1388334,I1388379,I1388396,I1388413,I1388444,I1388470,I1388478,I1388509,I1388526,I1388543,I1388569,I1388577,I1388594,I1388683,I1388709,I1388726,I1388734,I1388779,I1388796,I1388813,I1388830,I1388847,I1388864,I1388881,I1388912,I1388929,I1388974,I1388991,I1389008,I1389039,I1389065,I1389073,I1389104,I1389121,I1389138,I1389164,I1389172,I1389189,I1389278,I1389304,I1389321,I1389329,I1389374,I1389391,I1389408,I1389425,I1389442,I1389459,I1389476,I1389507,I1389524,I1389569,I1389586,I1389603,I1389634,I1389660,I1389668,I1389699,I1389716,I1389733,I1389759,I1389767,I1389784,I1389873,I1389899,I1389916,I1389924,I1389969,I1389986,I1390003,I1390020,I1390037,I1390054,I1390071,I1390102,I1390119,I1390164,I1390181,I1390198,I1390229,I1390255,I1390263,I1390294,I1390311,I1390328,I1390354,I1390362,I1390379,I1390468,I1390494,I1390511,I1390519,I1390564,I1390581,I1390598,I1390615,I1390632,I1390649,I1390666,I1390697,I1390714,I1390759,I1390776,I1390793,I1390824,I1390850,I1390858,I1390889,I1390906,I1390923,I1390949,I1390957,I1390974,I1391063,I1391089,I1391106,I1391114,I1391159,I1391176,I1391193,I1391210,I1391227,I1391244,I1391261,I1391292,I1391309,I1391354,I1391371,I1391388,I1391419,I1391445,I1391453,I1391484,I1391501,I1391518,I1391544,I1391552,I1391569,I1391658,I1391684,I1391701,I1391709,I1391754,I1391771,I1391788,I1391805,I1391822,I1391839,I1391856,I1391887,I1391904,I1391949,I1391966,I1391983,I1392014,I1392040,I1392048,I1392079,I1392096,I1392113,I1392139,I1392147,I1392164,I1392253,I1392279,I1392296,I1392304,I1392349,I1392366,I1392383,I1392400,I1392417,I1392434,I1392451,I1392482,I1392499,I1392544,I1392561,I1392578,I1392609,I1392635,I1392643,I1392674,I1392691,I1392708,I1392734,I1392742,I1392759,I1392848,I1392874,I1392891,I1392899,I1392944,I1392961,I1392978,I1392995,I1393012,I1393029,I1393046,I1393077,I1393094,I1393139,I1393156,I1393173,I1393204,I1393230,I1393238,I1393269,I1393286,I1393303,I1393329,I1393337,I1393354,I1393443,I1393469,I1393486,I1393494,I1393539,I1393556,I1393573,I1393590,I1393607,I1393624,I1393641,I1393672,I1393689,I1393734,I1393751,I1393768,I1393799,I1393825,I1393833,I1393864,I1393881,I1393898,I1393924,I1393932,I1393949,I1394038,I1394064,I1394081,I1394089,I1394134,I1394151,I1394168,I1394185,I1394202,I1394219,I1394236,I1394267,I1394284,I1394329,I1394346,I1394363,I1394394,I1394420,I1394428,I1394459,I1394476,I1394493,I1394519,I1394527,I1394544,I1394633,I1394659,I1394676,I1394684,I1394729,I1394746,I1394763,I1394780,I1394797,I1394814,I1394831,I1394862,I1394879,I1394924,I1394941,I1394958,I1394989,I1395015,I1395023,I1395054,I1395071,I1395088,I1395114,I1395122,I1395139,I1395228,I1395254,I1395271,I1395279,I1395324,I1395341,I1395358,I1395375,I1395392,I1395409,I1395426,I1395457,I1395474,I1395519,I1395536,I1395553,I1395584,I1395610,I1395618,I1395649,I1395666,I1395683,I1395709,I1395717,I1395734,I1395823,I1395849,I1395866,I1395874,I1395919,I1395936,I1395953,I1395970,I1395987,I1396004,I1396021,I1396052,I1396069,I1396114,I1396131,I1396148,I1396179,I1396205,I1396213,I1396244,I1396261,I1396278,I1396304,I1396312,I1396329,I1396418,I1396444,I1396461,I1396469,I1396514,I1396531,I1396548,I1396565,I1396582,I1396599,I1396616,I1396647,I1396664,I1396709,I1396726,I1396743,I1396774,I1396800,I1396808,I1396839,I1396856,I1396873,I1396899,I1396907,I1396924,I1397013,I1397039,I1397056,I1397064,I1397109,I1397126,I1397143,I1397160,I1397177,I1397194,I1397211,I1397242,I1397259,I1397304,I1397321,I1397338,I1397369,I1397395,I1397403,I1397434,I1397451,I1397468,I1397494,I1397502,I1397519,I1397608,I1397634,I1397651,I1397659,I1397704,I1397721,I1397738,I1397755,I1397772,I1397789,I1397806,I1397837,I1397854,I1397899,I1397916,I1397933,I1397964,I1397990,I1397998,I1398029,I1398046,I1398063,I1398089,I1398097,I1398114,I1398203,I1398229,I1398246,I1398254,I1398299,I1398316,I1398333,I1398350,I1398367,I1398384,I1398401,I1398432,I1398449,I1398494,I1398511,I1398528,I1398559,I1398585,I1398593,I1398624,I1398641,I1398658,I1398684,I1398692,I1398709,I1398798,I1398824,I1398841,I1398849,I1398894,I1398911,I1398928,I1398945,I1398962,I1398979,I1398996,I1399027,I1399044,I1399089,I1399106,I1399123,I1399154,I1399180,I1399188,I1399219,I1399236,I1399253,I1399279,I1399287,I1399304,I1399393,I1399419,I1399436,I1399444,I1399489,I1399506,I1399523,I1399540,I1399557,I1399574,I1399591,I1399622,I1399639,I1399684,I1399701,I1399718,I1399749,I1399775,I1399783,I1399814,I1399831,I1399848,I1399874,I1399882,I1399899,I1399988,I1400014,I1400031,I1400039,I1400084,I1400101,I1400118,I1400135,I1400152,I1400169,I1400186,I1400217,I1400234,I1400279,I1400296,I1400313,I1400344,I1400370,I1400378,I1400409,I1400426,I1400443,I1400469,I1400477,I1400494,I1400583,I1400609,I1400626,I1400634,I1400679,I1400696,I1400713,I1400730,I1400747,I1400764,I1400781,I1400812,I1400829,I1400874,I1400891,I1400908,I1400939,I1400965,I1400973,I1401004,I1401021,I1401038,I1401064,I1401072,I1401089,I1401178,I1401204,I1401221,I1401229,I1401274,I1401291,I1401308,I1401325,I1401342,I1401359,I1401376,I1401407,I1401424,I1401469,I1401486,I1401503,I1401534,I1401560,I1401568,I1401599,I1401616,I1401633,I1401659,I1401667,I1401684,I1401773,I1401799,I1401816,I1401824,I1401869,I1401886,I1401903,I1401920,I1401937,I1401954,I1401971,I1402002,I1402019,I1402064,I1402081,I1402098,I1402129,I1402155,I1402163,I1402194,I1402211,I1402228,I1402254,I1402262,I1402279,I1402368,I1402394,I1402411,I1402419,I1402464,I1402481,I1402498,I1402515,I1402532,I1402549,I1402566,I1402597,I1402614,I1402659,I1402676,I1402693,I1402724,I1402750,I1402758,I1402789,I1402806,I1402823,I1402849,I1402857,I1402874,I1402963,I1402989,I1403006,I1403014,I1403059,I1403076,I1403093,I1403110,I1403127,I1403144,I1403161,I1403192,I1403209,I1403254,I1403271,I1403288,I1403319,I1403345,I1403353,I1403384,I1403401,I1403418,I1403444,I1403452,I1403469,I1403558,I1403584,I1403601,I1403609,I1403654,I1403671,I1403688,I1403705,I1403722,I1403739,I1403756,I1403787,I1403804,I1403849,I1403866,I1403883,I1403914,I1403940,I1403948,I1403979,I1403996,I1404013,I1404039,I1404047,I1404064,I1404153,I1404179,I1404196,I1404204,I1404249,I1404266,I1404283,I1404300,I1404317,I1404334,I1404351,I1404382,I1404399,I1404444,I1404461,I1404478,I1404509,I1404535,I1404543,I1404574,I1404591,I1404608,I1404634,I1404642,I1404659,I1404748,I1404774,I1404791,I1404799,I1404844,I1404861,I1404878,I1404895,I1404912,I1404929,I1404946,I1404977,I1404994,I1405039,I1405056,I1405073,I1405104,I1405130,I1405138,I1405169,I1405186,I1405203,I1405229,I1405237,I1405254,I1405343,I1405369,I1405386,I1405394,I1405439,I1405456,I1405473,I1405490,I1405507,I1405524,I1405541,I1405572,I1405589,I1405634,I1405651,I1405668,I1405699,I1405725,I1405733,I1405764,I1405781,I1405798,I1405824,I1405832,I1405849,I1405938,I1405964,I1405981,I1405989,I1406034,I1406051,I1406068,I1406085,I1406102,I1406119,I1406136,I1406167,I1406184,I1406229,I1406246,I1406263,I1406294,I1406320,I1406328,I1406359,I1406376,I1406393,I1406419,I1406427,I1406444,I1406533,I1406559,I1406576,I1406584,I1406629,I1406646,I1406663,I1406680,I1406697,I1406714,I1406731,I1406762,I1406779,I1406824,I1406841,I1406858,I1406889,I1406915,I1406923,I1406954,I1406971,I1406988,I1407014,I1407022,I1407039,I1407128,I1407154,I1407171,I1407179,I1407224,I1407241,I1407258,I1407275,I1407292,I1407309,I1407326,I1407357,I1407374,I1407419,I1407436,I1407453,I1407484,I1407510,I1407518,I1407549,I1407566,I1407583,I1407609,I1407617,I1407634,I1407723,I1407749,I1407766,I1407774,I1407819,I1407836,I1407853,I1407870,I1407887,I1407904,I1407921,I1407952,I1407969,I1408014,I1408031,I1408048,I1408079,I1408105,I1408113,I1408144,I1408161,I1408178,I1408204,I1408212,I1408229;
not I_0 (I3602,I3570);
DFFARX1 I_1 (I1238388,I3563,I3602,I3628,);
nand I_2 (I3636,I3628,I1238388);
not I_3 (I3653,I3636);
DFFARX1 I_4 (I3653,I3563,I3602,I3594,);
DFFARX1 I_5 (I1238403,I3563,I3602,I3693,);
not I_6 (I3701,I3693);
not I_7 (I3718,I1238400);
not I_8 (I3735,I1238409);
nand I_9 (I3752,I3701,I3735);
nor I_10 (I3769,I3752,I1238400);
DFFARX1 I_11 (I3769,I3563,I3602,I3573,);
nor I_12 (I3800,I1238409,I1238400);
nand I_13 (I3817,I3693,I3800);
nor I_14 (I3834,I1238397,I1238406);
nor I_15 (I3576,I3752,I1238397);
not I_16 (I3865,I1238397);
not I_17 (I3882,I1238394);
nand I_18 (I3899,I3882,I1238385);
nand I_19 (I3916,I3718,I3899);
not I_20 (I3933,I3916);
nor I_21 (I3950,I1238394,I1238406);
nor I_22 (I3585,I3933,I3950);
nor I_23 (I3981,I1238391,I1238394);
and I_24 (I3998,I3981,I3834);
nor I_25 (I4015,I3916,I3998);
DFFARX1 I_26 (I4015,I3563,I3602,I3591,);
nor I_27 (I4046,I3636,I3998);
DFFARX1 I_28 (I4046,I3563,I3602,I3588,);
nor I_29 (I4077,I1238391,I1238385);
DFFARX1 I_30 (I4077,I3563,I3602,I4103,);
nor I_31 (I4111,I4103,I1238409);
nand I_32 (I4128,I4111,I3718);
nand I_33 (I3582,I4128,I3817);
nand I_34 (I3579,I4111,I3865);
not I_35 (I4197,I3570);
DFFARX1 I_36 (I242851,I3563,I4197,I4223,);
nand I_37 (I4231,I4223,I242851);
not I_38 (I4248,I4231);
DFFARX1 I_39 (I4248,I3563,I4197,I4189,);
DFFARX1 I_40 (I242857,I3563,I4197,I4288,);
not I_41 (I4296,I4288);
not I_42 (I4313,I242866);
not I_43 (I4330,I242860);
nand I_44 (I4347,I4296,I4330);
nor I_45 (I4364,I4347,I242866);
DFFARX1 I_46 (I4364,I3563,I4197,I4168,);
nor I_47 (I4395,I242860,I242866);
nand I_48 (I4412,I4288,I4395);
nor I_49 (I4429,I242863,I242869);
nor I_50 (I4171,I4347,I242863);
not I_51 (I4460,I242863);
not I_52 (I4477,I242872);
nand I_53 (I4494,I4477,I242848);
nand I_54 (I4511,I4313,I4494);
not I_55 (I4528,I4511);
nor I_56 (I4545,I242872,I242869);
nor I_57 (I4180,I4528,I4545);
nor I_58 (I4576,I242854,I242872);
and I_59 (I4593,I4576,I4429);
nor I_60 (I4610,I4511,I4593);
DFFARX1 I_61 (I4610,I3563,I4197,I4186,);
nor I_62 (I4641,I4231,I4593);
DFFARX1 I_63 (I4641,I3563,I4197,I4183,);
nor I_64 (I4672,I242854,I242848);
DFFARX1 I_65 (I4672,I3563,I4197,I4698,);
nor I_66 (I4706,I4698,I242860);
nand I_67 (I4723,I4706,I4313);
nand I_68 (I4177,I4723,I4412);
nand I_69 (I4174,I4706,I4460);
not I_70 (I4792,I3570);
DFFARX1 I_71 (I1234342,I3563,I4792,I4818,);
nand I_72 (I4826,I4818,I1234342);
not I_73 (I4843,I4826);
DFFARX1 I_74 (I4843,I3563,I4792,I4784,);
DFFARX1 I_75 (I1234357,I3563,I4792,I4883,);
not I_76 (I4891,I4883);
not I_77 (I4908,I1234354);
not I_78 (I4925,I1234363);
nand I_79 (I4942,I4891,I4925);
nor I_80 (I4959,I4942,I1234354);
DFFARX1 I_81 (I4959,I3563,I4792,I4763,);
nor I_82 (I4990,I1234363,I1234354);
nand I_83 (I5007,I4883,I4990);
nor I_84 (I5024,I1234351,I1234360);
nor I_85 (I4766,I4942,I1234351);
not I_86 (I5055,I1234351);
not I_87 (I5072,I1234348);
nand I_88 (I5089,I5072,I1234339);
nand I_89 (I5106,I4908,I5089);
not I_90 (I5123,I5106);
nor I_91 (I5140,I1234348,I1234360);
nor I_92 (I4775,I5123,I5140);
nor I_93 (I5171,I1234345,I1234348);
and I_94 (I5188,I5171,I5024);
nor I_95 (I5205,I5106,I5188);
DFFARX1 I_96 (I5205,I3563,I4792,I4781,);
nor I_97 (I5236,I4826,I5188);
DFFARX1 I_98 (I5236,I3563,I4792,I4778,);
nor I_99 (I5267,I1234345,I1234339);
DFFARX1 I_100 (I5267,I3563,I4792,I5293,);
nor I_101 (I5301,I5293,I1234363);
nand I_102 (I5318,I5301,I4908);
nand I_103 (I4772,I5318,I5007);
nand I_104 (I4769,I5301,I5055);
not I_105 (I5387,I3570);
DFFARX1 I_106 (I1056763,I3563,I5387,I5413,);
nand I_107 (I5421,I5413,I1056775);
not I_108 (I5438,I5421);
DFFARX1 I_109 (I5438,I3563,I5387,I5379,);
DFFARX1 I_110 (I1056760,I3563,I5387,I5478,);
not I_111 (I5486,I5478);
not I_112 (I5503,I1056763);
not I_113 (I5520,I1056757);
nand I_114 (I5537,I5486,I5520);
nor I_115 (I5554,I5537,I1056763);
DFFARX1 I_116 (I5554,I3563,I5387,I5358,);
nor I_117 (I5585,I1056757,I1056763);
nand I_118 (I5602,I5478,I5585);
nor I_119 (I5619,I1056766,I1056760);
nor I_120 (I5361,I5537,I1056766);
not I_121 (I5650,I1056766);
not I_122 (I5667,I1056772);
nand I_123 (I5684,I5667,I1056757);
nand I_124 (I5701,I5503,I5684);
not I_125 (I5718,I5701);
nor I_126 (I5735,I1056772,I1056760);
nor I_127 (I5370,I5718,I5735);
nor I_128 (I5766,I1056769,I1056772);
and I_129 (I5783,I5766,I5619);
nor I_130 (I5800,I5701,I5783);
DFFARX1 I_131 (I5800,I3563,I5387,I5376,);
nor I_132 (I5831,I5421,I5783);
DFFARX1 I_133 (I5831,I3563,I5387,I5373,);
nor I_134 (I5862,I1056769,I1056778);
DFFARX1 I_135 (I5862,I3563,I5387,I5888,);
nor I_136 (I5896,I5888,I1056757);
nand I_137 (I5913,I5896,I5503);
nand I_138 (I5367,I5913,I5602);
nand I_139 (I5364,I5896,I5650);
not I_140 (I5982,I3570);
DFFARX1 I_141 (I368646,I3563,I5982,I6008,);
nand I_142 (I6016,I6008,I368637);
not I_143 (I6033,I6016);
DFFARX1 I_144 (I6033,I3563,I5982,I5974,);
DFFARX1 I_145 (I368640,I3563,I5982,I6073,);
not I_146 (I6081,I6073);
not I_147 (I6098,I368634);
not I_148 (I6115,I368643);
nand I_149 (I6132,I6081,I6115);
nor I_150 (I6149,I6132,I368634);
DFFARX1 I_151 (I6149,I3563,I5982,I5953,);
nor I_152 (I6180,I368643,I368634);
nand I_153 (I6197,I6073,I6180);
nor I_154 (I6214,I368631,I368649);
nor I_155 (I5956,I6132,I368631);
not I_156 (I6245,I368631);
not I_157 (I6262,I368631);
nand I_158 (I6279,I6262,I368655);
nand I_159 (I6296,I6098,I6279);
not I_160 (I6313,I6296);
nor I_161 (I6330,I368631,I368649);
nor I_162 (I5965,I6313,I6330);
nor I_163 (I6361,I368652,I368631);
and I_164 (I6378,I6361,I6214);
nor I_165 (I6395,I6296,I6378);
DFFARX1 I_166 (I6395,I3563,I5982,I5971,);
nor I_167 (I6426,I6016,I6378);
DFFARX1 I_168 (I6426,I3563,I5982,I5968,);
nor I_169 (I6457,I368652,I368658);
DFFARX1 I_170 (I6457,I3563,I5982,I6483,);
nor I_171 (I6491,I6483,I368643);
nand I_172 (I6508,I6491,I6098);
nand I_173 (I5962,I6508,I6197);
nand I_174 (I5959,I6491,I6245);
not I_175 (I6577,I3570);
DFFARX1 I_176 (I332810,I3563,I6577,I6603,);
nand I_177 (I6611,I6603,I332801);
not I_178 (I6628,I6611);
DFFARX1 I_179 (I6628,I3563,I6577,I6569,);
DFFARX1 I_180 (I332804,I3563,I6577,I6668,);
not I_181 (I6676,I6668);
not I_182 (I6693,I332798);
not I_183 (I6710,I332807);
nand I_184 (I6727,I6676,I6710);
nor I_185 (I6744,I6727,I332798);
DFFARX1 I_186 (I6744,I3563,I6577,I6548,);
nor I_187 (I6775,I332807,I332798);
nand I_188 (I6792,I6668,I6775);
nor I_189 (I6809,I332795,I332813);
nor I_190 (I6551,I6727,I332795);
not I_191 (I6840,I332795);
not I_192 (I6857,I332795);
nand I_193 (I6874,I6857,I332819);
nand I_194 (I6891,I6693,I6874);
not I_195 (I6908,I6891);
nor I_196 (I6925,I332795,I332813);
nor I_197 (I6560,I6908,I6925);
nor I_198 (I6956,I332816,I332795);
and I_199 (I6973,I6956,I6809);
nor I_200 (I6990,I6891,I6973);
DFFARX1 I_201 (I6990,I3563,I6577,I6566,);
nor I_202 (I7021,I6611,I6973);
DFFARX1 I_203 (I7021,I3563,I6577,I6563,);
nor I_204 (I7052,I332816,I332822);
DFFARX1 I_205 (I7052,I3563,I6577,I7078,);
nor I_206 (I7086,I7078,I332807);
nand I_207 (I7103,I7086,I6693);
nand I_208 (I6557,I7103,I6792);
nand I_209 (I6554,I7086,I6840);
not I_210 (I7172,I3570);
DFFARX1 I_211 (I1193882,I3563,I7172,I7198,);
nand I_212 (I7206,I7198,I1193882);
not I_213 (I7223,I7206);
DFFARX1 I_214 (I7223,I3563,I7172,I7164,);
DFFARX1 I_215 (I1193897,I3563,I7172,I7263,);
not I_216 (I7271,I7263);
not I_217 (I7288,I1193894);
not I_218 (I7305,I1193903);
nand I_219 (I7322,I7271,I7305);
nor I_220 (I7339,I7322,I1193894);
DFFARX1 I_221 (I7339,I3563,I7172,I7143,);
nor I_222 (I7370,I1193903,I1193894);
nand I_223 (I7387,I7263,I7370);
nor I_224 (I7404,I1193891,I1193900);
nor I_225 (I7146,I7322,I1193891);
not I_226 (I7435,I1193891);
not I_227 (I7452,I1193888);
nand I_228 (I7469,I7452,I1193879);
nand I_229 (I7486,I7288,I7469);
not I_230 (I7503,I7486);
nor I_231 (I7520,I1193888,I1193900);
nor I_232 (I7155,I7503,I7520);
nor I_233 (I7551,I1193885,I1193888);
and I_234 (I7568,I7551,I7404);
nor I_235 (I7585,I7486,I7568);
DFFARX1 I_236 (I7585,I3563,I7172,I7161,);
nor I_237 (I7616,I7206,I7568);
DFFARX1 I_238 (I7616,I3563,I7172,I7158,);
nor I_239 (I7647,I1193885,I1193879);
DFFARX1 I_240 (I7647,I3563,I7172,I7673,);
nor I_241 (I7681,I7673,I1193903);
nand I_242 (I7698,I7681,I7288);
nand I_243 (I7152,I7698,I7387);
nand I_244 (I7149,I7681,I7435);
not I_245 (I7767,I3570);
DFFARX1 I_246 (I86171,I3563,I7767,I7793,);
nand I_247 (I7801,I7793,I86162);
not I_248 (I7818,I7801);
DFFARX1 I_249 (I7818,I3563,I7767,I7759,);
DFFARX1 I_250 (I86183,I3563,I7767,I7858,);
not I_251 (I7866,I7858);
not I_252 (I7883,I86159);
not I_253 (I7900,I86159);
nand I_254 (I7917,I7866,I7900);
nor I_255 (I7934,I7917,I86159);
DFFARX1 I_256 (I7934,I3563,I7767,I7738,);
nor I_257 (I7965,I86159,I86159);
nand I_258 (I7982,I7858,I7965);
nor I_259 (I7999,I86168,I86162);
nor I_260 (I7741,I7917,I86168);
not I_261 (I8030,I86168);
not I_262 (I8047,I86180);
nand I_263 (I8064,I8047,I86177);
nand I_264 (I8081,I7883,I8064);
not I_265 (I8098,I8081);
nor I_266 (I8115,I86180,I86162);
nor I_267 (I7750,I8098,I8115);
nor I_268 (I8146,I86174,I86180);
and I_269 (I8163,I8146,I7999);
nor I_270 (I8180,I8081,I8163);
DFFARX1 I_271 (I8180,I3563,I7767,I7756,);
nor I_272 (I8211,I7801,I8163);
DFFARX1 I_273 (I8211,I3563,I7767,I7753,);
nor I_274 (I8242,I86174,I86165);
DFFARX1 I_275 (I8242,I3563,I7767,I8268,);
nor I_276 (I8276,I8268,I86159);
nand I_277 (I8293,I8276,I7883);
nand I_278 (I7747,I8293,I7982);
nand I_279 (I7744,I8276,I8030);
not I_280 (I8362,I3570);
DFFARX1 I_281 (I39798,I3563,I8362,I8388,);
nand I_282 (I8396,I8388,I39792);
not I_283 (I8413,I8396);
DFFARX1 I_284 (I8413,I3563,I8362,I8354,);
DFFARX1 I_285 (I39807,I3563,I8362,I8453,);
not I_286 (I8461,I8453);
not I_287 (I8478,I39801);
not I_288 (I8495,I39783);
nand I_289 (I8512,I8461,I8495);
nor I_290 (I8529,I8512,I39801);
DFFARX1 I_291 (I8529,I3563,I8362,I8333,);
nor I_292 (I8560,I39783,I39801);
nand I_293 (I8577,I8453,I8560);
nor I_294 (I8594,I39789,I39795);
nor I_295 (I8336,I8512,I39789);
not I_296 (I8625,I39789);
not I_297 (I8642,I39786);
nand I_298 (I8659,I8642,I39804);
nand I_299 (I8676,I8478,I8659);
not I_300 (I8693,I8676);
nor I_301 (I8710,I39786,I39795);
nor I_302 (I8345,I8693,I8710);
nor I_303 (I8741,I39783,I39786);
and I_304 (I8758,I8741,I8594);
nor I_305 (I8775,I8676,I8758);
DFFARX1 I_306 (I8775,I3563,I8362,I8351,);
nor I_307 (I8806,I8396,I8758);
DFFARX1 I_308 (I8806,I3563,I8362,I8348,);
nor I_309 (I8837,I39783,I39786);
DFFARX1 I_310 (I8837,I3563,I8362,I8863,);
nor I_311 (I8871,I8863,I39783);
nand I_312 (I8888,I8871,I8478);
nand I_313 (I8342,I8888,I8577);
nand I_314 (I8339,I8871,I8625);
not I_315 (I8957,I3570);
DFFARX1 I_316 (I637030,I3563,I8957,I8983,);
nand I_317 (I8991,I8983,I637048);
not I_318 (I9008,I8991);
DFFARX1 I_319 (I9008,I3563,I8957,I8949,);
DFFARX1 I_320 (I637042,I3563,I8957,I9048,);
not I_321 (I9056,I9048);
not I_322 (I9073,I637033);
not I_323 (I9090,I637030);
nand I_324 (I9107,I9056,I9090);
nor I_325 (I9124,I9107,I637033);
DFFARX1 I_326 (I9124,I3563,I8957,I8928,);
nor I_327 (I9155,I637030,I637033);
nand I_328 (I9172,I9048,I9155);
nor I_329 (I9189,I637039,I637027);
nor I_330 (I8931,I9107,I637039);
not I_331 (I9220,I637039);
not I_332 (I9237,I637045);
nand I_333 (I9254,I9237,I637051);
nand I_334 (I9271,I9073,I9254);
not I_335 (I9288,I9271);
nor I_336 (I9305,I637045,I637027);
nor I_337 (I8940,I9288,I9305);
nor I_338 (I9336,I637027,I637045);
and I_339 (I9353,I9336,I9189);
nor I_340 (I9370,I9271,I9353);
DFFARX1 I_341 (I9370,I3563,I8957,I8946,);
nor I_342 (I9401,I8991,I9353);
DFFARX1 I_343 (I9401,I3563,I8957,I8943,);
nor I_344 (I9432,I637027,I637036);
DFFARX1 I_345 (I9432,I3563,I8957,I9458,);
nor I_346 (I9466,I9458,I637030);
nand I_347 (I9483,I9466,I9073);
nand I_348 (I8937,I9483,I9172);
nand I_349 (I8934,I9466,I9220);
not I_350 (I9552,I3570);
DFFARX1 I_351 (I174426,I3563,I9552,I9578,);
nand I_352 (I9586,I9578,I174426);
not I_353 (I9603,I9586);
DFFARX1 I_354 (I9603,I3563,I9552,I9544,);
DFFARX1 I_355 (I174432,I3563,I9552,I9643,);
not I_356 (I9651,I9643);
not I_357 (I9668,I174441);
not I_358 (I9685,I174435);
nand I_359 (I9702,I9651,I9685);
nor I_360 (I9719,I9702,I174441);
DFFARX1 I_361 (I9719,I3563,I9552,I9523,);
nor I_362 (I9750,I174435,I174441);
nand I_363 (I9767,I9643,I9750);
nor I_364 (I9784,I174438,I174444);
nor I_365 (I9526,I9702,I174438);
not I_366 (I9815,I174438);
not I_367 (I9832,I174447);
nand I_368 (I9849,I9832,I174423);
nand I_369 (I9866,I9668,I9849);
not I_370 (I9883,I9866);
nor I_371 (I9900,I174447,I174444);
nor I_372 (I9535,I9883,I9900);
nor I_373 (I9931,I174429,I174447);
and I_374 (I9948,I9931,I9784);
nor I_375 (I9965,I9866,I9948);
DFFARX1 I_376 (I9965,I3563,I9552,I9541,);
nor I_377 (I9996,I9586,I9948);
DFFARX1 I_378 (I9996,I3563,I9552,I9538,);
nor I_379 (I10027,I174429,I174423);
DFFARX1 I_380 (I10027,I3563,I9552,I10053,);
nor I_381 (I10061,I10053,I174435);
nand I_382 (I10078,I10061,I9668);
nand I_383 (I9532,I10078,I9767);
nand I_384 (I9529,I10061,I9815);
not I_385 (I10147,I3570);
DFFARX1 I_386 (I916834,I3563,I10147,I10173,);
nand I_387 (I10181,I10173,I916825);
not I_388 (I10198,I10181);
DFFARX1 I_389 (I10198,I3563,I10147,I10139,);
DFFARX1 I_390 (I916828,I3563,I10147,I10238,);
not I_391 (I10246,I10238);
not I_392 (I10263,I916840);
not I_393 (I10280,I916819);
nand I_394 (I10297,I10246,I10280);
nor I_395 (I10314,I10297,I916840);
DFFARX1 I_396 (I10314,I3563,I10147,I10118,);
nor I_397 (I10345,I916819,I916840);
nand I_398 (I10362,I10238,I10345);
nor I_399 (I10379,I916831,I916837);
nor I_400 (I10121,I10297,I916831);
not I_401 (I10410,I916831);
not I_402 (I10427,I916822);
nand I_403 (I10444,I10427,I916813);
nand I_404 (I10461,I10263,I10444);
not I_405 (I10478,I10461);
nor I_406 (I10495,I916822,I916837);
nor I_407 (I10130,I10478,I10495);
nor I_408 (I10526,I916813,I916822);
and I_409 (I10543,I10526,I10379);
nor I_410 (I10560,I10461,I10543);
DFFARX1 I_411 (I10560,I3563,I10147,I10136,);
nor I_412 (I10591,I10181,I10543);
DFFARX1 I_413 (I10591,I3563,I10147,I10133,);
nor I_414 (I10622,I916813,I916816);
DFFARX1 I_415 (I10622,I3563,I10147,I10648,);
nor I_416 (I10656,I10648,I916819);
nand I_417 (I10673,I10656,I10263);
nand I_418 (I10127,I10673,I10362);
nand I_419 (I10124,I10656,I10410);
not I_420 (I10742,I3570);
DFFARX1 I_421 (I708145,I3563,I10742,I10768,);
nand I_422 (I10776,I10768,I708124);
not I_423 (I10793,I10776);
DFFARX1 I_424 (I10793,I3563,I10742,I10734,);
DFFARX1 I_425 (I708133,I3563,I10742,I10833,);
not I_426 (I10841,I10833);
not I_427 (I10858,I708139);
not I_428 (I10875,I708136);
nand I_429 (I10892,I10841,I10875);
nor I_430 (I10909,I10892,I708139);
DFFARX1 I_431 (I10909,I3563,I10742,I10713,);
nor I_432 (I10940,I708136,I708139);
nand I_433 (I10957,I10833,I10940);
nor I_434 (I10974,I708127,I708121);
nor I_435 (I10716,I10892,I708127);
not I_436 (I11005,I708127);
not I_437 (I11022,I708142);
nand I_438 (I11039,I11022,I708124);
nand I_439 (I11056,I10858,I11039);
not I_440 (I11073,I11056);
nor I_441 (I11090,I708142,I708121);
nor I_442 (I10725,I11073,I11090);
nor I_443 (I11121,I708130,I708142);
and I_444 (I11138,I11121,I10974);
nor I_445 (I11155,I11056,I11138);
DFFARX1 I_446 (I11155,I3563,I10742,I10731,);
nor I_447 (I11186,I10776,I11138);
DFFARX1 I_448 (I11186,I3563,I10742,I10728,);
nor I_449 (I11217,I708130,I708121);
DFFARX1 I_450 (I11217,I3563,I10742,I11243,);
nor I_451 (I11251,I11243,I708136);
nand I_452 (I11268,I11251,I10858);
nand I_453 (I10722,I11268,I10957);
nand I_454 (I10719,I11251,I11005);
not I_455 (I11337,I3570);
DFFARX1 I_456 (I920710,I3563,I11337,I11363,);
nand I_457 (I11371,I11363,I920701);
not I_458 (I11388,I11371);
DFFARX1 I_459 (I11388,I3563,I11337,I11329,);
DFFARX1 I_460 (I920704,I3563,I11337,I11428,);
not I_461 (I11436,I11428);
not I_462 (I11453,I920716);
not I_463 (I11470,I920695);
nand I_464 (I11487,I11436,I11470);
nor I_465 (I11504,I11487,I920716);
DFFARX1 I_466 (I11504,I3563,I11337,I11308,);
nor I_467 (I11535,I920695,I920716);
nand I_468 (I11552,I11428,I11535);
nor I_469 (I11569,I920707,I920713);
nor I_470 (I11311,I11487,I920707);
not I_471 (I11600,I920707);
not I_472 (I11617,I920698);
nand I_473 (I11634,I11617,I920689);
nand I_474 (I11651,I11453,I11634);
not I_475 (I11668,I11651);
nor I_476 (I11685,I920698,I920713);
nor I_477 (I11320,I11668,I11685);
nor I_478 (I11716,I920689,I920698);
and I_479 (I11733,I11716,I11569);
nor I_480 (I11750,I11651,I11733);
DFFARX1 I_481 (I11750,I3563,I11337,I11326,);
nor I_482 (I11781,I11371,I11733);
DFFARX1 I_483 (I11781,I3563,I11337,I11323,);
nor I_484 (I11812,I920689,I920692);
DFFARX1 I_485 (I11812,I3563,I11337,I11838,);
nor I_486 (I11846,I11838,I920695);
nand I_487 (I11863,I11846,I11453);
nand I_488 (I11317,I11863,I11552);
nand I_489 (I11314,I11846,I11600);
not I_490 (I11932,I3570);
DFFARX1 I_491 (I1226828,I3563,I11932,I11958,);
nand I_492 (I11966,I11958,I1226828);
not I_493 (I11983,I11966);
DFFARX1 I_494 (I11983,I3563,I11932,I11924,);
DFFARX1 I_495 (I1226843,I3563,I11932,I12023,);
not I_496 (I12031,I12023);
not I_497 (I12048,I1226840);
not I_498 (I12065,I1226849);
nand I_499 (I12082,I12031,I12065);
nor I_500 (I12099,I12082,I1226840);
DFFARX1 I_501 (I12099,I3563,I11932,I11903,);
nor I_502 (I12130,I1226849,I1226840);
nand I_503 (I12147,I12023,I12130);
nor I_504 (I12164,I1226837,I1226846);
nor I_505 (I11906,I12082,I1226837);
not I_506 (I12195,I1226837);
not I_507 (I12212,I1226834);
nand I_508 (I12229,I12212,I1226825);
nand I_509 (I12246,I12048,I12229);
not I_510 (I12263,I12246);
nor I_511 (I12280,I1226834,I1226846);
nor I_512 (I11915,I12263,I12280);
nor I_513 (I12311,I1226831,I1226834);
and I_514 (I12328,I12311,I12164);
nor I_515 (I12345,I12246,I12328);
DFFARX1 I_516 (I12345,I3563,I11932,I11921,);
nor I_517 (I12376,I11966,I12328);
DFFARX1 I_518 (I12376,I3563,I11932,I11918,);
nor I_519 (I12407,I1226831,I1226825);
DFFARX1 I_520 (I12407,I3563,I11932,I12433,);
nor I_521 (I12441,I12433,I1226849);
nand I_522 (I12458,I12441,I12048);
nand I_523 (I11912,I12458,I12147);
nand I_524 (I11909,I12441,I12195);
not I_525 (I12527,I3570);
DFFARX1 I_526 (I1288912,I3563,I12527,I12553,);
nand I_527 (I12561,I12553,I1288918);
not I_528 (I12578,I12561);
DFFARX1 I_529 (I12578,I3563,I12527,I12519,);
DFFARX1 I_530 (I1288921,I3563,I12527,I12618,);
not I_531 (I12626,I12618);
not I_532 (I12643,I1288909);
not I_533 (I12660,I1288927);
nand I_534 (I12677,I12626,I12660);
nor I_535 (I12694,I12677,I1288909);
DFFARX1 I_536 (I12694,I3563,I12527,I12498,);
nor I_537 (I12725,I1288927,I1288909);
nand I_538 (I12742,I12618,I12725);
nor I_539 (I12759,I1288924,I1288933);
nor I_540 (I12501,I12677,I1288924);
not I_541 (I12790,I1288924);
not I_542 (I12807,I1288912);
nand I_543 (I12824,I12807,I1288930);
nand I_544 (I12841,I12643,I12824);
not I_545 (I12858,I12841);
nor I_546 (I12875,I1288912,I1288933);
nor I_547 (I12510,I12858,I12875);
nor I_548 (I12906,I1288915,I1288912);
and I_549 (I12923,I12906,I12759);
nor I_550 (I12940,I12841,I12923);
DFFARX1 I_551 (I12940,I3563,I12527,I12516,);
nor I_552 (I12971,I12561,I12923);
DFFARX1 I_553 (I12971,I3563,I12527,I12513,);
nor I_554 (I13002,I1288915,I1288909);
DFFARX1 I_555 (I13002,I3563,I12527,I13028,);
nor I_556 (I13036,I13028,I1288927);
nand I_557 (I13053,I13036,I12643);
nand I_558 (I12507,I13053,I12742);
nand I_559 (I12504,I13036,I12790);
not I_560 (I13122,I3570);
DFFARX1 I_561 (I1195038,I3563,I13122,I13148,);
nand I_562 (I13156,I13148,I1195038);
not I_563 (I13173,I13156);
DFFARX1 I_564 (I13173,I3563,I13122,I13114,);
DFFARX1 I_565 (I1195053,I3563,I13122,I13213,);
not I_566 (I13221,I13213);
not I_567 (I13238,I1195050);
not I_568 (I13255,I1195059);
nand I_569 (I13272,I13221,I13255);
nor I_570 (I13289,I13272,I1195050);
DFFARX1 I_571 (I13289,I3563,I13122,I13093,);
nor I_572 (I13320,I1195059,I1195050);
nand I_573 (I13337,I13213,I13320);
nor I_574 (I13354,I1195047,I1195056);
nor I_575 (I13096,I13272,I1195047);
not I_576 (I13385,I1195047);
not I_577 (I13402,I1195044);
nand I_578 (I13419,I13402,I1195035);
nand I_579 (I13436,I13238,I13419);
not I_580 (I13453,I13436);
nor I_581 (I13470,I1195044,I1195056);
nor I_582 (I13105,I13453,I13470);
nor I_583 (I13501,I1195041,I1195044);
and I_584 (I13518,I13501,I13354);
nor I_585 (I13535,I13436,I13518);
DFFARX1 I_586 (I13535,I3563,I13122,I13111,);
nor I_587 (I13566,I13156,I13518);
DFFARX1 I_588 (I13566,I3563,I13122,I13108,);
nor I_589 (I13597,I1195041,I1195035);
DFFARX1 I_590 (I13597,I3563,I13122,I13623,);
nor I_591 (I13631,I13623,I1195059);
nand I_592 (I13648,I13631,I13238);
nand I_593 (I13102,I13648,I13337);
nand I_594 (I13099,I13631,I13385);
not I_595 (I13717,I3570);
DFFARX1 I_596 (I426231,I3563,I13717,I13743,);
nand I_597 (I13751,I13743,I426213);
not I_598 (I13768,I13751);
DFFARX1 I_599 (I13768,I3563,I13717,I13709,);
DFFARX1 I_600 (I426225,I3563,I13717,I13808,);
not I_601 (I13816,I13808);
not I_602 (I13833,I426210);
not I_603 (I13850,I426219);
nand I_604 (I13867,I13816,I13850);
nor I_605 (I13884,I13867,I426210);
DFFARX1 I_606 (I13884,I3563,I13717,I13688,);
nor I_607 (I13915,I426219,I426210);
nand I_608 (I13932,I13808,I13915);
nor I_609 (I13949,I426216,I426237);
nor I_610 (I13691,I13867,I426216);
not I_611 (I13980,I426216);
not I_612 (I13997,I426228);
nand I_613 (I14014,I13997,I426234);
nand I_614 (I14031,I13833,I14014);
not I_615 (I14048,I14031);
nor I_616 (I14065,I426228,I426237);
nor I_617 (I13700,I14048,I14065);
nor I_618 (I14096,I426210,I426228);
and I_619 (I14113,I14096,I13949);
nor I_620 (I14130,I14031,I14113);
DFFARX1 I_621 (I14130,I3563,I13717,I13706,);
nor I_622 (I14161,I13751,I14113);
DFFARX1 I_623 (I14161,I3563,I13717,I13703,);
nor I_624 (I14192,I426210,I426222);
DFFARX1 I_625 (I14192,I3563,I13717,I14218,);
nor I_626 (I14226,I14218,I426219);
nand I_627 (I14243,I14226,I13833);
nand I_628 (I13697,I14243,I13932);
nand I_629 (I13694,I14226,I13980);
not I_630 (I14312,I3570);
DFFARX1 I_631 (I540586,I3563,I14312,I14338,);
nand I_632 (I14346,I14338,I540607);
not I_633 (I14363,I14346);
DFFARX1 I_634 (I14363,I3563,I14312,I14304,);
DFFARX1 I_635 (I540604,I3563,I14312,I14403,);
not I_636 (I14411,I14403);
not I_637 (I14428,I540586);
not I_638 (I14445,I540598);
nand I_639 (I14462,I14411,I14445);
nor I_640 (I14479,I14462,I540586);
DFFARX1 I_641 (I14479,I3563,I14312,I14283,);
nor I_642 (I14510,I540598,I540586);
nand I_643 (I14527,I14403,I14510);
nor I_644 (I14544,I540601,I540610);
nor I_645 (I14286,I14462,I540601);
not I_646 (I14575,I540601);
not I_647 (I14592,I540589);
nand I_648 (I14609,I14592,I540592);
nand I_649 (I14626,I14428,I14609);
not I_650 (I14643,I14626);
nor I_651 (I14660,I540589,I540610);
nor I_652 (I14295,I14643,I14660);
nor I_653 (I14691,I540589,I540589);
and I_654 (I14708,I14691,I14544);
nor I_655 (I14725,I14626,I14708);
DFFARX1 I_656 (I14725,I3563,I14312,I14301,);
nor I_657 (I14756,I14346,I14708);
DFFARX1 I_658 (I14756,I3563,I14312,I14298,);
nor I_659 (I14787,I540589,I540595);
DFFARX1 I_660 (I14787,I3563,I14312,I14813,);
nor I_661 (I14821,I14813,I540598);
nand I_662 (I14838,I14821,I14428);
nand I_663 (I14292,I14838,I14527);
nand I_664 (I14289,I14821,I14575);
not I_665 (I14907,I3570);
DFFARX1 I_666 (I1075837,I3563,I14907,I14933,);
nand I_667 (I14941,I14933,I1075849);
not I_668 (I14958,I14941);
DFFARX1 I_669 (I14958,I3563,I14907,I14899,);
DFFARX1 I_670 (I1075834,I3563,I14907,I14998,);
not I_671 (I15006,I14998);
not I_672 (I15023,I1075837);
not I_673 (I15040,I1075831);
nand I_674 (I15057,I15006,I15040);
nor I_675 (I15074,I15057,I1075837);
DFFARX1 I_676 (I15074,I3563,I14907,I14878,);
nor I_677 (I15105,I1075831,I1075837);
nand I_678 (I15122,I14998,I15105);
nor I_679 (I15139,I1075840,I1075834);
nor I_680 (I14881,I15057,I1075840);
not I_681 (I15170,I1075840);
not I_682 (I15187,I1075846);
nand I_683 (I15204,I15187,I1075831);
nand I_684 (I15221,I15023,I15204);
not I_685 (I15238,I15221);
nor I_686 (I15255,I1075846,I1075834);
nor I_687 (I14890,I15238,I15255);
nor I_688 (I15286,I1075843,I1075846);
and I_689 (I15303,I15286,I15139);
nor I_690 (I15320,I15221,I15303);
DFFARX1 I_691 (I15320,I3563,I14907,I14896,);
nor I_692 (I15351,I14941,I15303);
DFFARX1 I_693 (I15351,I3563,I14907,I14893,);
nor I_694 (I15382,I1075843,I1075852);
DFFARX1 I_695 (I15382,I3563,I14907,I15408,);
nor I_696 (I15416,I15408,I1075831);
nand I_697 (I15433,I15416,I15023);
nand I_698 (I14887,I15433,I15122);
nand I_699 (I14884,I15416,I15170);
not I_700 (I15502,I3570);
DFFARX1 I_701 (I1146486,I3563,I15502,I15528,);
nand I_702 (I15536,I15528,I1146486);
not I_703 (I15553,I15536);
DFFARX1 I_704 (I15553,I3563,I15502,I15494,);
DFFARX1 I_705 (I1146501,I3563,I15502,I15593,);
not I_706 (I15601,I15593);
not I_707 (I15618,I1146498);
not I_708 (I15635,I1146507);
nand I_709 (I15652,I15601,I15635);
nor I_710 (I15669,I15652,I1146498);
DFFARX1 I_711 (I15669,I3563,I15502,I15473,);
nor I_712 (I15700,I1146507,I1146498);
nand I_713 (I15717,I15593,I15700);
nor I_714 (I15734,I1146495,I1146504);
nor I_715 (I15476,I15652,I1146495);
not I_716 (I15765,I1146495);
not I_717 (I15782,I1146492);
nand I_718 (I15799,I15782,I1146483);
nand I_719 (I15816,I15618,I15799);
not I_720 (I15833,I15816);
nor I_721 (I15850,I1146492,I1146504);
nor I_722 (I15485,I15833,I15850);
nor I_723 (I15881,I1146489,I1146492);
and I_724 (I15898,I15881,I15734);
nor I_725 (I15915,I15816,I15898);
DFFARX1 I_726 (I15915,I3563,I15502,I15491,);
nor I_727 (I15946,I15536,I15898);
DFFARX1 I_728 (I15946,I3563,I15502,I15488,);
nor I_729 (I15977,I1146489,I1146483);
DFFARX1 I_730 (I15977,I3563,I15502,I16003,);
nor I_731 (I16011,I16003,I1146507);
nand I_732 (I16028,I16011,I15618);
nand I_733 (I15482,I16028,I15717);
nand I_734 (I15479,I16011,I15765);
not I_735 (I16100,I3570);
DFFARX1 I_736 (I1161535,I3563,I16100,I16126,);
DFFARX1 I_737 (I16126,I3563,I16100,I16143,);
not I_738 (I16151,I16143);
nand I_739 (I16168,I1161523,I1161514);
and I_740 (I16185,I16168,I1161511);
DFFARX1 I_741 (I16185,I3563,I16100,I16211,);
DFFARX1 I_742 (I16211,I3563,I16100,I16092,);
DFFARX1 I_743 (I16211,I3563,I16100,I16083,);
DFFARX1 I_744 (I1161517,I3563,I16100,I16256,);
nand I_745 (I16264,I16256,I1161529);
not I_746 (I16281,I16264);
nor I_747 (I16080,I16126,I16281);
DFFARX1 I_748 (I1161526,I3563,I16100,I16321,);
not I_749 (I16329,I16321);
nor I_750 (I16086,I16329,I16151);
nand I_751 (I16074,I16329,I16264);
nand I_752 (I16374,I1161520,I1161514);
and I_753 (I16391,I16374,I1161532);
DFFARX1 I_754 (I16391,I3563,I16100,I16417,);
nor I_755 (I16425,I16417,I16126);
DFFARX1 I_756 (I16425,I3563,I16100,I16068,);
not I_757 (I16456,I16417);
nor I_758 (I16473,I1161511,I1161514);
not I_759 (I16490,I16473);
nor I_760 (I16507,I16264,I16490);
nor I_761 (I16524,I16456,I16507);
DFFARX1 I_762 (I16524,I3563,I16100,I16089,);
nor I_763 (I16555,I16417,I16490);
nor I_764 (I16077,I16281,I16555);
nor I_765 (I16071,I16417,I16473);
not I_766 (I16627,I3570);
DFFARX1 I_767 (I1270345,I3563,I16627,I16653,);
DFFARX1 I_768 (I16653,I3563,I16627,I16670,);
not I_769 (I16678,I16670);
nand I_770 (I16695,I1270363,I1270357);
and I_771 (I16712,I16695,I1270366);
DFFARX1 I_772 (I16712,I3563,I16627,I16738,);
DFFARX1 I_773 (I16738,I3563,I16627,I16619,);
DFFARX1 I_774 (I16738,I3563,I16627,I16610,);
DFFARX1 I_775 (I1270351,I3563,I16627,I16783,);
nand I_776 (I16791,I16783,I1270360);
not I_777 (I16808,I16791);
nor I_778 (I16607,I16653,I16808);
DFFARX1 I_779 (I1270348,I3563,I16627,I16848,);
not I_780 (I16856,I16848);
nor I_781 (I16613,I16856,I16678);
nand I_782 (I16601,I16856,I16791);
nand I_783 (I16901,I1270369,I1270354);
and I_784 (I16918,I16901,I1270348);
DFFARX1 I_785 (I16918,I3563,I16627,I16944,);
nor I_786 (I16952,I16944,I16653);
DFFARX1 I_787 (I16952,I3563,I16627,I16595,);
not I_788 (I16983,I16944);
nor I_789 (I17000,I1270345,I1270354);
not I_790 (I17017,I17000);
nor I_791 (I17034,I16791,I17017);
nor I_792 (I17051,I16983,I17034);
DFFARX1 I_793 (I17051,I3563,I16627,I16616,);
nor I_794 (I17082,I16944,I17017);
nor I_795 (I16604,I16808,I17082);
nor I_796 (I16598,I16944,I17000);
not I_797 (I17154,I3570);
DFFARX1 I_798 (I264274,I3563,I17154,I17180,);
DFFARX1 I_799 (I17180,I3563,I17154,I17197,);
not I_800 (I17205,I17197);
nand I_801 (I17222,I264292,I264277);
and I_802 (I17239,I17222,I264280);
DFFARX1 I_803 (I17239,I3563,I17154,I17265,);
DFFARX1 I_804 (I17265,I3563,I17154,I17146,);
DFFARX1 I_805 (I17265,I3563,I17154,I17137,);
DFFARX1 I_806 (I264268,I3563,I17154,I17310,);
nand I_807 (I17318,I17310,I264271);
not I_808 (I17335,I17318);
nor I_809 (I17134,I17180,I17335);
DFFARX1 I_810 (I264283,I3563,I17154,I17375,);
not I_811 (I17383,I17375);
nor I_812 (I17140,I17383,I17205);
nand I_813 (I17128,I17383,I17318);
nand I_814 (I17428,I264289,I264286);
and I_815 (I17445,I17428,I264271);
DFFARX1 I_816 (I17445,I3563,I17154,I17471,);
nor I_817 (I17479,I17471,I17180);
DFFARX1 I_818 (I17479,I3563,I17154,I17122,);
not I_819 (I17510,I17471);
nor I_820 (I17527,I264268,I264286);
not I_821 (I17544,I17527);
nor I_822 (I17561,I17318,I17544);
nor I_823 (I17578,I17510,I17561);
DFFARX1 I_824 (I17578,I3563,I17154,I17143,);
nor I_825 (I17609,I17471,I17544);
nor I_826 (I17131,I17335,I17609);
nor I_827 (I17125,I17471,I17527);
not I_828 (I17681,I3570);
DFFARX1 I_829 (I604674,I3563,I17681,I17707,);
DFFARX1 I_830 (I17707,I3563,I17681,I17724,);
not I_831 (I17732,I17724);
nand I_832 (I17749,I604659,I604677);
and I_833 (I17766,I17749,I604671);
DFFARX1 I_834 (I17766,I3563,I17681,I17792,);
DFFARX1 I_835 (I17792,I3563,I17681,I17673,);
DFFARX1 I_836 (I17792,I3563,I17681,I17664,);
DFFARX1 I_837 (I604668,I3563,I17681,I17837,);
nand I_838 (I17845,I17837,I604659);
not I_839 (I17862,I17845);
nor I_840 (I17661,I17707,I17862);
DFFARX1 I_841 (I604662,I3563,I17681,I17902,);
not I_842 (I17910,I17902);
nor I_843 (I17667,I17910,I17732);
nand I_844 (I17655,I17910,I17845);
nand I_845 (I17955,I604683,I604665);
and I_846 (I17972,I17955,I604680);
DFFARX1 I_847 (I17972,I3563,I17681,I17998,);
nor I_848 (I18006,I17998,I17707);
DFFARX1 I_849 (I18006,I3563,I17681,I17649,);
not I_850 (I18037,I17998);
nor I_851 (I18054,I604662,I604665);
not I_852 (I18071,I18054);
nor I_853 (I18088,I17845,I18071);
nor I_854 (I18105,I18037,I18088);
DFFARX1 I_855 (I18105,I3563,I17681,I17670,);
nor I_856 (I18136,I17998,I18071);
nor I_857 (I17658,I17862,I18136);
nor I_858 (I17652,I17998,I18054);
not I_859 (I18208,I3570);
DFFARX1 I_860 (I838469,I3563,I18208,I18234,);
DFFARX1 I_861 (I18234,I3563,I18208,I18251,);
not I_862 (I18259,I18251);
nand I_863 (I18276,I838460,I838481);
and I_864 (I18293,I18276,I838463);
DFFARX1 I_865 (I18293,I3563,I18208,I18319,);
DFFARX1 I_866 (I18319,I3563,I18208,I18200,);
DFFARX1 I_867 (I18319,I3563,I18208,I18191,);
DFFARX1 I_868 (I838463,I3563,I18208,I18364,);
nand I_869 (I18372,I18364,I838478);
not I_870 (I18389,I18372);
nor I_871 (I18188,I18234,I18389);
DFFARX1 I_872 (I838472,I3563,I18208,I18429,);
not I_873 (I18437,I18429);
nor I_874 (I18194,I18437,I18259);
nand I_875 (I18182,I18437,I18372);
nand I_876 (I18482,I838466,I838475);
and I_877 (I18499,I18482,I838460);
DFFARX1 I_878 (I18499,I3563,I18208,I18525,);
nor I_879 (I18533,I18525,I18234);
DFFARX1 I_880 (I18533,I3563,I18208,I18176,);
not I_881 (I18564,I18525);
nor I_882 (I18581,I838466,I838475);
not I_883 (I18598,I18581);
nor I_884 (I18615,I18372,I18598);
nor I_885 (I18632,I18564,I18615);
DFFARX1 I_886 (I18632,I3563,I18208,I18197,);
nor I_887 (I18663,I18525,I18598);
nor I_888 (I18185,I18389,I18663);
nor I_889 (I18179,I18525,I18581);
not I_890 (I18735,I3570);
DFFARX1 I_891 (I97229,I3563,I18735,I18761,);
DFFARX1 I_892 (I18761,I3563,I18735,I18778,);
not I_893 (I18786,I18778);
nand I_894 (I18803,I97229,I97244);
and I_895 (I18820,I18803,I97247);
DFFARX1 I_896 (I18820,I3563,I18735,I18846,);
DFFARX1 I_897 (I18846,I3563,I18735,I18727,);
DFFARX1 I_898 (I18846,I3563,I18735,I18718,);
DFFARX1 I_899 (I97241,I3563,I18735,I18891,);
nand I_900 (I18899,I18891,I97250);
not I_901 (I18916,I18899);
nor I_902 (I18715,I18761,I18916);
DFFARX1 I_903 (I97226,I3563,I18735,I18956,);
not I_904 (I18964,I18956);
nor I_905 (I18721,I18964,I18786);
nand I_906 (I18709,I18964,I18899);
nand I_907 (I19009,I97226,I97232);
and I_908 (I19026,I19009,I97235);
DFFARX1 I_909 (I19026,I3563,I18735,I19052,);
nor I_910 (I19060,I19052,I18761);
DFFARX1 I_911 (I19060,I3563,I18735,I18703,);
not I_912 (I19091,I19052);
nor I_913 (I19108,I97238,I97232);
not I_914 (I19125,I19108);
nor I_915 (I19142,I18899,I19125);
nor I_916 (I19159,I19091,I19142);
DFFARX1 I_917 (I19159,I3563,I18735,I18724,);
nor I_918 (I19190,I19052,I19125);
nor I_919 (I18712,I18916,I19190);
nor I_920 (I18706,I19052,I19108);
not I_921 (I19262,I3570);
DFFARX1 I_922 (I880629,I3563,I19262,I19288,);
DFFARX1 I_923 (I19288,I3563,I19262,I19305,);
not I_924 (I19313,I19305);
nand I_925 (I19330,I880620,I880641);
and I_926 (I19347,I19330,I880623);
DFFARX1 I_927 (I19347,I3563,I19262,I19373,);
DFFARX1 I_928 (I19373,I3563,I19262,I19254,);
DFFARX1 I_929 (I19373,I3563,I19262,I19245,);
DFFARX1 I_930 (I880623,I3563,I19262,I19418,);
nand I_931 (I19426,I19418,I880638);
not I_932 (I19443,I19426);
nor I_933 (I19242,I19288,I19443);
DFFARX1 I_934 (I880632,I3563,I19262,I19483,);
not I_935 (I19491,I19483);
nor I_936 (I19248,I19491,I19313);
nand I_937 (I19236,I19491,I19426);
nand I_938 (I19536,I880626,I880635);
and I_939 (I19553,I19536,I880620);
DFFARX1 I_940 (I19553,I3563,I19262,I19579,);
nor I_941 (I19587,I19579,I19288);
DFFARX1 I_942 (I19587,I3563,I19262,I19230,);
not I_943 (I19618,I19579);
nor I_944 (I19635,I880626,I880635);
not I_945 (I19652,I19635);
nor I_946 (I19669,I19426,I19652);
nor I_947 (I19686,I19618,I19669);
DFFARX1 I_948 (I19686,I3563,I19262,I19251,);
nor I_949 (I19717,I19579,I19652);
nor I_950 (I19239,I19443,I19717);
nor I_951 (I19233,I19579,I19635);
not I_952 (I19789,I3570);
DFFARX1 I_953 (I83000,I3563,I19789,I19815,);
DFFARX1 I_954 (I19815,I3563,I19789,I19832,);
not I_955 (I19840,I19832);
nand I_956 (I19857,I83000,I83015);
and I_957 (I19874,I19857,I83018);
DFFARX1 I_958 (I19874,I3563,I19789,I19900,);
DFFARX1 I_959 (I19900,I3563,I19789,I19781,);
DFFARX1 I_960 (I19900,I3563,I19789,I19772,);
DFFARX1 I_961 (I83012,I3563,I19789,I19945,);
nand I_962 (I19953,I19945,I83021);
not I_963 (I19970,I19953);
nor I_964 (I19769,I19815,I19970);
DFFARX1 I_965 (I82997,I3563,I19789,I20010,);
not I_966 (I20018,I20010);
nor I_967 (I19775,I20018,I19840);
nand I_968 (I19763,I20018,I19953);
nand I_969 (I20063,I82997,I83003);
and I_970 (I20080,I20063,I83006);
DFFARX1 I_971 (I20080,I3563,I19789,I20106,);
nor I_972 (I20114,I20106,I19815);
DFFARX1 I_973 (I20114,I3563,I19789,I19757,);
not I_974 (I20145,I20106);
nor I_975 (I20162,I83009,I83003);
not I_976 (I20179,I20162);
nor I_977 (I20196,I19953,I20179);
nor I_978 (I20213,I20145,I20196);
DFFARX1 I_979 (I20213,I3563,I19789,I19778,);
nor I_980 (I20244,I20106,I20179);
nor I_981 (I19766,I19970,I20244);
nor I_982 (I19760,I20106,I20162);
not I_983 (I20316,I3570);
DFFARX1 I_984 (I479522,I3563,I20316,I20342,);
DFFARX1 I_985 (I20342,I3563,I20316,I20359,);
not I_986 (I20367,I20359);
nand I_987 (I20384,I479522,I479525);
and I_988 (I20401,I20384,I479546);
DFFARX1 I_989 (I20401,I3563,I20316,I20427,);
DFFARX1 I_990 (I20427,I3563,I20316,I20308,);
DFFARX1 I_991 (I20427,I3563,I20316,I20299,);
DFFARX1 I_992 (I479534,I3563,I20316,I20472,);
nand I_993 (I20480,I20472,I479537);
not I_994 (I20497,I20480);
nor I_995 (I20296,I20342,I20497);
DFFARX1 I_996 (I479543,I3563,I20316,I20537,);
not I_997 (I20545,I20537);
nor I_998 (I20302,I20545,I20367);
nand I_999 (I20290,I20545,I20480);
nand I_1000 (I20590,I479540,I479528);
and I_1001 (I20607,I20590,I479531);
DFFARX1 I_1002 (I20607,I3563,I20316,I20633,);
nor I_1003 (I20641,I20633,I20342);
DFFARX1 I_1004 (I20641,I3563,I20316,I20284,);
not I_1005 (I20672,I20633);
nor I_1006 (I20689,I479549,I479528);
not I_1007 (I20706,I20689);
nor I_1008 (I20723,I20480,I20706);
nor I_1009 (I20740,I20672,I20723);
DFFARX1 I_1010 (I20740,I3563,I20316,I20305,);
nor I_1011 (I20771,I20633,I20706);
nor I_1012 (I20293,I20497,I20771);
nor I_1013 (I20287,I20633,I20689);
not I_1014 (I20843,I3570);
DFFARX1 I_1015 (I1330933,I3563,I20843,I20869,);
DFFARX1 I_1016 (I20869,I3563,I20843,I20886,);
not I_1017 (I20894,I20886);
nand I_1018 (I20911,I1330936,I1330942);
and I_1019 (I20928,I20911,I1330951);
DFFARX1 I_1020 (I20928,I3563,I20843,I20954,);
DFFARX1 I_1021 (I20954,I3563,I20843,I20835,);
DFFARX1 I_1022 (I20954,I3563,I20843,I20826,);
DFFARX1 I_1023 (I1330954,I3563,I20843,I20999,);
nand I_1024 (I21007,I20999,I1330945);
not I_1025 (I21024,I21007);
nor I_1026 (I20823,I20869,I21024);
DFFARX1 I_1027 (I1330933,I3563,I20843,I21064,);
not I_1028 (I21072,I21064);
nor I_1029 (I20829,I21072,I20894);
nand I_1030 (I20817,I21072,I21007);
nand I_1031 (I21117,I1330960,I1330939);
and I_1032 (I21134,I21117,I1330948);
DFFARX1 I_1033 (I21134,I3563,I20843,I21160,);
nor I_1034 (I21168,I21160,I20869);
DFFARX1 I_1035 (I21168,I3563,I20843,I20811,);
not I_1036 (I21199,I21160);
nor I_1037 (I21216,I1330957,I1330939);
not I_1038 (I21233,I21216);
nor I_1039 (I21250,I21007,I21233);
nor I_1040 (I21267,I21199,I21250);
DFFARX1 I_1041 (I21267,I3563,I20843,I20832,);
nor I_1042 (I21298,I21160,I21233);
nor I_1043 (I20820,I21024,I21298);
nor I_1044 (I20814,I21160,I21216);
not I_1045 (I21370,I3570);
DFFARX1 I_1046 (I1200261,I3563,I21370,I21396,);
DFFARX1 I_1047 (I21396,I3563,I21370,I21413,);
not I_1048 (I21421,I21413);
nand I_1049 (I21438,I1200249,I1200240);
and I_1050 (I21455,I21438,I1200237);
DFFARX1 I_1051 (I21455,I3563,I21370,I21481,);
DFFARX1 I_1052 (I21481,I3563,I21370,I21362,);
DFFARX1 I_1053 (I21481,I3563,I21370,I21353,);
DFFARX1 I_1054 (I1200243,I3563,I21370,I21526,);
nand I_1055 (I21534,I21526,I1200255);
not I_1056 (I21551,I21534);
nor I_1057 (I21350,I21396,I21551);
DFFARX1 I_1058 (I1200252,I3563,I21370,I21591,);
not I_1059 (I21599,I21591);
nor I_1060 (I21356,I21599,I21421);
nand I_1061 (I21344,I21599,I21534);
nand I_1062 (I21644,I1200246,I1200240);
and I_1063 (I21661,I21644,I1200258);
DFFARX1 I_1064 (I21661,I3563,I21370,I21687,);
nor I_1065 (I21695,I21687,I21396);
DFFARX1 I_1066 (I21695,I3563,I21370,I21338,);
not I_1067 (I21726,I21687);
nor I_1068 (I21743,I1200237,I1200240);
not I_1069 (I21760,I21743);
nor I_1070 (I21777,I21534,I21760);
nor I_1071 (I21794,I21726,I21777);
DFFARX1 I_1072 (I21794,I3563,I21370,I21359,);
nor I_1073 (I21825,I21687,I21760);
nor I_1074 (I21347,I21551,I21825);
nor I_1075 (I21341,I21687,I21743);
not I_1076 (I21897,I3570);
DFFARX1 I_1077 (I870616,I3563,I21897,I21923,);
DFFARX1 I_1078 (I21923,I3563,I21897,I21940,);
not I_1079 (I21948,I21940);
nand I_1080 (I21965,I870607,I870628);
and I_1081 (I21982,I21965,I870610);
DFFARX1 I_1082 (I21982,I3563,I21897,I22008,);
DFFARX1 I_1083 (I22008,I3563,I21897,I21889,);
DFFARX1 I_1084 (I22008,I3563,I21897,I21880,);
DFFARX1 I_1085 (I870610,I3563,I21897,I22053,);
nand I_1086 (I22061,I22053,I870625);
not I_1087 (I22078,I22061);
nor I_1088 (I21877,I21923,I22078);
DFFARX1 I_1089 (I870619,I3563,I21897,I22118,);
not I_1090 (I22126,I22118);
nor I_1091 (I21883,I22126,I21948);
nand I_1092 (I21871,I22126,I22061);
nand I_1093 (I22171,I870613,I870622);
and I_1094 (I22188,I22171,I870607);
DFFARX1 I_1095 (I22188,I3563,I21897,I22214,);
nor I_1096 (I22222,I22214,I21923);
DFFARX1 I_1097 (I22222,I3563,I21897,I21865,);
not I_1098 (I22253,I22214);
nor I_1099 (I22270,I870613,I870622);
not I_1100 (I22287,I22270);
nor I_1101 (I22304,I22061,I22287);
nor I_1102 (I22321,I22253,I22304);
DFFARX1 I_1103 (I22321,I3563,I21897,I21886,);
nor I_1104 (I22352,I22214,I22287);
nor I_1105 (I21874,I22078,I22352);
nor I_1106 (I21868,I22214,I22270);
not I_1107 (I22424,I3570);
DFFARX1 I_1108 (I750899,I3563,I22424,I22450,);
DFFARX1 I_1109 (I22450,I3563,I22424,I22467,);
not I_1110 (I22475,I22467);
nand I_1111 (I22492,I750914,I750917);
and I_1112 (I22509,I22492,I750896);
DFFARX1 I_1113 (I22509,I3563,I22424,I22535,);
DFFARX1 I_1114 (I22535,I3563,I22424,I22416,);
DFFARX1 I_1115 (I22535,I3563,I22424,I22407,);
DFFARX1 I_1116 (I750902,I3563,I22424,I22580,);
nand I_1117 (I22588,I22580,I750908);
not I_1118 (I22605,I22588);
nor I_1119 (I22404,I22450,I22605);
DFFARX1 I_1120 (I750896,I3563,I22424,I22645,);
not I_1121 (I22653,I22645);
nor I_1122 (I22410,I22653,I22475);
nand I_1123 (I22398,I22653,I22588);
nand I_1124 (I22698,I750911,I750893);
and I_1125 (I22715,I22698,I750905);
DFFARX1 I_1126 (I22715,I3563,I22424,I22741,);
nor I_1127 (I22749,I22741,I22450);
DFFARX1 I_1128 (I22749,I3563,I22424,I22392,);
not I_1129 (I22780,I22741);
nor I_1130 (I22797,I750893,I750893);
not I_1131 (I22814,I22797);
nor I_1132 (I22831,I22588,I22814);
nor I_1133 (I22848,I22780,I22831);
DFFARX1 I_1134 (I22848,I3563,I22424,I22413,);
nor I_1135 (I22879,I22741,I22814);
nor I_1136 (I22401,I22605,I22879);
nor I_1137 (I22395,I22741,I22797);
not I_1138 (I22951,I3570);
DFFARX1 I_1139 (I650914,I3563,I22951,I22977,);
DFFARX1 I_1140 (I22977,I3563,I22951,I22994,);
not I_1141 (I23002,I22994);
nand I_1142 (I23019,I650899,I650917);
and I_1143 (I23036,I23019,I650911);
DFFARX1 I_1144 (I23036,I3563,I22951,I23062,);
DFFARX1 I_1145 (I23062,I3563,I22951,I22943,);
DFFARX1 I_1146 (I23062,I3563,I22951,I22934,);
DFFARX1 I_1147 (I650908,I3563,I22951,I23107,);
nand I_1148 (I23115,I23107,I650899);
not I_1149 (I23132,I23115);
nor I_1150 (I22931,I22977,I23132);
DFFARX1 I_1151 (I650902,I3563,I22951,I23172,);
not I_1152 (I23180,I23172);
nor I_1153 (I22937,I23180,I23002);
nand I_1154 (I22925,I23180,I23115);
nand I_1155 (I23225,I650923,I650905);
and I_1156 (I23242,I23225,I650920);
DFFARX1 I_1157 (I23242,I3563,I22951,I23268,);
nor I_1158 (I23276,I23268,I22977);
DFFARX1 I_1159 (I23276,I3563,I22951,I22919,);
not I_1160 (I23307,I23268);
nor I_1161 (I23324,I650902,I650905);
not I_1162 (I23341,I23324);
nor I_1163 (I23358,I23115,I23341);
nor I_1164 (I23375,I23307,I23358);
DFFARX1 I_1165 (I23375,I3563,I22951,I22940,);
nor I_1166 (I23406,I23268,I23341);
nor I_1167 (I22928,I23132,I23406);
nor I_1168 (I22922,I23268,I23324);
not I_1169 (I23478,I3570);
DFFARX1 I_1170 (I431106,I3563,I23478,I23504,);
DFFARX1 I_1171 (I23504,I3563,I23478,I23521,);
not I_1172 (I23529,I23521);
nand I_1173 (I23546,I431106,I431109);
and I_1174 (I23563,I23546,I431130);
DFFARX1 I_1175 (I23563,I3563,I23478,I23589,);
DFFARX1 I_1176 (I23589,I3563,I23478,I23470,);
DFFARX1 I_1177 (I23589,I3563,I23478,I23461,);
DFFARX1 I_1178 (I431118,I3563,I23478,I23634,);
nand I_1179 (I23642,I23634,I431121);
not I_1180 (I23659,I23642);
nor I_1181 (I23458,I23504,I23659);
DFFARX1 I_1182 (I431127,I3563,I23478,I23699,);
not I_1183 (I23707,I23699);
nor I_1184 (I23464,I23707,I23529);
nand I_1185 (I23452,I23707,I23642);
nand I_1186 (I23752,I431124,I431112);
and I_1187 (I23769,I23752,I431115);
DFFARX1 I_1188 (I23769,I3563,I23478,I23795,);
nor I_1189 (I23803,I23795,I23504);
DFFARX1 I_1190 (I23803,I3563,I23478,I23446,);
not I_1191 (I23834,I23795);
nor I_1192 (I23851,I431133,I431112);
not I_1193 (I23868,I23851);
nor I_1194 (I23885,I23642,I23868);
nor I_1195 (I23902,I23834,I23885);
DFFARX1 I_1196 (I23902,I3563,I23478,I23467,);
nor I_1197 (I23933,I23795,I23868);
nor I_1198 (I23455,I23659,I23933);
nor I_1199 (I23449,I23795,I23851);
not I_1200 (I24005,I3570);
DFFARX1 I_1201 (I248209,I3563,I24005,I24031,);
DFFARX1 I_1202 (I24031,I3563,I24005,I24048,);
not I_1203 (I24056,I24048);
nand I_1204 (I24073,I248227,I248212);
and I_1205 (I24090,I24073,I248215);
DFFARX1 I_1206 (I24090,I3563,I24005,I24116,);
DFFARX1 I_1207 (I24116,I3563,I24005,I23997,);
DFFARX1 I_1208 (I24116,I3563,I24005,I23988,);
DFFARX1 I_1209 (I248203,I3563,I24005,I24161,);
nand I_1210 (I24169,I24161,I248206);
not I_1211 (I24186,I24169);
nor I_1212 (I23985,I24031,I24186);
DFFARX1 I_1213 (I248218,I3563,I24005,I24226,);
not I_1214 (I24234,I24226);
nor I_1215 (I23991,I24234,I24056);
nand I_1216 (I23979,I24234,I24169);
nand I_1217 (I24279,I248224,I248221);
and I_1218 (I24296,I24279,I248206);
DFFARX1 I_1219 (I24296,I3563,I24005,I24322,);
nor I_1220 (I24330,I24322,I24031);
DFFARX1 I_1221 (I24330,I3563,I24005,I23973,);
not I_1222 (I24361,I24322);
nor I_1223 (I24378,I248203,I248221);
not I_1224 (I24395,I24378);
nor I_1225 (I24412,I24169,I24395);
nor I_1226 (I24429,I24361,I24412);
DFFARX1 I_1227 (I24429,I3563,I24005,I23994,);
nor I_1228 (I24460,I24322,I24395);
nor I_1229 (I23982,I24186,I24460);
nor I_1230 (I23976,I24322,I24378);
not I_1231 (I24532,I3570);
DFFARX1 I_1232 (I516514,I3563,I24532,I24558,);
DFFARX1 I_1233 (I24558,I3563,I24532,I24575,);
not I_1234 (I24583,I24575);
nand I_1235 (I24600,I516514,I516517);
and I_1236 (I24617,I24600,I516538);
DFFARX1 I_1237 (I24617,I3563,I24532,I24643,);
DFFARX1 I_1238 (I24643,I3563,I24532,I24524,);
DFFARX1 I_1239 (I24643,I3563,I24532,I24515,);
DFFARX1 I_1240 (I516526,I3563,I24532,I24688,);
nand I_1241 (I24696,I24688,I516529);
not I_1242 (I24713,I24696);
nor I_1243 (I24512,I24558,I24713);
DFFARX1 I_1244 (I516535,I3563,I24532,I24753,);
not I_1245 (I24761,I24753);
nor I_1246 (I24518,I24761,I24583);
nand I_1247 (I24506,I24761,I24696);
nand I_1248 (I24806,I516532,I516520);
and I_1249 (I24823,I24806,I516523);
DFFARX1 I_1250 (I24823,I3563,I24532,I24849,);
nor I_1251 (I24857,I24849,I24558);
DFFARX1 I_1252 (I24857,I3563,I24532,I24500,);
not I_1253 (I24888,I24849);
nor I_1254 (I24905,I516541,I516520);
not I_1255 (I24922,I24905);
nor I_1256 (I24939,I24696,I24922);
nor I_1257 (I24956,I24888,I24939);
DFFARX1 I_1258 (I24956,I3563,I24532,I24521,);
nor I_1259 (I24987,I24849,I24922);
nor I_1260 (I24509,I24713,I24987);
nor I_1261 (I24503,I24849,I24905);
not I_1262 (I25059,I3570);
DFFARX1 I_1263 (I1163847,I3563,I25059,I25085,);
DFFARX1 I_1264 (I25085,I3563,I25059,I25102,);
not I_1265 (I25110,I25102);
nand I_1266 (I25127,I1163835,I1163826);
and I_1267 (I25144,I25127,I1163823);
DFFARX1 I_1268 (I25144,I3563,I25059,I25170,);
DFFARX1 I_1269 (I25170,I3563,I25059,I25051,);
DFFARX1 I_1270 (I25170,I3563,I25059,I25042,);
DFFARX1 I_1271 (I1163829,I3563,I25059,I25215,);
nand I_1272 (I25223,I25215,I1163841);
not I_1273 (I25240,I25223);
nor I_1274 (I25039,I25085,I25240);
DFFARX1 I_1275 (I1163838,I3563,I25059,I25280,);
not I_1276 (I25288,I25280);
nor I_1277 (I25045,I25288,I25110);
nand I_1278 (I25033,I25288,I25223);
nand I_1279 (I25333,I1163832,I1163826);
and I_1280 (I25350,I25333,I1163844);
DFFARX1 I_1281 (I25350,I3563,I25059,I25376,);
nor I_1282 (I25384,I25376,I25085);
DFFARX1 I_1283 (I25384,I3563,I25059,I25027,);
not I_1284 (I25415,I25376);
nor I_1285 (I25432,I1163823,I1163826);
not I_1286 (I25449,I25432);
nor I_1287 (I25466,I25223,I25449);
nor I_1288 (I25483,I25415,I25466);
DFFARX1 I_1289 (I25483,I3563,I25059,I25048,);
nor I_1290 (I25514,I25376,I25449);
nor I_1291 (I25036,I25240,I25514);
nor I_1292 (I25030,I25376,I25432);
not I_1293 (I25586,I3570);
DFFARX1 I_1294 (I1320136,I3563,I25586,I25612,);
DFFARX1 I_1295 (I25612,I3563,I25586,I25629,);
not I_1296 (I25637,I25629);
nand I_1297 (I25654,I1320139,I1320133);
and I_1298 (I25671,I25654,I1320142);
DFFARX1 I_1299 (I25671,I3563,I25586,I25697,);
DFFARX1 I_1300 (I25697,I3563,I25586,I25578,);
DFFARX1 I_1301 (I25697,I3563,I25586,I25569,);
DFFARX1 I_1302 (I1320130,I3563,I25586,I25742,);
nand I_1303 (I25750,I25742,I1320145);
not I_1304 (I25767,I25750);
nor I_1305 (I25566,I25612,I25767);
DFFARX1 I_1306 (I1320121,I3563,I25586,I25807,);
not I_1307 (I25815,I25807);
nor I_1308 (I25572,I25815,I25637);
nand I_1309 (I25560,I25815,I25750);
nand I_1310 (I25860,I1320124,I1320124);
and I_1311 (I25877,I25860,I1320121);
DFFARX1 I_1312 (I25877,I3563,I25586,I25903,);
nor I_1313 (I25911,I25903,I25612);
DFFARX1 I_1314 (I25911,I3563,I25586,I25554,);
not I_1315 (I25942,I25903);
nor I_1316 (I25959,I1320127,I1320124);
not I_1317 (I25976,I25959);
nor I_1318 (I25993,I25750,I25976);
nor I_1319 (I26010,I25942,I25993);
DFFARX1 I_1320 (I26010,I3563,I25586,I25575,);
nor I_1321 (I26041,I25903,I25976);
nor I_1322 (I25563,I25767,I26041);
nor I_1323 (I25557,I25903,I25959);
not I_1324 (I26113,I3570);
DFFARX1 I_1325 (I138335,I3563,I26113,I26139,);
DFFARX1 I_1326 (I26139,I3563,I26113,I26156,);
not I_1327 (I26164,I26156);
nand I_1328 (I26181,I138335,I138350);
and I_1329 (I26198,I26181,I138353);
DFFARX1 I_1330 (I26198,I3563,I26113,I26224,);
DFFARX1 I_1331 (I26224,I3563,I26113,I26105,);
DFFARX1 I_1332 (I26224,I3563,I26113,I26096,);
DFFARX1 I_1333 (I138347,I3563,I26113,I26269,);
nand I_1334 (I26277,I26269,I138356);
not I_1335 (I26294,I26277);
nor I_1336 (I26093,I26139,I26294);
DFFARX1 I_1337 (I138332,I3563,I26113,I26334,);
not I_1338 (I26342,I26334);
nor I_1339 (I26099,I26342,I26164);
nand I_1340 (I26087,I26342,I26277);
nand I_1341 (I26387,I138332,I138338);
and I_1342 (I26404,I26387,I138341);
DFFARX1 I_1343 (I26404,I3563,I26113,I26430,);
nor I_1344 (I26438,I26430,I26139);
DFFARX1 I_1345 (I26438,I3563,I26113,I26081,);
not I_1346 (I26469,I26430);
nor I_1347 (I26486,I138344,I138338);
not I_1348 (I26503,I26486);
nor I_1349 (I26520,I26277,I26503);
nor I_1350 (I26537,I26469,I26520);
DFFARX1 I_1351 (I26537,I3563,I26113,I26102,);
nor I_1352 (I26568,I26430,I26503);
nor I_1353 (I26090,I26294,I26568);
nor I_1354 (I26084,I26430,I26486);
not I_1355 (I26640,I3570);
DFFARX1 I_1356 (I627216,I3563,I26640,I26666,);
DFFARX1 I_1357 (I26666,I3563,I26640,I26683,);
not I_1358 (I26691,I26683);
nand I_1359 (I26708,I627201,I627219);
and I_1360 (I26725,I26708,I627213);
DFFARX1 I_1361 (I26725,I3563,I26640,I26751,);
DFFARX1 I_1362 (I26751,I3563,I26640,I26632,);
DFFARX1 I_1363 (I26751,I3563,I26640,I26623,);
DFFARX1 I_1364 (I627210,I3563,I26640,I26796,);
nand I_1365 (I26804,I26796,I627201);
not I_1366 (I26821,I26804);
nor I_1367 (I26620,I26666,I26821);
DFFARX1 I_1368 (I627204,I3563,I26640,I26861,);
not I_1369 (I26869,I26861);
nor I_1370 (I26626,I26869,I26691);
nand I_1371 (I26614,I26869,I26804);
nand I_1372 (I26914,I627225,I627207);
and I_1373 (I26931,I26914,I627222);
DFFARX1 I_1374 (I26931,I3563,I26640,I26957,);
nor I_1375 (I26965,I26957,I26666);
DFFARX1 I_1376 (I26965,I3563,I26640,I26608,);
not I_1377 (I26996,I26957);
nor I_1378 (I27013,I627204,I627207);
not I_1379 (I27030,I27013);
nor I_1380 (I27047,I26804,I27030);
nor I_1381 (I27064,I26996,I27047);
DFFARX1 I_1382 (I27064,I3563,I26640,I26629,);
nor I_1383 (I27095,I26957,I27030);
nor I_1384 (I26617,I26821,I27095);
nor I_1385 (I26611,I26957,I27013);
not I_1386 (I27167,I3570);
DFFARX1 I_1387 (I745119,I3563,I27167,I27193,);
DFFARX1 I_1388 (I27193,I3563,I27167,I27210,);
not I_1389 (I27218,I27210);
nand I_1390 (I27235,I745134,I745137);
and I_1391 (I27252,I27235,I745116);
DFFARX1 I_1392 (I27252,I3563,I27167,I27278,);
DFFARX1 I_1393 (I27278,I3563,I27167,I27159,);
DFFARX1 I_1394 (I27278,I3563,I27167,I27150,);
DFFARX1 I_1395 (I745122,I3563,I27167,I27323,);
nand I_1396 (I27331,I27323,I745128);
not I_1397 (I27348,I27331);
nor I_1398 (I27147,I27193,I27348);
DFFARX1 I_1399 (I745116,I3563,I27167,I27388,);
not I_1400 (I27396,I27388);
nor I_1401 (I27153,I27396,I27218);
nand I_1402 (I27141,I27396,I27331);
nand I_1403 (I27441,I745131,I745113);
and I_1404 (I27458,I27441,I745125);
DFFARX1 I_1405 (I27458,I3563,I27167,I27484,);
nor I_1406 (I27492,I27484,I27193);
DFFARX1 I_1407 (I27492,I3563,I27167,I27135,);
not I_1408 (I27523,I27484);
nor I_1409 (I27540,I745113,I745113);
not I_1410 (I27557,I27540);
nor I_1411 (I27574,I27331,I27557);
nor I_1412 (I27591,I27523,I27574);
DFFARX1 I_1413 (I27591,I3563,I27167,I27156,);
nor I_1414 (I27622,I27484,I27557);
nor I_1415 (I27144,I27348,I27622);
nor I_1416 (I27138,I27484,I27540);
not I_1417 (I27694,I3570);
DFFARX1 I_1418 (I58231,I3563,I27694,I27720,);
DFFARX1 I_1419 (I27720,I3563,I27694,I27737,);
not I_1420 (I27745,I27737);
nand I_1421 (I27762,I58231,I58246);
and I_1422 (I27779,I27762,I58249);
DFFARX1 I_1423 (I27779,I3563,I27694,I27805,);
DFFARX1 I_1424 (I27805,I3563,I27694,I27686,);
DFFARX1 I_1425 (I27805,I3563,I27694,I27677,);
DFFARX1 I_1426 (I58243,I3563,I27694,I27850,);
nand I_1427 (I27858,I27850,I58252);
not I_1428 (I27875,I27858);
nor I_1429 (I27674,I27720,I27875);
DFFARX1 I_1430 (I58228,I3563,I27694,I27915,);
not I_1431 (I27923,I27915);
nor I_1432 (I27680,I27923,I27745);
nand I_1433 (I27668,I27923,I27858);
nand I_1434 (I27968,I58228,I58234);
and I_1435 (I27985,I27968,I58237);
DFFARX1 I_1436 (I27985,I3563,I27694,I28011,);
nor I_1437 (I28019,I28011,I27720);
DFFARX1 I_1438 (I28019,I3563,I27694,I27662,);
not I_1439 (I28050,I28011);
nor I_1440 (I28067,I58240,I58234);
not I_1441 (I28084,I28067);
nor I_1442 (I28101,I27858,I28084);
nor I_1443 (I28118,I28050,I28101);
DFFARX1 I_1444 (I28118,I3563,I27694,I27683,);
nor I_1445 (I28149,I28011,I28084);
nor I_1446 (I27671,I27875,I28149);
nor I_1447 (I27665,I28011,I28067);
not I_1448 (I28221,I3570);
DFFARX1 I_1449 (I1274153,I3563,I28221,I28247,);
DFFARX1 I_1450 (I28247,I3563,I28221,I28264,);
not I_1451 (I28272,I28264);
nand I_1452 (I28289,I1274171,I1274165);
and I_1453 (I28306,I28289,I1274174);
DFFARX1 I_1454 (I28306,I3563,I28221,I28332,);
DFFARX1 I_1455 (I28332,I3563,I28221,I28213,);
DFFARX1 I_1456 (I28332,I3563,I28221,I28204,);
DFFARX1 I_1457 (I1274159,I3563,I28221,I28377,);
nand I_1458 (I28385,I28377,I1274168);
not I_1459 (I28402,I28385);
nor I_1460 (I28201,I28247,I28402);
DFFARX1 I_1461 (I1274156,I3563,I28221,I28442,);
not I_1462 (I28450,I28442);
nor I_1463 (I28207,I28450,I28272);
nand I_1464 (I28195,I28450,I28385);
nand I_1465 (I28495,I1274177,I1274162);
and I_1466 (I28512,I28495,I1274156);
DFFARX1 I_1467 (I28512,I3563,I28221,I28538,);
nor I_1468 (I28546,I28538,I28247);
DFFARX1 I_1469 (I28546,I3563,I28221,I28189,);
not I_1470 (I28577,I28538);
nor I_1471 (I28594,I1274153,I1274162);
not I_1472 (I28611,I28594);
nor I_1473 (I28628,I28385,I28611);
nor I_1474 (I28645,I28577,I28628);
DFFARX1 I_1475 (I28645,I3563,I28221,I28210,);
nor I_1476 (I28676,I28538,I28611);
nor I_1477 (I28198,I28402,I28676);
nor I_1478 (I28192,I28538,I28594);
not I_1479 (I28748,I3570);
DFFARX1 I_1480 (I1165003,I3563,I28748,I28774,);
DFFARX1 I_1481 (I28774,I3563,I28748,I28791,);
not I_1482 (I28799,I28791);
nand I_1483 (I28816,I1164991,I1164982);
and I_1484 (I28833,I28816,I1164979);
DFFARX1 I_1485 (I28833,I3563,I28748,I28859,);
DFFARX1 I_1486 (I28859,I3563,I28748,I28740,);
DFFARX1 I_1487 (I28859,I3563,I28748,I28731,);
DFFARX1 I_1488 (I1164985,I3563,I28748,I28904,);
nand I_1489 (I28912,I28904,I1164997);
not I_1490 (I28929,I28912);
nor I_1491 (I28728,I28774,I28929);
DFFARX1 I_1492 (I1164994,I3563,I28748,I28969,);
not I_1493 (I28977,I28969);
nor I_1494 (I28734,I28977,I28799);
nand I_1495 (I28722,I28977,I28912);
nand I_1496 (I29022,I1164988,I1164982);
and I_1497 (I29039,I29022,I1165000);
DFFARX1 I_1498 (I29039,I3563,I28748,I29065,);
nor I_1499 (I29073,I29065,I28774);
DFFARX1 I_1500 (I29073,I3563,I28748,I28716,);
not I_1501 (I29104,I29065);
nor I_1502 (I29121,I1164979,I1164982);
not I_1503 (I29138,I29121);
nor I_1504 (I29155,I28912,I29138);
nor I_1505 (I29172,I29104,I29155);
DFFARX1 I_1506 (I29172,I3563,I28748,I28737,);
nor I_1507 (I29203,I29065,I29138);
nor I_1508 (I28725,I28929,I29203);
nor I_1509 (I28719,I29065,I29121);
not I_1510 (I29275,I3570);
DFFARX1 I_1511 (I903817,I3563,I29275,I29301,);
DFFARX1 I_1512 (I29301,I3563,I29275,I29318,);
not I_1513 (I29326,I29318);
nand I_1514 (I29343,I903808,I903829);
and I_1515 (I29360,I29343,I903811);
DFFARX1 I_1516 (I29360,I3563,I29275,I29386,);
DFFARX1 I_1517 (I29386,I3563,I29275,I29267,);
DFFARX1 I_1518 (I29386,I3563,I29275,I29258,);
DFFARX1 I_1519 (I903811,I3563,I29275,I29431,);
nand I_1520 (I29439,I29431,I903826);
not I_1521 (I29456,I29439);
nor I_1522 (I29255,I29301,I29456);
DFFARX1 I_1523 (I903820,I3563,I29275,I29496,);
not I_1524 (I29504,I29496);
nor I_1525 (I29261,I29504,I29326);
nand I_1526 (I29249,I29504,I29439);
nand I_1527 (I29549,I903814,I903823);
and I_1528 (I29566,I29549,I903808);
DFFARX1 I_1529 (I29566,I3563,I29275,I29592,);
nor I_1530 (I29600,I29592,I29301);
DFFARX1 I_1531 (I29600,I3563,I29275,I29243,);
not I_1532 (I29631,I29592);
nor I_1533 (I29648,I903814,I903823);
not I_1534 (I29665,I29648);
nor I_1535 (I29682,I29439,I29665);
nor I_1536 (I29699,I29631,I29682);
DFFARX1 I_1537 (I29699,I3563,I29275,I29264,);
nor I_1538 (I29730,I29592,I29665);
nor I_1539 (I29252,I29456,I29730);
nor I_1540 (I29246,I29592,I29648);
not I_1541 (I29802,I3570);
DFFARX1 I_1542 (I302256,I3563,I29802,I29828,);
DFFARX1 I_1543 (I29828,I3563,I29802,I29845,);
not I_1544 (I29853,I29845);
nand I_1545 (I29870,I302253,I302247);
and I_1546 (I29887,I29870,I302241);
DFFARX1 I_1547 (I29887,I3563,I29802,I29913,);
DFFARX1 I_1548 (I29913,I3563,I29802,I29794,);
DFFARX1 I_1549 (I29913,I3563,I29802,I29785,);
DFFARX1 I_1550 (I302229,I3563,I29802,I29958,);
nand I_1551 (I29966,I29958,I302238);
not I_1552 (I29983,I29966);
nor I_1553 (I29782,I29828,I29983);
DFFARX1 I_1554 (I302235,I3563,I29802,I30023,);
not I_1555 (I30031,I30023);
nor I_1556 (I29788,I30031,I29853);
nand I_1557 (I29776,I30031,I29966);
nand I_1558 (I30076,I302232,I302250);
and I_1559 (I30093,I30076,I302229);
DFFARX1 I_1560 (I30093,I3563,I29802,I30119,);
nor I_1561 (I30127,I30119,I29828);
DFFARX1 I_1562 (I30127,I3563,I29802,I29770,);
not I_1563 (I30158,I30119);
nor I_1564 (I30175,I302244,I302250);
not I_1565 (I30192,I30175);
nor I_1566 (I30209,I29966,I30192);
nor I_1567 (I30226,I30158,I30209);
DFFARX1 I_1568 (I30226,I3563,I29802,I29791,);
nor I_1569 (I30257,I30119,I30192);
nor I_1570 (I29779,I29983,I30257);
nor I_1571 (I29773,I30119,I30175);
not I_1572 (I30329,I3570);
DFFARX1 I_1573 (I523586,I3563,I30329,I30355,);
DFFARX1 I_1574 (I30355,I3563,I30329,I30372,);
not I_1575 (I30380,I30372);
nand I_1576 (I30397,I523586,I523589);
and I_1577 (I30414,I30397,I523610);
DFFARX1 I_1578 (I30414,I3563,I30329,I30440,);
DFFARX1 I_1579 (I30440,I3563,I30329,I30321,);
DFFARX1 I_1580 (I30440,I3563,I30329,I30312,);
DFFARX1 I_1581 (I523598,I3563,I30329,I30485,);
nand I_1582 (I30493,I30485,I523601);
not I_1583 (I30510,I30493);
nor I_1584 (I30309,I30355,I30510);
DFFARX1 I_1585 (I523607,I3563,I30329,I30550,);
not I_1586 (I30558,I30550);
nor I_1587 (I30315,I30558,I30380);
nand I_1588 (I30303,I30558,I30493);
nand I_1589 (I30603,I523604,I523592);
and I_1590 (I30620,I30603,I523595);
DFFARX1 I_1591 (I30620,I3563,I30329,I30646,);
nor I_1592 (I30654,I30646,I30355);
DFFARX1 I_1593 (I30654,I3563,I30329,I30297,);
not I_1594 (I30685,I30646);
nor I_1595 (I30702,I523613,I523592);
not I_1596 (I30719,I30702);
nor I_1597 (I30736,I30493,I30719);
nor I_1598 (I30753,I30685,I30736);
DFFARX1 I_1599 (I30753,I3563,I30329,I30318,);
nor I_1600 (I30784,I30646,I30719);
nor I_1601 (I30306,I30510,I30784);
nor I_1602 (I30300,I30646,I30702);
not I_1603 (I30856,I3570);
DFFARX1 I_1604 (I104080,I3563,I30856,I30882,);
DFFARX1 I_1605 (I30882,I3563,I30856,I30899,);
not I_1606 (I30907,I30899);
nand I_1607 (I30924,I104080,I104095);
and I_1608 (I30941,I30924,I104098);
DFFARX1 I_1609 (I30941,I3563,I30856,I30967,);
DFFARX1 I_1610 (I30967,I3563,I30856,I30848,);
DFFARX1 I_1611 (I30967,I3563,I30856,I30839,);
DFFARX1 I_1612 (I104092,I3563,I30856,I31012,);
nand I_1613 (I31020,I31012,I104101);
not I_1614 (I31037,I31020);
nor I_1615 (I30836,I30882,I31037);
DFFARX1 I_1616 (I104077,I3563,I30856,I31077,);
not I_1617 (I31085,I31077);
nor I_1618 (I30842,I31085,I30907);
nand I_1619 (I30830,I31085,I31020);
nand I_1620 (I31130,I104077,I104083);
and I_1621 (I31147,I31130,I104086);
DFFARX1 I_1622 (I31147,I3563,I30856,I31173,);
nor I_1623 (I31181,I31173,I30882);
DFFARX1 I_1624 (I31181,I3563,I30856,I30824,);
not I_1625 (I31212,I31173);
nor I_1626 (I31229,I104089,I104083);
not I_1627 (I31246,I31229);
nor I_1628 (I31263,I31020,I31246);
nor I_1629 (I31280,I31212,I31263);
DFFARX1 I_1630 (I31280,I3563,I30856,I30845,);
nor I_1631 (I31311,I31173,I31246);
nor I_1632 (I30833,I31037,I31311);
nor I_1633 (I30827,I31173,I31229);
not I_1634 (I31383,I3570);
DFFARX1 I_1635 (I380252,I3563,I31383,I31409,);
DFFARX1 I_1636 (I31409,I3563,I31383,I31426,);
not I_1637 (I31434,I31426);
nand I_1638 (I31451,I380249,I380243);
and I_1639 (I31468,I31451,I380237);
DFFARX1 I_1640 (I31468,I3563,I31383,I31494,);
DFFARX1 I_1641 (I31494,I3563,I31383,I31375,);
DFFARX1 I_1642 (I31494,I3563,I31383,I31366,);
DFFARX1 I_1643 (I380225,I3563,I31383,I31539,);
nand I_1644 (I31547,I31539,I380234);
not I_1645 (I31564,I31547);
nor I_1646 (I31363,I31409,I31564);
DFFARX1 I_1647 (I380231,I3563,I31383,I31604,);
not I_1648 (I31612,I31604);
nor I_1649 (I31369,I31612,I31434);
nand I_1650 (I31357,I31612,I31547);
nand I_1651 (I31657,I380228,I380246);
and I_1652 (I31674,I31657,I380225);
DFFARX1 I_1653 (I31674,I3563,I31383,I31700,);
nor I_1654 (I31708,I31700,I31409);
DFFARX1 I_1655 (I31708,I3563,I31383,I31351,);
not I_1656 (I31739,I31700);
nor I_1657 (I31756,I380240,I380246);
not I_1658 (I31773,I31756);
nor I_1659 (I31790,I31547,I31773);
nor I_1660 (I31807,I31739,I31790);
DFFARX1 I_1661 (I31807,I3563,I31383,I31372,);
nor I_1662 (I31838,I31700,I31773);
nor I_1663 (I31360,I31564,I31838);
nor I_1664 (I31354,I31700,I31756);
not I_1665 (I31910,I3570);
DFFARX1 I_1666 (I877994,I3563,I31910,I31936,);
DFFARX1 I_1667 (I31936,I3563,I31910,I31953,);
not I_1668 (I31961,I31953);
nand I_1669 (I31978,I877985,I878006);
and I_1670 (I31995,I31978,I877988);
DFFARX1 I_1671 (I31995,I3563,I31910,I32021,);
DFFARX1 I_1672 (I32021,I3563,I31910,I31902,);
DFFARX1 I_1673 (I32021,I3563,I31910,I31893,);
DFFARX1 I_1674 (I877988,I3563,I31910,I32066,);
nand I_1675 (I32074,I32066,I878003);
not I_1676 (I32091,I32074);
nor I_1677 (I31890,I31936,I32091);
DFFARX1 I_1678 (I877997,I3563,I31910,I32131,);
not I_1679 (I32139,I32131);
nor I_1680 (I31896,I32139,I31961);
nand I_1681 (I31884,I32139,I32074);
nand I_1682 (I32184,I877991,I878000);
and I_1683 (I32201,I32184,I877985);
DFFARX1 I_1684 (I32201,I3563,I31910,I32227,);
nor I_1685 (I32235,I32227,I31936);
DFFARX1 I_1686 (I32235,I3563,I31910,I31878,);
not I_1687 (I32266,I32227);
nor I_1688 (I32283,I877991,I878000);
not I_1689 (I32300,I32283);
nor I_1690 (I32317,I32074,I32300);
nor I_1691 (I32334,I32266,I32317);
DFFARX1 I_1692 (I32334,I3563,I31910,I31899,);
nor I_1693 (I32365,I32227,I32300);
nor I_1694 (I31887,I32091,I32365);
nor I_1695 (I31881,I32227,I32283);
not I_1696 (I32437,I3570);
DFFARX1 I_1697 (I280934,I3563,I32437,I32463,);
DFFARX1 I_1698 (I32463,I3563,I32437,I32480,);
not I_1699 (I32488,I32480);
nand I_1700 (I32505,I280952,I280937);
and I_1701 (I32522,I32505,I280940);
DFFARX1 I_1702 (I32522,I3563,I32437,I32548,);
DFFARX1 I_1703 (I32548,I3563,I32437,I32429,);
DFFARX1 I_1704 (I32548,I3563,I32437,I32420,);
DFFARX1 I_1705 (I280928,I3563,I32437,I32593,);
nand I_1706 (I32601,I32593,I280931);
not I_1707 (I32618,I32601);
nor I_1708 (I32417,I32463,I32618);
DFFARX1 I_1709 (I280943,I3563,I32437,I32658,);
not I_1710 (I32666,I32658);
nor I_1711 (I32423,I32666,I32488);
nand I_1712 (I32411,I32666,I32601);
nand I_1713 (I32711,I280949,I280946);
and I_1714 (I32728,I32711,I280931);
DFFARX1 I_1715 (I32728,I3563,I32437,I32754,);
nor I_1716 (I32762,I32754,I32463);
DFFARX1 I_1717 (I32762,I3563,I32437,I32405,);
not I_1718 (I32793,I32754);
nor I_1719 (I32810,I280928,I280946);
not I_1720 (I32827,I32810);
nor I_1721 (I32844,I32601,I32827);
nor I_1722 (I32861,I32793,I32844);
DFFARX1 I_1723 (I32861,I3563,I32437,I32426,);
nor I_1724 (I32892,I32754,I32827);
nor I_1725 (I32414,I32618,I32892);
nor I_1726 (I32408,I32754,I32810);
not I_1727 (I32964,I3570);
DFFARX1 I_1728 (I255349,I3563,I32964,I32990,);
DFFARX1 I_1729 (I32990,I3563,I32964,I33007,);
not I_1730 (I33015,I33007);
nand I_1731 (I33032,I255367,I255352);
and I_1732 (I33049,I33032,I255355);
DFFARX1 I_1733 (I33049,I3563,I32964,I33075,);
DFFARX1 I_1734 (I33075,I3563,I32964,I32956,);
DFFARX1 I_1735 (I33075,I3563,I32964,I32947,);
DFFARX1 I_1736 (I255343,I3563,I32964,I33120,);
nand I_1737 (I33128,I33120,I255346);
not I_1738 (I33145,I33128);
nor I_1739 (I32944,I32990,I33145);
DFFARX1 I_1740 (I255358,I3563,I32964,I33185,);
not I_1741 (I33193,I33185);
nor I_1742 (I32950,I33193,I33015);
nand I_1743 (I32938,I33193,I33128);
nand I_1744 (I33238,I255364,I255361);
and I_1745 (I33255,I33238,I255346);
DFFARX1 I_1746 (I33255,I3563,I32964,I33281,);
nor I_1747 (I33289,I33281,I32990);
DFFARX1 I_1748 (I33289,I3563,I32964,I32932,);
not I_1749 (I33320,I33281);
nor I_1750 (I33337,I255343,I255361);
not I_1751 (I33354,I33337);
nor I_1752 (I33371,I33128,I33354);
nor I_1753 (I33388,I33320,I33371);
DFFARX1 I_1754 (I33388,I3563,I32964,I32953,);
nor I_1755 (I33419,I33281,I33354);
nor I_1756 (I32941,I33145,I33419);
nor I_1757 (I32935,I33281,I33337);
not I_1758 (I33491,I3570);
DFFARX1 I_1759 (I942677,I3563,I33491,I33517,);
DFFARX1 I_1760 (I33517,I3563,I33491,I33534,);
not I_1761 (I33542,I33534);
nand I_1762 (I33559,I942653,I942680);
and I_1763 (I33576,I33559,I942665);
DFFARX1 I_1764 (I33576,I3563,I33491,I33602,);
DFFARX1 I_1765 (I33602,I3563,I33491,I33483,);
DFFARX1 I_1766 (I33602,I3563,I33491,I33474,);
DFFARX1 I_1767 (I942671,I3563,I33491,I33647,);
nand I_1768 (I33655,I33647,I942656);
not I_1769 (I33672,I33655);
nor I_1770 (I33471,I33517,I33672);
DFFARX1 I_1771 (I942674,I3563,I33491,I33712,);
not I_1772 (I33720,I33712);
nor I_1773 (I33477,I33720,I33542);
nand I_1774 (I33465,I33720,I33655);
nand I_1775 (I33765,I942659,I942662);
and I_1776 (I33782,I33765,I942653);
DFFARX1 I_1777 (I33782,I3563,I33491,I33808,);
nor I_1778 (I33816,I33808,I33517);
DFFARX1 I_1779 (I33816,I3563,I33491,I33459,);
not I_1780 (I33847,I33808);
nor I_1781 (I33864,I942668,I942662);
not I_1782 (I33881,I33864);
nor I_1783 (I33898,I33655,I33881);
nor I_1784 (I33915,I33847,I33898);
DFFARX1 I_1785 (I33915,I3563,I33491,I33480,);
nor I_1786 (I33946,I33808,I33881);
nor I_1787 (I33468,I33672,I33946);
nor I_1788 (I33462,I33808,I33864);
not I_1789 (I34018,I3570);
DFFARX1 I_1790 (I1317824,I3563,I34018,I34044,);
DFFARX1 I_1791 (I34044,I3563,I34018,I34061,);
not I_1792 (I34069,I34061);
nand I_1793 (I34086,I1317827,I1317821);
and I_1794 (I34103,I34086,I1317830);
DFFARX1 I_1795 (I34103,I3563,I34018,I34129,);
DFFARX1 I_1796 (I34129,I3563,I34018,I34010,);
DFFARX1 I_1797 (I34129,I3563,I34018,I34001,);
DFFARX1 I_1798 (I1317818,I3563,I34018,I34174,);
nand I_1799 (I34182,I34174,I1317833);
not I_1800 (I34199,I34182);
nor I_1801 (I33998,I34044,I34199);
DFFARX1 I_1802 (I1317809,I3563,I34018,I34239,);
not I_1803 (I34247,I34239);
nor I_1804 (I34004,I34247,I34069);
nand I_1805 (I33992,I34247,I34182);
nand I_1806 (I34292,I1317812,I1317812);
and I_1807 (I34309,I34292,I1317809);
DFFARX1 I_1808 (I34309,I3563,I34018,I34335,);
nor I_1809 (I34343,I34335,I34044);
DFFARX1 I_1810 (I34343,I3563,I34018,I33986,);
not I_1811 (I34374,I34335);
nor I_1812 (I34391,I1317815,I1317812);
not I_1813 (I34408,I34391);
nor I_1814 (I34425,I34182,I34408);
nor I_1815 (I34442,I34374,I34425);
DFFARX1 I_1816 (I34442,I3563,I34018,I34007,);
nor I_1817 (I34473,I34335,I34408);
nor I_1818 (I33995,I34199,I34473);
nor I_1819 (I33989,I34335,I34391);
not I_1820 (I34545,I3570);
DFFARX1 I_1821 (I519778,I3563,I34545,I34571,);
DFFARX1 I_1822 (I34571,I3563,I34545,I34588,);
not I_1823 (I34596,I34588);
nand I_1824 (I34613,I519778,I519781);
and I_1825 (I34630,I34613,I519802);
DFFARX1 I_1826 (I34630,I3563,I34545,I34656,);
DFFARX1 I_1827 (I34656,I3563,I34545,I34537,);
DFFARX1 I_1828 (I34656,I3563,I34545,I34528,);
DFFARX1 I_1829 (I519790,I3563,I34545,I34701,);
nand I_1830 (I34709,I34701,I519793);
not I_1831 (I34726,I34709);
nor I_1832 (I34525,I34571,I34726);
DFFARX1 I_1833 (I519799,I3563,I34545,I34766,);
not I_1834 (I34774,I34766);
nor I_1835 (I34531,I34774,I34596);
nand I_1836 (I34519,I34774,I34709);
nand I_1837 (I34819,I519796,I519784);
and I_1838 (I34836,I34819,I519787);
DFFARX1 I_1839 (I34836,I3563,I34545,I34862,);
nor I_1840 (I34870,I34862,I34571);
DFFARX1 I_1841 (I34870,I3563,I34545,I34513,);
not I_1842 (I34901,I34862);
nor I_1843 (I34918,I519805,I519784);
not I_1844 (I34935,I34918);
nor I_1845 (I34952,I34709,I34935);
nor I_1846 (I34969,I34901,I34952);
DFFARX1 I_1847 (I34969,I3563,I34545,I34534,);
nor I_1848 (I35000,I34862,I34935);
nor I_1849 (I34522,I34726,I35000);
nor I_1850 (I34516,I34862,I34918);
not I_1851 (I35072,I3570);
DFFARX1 I_1852 (I616812,I3563,I35072,I35098,);
DFFARX1 I_1853 (I35098,I3563,I35072,I35115,);
not I_1854 (I35123,I35115);
nand I_1855 (I35140,I616797,I616815);
and I_1856 (I35157,I35140,I616809);
DFFARX1 I_1857 (I35157,I3563,I35072,I35183,);
DFFARX1 I_1858 (I35183,I3563,I35072,I35064,);
DFFARX1 I_1859 (I35183,I3563,I35072,I35055,);
DFFARX1 I_1860 (I616806,I3563,I35072,I35228,);
nand I_1861 (I35236,I35228,I616797);
not I_1862 (I35253,I35236);
nor I_1863 (I35052,I35098,I35253);
DFFARX1 I_1864 (I616800,I3563,I35072,I35293,);
not I_1865 (I35301,I35293);
nor I_1866 (I35058,I35301,I35123);
nand I_1867 (I35046,I35301,I35236);
nand I_1868 (I35346,I616821,I616803);
and I_1869 (I35363,I35346,I616818);
DFFARX1 I_1870 (I35363,I3563,I35072,I35389,);
nor I_1871 (I35397,I35389,I35098);
DFFARX1 I_1872 (I35397,I3563,I35072,I35040,);
not I_1873 (I35428,I35389);
nor I_1874 (I35445,I616800,I616803);
not I_1875 (I35462,I35445);
nor I_1876 (I35479,I35236,I35462);
nor I_1877 (I35496,I35428,I35479);
DFFARX1 I_1878 (I35496,I3563,I35072,I35061,);
nor I_1879 (I35527,I35389,I35462);
nor I_1880 (I35049,I35253,I35527);
nor I_1881 (I35043,I35389,I35445);
not I_1882 (I35599,I3570);
DFFARX1 I_1883 (I1097955,I3563,I35599,I35625,);
DFFARX1 I_1884 (I35625,I3563,I35599,I35642,);
not I_1885 (I35650,I35642);
nand I_1886 (I35667,I1097943,I1097934);
and I_1887 (I35684,I35667,I1097931);
DFFARX1 I_1888 (I35684,I3563,I35599,I35710,);
DFFARX1 I_1889 (I35710,I3563,I35599,I35591,);
DFFARX1 I_1890 (I35710,I3563,I35599,I35582,);
DFFARX1 I_1891 (I1097937,I3563,I35599,I35755,);
nand I_1892 (I35763,I35755,I1097949);
not I_1893 (I35780,I35763);
nor I_1894 (I35579,I35625,I35780);
DFFARX1 I_1895 (I1097946,I3563,I35599,I35820,);
not I_1896 (I35828,I35820);
nor I_1897 (I35585,I35828,I35650);
nand I_1898 (I35573,I35828,I35763);
nand I_1899 (I35873,I1097940,I1097934);
and I_1900 (I35890,I35873,I1097952);
DFFARX1 I_1901 (I35890,I3563,I35599,I35916,);
nor I_1902 (I35924,I35916,I35625);
DFFARX1 I_1903 (I35924,I3563,I35599,I35567,);
not I_1904 (I35955,I35916);
nor I_1905 (I35972,I1097931,I1097934);
not I_1906 (I35989,I35972);
nor I_1907 (I36006,I35763,I35989);
nor I_1908 (I36023,I35955,I36006);
DFFARX1 I_1909 (I36023,I3563,I35599,I35588,);
nor I_1910 (I36054,I35916,I35989);
nor I_1911 (I35576,I35780,I36054);
nor I_1912 (I35570,I35916,I35972);
not I_1913 (I36126,I3570);
DFFARX1 I_1914 (I1283945,I3563,I36126,I36152,);
DFFARX1 I_1915 (I36152,I3563,I36126,I36169,);
not I_1916 (I36177,I36169);
nand I_1917 (I36194,I1283963,I1283957);
and I_1918 (I36211,I36194,I1283966);
DFFARX1 I_1919 (I36211,I3563,I36126,I36237,);
DFFARX1 I_1920 (I36237,I3563,I36126,I36118,);
DFFARX1 I_1921 (I36237,I3563,I36126,I36109,);
DFFARX1 I_1922 (I1283951,I3563,I36126,I36282,);
nand I_1923 (I36290,I36282,I1283960);
not I_1924 (I36307,I36290);
nor I_1925 (I36106,I36152,I36307);
DFFARX1 I_1926 (I1283948,I3563,I36126,I36347,);
not I_1927 (I36355,I36347);
nor I_1928 (I36112,I36355,I36177);
nand I_1929 (I36100,I36355,I36290);
nand I_1930 (I36400,I1283969,I1283954);
and I_1931 (I36417,I36400,I1283948);
DFFARX1 I_1932 (I36417,I3563,I36126,I36443,);
nor I_1933 (I36451,I36443,I36152);
DFFARX1 I_1934 (I36451,I3563,I36126,I36094,);
not I_1935 (I36482,I36443);
nor I_1936 (I36499,I1283945,I1283954);
not I_1937 (I36516,I36499);
nor I_1938 (I36533,I36290,I36516);
nor I_1939 (I36550,I36482,I36533);
DFFARX1 I_1940 (I36550,I3563,I36126,I36115,);
nor I_1941 (I36581,I36443,I36516);
nor I_1942 (I36103,I36307,I36581);
nor I_1943 (I36097,I36443,I36499);
not I_1944 (I36653,I3570);
DFFARX1 I_1945 (I475714,I3563,I36653,I36679,);
DFFARX1 I_1946 (I36679,I3563,I36653,I36696,);
not I_1947 (I36704,I36696);
nand I_1948 (I36721,I475714,I475717);
and I_1949 (I36738,I36721,I475738);
DFFARX1 I_1950 (I36738,I3563,I36653,I36764,);
DFFARX1 I_1951 (I36764,I3563,I36653,I36645,);
DFFARX1 I_1952 (I36764,I3563,I36653,I36636,);
DFFARX1 I_1953 (I475726,I3563,I36653,I36809,);
nand I_1954 (I36817,I36809,I475729);
not I_1955 (I36834,I36817);
nor I_1956 (I36633,I36679,I36834);
DFFARX1 I_1957 (I475735,I3563,I36653,I36874,);
not I_1958 (I36882,I36874);
nor I_1959 (I36639,I36882,I36704);
nand I_1960 (I36627,I36882,I36817);
nand I_1961 (I36927,I475732,I475720);
and I_1962 (I36944,I36927,I475723);
DFFARX1 I_1963 (I36944,I3563,I36653,I36970,);
nor I_1964 (I36978,I36970,I36679);
DFFARX1 I_1965 (I36978,I3563,I36653,I36621,);
not I_1966 (I37009,I36970);
nor I_1967 (I37026,I475741,I475720);
not I_1968 (I37043,I37026);
nor I_1969 (I37060,I36817,I37043);
nor I_1970 (I37077,I37009,I37060);
DFFARX1 I_1971 (I37077,I3563,I36653,I36642,);
nor I_1972 (I37108,I36970,I37043);
nor I_1973 (I36630,I36834,I37108);
nor I_1974 (I36624,I36970,I37026);
not I_1975 (I37180,I3570);
DFFARX1 I_1976 (I203584,I3563,I37180,I37206,);
DFFARX1 I_1977 (I37206,I3563,I37180,I37223,);
not I_1978 (I37231,I37223);
nand I_1979 (I37248,I203602,I203587);
and I_1980 (I37265,I37248,I203590);
DFFARX1 I_1981 (I37265,I3563,I37180,I37291,);
DFFARX1 I_1982 (I37291,I3563,I37180,I37172,);
DFFARX1 I_1983 (I37291,I3563,I37180,I37163,);
DFFARX1 I_1984 (I203578,I3563,I37180,I37336,);
nand I_1985 (I37344,I37336,I203581);
not I_1986 (I37361,I37344);
nor I_1987 (I37160,I37206,I37361);
DFFARX1 I_1988 (I203593,I3563,I37180,I37401,);
not I_1989 (I37409,I37401);
nor I_1990 (I37166,I37409,I37231);
nand I_1991 (I37154,I37409,I37344);
nand I_1992 (I37454,I203599,I203596);
and I_1993 (I37471,I37454,I203581);
DFFARX1 I_1994 (I37471,I3563,I37180,I37497,);
nor I_1995 (I37505,I37497,I37206);
DFFARX1 I_1996 (I37505,I3563,I37180,I37148,);
not I_1997 (I37536,I37497);
nor I_1998 (I37553,I203578,I203596);
not I_1999 (I37570,I37553);
nor I_2000 (I37587,I37344,I37570);
nor I_2001 (I37604,I37536,I37587);
DFFARX1 I_2002 (I37604,I3563,I37180,I37169,);
nor I_2003 (I37635,I37497,I37570);
nor I_2004 (I37157,I37361,I37635);
nor I_2005 (I37151,I37497,I37553);
not I_2006 (I37707,I3570);
DFFARX1 I_2007 (I1351163,I3563,I37707,I37733,);
DFFARX1 I_2008 (I37733,I3563,I37707,I37750,);
not I_2009 (I37758,I37750);
nand I_2010 (I37775,I1351166,I1351172);
and I_2011 (I37792,I37775,I1351181);
DFFARX1 I_2012 (I37792,I3563,I37707,I37818,);
DFFARX1 I_2013 (I37818,I3563,I37707,I37699,);
DFFARX1 I_2014 (I37818,I3563,I37707,I37690,);
DFFARX1 I_2015 (I1351184,I3563,I37707,I37863,);
nand I_2016 (I37871,I37863,I1351175);
not I_2017 (I37888,I37871);
nor I_2018 (I37687,I37733,I37888);
DFFARX1 I_2019 (I1351163,I3563,I37707,I37928,);
not I_2020 (I37936,I37928);
nor I_2021 (I37693,I37936,I37758);
nand I_2022 (I37681,I37936,I37871);
nand I_2023 (I37981,I1351190,I1351169);
and I_2024 (I37998,I37981,I1351178);
DFFARX1 I_2025 (I37998,I3563,I37707,I38024,);
nor I_2026 (I38032,I38024,I37733);
DFFARX1 I_2027 (I38032,I3563,I37707,I37675,);
not I_2028 (I38063,I38024);
nor I_2029 (I38080,I1351187,I1351169);
not I_2030 (I38097,I38080);
nor I_2031 (I38114,I37871,I38097);
nor I_2032 (I38131,I38063,I38114);
DFFARX1 I_2033 (I38131,I3563,I37707,I37696,);
nor I_2034 (I38162,I38024,I38097);
nor I_2035 (I37684,I37888,I38162);
nor I_2036 (I37678,I38024,I38080);
not I_2037 (I38234,I3570);
DFFARX1 I_2038 (I509986,I3563,I38234,I38260,);
DFFARX1 I_2039 (I38260,I3563,I38234,I38277,);
not I_2040 (I38285,I38277);
nand I_2041 (I38302,I509986,I509989);
and I_2042 (I38319,I38302,I510010);
DFFARX1 I_2043 (I38319,I3563,I38234,I38345,);
DFFARX1 I_2044 (I38345,I3563,I38234,I38226,);
DFFARX1 I_2045 (I38345,I3563,I38234,I38217,);
DFFARX1 I_2046 (I509998,I3563,I38234,I38390,);
nand I_2047 (I38398,I38390,I510001);
not I_2048 (I38415,I38398);
nor I_2049 (I38214,I38260,I38415);
DFFARX1 I_2050 (I510007,I3563,I38234,I38455,);
not I_2051 (I38463,I38455);
nor I_2052 (I38220,I38463,I38285);
nand I_2053 (I38208,I38463,I38398);
nand I_2054 (I38508,I510004,I509992);
and I_2055 (I38525,I38508,I509995);
DFFARX1 I_2056 (I38525,I3563,I38234,I38551,);
nor I_2057 (I38559,I38551,I38260);
DFFARX1 I_2058 (I38559,I3563,I38234,I38202,);
not I_2059 (I38590,I38551);
nor I_2060 (I38607,I510013,I509992);
not I_2061 (I38624,I38607);
nor I_2062 (I38641,I38398,I38624);
nor I_2063 (I38658,I38590,I38641);
DFFARX1 I_2064 (I38658,I3563,I38234,I38223,);
nor I_2065 (I38689,I38551,I38624);
nor I_2066 (I38211,I38415,I38689);
nor I_2067 (I38205,I38551,I38607);
not I_2068 (I38761,I3570);
DFFARX1 I_2069 (I329133,I3563,I38761,I38787,);
DFFARX1 I_2070 (I38787,I3563,I38761,I38804,);
not I_2071 (I38812,I38804);
nand I_2072 (I38829,I329130,I329124);
and I_2073 (I38846,I38829,I329118);
DFFARX1 I_2074 (I38846,I3563,I38761,I38872,);
DFFARX1 I_2075 (I38872,I3563,I38761,I38753,);
DFFARX1 I_2076 (I38872,I3563,I38761,I38744,);
DFFARX1 I_2077 (I329106,I3563,I38761,I38917,);
nand I_2078 (I38925,I38917,I329115);
not I_2079 (I38942,I38925);
nor I_2080 (I38741,I38787,I38942);
DFFARX1 I_2081 (I329112,I3563,I38761,I38982,);
not I_2082 (I38990,I38982);
nor I_2083 (I38747,I38990,I38812);
nand I_2084 (I38735,I38990,I38925);
nand I_2085 (I39035,I329109,I329127);
and I_2086 (I39052,I39035,I329106);
DFFARX1 I_2087 (I39052,I3563,I38761,I39078,);
nor I_2088 (I39086,I39078,I38787);
DFFARX1 I_2089 (I39086,I3563,I38761,I38729,);
not I_2090 (I39117,I39078);
nor I_2091 (I39134,I329121,I329127);
not I_2092 (I39151,I39134);
nor I_2093 (I39168,I38925,I39151);
nor I_2094 (I39185,I39117,I39168);
DFFARX1 I_2095 (I39185,I3563,I38761,I38750,);
nor I_2096 (I39216,I39078,I39151);
nor I_2097 (I38738,I38942,I39216);
nor I_2098 (I38732,I39078,I39134);
not I_2099 (I39288,I3570);
DFFARX1 I_2100 (I876940,I3563,I39288,I39314,);
DFFARX1 I_2101 (I39314,I3563,I39288,I39331,);
not I_2102 (I39339,I39331);
nand I_2103 (I39356,I876931,I876952);
and I_2104 (I39373,I39356,I876934);
DFFARX1 I_2105 (I39373,I3563,I39288,I39399,);
DFFARX1 I_2106 (I39399,I3563,I39288,I39280,);
DFFARX1 I_2107 (I39399,I3563,I39288,I39271,);
DFFARX1 I_2108 (I876934,I3563,I39288,I39444,);
nand I_2109 (I39452,I39444,I876949);
not I_2110 (I39469,I39452);
nor I_2111 (I39268,I39314,I39469);
DFFARX1 I_2112 (I876943,I3563,I39288,I39509,);
not I_2113 (I39517,I39509);
nor I_2114 (I39274,I39517,I39339);
nand I_2115 (I39262,I39517,I39452);
nand I_2116 (I39562,I876937,I876946);
and I_2117 (I39579,I39562,I876931);
DFFARX1 I_2118 (I39579,I3563,I39288,I39605,);
nor I_2119 (I39613,I39605,I39314);
DFFARX1 I_2120 (I39613,I3563,I39288,I39256,);
not I_2121 (I39644,I39605);
nor I_2122 (I39661,I876937,I876946);
not I_2123 (I39678,I39661);
nor I_2124 (I39695,I39452,I39678);
nor I_2125 (I39712,I39644,I39695);
DFFARX1 I_2126 (I39712,I3563,I39288,I39277,);
nor I_2127 (I39743,I39605,I39678);
nor I_2128 (I39265,I39469,I39743);
nor I_2129 (I39259,I39605,I39661);
not I_2130 (I39815,I3570);
DFFARX1 I_2131 (I1084252,I3563,I39815,I39841,);
DFFARX1 I_2132 (I39841,I3563,I39815,I39858,);
not I_2133 (I39866,I39858);
nand I_2134 (I39883,I1084246,I1084267);
and I_2135 (I39900,I39883,I1084252);
DFFARX1 I_2136 (I39900,I3563,I39815,I39926,);
DFFARX1 I_2137 (I39926,I3563,I39815,I39807,);
DFFARX1 I_2138 (I39926,I3563,I39815,I39798,);
DFFARX1 I_2139 (I1084249,I3563,I39815,I39971,);
nand I_2140 (I39979,I39971,I1084258);
not I_2141 (I39996,I39979);
nor I_2142 (I39795,I39841,I39996);
DFFARX1 I_2143 (I1084246,I3563,I39815,I40036,);
not I_2144 (I40044,I40036);
nor I_2145 (I39801,I40044,I39866);
nand I_2146 (I39789,I40044,I39979);
nand I_2147 (I40089,I1084249,I1084264);
and I_2148 (I40106,I40089,I1084255);
DFFARX1 I_2149 (I40106,I3563,I39815,I40132,);
nor I_2150 (I40140,I40132,I39841);
DFFARX1 I_2151 (I40140,I3563,I39815,I39783,);
not I_2152 (I40171,I40132);
nor I_2153 (I40188,I1084261,I1084264);
not I_2154 (I40205,I40188);
nor I_2155 (I40222,I39979,I40205);
nor I_2156 (I40239,I40171,I40222);
DFFARX1 I_2157 (I40239,I3563,I39815,I39804,);
nor I_2158 (I40270,I40132,I40205);
nor I_2159 (I39792,I39996,I40270);
nor I_2160 (I39786,I40132,I40188);
not I_2161 (I40342,I3570);
DFFARX1 I_2162 (I1162691,I3563,I40342,I40368,);
DFFARX1 I_2163 (I40368,I3563,I40342,I40385,);
not I_2164 (I40393,I40385);
nand I_2165 (I40410,I1162679,I1162670);
and I_2166 (I40427,I40410,I1162667);
DFFARX1 I_2167 (I40427,I3563,I40342,I40453,);
DFFARX1 I_2168 (I40453,I3563,I40342,I40334,);
DFFARX1 I_2169 (I40453,I3563,I40342,I40325,);
DFFARX1 I_2170 (I1162673,I3563,I40342,I40498,);
nand I_2171 (I40506,I40498,I1162685);
not I_2172 (I40523,I40506);
nor I_2173 (I40322,I40368,I40523);
DFFARX1 I_2174 (I1162682,I3563,I40342,I40563,);
not I_2175 (I40571,I40563);
nor I_2176 (I40328,I40571,I40393);
nand I_2177 (I40316,I40571,I40506);
nand I_2178 (I40616,I1162676,I1162670);
and I_2179 (I40633,I40616,I1162688);
DFFARX1 I_2180 (I40633,I3563,I40342,I40659,);
nor I_2181 (I40667,I40659,I40368);
DFFARX1 I_2182 (I40667,I3563,I40342,I40310,);
not I_2183 (I40698,I40659);
nor I_2184 (I40715,I1162667,I1162670);
not I_2185 (I40732,I40715);
nor I_2186 (I40749,I40506,I40732);
nor I_2187 (I40766,I40698,I40749);
DFFARX1 I_2188 (I40766,I3563,I40342,I40331,);
nor I_2189 (I40797,I40659,I40732);
nor I_2190 (I40319,I40523,I40797);
nor I_2191 (I40313,I40659,I40715);
not I_2192 (I40869,I3570);
DFFARX1 I_2193 (I1232051,I3563,I40869,I40895,);
DFFARX1 I_2194 (I40895,I3563,I40869,I40912,);
not I_2195 (I40920,I40912);
nand I_2196 (I40937,I1232039,I1232030);
and I_2197 (I40954,I40937,I1232027);
DFFARX1 I_2198 (I40954,I3563,I40869,I40980,);
DFFARX1 I_2199 (I40980,I3563,I40869,I40861,);
DFFARX1 I_2200 (I40980,I3563,I40869,I40852,);
DFFARX1 I_2201 (I1232033,I3563,I40869,I41025,);
nand I_2202 (I41033,I41025,I1232045);
not I_2203 (I41050,I41033);
nor I_2204 (I40849,I40895,I41050);
DFFARX1 I_2205 (I1232042,I3563,I40869,I41090,);
not I_2206 (I41098,I41090);
nor I_2207 (I40855,I41098,I40920);
nand I_2208 (I40843,I41098,I41033);
nand I_2209 (I41143,I1232036,I1232030);
and I_2210 (I41160,I41143,I1232048);
DFFARX1 I_2211 (I41160,I3563,I40869,I41186,);
nor I_2212 (I41194,I41186,I40895);
DFFARX1 I_2213 (I41194,I3563,I40869,I40837,);
not I_2214 (I41225,I41186);
nor I_2215 (I41242,I1232027,I1232030);
not I_2216 (I41259,I41242);
nor I_2217 (I41276,I41033,I41259);
nor I_2218 (I41293,I41225,I41276);
DFFARX1 I_2219 (I41293,I3563,I40869,I40858,);
nor I_2220 (I41324,I41186,I41259);
nor I_2221 (I40846,I41050,I41324);
nor I_2222 (I40840,I41186,I41242);
not I_2223 (I41396,I3570);
DFFARX1 I_2224 (I387630,I3563,I41396,I41422,);
DFFARX1 I_2225 (I41422,I3563,I41396,I41439,);
not I_2226 (I41447,I41439);
nand I_2227 (I41464,I387627,I387621);
and I_2228 (I41481,I41464,I387615);
DFFARX1 I_2229 (I41481,I3563,I41396,I41507,);
DFFARX1 I_2230 (I41507,I3563,I41396,I41388,);
DFFARX1 I_2231 (I41507,I3563,I41396,I41379,);
DFFARX1 I_2232 (I387603,I3563,I41396,I41552,);
nand I_2233 (I41560,I41552,I387612);
not I_2234 (I41577,I41560);
nor I_2235 (I41376,I41422,I41577);
DFFARX1 I_2236 (I387609,I3563,I41396,I41617,);
not I_2237 (I41625,I41617);
nor I_2238 (I41382,I41625,I41447);
nand I_2239 (I41370,I41625,I41560);
nand I_2240 (I41670,I387606,I387624);
and I_2241 (I41687,I41670,I387603);
DFFARX1 I_2242 (I41687,I3563,I41396,I41713,);
nor I_2243 (I41721,I41713,I41422);
DFFARX1 I_2244 (I41721,I3563,I41396,I41364,);
not I_2245 (I41752,I41713);
nor I_2246 (I41769,I387618,I387624);
not I_2247 (I41786,I41769);
nor I_2248 (I41803,I41560,I41786);
nor I_2249 (I41820,I41752,I41803);
DFFARX1 I_2250 (I41820,I3563,I41396,I41385,);
nor I_2251 (I41851,I41713,I41786);
nor I_2252 (I41373,I41577,I41851);
nor I_2253 (I41367,I41713,I41769);
not I_2254 (I41923,I3570);
DFFARX1 I_2255 (I949783,I3563,I41923,I41949,);
DFFARX1 I_2256 (I41949,I3563,I41923,I41966,);
not I_2257 (I41974,I41966);
nand I_2258 (I41991,I949759,I949786);
and I_2259 (I42008,I41991,I949771);
DFFARX1 I_2260 (I42008,I3563,I41923,I42034,);
DFFARX1 I_2261 (I42034,I3563,I41923,I41915,);
DFFARX1 I_2262 (I42034,I3563,I41923,I41906,);
DFFARX1 I_2263 (I949777,I3563,I41923,I42079,);
nand I_2264 (I42087,I42079,I949762);
not I_2265 (I42104,I42087);
nor I_2266 (I41903,I41949,I42104);
DFFARX1 I_2267 (I949780,I3563,I41923,I42144,);
not I_2268 (I42152,I42144);
nor I_2269 (I41909,I42152,I41974);
nand I_2270 (I41897,I42152,I42087);
nand I_2271 (I42197,I949765,I949768);
and I_2272 (I42214,I42197,I949759);
DFFARX1 I_2273 (I42214,I3563,I41923,I42240,);
nor I_2274 (I42248,I42240,I41949);
DFFARX1 I_2275 (I42248,I3563,I41923,I41891,);
not I_2276 (I42279,I42240);
nor I_2277 (I42296,I949774,I949768);
not I_2278 (I42313,I42296);
nor I_2279 (I42330,I42087,I42313);
nor I_2280 (I42347,I42279,I42330);
DFFARX1 I_2281 (I42347,I3563,I41923,I41912,);
nor I_2282 (I42378,I42240,I42313);
nor I_2283 (I41900,I42104,I42378);
nor I_2284 (I41894,I42240,I42296);
not I_2285 (I42450,I3570);
DFFARX1 I_2286 (I362334,I3563,I42450,I42476,);
DFFARX1 I_2287 (I42476,I3563,I42450,I42493,);
not I_2288 (I42501,I42493);
nand I_2289 (I42518,I362331,I362325);
and I_2290 (I42535,I42518,I362319);
DFFARX1 I_2291 (I42535,I3563,I42450,I42561,);
DFFARX1 I_2292 (I42561,I3563,I42450,I42442,);
DFFARX1 I_2293 (I42561,I3563,I42450,I42433,);
DFFARX1 I_2294 (I362307,I3563,I42450,I42606,);
nand I_2295 (I42614,I42606,I362316);
not I_2296 (I42631,I42614);
nor I_2297 (I42430,I42476,I42631);
DFFARX1 I_2298 (I362313,I3563,I42450,I42671,);
not I_2299 (I42679,I42671);
nor I_2300 (I42436,I42679,I42501);
nand I_2301 (I42424,I42679,I42614);
nand I_2302 (I42724,I362310,I362328);
and I_2303 (I42741,I42724,I362307);
DFFARX1 I_2304 (I42741,I3563,I42450,I42767,);
nor I_2305 (I42775,I42767,I42476);
DFFARX1 I_2306 (I42775,I3563,I42450,I42418,);
not I_2307 (I42806,I42767);
nor I_2308 (I42823,I362322,I362328);
not I_2309 (I42840,I42823);
nor I_2310 (I42857,I42614,I42840);
nor I_2311 (I42874,I42806,I42857);
DFFARX1 I_2312 (I42874,I3563,I42450,I42439,);
nor I_2313 (I42905,I42767,I42840);
nor I_2314 (I42427,I42631,I42905);
nor I_2315 (I42421,I42767,I42823);
not I_2316 (I42977,I3570);
DFFARX1 I_2317 (I1117029,I3563,I42977,I43003,);
DFFARX1 I_2318 (I43003,I3563,I42977,I43020,);
not I_2319 (I43028,I43020);
nand I_2320 (I43045,I1117017,I1117008);
and I_2321 (I43062,I43045,I1117005);
DFFARX1 I_2322 (I43062,I3563,I42977,I43088,);
DFFARX1 I_2323 (I43088,I3563,I42977,I42969,);
DFFARX1 I_2324 (I43088,I3563,I42977,I42960,);
DFFARX1 I_2325 (I1117011,I3563,I42977,I43133,);
nand I_2326 (I43141,I43133,I1117023);
not I_2327 (I43158,I43141);
nor I_2328 (I42957,I43003,I43158);
DFFARX1 I_2329 (I1117020,I3563,I42977,I43198,);
not I_2330 (I43206,I43198);
nor I_2331 (I42963,I43206,I43028);
nand I_2332 (I42951,I43206,I43141);
nand I_2333 (I43251,I1117014,I1117008);
and I_2334 (I43268,I43251,I1117026);
DFFARX1 I_2335 (I43268,I3563,I42977,I43294,);
nor I_2336 (I43302,I43294,I43003);
DFFARX1 I_2337 (I43302,I3563,I42977,I42945,);
not I_2338 (I43333,I43294);
nor I_2339 (I43350,I1117005,I1117008);
not I_2340 (I43367,I43350);
nor I_2341 (I43384,I43141,I43367);
nor I_2342 (I43401,I43333,I43384);
DFFARX1 I_2343 (I43401,I3563,I42977,I42966,);
nor I_2344 (I43432,I43294,I43367);
nor I_2345 (I42954,I43158,I43432);
nor I_2346 (I42948,I43294,I43350);
not I_2347 (I43504,I3570);
DFFARX1 I_2348 (I1192747,I3563,I43504,I43530,);
DFFARX1 I_2349 (I43530,I3563,I43504,I43547,);
not I_2350 (I43555,I43547);
nand I_2351 (I43572,I1192735,I1192726);
and I_2352 (I43589,I43572,I1192723);
DFFARX1 I_2353 (I43589,I3563,I43504,I43615,);
DFFARX1 I_2354 (I43615,I3563,I43504,I43496,);
DFFARX1 I_2355 (I43615,I3563,I43504,I43487,);
DFFARX1 I_2356 (I1192729,I3563,I43504,I43660,);
nand I_2357 (I43668,I43660,I1192741);
not I_2358 (I43685,I43668);
nor I_2359 (I43484,I43530,I43685);
DFFARX1 I_2360 (I1192738,I3563,I43504,I43725,);
not I_2361 (I43733,I43725);
nor I_2362 (I43490,I43733,I43555);
nand I_2363 (I43478,I43733,I43668);
nand I_2364 (I43778,I1192732,I1192726);
and I_2365 (I43795,I43778,I1192744);
DFFARX1 I_2366 (I43795,I3563,I43504,I43821,);
nor I_2367 (I43829,I43821,I43530);
DFFARX1 I_2368 (I43829,I3563,I43504,I43472,);
not I_2369 (I43860,I43821);
nor I_2370 (I43877,I1192723,I1192726);
not I_2371 (I43894,I43877);
nor I_2372 (I43911,I43668,I43894);
nor I_2373 (I43928,I43860,I43911);
DFFARX1 I_2374 (I43928,I3563,I43504,I43493,);
nor I_2375 (I43959,I43821,I43894);
nor I_2376 (I43481,I43685,I43959);
nor I_2377 (I43475,I43821,I43877);
not I_2378 (I44031,I3570);
DFFARX1 I_2379 (I495842,I3563,I44031,I44057,);
DFFARX1 I_2380 (I44057,I3563,I44031,I44074,);
not I_2381 (I44082,I44074);
nand I_2382 (I44099,I495842,I495845);
and I_2383 (I44116,I44099,I495866);
DFFARX1 I_2384 (I44116,I3563,I44031,I44142,);
DFFARX1 I_2385 (I44142,I3563,I44031,I44023,);
DFFARX1 I_2386 (I44142,I3563,I44031,I44014,);
DFFARX1 I_2387 (I495854,I3563,I44031,I44187,);
nand I_2388 (I44195,I44187,I495857);
not I_2389 (I44212,I44195);
nor I_2390 (I44011,I44057,I44212);
DFFARX1 I_2391 (I495863,I3563,I44031,I44252,);
not I_2392 (I44260,I44252);
nor I_2393 (I44017,I44260,I44082);
nand I_2394 (I44005,I44260,I44195);
nand I_2395 (I44305,I495860,I495848);
and I_2396 (I44322,I44305,I495851);
DFFARX1 I_2397 (I44322,I3563,I44031,I44348,);
nor I_2398 (I44356,I44348,I44057);
DFFARX1 I_2399 (I44356,I3563,I44031,I43999,);
not I_2400 (I44387,I44348);
nor I_2401 (I44404,I495869,I495848);
not I_2402 (I44421,I44404);
nor I_2403 (I44438,I44195,I44421);
nor I_2404 (I44455,I44387,I44438);
DFFARX1 I_2405 (I44455,I3563,I44031,I44020,);
nor I_2406 (I44486,I44348,I44421);
nor I_2407 (I44008,I44212,I44486);
nor I_2408 (I44002,I44348,I44404);
not I_2409 (I44558,I3570);
DFFARX1 I_2410 (I421858,I3563,I44558,I44584,);
DFFARX1 I_2411 (I44584,I3563,I44558,I44601,);
not I_2412 (I44609,I44601);
nand I_2413 (I44626,I421858,I421861);
and I_2414 (I44643,I44626,I421882);
DFFARX1 I_2415 (I44643,I3563,I44558,I44669,);
DFFARX1 I_2416 (I44669,I3563,I44558,I44550,);
DFFARX1 I_2417 (I44669,I3563,I44558,I44541,);
DFFARX1 I_2418 (I421870,I3563,I44558,I44714,);
nand I_2419 (I44722,I44714,I421873);
not I_2420 (I44739,I44722);
nor I_2421 (I44538,I44584,I44739);
DFFARX1 I_2422 (I421879,I3563,I44558,I44779,);
not I_2423 (I44787,I44779);
nor I_2424 (I44544,I44787,I44609);
nand I_2425 (I44532,I44787,I44722);
nand I_2426 (I44832,I421876,I421864);
and I_2427 (I44849,I44832,I421867);
DFFARX1 I_2428 (I44849,I3563,I44558,I44875,);
nor I_2429 (I44883,I44875,I44584);
DFFARX1 I_2430 (I44883,I3563,I44558,I44526,);
not I_2431 (I44914,I44875);
nor I_2432 (I44931,I421885,I421864);
not I_2433 (I44948,I44931);
nor I_2434 (I44965,I44722,I44948);
nor I_2435 (I44982,I44914,I44965);
DFFARX1 I_2436 (I44982,I3563,I44558,I44547,);
nor I_2437 (I45013,I44875,I44948);
nor I_2438 (I44535,I44739,I45013);
nor I_2439 (I44529,I44875,I44931);
not I_2440 (I45085,I3570);
DFFARX1 I_2441 (I871143,I3563,I45085,I45111,);
DFFARX1 I_2442 (I45111,I3563,I45085,I45128,);
not I_2443 (I45136,I45128);
nand I_2444 (I45153,I871134,I871155);
and I_2445 (I45170,I45153,I871137);
DFFARX1 I_2446 (I45170,I3563,I45085,I45196,);
DFFARX1 I_2447 (I45196,I3563,I45085,I45077,);
DFFARX1 I_2448 (I45196,I3563,I45085,I45068,);
DFFARX1 I_2449 (I871137,I3563,I45085,I45241,);
nand I_2450 (I45249,I45241,I871152);
not I_2451 (I45266,I45249);
nor I_2452 (I45065,I45111,I45266);
DFFARX1 I_2453 (I871146,I3563,I45085,I45306,);
not I_2454 (I45314,I45306);
nor I_2455 (I45071,I45314,I45136);
nand I_2456 (I45059,I45314,I45249);
nand I_2457 (I45359,I871140,I871149);
and I_2458 (I45376,I45359,I871134);
DFFARX1 I_2459 (I45376,I3563,I45085,I45402,);
nor I_2460 (I45410,I45402,I45111);
DFFARX1 I_2461 (I45410,I3563,I45085,I45053,);
not I_2462 (I45441,I45402);
nor I_2463 (I45458,I871140,I871149);
not I_2464 (I45475,I45458);
nor I_2465 (I45492,I45249,I45475);
nor I_2466 (I45509,I45441,I45492);
DFFARX1 I_2467 (I45509,I3563,I45085,I45074,);
nor I_2468 (I45540,I45402,I45475);
nor I_2469 (I45062,I45266,I45540);
nor I_2470 (I45056,I45402,I45458);
not I_2471 (I45612,I3570);
DFFARX1 I_2472 (I829510,I3563,I45612,I45638,);
DFFARX1 I_2473 (I45638,I3563,I45612,I45655,);
not I_2474 (I45663,I45655);
nand I_2475 (I45680,I829501,I829522);
and I_2476 (I45697,I45680,I829504);
DFFARX1 I_2477 (I45697,I3563,I45612,I45723,);
DFFARX1 I_2478 (I45723,I3563,I45612,I45604,);
DFFARX1 I_2479 (I45723,I3563,I45612,I45595,);
DFFARX1 I_2480 (I829504,I3563,I45612,I45768,);
nand I_2481 (I45776,I45768,I829519);
not I_2482 (I45793,I45776);
nor I_2483 (I45592,I45638,I45793);
DFFARX1 I_2484 (I829513,I3563,I45612,I45833,);
not I_2485 (I45841,I45833);
nor I_2486 (I45598,I45841,I45663);
nand I_2487 (I45586,I45841,I45776);
nand I_2488 (I45886,I829507,I829516);
and I_2489 (I45903,I45886,I829501);
DFFARX1 I_2490 (I45903,I3563,I45612,I45929,);
nor I_2491 (I45937,I45929,I45638);
DFFARX1 I_2492 (I45937,I3563,I45612,I45580,);
not I_2493 (I45968,I45929);
nor I_2494 (I45985,I829507,I829516);
not I_2495 (I46002,I45985);
nor I_2496 (I46019,I45776,I46002);
nor I_2497 (I46036,I45968,I46019);
DFFARX1 I_2498 (I46036,I3563,I45612,I45601,);
nor I_2499 (I46067,I45929,I46002);
nor I_2500 (I45589,I45793,I46067);
nor I_2501 (I45583,I45929,I45985);
not I_2502 (I46139,I3570);
DFFARX1 I_2503 (I1111249,I3563,I46139,I46165,);
DFFARX1 I_2504 (I46165,I3563,I46139,I46182,);
not I_2505 (I46190,I46182);
nand I_2506 (I46207,I1111237,I1111228);
and I_2507 (I46224,I46207,I1111225);
DFFARX1 I_2508 (I46224,I3563,I46139,I46250,);
DFFARX1 I_2509 (I46250,I3563,I46139,I46131,);
DFFARX1 I_2510 (I46250,I3563,I46139,I46122,);
DFFARX1 I_2511 (I1111231,I3563,I46139,I46295,);
nand I_2512 (I46303,I46295,I1111243);
not I_2513 (I46320,I46303);
nor I_2514 (I46119,I46165,I46320);
DFFARX1 I_2515 (I1111240,I3563,I46139,I46360,);
not I_2516 (I46368,I46360);
nor I_2517 (I46125,I46368,I46190);
nand I_2518 (I46113,I46368,I46303);
nand I_2519 (I46413,I1111234,I1111228);
and I_2520 (I46430,I46413,I1111246);
DFFARX1 I_2521 (I46430,I3563,I46139,I46456,);
nor I_2522 (I46464,I46456,I46165);
DFFARX1 I_2523 (I46464,I3563,I46139,I46107,);
not I_2524 (I46495,I46456);
nor I_2525 (I46512,I1111225,I1111228);
not I_2526 (I46529,I46512);
nor I_2527 (I46546,I46303,I46529);
nor I_2528 (I46563,I46495,I46546);
DFFARX1 I_2529 (I46563,I3563,I46139,I46128,);
nor I_2530 (I46594,I46456,I46529);
nor I_2531 (I46116,I46320,I46594);
nor I_2532 (I46110,I46456,I46512);
not I_2533 (I46666,I3570);
DFFARX1 I_2534 (I594848,I3563,I46666,I46692,);
DFFARX1 I_2535 (I46692,I3563,I46666,I46709,);
not I_2536 (I46717,I46709);
nand I_2537 (I46734,I594833,I594851);
and I_2538 (I46751,I46734,I594845);
DFFARX1 I_2539 (I46751,I3563,I46666,I46777,);
DFFARX1 I_2540 (I46777,I3563,I46666,I46658,);
DFFARX1 I_2541 (I46777,I3563,I46666,I46649,);
DFFARX1 I_2542 (I594842,I3563,I46666,I46822,);
nand I_2543 (I46830,I46822,I594833);
not I_2544 (I46847,I46830);
nor I_2545 (I46646,I46692,I46847);
DFFARX1 I_2546 (I594836,I3563,I46666,I46887,);
not I_2547 (I46895,I46887);
nor I_2548 (I46652,I46895,I46717);
nand I_2549 (I46640,I46895,I46830);
nand I_2550 (I46940,I594857,I594839);
and I_2551 (I46957,I46940,I594854);
DFFARX1 I_2552 (I46957,I3563,I46666,I46983,);
nor I_2553 (I46991,I46983,I46692);
DFFARX1 I_2554 (I46991,I3563,I46666,I46634,);
not I_2555 (I47022,I46983);
nor I_2556 (I47039,I594836,I594839);
not I_2557 (I47056,I47039);
nor I_2558 (I47073,I46830,I47056);
nor I_2559 (I47090,I47022,I47073);
DFFARX1 I_2560 (I47090,I3563,I46666,I46655,);
nor I_2561 (I47121,I46983,I47056);
nor I_2562 (I46643,I46847,I47121);
nor I_2563 (I46637,I46983,I47039);
not I_2564 (I47193,I3570);
DFFARX1 I_2565 (I901709,I3563,I47193,I47219,);
DFFARX1 I_2566 (I47219,I3563,I47193,I47236,);
not I_2567 (I47244,I47236);
nand I_2568 (I47261,I901700,I901721);
and I_2569 (I47278,I47261,I901703);
DFFARX1 I_2570 (I47278,I3563,I47193,I47304,);
DFFARX1 I_2571 (I47304,I3563,I47193,I47185,);
DFFARX1 I_2572 (I47304,I3563,I47193,I47176,);
DFFARX1 I_2573 (I901703,I3563,I47193,I47349,);
nand I_2574 (I47357,I47349,I901718);
not I_2575 (I47374,I47357);
nor I_2576 (I47173,I47219,I47374);
DFFARX1 I_2577 (I901712,I3563,I47193,I47414,);
not I_2578 (I47422,I47414);
nor I_2579 (I47179,I47422,I47244);
nand I_2580 (I47167,I47422,I47357);
nand I_2581 (I47467,I901706,I901715);
and I_2582 (I47484,I47467,I901700);
DFFARX1 I_2583 (I47484,I3563,I47193,I47510,);
nor I_2584 (I47518,I47510,I47219);
DFFARX1 I_2585 (I47518,I3563,I47193,I47161,);
not I_2586 (I47549,I47510);
nor I_2587 (I47566,I901706,I901715);
not I_2588 (I47583,I47566);
nor I_2589 (I47600,I47357,I47583);
nor I_2590 (I47617,I47549,I47600);
DFFARX1 I_2591 (I47617,I3563,I47193,I47182,);
nor I_2592 (I47648,I47510,I47583);
nor I_2593 (I47170,I47374,I47648);
nor I_2594 (I47164,I47510,I47566);
not I_2595 (I47720,I3570);
DFFARX1 I_2596 (I962057,I3563,I47720,I47746,);
DFFARX1 I_2597 (I47746,I3563,I47720,I47763,);
not I_2598 (I47771,I47763);
nand I_2599 (I47788,I962033,I962060);
and I_2600 (I47805,I47788,I962045);
DFFARX1 I_2601 (I47805,I3563,I47720,I47831,);
DFFARX1 I_2602 (I47831,I3563,I47720,I47712,);
DFFARX1 I_2603 (I47831,I3563,I47720,I47703,);
DFFARX1 I_2604 (I962051,I3563,I47720,I47876,);
nand I_2605 (I47884,I47876,I962036);
not I_2606 (I47901,I47884);
nor I_2607 (I47700,I47746,I47901);
DFFARX1 I_2608 (I962054,I3563,I47720,I47941,);
not I_2609 (I47949,I47941);
nor I_2610 (I47706,I47949,I47771);
nand I_2611 (I47694,I47949,I47884);
nand I_2612 (I47994,I962039,I962042);
and I_2613 (I48011,I47994,I962033);
DFFARX1 I_2614 (I48011,I3563,I47720,I48037,);
nor I_2615 (I48045,I48037,I47746);
DFFARX1 I_2616 (I48045,I3563,I47720,I47688,);
not I_2617 (I48076,I48037);
nor I_2618 (I48093,I962048,I962042);
not I_2619 (I48110,I48093);
nor I_2620 (I48127,I47884,I48110);
nor I_2621 (I48144,I48076,I48127);
DFFARX1 I_2622 (I48144,I3563,I47720,I47709,);
nor I_2623 (I48175,I48037,I48110);
nor I_2624 (I47697,I47901,I48175);
nor I_2625 (I47691,I48037,I48093);
not I_2626 (I48247,I3570);
DFFARX1 I_2627 (I1309732,I3563,I48247,I48273,);
DFFARX1 I_2628 (I48273,I3563,I48247,I48290,);
not I_2629 (I48298,I48290);
nand I_2630 (I48315,I1309735,I1309729);
and I_2631 (I48332,I48315,I1309738);
DFFARX1 I_2632 (I48332,I3563,I48247,I48358,);
DFFARX1 I_2633 (I48358,I3563,I48247,I48239,);
DFFARX1 I_2634 (I48358,I3563,I48247,I48230,);
DFFARX1 I_2635 (I1309726,I3563,I48247,I48403,);
nand I_2636 (I48411,I48403,I1309741);
not I_2637 (I48428,I48411);
nor I_2638 (I48227,I48273,I48428);
DFFARX1 I_2639 (I1309717,I3563,I48247,I48468,);
not I_2640 (I48476,I48468);
nor I_2641 (I48233,I48476,I48298);
nand I_2642 (I48221,I48476,I48411);
nand I_2643 (I48521,I1309720,I1309720);
and I_2644 (I48538,I48521,I1309717);
DFFARX1 I_2645 (I48538,I3563,I48247,I48564,);
nor I_2646 (I48572,I48564,I48273);
DFFARX1 I_2647 (I48572,I3563,I48247,I48215,);
not I_2648 (I48603,I48564);
nor I_2649 (I48620,I1309723,I1309720);
not I_2650 (I48637,I48620);
nor I_2651 (I48654,I48411,I48637);
nor I_2652 (I48671,I48603,I48654);
DFFARX1 I_2653 (I48671,I3563,I48247,I48236,);
nor I_2654 (I48702,I48564,I48637);
nor I_2655 (I48224,I48428,I48702);
nor I_2656 (I48218,I48564,I48620);
not I_2657 (I48774,I3570);
DFFARX1 I_2658 (I831618,I3563,I48774,I48800,);
DFFARX1 I_2659 (I48800,I3563,I48774,I48817,);
not I_2660 (I48825,I48817);
nand I_2661 (I48842,I831609,I831630);
and I_2662 (I48859,I48842,I831612);
DFFARX1 I_2663 (I48859,I3563,I48774,I48885,);
DFFARX1 I_2664 (I48885,I3563,I48774,I48766,);
DFFARX1 I_2665 (I48885,I3563,I48774,I48757,);
DFFARX1 I_2666 (I831612,I3563,I48774,I48930,);
nand I_2667 (I48938,I48930,I831627);
not I_2668 (I48955,I48938);
nor I_2669 (I48754,I48800,I48955);
DFFARX1 I_2670 (I831621,I3563,I48774,I48995,);
not I_2671 (I49003,I48995);
nor I_2672 (I48760,I49003,I48825);
nand I_2673 (I48748,I49003,I48938);
nand I_2674 (I49048,I831615,I831624);
and I_2675 (I49065,I49048,I831609);
DFFARX1 I_2676 (I49065,I3563,I48774,I49091,);
nor I_2677 (I49099,I49091,I48800);
DFFARX1 I_2678 (I49099,I3563,I48774,I48742,);
not I_2679 (I49130,I49091);
nor I_2680 (I49147,I831615,I831624);
not I_2681 (I49164,I49147);
nor I_2682 (I49181,I48938,I49164);
nor I_2683 (I49198,I49130,I49181);
DFFARX1 I_2684 (I49198,I3563,I48774,I48763,);
nor I_2685 (I49229,I49091,I49164);
nor I_2686 (I48751,I48955,I49229);
nor I_2687 (I48745,I49091,I49147);
not I_2688 (I49301,I3570);
DFFARX1 I_2689 (I1249673,I3563,I49301,I49327,);
DFFARX1 I_2690 (I49327,I3563,I49301,I49344,);
not I_2691 (I49352,I49344);
nand I_2692 (I49369,I1249691,I1249685);
and I_2693 (I49386,I49369,I1249694);
DFFARX1 I_2694 (I49386,I3563,I49301,I49412,);
DFFARX1 I_2695 (I49412,I3563,I49301,I49293,);
DFFARX1 I_2696 (I49412,I3563,I49301,I49284,);
DFFARX1 I_2697 (I1249679,I3563,I49301,I49457,);
nand I_2698 (I49465,I49457,I1249688);
not I_2699 (I49482,I49465);
nor I_2700 (I49281,I49327,I49482);
DFFARX1 I_2701 (I1249676,I3563,I49301,I49522,);
not I_2702 (I49530,I49522);
nor I_2703 (I49287,I49530,I49352);
nand I_2704 (I49275,I49530,I49465);
nand I_2705 (I49575,I1249697,I1249682);
and I_2706 (I49592,I49575,I1249676);
DFFARX1 I_2707 (I49592,I3563,I49301,I49618,);
nor I_2708 (I49626,I49618,I49327);
DFFARX1 I_2709 (I49626,I3563,I49301,I49269,);
not I_2710 (I49657,I49618);
nor I_2711 (I49674,I1249673,I1249682);
not I_2712 (I49691,I49674);
nor I_2713 (I49708,I49465,I49691);
nor I_2714 (I49725,I49657,I49708);
DFFARX1 I_2715 (I49725,I3563,I49301,I49290,);
nor I_2716 (I49756,I49618,I49691);
nor I_2717 (I49278,I49482,I49756);
nor I_2718 (I49272,I49618,I49674);
not I_2719 (I49828,I3570);
DFFARX1 I_2720 (I1131479,I3563,I49828,I49854,);
DFFARX1 I_2721 (I49854,I3563,I49828,I49871,);
not I_2722 (I49879,I49871);
nand I_2723 (I49896,I1131467,I1131458);
and I_2724 (I49913,I49896,I1131455);
DFFARX1 I_2725 (I49913,I3563,I49828,I49939,);
DFFARX1 I_2726 (I49939,I3563,I49828,I49820,);
DFFARX1 I_2727 (I49939,I3563,I49828,I49811,);
DFFARX1 I_2728 (I1131461,I3563,I49828,I49984,);
nand I_2729 (I49992,I49984,I1131473);
not I_2730 (I50009,I49992);
nor I_2731 (I49808,I49854,I50009);
DFFARX1 I_2732 (I1131470,I3563,I49828,I50049,);
not I_2733 (I50057,I50049);
nor I_2734 (I49814,I50057,I49879);
nand I_2735 (I49802,I50057,I49992);
nand I_2736 (I50102,I1131464,I1131458);
and I_2737 (I50119,I50102,I1131476);
DFFARX1 I_2738 (I50119,I3563,I49828,I50145,);
nor I_2739 (I50153,I50145,I49854);
DFFARX1 I_2740 (I50153,I3563,I49828,I49796,);
not I_2741 (I50184,I50145);
nor I_2742 (I50201,I1131455,I1131458);
not I_2743 (I50218,I50201);
nor I_2744 (I50235,I49992,I50218);
nor I_2745 (I50252,I50184,I50235);
DFFARX1 I_2746 (I50252,I3563,I49828,I49817,);
nor I_2747 (I50283,I50145,I50218);
nor I_2748 (I49805,I50009,I50283);
nor I_2749 (I49799,I50145,I50201);
not I_2750 (I50355,I3570);
DFFARX1 I_2751 (I509442,I3563,I50355,I50381,);
DFFARX1 I_2752 (I50381,I3563,I50355,I50398,);
not I_2753 (I50406,I50398);
nand I_2754 (I50423,I509442,I509445);
and I_2755 (I50440,I50423,I509466);
DFFARX1 I_2756 (I50440,I3563,I50355,I50466,);
DFFARX1 I_2757 (I50466,I3563,I50355,I50347,);
DFFARX1 I_2758 (I50466,I3563,I50355,I50338,);
DFFARX1 I_2759 (I509454,I3563,I50355,I50511,);
nand I_2760 (I50519,I50511,I509457);
not I_2761 (I50536,I50519);
nor I_2762 (I50335,I50381,I50536);
DFFARX1 I_2763 (I509463,I3563,I50355,I50576,);
not I_2764 (I50584,I50576);
nor I_2765 (I50341,I50584,I50406);
nand I_2766 (I50329,I50584,I50519);
nand I_2767 (I50629,I509460,I509448);
and I_2768 (I50646,I50629,I509451);
DFFARX1 I_2769 (I50646,I3563,I50355,I50672,);
nor I_2770 (I50680,I50672,I50381);
DFFARX1 I_2771 (I50680,I3563,I50355,I50323,);
not I_2772 (I50711,I50672);
nor I_2773 (I50728,I509469,I509448);
not I_2774 (I50745,I50728);
nor I_2775 (I50762,I50519,I50745);
nor I_2776 (I50779,I50711,I50762);
DFFARX1 I_2777 (I50779,I3563,I50355,I50344,);
nor I_2778 (I50810,I50672,I50745);
nor I_2779 (I50332,I50536,I50810);
nor I_2780 (I50326,I50672,I50728);
not I_2781 (I50882,I3570);
DFFARX1 I_2782 (I1388053,I3563,I50882,I50908,);
DFFARX1 I_2783 (I50908,I3563,I50882,I50925,);
not I_2784 (I50933,I50925);
nand I_2785 (I50950,I1388056,I1388062);
and I_2786 (I50967,I50950,I1388071);
DFFARX1 I_2787 (I50967,I3563,I50882,I50993,);
DFFARX1 I_2788 (I50993,I3563,I50882,I50874,);
DFFARX1 I_2789 (I50993,I3563,I50882,I50865,);
DFFARX1 I_2790 (I1388074,I3563,I50882,I51038,);
nand I_2791 (I51046,I51038,I1388065);
not I_2792 (I51063,I51046);
nor I_2793 (I50862,I50908,I51063);
DFFARX1 I_2794 (I1388053,I3563,I50882,I51103,);
not I_2795 (I51111,I51103);
nor I_2796 (I50868,I51111,I50933);
nand I_2797 (I50856,I51111,I51046);
nand I_2798 (I51156,I1388080,I1388059);
and I_2799 (I51173,I51156,I1388068);
DFFARX1 I_2800 (I51173,I3563,I50882,I51199,);
nor I_2801 (I51207,I51199,I50908);
DFFARX1 I_2802 (I51207,I3563,I50882,I50850,);
not I_2803 (I51238,I51199);
nor I_2804 (I51255,I1388077,I1388059);
not I_2805 (I51272,I51255);
nor I_2806 (I51289,I51046,I51272);
nor I_2807 (I51306,I51238,I51289);
DFFARX1 I_2808 (I51306,I3563,I50882,I50871,);
nor I_2809 (I51337,I51199,I51272);
nor I_2810 (I50859,I51063,I51337);
nor I_2811 (I50853,I51199,I51255);
not I_2812 (I51409,I3570);
DFFARX1 I_2813 (I263679,I3563,I51409,I51435,);
DFFARX1 I_2814 (I51435,I3563,I51409,I51452,);
not I_2815 (I51460,I51452);
nand I_2816 (I51477,I263697,I263682);
and I_2817 (I51494,I51477,I263685);
DFFARX1 I_2818 (I51494,I3563,I51409,I51520,);
DFFARX1 I_2819 (I51520,I3563,I51409,I51401,);
DFFARX1 I_2820 (I51520,I3563,I51409,I51392,);
DFFARX1 I_2821 (I263673,I3563,I51409,I51565,);
nand I_2822 (I51573,I51565,I263676);
not I_2823 (I51590,I51573);
nor I_2824 (I51389,I51435,I51590);
DFFARX1 I_2825 (I263688,I3563,I51409,I51630,);
not I_2826 (I51638,I51630);
nor I_2827 (I51395,I51638,I51460);
nand I_2828 (I51383,I51638,I51573);
nand I_2829 (I51683,I263694,I263691);
and I_2830 (I51700,I51683,I263676);
DFFARX1 I_2831 (I51700,I3563,I51409,I51726,);
nor I_2832 (I51734,I51726,I51435);
DFFARX1 I_2833 (I51734,I3563,I51409,I51377,);
not I_2834 (I51765,I51726);
nor I_2835 (I51782,I263673,I263691);
not I_2836 (I51799,I51782);
nor I_2837 (I51816,I51573,I51799);
nor I_2838 (I51833,I51765,I51816);
DFFARX1 I_2839 (I51833,I3563,I51409,I51398,);
nor I_2840 (I51864,I51726,I51799);
nor I_2841 (I51386,I51590,I51864);
nor I_2842 (I51380,I51726,I51782);
not I_2843 (I51936,I3570);
DFFARX1 I_2844 (I773441,I3563,I51936,I51962,);
DFFARX1 I_2845 (I51962,I3563,I51936,I51979,);
not I_2846 (I51987,I51979);
nand I_2847 (I52004,I773456,I773459);
and I_2848 (I52021,I52004,I773438);
DFFARX1 I_2849 (I52021,I3563,I51936,I52047,);
DFFARX1 I_2850 (I52047,I3563,I51936,I51928,);
DFFARX1 I_2851 (I52047,I3563,I51936,I51919,);
DFFARX1 I_2852 (I773444,I3563,I51936,I52092,);
nand I_2853 (I52100,I52092,I773450);
not I_2854 (I52117,I52100);
nor I_2855 (I51916,I51962,I52117);
DFFARX1 I_2856 (I773438,I3563,I51936,I52157,);
not I_2857 (I52165,I52157);
nor I_2858 (I51922,I52165,I51987);
nand I_2859 (I51910,I52165,I52100);
nand I_2860 (I52210,I773453,I773435);
and I_2861 (I52227,I52210,I773447);
DFFARX1 I_2862 (I52227,I3563,I51936,I52253,);
nor I_2863 (I52261,I52253,I51962);
DFFARX1 I_2864 (I52261,I3563,I51936,I51904,);
not I_2865 (I52292,I52253);
nor I_2866 (I52309,I773435,I773435);
not I_2867 (I52326,I52309);
nor I_2868 (I52343,I52100,I52326);
nor I_2869 (I52360,I52292,I52343);
DFFARX1 I_2870 (I52360,I3563,I51936,I51925,);
nor I_2871 (I52391,I52253,I52326);
nor I_2872 (I51913,I52117,I52391);
nor I_2873 (I51907,I52253,I52309);
not I_2874 (I52463,I3570);
DFFARX1 I_2875 (I794249,I3563,I52463,I52489,);
DFFARX1 I_2876 (I52489,I3563,I52463,I52506,);
not I_2877 (I52514,I52506);
nand I_2878 (I52531,I794264,I794267);
and I_2879 (I52548,I52531,I794246);
DFFARX1 I_2880 (I52548,I3563,I52463,I52574,);
DFFARX1 I_2881 (I52574,I3563,I52463,I52455,);
DFFARX1 I_2882 (I52574,I3563,I52463,I52446,);
DFFARX1 I_2883 (I794252,I3563,I52463,I52619,);
nand I_2884 (I52627,I52619,I794258);
not I_2885 (I52644,I52627);
nor I_2886 (I52443,I52489,I52644);
DFFARX1 I_2887 (I794246,I3563,I52463,I52684,);
not I_2888 (I52692,I52684);
nor I_2889 (I52449,I52692,I52514);
nand I_2890 (I52437,I52692,I52627);
nand I_2891 (I52737,I794261,I794243);
and I_2892 (I52754,I52737,I794255);
DFFARX1 I_2893 (I52754,I3563,I52463,I52780,);
nor I_2894 (I52788,I52780,I52489);
DFFARX1 I_2895 (I52788,I3563,I52463,I52431,);
not I_2896 (I52819,I52780);
nor I_2897 (I52836,I794243,I794243);
not I_2898 (I52853,I52836);
nor I_2899 (I52870,I52627,I52853);
nor I_2900 (I52887,I52819,I52870);
DFFARX1 I_2901 (I52887,I3563,I52463,I52452,);
nor I_2902 (I52918,I52780,I52853);
nor I_2903 (I52440,I52644,I52918);
nor I_2904 (I52434,I52780,I52836);
not I_2905 (I52990,I3570);
DFFARX1 I_2906 (I452322,I3563,I52990,I53016,);
DFFARX1 I_2907 (I53016,I3563,I52990,I53033,);
not I_2908 (I53041,I53033);
nand I_2909 (I53058,I452322,I452325);
and I_2910 (I53075,I53058,I452346);
DFFARX1 I_2911 (I53075,I3563,I52990,I53101,);
DFFARX1 I_2912 (I53101,I3563,I52990,I52982,);
DFFARX1 I_2913 (I53101,I3563,I52990,I52973,);
DFFARX1 I_2914 (I452334,I3563,I52990,I53146,);
nand I_2915 (I53154,I53146,I452337);
not I_2916 (I53171,I53154);
nor I_2917 (I52970,I53016,I53171);
DFFARX1 I_2918 (I452343,I3563,I52990,I53211,);
not I_2919 (I53219,I53211);
nor I_2920 (I52976,I53219,I53041);
nand I_2921 (I52964,I53219,I53154);
nand I_2922 (I53264,I452340,I452328);
and I_2923 (I53281,I53264,I452331);
DFFARX1 I_2924 (I53281,I3563,I52990,I53307,);
nor I_2925 (I53315,I53307,I53016);
DFFARX1 I_2926 (I53315,I3563,I52990,I52958,);
not I_2927 (I53346,I53307);
nor I_2928 (I53363,I452349,I452328);
not I_2929 (I53380,I53363);
nor I_2930 (I53397,I53154,I53380);
nor I_2931 (I53414,I53346,I53397);
DFFARX1 I_2932 (I53414,I3563,I52990,I52979,);
nor I_2933 (I53445,I53307,I53380);
nor I_2934 (I52967,I53171,I53445);
nor I_2935 (I52961,I53307,I53363);
not I_2936 (I53517,I3570);
DFFARX1 I_2937 (I1281769,I3563,I53517,I53543,);
DFFARX1 I_2938 (I53543,I3563,I53517,I53560,);
not I_2939 (I53568,I53560);
nand I_2940 (I53585,I1281787,I1281781);
and I_2941 (I53602,I53585,I1281790);
DFFARX1 I_2942 (I53602,I3563,I53517,I53628,);
DFFARX1 I_2943 (I53628,I3563,I53517,I53509,);
DFFARX1 I_2944 (I53628,I3563,I53517,I53500,);
DFFARX1 I_2945 (I1281775,I3563,I53517,I53673,);
nand I_2946 (I53681,I53673,I1281784);
not I_2947 (I53698,I53681);
nor I_2948 (I53497,I53543,I53698);
DFFARX1 I_2949 (I1281772,I3563,I53517,I53738,);
not I_2950 (I53746,I53738);
nor I_2951 (I53503,I53746,I53568);
nand I_2952 (I53491,I53746,I53681);
nand I_2953 (I53791,I1281793,I1281778);
and I_2954 (I53808,I53791,I1281772);
DFFARX1 I_2955 (I53808,I3563,I53517,I53834,);
nor I_2956 (I53842,I53834,I53543);
DFFARX1 I_2957 (I53842,I3563,I53517,I53485,);
not I_2958 (I53873,I53834);
nor I_2959 (I53890,I1281769,I1281778);
not I_2960 (I53907,I53890);
nor I_2961 (I53924,I53681,I53907);
nor I_2962 (I53941,I53873,I53924);
DFFARX1 I_2963 (I53941,I3563,I53517,I53506,);
nor I_2964 (I53972,I53834,I53907);
nor I_2965 (I53494,I53698,I53972);
nor I_2966 (I53488,I53834,I53890);
not I_2967 (I54044,I3570);
DFFARX1 I_2968 (I876413,I3563,I54044,I54070,);
DFFARX1 I_2969 (I54070,I3563,I54044,I54087,);
not I_2970 (I54095,I54087);
nand I_2971 (I54112,I876404,I876425);
and I_2972 (I54129,I54112,I876407);
DFFARX1 I_2973 (I54129,I3563,I54044,I54155,);
DFFARX1 I_2974 (I54155,I3563,I54044,I54036,);
DFFARX1 I_2975 (I54155,I3563,I54044,I54027,);
DFFARX1 I_2976 (I876407,I3563,I54044,I54200,);
nand I_2977 (I54208,I54200,I876422);
not I_2978 (I54225,I54208);
nor I_2979 (I54024,I54070,I54225);
DFFARX1 I_2980 (I876416,I3563,I54044,I54265,);
not I_2981 (I54273,I54265);
nor I_2982 (I54030,I54273,I54095);
nand I_2983 (I54018,I54273,I54208);
nand I_2984 (I54318,I876410,I876419);
and I_2985 (I54335,I54318,I876404);
DFFARX1 I_2986 (I54335,I3563,I54044,I54361,);
nor I_2987 (I54369,I54361,I54070);
DFFARX1 I_2988 (I54369,I3563,I54044,I54012,);
not I_2989 (I54400,I54361);
nor I_2990 (I54417,I876410,I876419);
not I_2991 (I54434,I54417);
nor I_2992 (I54451,I54208,I54434);
nor I_2993 (I54468,I54400,I54451);
DFFARX1 I_2994 (I54468,I3563,I54044,I54033,);
nor I_2995 (I54499,I54361,I54434);
nor I_2996 (I54021,I54225,I54499);
nor I_2997 (I54015,I54361,I54417);
not I_2998 (I54571,I3570);
DFFARX1 I_2999 (I836888,I3563,I54571,I54597,);
DFFARX1 I_3000 (I54597,I3563,I54571,I54614,);
not I_3001 (I54622,I54614);
nand I_3002 (I54639,I836879,I836900);
and I_3003 (I54656,I54639,I836882);
DFFARX1 I_3004 (I54656,I3563,I54571,I54682,);
DFFARX1 I_3005 (I54682,I3563,I54571,I54563,);
DFFARX1 I_3006 (I54682,I3563,I54571,I54554,);
DFFARX1 I_3007 (I836882,I3563,I54571,I54727,);
nand I_3008 (I54735,I54727,I836897);
not I_3009 (I54752,I54735);
nor I_3010 (I54551,I54597,I54752);
DFFARX1 I_3011 (I836891,I3563,I54571,I54792,);
not I_3012 (I54800,I54792);
nor I_3013 (I54557,I54800,I54622);
nand I_3014 (I54545,I54800,I54735);
nand I_3015 (I54845,I836885,I836894);
and I_3016 (I54862,I54845,I836879);
DFFARX1 I_3017 (I54862,I3563,I54571,I54888,);
nor I_3018 (I54896,I54888,I54597);
DFFARX1 I_3019 (I54896,I3563,I54571,I54539,);
not I_3020 (I54927,I54888);
nor I_3021 (I54944,I836885,I836894);
not I_3022 (I54961,I54944);
nor I_3023 (I54978,I54735,I54961);
nor I_3024 (I54995,I54927,I54978);
DFFARX1 I_3025 (I54995,I3563,I54571,I54560,);
nor I_3026 (I55026,I54888,I54961);
nor I_3027 (I54548,I54752,I55026);
nor I_3028 (I54542,I54888,I54944);
not I_3029 (I55098,I3570);
DFFARX1 I_3030 (I296459,I3563,I55098,I55124,);
DFFARX1 I_3031 (I55124,I3563,I55098,I55141,);
not I_3032 (I55149,I55141);
nand I_3033 (I55166,I296456,I296450);
and I_3034 (I55183,I55166,I296444);
DFFARX1 I_3035 (I55183,I3563,I55098,I55209,);
DFFARX1 I_3036 (I55209,I3563,I55098,I55090,);
DFFARX1 I_3037 (I55209,I3563,I55098,I55081,);
DFFARX1 I_3038 (I296432,I3563,I55098,I55254,);
nand I_3039 (I55262,I55254,I296441);
not I_3040 (I55279,I55262);
nor I_3041 (I55078,I55124,I55279);
DFFARX1 I_3042 (I296438,I3563,I55098,I55319,);
not I_3043 (I55327,I55319);
nor I_3044 (I55084,I55327,I55149);
nand I_3045 (I55072,I55327,I55262);
nand I_3046 (I55372,I296435,I296453);
and I_3047 (I55389,I55372,I296432);
DFFARX1 I_3048 (I55389,I3563,I55098,I55415,);
nor I_3049 (I55423,I55415,I55124);
DFFARX1 I_3050 (I55423,I3563,I55098,I55066,);
not I_3051 (I55454,I55415);
nor I_3052 (I55471,I296447,I296453);
not I_3053 (I55488,I55471);
nor I_3054 (I55505,I55262,I55488);
nor I_3055 (I55522,I55454,I55505);
DFFARX1 I_3056 (I55522,I3563,I55098,I55087,);
nor I_3057 (I55553,I55415,I55488);
nor I_3058 (I55075,I55279,I55553);
nor I_3059 (I55069,I55415,I55471);
not I_3060 (I55625,I3570);
DFFARX1 I_3061 (I634730,I3563,I55625,I55651,);
DFFARX1 I_3062 (I55651,I3563,I55625,I55668,);
not I_3063 (I55676,I55668);
nand I_3064 (I55693,I634715,I634733);
and I_3065 (I55710,I55693,I634727);
DFFARX1 I_3066 (I55710,I3563,I55625,I55736,);
DFFARX1 I_3067 (I55736,I3563,I55625,I55617,);
DFFARX1 I_3068 (I55736,I3563,I55625,I55608,);
DFFARX1 I_3069 (I634724,I3563,I55625,I55781,);
nand I_3070 (I55789,I55781,I634715);
not I_3071 (I55806,I55789);
nor I_3072 (I55605,I55651,I55806);
DFFARX1 I_3073 (I634718,I3563,I55625,I55846,);
not I_3074 (I55854,I55846);
nor I_3075 (I55611,I55854,I55676);
nand I_3076 (I55599,I55854,I55789);
nand I_3077 (I55899,I634739,I634721);
and I_3078 (I55916,I55899,I634736);
DFFARX1 I_3079 (I55916,I3563,I55625,I55942,);
nor I_3080 (I55950,I55942,I55651);
DFFARX1 I_3081 (I55950,I3563,I55625,I55593,);
not I_3082 (I55981,I55942);
nor I_3083 (I55998,I634718,I634721);
not I_3084 (I56015,I55998);
nor I_3085 (I56032,I55789,I56015);
nor I_3086 (I56049,I55981,I56032);
DFFARX1 I_3087 (I56049,I3563,I55625,I55614,);
nor I_3088 (I56080,I55942,I56015);
nor I_3089 (I55602,I55806,I56080);
nor I_3090 (I55596,I55942,I55998);
not I_3091 (I56152,I3570);
DFFARX1 I_3092 (I733559,I3563,I56152,I56178,);
DFFARX1 I_3093 (I56178,I3563,I56152,I56195,);
not I_3094 (I56203,I56195);
nand I_3095 (I56220,I733574,I733577);
and I_3096 (I56237,I56220,I733556);
DFFARX1 I_3097 (I56237,I3563,I56152,I56263,);
DFFARX1 I_3098 (I56263,I3563,I56152,I56144,);
DFFARX1 I_3099 (I56263,I3563,I56152,I56135,);
DFFARX1 I_3100 (I733562,I3563,I56152,I56308,);
nand I_3101 (I56316,I56308,I733568);
not I_3102 (I56333,I56316);
nor I_3103 (I56132,I56178,I56333);
DFFARX1 I_3104 (I733556,I3563,I56152,I56373,);
not I_3105 (I56381,I56373);
nor I_3106 (I56138,I56381,I56203);
nand I_3107 (I56126,I56381,I56316);
nand I_3108 (I56426,I733571,I733553);
and I_3109 (I56443,I56426,I733565);
DFFARX1 I_3110 (I56443,I3563,I56152,I56469,);
nor I_3111 (I56477,I56469,I56178);
DFFARX1 I_3112 (I56477,I3563,I56152,I56120,);
not I_3113 (I56508,I56469);
nor I_3114 (I56525,I733553,I733553);
not I_3115 (I56542,I56525);
nor I_3116 (I56559,I56316,I56542);
nor I_3117 (I56576,I56508,I56559);
DFFARX1 I_3118 (I56576,I3563,I56152,I56141,);
nor I_3119 (I56607,I56469,I56542);
nor I_3120 (I56129,I56333,I56607);
nor I_3121 (I56123,I56469,I56525);
not I_3122 (I56679,I3570);
DFFARX1 I_3123 (I1185811,I3563,I56679,I56705,);
DFFARX1 I_3124 (I56705,I3563,I56679,I56722,);
not I_3125 (I56730,I56722);
nand I_3126 (I56747,I1185799,I1185790);
and I_3127 (I56764,I56747,I1185787);
DFFARX1 I_3128 (I56764,I3563,I56679,I56790,);
DFFARX1 I_3129 (I56790,I3563,I56679,I56671,);
DFFARX1 I_3130 (I56790,I3563,I56679,I56662,);
DFFARX1 I_3131 (I1185793,I3563,I56679,I56835,);
nand I_3132 (I56843,I56835,I1185805);
not I_3133 (I56860,I56843);
nor I_3134 (I56659,I56705,I56860);
DFFARX1 I_3135 (I1185802,I3563,I56679,I56900,);
not I_3136 (I56908,I56900);
nor I_3137 (I56665,I56908,I56730);
nand I_3138 (I56653,I56908,I56843);
nand I_3139 (I56953,I1185796,I1185790);
and I_3140 (I56970,I56953,I1185808);
DFFARX1 I_3141 (I56970,I3563,I56679,I56996,);
nor I_3142 (I57004,I56996,I56705);
DFFARX1 I_3143 (I57004,I3563,I56679,I56647,);
not I_3144 (I57035,I56996);
nor I_3145 (I57052,I1185787,I1185790);
not I_3146 (I57069,I57052);
nor I_3147 (I57086,I56843,I57069);
nor I_3148 (I57103,I57035,I57086);
DFFARX1 I_3149 (I57103,I3563,I56679,I56668,);
nor I_3150 (I57134,I56996,I57069);
nor I_3151 (I56656,I56860,I57134);
nor I_3152 (I56650,I56996,I57052);
not I_3153 (I57206,I3570);
DFFARX1 I_3154 (I1212977,I3563,I57206,I57232,);
DFFARX1 I_3155 (I57232,I3563,I57206,I57249,);
not I_3156 (I57257,I57249);
nand I_3157 (I57274,I1212965,I1212956);
and I_3158 (I57291,I57274,I1212953);
DFFARX1 I_3159 (I57291,I3563,I57206,I57317,);
DFFARX1 I_3160 (I57317,I3563,I57206,I57198,);
DFFARX1 I_3161 (I57317,I3563,I57206,I57189,);
DFFARX1 I_3162 (I1212959,I3563,I57206,I57362,);
nand I_3163 (I57370,I57362,I1212971);
not I_3164 (I57387,I57370);
nor I_3165 (I57186,I57232,I57387);
DFFARX1 I_3166 (I1212968,I3563,I57206,I57427,);
not I_3167 (I57435,I57427);
nor I_3168 (I57192,I57435,I57257);
nand I_3169 (I57180,I57435,I57370);
nand I_3170 (I57480,I1212962,I1212956);
and I_3171 (I57497,I57480,I1212974);
DFFARX1 I_3172 (I57497,I3563,I57206,I57523,);
nor I_3173 (I57531,I57523,I57232);
DFFARX1 I_3174 (I57531,I3563,I57206,I57174,);
not I_3175 (I57562,I57523);
nor I_3176 (I57579,I1212953,I1212956);
not I_3177 (I57596,I57579);
nor I_3178 (I57613,I57370,I57596);
nor I_3179 (I57630,I57562,I57613);
DFFARX1 I_3180 (I57630,I3563,I57206,I57195,);
nor I_3181 (I57661,I57523,I57596);
nor I_3182 (I57183,I57387,I57661);
nor I_3183 (I57177,I57523,I57579);
not I_3184 (I57733,I3570);
DFFARX1 I_3185 (I1233207,I3563,I57733,I57759,);
DFFARX1 I_3186 (I57759,I3563,I57733,I57776,);
not I_3187 (I57784,I57776);
nand I_3188 (I57801,I1233195,I1233186);
and I_3189 (I57818,I57801,I1233183);
DFFARX1 I_3190 (I57818,I3563,I57733,I57844,);
DFFARX1 I_3191 (I57844,I3563,I57733,I57725,);
DFFARX1 I_3192 (I57844,I3563,I57733,I57716,);
DFFARX1 I_3193 (I1233189,I3563,I57733,I57889,);
nand I_3194 (I57897,I57889,I1233201);
not I_3195 (I57914,I57897);
nor I_3196 (I57713,I57759,I57914);
DFFARX1 I_3197 (I1233198,I3563,I57733,I57954,);
not I_3198 (I57962,I57954);
nor I_3199 (I57719,I57962,I57784);
nand I_3200 (I57707,I57962,I57897);
nand I_3201 (I58007,I1233192,I1233186);
and I_3202 (I58024,I58007,I1233204);
DFFARX1 I_3203 (I58024,I3563,I57733,I58050,);
nor I_3204 (I58058,I58050,I57759);
DFFARX1 I_3205 (I58058,I3563,I57733,I57701,);
not I_3206 (I58089,I58050);
nor I_3207 (I58106,I1233183,I1233186);
not I_3208 (I58123,I58106);
nor I_3209 (I58140,I57897,I58123);
nor I_3210 (I58157,I58089,I58140);
DFFARX1 I_3211 (I58157,I3563,I57733,I57722,);
nor I_3212 (I58188,I58050,I58123);
nor I_3213 (I57710,I57914,I58188);
nor I_3214 (I57704,I58050,I58106);
not I_3215 (I58260,I3570);
DFFARX1 I_3216 (I353902,I3563,I58260,I58286,);
not I_3217 (I58294,I58286);
nand I_3218 (I58311,I353884,I353899);
and I_3219 (I58328,I58311,I353875);
DFFARX1 I_3220 (I58328,I3563,I58260,I58354,);
DFFARX1 I_3221 (I353878,I3563,I58260,I58371,);
and I_3222 (I58379,I58371,I353893);
nor I_3223 (I58396,I58354,I58379);
DFFARX1 I_3224 (I58396,I3563,I58260,I58228,);
nand I_3225 (I58427,I58371,I353893);
nand I_3226 (I58444,I58294,I58427);
not I_3227 (I58240,I58444);
DFFARX1 I_3228 (I353896,I3563,I58260,I58484,);
DFFARX1 I_3229 (I58484,I3563,I58260,I58249,);
nand I_3230 (I58506,I353875,I353887);
and I_3231 (I58523,I58506,I353881);
DFFARX1 I_3232 (I58523,I3563,I58260,I58549,);
DFFARX1 I_3233 (I58549,I3563,I58260,I58566,);
not I_3234 (I58252,I58566);
not I_3235 (I58588,I58549);
nand I_3236 (I58237,I58588,I58427);
nor I_3237 (I58619,I353890,I353887);
not I_3238 (I58636,I58619);
nor I_3239 (I58653,I58588,I58636);
nor I_3240 (I58670,I58294,I58653);
DFFARX1 I_3241 (I58670,I3563,I58260,I58246,);
nor I_3242 (I58701,I58354,I58636);
nor I_3243 (I58234,I58549,I58701);
nor I_3244 (I58243,I58484,I58619);
nor I_3245 (I58231,I58354,I58619);
not I_3246 (I58787,I3570);
DFFARX1 I_3247 (I217870,I3563,I58787,I58813,);
not I_3248 (I58821,I58813);
nand I_3249 (I58838,I217864,I217858);
and I_3250 (I58855,I58838,I217879);
DFFARX1 I_3251 (I58855,I3563,I58787,I58881,);
DFFARX1 I_3252 (I217876,I3563,I58787,I58898,);
and I_3253 (I58906,I58898,I217873);
nor I_3254 (I58923,I58881,I58906);
DFFARX1 I_3255 (I58923,I3563,I58787,I58755,);
nand I_3256 (I58954,I58898,I217873);
nand I_3257 (I58971,I58821,I58954);
not I_3258 (I58767,I58971);
DFFARX1 I_3259 (I217858,I3563,I58787,I59011,);
DFFARX1 I_3260 (I59011,I3563,I58787,I58776,);
nand I_3261 (I59033,I217861,I217861);
and I_3262 (I59050,I59033,I217882);
DFFARX1 I_3263 (I59050,I3563,I58787,I59076,);
DFFARX1 I_3264 (I59076,I3563,I58787,I59093,);
not I_3265 (I58779,I59093);
not I_3266 (I59115,I59076);
nand I_3267 (I58764,I59115,I58954);
nor I_3268 (I59146,I217867,I217861);
not I_3269 (I59163,I59146);
nor I_3270 (I59180,I59115,I59163);
nor I_3271 (I59197,I58821,I59180);
DFFARX1 I_3272 (I59197,I3563,I58787,I58773,);
nor I_3273 (I59228,I58881,I59163);
nor I_3274 (I58761,I59076,I59228);
nor I_3275 (I58770,I59011,I59146);
nor I_3276 (I58758,I58881,I59146);
not I_3277 (I59314,I3570);
DFFARX1 I_3278 (I1380925,I3563,I59314,I59340,);
not I_3279 (I59348,I59340);
nand I_3280 (I59365,I1380919,I1380940);
and I_3281 (I59382,I59365,I1380916);
DFFARX1 I_3282 (I59382,I3563,I59314,I59408,);
DFFARX1 I_3283 (I1380937,I3563,I59314,I59425,);
and I_3284 (I59433,I59425,I1380934);
nor I_3285 (I59450,I59408,I59433);
DFFARX1 I_3286 (I59450,I3563,I59314,I59282,);
nand I_3287 (I59481,I59425,I1380934);
nand I_3288 (I59498,I59348,I59481);
not I_3289 (I59294,I59498);
DFFARX1 I_3290 (I1380922,I3563,I59314,I59538,);
DFFARX1 I_3291 (I59538,I3563,I59314,I59303,);
nand I_3292 (I59560,I1380931,I1380928);
and I_3293 (I59577,I59560,I1380913);
DFFARX1 I_3294 (I59577,I3563,I59314,I59603,);
DFFARX1 I_3295 (I59603,I3563,I59314,I59620,);
not I_3296 (I59306,I59620);
not I_3297 (I59642,I59603);
nand I_3298 (I59291,I59642,I59481);
nor I_3299 (I59673,I1380913,I1380928);
not I_3300 (I59690,I59673);
nor I_3301 (I59707,I59642,I59690);
nor I_3302 (I59724,I59348,I59707);
DFFARX1 I_3303 (I59724,I3563,I59314,I59300,);
nor I_3304 (I59755,I59408,I59690);
nor I_3305 (I59288,I59603,I59755);
nor I_3306 (I59297,I59538,I59673);
nor I_3307 (I59285,I59408,I59673);
not I_3308 (I59841,I3570);
DFFARX1 I_3309 (I650330,I3563,I59841,I59867,);
not I_3310 (I59875,I59867);
nand I_3311 (I59892,I650342,I650327);
and I_3312 (I59909,I59892,I650321);
DFFARX1 I_3313 (I59909,I3563,I59841,I59935,);
DFFARX1 I_3314 (I650336,I3563,I59841,I59952,);
and I_3315 (I59960,I59952,I650324);
nor I_3316 (I59977,I59935,I59960);
DFFARX1 I_3317 (I59977,I3563,I59841,I59809,);
nand I_3318 (I60008,I59952,I650324);
nand I_3319 (I60025,I59875,I60008);
not I_3320 (I59821,I60025);
DFFARX1 I_3321 (I650333,I3563,I59841,I60065,);
DFFARX1 I_3322 (I60065,I3563,I59841,I59830,);
nand I_3323 (I60087,I650339,I650345);
and I_3324 (I60104,I60087,I650321);
DFFARX1 I_3325 (I60104,I3563,I59841,I60130,);
DFFARX1 I_3326 (I60130,I3563,I59841,I60147,);
not I_3327 (I59833,I60147);
not I_3328 (I60169,I60130);
nand I_3329 (I59818,I60169,I60008);
nor I_3330 (I60200,I650324,I650345);
not I_3331 (I60217,I60200);
nor I_3332 (I60234,I60169,I60217);
nor I_3333 (I60251,I59875,I60234);
DFFARX1 I_3334 (I60251,I3563,I59841,I59827,);
nor I_3335 (I60282,I59935,I60217);
nor I_3336 (I59815,I60130,I60282);
nor I_3337 (I59824,I60065,I60200);
nor I_3338 (I59812,I59935,I60200);
not I_3339 (I60368,I3570);
DFFARX1 I_3340 (I771135,I3563,I60368,I60394,);
not I_3341 (I60402,I60394);
nand I_3342 (I60419,I771126,I771144);
and I_3343 (I60436,I60419,I771123);
DFFARX1 I_3344 (I60436,I3563,I60368,I60462,);
DFFARX1 I_3345 (I771126,I3563,I60368,I60479,);
and I_3346 (I60487,I60479,I771129);
nor I_3347 (I60504,I60462,I60487);
DFFARX1 I_3348 (I60504,I3563,I60368,I60336,);
nand I_3349 (I60535,I60479,I771129);
nand I_3350 (I60552,I60402,I60535);
not I_3351 (I60348,I60552);
DFFARX1 I_3352 (I771123,I3563,I60368,I60592,);
DFFARX1 I_3353 (I60592,I3563,I60368,I60357,);
nand I_3354 (I60614,I771141,I771132);
and I_3355 (I60631,I60614,I771147);
DFFARX1 I_3356 (I60631,I3563,I60368,I60657,);
DFFARX1 I_3357 (I60657,I3563,I60368,I60674,);
not I_3358 (I60360,I60674);
not I_3359 (I60696,I60657);
nand I_3360 (I60345,I60696,I60535);
nor I_3361 (I60727,I771138,I771132);
not I_3362 (I60744,I60727);
nor I_3363 (I60761,I60696,I60744);
nor I_3364 (I60778,I60402,I60761);
DFFARX1 I_3365 (I60778,I3563,I60368,I60354,);
nor I_3366 (I60809,I60462,I60744);
nor I_3367 (I60342,I60657,I60809);
nor I_3368 (I60351,I60592,I60727);
nor I_3369 (I60339,I60462,I60727);
not I_3370 (I60895,I3570);
DFFARX1 I_3371 (I578080,I3563,I60895,I60921,);
not I_3372 (I60929,I60921);
nand I_3373 (I60946,I578092,I578077);
and I_3374 (I60963,I60946,I578071);
DFFARX1 I_3375 (I60963,I3563,I60895,I60989,);
DFFARX1 I_3376 (I578086,I3563,I60895,I61006,);
and I_3377 (I61014,I61006,I578074);
nor I_3378 (I61031,I60989,I61014);
DFFARX1 I_3379 (I61031,I3563,I60895,I60863,);
nand I_3380 (I61062,I61006,I578074);
nand I_3381 (I61079,I60929,I61062);
not I_3382 (I60875,I61079);
DFFARX1 I_3383 (I578083,I3563,I60895,I61119,);
DFFARX1 I_3384 (I61119,I3563,I60895,I60884,);
nand I_3385 (I61141,I578089,I578095);
and I_3386 (I61158,I61141,I578071);
DFFARX1 I_3387 (I61158,I3563,I60895,I61184,);
DFFARX1 I_3388 (I61184,I3563,I60895,I61201,);
not I_3389 (I60887,I61201);
not I_3390 (I61223,I61184);
nand I_3391 (I60872,I61223,I61062);
nor I_3392 (I61254,I578074,I578095);
not I_3393 (I61271,I61254);
nor I_3394 (I61288,I61223,I61271);
nor I_3395 (I61305,I60929,I61288);
DFFARX1 I_3396 (I61305,I3563,I60895,I60881,);
nor I_3397 (I61336,I60989,I61271);
nor I_3398 (I60869,I61184,I61336);
nor I_3399 (I60878,I61119,I61254);
nor I_3400 (I60866,I60989,I61254);
not I_3401 (I61422,I3570);
DFFARX1 I_3402 (I341781,I3563,I61422,I61448,);
not I_3403 (I61456,I61448);
nand I_3404 (I61473,I341763,I341778);
and I_3405 (I61490,I61473,I341754);
DFFARX1 I_3406 (I61490,I3563,I61422,I61516,);
DFFARX1 I_3407 (I341757,I3563,I61422,I61533,);
and I_3408 (I61541,I61533,I341772);
nor I_3409 (I61558,I61516,I61541);
DFFARX1 I_3410 (I61558,I3563,I61422,I61390,);
nand I_3411 (I61589,I61533,I341772);
nand I_3412 (I61606,I61456,I61589);
not I_3413 (I61402,I61606);
DFFARX1 I_3414 (I341775,I3563,I61422,I61646,);
DFFARX1 I_3415 (I61646,I3563,I61422,I61411,);
nand I_3416 (I61668,I341754,I341766);
and I_3417 (I61685,I61668,I341760);
DFFARX1 I_3418 (I61685,I3563,I61422,I61711,);
DFFARX1 I_3419 (I61711,I3563,I61422,I61728,);
not I_3420 (I61414,I61728);
not I_3421 (I61750,I61711);
nand I_3422 (I61399,I61750,I61589);
nor I_3423 (I61781,I341769,I341766);
not I_3424 (I61798,I61781);
nor I_3425 (I61815,I61750,I61798);
nor I_3426 (I61832,I61456,I61815);
DFFARX1 I_3427 (I61832,I3563,I61422,I61408,);
nor I_3428 (I61863,I61516,I61798);
nor I_3429 (I61396,I61711,I61863);
nor I_3430 (I61405,I61646,I61781);
nor I_3431 (I61393,I61516,I61781);
not I_3432 (I61949,I3570);
DFFARX1 I_3433 (I589062,I3563,I61949,I61975,);
not I_3434 (I61983,I61975);
nand I_3435 (I62000,I589074,I589059);
and I_3436 (I62017,I62000,I589053);
DFFARX1 I_3437 (I62017,I3563,I61949,I62043,);
DFFARX1 I_3438 (I589068,I3563,I61949,I62060,);
and I_3439 (I62068,I62060,I589056);
nor I_3440 (I62085,I62043,I62068);
DFFARX1 I_3441 (I62085,I3563,I61949,I61917,);
nand I_3442 (I62116,I62060,I589056);
nand I_3443 (I62133,I61983,I62116);
not I_3444 (I61929,I62133);
DFFARX1 I_3445 (I589065,I3563,I61949,I62173,);
DFFARX1 I_3446 (I62173,I3563,I61949,I61938,);
nand I_3447 (I62195,I589071,I589077);
and I_3448 (I62212,I62195,I589053);
DFFARX1 I_3449 (I62212,I3563,I61949,I62238,);
DFFARX1 I_3450 (I62238,I3563,I61949,I62255,);
not I_3451 (I61941,I62255);
not I_3452 (I62277,I62238);
nand I_3453 (I61926,I62277,I62116);
nor I_3454 (I62308,I589056,I589077);
not I_3455 (I62325,I62308);
nor I_3456 (I62342,I62277,I62325);
nor I_3457 (I62359,I61983,I62342);
DFFARX1 I_3458 (I62359,I3563,I61949,I61935,);
nor I_3459 (I62390,I62043,I62325);
nor I_3460 (I61923,I62238,I62390);
nor I_3461 (I61932,I62173,I62308);
nor I_3462 (I61920,I62043,I62308);
not I_3463 (I62476,I3570);
DFFARX1 I_3464 (I649752,I3563,I62476,I62502,);
not I_3465 (I62510,I62502);
nand I_3466 (I62527,I649764,I649749);
and I_3467 (I62544,I62527,I649743);
DFFARX1 I_3468 (I62544,I3563,I62476,I62570,);
DFFARX1 I_3469 (I649758,I3563,I62476,I62587,);
and I_3470 (I62595,I62587,I649746);
nor I_3471 (I62612,I62570,I62595);
DFFARX1 I_3472 (I62612,I3563,I62476,I62444,);
nand I_3473 (I62643,I62587,I649746);
nand I_3474 (I62660,I62510,I62643);
not I_3475 (I62456,I62660);
DFFARX1 I_3476 (I649755,I3563,I62476,I62700,);
DFFARX1 I_3477 (I62700,I3563,I62476,I62465,);
nand I_3478 (I62722,I649761,I649767);
and I_3479 (I62739,I62722,I649743);
DFFARX1 I_3480 (I62739,I3563,I62476,I62765,);
DFFARX1 I_3481 (I62765,I3563,I62476,I62782,);
not I_3482 (I62468,I62782);
not I_3483 (I62804,I62765);
nand I_3484 (I62453,I62804,I62643);
nor I_3485 (I62835,I649746,I649767);
not I_3486 (I62852,I62835);
nor I_3487 (I62869,I62804,I62852);
nor I_3488 (I62886,I62510,I62869);
DFFARX1 I_3489 (I62886,I3563,I62476,I62462,);
nor I_3490 (I62917,I62570,I62852);
nor I_3491 (I62450,I62765,I62917);
nor I_3492 (I62459,I62700,I62835);
nor I_3493 (I62447,I62570,I62835);
not I_3494 (I63003,I3570);
DFFARX1 I_3495 (I407129,I3563,I63003,I63029,);
not I_3496 (I63037,I63029);
nand I_3497 (I63054,I407111,I407126);
and I_3498 (I63071,I63054,I407102);
DFFARX1 I_3499 (I63071,I3563,I63003,I63097,);
DFFARX1 I_3500 (I407105,I3563,I63003,I63114,);
and I_3501 (I63122,I63114,I407120);
nor I_3502 (I63139,I63097,I63122);
DFFARX1 I_3503 (I63139,I3563,I63003,I62971,);
nand I_3504 (I63170,I63114,I407120);
nand I_3505 (I63187,I63037,I63170);
not I_3506 (I62983,I63187);
DFFARX1 I_3507 (I407123,I3563,I63003,I63227,);
DFFARX1 I_3508 (I63227,I3563,I63003,I62992,);
nand I_3509 (I63249,I407102,I407114);
and I_3510 (I63266,I63249,I407108);
DFFARX1 I_3511 (I63266,I3563,I63003,I63292,);
DFFARX1 I_3512 (I63292,I3563,I63003,I63309,);
not I_3513 (I62995,I63309);
not I_3514 (I63331,I63292);
nand I_3515 (I62980,I63331,I63170);
nor I_3516 (I63362,I407117,I407114);
not I_3517 (I63379,I63362);
nor I_3518 (I63396,I63331,I63379);
nor I_3519 (I63413,I63037,I63396);
DFFARX1 I_3520 (I63413,I3563,I63003,I62989,);
nor I_3521 (I63444,I63097,I63379);
nor I_3522 (I62977,I63292,I63444);
nor I_3523 (I62986,I63227,I63362);
nor I_3524 (I62974,I63097,I63362);
not I_3525 (I63530,I3570);
DFFARX1 I_3526 (I1532,I3563,I63530,I63556,);
not I_3527 (I63564,I63556);
nand I_3528 (I63581,I3532,I2412);
and I_3529 (I63598,I63581,I1388);
DFFARX1 I_3530 (I63598,I3563,I63530,I63624,);
DFFARX1 I_3531 (I1460,I3563,I63530,I63641,);
and I_3532 (I63649,I63641,I2788);
nor I_3533 (I63666,I63624,I63649);
DFFARX1 I_3534 (I63666,I3563,I63530,I63498,);
nand I_3535 (I63697,I63641,I2788);
nand I_3536 (I63714,I63564,I63697);
not I_3537 (I63510,I63714);
DFFARX1 I_3538 (I1996,I3563,I63530,I63754,);
DFFARX1 I_3539 (I63754,I3563,I63530,I63519,);
nand I_3540 (I63776,I2924,I2604);
and I_3541 (I63793,I63776,I2476);
DFFARX1 I_3542 (I63793,I3563,I63530,I63819,);
DFFARX1 I_3543 (I63819,I3563,I63530,I63836,);
not I_3544 (I63522,I63836);
not I_3545 (I63858,I63819);
nand I_3546 (I63507,I63858,I63697);
nor I_3547 (I63889,I3004,I2604);
not I_3548 (I63906,I63889);
nor I_3549 (I63923,I63858,I63906);
nor I_3550 (I63940,I63564,I63923);
DFFARX1 I_3551 (I63940,I3563,I63530,I63516,);
nor I_3552 (I63971,I63624,I63906);
nor I_3553 (I63504,I63819,I63971);
nor I_3554 (I63513,I63754,I63889);
nor I_3555 (I63501,I63624,I63889);
not I_3556 (I64057,I3570);
DFFARX1 I_3557 (I1009846,I3563,I64057,I64083,);
not I_3558 (I64091,I64083);
nand I_3559 (I64108,I1009864,I1009858);
and I_3560 (I64125,I64108,I1009837);
DFFARX1 I_3561 (I64125,I3563,I64057,I64151,);
DFFARX1 I_3562 (I1009855,I3563,I64057,I64168,);
and I_3563 (I64176,I64168,I1009840);
nor I_3564 (I64193,I64151,I64176);
DFFARX1 I_3565 (I64193,I3563,I64057,I64025,);
nand I_3566 (I64224,I64168,I1009840);
nand I_3567 (I64241,I64091,I64224);
not I_3568 (I64037,I64241);
DFFARX1 I_3569 (I1009852,I3563,I64057,I64281,);
DFFARX1 I_3570 (I64281,I3563,I64057,I64046,);
nand I_3571 (I64303,I1009861,I1009849);
and I_3572 (I64320,I64303,I1009843);
DFFARX1 I_3573 (I64320,I3563,I64057,I64346,);
DFFARX1 I_3574 (I64346,I3563,I64057,I64363,);
not I_3575 (I64049,I64363);
not I_3576 (I64385,I64346);
nand I_3577 (I64034,I64385,I64224);
nor I_3578 (I64416,I1009837,I1009849);
not I_3579 (I64433,I64416);
nor I_3580 (I64450,I64385,I64433);
nor I_3581 (I64467,I64091,I64450);
DFFARX1 I_3582 (I64467,I3563,I64057,I64043,);
nor I_3583 (I64498,I64151,I64433);
nor I_3584 (I64031,I64346,I64498);
nor I_3585 (I64040,I64281,I64416);
nor I_3586 (I64028,I64151,I64416);
not I_3587 (I64584,I3570);
DFFARX1 I_3588 (I361807,I3563,I64584,I64610,);
not I_3589 (I64618,I64610);
nand I_3590 (I64635,I361789,I361804);
and I_3591 (I64652,I64635,I361780);
DFFARX1 I_3592 (I64652,I3563,I64584,I64678,);
DFFARX1 I_3593 (I361783,I3563,I64584,I64695,);
and I_3594 (I64703,I64695,I361798);
nor I_3595 (I64720,I64678,I64703);
DFFARX1 I_3596 (I64720,I3563,I64584,I64552,);
nand I_3597 (I64751,I64695,I361798);
nand I_3598 (I64768,I64618,I64751);
not I_3599 (I64564,I64768);
DFFARX1 I_3600 (I361801,I3563,I64584,I64808,);
DFFARX1 I_3601 (I64808,I3563,I64584,I64573,);
nand I_3602 (I64830,I361780,I361792);
and I_3603 (I64847,I64830,I361786);
DFFARX1 I_3604 (I64847,I3563,I64584,I64873,);
DFFARX1 I_3605 (I64873,I3563,I64584,I64890,);
not I_3606 (I64576,I64890);
not I_3607 (I64912,I64873);
nand I_3608 (I64561,I64912,I64751);
nor I_3609 (I64943,I361795,I361792);
not I_3610 (I64960,I64943);
nor I_3611 (I64977,I64912,I64960);
nor I_3612 (I64994,I64618,I64977);
DFFARX1 I_3613 (I64994,I3563,I64584,I64570,);
nor I_3614 (I65025,I64678,I64960);
nor I_3615 (I64558,I64873,I65025);
nor I_3616 (I64567,I64808,I64943);
nor I_3617 (I64555,I64678,I64943);
not I_3618 (I65111,I3570);
DFFARX1 I_3619 (I617384,I3563,I65111,I65137,);
not I_3620 (I65145,I65137);
nand I_3621 (I65162,I617396,I617381);
and I_3622 (I65179,I65162,I617375);
DFFARX1 I_3623 (I65179,I3563,I65111,I65205,);
DFFARX1 I_3624 (I617390,I3563,I65111,I65222,);
and I_3625 (I65230,I65222,I617378);
nor I_3626 (I65247,I65205,I65230);
DFFARX1 I_3627 (I65247,I3563,I65111,I65079,);
nand I_3628 (I65278,I65222,I617378);
nand I_3629 (I65295,I65145,I65278);
not I_3630 (I65091,I65295);
DFFARX1 I_3631 (I617387,I3563,I65111,I65335,);
DFFARX1 I_3632 (I65335,I3563,I65111,I65100,);
nand I_3633 (I65357,I617393,I617399);
and I_3634 (I65374,I65357,I617375);
DFFARX1 I_3635 (I65374,I3563,I65111,I65400,);
DFFARX1 I_3636 (I65400,I3563,I65111,I65417,);
not I_3637 (I65103,I65417);
not I_3638 (I65439,I65400);
nand I_3639 (I65088,I65439,I65278);
nor I_3640 (I65470,I617378,I617399);
not I_3641 (I65487,I65470);
nor I_3642 (I65504,I65439,I65487);
nor I_3643 (I65521,I65145,I65504);
DFFARX1 I_3644 (I65521,I3563,I65111,I65097,);
nor I_3645 (I65552,I65205,I65487);
nor I_3646 (I65085,I65400,I65552);
nor I_3647 (I65094,I65335,I65470);
nor I_3648 (I65082,I65205,I65470);
not I_3649 (I65638,I3570);
DFFARX1 I_3650 (I437652,I3563,I65638,I65664,);
not I_3651 (I65672,I65664);
nand I_3652 (I65689,I437646,I437637);
and I_3653 (I65706,I65689,I437658);
DFFARX1 I_3654 (I65706,I3563,I65638,I65732,);
DFFARX1 I_3655 (I437640,I3563,I65638,I65749,);
and I_3656 (I65757,I65749,I437634);
nor I_3657 (I65774,I65732,I65757);
DFFARX1 I_3658 (I65774,I3563,I65638,I65606,);
nand I_3659 (I65805,I65749,I437634);
nand I_3660 (I65822,I65672,I65805);
not I_3661 (I65618,I65822);
DFFARX1 I_3662 (I437634,I3563,I65638,I65862,);
DFFARX1 I_3663 (I65862,I3563,I65638,I65627,);
nand I_3664 (I65884,I437661,I437643);
and I_3665 (I65901,I65884,I437649);
DFFARX1 I_3666 (I65901,I3563,I65638,I65927,);
DFFARX1 I_3667 (I65927,I3563,I65638,I65944,);
not I_3668 (I65630,I65944);
not I_3669 (I65966,I65927);
nand I_3670 (I65615,I65966,I65805);
nor I_3671 (I65997,I437655,I437643);
not I_3672 (I66014,I65997);
nor I_3673 (I66031,I65966,I66014);
nor I_3674 (I66048,I65672,I66031);
DFFARX1 I_3675 (I66048,I3563,I65638,I65624,);
nor I_3676 (I66079,I65732,I66014);
nor I_3677 (I65612,I65927,I66079);
nor I_3678 (I65621,I65862,I65997);
nor I_3679 (I65609,I65732,I65997);
not I_3680 (I66165,I3570);
DFFARX1 I_3681 (I1286671,I3563,I66165,I66191,);
not I_3682 (I66199,I66191);
nand I_3683 (I66216,I1286665,I1286686);
and I_3684 (I66233,I66216,I1286677);
DFFARX1 I_3685 (I66233,I3563,I66165,I66259,);
DFFARX1 I_3686 (I1286668,I3563,I66165,I66276,);
and I_3687 (I66284,I66276,I1286680);
nor I_3688 (I66301,I66259,I66284);
DFFARX1 I_3689 (I66301,I3563,I66165,I66133,);
nand I_3690 (I66332,I66276,I1286680);
nand I_3691 (I66349,I66199,I66332);
not I_3692 (I66145,I66349);
DFFARX1 I_3693 (I1286668,I3563,I66165,I66389,);
DFFARX1 I_3694 (I66389,I3563,I66165,I66154,);
nand I_3695 (I66411,I1286689,I1286674);
and I_3696 (I66428,I66411,I1286665);
DFFARX1 I_3697 (I66428,I3563,I66165,I66454,);
DFFARX1 I_3698 (I66454,I3563,I66165,I66471,);
not I_3699 (I66157,I66471);
not I_3700 (I66493,I66454);
nand I_3701 (I66142,I66493,I66332);
nor I_3702 (I66524,I1286683,I1286674);
not I_3703 (I66541,I66524);
nor I_3704 (I66558,I66493,I66541);
nor I_3705 (I66575,I66199,I66558);
DFFARX1 I_3706 (I66575,I3563,I66165,I66151,);
nor I_3707 (I66606,I66259,I66541);
nor I_3708 (I66139,I66454,I66606);
nor I_3709 (I66148,I66389,I66524);
nor I_3710 (I66136,I66259,I66524);
not I_3711 (I66692,I3570);
DFFARX1 I_3712 (I226795,I3563,I66692,I66718,);
not I_3713 (I66726,I66718);
nand I_3714 (I66743,I226789,I226783);
and I_3715 (I66760,I66743,I226804);
DFFARX1 I_3716 (I66760,I3563,I66692,I66786,);
DFFARX1 I_3717 (I226801,I3563,I66692,I66803,);
and I_3718 (I66811,I66803,I226798);
nor I_3719 (I66828,I66786,I66811);
DFFARX1 I_3720 (I66828,I3563,I66692,I66660,);
nand I_3721 (I66859,I66803,I226798);
nand I_3722 (I66876,I66726,I66859);
not I_3723 (I66672,I66876);
DFFARX1 I_3724 (I226783,I3563,I66692,I66916,);
DFFARX1 I_3725 (I66916,I3563,I66692,I66681,);
nand I_3726 (I66938,I226786,I226786);
and I_3727 (I66955,I66938,I226807);
DFFARX1 I_3728 (I66955,I3563,I66692,I66981,);
DFFARX1 I_3729 (I66981,I3563,I66692,I66998,);
not I_3730 (I66684,I66998);
not I_3731 (I67020,I66981);
nand I_3732 (I66669,I67020,I66859);
nor I_3733 (I67051,I226792,I226786);
not I_3734 (I67068,I67051);
nor I_3735 (I67085,I67020,I67068);
nor I_3736 (I67102,I66726,I67085);
DFFARX1 I_3737 (I67102,I3563,I66692,I66678,);
nor I_3738 (I67133,I66786,I67068);
nor I_3739 (I66666,I66981,I67133);
nor I_3740 (I66675,I66916,I67051);
nor I_3741 (I66663,I66786,I67051);
not I_3742 (I67219,I3570);
DFFARX1 I_3743 (I891169,I3563,I67219,I67245,);
not I_3744 (I67253,I67245);
nand I_3745 (I67270,I891166,I891181);
and I_3746 (I67287,I67270,I891163);
DFFARX1 I_3747 (I67287,I3563,I67219,I67313,);
DFFARX1 I_3748 (I891160,I3563,I67219,I67330,);
and I_3749 (I67338,I67330,I891160);
nor I_3750 (I67355,I67313,I67338);
DFFARX1 I_3751 (I67355,I3563,I67219,I67187,);
nand I_3752 (I67386,I67330,I891160);
nand I_3753 (I67403,I67253,I67386);
not I_3754 (I67199,I67403);
DFFARX1 I_3755 (I891163,I3563,I67219,I67443,);
DFFARX1 I_3756 (I67443,I3563,I67219,I67208,);
nand I_3757 (I67465,I891175,I891166);
and I_3758 (I67482,I67465,I891178);
DFFARX1 I_3759 (I67482,I3563,I67219,I67508,);
DFFARX1 I_3760 (I67508,I3563,I67219,I67525,);
not I_3761 (I67211,I67525);
not I_3762 (I67547,I67508);
nand I_3763 (I67196,I67547,I67386);
nor I_3764 (I67578,I891172,I891166);
not I_3765 (I67595,I67578);
nor I_3766 (I67612,I67547,I67595);
nor I_3767 (I67629,I67253,I67612);
DFFARX1 I_3768 (I67629,I3563,I67219,I67205,);
nor I_3769 (I67660,I67313,I67595);
nor I_3770 (I67193,I67508,I67660);
nor I_3771 (I67202,I67443,I67578);
nor I_3772 (I67190,I67313,I67578);
not I_3773 (I67746,I3570);
DFFARX1 I_3774 (I1137241,I3563,I67746,I67772,);
not I_3775 (I67780,I67772);
nand I_3776 (I67797,I1137256,I1137235);
and I_3777 (I67814,I67797,I1137238);
DFFARX1 I_3778 (I67814,I3563,I67746,I67840,);
DFFARX1 I_3779 (I1137259,I3563,I67746,I67857,);
and I_3780 (I67865,I67857,I1137238);
nor I_3781 (I67882,I67840,I67865);
DFFARX1 I_3782 (I67882,I3563,I67746,I67714,);
nand I_3783 (I67913,I67857,I1137238);
nand I_3784 (I67930,I67780,I67913);
not I_3785 (I67726,I67930);
DFFARX1 I_3786 (I1137235,I3563,I67746,I67970,);
DFFARX1 I_3787 (I67970,I3563,I67746,I67735,);
nand I_3788 (I67992,I1137247,I1137244);
and I_3789 (I68009,I67992,I1137250);
DFFARX1 I_3790 (I68009,I3563,I67746,I68035,);
DFFARX1 I_3791 (I68035,I3563,I67746,I68052,);
not I_3792 (I67738,I68052);
not I_3793 (I68074,I68035);
nand I_3794 (I67723,I68074,I67913);
nor I_3795 (I68105,I1137253,I1137244);
not I_3796 (I68122,I68105);
nor I_3797 (I68139,I68074,I68122);
nor I_3798 (I68156,I67780,I68139);
DFFARX1 I_3799 (I68156,I3563,I67746,I67732,);
nor I_3800 (I68187,I67840,I68122);
nor I_3801 (I67720,I68035,I68187);
nor I_3802 (I67729,I67970,I68105);
nor I_3803 (I67717,I67840,I68105);
not I_3804 (I68273,I3570);
DFFARX1 I_3805 (I849009,I3563,I68273,I68299,);
not I_3806 (I68307,I68299);
nand I_3807 (I68324,I849006,I849021);
and I_3808 (I68341,I68324,I849003);
DFFARX1 I_3809 (I68341,I3563,I68273,I68367,);
DFFARX1 I_3810 (I849000,I3563,I68273,I68384,);
and I_3811 (I68392,I68384,I849000);
nor I_3812 (I68409,I68367,I68392);
DFFARX1 I_3813 (I68409,I3563,I68273,I68241,);
nand I_3814 (I68440,I68384,I849000);
nand I_3815 (I68457,I68307,I68440);
not I_3816 (I68253,I68457);
DFFARX1 I_3817 (I849003,I3563,I68273,I68497,);
DFFARX1 I_3818 (I68497,I3563,I68273,I68262,);
nand I_3819 (I68519,I849015,I849006);
and I_3820 (I68536,I68519,I849018);
DFFARX1 I_3821 (I68536,I3563,I68273,I68562,);
DFFARX1 I_3822 (I68562,I3563,I68273,I68579,);
not I_3823 (I68265,I68579);
not I_3824 (I68601,I68562);
nand I_3825 (I68250,I68601,I68440);
nor I_3826 (I68632,I849012,I849006);
not I_3827 (I68649,I68632);
nor I_3828 (I68666,I68601,I68649);
nor I_3829 (I68683,I68307,I68666);
DFFARX1 I_3830 (I68683,I3563,I68273,I68259,);
nor I_3831 (I68714,I68367,I68649);
nor I_3832 (I68247,I68562,I68714);
nor I_3833 (I68256,I68497,I68632);
nor I_3834 (I68244,I68367,I68632);
not I_3835 (I68800,I3570);
DFFARX1 I_3836 (I1258383,I3563,I68800,I68826,);
not I_3837 (I68834,I68826);
nand I_3838 (I68851,I1258377,I1258398);
and I_3839 (I68868,I68851,I1258389);
DFFARX1 I_3840 (I68868,I3563,I68800,I68894,);
DFFARX1 I_3841 (I1258380,I3563,I68800,I68911,);
and I_3842 (I68919,I68911,I1258392);
nor I_3843 (I68936,I68894,I68919);
DFFARX1 I_3844 (I68936,I3563,I68800,I68768,);
nand I_3845 (I68967,I68911,I1258392);
nand I_3846 (I68984,I68834,I68967);
not I_3847 (I68780,I68984);
DFFARX1 I_3848 (I1258380,I3563,I68800,I69024,);
DFFARX1 I_3849 (I69024,I3563,I68800,I68789,);
nand I_3850 (I69046,I1258401,I1258386);
and I_3851 (I69063,I69046,I1258377);
DFFARX1 I_3852 (I69063,I3563,I68800,I69089,);
DFFARX1 I_3853 (I69089,I3563,I68800,I69106,);
not I_3854 (I68792,I69106);
not I_3855 (I69128,I69089);
nand I_3856 (I68777,I69128,I68967);
nor I_3857 (I69159,I1258395,I1258386);
not I_3858 (I69176,I69159);
nor I_3859 (I69193,I69128,I69176);
nor I_3860 (I69210,I68834,I69193);
DFFARX1 I_3861 (I69210,I3563,I68800,I68786,);
nor I_3862 (I69241,I68894,I69176);
nor I_3863 (I68774,I69089,I69241);
nor I_3864 (I68783,I69024,I69159);
nor I_3865 (I68771,I68894,I69159);
not I_3866 (I69327,I3570);
DFFARX1 I_3867 (I1005324,I3563,I69327,I69353,);
not I_3868 (I69361,I69353);
nand I_3869 (I69378,I1005342,I1005336);
and I_3870 (I69395,I69378,I1005315);
DFFARX1 I_3871 (I69395,I3563,I69327,I69421,);
DFFARX1 I_3872 (I1005333,I3563,I69327,I69438,);
and I_3873 (I69446,I69438,I1005318);
nor I_3874 (I69463,I69421,I69446);
DFFARX1 I_3875 (I69463,I3563,I69327,I69295,);
nand I_3876 (I69494,I69438,I1005318);
nand I_3877 (I69511,I69361,I69494);
not I_3878 (I69307,I69511);
DFFARX1 I_3879 (I1005330,I3563,I69327,I69551,);
DFFARX1 I_3880 (I69551,I3563,I69327,I69316,);
nand I_3881 (I69573,I1005339,I1005327);
and I_3882 (I69590,I69573,I1005321);
DFFARX1 I_3883 (I69590,I3563,I69327,I69616,);
DFFARX1 I_3884 (I69616,I3563,I69327,I69633,);
not I_3885 (I69319,I69633);
not I_3886 (I69655,I69616);
nand I_3887 (I69304,I69655,I69494);
nor I_3888 (I69686,I1005315,I1005327);
not I_3889 (I69703,I69686);
nor I_3890 (I69720,I69655,I69703);
nor I_3891 (I69737,I69361,I69720);
DFFARX1 I_3892 (I69737,I3563,I69327,I69313,);
nor I_3893 (I69768,I69421,I69703);
nor I_3894 (I69301,I69616,I69768);
nor I_3895 (I69310,I69551,I69686);
nor I_3896 (I69298,I69421,I69686);
not I_3897 (I69854,I3570);
DFFARX1 I_3898 (I1355340,I3563,I69854,I69880,);
not I_3899 (I69888,I69880);
nand I_3900 (I69905,I1355334,I1355355);
and I_3901 (I69922,I69905,I1355331);
DFFARX1 I_3902 (I69922,I3563,I69854,I69948,);
DFFARX1 I_3903 (I1355352,I3563,I69854,I69965,);
and I_3904 (I69973,I69965,I1355349);
nor I_3905 (I69990,I69948,I69973);
DFFARX1 I_3906 (I69990,I3563,I69854,I69822,);
nand I_3907 (I70021,I69965,I1355349);
nand I_3908 (I70038,I69888,I70021);
not I_3909 (I69834,I70038);
DFFARX1 I_3910 (I1355337,I3563,I69854,I70078,);
DFFARX1 I_3911 (I70078,I3563,I69854,I69843,);
nand I_3912 (I70100,I1355346,I1355343);
and I_3913 (I70117,I70100,I1355328);
DFFARX1 I_3914 (I70117,I3563,I69854,I70143,);
DFFARX1 I_3915 (I70143,I3563,I69854,I70160,);
not I_3916 (I69846,I70160);
not I_3917 (I70182,I70143);
nand I_3918 (I69831,I70182,I70021);
nor I_3919 (I70213,I1355328,I1355343);
not I_3920 (I70230,I70213);
nor I_3921 (I70247,I70182,I70230);
nor I_3922 (I70264,I69888,I70247);
DFFARX1 I_3923 (I70264,I3563,I69854,I69840,);
nor I_3924 (I70295,I69948,I70230);
nor I_3925 (I69828,I70143,I70295);
nor I_3926 (I69837,I70078,I70213);
nor I_3927 (I69825,I69948,I70213);
not I_3928 (I70381,I3570);
DFFARX1 I_3929 (I1034394,I3563,I70381,I70407,);
not I_3930 (I70415,I70407);
nand I_3931 (I70432,I1034412,I1034406);
and I_3932 (I70449,I70432,I1034385);
DFFARX1 I_3933 (I70449,I3563,I70381,I70475,);
DFFARX1 I_3934 (I1034403,I3563,I70381,I70492,);
and I_3935 (I70500,I70492,I1034388);
nor I_3936 (I70517,I70475,I70500);
DFFARX1 I_3937 (I70517,I3563,I70381,I70349,);
nand I_3938 (I70548,I70492,I1034388);
nand I_3939 (I70565,I70415,I70548);
not I_3940 (I70361,I70565);
DFFARX1 I_3941 (I1034400,I3563,I70381,I70605,);
DFFARX1 I_3942 (I70605,I3563,I70381,I70370,);
nand I_3943 (I70627,I1034409,I1034397);
and I_3944 (I70644,I70627,I1034391);
DFFARX1 I_3945 (I70644,I3563,I70381,I70670,);
DFFARX1 I_3946 (I70670,I3563,I70381,I70687,);
not I_3947 (I70373,I70687);
not I_3948 (I70709,I70670);
nand I_3949 (I70358,I70709,I70548);
nor I_3950 (I70740,I1034385,I1034397);
not I_3951 (I70757,I70740);
nor I_3952 (I70774,I70709,I70757);
nor I_3953 (I70791,I70415,I70774);
DFFARX1 I_3954 (I70791,I3563,I70381,I70367,);
nor I_3955 (I70822,I70475,I70757);
nor I_3956 (I70355,I70670,I70822);
nor I_3957 (I70364,I70605,I70740);
nor I_3958 (I70352,I70475,I70740);
not I_3959 (I70908,I3570);
DFFARX1 I_3960 (I1308582,I3563,I70908,I70934,);
not I_3961 (I70942,I70934);
nand I_3962 (I70959,I1308585,I1308579);
and I_3963 (I70976,I70959,I1308576);
DFFARX1 I_3964 (I70976,I3563,I70908,I71002,);
DFFARX1 I_3965 (I1308561,I3563,I70908,I71019,);
and I_3966 (I71027,I71019,I1308570);
nor I_3967 (I71044,I71002,I71027);
DFFARX1 I_3968 (I71044,I3563,I70908,I70876,);
nand I_3969 (I71075,I71019,I1308570);
nand I_3970 (I71092,I70942,I71075);
not I_3971 (I70888,I71092);
DFFARX1 I_3972 (I1308561,I3563,I70908,I71132,);
DFFARX1 I_3973 (I71132,I3563,I70908,I70897,);
nand I_3974 (I71154,I1308564,I1308567);
and I_3975 (I71171,I71154,I1308573);
DFFARX1 I_3976 (I71171,I3563,I70908,I71197,);
DFFARX1 I_3977 (I71197,I3563,I70908,I71214,);
not I_3978 (I70900,I71214);
not I_3979 (I71236,I71197);
nand I_3980 (I70885,I71236,I71075);
nor I_3981 (I71267,I1308564,I1308567);
not I_3982 (I71284,I71267);
nor I_3983 (I71301,I71236,I71284);
nor I_3984 (I71318,I70942,I71301);
DFFARX1 I_3985 (I71318,I3563,I70908,I70894,);
nor I_3986 (I71349,I71002,I71284);
nor I_3987 (I70882,I71197,I71349);
nor I_3988 (I70891,I71132,I71267);
nor I_3989 (I70879,I71002,I71267);
not I_3990 (I71435,I3570);
DFFARX1 I_3991 (I1127415,I3563,I71435,I71461,);
not I_3992 (I71469,I71461);
nand I_3993 (I71486,I1127430,I1127409);
and I_3994 (I71503,I71486,I1127412);
DFFARX1 I_3995 (I71503,I3563,I71435,I71529,);
DFFARX1 I_3996 (I1127433,I3563,I71435,I71546,);
and I_3997 (I71554,I71546,I1127412);
nor I_3998 (I71571,I71529,I71554);
DFFARX1 I_3999 (I71571,I3563,I71435,I71403,);
nand I_4000 (I71602,I71546,I1127412);
nand I_4001 (I71619,I71469,I71602);
not I_4002 (I71415,I71619);
DFFARX1 I_4003 (I1127409,I3563,I71435,I71659,);
DFFARX1 I_4004 (I71659,I3563,I71435,I71424,);
nand I_4005 (I71681,I1127421,I1127418);
and I_4006 (I71698,I71681,I1127424);
DFFARX1 I_4007 (I71698,I3563,I71435,I71724,);
DFFARX1 I_4008 (I71724,I3563,I71435,I71741,);
not I_4009 (I71427,I71741);
not I_4010 (I71763,I71724);
nand I_4011 (I71412,I71763,I71602);
nor I_4012 (I71794,I1127427,I1127418);
not I_4013 (I71811,I71794);
nor I_4014 (I71828,I71763,I71811);
nor I_4015 (I71845,I71469,I71828);
DFFARX1 I_4016 (I71845,I3563,I71435,I71421,);
nor I_4017 (I71876,I71529,I71811);
nor I_4018 (I71409,I71724,I71876);
nor I_4019 (I71418,I71659,I71794);
nor I_4020 (I71406,I71529,I71794);
not I_4021 (I71962,I3570);
DFFARX1 I_4022 (I358645,I3563,I71962,I71988,);
not I_4023 (I71996,I71988);
nand I_4024 (I72013,I358627,I358642);
and I_4025 (I72030,I72013,I358618);
DFFARX1 I_4026 (I72030,I3563,I71962,I72056,);
DFFARX1 I_4027 (I358621,I3563,I71962,I72073,);
and I_4028 (I72081,I72073,I358636);
nor I_4029 (I72098,I72056,I72081);
DFFARX1 I_4030 (I72098,I3563,I71962,I71930,);
nand I_4031 (I72129,I72073,I358636);
nand I_4032 (I72146,I71996,I72129);
not I_4033 (I71942,I72146);
DFFARX1 I_4034 (I358639,I3563,I71962,I72186,);
DFFARX1 I_4035 (I72186,I3563,I71962,I71951,);
nand I_4036 (I72208,I358618,I358630);
and I_4037 (I72225,I72208,I358624);
DFFARX1 I_4038 (I72225,I3563,I71962,I72251,);
DFFARX1 I_4039 (I72251,I3563,I71962,I72268,);
not I_4040 (I71954,I72268);
not I_4041 (I72290,I72251);
nand I_4042 (I71939,I72290,I72129);
nor I_4043 (I72321,I358633,I358630);
not I_4044 (I72338,I72321);
nor I_4045 (I72355,I72290,I72338);
nor I_4046 (I72372,I71996,I72355);
DFFARX1 I_4047 (I72372,I3563,I71962,I71948,);
nor I_4048 (I72403,I72056,I72338);
nor I_4049 (I71936,I72251,I72403);
nor I_4050 (I71945,I72186,I72321);
nor I_4051 (I71933,I72056,I72321);
not I_4052 (I72489,I3570);
DFFARX1 I_4053 (I6563,I3563,I72489,I72515,);
not I_4054 (I72523,I72515);
nand I_4055 (I72540,I6548,I6548);
and I_4056 (I72557,I72540,I6569);
DFFARX1 I_4057 (I72557,I3563,I72489,I72583,);
DFFARX1 I_4058 (I6551,I3563,I72489,I72600,);
and I_4059 (I72608,I72600,I6560);
nor I_4060 (I72625,I72583,I72608);
DFFARX1 I_4061 (I72625,I3563,I72489,I72457,);
nand I_4062 (I72656,I72600,I6560);
nand I_4063 (I72673,I72523,I72656);
not I_4064 (I72469,I72673);
DFFARX1 I_4065 (I6554,I3563,I72489,I72713,);
DFFARX1 I_4066 (I72713,I3563,I72489,I72478,);
nand I_4067 (I72735,I6557,I6566);
and I_4068 (I72752,I72735,I6551);
DFFARX1 I_4069 (I72752,I3563,I72489,I72778,);
DFFARX1 I_4070 (I72778,I3563,I72489,I72795,);
not I_4071 (I72481,I72795);
not I_4072 (I72817,I72778);
nand I_4073 (I72466,I72817,I72656);
nor I_4074 (I72848,I6554,I6566);
not I_4075 (I72865,I72848);
nor I_4076 (I72882,I72817,I72865);
nor I_4077 (I72899,I72523,I72882);
DFFARX1 I_4078 (I72899,I3563,I72489,I72475,);
nor I_4079 (I72930,I72583,I72865);
nor I_4080 (I72463,I72778,I72930);
nor I_4081 (I72472,I72713,I72848);
nor I_4082 (I72460,I72583,I72848);
not I_4083 (I73016,I3570);
DFFARX1 I_4084 (I208350,I3563,I73016,I73042,);
not I_4085 (I73050,I73042);
nand I_4086 (I73067,I208344,I208338);
and I_4087 (I73084,I73067,I208359);
DFFARX1 I_4088 (I73084,I3563,I73016,I73110,);
DFFARX1 I_4089 (I208356,I3563,I73016,I73127,);
and I_4090 (I73135,I73127,I208353);
nor I_4091 (I73152,I73110,I73135);
DFFARX1 I_4092 (I73152,I3563,I73016,I72984,);
nand I_4093 (I73183,I73127,I208353);
nand I_4094 (I73200,I73050,I73183);
not I_4095 (I72996,I73200);
DFFARX1 I_4096 (I208338,I3563,I73016,I73240,);
DFFARX1 I_4097 (I73240,I3563,I73016,I73005,);
nand I_4098 (I73262,I208341,I208341);
and I_4099 (I73279,I73262,I208362);
DFFARX1 I_4100 (I73279,I3563,I73016,I73305,);
DFFARX1 I_4101 (I73305,I3563,I73016,I73322,);
not I_4102 (I73008,I73322);
not I_4103 (I73344,I73305);
nand I_4104 (I72993,I73344,I73183);
nor I_4105 (I73375,I208347,I208341);
not I_4106 (I73392,I73375);
nor I_4107 (I73409,I73344,I73392);
nor I_4108 (I73426,I73050,I73409);
DFFARX1 I_4109 (I73426,I3563,I73016,I73002,);
nor I_4110 (I73457,I73110,I73392);
nor I_4111 (I72990,I73305,I73457);
nor I_4112 (I72999,I73240,I73375);
nor I_4113 (I72987,I73110,I73375);
not I_4114 (I73543,I3570);
DFFARX1 I_4115 (I887480,I3563,I73543,I73569,);
not I_4116 (I73577,I73569);
nand I_4117 (I73594,I887477,I887492);
and I_4118 (I73611,I73594,I887474);
DFFARX1 I_4119 (I73611,I3563,I73543,I73637,);
DFFARX1 I_4120 (I887471,I3563,I73543,I73654,);
and I_4121 (I73662,I73654,I887471);
nor I_4122 (I73679,I73637,I73662);
DFFARX1 I_4123 (I73679,I3563,I73543,I73511,);
nand I_4124 (I73710,I73654,I887471);
nand I_4125 (I73727,I73577,I73710);
not I_4126 (I73523,I73727);
DFFARX1 I_4127 (I887474,I3563,I73543,I73767,);
DFFARX1 I_4128 (I73767,I3563,I73543,I73532,);
nand I_4129 (I73789,I887486,I887477);
and I_4130 (I73806,I73789,I887489);
DFFARX1 I_4131 (I73806,I3563,I73543,I73832,);
DFFARX1 I_4132 (I73832,I3563,I73543,I73849,);
not I_4133 (I73535,I73849);
not I_4134 (I73871,I73832);
nand I_4135 (I73520,I73871,I73710);
nor I_4136 (I73902,I887483,I887477);
not I_4137 (I73919,I73902);
nor I_4138 (I73936,I73871,I73919);
nor I_4139 (I73953,I73577,I73936);
DFFARX1 I_4140 (I73953,I3563,I73543,I73529,);
nor I_4141 (I73984,I73637,I73919);
nor I_4142 (I73517,I73832,I73984);
nor I_4143 (I73526,I73767,I73902);
nor I_4144 (I73514,I73637,I73902);
not I_4145 (I74070,I3570);
DFFARX1 I_4146 (I526309,I3563,I74070,I74096,);
not I_4147 (I74104,I74096);
nand I_4148 (I74121,I526330,I526324);
and I_4149 (I74138,I74121,I526306);
DFFARX1 I_4150 (I74138,I3563,I74070,I74164,);
DFFARX1 I_4151 (I526309,I3563,I74070,I74181,);
and I_4152 (I74189,I74181,I526318);
nor I_4153 (I74206,I74164,I74189);
DFFARX1 I_4154 (I74206,I3563,I74070,I74038,);
nand I_4155 (I74237,I74181,I526318);
nand I_4156 (I74254,I74104,I74237);
not I_4157 (I74050,I74254);
DFFARX1 I_4158 (I526315,I3563,I74070,I74294,);
DFFARX1 I_4159 (I74294,I3563,I74070,I74059,);
nand I_4160 (I74316,I526321,I526312);
and I_4161 (I74333,I74316,I526306);
DFFARX1 I_4162 (I74333,I3563,I74070,I74359,);
DFFARX1 I_4163 (I74359,I3563,I74070,I74376,);
not I_4164 (I74062,I74376);
not I_4165 (I74398,I74359);
nand I_4166 (I74047,I74398,I74237);
nor I_4167 (I74429,I526327,I526312);
not I_4168 (I74446,I74429);
nor I_4169 (I74463,I74398,I74446);
nor I_4170 (I74480,I74104,I74463);
DFFARX1 I_4171 (I74480,I3563,I74070,I74056,);
nor I_4172 (I74511,I74164,I74446);
nor I_4173 (I74044,I74359,I74511);
nor I_4174 (I74053,I74294,I74429);
nor I_4175 (I74041,I74164,I74429);
not I_4176 (I74597,I3570);
DFFARX1 I_4177 (I206565,I3563,I74597,I74623,);
not I_4178 (I74631,I74623);
nand I_4179 (I74648,I206559,I206553);
and I_4180 (I74665,I74648,I206574);
DFFARX1 I_4181 (I74665,I3563,I74597,I74691,);
DFFARX1 I_4182 (I206571,I3563,I74597,I74708,);
and I_4183 (I74716,I74708,I206568);
nor I_4184 (I74733,I74691,I74716);
DFFARX1 I_4185 (I74733,I3563,I74597,I74565,);
nand I_4186 (I74764,I74708,I206568);
nand I_4187 (I74781,I74631,I74764);
not I_4188 (I74577,I74781);
DFFARX1 I_4189 (I206553,I3563,I74597,I74821,);
DFFARX1 I_4190 (I74821,I3563,I74597,I74586,);
nand I_4191 (I74843,I206556,I206556);
and I_4192 (I74860,I74843,I206577);
DFFARX1 I_4193 (I74860,I3563,I74597,I74886,);
DFFARX1 I_4194 (I74886,I3563,I74597,I74903,);
not I_4195 (I74589,I74903);
not I_4196 (I74925,I74886);
nand I_4197 (I74574,I74925,I74764);
nor I_4198 (I74956,I206562,I206556);
not I_4199 (I74973,I74956);
nor I_4200 (I74990,I74925,I74973);
nor I_4201 (I75007,I74631,I74990);
DFFARX1 I_4202 (I75007,I3563,I74597,I74583,);
nor I_4203 (I75038,I74691,I74973);
nor I_4204 (I74571,I74886,I75038);
nor I_4205 (I74580,I74821,I74956);
nor I_4206 (I74568,I74691,I74956);
not I_4207 (I75124,I3570);
DFFARX1 I_4208 (I2620,I3563,I75124,I75150,);
not I_4209 (I75158,I75150);
nand I_4210 (I75175,I3500,I2556);
and I_4211 (I75192,I75175,I1916);
DFFARX1 I_4212 (I75192,I3563,I75124,I75218,);
DFFARX1 I_4213 (I3396,I3563,I75124,I75235,);
and I_4214 (I75243,I75235,I2396);
nor I_4215 (I75260,I75218,I75243);
DFFARX1 I_4216 (I75260,I3563,I75124,I75092,);
nand I_4217 (I75291,I75235,I2396);
nand I_4218 (I75308,I75158,I75291);
not I_4219 (I75104,I75308);
DFFARX1 I_4220 (I2004,I3563,I75124,I75348,);
DFFARX1 I_4221 (I75348,I3563,I75124,I75113,);
nand I_4222 (I75370,I2044,I2380);
and I_4223 (I75387,I75370,I1540);
DFFARX1 I_4224 (I75387,I3563,I75124,I75413,);
DFFARX1 I_4225 (I75413,I3563,I75124,I75430,);
not I_4226 (I75116,I75430);
not I_4227 (I75452,I75413);
nand I_4228 (I75101,I75452,I75291);
nor I_4229 (I75483,I3356,I2380);
not I_4230 (I75500,I75483);
nor I_4231 (I75517,I75452,I75500);
nor I_4232 (I75534,I75158,I75517);
DFFARX1 I_4233 (I75534,I3563,I75124,I75110,);
nor I_4234 (I75565,I75218,I75500);
nor I_4235 (I75098,I75413,I75565);
nor I_4236 (I75107,I75348,I75483);
nor I_4237 (I75095,I75218,I75483);
not I_4238 (I75651,I3570);
DFFARX1 I_4239 (I471380,I3563,I75651,I75677,);
not I_4240 (I75685,I75677);
nand I_4241 (I75702,I471374,I471365);
and I_4242 (I75719,I75702,I471386);
DFFARX1 I_4243 (I75719,I3563,I75651,I75745,);
DFFARX1 I_4244 (I471368,I3563,I75651,I75762,);
and I_4245 (I75770,I75762,I471362);
nor I_4246 (I75787,I75745,I75770);
DFFARX1 I_4247 (I75787,I3563,I75651,I75619,);
nand I_4248 (I75818,I75762,I471362);
nand I_4249 (I75835,I75685,I75818);
not I_4250 (I75631,I75835);
DFFARX1 I_4251 (I471362,I3563,I75651,I75875,);
DFFARX1 I_4252 (I75875,I3563,I75651,I75640,);
nand I_4253 (I75897,I471389,I471371);
and I_4254 (I75914,I75897,I471377);
DFFARX1 I_4255 (I75914,I3563,I75651,I75940,);
DFFARX1 I_4256 (I75940,I3563,I75651,I75957,);
not I_4257 (I75643,I75957);
not I_4258 (I75979,I75940);
nand I_4259 (I75628,I75979,I75818);
nor I_4260 (I76010,I471383,I471371);
not I_4261 (I76027,I76010);
nor I_4262 (I76044,I75979,I76027);
nor I_4263 (I76061,I75685,I76044);
DFFARX1 I_4264 (I76061,I3563,I75651,I75637,);
nor I_4265 (I76092,I75745,I76027);
nor I_4266 (I75625,I75940,I76092);
nor I_4267 (I75634,I75875,I76010);
nor I_4268 (I75622,I75745,I76010);
not I_4269 (I76178,I3570);
DFFARX1 I_4270 (I254760,I3563,I76178,I76204,);
not I_4271 (I76212,I76204);
nand I_4272 (I76229,I254754,I254748);
and I_4273 (I76246,I76229,I254769);
DFFARX1 I_4274 (I76246,I3563,I76178,I76272,);
DFFARX1 I_4275 (I254766,I3563,I76178,I76289,);
and I_4276 (I76297,I76289,I254763);
nor I_4277 (I76314,I76272,I76297);
DFFARX1 I_4278 (I76314,I3563,I76178,I76146,);
nand I_4279 (I76345,I76289,I254763);
nand I_4280 (I76362,I76212,I76345);
not I_4281 (I76158,I76362);
DFFARX1 I_4282 (I254748,I3563,I76178,I76402,);
DFFARX1 I_4283 (I76402,I3563,I76178,I76167,);
nand I_4284 (I76424,I254751,I254751);
and I_4285 (I76441,I76424,I254772);
DFFARX1 I_4286 (I76441,I3563,I76178,I76467,);
DFFARX1 I_4287 (I76467,I3563,I76178,I76484,);
not I_4288 (I76170,I76484);
not I_4289 (I76506,I76467);
nand I_4290 (I76155,I76506,I76345);
nor I_4291 (I76537,I254757,I254751);
not I_4292 (I76554,I76537);
nor I_4293 (I76571,I76506,I76554);
nor I_4294 (I76588,I76212,I76571);
DFFARX1 I_4295 (I76588,I3563,I76178,I76164,);
nor I_4296 (I76619,I76272,I76554);
nor I_4297 (I76152,I76467,I76619);
nor I_4298 (I76161,I76402,I76537);
nor I_4299 (I76149,I76272,I76537);
not I_4300 (I76705,I3570);
DFFARX1 I_4301 (I379725,I3563,I76705,I76731,);
not I_4302 (I76739,I76731);
nand I_4303 (I76756,I379707,I379722);
and I_4304 (I76773,I76756,I379698);
DFFARX1 I_4305 (I76773,I3563,I76705,I76799,);
DFFARX1 I_4306 (I379701,I3563,I76705,I76816,);
and I_4307 (I76824,I76816,I379716);
nor I_4308 (I76841,I76799,I76824);
DFFARX1 I_4309 (I76841,I3563,I76705,I76673,);
nand I_4310 (I76872,I76816,I379716);
nand I_4311 (I76889,I76739,I76872);
not I_4312 (I76685,I76889);
DFFARX1 I_4313 (I379719,I3563,I76705,I76929,);
DFFARX1 I_4314 (I76929,I3563,I76705,I76694,);
nand I_4315 (I76951,I379698,I379710);
and I_4316 (I76968,I76951,I379704);
DFFARX1 I_4317 (I76968,I3563,I76705,I76994,);
DFFARX1 I_4318 (I76994,I3563,I76705,I77011,);
not I_4319 (I76697,I77011);
not I_4320 (I77033,I76994);
nand I_4321 (I76682,I77033,I76872);
nor I_4322 (I77064,I379713,I379710);
not I_4323 (I77081,I77064);
nor I_4324 (I77098,I77033,I77081);
nor I_4325 (I77115,I76739,I77098);
DFFARX1 I_4326 (I77115,I3563,I76705,I76691,);
nor I_4327 (I77146,I76799,I77081);
nor I_4328 (I76679,I76994,I77146);
nor I_4329 (I76688,I76929,I77064);
nor I_4330 (I76676,I76799,I77064);
not I_4331 (I77232,I3570);
DFFARX1 I_4332 (I1174811,I3563,I77232,I77258,);
not I_4333 (I77266,I77258);
nand I_4334 (I77283,I1174826,I1174805);
and I_4335 (I77300,I77283,I1174808);
DFFARX1 I_4336 (I77300,I3563,I77232,I77326,);
DFFARX1 I_4337 (I1174829,I3563,I77232,I77343,);
and I_4338 (I77351,I77343,I1174808);
nor I_4339 (I77368,I77326,I77351);
DFFARX1 I_4340 (I77368,I3563,I77232,I77200,);
nand I_4341 (I77399,I77343,I1174808);
nand I_4342 (I77416,I77266,I77399);
not I_4343 (I77212,I77416);
DFFARX1 I_4344 (I1174805,I3563,I77232,I77456,);
DFFARX1 I_4345 (I77456,I3563,I77232,I77221,);
nand I_4346 (I77478,I1174817,I1174814);
and I_4347 (I77495,I77478,I1174820);
DFFARX1 I_4348 (I77495,I3563,I77232,I77521,);
DFFARX1 I_4349 (I77521,I3563,I77232,I77538,);
not I_4350 (I77224,I77538);
not I_4351 (I77560,I77521);
nand I_4352 (I77209,I77560,I77399);
nor I_4353 (I77591,I1174823,I1174814);
not I_4354 (I77608,I77591);
nor I_4355 (I77625,I77560,I77608);
nor I_4356 (I77642,I77266,I77625);
DFFARX1 I_4357 (I77642,I3563,I77232,I77218,);
nor I_4358 (I77673,I77326,I77608);
nor I_4359 (I77206,I77521,I77673);
nor I_4360 (I77215,I77456,I77591);
nor I_4361 (I77203,I77326,I77591);
not I_4362 (I77759,I3570);
DFFARX1 I_4363 (I555464,I3563,I77759,I77785,);
not I_4364 (I77793,I77785);
nand I_4365 (I77810,I555485,I555479);
and I_4366 (I77827,I77810,I555461);
DFFARX1 I_4367 (I77827,I3563,I77759,I77853,);
DFFARX1 I_4368 (I555464,I3563,I77759,I77870,);
and I_4369 (I77878,I77870,I555473);
nor I_4370 (I77895,I77853,I77878);
DFFARX1 I_4371 (I77895,I3563,I77759,I77727,);
nand I_4372 (I77926,I77870,I555473);
nand I_4373 (I77943,I77793,I77926);
not I_4374 (I77739,I77943);
DFFARX1 I_4375 (I555470,I3563,I77759,I77983,);
DFFARX1 I_4376 (I77983,I3563,I77759,I77748,);
nand I_4377 (I78005,I555476,I555467);
and I_4378 (I78022,I78005,I555461);
DFFARX1 I_4379 (I78022,I3563,I77759,I78048,);
DFFARX1 I_4380 (I78048,I3563,I77759,I78065,);
not I_4381 (I77751,I78065);
not I_4382 (I78087,I78048);
nand I_4383 (I77736,I78087,I77926);
nor I_4384 (I78118,I555482,I555467);
not I_4385 (I78135,I78118);
nor I_4386 (I78152,I78087,I78135);
nor I_4387 (I78169,I77793,I78152);
DFFARX1 I_4388 (I78169,I3563,I77759,I77745,);
nor I_4389 (I78200,I77853,I78135);
nor I_4390 (I77733,I78048,I78200);
nor I_4391 (I77742,I77983,I78118);
nor I_4392 (I77730,I77853,I78118);
not I_4393 (I78286,I3570);
DFFARX1 I_4394 (I307526,I3563,I78286,I78312,);
not I_4395 (I78320,I78312);
nand I_4396 (I78337,I307508,I307523);
and I_4397 (I78354,I78337,I307499);
DFFARX1 I_4398 (I78354,I3563,I78286,I78380,);
DFFARX1 I_4399 (I307502,I3563,I78286,I78397,);
and I_4400 (I78405,I78397,I307517);
nor I_4401 (I78422,I78380,I78405);
DFFARX1 I_4402 (I78422,I3563,I78286,I78254,);
nand I_4403 (I78453,I78397,I307517);
nand I_4404 (I78470,I78320,I78453);
not I_4405 (I78266,I78470);
DFFARX1 I_4406 (I307520,I3563,I78286,I78510,);
DFFARX1 I_4407 (I78510,I3563,I78286,I78275,);
nand I_4408 (I78532,I307499,I307511);
and I_4409 (I78549,I78532,I307505);
DFFARX1 I_4410 (I78549,I3563,I78286,I78575,);
DFFARX1 I_4411 (I78575,I3563,I78286,I78592,);
not I_4412 (I78278,I78592);
not I_4413 (I78614,I78575);
nand I_4414 (I78263,I78614,I78453);
nor I_4415 (I78645,I307514,I307511);
not I_4416 (I78662,I78645);
nor I_4417 (I78679,I78614,I78662);
nor I_4418 (I78696,I78320,I78679);
DFFARX1 I_4419 (I78696,I3563,I78286,I78272,);
nor I_4420 (I78727,I78380,I78662);
nor I_4421 (I78260,I78575,I78727);
nor I_4422 (I78269,I78510,I78645);
nor I_4423 (I78257,I78380,I78645);
not I_4424 (I78813,I3570);
DFFARX1 I_4425 (I573314,I3563,I78813,I78839,);
not I_4426 (I78847,I78839);
nand I_4427 (I78864,I573335,I573329);
and I_4428 (I78881,I78864,I573311);
DFFARX1 I_4429 (I78881,I3563,I78813,I78907,);
DFFARX1 I_4430 (I573314,I3563,I78813,I78924,);
and I_4431 (I78932,I78924,I573323);
nor I_4432 (I78949,I78907,I78932);
DFFARX1 I_4433 (I78949,I3563,I78813,I78781,);
nand I_4434 (I78980,I78924,I573323);
nand I_4435 (I78997,I78847,I78980);
not I_4436 (I78793,I78997);
DFFARX1 I_4437 (I573320,I3563,I78813,I79037,);
DFFARX1 I_4438 (I79037,I3563,I78813,I78802,);
nand I_4439 (I79059,I573326,I573317);
and I_4440 (I79076,I79059,I573311);
DFFARX1 I_4441 (I79076,I3563,I78813,I79102,);
DFFARX1 I_4442 (I79102,I3563,I78813,I79119,);
not I_4443 (I78805,I79119);
not I_4444 (I79141,I79102);
nand I_4445 (I78790,I79141,I78980);
nor I_4446 (I79172,I573332,I573317);
not I_4447 (I79189,I79172);
nor I_4448 (I79206,I79141,I79189);
nor I_4449 (I79223,I78847,I79206);
DFFARX1 I_4450 (I79223,I3563,I78813,I78799,);
nor I_4451 (I79254,I78907,I79189);
nor I_4452 (I78787,I79102,I79254);
nor I_4453 (I78796,I79037,I79172);
nor I_4454 (I78784,I78907,I79172);
not I_4455 (I79340,I3570);
DFFARX1 I_4456 (I994988,I3563,I79340,I79366,);
not I_4457 (I79374,I79366);
nand I_4458 (I79391,I995006,I995000);
and I_4459 (I79408,I79391,I994979);
DFFARX1 I_4460 (I79408,I3563,I79340,I79434,);
DFFARX1 I_4461 (I994997,I3563,I79340,I79451,);
and I_4462 (I79459,I79451,I994982);
nor I_4463 (I79476,I79434,I79459);
DFFARX1 I_4464 (I79476,I3563,I79340,I79308,);
nand I_4465 (I79507,I79451,I994982);
nand I_4466 (I79524,I79374,I79507);
not I_4467 (I79320,I79524);
DFFARX1 I_4468 (I994994,I3563,I79340,I79564,);
DFFARX1 I_4469 (I79564,I3563,I79340,I79329,);
nand I_4470 (I79586,I995003,I994991);
and I_4471 (I79603,I79586,I994985);
DFFARX1 I_4472 (I79603,I3563,I79340,I79629,);
DFFARX1 I_4473 (I79629,I3563,I79340,I79646,);
not I_4474 (I79332,I79646);
not I_4475 (I79668,I79629);
nand I_4476 (I79317,I79668,I79507);
nor I_4477 (I79699,I994979,I994991);
not I_4478 (I79716,I79699);
nor I_4479 (I79733,I79668,I79716);
nor I_4480 (I79750,I79374,I79733);
DFFARX1 I_4481 (I79750,I3563,I79340,I79326,);
nor I_4482 (I79781,I79434,I79716);
nor I_4483 (I79314,I79629,I79781);
nor I_4484 (I79323,I79564,I79699);
nor I_4485 (I79311,I79434,I79699);
not I_4486 (I79867,I3570);
DFFARX1 I_4487 (I336511,I3563,I79867,I79893,);
not I_4488 (I79901,I79893);
nand I_4489 (I79918,I336493,I336508);
and I_4490 (I79935,I79918,I336484);
DFFARX1 I_4491 (I79935,I3563,I79867,I79961,);
DFFARX1 I_4492 (I336487,I3563,I79867,I79978,);
and I_4493 (I79986,I79978,I336502);
nor I_4494 (I80003,I79961,I79986);
DFFARX1 I_4495 (I80003,I3563,I79867,I79835,);
nand I_4496 (I80034,I79978,I336502);
nand I_4497 (I80051,I79901,I80034);
not I_4498 (I79847,I80051);
DFFARX1 I_4499 (I336505,I3563,I79867,I80091,);
DFFARX1 I_4500 (I80091,I3563,I79867,I79856,);
nand I_4501 (I80113,I336484,I336496);
and I_4502 (I80130,I80113,I336490);
DFFARX1 I_4503 (I80130,I3563,I79867,I80156,);
DFFARX1 I_4504 (I80156,I3563,I79867,I80173,);
not I_4505 (I79859,I80173);
not I_4506 (I80195,I80156);
nand I_4507 (I79844,I80195,I80034);
nor I_4508 (I80226,I336499,I336496);
not I_4509 (I80243,I80226);
nor I_4510 (I80260,I80195,I80243);
nor I_4511 (I80277,I79901,I80260);
DFFARX1 I_4512 (I80277,I3563,I79867,I79853,);
nor I_4513 (I80308,I79961,I80243);
nor I_4514 (I79841,I80156,I80308);
nor I_4515 (I79850,I80091,I80226);
nor I_4516 (I79838,I79961,I80226);
not I_4517 (I80394,I3570);
DFFARX1 I_4518 (I788475,I3563,I80394,I80420,);
not I_4519 (I80428,I80420);
nand I_4520 (I80445,I788466,I788484);
and I_4521 (I80462,I80445,I788463);
DFFARX1 I_4522 (I80462,I3563,I80394,I80488,);
DFFARX1 I_4523 (I788466,I3563,I80394,I80505,);
and I_4524 (I80513,I80505,I788469);
nor I_4525 (I80530,I80488,I80513);
DFFARX1 I_4526 (I80530,I3563,I80394,I80362,);
nand I_4527 (I80561,I80505,I788469);
nand I_4528 (I80578,I80428,I80561);
not I_4529 (I80374,I80578);
DFFARX1 I_4530 (I788463,I3563,I80394,I80618,);
DFFARX1 I_4531 (I80618,I3563,I80394,I80383,);
nand I_4532 (I80640,I788481,I788472);
and I_4533 (I80657,I80640,I788487);
DFFARX1 I_4534 (I80657,I3563,I80394,I80683,);
DFFARX1 I_4535 (I80683,I3563,I80394,I80700,);
not I_4536 (I80386,I80700);
not I_4537 (I80722,I80683);
nand I_4538 (I80371,I80722,I80561);
nor I_4539 (I80753,I788478,I788472);
not I_4540 (I80770,I80753);
nor I_4541 (I80787,I80722,I80770);
nor I_4542 (I80804,I80428,I80787);
DFFARX1 I_4543 (I80804,I3563,I80394,I80380,);
nor I_4544 (I80835,I80488,I80770);
nor I_4545 (I80368,I80683,I80835);
nor I_4546 (I80377,I80618,I80753);
nor I_4547 (I80365,I80488,I80753);
not I_4548 (I80921,I3570);
DFFARX1 I_4549 (I176220,I3563,I80921,I80947,);
not I_4550 (I80955,I80947);
nand I_4551 (I80972,I176214,I176208);
and I_4552 (I80989,I80972,I176229);
DFFARX1 I_4553 (I80989,I3563,I80921,I81015,);
DFFARX1 I_4554 (I176226,I3563,I80921,I81032,);
and I_4555 (I81040,I81032,I176223);
nor I_4556 (I81057,I81015,I81040);
DFFARX1 I_4557 (I81057,I3563,I80921,I80889,);
nand I_4558 (I81088,I81032,I176223);
nand I_4559 (I81105,I80955,I81088);
not I_4560 (I80901,I81105);
DFFARX1 I_4561 (I176208,I3563,I80921,I81145,);
DFFARX1 I_4562 (I81145,I3563,I80921,I80910,);
nand I_4563 (I81167,I176211,I176211);
and I_4564 (I81184,I81167,I176232);
DFFARX1 I_4565 (I81184,I3563,I80921,I81210,);
DFFARX1 I_4566 (I81210,I3563,I80921,I81227,);
not I_4567 (I80913,I81227);
not I_4568 (I81249,I81210);
nand I_4569 (I80898,I81249,I81088);
nor I_4570 (I81280,I176217,I176211);
not I_4571 (I81297,I81280);
nor I_4572 (I81314,I81249,I81297);
nor I_4573 (I81331,I80955,I81314);
DFFARX1 I_4574 (I81331,I3563,I80921,I80907,);
nor I_4575 (I81362,I81015,I81297);
nor I_4576 (I80895,I81210,I81362);
nor I_4577 (I80904,I81145,I81280);
nor I_4578 (I80892,I81015,I81280);
not I_4579 (I81448,I3570);
DFFARX1 I_4580 (I705243,I3563,I81448,I81474,);
not I_4581 (I81482,I81474);
nand I_4582 (I81499,I705234,I705252);
and I_4583 (I81516,I81499,I705231);
DFFARX1 I_4584 (I81516,I3563,I81448,I81542,);
DFFARX1 I_4585 (I705234,I3563,I81448,I81559,);
and I_4586 (I81567,I81559,I705237);
nor I_4587 (I81584,I81542,I81567);
DFFARX1 I_4588 (I81584,I3563,I81448,I81416,);
nand I_4589 (I81615,I81559,I705237);
nand I_4590 (I81632,I81482,I81615);
not I_4591 (I81428,I81632);
DFFARX1 I_4592 (I705231,I3563,I81448,I81672,);
DFFARX1 I_4593 (I81672,I3563,I81448,I81437,);
nand I_4594 (I81694,I705249,I705240);
and I_4595 (I81711,I81694,I705255);
DFFARX1 I_4596 (I81711,I3563,I81448,I81737,);
DFFARX1 I_4597 (I81737,I3563,I81448,I81754,);
not I_4598 (I81440,I81754);
not I_4599 (I81776,I81737);
nand I_4600 (I81425,I81776,I81615);
nor I_4601 (I81807,I705246,I705240);
not I_4602 (I81824,I81807);
nor I_4603 (I81841,I81776,I81824);
nor I_4604 (I81858,I81482,I81841);
DFFARX1 I_4605 (I81858,I3563,I81448,I81434,);
nor I_4606 (I81889,I81542,I81824);
nor I_4607 (I81422,I81737,I81889);
nor I_4608 (I81431,I81672,I81807);
nor I_4609 (I81419,I81542,I81807);
not I_4610 (I81975,I3570);
DFFARX1 I_4611 (I556059,I3563,I81975,I82001,);
not I_4612 (I82009,I82001);
nand I_4613 (I82026,I556080,I556074);
and I_4614 (I82043,I82026,I556056);
DFFARX1 I_4615 (I82043,I3563,I81975,I82069,);
DFFARX1 I_4616 (I556059,I3563,I81975,I82086,);
and I_4617 (I82094,I82086,I556068);
nor I_4618 (I82111,I82069,I82094);
DFFARX1 I_4619 (I82111,I3563,I81975,I81943,);
nand I_4620 (I82142,I82086,I556068);
nand I_4621 (I82159,I82009,I82142);
not I_4622 (I81955,I82159);
DFFARX1 I_4623 (I556065,I3563,I81975,I82199,);
DFFARX1 I_4624 (I82199,I3563,I81975,I81964,);
nand I_4625 (I82221,I556071,I556062);
and I_4626 (I82238,I82221,I556056);
DFFARX1 I_4627 (I82238,I3563,I81975,I82264,);
DFFARX1 I_4628 (I82264,I3563,I81975,I82281,);
not I_4629 (I81967,I82281);
not I_4630 (I82303,I82264);
nand I_4631 (I81952,I82303,I82142);
nor I_4632 (I82334,I556077,I556062);
not I_4633 (I82351,I82334);
nor I_4634 (I82368,I82303,I82351);
nor I_4635 (I82385,I82009,I82368);
DFFARX1 I_4636 (I82385,I3563,I81975,I81961,);
nor I_4637 (I82416,I82069,I82351);
nor I_4638 (I81949,I82264,I82416);
nor I_4639 (I81958,I82199,I82334);
nor I_4640 (I81946,I82069,I82334);
not I_4641 (I82502,I3570);
DFFARX1 I_4642 (I342308,I3563,I82502,I82528,);
not I_4643 (I82536,I82528);
nand I_4644 (I82553,I342290,I342305);
and I_4645 (I82570,I82553,I342281);
DFFARX1 I_4646 (I82570,I3563,I82502,I82596,);
DFFARX1 I_4647 (I342284,I3563,I82502,I82613,);
and I_4648 (I82621,I82613,I342299);
nor I_4649 (I82638,I82596,I82621);
DFFARX1 I_4650 (I82638,I3563,I82502,I82470,);
nand I_4651 (I82669,I82613,I342299);
nand I_4652 (I82686,I82536,I82669);
not I_4653 (I82482,I82686);
DFFARX1 I_4654 (I342302,I3563,I82502,I82726,);
DFFARX1 I_4655 (I82726,I3563,I82502,I82491,);
nand I_4656 (I82748,I342281,I342293);
and I_4657 (I82765,I82748,I342287);
DFFARX1 I_4658 (I82765,I3563,I82502,I82791,);
DFFARX1 I_4659 (I82791,I3563,I82502,I82808,);
not I_4660 (I82494,I82808);
not I_4661 (I82830,I82791);
nand I_4662 (I82479,I82830,I82669);
nor I_4663 (I82861,I342296,I342293);
not I_4664 (I82878,I82861);
nor I_4665 (I82895,I82830,I82878);
nor I_4666 (I82912,I82536,I82895);
DFFARX1 I_4667 (I82912,I3563,I82502,I82488,);
nor I_4668 (I82943,I82596,I82878);
nor I_4669 (I82476,I82791,I82943);
nor I_4670 (I82485,I82726,I82861);
nor I_4671 (I82473,I82596,I82861);
not I_4672 (I83029,I3570);
DFFARX1 I_4673 (I858495,I3563,I83029,I83055,);
not I_4674 (I83063,I83055);
nand I_4675 (I83080,I858492,I858507);
and I_4676 (I83097,I83080,I858489);
DFFARX1 I_4677 (I83097,I3563,I83029,I83123,);
DFFARX1 I_4678 (I858486,I3563,I83029,I83140,);
and I_4679 (I83148,I83140,I858486);
nor I_4680 (I83165,I83123,I83148);
DFFARX1 I_4681 (I83165,I3563,I83029,I82997,);
nand I_4682 (I83196,I83140,I858486);
nand I_4683 (I83213,I83063,I83196);
not I_4684 (I83009,I83213);
DFFARX1 I_4685 (I858489,I3563,I83029,I83253,);
DFFARX1 I_4686 (I83253,I3563,I83029,I83018,);
nand I_4687 (I83275,I858501,I858492);
and I_4688 (I83292,I83275,I858504);
DFFARX1 I_4689 (I83292,I3563,I83029,I83318,);
DFFARX1 I_4690 (I83318,I3563,I83029,I83335,);
not I_4691 (I83021,I83335);
not I_4692 (I83357,I83318);
nand I_4693 (I83006,I83357,I83196);
nor I_4694 (I83388,I858498,I858492);
not I_4695 (I83405,I83388);
nor I_4696 (I83422,I83357,I83405);
nor I_4697 (I83439,I83063,I83422);
DFFARX1 I_4698 (I83439,I3563,I83029,I83015,);
nor I_4699 (I83470,I83123,I83405);
nor I_4700 (I83003,I83318,I83470);
nor I_4701 (I83012,I83253,I83388);
nor I_4702 (I83000,I83123,I83388);
not I_4703 (I83556,I3570);
DFFARX1 I_4704 (I624898,I3563,I83556,I83582,);
not I_4705 (I83590,I83582);
nand I_4706 (I83607,I624910,I624895);
and I_4707 (I83624,I83607,I624889);
DFFARX1 I_4708 (I83624,I3563,I83556,I83650,);
DFFARX1 I_4709 (I624904,I3563,I83556,I83667,);
and I_4710 (I83675,I83667,I624892);
nor I_4711 (I83692,I83650,I83675);
DFFARX1 I_4712 (I83692,I3563,I83556,I83524,);
nand I_4713 (I83723,I83667,I624892);
nand I_4714 (I83740,I83590,I83723);
not I_4715 (I83536,I83740);
DFFARX1 I_4716 (I624901,I3563,I83556,I83780,);
DFFARX1 I_4717 (I83780,I3563,I83556,I83545,);
nand I_4718 (I83802,I624907,I624913);
and I_4719 (I83819,I83802,I624889);
DFFARX1 I_4720 (I83819,I3563,I83556,I83845,);
DFFARX1 I_4721 (I83845,I3563,I83556,I83862,);
not I_4722 (I83548,I83862);
not I_4723 (I83884,I83845);
nand I_4724 (I83533,I83884,I83723);
nor I_4725 (I83915,I624892,I624913);
not I_4726 (I83932,I83915);
nor I_4727 (I83949,I83884,I83932);
nor I_4728 (I83966,I83590,I83949);
DFFARX1 I_4729 (I83966,I3563,I83556,I83542,);
nor I_4730 (I83997,I83650,I83932);
nor I_4731 (I83530,I83845,I83997);
nor I_4732 (I83539,I83780,I83915);
nor I_4733 (I83527,I83650,I83915);
not I_4734 (I84083,I3570);
DFFARX1 I_4735 (I1347010,I3563,I84083,I84109,);
not I_4736 (I84117,I84109);
nand I_4737 (I84134,I1347004,I1347025);
and I_4738 (I84151,I84134,I1347001);
DFFARX1 I_4739 (I84151,I3563,I84083,I84177,);
DFFARX1 I_4740 (I1347022,I3563,I84083,I84194,);
and I_4741 (I84202,I84194,I1347019);
nor I_4742 (I84219,I84177,I84202);
DFFARX1 I_4743 (I84219,I3563,I84083,I84051,);
nand I_4744 (I84250,I84194,I1347019);
nand I_4745 (I84267,I84117,I84250);
not I_4746 (I84063,I84267);
DFFARX1 I_4747 (I1347007,I3563,I84083,I84307,);
DFFARX1 I_4748 (I84307,I3563,I84083,I84072,);
nand I_4749 (I84329,I1347016,I1347013);
and I_4750 (I84346,I84329,I1346998);
DFFARX1 I_4751 (I84346,I3563,I84083,I84372,);
DFFARX1 I_4752 (I84372,I3563,I84083,I84389,);
not I_4753 (I84075,I84389);
not I_4754 (I84411,I84372);
nand I_4755 (I84060,I84411,I84250);
nor I_4756 (I84442,I1346998,I1347013);
not I_4757 (I84459,I84442);
nor I_4758 (I84476,I84411,I84459);
nor I_4759 (I84493,I84117,I84476);
DFFARX1 I_4760 (I84493,I3563,I84083,I84069,);
nor I_4761 (I84524,I84177,I84459);
nor I_4762 (I84057,I84372,I84524);
nor I_4763 (I84066,I84307,I84442);
nor I_4764 (I84054,I84177,I84442);
not I_4765 (I84610,I3570);
DFFARX1 I_4766 (I205970,I3563,I84610,I84636,);
not I_4767 (I84644,I84636);
nand I_4768 (I84661,I205964,I205958);
and I_4769 (I84678,I84661,I205979);
DFFARX1 I_4770 (I84678,I3563,I84610,I84704,);
DFFARX1 I_4771 (I205976,I3563,I84610,I84721,);
and I_4772 (I84729,I84721,I205973);
nor I_4773 (I84746,I84704,I84729);
DFFARX1 I_4774 (I84746,I3563,I84610,I84578,);
nand I_4775 (I84777,I84721,I205973);
nand I_4776 (I84794,I84644,I84777);
not I_4777 (I84590,I84794);
DFFARX1 I_4778 (I205958,I3563,I84610,I84834,);
DFFARX1 I_4779 (I84834,I3563,I84610,I84599,);
nand I_4780 (I84856,I205961,I205961);
and I_4781 (I84873,I84856,I205982);
DFFARX1 I_4782 (I84873,I3563,I84610,I84899,);
DFFARX1 I_4783 (I84899,I3563,I84610,I84916,);
not I_4784 (I84602,I84916);
not I_4785 (I84938,I84899);
nand I_4786 (I84587,I84938,I84777);
nor I_4787 (I84969,I205967,I205961);
not I_4788 (I84986,I84969);
nor I_4789 (I85003,I84938,I84986);
nor I_4790 (I85020,I84644,I85003);
DFFARX1 I_4791 (I85020,I3563,I84610,I84596,);
nor I_4792 (I85051,I84704,I84986);
nor I_4793 (I84584,I84899,I85051);
nor I_4794 (I84593,I84834,I84969);
nor I_4795 (I84581,I84704,I84969);
not I_4796 (I85137,I3570);
DFFARX1 I_4797 (I1204867,I3563,I85137,I85163,);
not I_4798 (I85171,I85163);
nand I_4799 (I85188,I1204882,I1204861);
and I_4800 (I85205,I85188,I1204864);
DFFARX1 I_4801 (I85205,I3563,I85137,I85231,);
DFFARX1 I_4802 (I1204885,I3563,I85137,I85248,);
and I_4803 (I85256,I85248,I1204864);
nor I_4804 (I85273,I85231,I85256);
DFFARX1 I_4805 (I85273,I3563,I85137,I85105,);
nand I_4806 (I85304,I85248,I1204864);
nand I_4807 (I85321,I85171,I85304);
not I_4808 (I85117,I85321);
DFFARX1 I_4809 (I1204861,I3563,I85137,I85361,);
DFFARX1 I_4810 (I85361,I3563,I85137,I85126,);
nand I_4811 (I85383,I1204873,I1204870);
and I_4812 (I85400,I85383,I1204876);
DFFARX1 I_4813 (I85400,I3563,I85137,I85426,);
DFFARX1 I_4814 (I85426,I3563,I85137,I85443,);
not I_4815 (I85129,I85443);
not I_4816 (I85465,I85426);
nand I_4817 (I85114,I85465,I85304);
nor I_4818 (I85496,I1204879,I1204870);
not I_4819 (I85513,I85496);
nor I_4820 (I85530,I85465,I85513);
nor I_4821 (I85547,I85171,I85530);
DFFARX1 I_4822 (I85547,I3563,I85137,I85123,);
nor I_4823 (I85578,I85231,I85513);
nor I_4824 (I85111,I85426,I85578);
nor I_4825 (I85120,I85361,I85496);
nor I_4826 (I85108,I85231,I85496);
not I_4827 (I85664,I3570);
DFFARX1 I_4828 (I755529,I3563,I85664,I85690,);
not I_4829 (I85698,I85690);
nand I_4830 (I85715,I755520,I755538);
and I_4831 (I85732,I85715,I755517);
DFFARX1 I_4832 (I85732,I3563,I85664,I85758,);
DFFARX1 I_4833 (I755520,I3563,I85664,I85775,);
and I_4834 (I85783,I85775,I755523);
nor I_4835 (I85800,I85758,I85783);
DFFARX1 I_4836 (I85800,I3563,I85664,I85632,);
nand I_4837 (I85831,I85775,I755523);
nand I_4838 (I85848,I85698,I85831);
not I_4839 (I85644,I85848);
DFFARX1 I_4840 (I755517,I3563,I85664,I85888,);
DFFARX1 I_4841 (I85888,I3563,I85664,I85653,);
nand I_4842 (I85910,I755535,I755526);
and I_4843 (I85927,I85910,I755541);
DFFARX1 I_4844 (I85927,I3563,I85664,I85953,);
DFFARX1 I_4845 (I85953,I3563,I85664,I85970,);
not I_4846 (I85656,I85970);
not I_4847 (I85992,I85953);
nand I_4848 (I85641,I85992,I85831);
nor I_4849 (I86023,I755532,I755526);
not I_4850 (I86040,I86023);
nor I_4851 (I86057,I85992,I86040);
nor I_4852 (I86074,I85698,I86057);
DFFARX1 I_4853 (I86074,I3563,I85664,I85650,);
nor I_4854 (I86105,I85758,I86040);
nor I_4855 (I85638,I85953,I86105);
nor I_4856 (I85647,I85888,I86023);
nor I_4857 (I85635,I85758,I86023);
not I_4858 (I86191,I3570);
DFFARX1 I_4859 (I1189261,I3563,I86191,I86217,);
not I_4860 (I86225,I86217);
nand I_4861 (I86242,I1189276,I1189255);
and I_4862 (I86259,I86242,I1189258);
DFFARX1 I_4863 (I86259,I3563,I86191,I86285,);
DFFARX1 I_4864 (I1189279,I3563,I86191,I86302,);
and I_4865 (I86310,I86302,I1189258);
nor I_4866 (I86327,I86285,I86310);
DFFARX1 I_4867 (I86327,I3563,I86191,I86159,);
nand I_4868 (I86358,I86302,I1189258);
nand I_4869 (I86375,I86225,I86358);
not I_4870 (I86171,I86375);
DFFARX1 I_4871 (I1189255,I3563,I86191,I86415,);
DFFARX1 I_4872 (I86415,I3563,I86191,I86180,);
nand I_4873 (I86437,I1189267,I1189264);
and I_4874 (I86454,I86437,I1189270);
DFFARX1 I_4875 (I86454,I3563,I86191,I86480,);
DFFARX1 I_4876 (I86480,I3563,I86191,I86497,);
not I_4877 (I86183,I86497);
not I_4878 (I86519,I86480);
nand I_4879 (I86168,I86519,I86358);
nor I_4880 (I86550,I1189273,I1189264);
not I_4881 (I86567,I86550);
nor I_4882 (I86584,I86519,I86567);
nor I_4883 (I86601,I86225,I86584);
DFFARX1 I_4884 (I86601,I3563,I86191,I86177,);
nor I_4885 (I86632,I86285,I86567);
nor I_4886 (I86165,I86480,I86632);
nor I_4887 (I86174,I86415,I86550);
nor I_4888 (I86162,I86285,I86550);
not I_4889 (I86718,I3570);
DFFARX1 I_4890 (I1088176,I3563,I86718,I86744,);
not I_4891 (I86752,I86744);
nand I_4892 (I86769,I1088173,I1088179);
and I_4893 (I86786,I86769,I1088176);
DFFARX1 I_4894 (I86786,I3563,I86718,I86812,);
DFFARX1 I_4895 (I1088179,I3563,I86718,I86829,);
and I_4896 (I86837,I86829,I1088173);
nor I_4897 (I86854,I86812,I86837);
DFFARX1 I_4898 (I86854,I3563,I86718,I86686,);
nand I_4899 (I86885,I86829,I1088173);
nand I_4900 (I86902,I86752,I86885);
not I_4901 (I86698,I86902);
DFFARX1 I_4902 (I1088182,I3563,I86718,I86942,);
DFFARX1 I_4903 (I86942,I3563,I86718,I86707,);
nand I_4904 (I86964,I1088185,I1088194);
and I_4905 (I86981,I86964,I1088188);
DFFARX1 I_4906 (I86981,I3563,I86718,I87007,);
DFFARX1 I_4907 (I87007,I3563,I86718,I87024,);
not I_4908 (I86710,I87024);
not I_4909 (I87046,I87007);
nand I_4910 (I86695,I87046,I86885);
nor I_4911 (I87077,I1088191,I1088194);
not I_4912 (I87094,I87077);
nor I_4913 (I87111,I87046,I87094);
nor I_4914 (I87128,I86752,I87111);
DFFARX1 I_4915 (I87128,I3563,I86718,I86704,);
nor I_4916 (I87159,I86812,I87094);
nor I_4917 (I86692,I87007,I87159);
nor I_4918 (I86701,I86942,I87077);
nor I_4919 (I86689,I86812,I87077);
not I_4920 (I87245,I3570);
DFFARX1 I_4921 (I446900,I3563,I87245,I87271,);
not I_4922 (I87279,I87271);
nand I_4923 (I87296,I446894,I446885);
and I_4924 (I87313,I87296,I446906);
DFFARX1 I_4925 (I87313,I3563,I87245,I87339,);
DFFARX1 I_4926 (I446888,I3563,I87245,I87356,);
and I_4927 (I87364,I87356,I446882);
nor I_4928 (I87381,I87339,I87364);
DFFARX1 I_4929 (I87381,I3563,I87245,I87213,);
nand I_4930 (I87412,I87356,I446882);
nand I_4931 (I87429,I87279,I87412);
not I_4932 (I87225,I87429);
DFFARX1 I_4933 (I446882,I3563,I87245,I87469,);
DFFARX1 I_4934 (I87469,I3563,I87245,I87234,);
nand I_4935 (I87491,I446909,I446891);
and I_4936 (I87508,I87491,I446897);
DFFARX1 I_4937 (I87508,I3563,I87245,I87534,);
DFFARX1 I_4938 (I87534,I3563,I87245,I87551,);
not I_4939 (I87237,I87551);
not I_4940 (I87573,I87534);
nand I_4941 (I87222,I87573,I87412);
nor I_4942 (I87604,I446903,I446891);
not I_4943 (I87621,I87604);
nor I_4944 (I87638,I87573,I87621);
nor I_4945 (I87655,I87279,I87638);
DFFARX1 I_4946 (I87655,I3563,I87245,I87231,);
nor I_4947 (I87686,I87339,I87621);
nor I_4948 (I87219,I87534,I87686);
nor I_4949 (I87228,I87469,I87604);
nor I_4950 (I87216,I87339,I87604);
not I_4951 (I87772,I3570);
DFFARX1 I_4952 (I468660,I3563,I87772,I87798,);
not I_4953 (I87806,I87798);
nand I_4954 (I87823,I468654,I468645);
and I_4955 (I87840,I87823,I468666);
DFFARX1 I_4956 (I87840,I3563,I87772,I87866,);
DFFARX1 I_4957 (I468648,I3563,I87772,I87883,);
and I_4958 (I87891,I87883,I468642);
nor I_4959 (I87908,I87866,I87891);
DFFARX1 I_4960 (I87908,I3563,I87772,I87740,);
nand I_4961 (I87939,I87883,I468642);
nand I_4962 (I87956,I87806,I87939);
not I_4963 (I87752,I87956);
DFFARX1 I_4964 (I468642,I3563,I87772,I87996,);
DFFARX1 I_4965 (I87996,I3563,I87772,I87761,);
nand I_4966 (I88018,I468669,I468651);
and I_4967 (I88035,I88018,I468657);
DFFARX1 I_4968 (I88035,I3563,I87772,I88061,);
DFFARX1 I_4969 (I88061,I3563,I87772,I88078,);
not I_4970 (I87764,I88078);
not I_4971 (I88100,I88061);
nand I_4972 (I87749,I88100,I87939);
nor I_4973 (I88131,I468663,I468651);
not I_4974 (I88148,I88131);
nor I_4975 (I88165,I88100,I88148);
nor I_4976 (I88182,I87806,I88165);
DFFARX1 I_4977 (I88182,I3563,I87772,I87758,);
nor I_4978 (I88213,I87866,I88148);
nor I_4979 (I87746,I88061,I88213);
nor I_4980 (I87755,I87996,I88131);
nor I_4981 (I87743,I87866,I88131);
not I_4982 (I88299,I3570);
DFFARX1 I_4983 (I803503,I3563,I88299,I88325,);
not I_4984 (I88333,I88325);
nand I_4985 (I88350,I803494,I803512);
and I_4986 (I88367,I88350,I803491);
DFFARX1 I_4987 (I88367,I3563,I88299,I88393,);
DFFARX1 I_4988 (I803494,I3563,I88299,I88410,);
and I_4989 (I88418,I88410,I803497);
nor I_4990 (I88435,I88393,I88418);
DFFARX1 I_4991 (I88435,I3563,I88299,I88267,);
nand I_4992 (I88466,I88410,I803497);
nand I_4993 (I88483,I88333,I88466);
not I_4994 (I88279,I88483);
DFFARX1 I_4995 (I803491,I3563,I88299,I88523,);
DFFARX1 I_4996 (I88523,I3563,I88299,I88288,);
nand I_4997 (I88545,I803509,I803500);
and I_4998 (I88562,I88545,I803515);
DFFARX1 I_4999 (I88562,I3563,I88299,I88588,);
DFFARX1 I_5000 (I88588,I3563,I88299,I88605,);
not I_5001 (I88291,I88605);
not I_5002 (I88627,I88588);
nand I_5003 (I88276,I88627,I88466);
nor I_5004 (I88658,I803506,I803500);
not I_5005 (I88675,I88658);
nor I_5006 (I88692,I88627,I88675);
nor I_5007 (I88709,I88333,I88692);
DFFARX1 I_5008 (I88709,I3563,I88299,I88285,);
nor I_5009 (I88740,I88393,I88675);
nor I_5010 (I88273,I88588,I88740);
nor I_5011 (I88282,I88523,I88658);
nor I_5012 (I88270,I88393,I88658);
not I_5013 (I88826,I3570);
DFFARX1 I_5014 (I364442,I3563,I88826,I88852,);
not I_5015 (I88860,I88852);
nand I_5016 (I88877,I364424,I364439);
and I_5017 (I88894,I88877,I364415);
DFFARX1 I_5018 (I88894,I3563,I88826,I88920,);
DFFARX1 I_5019 (I364418,I3563,I88826,I88937,);
and I_5020 (I88945,I88937,I364433);
nor I_5021 (I88962,I88920,I88945);
DFFARX1 I_5022 (I88962,I3563,I88826,I88794,);
nand I_5023 (I88993,I88937,I364433);
nand I_5024 (I89010,I88860,I88993);
not I_5025 (I88806,I89010);
DFFARX1 I_5026 (I364436,I3563,I88826,I89050,);
DFFARX1 I_5027 (I89050,I3563,I88826,I88815,);
nand I_5028 (I89072,I364415,I364427);
and I_5029 (I89089,I89072,I364421);
DFFARX1 I_5030 (I89089,I3563,I88826,I89115,);
DFFARX1 I_5031 (I89115,I3563,I88826,I89132,);
not I_5032 (I88818,I89132);
not I_5033 (I89154,I89115);
nand I_5034 (I88803,I89154,I88993);
nor I_5035 (I89185,I364430,I364427);
not I_5036 (I89202,I89185);
nor I_5037 (I89219,I89154,I89202);
nor I_5038 (I89236,I88860,I89219);
DFFARX1 I_5039 (I89236,I3563,I88826,I88812,);
nor I_5040 (I89267,I88920,I89202);
nor I_5041 (I88800,I89115,I89267);
nor I_5042 (I88809,I89050,I89185);
nor I_5043 (I88797,I88920,I89185);
not I_5044 (I89353,I3570);
DFFARX1 I_5045 (I38753,I3563,I89353,I89379,);
not I_5046 (I89387,I89379);
nand I_5047 (I89404,I38741,I38747);
and I_5048 (I89421,I89404,I38750);
DFFARX1 I_5049 (I89421,I3563,I89353,I89447,);
DFFARX1 I_5050 (I38732,I3563,I89353,I89464,);
and I_5051 (I89472,I89464,I38738);
nor I_5052 (I89489,I89447,I89472);
DFFARX1 I_5053 (I89489,I3563,I89353,I89321,);
nand I_5054 (I89520,I89464,I38738);
nand I_5055 (I89537,I89387,I89520);
not I_5056 (I89333,I89537);
DFFARX1 I_5057 (I38732,I3563,I89353,I89577,);
DFFARX1 I_5058 (I89577,I3563,I89353,I89342,);
nand I_5059 (I89599,I38735,I38729);
and I_5060 (I89616,I89599,I38744);
DFFARX1 I_5061 (I89616,I3563,I89353,I89642,);
DFFARX1 I_5062 (I89642,I3563,I89353,I89659,);
not I_5063 (I89345,I89659);
not I_5064 (I89681,I89642);
nand I_5065 (I89330,I89681,I89520);
nor I_5066 (I89712,I38729,I38729);
not I_5067 (I89729,I89712);
nor I_5068 (I89746,I89681,I89729);
nor I_5069 (I89763,I89387,I89746);
DFFARX1 I_5070 (I89763,I3563,I89353,I89339,);
nor I_5071 (I89794,I89447,I89729);
nor I_5072 (I89327,I89642,I89794);
nor I_5073 (I89336,I89577,I89712);
nor I_5074 (I89324,I89447,I89712);
not I_5075 (I89880,I3570);
DFFARX1 I_5076 (I749171,I3563,I89880,I89906,);
not I_5077 (I89914,I89906);
nand I_5078 (I89931,I749162,I749180);
and I_5079 (I89948,I89931,I749159);
DFFARX1 I_5080 (I89948,I3563,I89880,I89974,);
DFFARX1 I_5081 (I749162,I3563,I89880,I89991,);
and I_5082 (I89999,I89991,I749165);
nor I_5083 (I90016,I89974,I89999);
DFFARX1 I_5084 (I90016,I3563,I89880,I89848,);
nand I_5085 (I90047,I89991,I749165);
nand I_5086 (I90064,I89914,I90047);
not I_5087 (I89860,I90064);
DFFARX1 I_5088 (I749159,I3563,I89880,I90104,);
DFFARX1 I_5089 (I90104,I3563,I89880,I89869,);
nand I_5090 (I90126,I749177,I749168);
and I_5091 (I90143,I90126,I749183);
DFFARX1 I_5092 (I90143,I3563,I89880,I90169,);
DFFARX1 I_5093 (I90169,I3563,I89880,I90186,);
not I_5094 (I89872,I90186);
not I_5095 (I90208,I90169);
nand I_5096 (I89857,I90208,I90047);
nor I_5097 (I90239,I749174,I749168);
not I_5098 (I90256,I90239);
nor I_5099 (I90273,I90208,I90256);
nor I_5100 (I90290,I89914,I90273);
DFFARX1 I_5101 (I90290,I3563,I89880,I89866,);
nor I_5102 (I90321,I89974,I90256);
nor I_5103 (I89854,I90169,I90321);
nor I_5104 (I89863,I90104,I90239);
nor I_5105 (I89851,I89974,I90239);
not I_5106 (I90407,I3570);
DFFARX1 I_5107 (I257735,I3563,I90407,I90433,);
not I_5108 (I90441,I90433);
nand I_5109 (I90458,I257729,I257723);
and I_5110 (I90475,I90458,I257744);
DFFARX1 I_5111 (I90475,I3563,I90407,I90501,);
DFFARX1 I_5112 (I257741,I3563,I90407,I90518,);
and I_5113 (I90526,I90518,I257738);
nor I_5114 (I90543,I90501,I90526);
DFFARX1 I_5115 (I90543,I3563,I90407,I90375,);
nand I_5116 (I90574,I90518,I257738);
nand I_5117 (I90591,I90441,I90574);
not I_5118 (I90387,I90591);
DFFARX1 I_5119 (I257723,I3563,I90407,I90631,);
DFFARX1 I_5120 (I90631,I3563,I90407,I90396,);
nand I_5121 (I90653,I257726,I257726);
and I_5122 (I90670,I90653,I257747);
DFFARX1 I_5123 (I90670,I3563,I90407,I90696,);
DFFARX1 I_5124 (I90696,I3563,I90407,I90713,);
not I_5125 (I90399,I90713);
not I_5126 (I90735,I90696);
nand I_5127 (I90384,I90735,I90574);
nor I_5128 (I90766,I257732,I257726);
not I_5129 (I90783,I90766);
nor I_5130 (I90800,I90735,I90783);
nor I_5131 (I90817,I90441,I90800);
DFFARX1 I_5132 (I90817,I3563,I90407,I90393,);
nor I_5133 (I90848,I90501,I90783);
nor I_5134 (I90381,I90696,I90848);
nor I_5135 (I90390,I90631,I90766);
nor I_5136 (I90378,I90501,I90766);
not I_5137 (I90934,I3570);
DFFARX1 I_5138 (I654954,I3563,I90934,I90960,);
not I_5139 (I90968,I90960);
nand I_5140 (I90985,I654966,I654951);
and I_5141 (I91002,I90985,I654945);
DFFARX1 I_5142 (I91002,I3563,I90934,I91028,);
DFFARX1 I_5143 (I654960,I3563,I90934,I91045,);
and I_5144 (I91053,I91045,I654948);
nor I_5145 (I91070,I91028,I91053);
DFFARX1 I_5146 (I91070,I3563,I90934,I90902,);
nand I_5147 (I91101,I91045,I654948);
nand I_5148 (I91118,I90968,I91101);
not I_5149 (I90914,I91118);
DFFARX1 I_5150 (I654957,I3563,I90934,I91158,);
DFFARX1 I_5151 (I91158,I3563,I90934,I90923,);
nand I_5152 (I91180,I654963,I654969);
and I_5153 (I91197,I91180,I654945);
DFFARX1 I_5154 (I91197,I3563,I90934,I91223,);
DFFARX1 I_5155 (I91223,I3563,I90934,I91240,);
not I_5156 (I90926,I91240);
not I_5157 (I91262,I91223);
nand I_5158 (I90911,I91262,I91101);
nor I_5159 (I91293,I654948,I654969);
not I_5160 (I91310,I91293);
nor I_5161 (I91327,I91262,I91310);
nor I_5162 (I91344,I90968,I91327);
DFFARX1 I_5163 (I91344,I3563,I90934,I90920,);
nor I_5164 (I91375,I91028,I91310);
nor I_5165 (I90908,I91223,I91375);
nor I_5166 (I90917,I91158,I91293);
nor I_5167 (I90905,I91028,I91293);
not I_5168 (I91461,I3570);
DFFARX1 I_5169 (I1271983,I3563,I91461,I91487,);
not I_5170 (I91495,I91487);
nand I_5171 (I91512,I1271977,I1271998);
and I_5172 (I91529,I91512,I1271989);
DFFARX1 I_5173 (I91529,I3563,I91461,I91555,);
DFFARX1 I_5174 (I1271980,I3563,I91461,I91572,);
and I_5175 (I91580,I91572,I1271992);
nor I_5176 (I91597,I91555,I91580);
DFFARX1 I_5177 (I91597,I3563,I91461,I91429,);
nand I_5178 (I91628,I91572,I1271992);
nand I_5179 (I91645,I91495,I91628);
not I_5180 (I91441,I91645);
DFFARX1 I_5181 (I1271980,I3563,I91461,I91685,);
DFFARX1 I_5182 (I91685,I3563,I91461,I91450,);
nand I_5183 (I91707,I1272001,I1271986);
and I_5184 (I91724,I91707,I1271977);
DFFARX1 I_5185 (I91724,I3563,I91461,I91750,);
DFFARX1 I_5186 (I91750,I3563,I91461,I91767,);
not I_5187 (I91453,I91767);
not I_5188 (I91789,I91750);
nand I_5189 (I91438,I91789,I91628);
nor I_5190 (I91820,I1271995,I1271986);
not I_5191 (I91837,I91820);
nor I_5192 (I91854,I91789,I91837);
nor I_5193 (I91871,I91495,I91854);
DFFARX1 I_5194 (I91871,I3563,I91461,I91447,);
nor I_5195 (I91902,I91555,I91837);
nor I_5196 (I91435,I91750,I91902);
nor I_5197 (I91444,I91685,I91820);
nor I_5198 (I91432,I91555,I91820);
not I_5199 (I91988,I3570);
DFFARX1 I_5200 (I25051,I3563,I91988,I92014,);
not I_5201 (I92022,I92014);
nand I_5202 (I92039,I25039,I25045);
and I_5203 (I92056,I92039,I25048);
DFFARX1 I_5204 (I92056,I3563,I91988,I92082,);
DFFARX1 I_5205 (I25030,I3563,I91988,I92099,);
and I_5206 (I92107,I92099,I25036);
nor I_5207 (I92124,I92082,I92107);
DFFARX1 I_5208 (I92124,I3563,I91988,I91956,);
nand I_5209 (I92155,I92099,I25036);
nand I_5210 (I92172,I92022,I92155);
not I_5211 (I91968,I92172);
DFFARX1 I_5212 (I25030,I3563,I91988,I92212,);
DFFARX1 I_5213 (I92212,I3563,I91988,I91977,);
nand I_5214 (I92234,I25033,I25027);
and I_5215 (I92251,I92234,I25042);
DFFARX1 I_5216 (I92251,I3563,I91988,I92277,);
DFFARX1 I_5217 (I92277,I3563,I91988,I92294,);
not I_5218 (I91980,I92294);
not I_5219 (I92316,I92277);
nand I_5220 (I91965,I92316,I92155);
nor I_5221 (I92347,I25027,I25027);
not I_5222 (I92364,I92347);
nor I_5223 (I92381,I92316,I92364);
nor I_5224 (I92398,I92022,I92381);
DFFARX1 I_5225 (I92398,I3563,I91988,I91974,);
nor I_5226 (I92429,I92082,I92364);
nor I_5227 (I91962,I92277,I92429);
nor I_5228 (I91971,I92212,I92347);
nor I_5229 (I91959,I92082,I92347);
not I_5230 (I92515,I3570);
DFFARX1 I_5231 (I508372,I3563,I92515,I92541,);
not I_5232 (I92549,I92541);
nand I_5233 (I92566,I508366,I508357);
and I_5234 (I92583,I92566,I508378);
DFFARX1 I_5235 (I92583,I3563,I92515,I92609,);
DFFARX1 I_5236 (I508360,I3563,I92515,I92626,);
and I_5237 (I92634,I92626,I508354);
nor I_5238 (I92651,I92609,I92634);
DFFARX1 I_5239 (I92651,I3563,I92515,I92483,);
nand I_5240 (I92682,I92626,I508354);
nand I_5241 (I92699,I92549,I92682);
not I_5242 (I92495,I92699);
DFFARX1 I_5243 (I508354,I3563,I92515,I92739,);
DFFARX1 I_5244 (I92739,I3563,I92515,I92504,);
nand I_5245 (I92761,I508381,I508363);
and I_5246 (I92778,I92761,I508369);
DFFARX1 I_5247 (I92778,I3563,I92515,I92804,);
DFFARX1 I_5248 (I92804,I3563,I92515,I92821,);
not I_5249 (I92507,I92821);
not I_5250 (I92843,I92804);
nand I_5251 (I92492,I92843,I92682);
nor I_5252 (I92874,I508375,I508363);
not I_5253 (I92891,I92874);
nor I_5254 (I92908,I92843,I92891);
nor I_5255 (I92925,I92549,I92908);
DFFARX1 I_5256 (I92925,I3563,I92515,I92501,);
nor I_5257 (I92956,I92609,I92891);
nor I_5258 (I92489,I92804,I92956);
nor I_5259 (I92498,I92739,I92874);
nor I_5260 (I92486,I92609,I92874);
not I_5261 (I93042,I3570);
DFFARX1 I_5262 (I219655,I3563,I93042,I93068,);
not I_5263 (I93076,I93068);
nand I_5264 (I93093,I219649,I219643);
and I_5265 (I93110,I93093,I219664);
DFFARX1 I_5266 (I93110,I3563,I93042,I93136,);
DFFARX1 I_5267 (I219661,I3563,I93042,I93153,);
and I_5268 (I93161,I93153,I219658);
nor I_5269 (I93178,I93136,I93161);
DFFARX1 I_5270 (I93178,I3563,I93042,I93010,);
nand I_5271 (I93209,I93153,I219658);
nand I_5272 (I93226,I93076,I93209);
not I_5273 (I93022,I93226);
DFFARX1 I_5274 (I219643,I3563,I93042,I93266,);
DFFARX1 I_5275 (I93266,I3563,I93042,I93031,);
nand I_5276 (I93288,I219646,I219646);
and I_5277 (I93305,I93288,I219667);
DFFARX1 I_5278 (I93305,I3563,I93042,I93331,);
DFFARX1 I_5279 (I93331,I3563,I93042,I93348,);
not I_5280 (I93034,I93348);
not I_5281 (I93370,I93331);
nand I_5282 (I93019,I93370,I93209);
nor I_5283 (I93401,I219652,I219646);
not I_5284 (I93418,I93401);
nor I_5285 (I93435,I93370,I93418);
nor I_5286 (I93452,I93076,I93435);
DFFARX1 I_5287 (I93452,I3563,I93042,I93028,);
nor I_5288 (I93483,I93136,I93418);
nor I_5289 (I93016,I93331,I93483);
nor I_5290 (I93025,I93266,I93401);
nor I_5291 (I93013,I93136,I93401);
not I_5292 (I93569,I3570);
DFFARX1 I_5293 (I1223363,I3563,I93569,I93595,);
not I_5294 (I93603,I93595);
nand I_5295 (I93620,I1223378,I1223357);
and I_5296 (I93637,I93620,I1223360);
DFFARX1 I_5297 (I93637,I3563,I93569,I93663,);
DFFARX1 I_5298 (I1223381,I3563,I93569,I93680,);
and I_5299 (I93688,I93680,I1223360);
nor I_5300 (I93705,I93663,I93688);
DFFARX1 I_5301 (I93705,I3563,I93569,I93537,);
nand I_5302 (I93736,I93680,I1223360);
nand I_5303 (I93753,I93603,I93736);
not I_5304 (I93549,I93753);
DFFARX1 I_5305 (I1223357,I3563,I93569,I93793,);
DFFARX1 I_5306 (I93793,I3563,I93569,I93558,);
nand I_5307 (I93815,I1223369,I1223366);
and I_5308 (I93832,I93815,I1223372);
DFFARX1 I_5309 (I93832,I3563,I93569,I93858,);
DFFARX1 I_5310 (I93858,I3563,I93569,I93875,);
not I_5311 (I93561,I93875);
not I_5312 (I93897,I93858);
nand I_5313 (I93546,I93897,I93736);
nor I_5314 (I93928,I1223375,I1223366);
not I_5315 (I93945,I93928);
nor I_5316 (I93962,I93897,I93945);
nor I_5317 (I93979,I93603,I93962);
DFFARX1 I_5318 (I93979,I3563,I93569,I93555,);
nor I_5319 (I94010,I93663,I93945);
nor I_5320 (I93543,I93858,I94010);
nor I_5321 (I93552,I93793,I93928);
nor I_5322 (I93540,I93663,I93928);
not I_5323 (I94096,I3570);
DFFARX1 I_5324 (I1007908,I3563,I94096,I94122,);
not I_5325 (I94130,I94122);
nand I_5326 (I94147,I1007926,I1007920);
and I_5327 (I94164,I94147,I1007899);
DFFARX1 I_5328 (I94164,I3563,I94096,I94190,);
DFFARX1 I_5329 (I1007917,I3563,I94096,I94207,);
and I_5330 (I94215,I94207,I1007902);
nor I_5331 (I94232,I94190,I94215);
DFFARX1 I_5332 (I94232,I3563,I94096,I94064,);
nand I_5333 (I94263,I94207,I1007902);
nand I_5334 (I94280,I94130,I94263);
not I_5335 (I94076,I94280);
DFFARX1 I_5336 (I1007914,I3563,I94096,I94320,);
DFFARX1 I_5337 (I94320,I3563,I94096,I94085,);
nand I_5338 (I94342,I1007923,I1007911);
and I_5339 (I94359,I94342,I1007905);
DFFARX1 I_5340 (I94359,I3563,I94096,I94385,);
DFFARX1 I_5341 (I94385,I3563,I94096,I94402,);
not I_5342 (I94088,I94402);
not I_5343 (I94424,I94385);
nand I_5344 (I94073,I94424,I94263);
nor I_5345 (I94455,I1007899,I1007911);
not I_5346 (I94472,I94455);
nor I_5347 (I94489,I94424,I94472);
nor I_5348 (I94506,I94130,I94489);
DFFARX1 I_5349 (I94506,I3563,I94096,I94082,);
nor I_5350 (I94537,I94190,I94472);
nor I_5351 (I94070,I94385,I94537);
nor I_5352 (I94079,I94320,I94455);
nor I_5353 (I94067,I94190,I94455);
not I_5354 (I94623,I3570);
DFFARX1 I_5355 (I1273615,I3563,I94623,I94649,);
not I_5356 (I94657,I94649);
nand I_5357 (I94674,I1273609,I1273630);
and I_5358 (I94691,I94674,I1273621);
DFFARX1 I_5359 (I94691,I3563,I94623,I94717,);
DFFARX1 I_5360 (I1273612,I3563,I94623,I94734,);
and I_5361 (I94742,I94734,I1273624);
nor I_5362 (I94759,I94717,I94742);
DFFARX1 I_5363 (I94759,I3563,I94623,I94591,);
nand I_5364 (I94790,I94734,I1273624);
nand I_5365 (I94807,I94657,I94790);
not I_5366 (I94603,I94807);
DFFARX1 I_5367 (I1273612,I3563,I94623,I94847,);
DFFARX1 I_5368 (I94847,I3563,I94623,I94612,);
nand I_5369 (I94869,I1273633,I1273618);
and I_5370 (I94886,I94869,I1273609);
DFFARX1 I_5371 (I94886,I3563,I94623,I94912,);
DFFARX1 I_5372 (I94912,I3563,I94623,I94929,);
not I_5373 (I94615,I94929);
not I_5374 (I94951,I94912);
nand I_5375 (I94600,I94951,I94790);
nor I_5376 (I94982,I1273627,I1273618);
not I_5377 (I94999,I94982);
nor I_5378 (I95016,I94951,I94999);
nor I_5379 (I95033,I94657,I95016);
DFFARX1 I_5380 (I95033,I3563,I94623,I94609,);
nor I_5381 (I95064,I94717,I94999);
nor I_5382 (I94597,I94912,I95064);
nor I_5383 (I94606,I94847,I94982);
nor I_5384 (I94594,I94717,I94982);
not I_5385 (I95150,I3570);
DFFARX1 I_5386 (I1125681,I3563,I95150,I95176,);
not I_5387 (I95184,I95176);
nand I_5388 (I95201,I1125696,I1125675);
and I_5389 (I95218,I95201,I1125678);
DFFARX1 I_5390 (I95218,I3563,I95150,I95244,);
DFFARX1 I_5391 (I1125699,I3563,I95150,I95261,);
and I_5392 (I95269,I95261,I1125678);
nor I_5393 (I95286,I95244,I95269);
DFFARX1 I_5394 (I95286,I3563,I95150,I95118,);
nand I_5395 (I95317,I95261,I1125678);
nand I_5396 (I95334,I95184,I95317);
not I_5397 (I95130,I95334);
DFFARX1 I_5398 (I1125675,I3563,I95150,I95374,);
DFFARX1 I_5399 (I95374,I3563,I95150,I95139,);
nand I_5400 (I95396,I1125687,I1125684);
and I_5401 (I95413,I95396,I1125690);
DFFARX1 I_5402 (I95413,I3563,I95150,I95439,);
DFFARX1 I_5403 (I95439,I3563,I95150,I95456,);
not I_5404 (I95142,I95456);
not I_5405 (I95478,I95439);
nand I_5406 (I95127,I95478,I95317);
nor I_5407 (I95509,I1125693,I1125684);
not I_5408 (I95526,I95509);
nor I_5409 (I95543,I95478,I95526);
nor I_5410 (I95560,I95184,I95543);
DFFARX1 I_5411 (I95560,I3563,I95150,I95136,);
nor I_5412 (I95591,I95244,I95526);
nor I_5413 (I95124,I95439,I95591);
nor I_5414 (I95133,I95374,I95509);
nor I_5415 (I95121,I95244,I95509);
not I_5416 (I95677,I3570);
DFFARX1 I_5417 (I166700,I3563,I95677,I95703,);
not I_5418 (I95711,I95703);
nand I_5419 (I95728,I166694,I166688);
and I_5420 (I95745,I95728,I166709);
DFFARX1 I_5421 (I95745,I3563,I95677,I95771,);
DFFARX1 I_5422 (I166706,I3563,I95677,I95788,);
and I_5423 (I95796,I95788,I166703);
nor I_5424 (I95813,I95771,I95796);
DFFARX1 I_5425 (I95813,I3563,I95677,I95645,);
nand I_5426 (I95844,I95788,I166703);
nand I_5427 (I95861,I95711,I95844);
not I_5428 (I95657,I95861);
DFFARX1 I_5429 (I166688,I3563,I95677,I95901,);
DFFARX1 I_5430 (I95901,I3563,I95677,I95666,);
nand I_5431 (I95923,I166691,I166691);
and I_5432 (I95940,I95923,I166712);
DFFARX1 I_5433 (I95940,I3563,I95677,I95966,);
DFFARX1 I_5434 (I95966,I3563,I95677,I95983,);
not I_5435 (I95669,I95983);
not I_5436 (I96005,I95966);
nand I_5437 (I95654,I96005,I95844);
nor I_5438 (I96036,I166697,I166691);
not I_5439 (I96053,I96036);
nor I_5440 (I96070,I96005,I96053);
nor I_5441 (I96087,I95711,I96070);
DFFARX1 I_5442 (I96087,I3563,I95677,I95663,);
nor I_5443 (I96118,I95771,I96053);
nor I_5444 (I95651,I95966,I96118);
nor I_5445 (I95660,I95901,I96036);
nor I_5446 (I95648,I95771,I96036);
not I_5447 (I96204,I3570);
DFFARX1 I_5448 (I807549,I3563,I96204,I96230,);
not I_5449 (I96238,I96230);
nand I_5450 (I96255,I807540,I807558);
and I_5451 (I96272,I96255,I807537);
DFFARX1 I_5452 (I96272,I3563,I96204,I96298,);
DFFARX1 I_5453 (I807540,I3563,I96204,I96315,);
and I_5454 (I96323,I96315,I807543);
nor I_5455 (I96340,I96298,I96323);
DFFARX1 I_5456 (I96340,I3563,I96204,I96172,);
nand I_5457 (I96371,I96315,I807543);
nand I_5458 (I96388,I96238,I96371);
not I_5459 (I96184,I96388);
DFFARX1 I_5460 (I807537,I3563,I96204,I96428,);
DFFARX1 I_5461 (I96428,I3563,I96204,I96193,);
nand I_5462 (I96450,I807555,I807546);
and I_5463 (I96467,I96450,I807561);
DFFARX1 I_5464 (I96467,I3563,I96204,I96493,);
DFFARX1 I_5465 (I96493,I3563,I96204,I96510,);
not I_5466 (I96196,I96510);
not I_5467 (I96532,I96493);
nand I_5468 (I96181,I96532,I96371);
nor I_5469 (I96563,I807552,I807546);
not I_5470 (I96580,I96563);
nor I_5471 (I96597,I96532,I96580);
nor I_5472 (I96614,I96238,I96597);
DFFARX1 I_5473 (I96614,I3563,I96204,I96190,);
nor I_5474 (I96645,I96298,I96580);
nor I_5475 (I96178,I96493,I96645);
nor I_5476 (I96187,I96428,I96563);
nor I_5477 (I96175,I96298,I96563);
not I_5478 (I96731,I3570);
DFFARX1 I_5479 (I601200,I3563,I96731,I96757,);
not I_5480 (I96765,I96757);
nand I_5481 (I96782,I601212,I601197);
and I_5482 (I96799,I96782,I601191);
DFFARX1 I_5483 (I96799,I3563,I96731,I96825,);
DFFARX1 I_5484 (I601206,I3563,I96731,I96842,);
and I_5485 (I96850,I96842,I601194);
nor I_5486 (I96867,I96825,I96850);
DFFARX1 I_5487 (I96867,I3563,I96731,I96699,);
nand I_5488 (I96898,I96842,I601194);
nand I_5489 (I96915,I96765,I96898);
not I_5490 (I96711,I96915);
DFFARX1 I_5491 (I601203,I3563,I96731,I96955,);
DFFARX1 I_5492 (I96955,I3563,I96731,I96720,);
nand I_5493 (I96977,I601209,I601215);
and I_5494 (I96994,I96977,I601191);
DFFARX1 I_5495 (I96994,I3563,I96731,I97020,);
DFFARX1 I_5496 (I97020,I3563,I96731,I97037,);
not I_5497 (I96723,I97037);
not I_5498 (I97059,I97020);
nand I_5499 (I96708,I97059,I96898);
nor I_5500 (I97090,I601194,I601215);
not I_5501 (I97107,I97090);
nor I_5502 (I97124,I97059,I97107);
nor I_5503 (I97141,I96765,I97124);
DFFARX1 I_5504 (I97141,I3563,I96731,I96717,);
nor I_5505 (I97172,I96825,I97107);
nor I_5506 (I96705,I97020,I97172);
nor I_5507 (I96714,I96955,I97090);
nor I_5508 (I96702,I96825,I97090);
not I_5509 (I97258,I3570);
DFFARX1 I_5510 (I175030,I3563,I97258,I97284,);
not I_5511 (I97292,I97284);
nand I_5512 (I97309,I175024,I175018);
and I_5513 (I97326,I97309,I175039);
DFFARX1 I_5514 (I97326,I3563,I97258,I97352,);
DFFARX1 I_5515 (I175036,I3563,I97258,I97369,);
and I_5516 (I97377,I97369,I175033);
nor I_5517 (I97394,I97352,I97377);
DFFARX1 I_5518 (I97394,I3563,I97258,I97226,);
nand I_5519 (I97425,I97369,I175033);
nand I_5520 (I97442,I97292,I97425);
not I_5521 (I97238,I97442);
DFFARX1 I_5522 (I175018,I3563,I97258,I97482,);
DFFARX1 I_5523 (I97482,I3563,I97258,I97247,);
nand I_5524 (I97504,I175021,I175021);
and I_5525 (I97521,I97504,I175042);
DFFARX1 I_5526 (I97521,I3563,I97258,I97547,);
DFFARX1 I_5527 (I97547,I3563,I97258,I97564,);
not I_5528 (I97250,I97564);
not I_5529 (I97586,I97547);
nand I_5530 (I97235,I97586,I97425);
nor I_5531 (I97617,I175027,I175021);
not I_5532 (I97634,I97617);
nor I_5533 (I97651,I97586,I97634);
nor I_5534 (I97668,I97292,I97651);
DFFARX1 I_5535 (I97668,I3563,I97258,I97244,);
nor I_5536 (I97699,I97352,I97634);
nor I_5537 (I97232,I97547,I97699);
nor I_5538 (I97241,I97482,I97617);
nor I_5539 (I97229,I97352,I97617);
not I_5540 (I97785,I3570);
DFFARX1 I_5541 (I49293,I3563,I97785,I97811,);
not I_5542 (I97819,I97811);
nand I_5543 (I97836,I49281,I49287);
and I_5544 (I97853,I97836,I49290);
DFFARX1 I_5545 (I97853,I3563,I97785,I97879,);
DFFARX1 I_5546 (I49272,I3563,I97785,I97896,);
and I_5547 (I97904,I97896,I49278);
nor I_5548 (I97921,I97879,I97904);
DFFARX1 I_5549 (I97921,I3563,I97785,I97753,);
nand I_5550 (I97952,I97896,I49278);
nand I_5551 (I97969,I97819,I97952);
not I_5552 (I97765,I97969);
DFFARX1 I_5553 (I49272,I3563,I97785,I98009,);
DFFARX1 I_5554 (I98009,I3563,I97785,I97774,);
nand I_5555 (I98031,I49275,I49269);
and I_5556 (I98048,I98031,I49284);
DFFARX1 I_5557 (I98048,I3563,I97785,I98074,);
DFFARX1 I_5558 (I98074,I3563,I97785,I98091,);
not I_5559 (I97777,I98091);
not I_5560 (I98113,I98074);
nand I_5561 (I97762,I98113,I97952);
nor I_5562 (I98144,I49269,I49269);
not I_5563 (I98161,I98144);
nor I_5564 (I98178,I98113,I98161);
nor I_5565 (I98195,I97819,I98178);
DFFARX1 I_5566 (I98195,I3563,I97785,I97771,);
nor I_5567 (I98226,I97879,I98161);
nor I_5568 (I97759,I98074,I98226);
nor I_5569 (I97768,I98009,I98144);
nor I_5570 (I97756,I97879,I98144);
not I_5571 (I98312,I3570);
DFFARX1 I_5572 (I832145,I3563,I98312,I98338,);
not I_5573 (I98346,I98338);
nand I_5574 (I98363,I832142,I832157);
and I_5575 (I98380,I98363,I832139);
DFFARX1 I_5576 (I98380,I3563,I98312,I98406,);
DFFARX1 I_5577 (I832136,I3563,I98312,I98423,);
and I_5578 (I98431,I98423,I832136);
nor I_5579 (I98448,I98406,I98431);
DFFARX1 I_5580 (I98448,I3563,I98312,I98280,);
nand I_5581 (I98479,I98423,I832136);
nand I_5582 (I98496,I98346,I98479);
not I_5583 (I98292,I98496);
DFFARX1 I_5584 (I832139,I3563,I98312,I98536,);
DFFARX1 I_5585 (I98536,I3563,I98312,I98301,);
nand I_5586 (I98558,I832151,I832142);
and I_5587 (I98575,I98558,I832154);
DFFARX1 I_5588 (I98575,I3563,I98312,I98601,);
DFFARX1 I_5589 (I98601,I3563,I98312,I98618,);
not I_5590 (I98304,I98618);
not I_5591 (I98640,I98601);
nand I_5592 (I98289,I98640,I98479);
nor I_5593 (I98671,I832148,I832142);
not I_5594 (I98688,I98671);
nor I_5595 (I98705,I98640,I98688);
nor I_5596 (I98722,I98346,I98705);
DFFARX1 I_5597 (I98722,I3563,I98312,I98298,);
nor I_5598 (I98753,I98406,I98688);
nor I_5599 (I98286,I98601,I98753);
nor I_5600 (I98295,I98536,I98671);
nor I_5601 (I98283,I98406,I98671);
not I_5602 (I98839,I3570);
DFFARX1 I_5603 (I285105,I3563,I98839,I98865,);
not I_5604 (I98873,I98865);
nand I_5605 (I98890,I285099,I285093);
and I_5606 (I98907,I98890,I285114);
DFFARX1 I_5607 (I98907,I3563,I98839,I98933,);
DFFARX1 I_5608 (I285111,I3563,I98839,I98950,);
and I_5609 (I98958,I98950,I285108);
nor I_5610 (I98975,I98933,I98958);
DFFARX1 I_5611 (I98975,I3563,I98839,I98807,);
nand I_5612 (I99006,I98950,I285108);
nand I_5613 (I99023,I98873,I99006);
not I_5614 (I98819,I99023);
DFFARX1 I_5615 (I285093,I3563,I98839,I99063,);
DFFARX1 I_5616 (I99063,I3563,I98839,I98828,);
nand I_5617 (I99085,I285096,I285096);
and I_5618 (I99102,I99085,I285117);
DFFARX1 I_5619 (I99102,I3563,I98839,I99128,);
DFFARX1 I_5620 (I99128,I3563,I98839,I99145,);
not I_5621 (I98831,I99145);
not I_5622 (I99167,I99128);
nand I_5623 (I98816,I99167,I99006);
nor I_5624 (I99198,I285102,I285096);
not I_5625 (I99215,I99198);
nor I_5626 (I99232,I99167,I99215);
nor I_5627 (I99249,I98873,I99232);
DFFARX1 I_5628 (I99249,I3563,I98839,I98825,);
nor I_5629 (I99280,I98933,I99215);
nor I_5630 (I98813,I99128,I99280);
nor I_5631 (I98822,I99063,I99198);
nor I_5632 (I98810,I98933,I99198);
not I_5633 (I99366,I3570);
DFFARX1 I_5634 (I1345820,I3563,I99366,I99392,);
not I_5635 (I99400,I99392);
nand I_5636 (I99417,I1345814,I1345835);
and I_5637 (I99434,I99417,I1345811);
DFFARX1 I_5638 (I99434,I3563,I99366,I99460,);
DFFARX1 I_5639 (I1345832,I3563,I99366,I99477,);
and I_5640 (I99485,I99477,I1345829);
nor I_5641 (I99502,I99460,I99485);
DFFARX1 I_5642 (I99502,I3563,I99366,I99334,);
nand I_5643 (I99533,I99477,I1345829);
nand I_5644 (I99550,I99400,I99533);
not I_5645 (I99346,I99550);
DFFARX1 I_5646 (I1345817,I3563,I99366,I99590,);
DFFARX1 I_5647 (I99590,I3563,I99366,I99355,);
nand I_5648 (I99612,I1345826,I1345823);
and I_5649 (I99629,I99612,I1345808);
DFFARX1 I_5650 (I99629,I3563,I99366,I99655,);
DFFARX1 I_5651 (I99655,I3563,I99366,I99672,);
not I_5652 (I99358,I99672);
not I_5653 (I99694,I99655);
nand I_5654 (I99343,I99694,I99533);
nor I_5655 (I99725,I1345808,I1345823);
not I_5656 (I99742,I99725);
nor I_5657 (I99759,I99694,I99742);
nor I_5658 (I99776,I99400,I99759);
DFFARX1 I_5659 (I99776,I3563,I99366,I99352,);
nor I_5660 (I99807,I99460,I99742);
nor I_5661 (I99340,I99655,I99807);
nor I_5662 (I99349,I99590,I99725);
nor I_5663 (I99337,I99460,I99725);
not I_5664 (I99893,I3570);
DFFARX1 I_5665 (I299621,I3563,I99893,I99919,);
not I_5666 (I99927,I99919);
nand I_5667 (I99944,I299603,I299618);
and I_5668 (I99961,I99944,I299594);
DFFARX1 I_5669 (I99961,I3563,I99893,I99987,);
DFFARX1 I_5670 (I299597,I3563,I99893,I100004,);
and I_5671 (I100012,I100004,I299612);
nor I_5672 (I100029,I99987,I100012);
DFFARX1 I_5673 (I100029,I3563,I99893,I99861,);
nand I_5674 (I100060,I100004,I299612);
nand I_5675 (I100077,I99927,I100060);
not I_5676 (I99873,I100077);
DFFARX1 I_5677 (I299615,I3563,I99893,I100117,);
DFFARX1 I_5678 (I100117,I3563,I99893,I99882,);
nand I_5679 (I100139,I299594,I299606);
and I_5680 (I100156,I100139,I299600);
DFFARX1 I_5681 (I100156,I3563,I99893,I100182,);
DFFARX1 I_5682 (I100182,I3563,I99893,I100199,);
not I_5683 (I99885,I100199);
not I_5684 (I100221,I100182);
nand I_5685 (I99870,I100221,I100060);
nor I_5686 (I100252,I299609,I299606);
not I_5687 (I100269,I100252);
nor I_5688 (I100286,I100221,I100269);
nor I_5689 (I100303,I99927,I100286);
DFFARX1 I_5690 (I100303,I3563,I99893,I99879,);
nor I_5691 (I100334,I99987,I100269);
nor I_5692 (I99867,I100182,I100334);
nor I_5693 (I99876,I100117,I100252);
nor I_5694 (I99864,I99987,I100252);
not I_5695 (I100420,I3570);
DFFARX1 I_5696 (I1401155,I3563,I100420,I100446,);
not I_5697 (I100454,I100446);
nand I_5698 (I100471,I1401149,I1401170);
and I_5699 (I100488,I100471,I1401146);
DFFARX1 I_5700 (I100488,I3563,I100420,I100514,);
DFFARX1 I_5701 (I1401167,I3563,I100420,I100531,);
and I_5702 (I100539,I100531,I1401164);
nor I_5703 (I100556,I100514,I100539);
DFFARX1 I_5704 (I100556,I3563,I100420,I100388,);
nand I_5705 (I100587,I100531,I1401164);
nand I_5706 (I100604,I100454,I100587);
not I_5707 (I100400,I100604);
DFFARX1 I_5708 (I1401152,I3563,I100420,I100644,);
DFFARX1 I_5709 (I100644,I3563,I100420,I100409,);
nand I_5710 (I100666,I1401161,I1401158);
and I_5711 (I100683,I100666,I1401143);
DFFARX1 I_5712 (I100683,I3563,I100420,I100709,);
DFFARX1 I_5713 (I100709,I3563,I100420,I100726,);
not I_5714 (I100412,I100726);
not I_5715 (I100748,I100709);
nand I_5716 (I100397,I100748,I100587);
nor I_5717 (I100779,I1401143,I1401158);
not I_5718 (I100796,I100779);
nor I_5719 (I100813,I100748,I100796);
nor I_5720 (I100830,I100454,I100813);
DFFARX1 I_5721 (I100830,I3563,I100420,I100406,);
nor I_5722 (I100861,I100514,I100796);
nor I_5723 (I100394,I100709,I100861);
nor I_5724 (I100403,I100644,I100779);
nor I_5725 (I100391,I100514,I100779);
not I_5726 (I100947,I3570);
DFFARX1 I_5727 (I692527,I3563,I100947,I100973,);
not I_5728 (I100981,I100973);
nand I_5729 (I100998,I692518,I692536);
and I_5730 (I101015,I100998,I692515);
DFFARX1 I_5731 (I101015,I3563,I100947,I101041,);
DFFARX1 I_5732 (I692518,I3563,I100947,I101058,);
and I_5733 (I101066,I101058,I692521);
nor I_5734 (I101083,I101041,I101066);
DFFARX1 I_5735 (I101083,I3563,I100947,I100915,);
nand I_5736 (I101114,I101058,I692521);
nand I_5737 (I101131,I100981,I101114);
not I_5738 (I100927,I101131);
DFFARX1 I_5739 (I692515,I3563,I100947,I101171,);
DFFARX1 I_5740 (I101171,I3563,I100947,I100936,);
nand I_5741 (I101193,I692533,I692524);
and I_5742 (I101210,I101193,I692539);
DFFARX1 I_5743 (I101210,I3563,I100947,I101236,);
DFFARX1 I_5744 (I101236,I3563,I100947,I101253,);
not I_5745 (I100939,I101253);
not I_5746 (I101275,I101236);
nand I_5747 (I100924,I101275,I101114);
nor I_5748 (I101306,I692530,I692524);
not I_5749 (I101323,I101306);
nor I_5750 (I101340,I101275,I101323);
nor I_5751 (I101357,I100981,I101340);
DFFARX1 I_5752 (I101357,I3563,I100947,I100933,);
nor I_5753 (I101388,I101041,I101323);
nor I_5754 (I100921,I101236,I101388);
nor I_5755 (I100930,I101171,I101306);
nor I_5756 (I100918,I101041,I101306);
not I_5757 (I101474,I3570);
DFFARX1 I_5758 (I826875,I3563,I101474,I101500,);
not I_5759 (I101508,I101500);
nand I_5760 (I101525,I826872,I826887);
and I_5761 (I101542,I101525,I826869);
DFFARX1 I_5762 (I101542,I3563,I101474,I101568,);
DFFARX1 I_5763 (I826866,I3563,I101474,I101585,);
and I_5764 (I101593,I101585,I826866);
nor I_5765 (I101610,I101568,I101593);
DFFARX1 I_5766 (I101610,I3563,I101474,I101442,);
nand I_5767 (I101641,I101585,I826866);
nand I_5768 (I101658,I101508,I101641);
not I_5769 (I101454,I101658);
DFFARX1 I_5770 (I826869,I3563,I101474,I101698,);
DFFARX1 I_5771 (I101698,I3563,I101474,I101463,);
nand I_5772 (I101720,I826881,I826872);
and I_5773 (I101737,I101720,I826884);
DFFARX1 I_5774 (I101737,I3563,I101474,I101763,);
DFFARX1 I_5775 (I101763,I3563,I101474,I101780,);
not I_5776 (I101466,I101780);
not I_5777 (I101802,I101763);
nand I_5778 (I101451,I101802,I101641);
nor I_5779 (I101833,I826878,I826872);
not I_5780 (I101850,I101833);
nor I_5781 (I101867,I101802,I101850);
nor I_5782 (I101884,I101508,I101867);
DFFARX1 I_5783 (I101884,I3563,I101474,I101460,);
nor I_5784 (I101915,I101568,I101850);
nor I_5785 (I101448,I101763,I101915);
nor I_5786 (I101457,I101698,I101833);
nor I_5787 (I101445,I101568,I101833);
not I_5788 (I102001,I3570);
DFFARX1 I_5789 (I28213,I3563,I102001,I102027,);
not I_5790 (I102035,I102027);
nand I_5791 (I102052,I28201,I28207);
and I_5792 (I102069,I102052,I28210);
DFFARX1 I_5793 (I102069,I3563,I102001,I102095,);
DFFARX1 I_5794 (I28192,I3563,I102001,I102112,);
and I_5795 (I102120,I102112,I28198);
nor I_5796 (I102137,I102095,I102120);
DFFARX1 I_5797 (I102137,I3563,I102001,I101969,);
nand I_5798 (I102168,I102112,I28198);
nand I_5799 (I102185,I102035,I102168);
not I_5800 (I101981,I102185);
DFFARX1 I_5801 (I28192,I3563,I102001,I102225,);
DFFARX1 I_5802 (I102225,I3563,I102001,I101990,);
nand I_5803 (I102247,I28195,I28189);
and I_5804 (I102264,I102247,I28204);
DFFARX1 I_5805 (I102264,I3563,I102001,I102290,);
DFFARX1 I_5806 (I102290,I3563,I102001,I102307,);
not I_5807 (I101993,I102307);
not I_5808 (I102329,I102290);
nand I_5809 (I101978,I102329,I102168);
nor I_5810 (I102360,I28189,I28189);
not I_5811 (I102377,I102360);
nor I_5812 (I102394,I102329,I102377);
nor I_5813 (I102411,I102035,I102394);
DFFARX1 I_5814 (I102411,I3563,I102001,I101987,);
nor I_5815 (I102442,I102095,I102377);
nor I_5816 (I101975,I102290,I102442);
nor I_5817 (I101984,I102225,I102360);
nor I_5818 (I101972,I102095,I102360);
not I_5819 (I102528,I3570);
DFFARX1 I_5820 (I484980,I3563,I102528,I102554,);
not I_5821 (I102562,I102554);
nand I_5822 (I102579,I484974,I484965);
and I_5823 (I102596,I102579,I484986);
DFFARX1 I_5824 (I102596,I3563,I102528,I102622,);
DFFARX1 I_5825 (I484968,I3563,I102528,I102639,);
and I_5826 (I102647,I102639,I484962);
nor I_5827 (I102664,I102622,I102647);
DFFARX1 I_5828 (I102664,I3563,I102528,I102496,);
nand I_5829 (I102695,I102639,I484962);
nand I_5830 (I102712,I102562,I102695);
not I_5831 (I102508,I102712);
DFFARX1 I_5832 (I484962,I3563,I102528,I102752,);
DFFARX1 I_5833 (I102752,I3563,I102528,I102517,);
nand I_5834 (I102774,I484989,I484971);
and I_5835 (I102791,I102774,I484977);
DFFARX1 I_5836 (I102791,I3563,I102528,I102817,);
DFFARX1 I_5837 (I102817,I3563,I102528,I102834,);
not I_5838 (I102520,I102834);
not I_5839 (I102856,I102817);
nand I_5840 (I102505,I102856,I102695);
nor I_5841 (I102887,I484983,I484971);
not I_5842 (I102904,I102887);
nor I_5843 (I102921,I102856,I102904);
nor I_5844 (I102938,I102562,I102921);
DFFARX1 I_5845 (I102938,I3563,I102528,I102514,);
nor I_5846 (I102969,I102622,I102904);
nor I_5847 (I102502,I102817,I102969);
nor I_5848 (I102511,I102752,I102887);
nor I_5849 (I102499,I102622,I102887);
not I_5850 (I103055,I3570);
DFFARX1 I_5851 (I1333325,I3563,I103055,I103081,);
not I_5852 (I103089,I103081);
nand I_5853 (I103106,I1333319,I1333340);
and I_5854 (I103123,I103106,I1333316);
DFFARX1 I_5855 (I103123,I3563,I103055,I103149,);
DFFARX1 I_5856 (I1333337,I3563,I103055,I103166,);
and I_5857 (I103174,I103166,I1333334);
nor I_5858 (I103191,I103149,I103174);
DFFARX1 I_5859 (I103191,I3563,I103055,I103023,);
nand I_5860 (I103222,I103166,I1333334);
nand I_5861 (I103239,I103089,I103222);
not I_5862 (I103035,I103239);
DFFARX1 I_5863 (I1333322,I3563,I103055,I103279,);
DFFARX1 I_5864 (I103279,I3563,I103055,I103044,);
nand I_5865 (I103301,I1333331,I1333328);
and I_5866 (I103318,I103301,I1333313);
DFFARX1 I_5867 (I103318,I3563,I103055,I103344,);
DFFARX1 I_5868 (I103344,I3563,I103055,I103361,);
not I_5869 (I103047,I103361);
not I_5870 (I103383,I103344);
nand I_5871 (I103032,I103383,I103222);
nor I_5872 (I103414,I1333313,I1333328);
not I_5873 (I103431,I103414);
nor I_5874 (I103448,I103383,I103431);
nor I_5875 (I103465,I103089,I103448);
DFFARX1 I_5876 (I103465,I3563,I103055,I103041,);
nor I_5877 (I103496,I103149,I103431);
nor I_5878 (I103029,I103344,I103496);
nor I_5879 (I103038,I103279,I103414);
nor I_5880 (I103026,I103149,I103414);
not I_5881 (I103582,I3570);
DFFARX1 I_5882 (I429492,I3563,I103582,I103608,);
not I_5883 (I103616,I103608);
nand I_5884 (I103633,I429486,I429477);
and I_5885 (I103650,I103633,I429498);
DFFARX1 I_5886 (I103650,I3563,I103582,I103676,);
DFFARX1 I_5887 (I429480,I3563,I103582,I103693,);
and I_5888 (I103701,I103693,I429474);
nor I_5889 (I103718,I103676,I103701);
DFFARX1 I_5890 (I103718,I3563,I103582,I103550,);
nand I_5891 (I103749,I103693,I429474);
nand I_5892 (I103766,I103616,I103749);
not I_5893 (I103562,I103766);
DFFARX1 I_5894 (I429474,I3563,I103582,I103806,);
DFFARX1 I_5895 (I103806,I3563,I103582,I103571,);
nand I_5896 (I103828,I429501,I429483);
and I_5897 (I103845,I103828,I429489);
DFFARX1 I_5898 (I103845,I3563,I103582,I103871,);
DFFARX1 I_5899 (I103871,I3563,I103582,I103888,);
not I_5900 (I103574,I103888);
not I_5901 (I103910,I103871);
nand I_5902 (I103559,I103910,I103749);
nor I_5903 (I103941,I429495,I429483);
not I_5904 (I103958,I103941);
nor I_5905 (I103975,I103910,I103958);
nor I_5906 (I103992,I103616,I103975);
DFFARX1 I_5907 (I103992,I3563,I103582,I103568,);
nor I_5908 (I104023,I103676,I103958);
nor I_5909 (I103556,I103871,I104023);
nor I_5910 (I103565,I103806,I103941);
nor I_5911 (I103553,I103676,I103941);
not I_5912 (I104109,I3570);
DFFARX1 I_5913 (I996280,I3563,I104109,I104135,);
not I_5914 (I104143,I104135);
nand I_5915 (I104160,I996298,I996292);
and I_5916 (I104177,I104160,I996271);
DFFARX1 I_5917 (I104177,I3563,I104109,I104203,);
DFFARX1 I_5918 (I996289,I3563,I104109,I104220,);
and I_5919 (I104228,I104220,I996274);
nor I_5920 (I104245,I104203,I104228);
DFFARX1 I_5921 (I104245,I3563,I104109,I104077,);
nand I_5922 (I104276,I104220,I996274);
nand I_5923 (I104293,I104143,I104276);
not I_5924 (I104089,I104293);
DFFARX1 I_5925 (I996286,I3563,I104109,I104333,);
DFFARX1 I_5926 (I104333,I3563,I104109,I104098,);
nand I_5927 (I104355,I996295,I996283);
and I_5928 (I104372,I104355,I996277);
DFFARX1 I_5929 (I104372,I3563,I104109,I104398,);
DFFARX1 I_5930 (I104398,I3563,I104109,I104415,);
not I_5931 (I104101,I104415);
not I_5932 (I104437,I104398);
nand I_5933 (I104086,I104437,I104276);
nor I_5934 (I104468,I996271,I996283);
not I_5935 (I104485,I104468);
nor I_5936 (I104502,I104437,I104485);
nor I_5937 (I104519,I104143,I104502);
DFFARX1 I_5938 (I104519,I3563,I104109,I104095,);
nor I_5939 (I104550,I104203,I104485);
nor I_5940 (I104083,I104398,I104550);
nor I_5941 (I104092,I104333,I104468);
nor I_5942 (I104080,I104203,I104468);
not I_5943 (I104636,I3570);
DFFARX1 I_5944 (I793677,I3563,I104636,I104662,);
not I_5945 (I104670,I104662);
nand I_5946 (I104687,I793668,I793686);
and I_5947 (I104704,I104687,I793665);
DFFARX1 I_5948 (I104704,I3563,I104636,I104730,);
DFFARX1 I_5949 (I793668,I3563,I104636,I104747,);
and I_5950 (I104755,I104747,I793671);
nor I_5951 (I104772,I104730,I104755);
DFFARX1 I_5952 (I104772,I3563,I104636,I104604,);
nand I_5953 (I104803,I104747,I793671);
nand I_5954 (I104820,I104670,I104803);
not I_5955 (I104616,I104820);
DFFARX1 I_5956 (I793665,I3563,I104636,I104860,);
DFFARX1 I_5957 (I104860,I3563,I104636,I104625,);
nand I_5958 (I104882,I793683,I793674);
and I_5959 (I104899,I104882,I793689);
DFFARX1 I_5960 (I104899,I3563,I104636,I104925,);
DFFARX1 I_5961 (I104925,I3563,I104636,I104942,);
not I_5962 (I104628,I104942);
not I_5963 (I104964,I104925);
nand I_5964 (I104613,I104964,I104803);
nor I_5965 (I104995,I793680,I793674);
not I_5966 (I105012,I104995);
nor I_5967 (I105029,I104964,I105012);
nor I_5968 (I105046,I104670,I105029);
DFFARX1 I_5969 (I105046,I3563,I104636,I104622,);
nor I_5970 (I105077,I104730,I105012);
nor I_5971 (I104610,I104925,I105077);
nor I_5972 (I104619,I104860,I104995);
nor I_5973 (I104607,I104730,I104995);
not I_5974 (I105163,I3570);
DFFARX1 I_5975 (I211920,I3563,I105163,I105189,);
not I_5976 (I105197,I105189);
nand I_5977 (I105214,I211914,I211908);
and I_5978 (I105231,I105214,I211929);
DFFARX1 I_5979 (I105231,I3563,I105163,I105257,);
DFFARX1 I_5980 (I211926,I3563,I105163,I105274,);
and I_5981 (I105282,I105274,I211923);
nor I_5982 (I105299,I105257,I105282);
DFFARX1 I_5983 (I105299,I3563,I105163,I105131,);
nand I_5984 (I105330,I105274,I211923);
nand I_5985 (I105347,I105197,I105330);
not I_5986 (I105143,I105347);
DFFARX1 I_5987 (I211908,I3563,I105163,I105387,);
DFFARX1 I_5988 (I105387,I3563,I105163,I105152,);
nand I_5989 (I105409,I211911,I211911);
and I_5990 (I105426,I105409,I211932);
DFFARX1 I_5991 (I105426,I3563,I105163,I105452,);
DFFARX1 I_5992 (I105452,I3563,I105163,I105469,);
not I_5993 (I105155,I105469);
not I_5994 (I105491,I105452);
nand I_5995 (I105140,I105491,I105330);
nor I_5996 (I105522,I211917,I211911);
not I_5997 (I105539,I105522);
nor I_5998 (I105556,I105491,I105539);
nor I_5999 (I105573,I105197,I105556);
DFFARX1 I_6000 (I105573,I3563,I105163,I105149,);
nor I_6001 (I105604,I105257,I105539);
nor I_6002 (I105137,I105452,I105604);
nor I_6003 (I105146,I105387,I105522);
nor I_6004 (I105134,I105257,I105522);
not I_6005 (I105690,I3570);
DFFARX1 I_6006 (I635880,I3563,I105690,I105716,);
not I_6007 (I105724,I105716);
nand I_6008 (I105741,I635892,I635877);
and I_6009 (I105758,I105741,I635871);
DFFARX1 I_6010 (I105758,I3563,I105690,I105784,);
DFFARX1 I_6011 (I635886,I3563,I105690,I105801,);
and I_6012 (I105809,I105801,I635874);
nor I_6013 (I105826,I105784,I105809);
DFFARX1 I_6014 (I105826,I3563,I105690,I105658,);
nand I_6015 (I105857,I105801,I635874);
nand I_6016 (I105874,I105724,I105857);
not I_6017 (I105670,I105874);
DFFARX1 I_6018 (I635883,I3563,I105690,I105914,);
DFFARX1 I_6019 (I105914,I3563,I105690,I105679,);
nand I_6020 (I105936,I635889,I635895);
and I_6021 (I105953,I105936,I635871);
DFFARX1 I_6022 (I105953,I3563,I105690,I105979,);
DFFARX1 I_6023 (I105979,I3563,I105690,I105996,);
not I_6024 (I105682,I105996);
not I_6025 (I106018,I105979);
nand I_6026 (I105667,I106018,I105857);
nor I_6027 (I106049,I635874,I635895);
not I_6028 (I106066,I106049);
nor I_6029 (I106083,I106018,I106066);
nor I_6030 (I106100,I105724,I106083);
DFFARX1 I_6031 (I106100,I3563,I105690,I105676,);
nor I_6032 (I106131,I105784,I106066);
nor I_6033 (I105664,I105979,I106131);
nor I_6034 (I105673,I105914,I106049);
nor I_6035 (I105661,I105784,I106049);
not I_6036 (I106217,I3570);
DFFARX1 I_6037 (I778071,I3563,I106217,I106243,);
not I_6038 (I106251,I106243);
nand I_6039 (I106268,I778062,I778080);
and I_6040 (I106285,I106268,I778059);
DFFARX1 I_6041 (I106285,I3563,I106217,I106311,);
DFFARX1 I_6042 (I778062,I3563,I106217,I106328,);
and I_6043 (I106336,I106328,I778065);
nor I_6044 (I106353,I106311,I106336);
DFFARX1 I_6045 (I106353,I3563,I106217,I106185,);
nand I_6046 (I106384,I106328,I778065);
nand I_6047 (I106401,I106251,I106384);
not I_6048 (I106197,I106401);
DFFARX1 I_6049 (I778059,I3563,I106217,I106441,);
DFFARX1 I_6050 (I106441,I3563,I106217,I106206,);
nand I_6051 (I106463,I778077,I778068);
and I_6052 (I106480,I106463,I778083);
DFFARX1 I_6053 (I106480,I3563,I106217,I106506,);
DFFARX1 I_6054 (I106506,I3563,I106217,I106523,);
not I_6055 (I106209,I106523);
not I_6056 (I106545,I106506);
nand I_6057 (I106194,I106545,I106384);
nor I_6058 (I106576,I778074,I778068);
not I_6059 (I106593,I106576);
nor I_6060 (I106610,I106545,I106593);
nor I_6061 (I106627,I106251,I106610);
DFFARX1 I_6062 (I106627,I3563,I106217,I106203,);
nor I_6063 (I106658,I106311,I106593);
nor I_6064 (I106191,I106506,I106658);
nor I_6065 (I106200,I106441,I106576);
nor I_6066 (I106188,I106311,I106576);
not I_6067 (I106744,I3570);
DFFARX1 I_6068 (I669985,I3563,I106744,I106770,);
not I_6069 (I106778,I106770);
nand I_6070 (I106795,I669976,I669994);
and I_6071 (I106812,I106795,I669973);
DFFARX1 I_6072 (I106812,I3563,I106744,I106838,);
DFFARX1 I_6073 (I669976,I3563,I106744,I106855,);
and I_6074 (I106863,I106855,I669979);
nor I_6075 (I106880,I106838,I106863);
DFFARX1 I_6076 (I106880,I3563,I106744,I106712,);
nand I_6077 (I106911,I106855,I669979);
nand I_6078 (I106928,I106778,I106911);
not I_6079 (I106724,I106928);
DFFARX1 I_6080 (I669973,I3563,I106744,I106968,);
DFFARX1 I_6081 (I106968,I3563,I106744,I106733,);
nand I_6082 (I106990,I669991,I669982);
and I_6083 (I107007,I106990,I669997);
DFFARX1 I_6084 (I107007,I3563,I106744,I107033,);
DFFARX1 I_6085 (I107033,I3563,I106744,I107050,);
not I_6086 (I106736,I107050);
not I_6087 (I107072,I107033);
nand I_6088 (I106721,I107072,I106911);
nor I_6089 (I107103,I669988,I669982);
not I_6090 (I107120,I107103);
nor I_6091 (I107137,I107072,I107120);
nor I_6092 (I107154,I106778,I107137);
DFFARX1 I_6093 (I107154,I3563,I106744,I106730,);
nor I_6094 (I107185,I106838,I107120);
nor I_6095 (I106718,I107033,I107185);
nor I_6096 (I106727,I106968,I107103);
nor I_6097 (I106715,I106838,I107103);
not I_6098 (I107271,I3570);
DFFARX1 I_6099 (I517620,I3563,I107271,I107297,);
not I_6100 (I107305,I107297);
nand I_6101 (I107322,I517614,I517605);
and I_6102 (I107339,I107322,I517626);
DFFARX1 I_6103 (I107339,I3563,I107271,I107365,);
DFFARX1 I_6104 (I517608,I3563,I107271,I107382,);
and I_6105 (I107390,I107382,I517602);
nor I_6106 (I107407,I107365,I107390);
DFFARX1 I_6107 (I107407,I3563,I107271,I107239,);
nand I_6108 (I107438,I107382,I517602);
nand I_6109 (I107455,I107305,I107438);
not I_6110 (I107251,I107455);
DFFARX1 I_6111 (I517602,I3563,I107271,I107495,);
DFFARX1 I_6112 (I107495,I3563,I107271,I107260,);
nand I_6113 (I107517,I517629,I517611);
and I_6114 (I107534,I107517,I517617);
DFFARX1 I_6115 (I107534,I3563,I107271,I107560,);
DFFARX1 I_6116 (I107560,I3563,I107271,I107577,);
not I_6117 (I107263,I107577);
not I_6118 (I107599,I107560);
nand I_6119 (I107248,I107599,I107438);
nor I_6120 (I107630,I517623,I517611);
not I_6121 (I107647,I107630);
nor I_6122 (I107664,I107599,I107647);
nor I_6123 (I107681,I107305,I107664);
DFFARX1 I_6124 (I107681,I3563,I107271,I107257,);
nor I_6125 (I107712,I107365,I107647);
nor I_6126 (I107245,I107560,I107712);
nor I_6127 (I107254,I107495,I107630);
nor I_6128 (I107242,I107365,I107630);
not I_6129 (I107798,I3570);
DFFARX1 I_6130 (I333876,I3563,I107798,I107824,);
not I_6131 (I107832,I107824);
nand I_6132 (I107849,I333858,I333873);
and I_6133 (I107866,I107849,I333849);
DFFARX1 I_6134 (I107866,I3563,I107798,I107892,);
DFFARX1 I_6135 (I333852,I3563,I107798,I107909,);
and I_6136 (I107917,I107909,I333867);
nor I_6137 (I107934,I107892,I107917);
DFFARX1 I_6138 (I107934,I3563,I107798,I107766,);
nand I_6139 (I107965,I107909,I333867);
nand I_6140 (I107982,I107832,I107965);
not I_6141 (I107778,I107982);
DFFARX1 I_6142 (I333870,I3563,I107798,I108022,);
DFFARX1 I_6143 (I108022,I3563,I107798,I107787,);
nand I_6144 (I108044,I333849,I333861);
and I_6145 (I108061,I108044,I333855);
DFFARX1 I_6146 (I108061,I3563,I107798,I108087,);
DFFARX1 I_6147 (I108087,I3563,I107798,I108104,);
not I_6148 (I107790,I108104);
not I_6149 (I108126,I108087);
nand I_6150 (I107775,I108126,I107965);
nor I_6151 (I108157,I333864,I333861);
not I_6152 (I108174,I108157);
nor I_6153 (I108191,I108126,I108174);
nor I_6154 (I108208,I107832,I108191);
DFFARX1 I_6155 (I108208,I3563,I107798,I107784,);
nor I_6156 (I108239,I107892,I108174);
nor I_6157 (I107772,I108087,I108239);
nor I_6158 (I107781,I108022,I108157);
nor I_6159 (I107769,I107892,I108157);
not I_6160 (I108325,I3570);
DFFARX1 I_6161 (I49820,I3563,I108325,I108351,);
not I_6162 (I108359,I108351);
nand I_6163 (I108376,I49808,I49814);
and I_6164 (I108393,I108376,I49817);
DFFARX1 I_6165 (I108393,I3563,I108325,I108419,);
DFFARX1 I_6166 (I49799,I3563,I108325,I108436,);
and I_6167 (I108444,I108436,I49805);
nor I_6168 (I108461,I108419,I108444);
DFFARX1 I_6169 (I108461,I3563,I108325,I108293,);
nand I_6170 (I108492,I108436,I49805);
nand I_6171 (I108509,I108359,I108492);
not I_6172 (I108305,I108509);
DFFARX1 I_6173 (I49799,I3563,I108325,I108549,);
DFFARX1 I_6174 (I108549,I3563,I108325,I108314,);
nand I_6175 (I108571,I49802,I49796);
and I_6176 (I108588,I108571,I49811);
DFFARX1 I_6177 (I108588,I3563,I108325,I108614,);
DFFARX1 I_6178 (I108614,I3563,I108325,I108631,);
not I_6179 (I108317,I108631);
not I_6180 (I108653,I108614);
nand I_6181 (I108302,I108653,I108492);
nor I_6182 (I108684,I49796,I49796);
not I_6183 (I108701,I108684);
nor I_6184 (I108718,I108653,I108701);
nor I_6185 (I108735,I108359,I108718);
DFFARX1 I_6186 (I108735,I3563,I108325,I108311,);
nor I_6187 (I108766,I108419,I108701);
nor I_6188 (I108299,I108614,I108766);
nor I_6189 (I108308,I108549,I108684);
nor I_6190 (I108296,I108419,I108684);
not I_6191 (I108852,I3570);
DFFARX1 I_6192 (I1031164,I3563,I108852,I108878,);
not I_6193 (I108886,I108878);
nand I_6194 (I108903,I1031182,I1031176);
and I_6195 (I108920,I108903,I1031155);
DFFARX1 I_6196 (I108920,I3563,I108852,I108946,);
DFFARX1 I_6197 (I1031173,I3563,I108852,I108963,);
and I_6198 (I108971,I108963,I1031158);
nor I_6199 (I108988,I108946,I108971);
DFFARX1 I_6200 (I108988,I3563,I108852,I108820,);
nand I_6201 (I109019,I108963,I1031158);
nand I_6202 (I109036,I108886,I109019);
not I_6203 (I108832,I109036);
DFFARX1 I_6204 (I1031170,I3563,I108852,I109076,);
DFFARX1 I_6205 (I109076,I3563,I108852,I108841,);
nand I_6206 (I109098,I1031179,I1031167);
and I_6207 (I109115,I109098,I1031161);
DFFARX1 I_6208 (I109115,I3563,I108852,I109141,);
DFFARX1 I_6209 (I109141,I3563,I108852,I109158,);
not I_6210 (I108844,I109158);
not I_6211 (I109180,I109141);
nand I_6212 (I108829,I109180,I109019);
nor I_6213 (I109211,I1031155,I1031167);
not I_6214 (I109228,I109211);
nor I_6215 (I109245,I109180,I109228);
nor I_6216 (I109262,I108886,I109245);
DFFARX1 I_6217 (I109262,I3563,I108852,I108838,);
nor I_6218 (I109293,I108946,I109228);
nor I_6219 (I108826,I109141,I109293);
nor I_6220 (I108835,I109076,I109211);
nor I_6221 (I108823,I108946,I109211);
not I_6222 (I109379,I3570);
DFFARX1 I_6223 (I1394015,I3563,I109379,I109405,);
not I_6224 (I109413,I109405);
nand I_6225 (I109430,I1394009,I1394030);
and I_6226 (I109447,I109430,I1394006);
DFFARX1 I_6227 (I109447,I3563,I109379,I109473,);
DFFARX1 I_6228 (I1394027,I3563,I109379,I109490,);
and I_6229 (I109498,I109490,I1394024);
nor I_6230 (I109515,I109473,I109498);
DFFARX1 I_6231 (I109515,I3563,I109379,I109347,);
nand I_6232 (I109546,I109490,I1394024);
nand I_6233 (I109563,I109413,I109546);
not I_6234 (I109359,I109563);
DFFARX1 I_6235 (I1394012,I3563,I109379,I109603,);
DFFARX1 I_6236 (I109603,I3563,I109379,I109368,);
nand I_6237 (I109625,I1394021,I1394018);
and I_6238 (I109642,I109625,I1394003);
DFFARX1 I_6239 (I109642,I3563,I109379,I109668,);
DFFARX1 I_6240 (I109668,I3563,I109379,I109685,);
not I_6241 (I109371,I109685);
not I_6242 (I109707,I109668);
nand I_6243 (I109356,I109707,I109546);
nor I_6244 (I109738,I1394003,I1394018);
not I_6245 (I109755,I109738);
nor I_6246 (I109772,I109707,I109755);
nor I_6247 (I109789,I109413,I109772);
DFFARX1 I_6248 (I109789,I3563,I109379,I109365,);
nor I_6249 (I109820,I109473,I109755);
nor I_6250 (I109353,I109668,I109820);
nor I_6251 (I109362,I109603,I109738);
nor I_6252 (I109350,I109473,I109738);
not I_6253 (I109906,I3570);
DFFARX1 I_6254 (I638770,I3563,I109906,I109932,);
not I_6255 (I109940,I109932);
nand I_6256 (I109957,I638782,I638767);
and I_6257 (I109974,I109957,I638761);
DFFARX1 I_6258 (I109974,I3563,I109906,I110000,);
DFFARX1 I_6259 (I638776,I3563,I109906,I110017,);
and I_6260 (I110025,I110017,I638764);
nor I_6261 (I110042,I110000,I110025);
DFFARX1 I_6262 (I110042,I3563,I109906,I109874,);
nand I_6263 (I110073,I110017,I638764);
nand I_6264 (I110090,I109940,I110073);
not I_6265 (I109886,I110090);
DFFARX1 I_6266 (I638773,I3563,I109906,I110130,);
DFFARX1 I_6267 (I110130,I3563,I109906,I109895,);
nand I_6268 (I110152,I638779,I638785);
and I_6269 (I110169,I110152,I638761);
DFFARX1 I_6270 (I110169,I3563,I109906,I110195,);
DFFARX1 I_6271 (I110195,I3563,I109906,I110212,);
not I_6272 (I109898,I110212);
not I_6273 (I110234,I110195);
nand I_6274 (I109883,I110234,I110073);
nor I_6275 (I110265,I638764,I638785);
not I_6276 (I110282,I110265);
nor I_6277 (I110299,I110234,I110282);
nor I_6278 (I110316,I109940,I110299);
DFFARX1 I_6279 (I110316,I3563,I109906,I109892,);
nor I_6280 (I110347,I110000,I110282);
nor I_6281 (I109880,I110195,I110347);
nor I_6282 (I109889,I110130,I110265);
nor I_6283 (I109877,I110000,I110265);
not I_6284 (I110433,I3570);
DFFARX1 I_6285 (I168485,I3563,I110433,I110459,);
not I_6286 (I110467,I110459);
nand I_6287 (I110484,I168479,I168473);
and I_6288 (I110501,I110484,I168494);
DFFARX1 I_6289 (I110501,I3563,I110433,I110527,);
DFFARX1 I_6290 (I168491,I3563,I110433,I110544,);
and I_6291 (I110552,I110544,I168488);
nor I_6292 (I110569,I110527,I110552);
DFFARX1 I_6293 (I110569,I3563,I110433,I110401,);
nand I_6294 (I110600,I110544,I168488);
nand I_6295 (I110617,I110467,I110600);
not I_6296 (I110413,I110617);
DFFARX1 I_6297 (I168473,I3563,I110433,I110657,);
DFFARX1 I_6298 (I110657,I3563,I110433,I110422,);
nand I_6299 (I110679,I168476,I168476);
and I_6300 (I110696,I110679,I168497);
DFFARX1 I_6301 (I110696,I3563,I110433,I110722,);
DFFARX1 I_6302 (I110722,I3563,I110433,I110739,);
not I_6303 (I110425,I110739);
not I_6304 (I110761,I110722);
nand I_6305 (I110410,I110761,I110600);
nor I_6306 (I110792,I168482,I168476);
not I_6307 (I110809,I110792);
nor I_6308 (I110826,I110761,I110809);
nor I_6309 (I110843,I110467,I110826);
DFFARX1 I_6310 (I110843,I3563,I110433,I110419,);
nor I_6311 (I110874,I110527,I110809);
nor I_6312 (I110407,I110722,I110874);
nor I_6313 (I110416,I110657,I110792);
nor I_6314 (I110404,I110527,I110792);
not I_6315 (I110960,I3570);
DFFARX1 I_6316 (I985944,I3563,I110960,I110986,);
not I_6317 (I110994,I110986);
nand I_6318 (I111011,I985962,I985956);
and I_6319 (I111028,I111011,I985935);
DFFARX1 I_6320 (I111028,I3563,I110960,I111054,);
DFFARX1 I_6321 (I985953,I3563,I110960,I111071,);
and I_6322 (I111079,I111071,I985938);
nor I_6323 (I111096,I111054,I111079);
DFFARX1 I_6324 (I111096,I3563,I110960,I110928,);
nand I_6325 (I111127,I111071,I985938);
nand I_6326 (I111144,I110994,I111127);
not I_6327 (I110940,I111144);
DFFARX1 I_6328 (I985950,I3563,I110960,I111184,);
DFFARX1 I_6329 (I111184,I3563,I110960,I110949,);
nand I_6330 (I111206,I985959,I985947);
and I_6331 (I111223,I111206,I985941);
DFFARX1 I_6332 (I111223,I3563,I110960,I111249,);
DFFARX1 I_6333 (I111249,I3563,I110960,I111266,);
not I_6334 (I110952,I111266);
not I_6335 (I111288,I111249);
nand I_6336 (I110937,I111288,I111127);
nor I_6337 (I111319,I985935,I985947);
not I_6338 (I111336,I111319);
nor I_6339 (I111353,I111288,I111336);
nor I_6340 (I111370,I110994,I111353);
DFFARX1 I_6341 (I111370,I3563,I110960,I110946,);
nor I_6342 (I111401,I111054,I111336);
nor I_6343 (I110934,I111249,I111401);
nor I_6344 (I110943,I111184,I111319);
nor I_6345 (I110931,I111054,I111319);
not I_6346 (I111487,I3570);
DFFARX1 I_6347 (I1178857,I3563,I111487,I111513,);
not I_6348 (I111521,I111513);
nand I_6349 (I111538,I1178872,I1178851);
and I_6350 (I111555,I111538,I1178854);
DFFARX1 I_6351 (I111555,I3563,I111487,I111581,);
DFFARX1 I_6352 (I1178875,I3563,I111487,I111598,);
and I_6353 (I111606,I111598,I1178854);
nor I_6354 (I111623,I111581,I111606);
DFFARX1 I_6355 (I111623,I3563,I111487,I111455,);
nand I_6356 (I111654,I111598,I1178854);
nand I_6357 (I111671,I111521,I111654);
not I_6358 (I111467,I111671);
DFFARX1 I_6359 (I1178851,I3563,I111487,I111711,);
DFFARX1 I_6360 (I111711,I3563,I111487,I111476,);
nand I_6361 (I111733,I1178863,I1178860);
and I_6362 (I111750,I111733,I1178866);
DFFARX1 I_6363 (I111750,I3563,I111487,I111776,);
DFFARX1 I_6364 (I111776,I3563,I111487,I111793,);
not I_6365 (I111479,I111793);
not I_6366 (I111815,I111776);
nand I_6367 (I111464,I111815,I111654);
nor I_6368 (I111846,I1178869,I1178860);
not I_6369 (I111863,I111846);
nor I_6370 (I111880,I111815,I111863);
nor I_6371 (I111897,I111521,I111880);
DFFARX1 I_6372 (I111897,I3563,I111487,I111473,);
nor I_6373 (I111928,I111581,I111863);
nor I_6374 (I111461,I111776,I111928);
nor I_6375 (I111470,I111711,I111846);
nor I_6376 (I111458,I111581,I111846);
not I_6377 (I112014,I3570);
DFFARX1 I_6378 (I1240125,I3563,I112014,I112040,);
not I_6379 (I112048,I112040);
nand I_6380 (I112065,I1240140,I1240119);
and I_6381 (I112082,I112065,I1240122);
DFFARX1 I_6382 (I112082,I3563,I112014,I112108,);
DFFARX1 I_6383 (I1240143,I3563,I112014,I112125,);
and I_6384 (I112133,I112125,I1240122);
nor I_6385 (I112150,I112108,I112133);
DFFARX1 I_6386 (I112150,I3563,I112014,I111982,);
nand I_6387 (I112181,I112125,I1240122);
nand I_6388 (I112198,I112048,I112181);
not I_6389 (I111994,I112198);
DFFARX1 I_6390 (I1240119,I3563,I112014,I112238,);
DFFARX1 I_6391 (I112238,I3563,I112014,I112003,);
nand I_6392 (I112260,I1240131,I1240128);
and I_6393 (I112277,I112260,I1240134);
DFFARX1 I_6394 (I112277,I3563,I112014,I112303,);
DFFARX1 I_6395 (I112303,I3563,I112014,I112320,);
not I_6396 (I112006,I112320);
not I_6397 (I112342,I112303);
nand I_6398 (I111991,I112342,I112181);
nor I_6399 (I112373,I1240137,I1240128);
not I_6400 (I112390,I112373);
nor I_6401 (I112407,I112342,I112390);
nor I_6402 (I112424,I112048,I112407);
DFFARX1 I_6403 (I112424,I3563,I112014,I112000,);
nor I_6404 (I112455,I112108,I112390);
nor I_6405 (I111988,I112303,I112455);
nor I_6406 (I111997,I112238,I112373);
nor I_6407 (I111985,I112108,I112373);
not I_6408 (I112541,I3570);
DFFARX1 I_6409 (I787897,I3563,I112541,I112567,);
not I_6410 (I112575,I112567);
nand I_6411 (I112592,I787888,I787906);
and I_6412 (I112609,I112592,I787885);
DFFARX1 I_6413 (I112609,I3563,I112541,I112635,);
DFFARX1 I_6414 (I787888,I3563,I112541,I112652,);
and I_6415 (I112660,I112652,I787891);
nor I_6416 (I112677,I112635,I112660);
DFFARX1 I_6417 (I112677,I3563,I112541,I112509,);
nand I_6418 (I112708,I112652,I787891);
nand I_6419 (I112725,I112575,I112708);
not I_6420 (I112521,I112725);
DFFARX1 I_6421 (I787885,I3563,I112541,I112765,);
DFFARX1 I_6422 (I112765,I3563,I112541,I112530,);
nand I_6423 (I112787,I787903,I787894);
and I_6424 (I112804,I112787,I787909);
DFFARX1 I_6425 (I112804,I3563,I112541,I112830,);
DFFARX1 I_6426 (I112830,I3563,I112541,I112847,);
not I_6427 (I112533,I112847);
not I_6428 (I112869,I112830);
nand I_6429 (I112518,I112869,I112708);
nor I_6430 (I112900,I787900,I787894);
not I_6431 (I112917,I112900);
nor I_6432 (I112934,I112869,I112917);
nor I_6433 (I112951,I112575,I112934);
DFFARX1 I_6434 (I112951,I3563,I112541,I112527,);
nor I_6435 (I112982,I112635,I112917);
nor I_6436 (I112515,I112830,I112982);
nor I_6437 (I112524,I112765,I112900);
nor I_6438 (I112512,I112635,I112900);
not I_6439 (I113068,I3570);
DFFARX1 I_6440 (I277370,I3563,I113068,I113094,);
not I_6441 (I113102,I113094);
nand I_6442 (I113119,I277364,I277358);
and I_6443 (I113136,I113119,I277379);
DFFARX1 I_6444 (I113136,I3563,I113068,I113162,);
DFFARX1 I_6445 (I277376,I3563,I113068,I113179,);
and I_6446 (I113187,I113179,I277373);
nor I_6447 (I113204,I113162,I113187);
DFFARX1 I_6448 (I113204,I3563,I113068,I113036,);
nand I_6449 (I113235,I113179,I277373);
nand I_6450 (I113252,I113102,I113235);
not I_6451 (I113048,I113252);
DFFARX1 I_6452 (I277358,I3563,I113068,I113292,);
DFFARX1 I_6453 (I113292,I3563,I113068,I113057,);
nand I_6454 (I113314,I277361,I277361);
and I_6455 (I113331,I113314,I277382);
DFFARX1 I_6456 (I113331,I3563,I113068,I113357,);
DFFARX1 I_6457 (I113357,I3563,I113068,I113374,);
not I_6458 (I113060,I113374);
not I_6459 (I113396,I113357);
nand I_6460 (I113045,I113396,I113235);
nor I_6461 (I113427,I277367,I277361);
not I_6462 (I113444,I113427);
nor I_6463 (I113461,I113396,I113444);
nor I_6464 (I113478,I113102,I113461);
DFFARX1 I_6465 (I113478,I3563,I113068,I113054,);
nor I_6466 (I113509,I113162,I113444);
nor I_6467 (I113042,I113357,I113509);
nor I_6468 (I113051,I113292,I113427);
nor I_6469 (I113039,I113162,I113427);
not I_6470 (I113595,I3570);
DFFARX1 I_6471 (I1329777,I3563,I113595,I113621,);
not I_6472 (I113629,I113621);
nand I_6473 (I113646,I1329783,I1329801);
and I_6474 (I113663,I113646,I1329798);
DFFARX1 I_6475 (I113663,I3563,I113595,I113689,);
DFFARX1 I_6476 (I1329795,I3563,I113595,I113706,);
and I_6477 (I113714,I113706,I1329789);
nor I_6478 (I113731,I113689,I113714);
DFFARX1 I_6479 (I113731,I3563,I113595,I113563,);
nand I_6480 (I113762,I113706,I1329789);
nand I_6481 (I113779,I113629,I113762);
not I_6482 (I113575,I113779);
DFFARX1 I_6483 (I1329777,I3563,I113595,I113819,);
DFFARX1 I_6484 (I113819,I3563,I113595,I113584,);
nand I_6485 (I113841,I1329792,I1329780);
and I_6486 (I113858,I113841,I1329804);
DFFARX1 I_6487 (I113858,I3563,I113595,I113884,);
DFFARX1 I_6488 (I113884,I3563,I113595,I113901,);
not I_6489 (I113587,I113901);
not I_6490 (I113923,I113884);
nand I_6491 (I113572,I113923,I113762);
nor I_6492 (I113954,I1329786,I1329780);
not I_6493 (I113971,I113954);
nor I_6494 (I113988,I113923,I113971);
nor I_6495 (I114005,I113629,I113988);
DFFARX1 I_6496 (I114005,I3563,I113595,I113581,);
nor I_6497 (I114036,I113689,I113971);
nor I_6498 (I113569,I113884,I114036);
nor I_6499 (I113578,I113819,I113954);
nor I_6500 (I113566,I113689,I113954);
not I_6501 (I114122,I3570);
DFFARX1 I_6502 (I633568,I3563,I114122,I114148,);
not I_6503 (I114156,I114148);
nand I_6504 (I114173,I633580,I633565);
and I_6505 (I114190,I114173,I633559);
DFFARX1 I_6506 (I114190,I3563,I114122,I114216,);
DFFARX1 I_6507 (I633574,I3563,I114122,I114233,);
and I_6508 (I114241,I114233,I633562);
nor I_6509 (I114258,I114216,I114241);
DFFARX1 I_6510 (I114258,I3563,I114122,I114090,);
nand I_6511 (I114289,I114233,I633562);
nand I_6512 (I114306,I114156,I114289);
not I_6513 (I114102,I114306);
DFFARX1 I_6514 (I633571,I3563,I114122,I114346,);
DFFARX1 I_6515 (I114346,I3563,I114122,I114111,);
nand I_6516 (I114368,I633577,I633583);
and I_6517 (I114385,I114368,I633559);
DFFARX1 I_6518 (I114385,I3563,I114122,I114411,);
DFFARX1 I_6519 (I114411,I3563,I114122,I114428,);
not I_6520 (I114114,I114428);
not I_6521 (I114450,I114411);
nand I_6522 (I114099,I114450,I114289);
nor I_6523 (I114481,I633562,I633583);
not I_6524 (I114498,I114481);
nor I_6525 (I114515,I114450,I114498);
nor I_6526 (I114532,I114156,I114515);
DFFARX1 I_6527 (I114532,I3563,I114122,I114108,);
nor I_6528 (I114563,I114216,I114498);
nor I_6529 (I114096,I114411,I114563);
nor I_6530 (I114105,I114346,I114481);
nor I_6531 (I114093,I114216,I114481);
not I_6532 (I114649,I3570);
DFFARX1 I_6533 (I908560,I3563,I114649,I114675,);
not I_6534 (I114683,I114675);
nand I_6535 (I114700,I908557,I908572);
and I_6536 (I114717,I114700,I908554);
DFFARX1 I_6537 (I114717,I3563,I114649,I114743,);
DFFARX1 I_6538 (I908551,I3563,I114649,I114760,);
and I_6539 (I114768,I114760,I908551);
nor I_6540 (I114785,I114743,I114768);
DFFARX1 I_6541 (I114785,I3563,I114649,I114617,);
nand I_6542 (I114816,I114760,I908551);
nand I_6543 (I114833,I114683,I114816);
not I_6544 (I114629,I114833);
DFFARX1 I_6545 (I908554,I3563,I114649,I114873,);
DFFARX1 I_6546 (I114873,I3563,I114649,I114638,);
nand I_6547 (I114895,I908566,I908557);
and I_6548 (I114912,I114895,I908569);
DFFARX1 I_6549 (I114912,I3563,I114649,I114938,);
DFFARX1 I_6550 (I114938,I3563,I114649,I114955,);
not I_6551 (I114641,I114955);
not I_6552 (I114977,I114938);
nand I_6553 (I114626,I114977,I114816);
nor I_6554 (I115008,I908563,I908557);
not I_6555 (I115025,I115008);
nor I_6556 (I115042,I114977,I115025);
nor I_6557 (I115059,I114683,I115042);
DFFARX1 I_6558 (I115059,I3563,I114649,I114635,);
nor I_6559 (I115090,I114743,I115025);
nor I_6560 (I114623,I114938,I115090);
nor I_6561 (I114632,I114873,I115008);
nor I_6562 (I114620,I114743,I115008);
not I_6563 (I115176,I3570);
DFFARX1 I_6564 (I365496,I3563,I115176,I115202,);
not I_6565 (I115210,I115202);
nand I_6566 (I115227,I365478,I365493);
and I_6567 (I115244,I115227,I365469);
DFFARX1 I_6568 (I115244,I3563,I115176,I115270,);
DFFARX1 I_6569 (I365472,I3563,I115176,I115287,);
and I_6570 (I115295,I115287,I365487);
nor I_6571 (I115312,I115270,I115295);
DFFARX1 I_6572 (I115312,I3563,I115176,I115144,);
nand I_6573 (I115343,I115287,I365487);
nand I_6574 (I115360,I115210,I115343);
not I_6575 (I115156,I115360);
DFFARX1 I_6576 (I365490,I3563,I115176,I115400,);
DFFARX1 I_6577 (I115400,I3563,I115176,I115165,);
nand I_6578 (I115422,I365469,I365481);
and I_6579 (I115439,I115422,I365475);
DFFARX1 I_6580 (I115439,I3563,I115176,I115465,);
DFFARX1 I_6581 (I115465,I3563,I115176,I115482,);
not I_6582 (I115168,I115482);
not I_6583 (I115504,I115465);
nand I_6584 (I115153,I115504,I115343);
nor I_6585 (I115535,I365484,I365481);
not I_6586 (I115552,I115535);
nor I_6587 (I115569,I115504,I115552);
nor I_6588 (I115586,I115210,I115569);
DFFARX1 I_6589 (I115586,I3563,I115176,I115162,);
nor I_6590 (I115617,I115270,I115552);
nor I_6591 (I115150,I115465,I115617);
nor I_6592 (I115159,I115400,I115535);
nor I_6593 (I115147,I115270,I115535);
not I_6594 (I115703,I3570);
DFFARX1 I_6595 (I466484,I3563,I115703,I115729,);
not I_6596 (I115737,I115729);
nand I_6597 (I115754,I466478,I466469);
and I_6598 (I115771,I115754,I466490);
DFFARX1 I_6599 (I115771,I3563,I115703,I115797,);
DFFARX1 I_6600 (I466472,I3563,I115703,I115814,);
and I_6601 (I115822,I115814,I466466);
nor I_6602 (I115839,I115797,I115822);
DFFARX1 I_6603 (I115839,I3563,I115703,I115671,);
nand I_6604 (I115870,I115814,I466466);
nand I_6605 (I115887,I115737,I115870);
not I_6606 (I115683,I115887);
DFFARX1 I_6607 (I466466,I3563,I115703,I115927,);
DFFARX1 I_6608 (I115927,I3563,I115703,I115692,);
nand I_6609 (I115949,I466493,I466475);
and I_6610 (I115966,I115949,I466481);
DFFARX1 I_6611 (I115966,I3563,I115703,I115992,);
DFFARX1 I_6612 (I115992,I3563,I115703,I116009,);
not I_6613 (I115695,I116009);
not I_6614 (I116031,I115992);
nand I_6615 (I115680,I116031,I115870);
nor I_6616 (I116062,I466487,I466475);
not I_6617 (I116079,I116062);
nor I_6618 (I116096,I116031,I116079);
nor I_6619 (I116113,I115737,I116096);
DFFARX1 I_6620 (I116113,I3563,I115703,I115689,);
nor I_6621 (I116144,I115797,I116079);
nor I_6622 (I115677,I115992,I116144);
nor I_6623 (I115686,I115927,I116062);
nor I_6624 (I115674,I115797,I116062);
not I_6625 (I116230,I3570);
DFFARX1 I_6626 (I361280,I3563,I116230,I116256,);
not I_6627 (I116264,I116256);
nand I_6628 (I116281,I361262,I361277);
and I_6629 (I116298,I116281,I361253);
DFFARX1 I_6630 (I116298,I3563,I116230,I116324,);
DFFARX1 I_6631 (I361256,I3563,I116230,I116341,);
and I_6632 (I116349,I116341,I361271);
nor I_6633 (I116366,I116324,I116349);
DFFARX1 I_6634 (I116366,I3563,I116230,I116198,);
nand I_6635 (I116397,I116341,I361271);
nand I_6636 (I116414,I116264,I116397);
not I_6637 (I116210,I116414);
DFFARX1 I_6638 (I361274,I3563,I116230,I116454,);
DFFARX1 I_6639 (I116454,I3563,I116230,I116219,);
nand I_6640 (I116476,I361253,I361265);
and I_6641 (I116493,I116476,I361259);
DFFARX1 I_6642 (I116493,I3563,I116230,I116519,);
DFFARX1 I_6643 (I116519,I3563,I116230,I116536,);
not I_6644 (I116222,I116536);
not I_6645 (I116558,I116519);
nand I_6646 (I116207,I116558,I116397);
nor I_6647 (I116589,I361268,I361265);
not I_6648 (I116606,I116589);
nor I_6649 (I116623,I116558,I116606);
nor I_6650 (I116640,I116264,I116623);
DFFARX1 I_6651 (I116640,I3563,I116230,I116216,);
nor I_6652 (I116671,I116324,I116606);
nor I_6653 (I116204,I116519,I116671);
nor I_6654 (I116213,I116454,I116589);
nor I_6655 (I116201,I116324,I116589);
not I_6656 (I116757,I3570);
DFFARX1 I_6657 (I1065736,I3563,I116757,I116783,);
not I_6658 (I116791,I116783);
nand I_6659 (I116808,I1065733,I1065739);
and I_6660 (I116825,I116808,I1065736);
DFFARX1 I_6661 (I116825,I3563,I116757,I116851,);
DFFARX1 I_6662 (I1065739,I3563,I116757,I116868,);
and I_6663 (I116876,I116868,I1065733);
nor I_6664 (I116893,I116851,I116876);
DFFARX1 I_6665 (I116893,I3563,I116757,I116725,);
nand I_6666 (I116924,I116868,I1065733);
nand I_6667 (I116941,I116791,I116924);
not I_6668 (I116737,I116941);
DFFARX1 I_6669 (I1065742,I3563,I116757,I116981,);
DFFARX1 I_6670 (I116981,I3563,I116757,I116746,);
nand I_6671 (I117003,I1065745,I1065754);
and I_6672 (I117020,I117003,I1065748);
DFFARX1 I_6673 (I117020,I3563,I116757,I117046,);
DFFARX1 I_6674 (I117046,I3563,I116757,I117063,);
not I_6675 (I116749,I117063);
not I_6676 (I117085,I117046);
nand I_6677 (I116734,I117085,I116924);
nor I_6678 (I117116,I1065751,I1065754);
not I_6679 (I117133,I117116);
nor I_6680 (I117150,I117085,I117133);
nor I_6681 (I117167,I116791,I117150);
DFFARX1 I_6682 (I117167,I3563,I116757,I116743,);
nor I_6683 (I117198,I116851,I117133);
nor I_6684 (I116731,I117046,I117198);
nor I_6685 (I116740,I116981,I117116);
nor I_6686 (I116728,I116851,I117116);
not I_6687 (I117284,I3570);
DFFARX1 I_6688 (I562604,I3563,I117284,I117310,);
not I_6689 (I117318,I117310);
nand I_6690 (I117335,I562625,I562619);
and I_6691 (I117352,I117335,I562601);
DFFARX1 I_6692 (I117352,I3563,I117284,I117378,);
DFFARX1 I_6693 (I562604,I3563,I117284,I117395,);
and I_6694 (I117403,I117395,I562613);
nor I_6695 (I117420,I117378,I117403);
DFFARX1 I_6696 (I117420,I3563,I117284,I117252,);
nand I_6697 (I117451,I117395,I562613);
nand I_6698 (I117468,I117318,I117451);
not I_6699 (I117264,I117468);
DFFARX1 I_6700 (I562610,I3563,I117284,I117508,);
DFFARX1 I_6701 (I117508,I3563,I117284,I117273,);
nand I_6702 (I117530,I562616,I562607);
and I_6703 (I117547,I117530,I562601);
DFFARX1 I_6704 (I117547,I3563,I117284,I117573,);
DFFARX1 I_6705 (I117573,I3563,I117284,I117590,);
not I_6706 (I117276,I117590);
not I_6707 (I117612,I117573);
nand I_6708 (I117261,I117612,I117451);
nor I_6709 (I117643,I562622,I562607);
not I_6710 (I117660,I117643);
nor I_6711 (I117677,I117612,I117660);
nor I_6712 (I117694,I117318,I117677);
DFFARX1 I_6713 (I117694,I3563,I117284,I117270,);
nor I_6714 (I117725,I117378,I117660);
nor I_6715 (I117258,I117573,I117725);
nor I_6716 (I117267,I117508,I117643);
nor I_6717 (I117255,I117378,I117643);
not I_6718 (I117811,I3570);
DFFARX1 I_6719 (I322809,I3563,I117811,I117837,);
not I_6720 (I117845,I117837);
nand I_6721 (I117862,I322791,I322806);
and I_6722 (I117879,I117862,I322782);
DFFARX1 I_6723 (I117879,I3563,I117811,I117905,);
DFFARX1 I_6724 (I322785,I3563,I117811,I117922,);
and I_6725 (I117930,I117922,I322800);
nor I_6726 (I117947,I117905,I117930);
DFFARX1 I_6727 (I117947,I3563,I117811,I117779,);
nand I_6728 (I117978,I117922,I322800);
nand I_6729 (I117995,I117845,I117978);
not I_6730 (I117791,I117995);
DFFARX1 I_6731 (I322803,I3563,I117811,I118035,);
DFFARX1 I_6732 (I118035,I3563,I117811,I117800,);
nand I_6733 (I118057,I322782,I322794);
and I_6734 (I118074,I118057,I322788);
DFFARX1 I_6735 (I118074,I3563,I117811,I118100,);
DFFARX1 I_6736 (I118100,I3563,I117811,I118117,);
not I_6737 (I117803,I118117);
not I_6738 (I118139,I118100);
nand I_6739 (I117788,I118139,I117978);
nor I_6740 (I118170,I322797,I322794);
not I_6741 (I118187,I118170);
nor I_6742 (I118204,I118139,I118187);
nor I_6743 (I118221,I117845,I118204);
DFFARX1 I_6744 (I118221,I3563,I117811,I117797,);
nor I_6745 (I118252,I117905,I118187);
nor I_6746 (I117785,I118100,I118252);
nor I_6747 (I117794,I118035,I118170);
nor I_6748 (I117782,I117905,I118170);
not I_6749 (I118338,I3570);
DFFARX1 I_6750 (I671141,I3563,I118338,I118364,);
not I_6751 (I118372,I118364);
nand I_6752 (I118389,I671132,I671150);
and I_6753 (I118406,I118389,I671129);
DFFARX1 I_6754 (I118406,I3563,I118338,I118432,);
DFFARX1 I_6755 (I671132,I3563,I118338,I118449,);
and I_6756 (I118457,I118449,I671135);
nor I_6757 (I118474,I118432,I118457);
DFFARX1 I_6758 (I118474,I3563,I118338,I118306,);
nand I_6759 (I118505,I118449,I671135);
nand I_6760 (I118522,I118372,I118505);
not I_6761 (I118318,I118522);
DFFARX1 I_6762 (I671129,I3563,I118338,I118562,);
DFFARX1 I_6763 (I118562,I3563,I118338,I118327,);
nand I_6764 (I118584,I671147,I671138);
and I_6765 (I118601,I118584,I671153);
DFFARX1 I_6766 (I118601,I3563,I118338,I118627,);
DFFARX1 I_6767 (I118627,I3563,I118338,I118644,);
not I_6768 (I118330,I118644);
not I_6769 (I118666,I118627);
nand I_6770 (I118315,I118666,I118505);
nor I_6771 (I118697,I671144,I671138);
not I_6772 (I118714,I118697);
nor I_6773 (I118731,I118666,I118714);
nor I_6774 (I118748,I118372,I118731);
DFFARX1 I_6775 (I118748,I3563,I118338,I118324,);
nor I_6776 (I118779,I118432,I118714);
nor I_6777 (I118312,I118627,I118779);
nor I_6778 (I118321,I118562,I118697);
nor I_6779 (I118309,I118432,I118697);
not I_6780 (I118865,I3570);
DFFARX1 I_6781 (I1265455,I3563,I118865,I118891,);
not I_6782 (I118899,I118891);
nand I_6783 (I118916,I1265449,I1265470);
and I_6784 (I118933,I118916,I1265461);
DFFARX1 I_6785 (I118933,I3563,I118865,I118959,);
DFFARX1 I_6786 (I1265452,I3563,I118865,I118976,);
and I_6787 (I118984,I118976,I1265464);
nor I_6788 (I119001,I118959,I118984);
DFFARX1 I_6789 (I119001,I3563,I118865,I118833,);
nand I_6790 (I119032,I118976,I1265464);
nand I_6791 (I119049,I118899,I119032);
not I_6792 (I118845,I119049);
DFFARX1 I_6793 (I1265452,I3563,I118865,I119089,);
DFFARX1 I_6794 (I119089,I3563,I118865,I118854,);
nand I_6795 (I119111,I1265473,I1265458);
and I_6796 (I119128,I119111,I1265449);
DFFARX1 I_6797 (I119128,I3563,I118865,I119154,);
DFFARX1 I_6798 (I119154,I3563,I118865,I119171,);
not I_6799 (I118857,I119171);
not I_6800 (I119193,I119154);
nand I_6801 (I118842,I119193,I119032);
nor I_6802 (I119224,I1265467,I1265458);
not I_6803 (I119241,I119224);
nor I_6804 (I119258,I119193,I119241);
nor I_6805 (I119275,I118899,I119258);
DFFARX1 I_6806 (I119275,I3563,I118865,I118851,);
nor I_6807 (I119306,I118959,I119241);
nor I_6808 (I118839,I119154,I119306);
nor I_6809 (I118848,I119089,I119224);
nor I_6810 (I118836,I118959,I119224);
not I_6811 (I119392,I3570);
DFFARX1 I_6812 (I822132,I3563,I119392,I119418,);
not I_6813 (I119426,I119418);
nand I_6814 (I119443,I822129,I822144);
and I_6815 (I119460,I119443,I822126);
DFFARX1 I_6816 (I119460,I3563,I119392,I119486,);
DFFARX1 I_6817 (I822123,I3563,I119392,I119503,);
and I_6818 (I119511,I119503,I822123);
nor I_6819 (I119528,I119486,I119511);
DFFARX1 I_6820 (I119528,I3563,I119392,I119360,);
nand I_6821 (I119559,I119503,I822123);
nand I_6822 (I119576,I119426,I119559);
not I_6823 (I119372,I119576);
DFFARX1 I_6824 (I822126,I3563,I119392,I119616,);
DFFARX1 I_6825 (I119616,I3563,I119392,I119381,);
nand I_6826 (I119638,I822138,I822129);
and I_6827 (I119655,I119638,I822141);
DFFARX1 I_6828 (I119655,I3563,I119392,I119681,);
DFFARX1 I_6829 (I119681,I3563,I119392,I119698,);
not I_6830 (I119384,I119698);
not I_6831 (I119720,I119681);
nand I_6832 (I119369,I119720,I119559);
nor I_6833 (I119751,I822135,I822129);
not I_6834 (I119768,I119751);
nor I_6835 (I119785,I119720,I119768);
nor I_6836 (I119802,I119426,I119785);
DFFARX1 I_6837 (I119802,I3563,I119392,I119378,);
nor I_6838 (I119833,I119486,I119768);
nor I_6839 (I119366,I119681,I119833);
nor I_6840 (I119375,I119616,I119751);
nor I_6841 (I119363,I119486,I119751);
not I_6842 (I119919,I3570);
DFFARX1 I_6843 (I510548,I3563,I119919,I119945,);
not I_6844 (I119953,I119945);
nand I_6845 (I119970,I510542,I510533);
and I_6846 (I119987,I119970,I510554);
DFFARX1 I_6847 (I119987,I3563,I119919,I120013,);
DFFARX1 I_6848 (I510536,I3563,I119919,I120030,);
and I_6849 (I120038,I120030,I510530);
nor I_6850 (I120055,I120013,I120038);
DFFARX1 I_6851 (I120055,I3563,I119919,I119887,);
nand I_6852 (I120086,I120030,I510530);
nand I_6853 (I120103,I119953,I120086);
not I_6854 (I119899,I120103);
DFFARX1 I_6855 (I510530,I3563,I119919,I120143,);
DFFARX1 I_6856 (I120143,I3563,I119919,I119908,);
nand I_6857 (I120165,I510557,I510539);
and I_6858 (I120182,I120165,I510545);
DFFARX1 I_6859 (I120182,I3563,I119919,I120208,);
DFFARX1 I_6860 (I120208,I3563,I119919,I120225,);
not I_6861 (I119911,I120225);
not I_6862 (I120247,I120208);
nand I_6863 (I119896,I120247,I120086);
nor I_6864 (I120278,I510551,I510539);
not I_6865 (I120295,I120278);
nor I_6866 (I120312,I120247,I120295);
nor I_6867 (I120329,I119953,I120312);
DFFARX1 I_6868 (I120329,I3563,I119919,I119905,);
nor I_6869 (I120360,I120013,I120295);
nor I_6870 (I119893,I120208,I120360);
nor I_6871 (I119902,I120143,I120278);
nor I_6872 (I119890,I120013,I120278);
not I_6873 (I120446,I3570);
DFFARX1 I_6874 (I377090,I3563,I120446,I120472,);
not I_6875 (I120480,I120472);
nand I_6876 (I120497,I377072,I377087);
and I_6877 (I120514,I120497,I377063);
DFFARX1 I_6878 (I120514,I3563,I120446,I120540,);
DFFARX1 I_6879 (I377066,I3563,I120446,I120557,);
and I_6880 (I120565,I120557,I377081);
nor I_6881 (I120582,I120540,I120565);
DFFARX1 I_6882 (I120582,I3563,I120446,I120414,);
nand I_6883 (I120613,I120557,I377081);
nand I_6884 (I120630,I120480,I120613);
not I_6885 (I120426,I120630);
DFFARX1 I_6886 (I377084,I3563,I120446,I120670,);
DFFARX1 I_6887 (I120670,I3563,I120446,I120435,);
nand I_6888 (I120692,I377063,I377075);
and I_6889 (I120709,I120692,I377069);
DFFARX1 I_6890 (I120709,I3563,I120446,I120735,);
DFFARX1 I_6891 (I120735,I3563,I120446,I120752,);
not I_6892 (I120438,I120752);
not I_6893 (I120774,I120735);
nand I_6894 (I120423,I120774,I120613);
nor I_6895 (I120805,I377078,I377075);
not I_6896 (I120822,I120805);
nor I_6897 (I120839,I120774,I120822);
nor I_6898 (I120856,I120480,I120839);
DFFARX1 I_6899 (I120856,I3563,I120446,I120432,);
nor I_6900 (I120887,I120540,I120822);
nor I_6901 (I120420,I120735,I120887);
nor I_6902 (I120429,I120670,I120805);
nor I_6903 (I120417,I120540,I120805);
not I_6904 (I120973,I3570);
DFFARX1 I_6905 (I725473,I3563,I120973,I120999,);
not I_6906 (I121007,I120999);
nand I_6907 (I121024,I725464,I725482);
and I_6908 (I121041,I121024,I725461);
DFFARX1 I_6909 (I121041,I3563,I120973,I121067,);
DFFARX1 I_6910 (I725464,I3563,I120973,I121084,);
and I_6911 (I121092,I121084,I725467);
nor I_6912 (I121109,I121067,I121092);
DFFARX1 I_6913 (I121109,I3563,I120973,I120941,);
nand I_6914 (I121140,I121084,I725467);
nand I_6915 (I121157,I121007,I121140);
not I_6916 (I120953,I121157);
DFFARX1 I_6917 (I725461,I3563,I120973,I121197,);
DFFARX1 I_6918 (I121197,I3563,I120973,I120962,);
nand I_6919 (I121219,I725479,I725470);
and I_6920 (I121236,I121219,I725485);
DFFARX1 I_6921 (I121236,I3563,I120973,I121262,);
DFFARX1 I_6922 (I121262,I3563,I120973,I121279,);
not I_6923 (I120965,I121279);
not I_6924 (I121301,I121262);
nand I_6925 (I120950,I121301,I121140);
nor I_6926 (I121332,I725476,I725470);
not I_6927 (I121349,I121332);
nor I_6928 (I121366,I121301,I121349);
nor I_6929 (I121383,I121007,I121366);
DFFARX1 I_6930 (I121383,I3563,I120973,I120959,);
nor I_6931 (I121414,I121067,I121349);
nor I_6932 (I120947,I121262,I121414);
nor I_6933 (I120956,I121197,I121332);
nor I_6934 (I120944,I121067,I121332);
not I_6935 (I121500,I3570);
DFFARX1 I_6936 (I783851,I3563,I121500,I121526,);
not I_6937 (I121534,I121526);
nand I_6938 (I121551,I783842,I783860);
and I_6939 (I121568,I121551,I783839);
DFFARX1 I_6940 (I121568,I3563,I121500,I121594,);
DFFARX1 I_6941 (I783842,I3563,I121500,I121611,);
and I_6942 (I121619,I121611,I783845);
nor I_6943 (I121636,I121594,I121619);
DFFARX1 I_6944 (I121636,I3563,I121500,I121468,);
nand I_6945 (I121667,I121611,I783845);
nand I_6946 (I121684,I121534,I121667);
not I_6947 (I121480,I121684);
DFFARX1 I_6948 (I783839,I3563,I121500,I121724,);
DFFARX1 I_6949 (I121724,I3563,I121500,I121489,);
nand I_6950 (I121746,I783857,I783848);
and I_6951 (I121763,I121746,I783863);
DFFARX1 I_6952 (I121763,I3563,I121500,I121789,);
DFFARX1 I_6953 (I121789,I3563,I121500,I121806,);
not I_6954 (I121492,I121806);
not I_6955 (I121828,I121789);
nand I_6956 (I121477,I121828,I121667);
nor I_6957 (I121859,I783854,I783848);
not I_6958 (I121876,I121859);
nor I_6959 (I121893,I121828,I121876);
nor I_6960 (I121910,I121534,I121893);
DFFARX1 I_6961 (I121910,I3563,I121500,I121486,);
nor I_6962 (I121941,I121594,I121876);
nor I_6963 (I121474,I121789,I121941);
nor I_6964 (I121483,I121724,I121859);
nor I_6965 (I121471,I121594,I121859);
not I_6966 (I122027,I3570);
DFFARX1 I_6967 (I430580,I3563,I122027,I122053,);
not I_6968 (I122061,I122053);
nand I_6969 (I122078,I430574,I430565);
and I_6970 (I122095,I122078,I430586);
DFFARX1 I_6971 (I122095,I3563,I122027,I122121,);
DFFARX1 I_6972 (I430568,I3563,I122027,I122138,);
and I_6973 (I122146,I122138,I430562);
nor I_6974 (I122163,I122121,I122146);
DFFARX1 I_6975 (I122163,I3563,I122027,I121995,);
nand I_6976 (I122194,I122138,I430562);
nand I_6977 (I122211,I122061,I122194);
not I_6978 (I122007,I122211);
DFFARX1 I_6979 (I430562,I3563,I122027,I122251,);
DFFARX1 I_6980 (I122251,I3563,I122027,I122016,);
nand I_6981 (I122273,I430589,I430571);
and I_6982 (I122290,I122273,I430577);
DFFARX1 I_6983 (I122290,I3563,I122027,I122316,);
DFFARX1 I_6984 (I122316,I3563,I122027,I122333,);
not I_6985 (I122019,I122333);
not I_6986 (I122355,I122316);
nand I_6987 (I122004,I122355,I122194);
nor I_6988 (I122386,I430583,I430571);
not I_6989 (I122403,I122386);
nor I_6990 (I122420,I122355,I122403);
nor I_6991 (I122437,I122061,I122420);
DFFARX1 I_6992 (I122437,I3563,I122027,I122013,);
nor I_6993 (I122468,I122121,I122403);
nor I_6994 (I122001,I122316,I122468);
nor I_6995 (I122010,I122251,I122386);
nor I_6996 (I121998,I122121,I122386);
not I_6997 (I122554,I3570);
DFFARX1 I_6998 (I957520,I3563,I122554,I122580,);
not I_6999 (I122588,I122580);
nand I_7000 (I122605,I957538,I957532);
and I_7001 (I122622,I122605,I957511);
DFFARX1 I_7002 (I122622,I3563,I122554,I122648,);
DFFARX1 I_7003 (I957529,I3563,I122554,I122665,);
and I_7004 (I122673,I122665,I957514);
nor I_7005 (I122690,I122648,I122673);
DFFARX1 I_7006 (I122690,I3563,I122554,I122522,);
nand I_7007 (I122721,I122665,I957514);
nand I_7008 (I122738,I122588,I122721);
not I_7009 (I122534,I122738);
DFFARX1 I_7010 (I957526,I3563,I122554,I122778,);
DFFARX1 I_7011 (I122778,I3563,I122554,I122543,);
nand I_7012 (I122800,I957535,I957523);
and I_7013 (I122817,I122800,I957517);
DFFARX1 I_7014 (I122817,I3563,I122554,I122843,);
DFFARX1 I_7015 (I122843,I3563,I122554,I122860,);
not I_7016 (I122546,I122860);
not I_7017 (I122882,I122843);
nand I_7018 (I122531,I122882,I122721);
nor I_7019 (I122913,I957511,I957523);
not I_7020 (I122930,I122913);
nor I_7021 (I122947,I122882,I122930);
nor I_7022 (I122964,I122588,I122947);
DFFARX1 I_7023 (I122964,I3563,I122554,I122540,);
nor I_7024 (I122995,I122648,I122930);
nor I_7025 (I122528,I122843,I122995);
nor I_7026 (I122537,I122778,I122913);
nor I_7027 (I122525,I122648,I122913);
not I_7028 (I123081,I3570);
DFFARX1 I_7029 (I1243015,I3563,I123081,I123107,);
not I_7030 (I123115,I123107);
nand I_7031 (I123132,I1243030,I1243009);
and I_7032 (I123149,I123132,I1243012);
DFFARX1 I_7033 (I123149,I3563,I123081,I123175,);
DFFARX1 I_7034 (I1243033,I3563,I123081,I123192,);
and I_7035 (I123200,I123192,I1243012);
nor I_7036 (I123217,I123175,I123200);
DFFARX1 I_7037 (I123217,I3563,I123081,I123049,);
nand I_7038 (I123248,I123192,I1243012);
nand I_7039 (I123265,I123115,I123248);
not I_7040 (I123061,I123265);
DFFARX1 I_7041 (I1243009,I3563,I123081,I123305,);
DFFARX1 I_7042 (I123305,I3563,I123081,I123070,);
nand I_7043 (I123327,I1243021,I1243018);
and I_7044 (I123344,I123327,I1243024);
DFFARX1 I_7045 (I123344,I3563,I123081,I123370,);
DFFARX1 I_7046 (I123370,I3563,I123081,I123387,);
not I_7047 (I123073,I123387);
not I_7048 (I123409,I123370);
nand I_7049 (I123058,I123409,I123248);
nor I_7050 (I123440,I1243027,I1243018);
not I_7051 (I123457,I123440);
nor I_7052 (I123474,I123409,I123457);
nor I_7053 (I123491,I123115,I123474);
DFFARX1 I_7054 (I123491,I3563,I123081,I123067,);
nor I_7055 (I123522,I123175,I123457);
nor I_7056 (I123055,I123370,I123522);
nor I_7057 (I123064,I123305,I123440);
nor I_7058 (I123052,I123175,I123440);
not I_7059 (I123608,I3570);
DFFARX1 I_7060 (I615072,I3563,I123608,I123634,);
not I_7061 (I123642,I123634);
nand I_7062 (I123659,I615084,I615069);
and I_7063 (I123676,I123659,I615063);
DFFARX1 I_7064 (I123676,I3563,I123608,I123702,);
DFFARX1 I_7065 (I615078,I3563,I123608,I123719,);
and I_7066 (I123727,I123719,I615066);
nor I_7067 (I123744,I123702,I123727);
DFFARX1 I_7068 (I123744,I3563,I123608,I123576,);
nand I_7069 (I123775,I123719,I615066);
nand I_7070 (I123792,I123642,I123775);
not I_7071 (I123588,I123792);
DFFARX1 I_7072 (I615075,I3563,I123608,I123832,);
DFFARX1 I_7073 (I123832,I3563,I123608,I123597,);
nand I_7074 (I123854,I615081,I615087);
and I_7075 (I123871,I123854,I615063);
DFFARX1 I_7076 (I123871,I3563,I123608,I123897,);
DFFARX1 I_7077 (I123897,I3563,I123608,I123914,);
not I_7078 (I123600,I123914);
not I_7079 (I123936,I123897);
nand I_7080 (I123585,I123936,I123775);
nor I_7081 (I123967,I615066,I615087);
not I_7082 (I123984,I123967);
nor I_7083 (I124001,I123936,I123984);
nor I_7084 (I124018,I123642,I124001);
DFFARX1 I_7085 (I124018,I3563,I123608,I123594,);
nor I_7086 (I124049,I123702,I123984);
nor I_7087 (I123582,I123897,I124049);
nor I_7088 (I123591,I123832,I123967);
nor I_7089 (I123579,I123702,I123967);
not I_7090 (I124135,I3570);
DFFARX1 I_7091 (I1169609,I3563,I124135,I124161,);
not I_7092 (I124169,I124161);
nand I_7093 (I124186,I1169624,I1169603);
and I_7094 (I124203,I124186,I1169606);
DFFARX1 I_7095 (I124203,I3563,I124135,I124229,);
DFFARX1 I_7096 (I1169627,I3563,I124135,I124246,);
and I_7097 (I124254,I124246,I1169606);
nor I_7098 (I124271,I124229,I124254);
DFFARX1 I_7099 (I124271,I3563,I124135,I124103,);
nand I_7100 (I124302,I124246,I1169606);
nand I_7101 (I124319,I124169,I124302);
not I_7102 (I124115,I124319);
DFFARX1 I_7103 (I1169603,I3563,I124135,I124359,);
DFFARX1 I_7104 (I124359,I3563,I124135,I124124,);
nand I_7105 (I124381,I1169615,I1169612);
and I_7106 (I124398,I124381,I1169618);
DFFARX1 I_7107 (I124398,I3563,I124135,I124424,);
DFFARX1 I_7108 (I124424,I3563,I124135,I124441,);
not I_7109 (I124127,I124441);
not I_7110 (I124463,I124424);
nand I_7111 (I124112,I124463,I124302);
nor I_7112 (I124494,I1169621,I1169612);
not I_7113 (I124511,I124494);
nor I_7114 (I124528,I124463,I124511);
nor I_7115 (I124545,I124169,I124528);
DFFARX1 I_7116 (I124545,I3563,I124135,I124121,);
nor I_7117 (I124576,I124229,I124511);
nor I_7118 (I124109,I124424,I124576);
nor I_7119 (I124118,I124359,I124494);
nor I_7120 (I124106,I124229,I124494);
not I_7121 (I124662,I3570);
DFFARX1 I_7122 (I898547,I3563,I124662,I124688,);
not I_7123 (I124696,I124688);
nand I_7124 (I124713,I898544,I898559);
and I_7125 (I124730,I124713,I898541);
DFFARX1 I_7126 (I124730,I3563,I124662,I124756,);
DFFARX1 I_7127 (I898538,I3563,I124662,I124773,);
and I_7128 (I124781,I124773,I898538);
nor I_7129 (I124798,I124756,I124781);
DFFARX1 I_7130 (I124798,I3563,I124662,I124630,);
nand I_7131 (I124829,I124773,I898538);
nand I_7132 (I124846,I124696,I124829);
not I_7133 (I124642,I124846);
DFFARX1 I_7134 (I898541,I3563,I124662,I124886,);
DFFARX1 I_7135 (I124886,I3563,I124662,I124651,);
nand I_7136 (I124908,I898553,I898544);
and I_7137 (I124925,I124908,I898556);
DFFARX1 I_7138 (I124925,I3563,I124662,I124951,);
DFFARX1 I_7139 (I124951,I3563,I124662,I124968,);
not I_7140 (I124654,I124968);
not I_7141 (I124990,I124951);
nand I_7142 (I124639,I124990,I124829);
nor I_7143 (I125021,I898550,I898544);
not I_7144 (I125038,I125021);
nor I_7145 (I125055,I124990,I125038);
nor I_7146 (I125072,I124696,I125055);
DFFARX1 I_7147 (I125072,I3563,I124662,I124648,);
nor I_7148 (I125103,I124756,I125038);
nor I_7149 (I124636,I124951,I125103);
nor I_7150 (I124645,I124886,I125021);
nor I_7151 (I124633,I124756,I125021);
not I_7152 (I125189,I3570);
DFFARX1 I_7153 (I44550,I3563,I125189,I125215,);
not I_7154 (I125223,I125215);
nand I_7155 (I125240,I44538,I44544);
and I_7156 (I125257,I125240,I44547);
DFFARX1 I_7157 (I125257,I3563,I125189,I125283,);
DFFARX1 I_7158 (I44529,I3563,I125189,I125300,);
and I_7159 (I125308,I125300,I44535);
nor I_7160 (I125325,I125283,I125308);
DFFARX1 I_7161 (I125325,I3563,I125189,I125157,);
nand I_7162 (I125356,I125300,I44535);
nand I_7163 (I125373,I125223,I125356);
not I_7164 (I125169,I125373);
DFFARX1 I_7165 (I44529,I3563,I125189,I125413,);
DFFARX1 I_7166 (I125413,I3563,I125189,I125178,);
nand I_7167 (I125435,I44532,I44526);
and I_7168 (I125452,I125435,I44541);
DFFARX1 I_7169 (I125452,I3563,I125189,I125478,);
DFFARX1 I_7170 (I125478,I3563,I125189,I125495,);
not I_7171 (I125181,I125495);
not I_7172 (I125517,I125478);
nand I_7173 (I125166,I125517,I125356);
nor I_7174 (I125548,I44526,I44526);
not I_7175 (I125565,I125548);
nor I_7176 (I125582,I125517,I125565);
nor I_7177 (I125599,I125223,I125582);
DFFARX1 I_7178 (I125599,I3563,I125189,I125175,);
nor I_7179 (I125630,I125283,I125565);
nor I_7180 (I125163,I125478,I125630);
nor I_7181 (I125172,I125413,I125548);
nor I_7182 (I125160,I125283,I125548);
not I_7183 (I125716,I3570);
DFFARX1 I_7184 (I639926,I3563,I125716,I125742,);
not I_7185 (I125750,I125742);
nand I_7186 (I125767,I639938,I639923);
and I_7187 (I125784,I125767,I639917);
DFFARX1 I_7188 (I125784,I3563,I125716,I125810,);
DFFARX1 I_7189 (I639932,I3563,I125716,I125827,);
and I_7190 (I125835,I125827,I639920);
nor I_7191 (I125852,I125810,I125835);
DFFARX1 I_7192 (I125852,I3563,I125716,I125684,);
nand I_7193 (I125883,I125827,I639920);
nand I_7194 (I125900,I125750,I125883);
not I_7195 (I125696,I125900);
DFFARX1 I_7196 (I639929,I3563,I125716,I125940,);
DFFARX1 I_7197 (I125940,I3563,I125716,I125705,);
nand I_7198 (I125962,I639935,I639941);
and I_7199 (I125979,I125962,I639917);
DFFARX1 I_7200 (I125979,I3563,I125716,I126005,);
DFFARX1 I_7201 (I126005,I3563,I125716,I126022,);
not I_7202 (I125708,I126022);
not I_7203 (I126044,I126005);
nand I_7204 (I125693,I126044,I125883);
nor I_7205 (I126075,I639920,I639941);
not I_7206 (I126092,I126075);
nor I_7207 (I126109,I126044,I126092);
nor I_7208 (I126126,I125750,I126109);
DFFARX1 I_7209 (I126126,I3563,I125716,I125702,);
nor I_7210 (I126157,I125810,I126092);
nor I_7211 (I125690,I126005,I126157);
nor I_7212 (I125699,I125940,I126075);
nor I_7213 (I125687,I125810,I126075);
not I_7214 (I126243,I3570);
DFFARX1 I_7215 (I823186,I3563,I126243,I126269,);
not I_7216 (I126277,I126269);
nand I_7217 (I126294,I823183,I823198);
and I_7218 (I126311,I126294,I823180);
DFFARX1 I_7219 (I126311,I3563,I126243,I126337,);
DFFARX1 I_7220 (I823177,I3563,I126243,I126354,);
and I_7221 (I126362,I126354,I823177);
nor I_7222 (I126379,I126337,I126362);
DFFARX1 I_7223 (I126379,I3563,I126243,I126211,);
nand I_7224 (I126410,I126354,I823177);
nand I_7225 (I126427,I126277,I126410);
not I_7226 (I126223,I126427);
DFFARX1 I_7227 (I823180,I3563,I126243,I126467,);
DFFARX1 I_7228 (I126467,I3563,I126243,I126232,);
nand I_7229 (I126489,I823192,I823183);
and I_7230 (I126506,I126489,I823195);
DFFARX1 I_7231 (I126506,I3563,I126243,I126532,);
DFFARX1 I_7232 (I126532,I3563,I126243,I126549,);
not I_7233 (I126235,I126549);
not I_7234 (I126571,I126532);
nand I_7235 (I126220,I126571,I126410);
nor I_7236 (I126602,I823189,I823183);
not I_7237 (I126619,I126602);
nor I_7238 (I126636,I126571,I126619);
nor I_7239 (I126653,I126277,I126636);
DFFARX1 I_7240 (I126653,I3563,I126243,I126229,);
nor I_7241 (I126684,I126337,I126619);
nor I_7242 (I126217,I126532,I126684);
nor I_7243 (I126226,I126467,I126602);
nor I_7244 (I126214,I126337,I126602);
not I_7245 (I126770,I3570);
DFFARX1 I_7246 (I483892,I3563,I126770,I126796,);
not I_7247 (I126804,I126796);
nand I_7248 (I126821,I483886,I483877);
and I_7249 (I126838,I126821,I483898);
DFFARX1 I_7250 (I126838,I3563,I126770,I126864,);
DFFARX1 I_7251 (I483880,I3563,I126770,I126881,);
and I_7252 (I126889,I126881,I483874);
nor I_7253 (I126906,I126864,I126889);
DFFARX1 I_7254 (I126906,I3563,I126770,I126738,);
nand I_7255 (I126937,I126881,I483874);
nand I_7256 (I126954,I126804,I126937);
not I_7257 (I126750,I126954);
DFFARX1 I_7258 (I483874,I3563,I126770,I126994,);
DFFARX1 I_7259 (I126994,I3563,I126770,I126759,);
nand I_7260 (I127016,I483901,I483883);
and I_7261 (I127033,I127016,I483889);
DFFARX1 I_7262 (I127033,I3563,I126770,I127059,);
DFFARX1 I_7263 (I127059,I3563,I126770,I127076,);
not I_7264 (I126762,I127076);
not I_7265 (I127098,I127059);
nand I_7266 (I126747,I127098,I126937);
nor I_7267 (I127129,I483895,I483883);
not I_7268 (I127146,I127129);
nor I_7269 (I127163,I127098,I127146);
nor I_7270 (I127180,I126804,I127163);
DFFARX1 I_7271 (I127180,I3563,I126770,I126756,);
nor I_7272 (I127211,I126864,I127146);
nor I_7273 (I126744,I127059,I127211);
nor I_7274 (I126753,I126994,I127129);
nor I_7275 (I126741,I126864,I127129);
not I_7276 (I127297,I3570);
DFFARX1 I_7277 (I1133195,I3563,I127297,I127323,);
not I_7278 (I127331,I127323);
nand I_7279 (I127348,I1133210,I1133189);
and I_7280 (I127365,I127348,I1133192);
DFFARX1 I_7281 (I127365,I3563,I127297,I127391,);
DFFARX1 I_7282 (I1133213,I3563,I127297,I127408,);
and I_7283 (I127416,I127408,I1133192);
nor I_7284 (I127433,I127391,I127416);
DFFARX1 I_7285 (I127433,I3563,I127297,I127265,);
nand I_7286 (I127464,I127408,I1133192);
nand I_7287 (I127481,I127331,I127464);
not I_7288 (I127277,I127481);
DFFARX1 I_7289 (I1133189,I3563,I127297,I127521,);
DFFARX1 I_7290 (I127521,I3563,I127297,I127286,);
nand I_7291 (I127543,I1133201,I1133198);
and I_7292 (I127560,I127543,I1133204);
DFFARX1 I_7293 (I127560,I3563,I127297,I127586,);
DFFARX1 I_7294 (I127586,I3563,I127297,I127603,);
not I_7295 (I127289,I127603);
not I_7296 (I127625,I127586);
nand I_7297 (I127274,I127625,I127464);
nor I_7298 (I127656,I1133207,I1133198);
not I_7299 (I127673,I127656);
nor I_7300 (I127690,I127625,I127673);
nor I_7301 (I127707,I127331,I127690);
DFFARX1 I_7302 (I127707,I3563,I127297,I127283,);
nor I_7303 (I127738,I127391,I127673);
nor I_7304 (I127271,I127586,I127738);
nor I_7305 (I127280,I127521,I127656);
nor I_7306 (I127268,I127391,I127656);
not I_7307 (I127824,I3570);
DFFARX1 I_7308 (I1024704,I3563,I127824,I127850,);
not I_7309 (I127858,I127850);
nand I_7310 (I127875,I1024722,I1024716);
and I_7311 (I127892,I127875,I1024695);
DFFARX1 I_7312 (I127892,I3563,I127824,I127918,);
DFFARX1 I_7313 (I1024713,I3563,I127824,I127935,);
and I_7314 (I127943,I127935,I1024698);
nor I_7315 (I127960,I127918,I127943);
DFFARX1 I_7316 (I127960,I3563,I127824,I127792,);
nand I_7317 (I127991,I127935,I1024698);
nand I_7318 (I128008,I127858,I127991);
not I_7319 (I127804,I128008);
DFFARX1 I_7320 (I1024710,I3563,I127824,I128048,);
DFFARX1 I_7321 (I128048,I3563,I127824,I127813,);
nand I_7322 (I128070,I1024719,I1024707);
and I_7323 (I128087,I128070,I1024701);
DFFARX1 I_7324 (I128087,I3563,I127824,I128113,);
DFFARX1 I_7325 (I128113,I3563,I127824,I128130,);
not I_7326 (I127816,I128130);
not I_7327 (I128152,I128113);
nand I_7328 (I127801,I128152,I127991);
nor I_7329 (I128183,I1024695,I1024707);
not I_7330 (I128200,I128183);
nor I_7331 (I128217,I128152,I128200);
nor I_7332 (I128234,I127858,I128217);
DFFARX1 I_7333 (I128234,I3563,I127824,I127810,);
nor I_7334 (I128265,I127918,I128200);
nor I_7335 (I127798,I128113,I128265);
nor I_7336 (I127807,I128048,I128183);
nor I_7337 (I127795,I127918,I128183);
not I_7338 (I128351,I3570);
DFFARX1 I_7339 (I608714,I3563,I128351,I128377,);
not I_7340 (I128385,I128377);
nand I_7341 (I128402,I608726,I608711);
and I_7342 (I128419,I128402,I608705);
DFFARX1 I_7343 (I128419,I3563,I128351,I128445,);
DFFARX1 I_7344 (I608720,I3563,I128351,I128462,);
and I_7345 (I128470,I128462,I608708);
nor I_7346 (I128487,I128445,I128470);
DFFARX1 I_7347 (I128487,I3563,I128351,I128319,);
nand I_7348 (I128518,I128462,I608708);
nand I_7349 (I128535,I128385,I128518);
not I_7350 (I128331,I128535);
DFFARX1 I_7351 (I608717,I3563,I128351,I128575,);
DFFARX1 I_7352 (I128575,I3563,I128351,I128340,);
nand I_7353 (I128597,I608723,I608729);
and I_7354 (I128614,I128597,I608705);
DFFARX1 I_7355 (I128614,I3563,I128351,I128640,);
DFFARX1 I_7356 (I128640,I3563,I128351,I128657,);
not I_7357 (I128343,I128657);
not I_7358 (I128679,I128640);
nand I_7359 (I128328,I128679,I128518);
nor I_7360 (I128710,I608708,I608729);
not I_7361 (I128727,I128710);
nor I_7362 (I128744,I128679,I128727);
nor I_7363 (I128761,I128385,I128744);
DFFARX1 I_7364 (I128761,I3563,I128351,I128337,);
nor I_7365 (I128792,I128445,I128727);
nor I_7366 (I128325,I128640,I128792);
nor I_7367 (I128334,I128575,I128710);
nor I_7368 (I128322,I128445,I128710);
not I_7369 (I128878,I3570);
DFFARX1 I_7370 (I360753,I3563,I128878,I128904,);
not I_7371 (I128912,I128904);
nand I_7372 (I128929,I360735,I360750);
and I_7373 (I128946,I128929,I360726);
DFFARX1 I_7374 (I128946,I3563,I128878,I128972,);
DFFARX1 I_7375 (I360729,I3563,I128878,I128989,);
and I_7376 (I128997,I128989,I360744);
nor I_7377 (I129014,I128972,I128997);
DFFARX1 I_7378 (I129014,I3563,I128878,I128846,);
nand I_7379 (I129045,I128989,I360744);
nand I_7380 (I129062,I128912,I129045);
not I_7381 (I128858,I129062);
DFFARX1 I_7382 (I360747,I3563,I128878,I129102,);
DFFARX1 I_7383 (I129102,I3563,I128878,I128867,);
nand I_7384 (I129124,I360726,I360738);
and I_7385 (I129141,I129124,I360732);
DFFARX1 I_7386 (I129141,I3563,I128878,I129167,);
DFFARX1 I_7387 (I129167,I3563,I128878,I129184,);
not I_7388 (I128870,I129184);
not I_7389 (I129206,I129167);
nand I_7390 (I128855,I129206,I129045);
nor I_7391 (I129237,I360741,I360738);
not I_7392 (I129254,I129237);
nor I_7393 (I129271,I129206,I129254);
nor I_7394 (I129288,I128912,I129271);
DFFARX1 I_7395 (I129288,I3563,I128878,I128864,);
nor I_7396 (I129319,I128972,I129254);
nor I_7397 (I128852,I129167,I129319);
nor I_7398 (I128861,I129102,I129237);
nor I_7399 (I128849,I128972,I129237);
not I_7400 (I129405,I3570);
DFFARX1 I_7401 (I635302,I3563,I129405,I129431,);
not I_7402 (I129439,I129431);
nand I_7403 (I129456,I635314,I635299);
and I_7404 (I129473,I129456,I635293);
DFFARX1 I_7405 (I129473,I3563,I129405,I129499,);
DFFARX1 I_7406 (I635308,I3563,I129405,I129516,);
and I_7407 (I129524,I129516,I635296);
nor I_7408 (I129541,I129499,I129524);
DFFARX1 I_7409 (I129541,I3563,I129405,I129373,);
nand I_7410 (I129572,I129516,I635296);
nand I_7411 (I129589,I129439,I129572);
not I_7412 (I129385,I129589);
DFFARX1 I_7413 (I635305,I3563,I129405,I129629,);
DFFARX1 I_7414 (I129629,I3563,I129405,I129394,);
nand I_7415 (I129651,I635311,I635317);
and I_7416 (I129668,I129651,I635293);
DFFARX1 I_7417 (I129668,I3563,I129405,I129694,);
DFFARX1 I_7418 (I129694,I3563,I129405,I129711,);
not I_7419 (I129397,I129711);
not I_7420 (I129733,I129694);
nand I_7421 (I129382,I129733,I129572);
nor I_7422 (I129764,I635296,I635317);
not I_7423 (I129781,I129764);
nor I_7424 (I129798,I129733,I129781);
nor I_7425 (I129815,I129439,I129798);
DFFARX1 I_7426 (I129815,I3563,I129405,I129391,);
nor I_7427 (I129846,I129499,I129781);
nor I_7428 (I129379,I129694,I129846);
nor I_7429 (I129388,I129629,I129764);
nor I_7430 (I129376,I129499,I129764);
not I_7431 (I129932,I3570);
DFFARX1 I_7432 (I974316,I3563,I129932,I129958,);
not I_7433 (I129966,I129958);
nand I_7434 (I129983,I974334,I974328);
and I_7435 (I130000,I129983,I974307);
DFFARX1 I_7436 (I130000,I3563,I129932,I130026,);
DFFARX1 I_7437 (I974325,I3563,I129932,I130043,);
and I_7438 (I130051,I130043,I974310);
nor I_7439 (I130068,I130026,I130051);
DFFARX1 I_7440 (I130068,I3563,I129932,I129900,);
nand I_7441 (I130099,I130043,I974310);
nand I_7442 (I130116,I129966,I130099);
not I_7443 (I129912,I130116);
DFFARX1 I_7444 (I974322,I3563,I129932,I130156,);
DFFARX1 I_7445 (I130156,I3563,I129932,I129921,);
nand I_7446 (I130178,I974331,I974319);
and I_7447 (I130195,I130178,I974313);
DFFARX1 I_7448 (I130195,I3563,I129932,I130221,);
DFFARX1 I_7449 (I130221,I3563,I129932,I130238,);
not I_7450 (I129924,I130238);
not I_7451 (I130260,I130221);
nand I_7452 (I129909,I130260,I130099);
nor I_7453 (I130291,I974307,I974319);
not I_7454 (I130308,I130291);
nor I_7455 (I130325,I130260,I130308);
nor I_7456 (I130342,I129966,I130325);
DFFARX1 I_7457 (I130342,I3563,I129932,I129918,);
nor I_7458 (I130373,I130026,I130308);
nor I_7459 (I129906,I130221,I130373);
nor I_7460 (I129915,I130156,I130291);
nor I_7461 (I129903,I130026,I130291);
not I_7462 (I130459,I3570);
DFFARX1 I_7463 (I953644,I3563,I130459,I130485,);
not I_7464 (I130493,I130485);
nand I_7465 (I130510,I953662,I953656);
and I_7466 (I130527,I130510,I953635);
DFFARX1 I_7467 (I130527,I3563,I130459,I130553,);
DFFARX1 I_7468 (I953653,I3563,I130459,I130570,);
and I_7469 (I130578,I130570,I953638);
nor I_7470 (I130595,I130553,I130578);
DFFARX1 I_7471 (I130595,I3563,I130459,I130427,);
nand I_7472 (I130626,I130570,I953638);
nand I_7473 (I130643,I130493,I130626);
not I_7474 (I130439,I130643);
DFFARX1 I_7475 (I953650,I3563,I130459,I130683,);
DFFARX1 I_7476 (I130683,I3563,I130459,I130448,);
nand I_7477 (I130705,I953659,I953647);
and I_7478 (I130722,I130705,I953641);
DFFARX1 I_7479 (I130722,I3563,I130459,I130748,);
DFFARX1 I_7480 (I130748,I3563,I130459,I130765,);
not I_7481 (I130451,I130765);
not I_7482 (I130787,I130748);
nand I_7483 (I130436,I130787,I130626);
nor I_7484 (I130818,I953635,I953647);
not I_7485 (I130835,I130818);
nor I_7486 (I130852,I130787,I130835);
nor I_7487 (I130869,I130493,I130852);
DFFARX1 I_7488 (I130869,I3563,I130459,I130445,);
nor I_7489 (I130900,I130553,I130835);
nor I_7490 (I130433,I130748,I130900);
nor I_7491 (I130442,I130683,I130818);
nor I_7492 (I130430,I130553,I130818);
not I_7493 (I130986,I3570);
DFFARX1 I_7494 (I46131,I3563,I130986,I131012,);
not I_7495 (I131020,I131012);
nand I_7496 (I131037,I46119,I46125);
and I_7497 (I131054,I131037,I46128);
DFFARX1 I_7498 (I131054,I3563,I130986,I131080,);
DFFARX1 I_7499 (I46110,I3563,I130986,I131097,);
and I_7500 (I131105,I131097,I46116);
nor I_7501 (I131122,I131080,I131105);
DFFARX1 I_7502 (I131122,I3563,I130986,I130954,);
nand I_7503 (I131153,I131097,I46116);
nand I_7504 (I131170,I131020,I131153);
not I_7505 (I130966,I131170);
DFFARX1 I_7506 (I46110,I3563,I130986,I131210,);
DFFARX1 I_7507 (I131210,I3563,I130986,I130975,);
nand I_7508 (I131232,I46113,I46107);
and I_7509 (I131249,I131232,I46122);
DFFARX1 I_7510 (I131249,I3563,I130986,I131275,);
DFFARX1 I_7511 (I131275,I3563,I130986,I131292,);
not I_7512 (I130978,I131292);
not I_7513 (I131314,I131275);
nand I_7514 (I130963,I131314,I131153);
nor I_7515 (I131345,I46107,I46107);
not I_7516 (I131362,I131345);
nor I_7517 (I131379,I131314,I131362);
nor I_7518 (I131396,I131020,I131379);
DFFARX1 I_7519 (I131396,I3563,I130986,I130972,);
nor I_7520 (I131427,I131080,I131362);
nor I_7521 (I130960,I131275,I131427);
nor I_7522 (I130969,I131210,I131345);
nor I_7523 (I130957,I131080,I131345);
not I_7524 (I131513,I3570);
DFFARX1 I_7525 (I1003386,I3563,I131513,I131539,);
not I_7526 (I131547,I131539);
nand I_7527 (I131564,I1003404,I1003398);
and I_7528 (I131581,I131564,I1003377);
DFFARX1 I_7529 (I131581,I3563,I131513,I131607,);
DFFARX1 I_7530 (I1003395,I3563,I131513,I131624,);
and I_7531 (I131632,I131624,I1003380);
nor I_7532 (I131649,I131607,I131632);
DFFARX1 I_7533 (I131649,I3563,I131513,I131481,);
nand I_7534 (I131680,I131624,I1003380);
nand I_7535 (I131697,I131547,I131680);
not I_7536 (I131493,I131697);
DFFARX1 I_7537 (I1003392,I3563,I131513,I131737,);
DFFARX1 I_7538 (I131737,I3563,I131513,I131502,);
nand I_7539 (I131759,I1003401,I1003389);
and I_7540 (I131776,I131759,I1003383);
DFFARX1 I_7541 (I131776,I3563,I131513,I131802,);
DFFARX1 I_7542 (I131802,I3563,I131513,I131819,);
not I_7543 (I131505,I131819);
not I_7544 (I131841,I131802);
nand I_7545 (I131490,I131841,I131680);
nor I_7546 (I131872,I1003377,I1003389);
not I_7547 (I131889,I131872);
nor I_7548 (I131906,I131841,I131889);
nor I_7549 (I131923,I131547,I131906);
DFFARX1 I_7550 (I131923,I3563,I131513,I131499,);
nor I_7551 (I131954,I131607,I131889);
nor I_7552 (I131487,I131802,I131954);
nor I_7553 (I131496,I131737,I131872);
nor I_7554 (I131484,I131607,I131872);
not I_7555 (I132040,I3570);
DFFARX1 I_7556 (I854806,I3563,I132040,I132066,);
not I_7557 (I132074,I132066);
nand I_7558 (I132091,I854803,I854818);
and I_7559 (I132108,I132091,I854800);
DFFARX1 I_7560 (I132108,I3563,I132040,I132134,);
DFFARX1 I_7561 (I854797,I3563,I132040,I132151,);
and I_7562 (I132159,I132151,I854797);
nor I_7563 (I132176,I132134,I132159);
DFFARX1 I_7564 (I132176,I3563,I132040,I132008,);
nand I_7565 (I132207,I132151,I854797);
nand I_7566 (I132224,I132074,I132207);
not I_7567 (I132020,I132224);
DFFARX1 I_7568 (I854800,I3563,I132040,I132264,);
DFFARX1 I_7569 (I132264,I3563,I132040,I132029,);
nand I_7570 (I132286,I854812,I854803);
and I_7571 (I132303,I132286,I854815);
DFFARX1 I_7572 (I132303,I3563,I132040,I132329,);
DFFARX1 I_7573 (I132329,I3563,I132040,I132346,);
not I_7574 (I132032,I132346);
not I_7575 (I132368,I132329);
nand I_7576 (I132017,I132368,I132207);
nor I_7577 (I132399,I854809,I854803);
not I_7578 (I132416,I132399);
nor I_7579 (I132433,I132368,I132416);
nor I_7580 (I132450,I132074,I132433);
DFFARX1 I_7581 (I132450,I3563,I132040,I132026,);
nor I_7582 (I132481,I132134,I132416);
nor I_7583 (I132014,I132329,I132481);
nor I_7584 (I132023,I132264,I132399);
nor I_7585 (I132011,I132134,I132399);
not I_7586 (I132567,I3570);
DFFARX1 I_7587 (I613916,I3563,I132567,I132593,);
not I_7588 (I132601,I132593);
nand I_7589 (I132618,I613928,I613913);
and I_7590 (I132635,I132618,I613907);
DFFARX1 I_7591 (I132635,I3563,I132567,I132661,);
DFFARX1 I_7592 (I613922,I3563,I132567,I132678,);
and I_7593 (I132686,I132678,I613910);
nor I_7594 (I132703,I132661,I132686);
DFFARX1 I_7595 (I132703,I3563,I132567,I132535,);
nand I_7596 (I132734,I132678,I613910);
nand I_7597 (I132751,I132601,I132734);
not I_7598 (I132547,I132751);
DFFARX1 I_7599 (I613919,I3563,I132567,I132791,);
DFFARX1 I_7600 (I132791,I3563,I132567,I132556,);
nand I_7601 (I132813,I613925,I613931);
and I_7602 (I132830,I132813,I613907);
DFFARX1 I_7603 (I132830,I3563,I132567,I132856,);
DFFARX1 I_7604 (I132856,I3563,I132567,I132873,);
not I_7605 (I132559,I132873);
not I_7606 (I132895,I132856);
nand I_7607 (I132544,I132895,I132734);
nor I_7608 (I132926,I613910,I613931);
not I_7609 (I132943,I132926);
nor I_7610 (I132960,I132895,I132943);
nor I_7611 (I132977,I132601,I132960);
DFFARX1 I_7612 (I132977,I3563,I132567,I132553,);
nor I_7613 (I133008,I132661,I132943);
nor I_7614 (I132541,I132856,I133008);
nor I_7615 (I132550,I132791,I132926);
nor I_7616 (I132538,I132661,I132926);
not I_7617 (I133094,I3570);
DFFARX1 I_7618 (I867981,I3563,I133094,I133120,);
not I_7619 (I133128,I133120);
nand I_7620 (I133145,I867978,I867993);
and I_7621 (I133162,I133145,I867975);
DFFARX1 I_7622 (I133162,I3563,I133094,I133188,);
DFFARX1 I_7623 (I867972,I3563,I133094,I133205,);
and I_7624 (I133213,I133205,I867972);
nor I_7625 (I133230,I133188,I133213);
DFFARX1 I_7626 (I133230,I3563,I133094,I133062,);
nand I_7627 (I133261,I133205,I867972);
nand I_7628 (I133278,I133128,I133261);
not I_7629 (I133074,I133278);
DFFARX1 I_7630 (I867975,I3563,I133094,I133318,);
DFFARX1 I_7631 (I133318,I3563,I133094,I133083,);
nand I_7632 (I133340,I867987,I867978);
and I_7633 (I133357,I133340,I867990);
DFFARX1 I_7634 (I133357,I3563,I133094,I133383,);
DFFARX1 I_7635 (I133383,I3563,I133094,I133400,);
not I_7636 (I133086,I133400);
not I_7637 (I133422,I133383);
nand I_7638 (I133071,I133422,I133261);
nor I_7639 (I133453,I867984,I867978);
not I_7640 (I133470,I133453);
nor I_7641 (I133487,I133422,I133470);
nor I_7642 (I133504,I133128,I133487);
DFFARX1 I_7643 (I133504,I3563,I133094,I133080,);
nor I_7644 (I133535,I133188,I133470);
nor I_7645 (I133068,I133383,I133535);
nor I_7646 (I133077,I133318,I133453);
nor I_7647 (I133065,I133188,I133453);
not I_7648 (I133621,I3570);
DFFARX1 I_7649 (I311742,I3563,I133621,I133647,);
not I_7650 (I133655,I133647);
nand I_7651 (I133672,I311724,I311739);
and I_7652 (I133689,I133672,I311715);
DFFARX1 I_7653 (I133689,I3563,I133621,I133715,);
DFFARX1 I_7654 (I311718,I3563,I133621,I133732,);
and I_7655 (I133740,I133732,I311733);
nor I_7656 (I133757,I133715,I133740);
DFFARX1 I_7657 (I133757,I3563,I133621,I133589,);
nand I_7658 (I133788,I133732,I311733);
nand I_7659 (I133805,I133655,I133788);
not I_7660 (I133601,I133805);
DFFARX1 I_7661 (I311736,I3563,I133621,I133845,);
DFFARX1 I_7662 (I133845,I3563,I133621,I133610,);
nand I_7663 (I133867,I311715,I311727);
and I_7664 (I133884,I133867,I311721);
DFFARX1 I_7665 (I133884,I3563,I133621,I133910,);
DFFARX1 I_7666 (I133910,I3563,I133621,I133927,);
not I_7667 (I133613,I133927);
not I_7668 (I133949,I133910);
nand I_7669 (I133598,I133949,I133788);
nor I_7670 (I133980,I311730,I311727);
not I_7671 (I133997,I133980);
nor I_7672 (I134014,I133949,I133997);
nor I_7673 (I134031,I133655,I134014);
DFFARX1 I_7674 (I134031,I3563,I133621,I133607,);
nor I_7675 (I134062,I133715,I133997);
nor I_7676 (I133595,I133910,I134062);
nor I_7677 (I133604,I133845,I133980);
nor I_7678 (I133592,I133715,I133980);
not I_7679 (I134148,I3570);
DFFARX1 I_7680 (I682123,I3563,I134148,I134174,);
not I_7681 (I134182,I134174);
nand I_7682 (I134199,I682114,I682132);
and I_7683 (I134216,I134199,I682111);
DFFARX1 I_7684 (I134216,I3563,I134148,I134242,);
DFFARX1 I_7685 (I682114,I3563,I134148,I134259,);
and I_7686 (I134267,I134259,I682117);
nor I_7687 (I134284,I134242,I134267);
DFFARX1 I_7688 (I134284,I3563,I134148,I134116,);
nand I_7689 (I134315,I134259,I682117);
nand I_7690 (I134332,I134182,I134315);
not I_7691 (I134128,I134332);
DFFARX1 I_7692 (I682111,I3563,I134148,I134372,);
DFFARX1 I_7693 (I134372,I3563,I134148,I134137,);
nand I_7694 (I134394,I682129,I682120);
and I_7695 (I134411,I134394,I682135);
DFFARX1 I_7696 (I134411,I3563,I134148,I134437,);
DFFARX1 I_7697 (I134437,I3563,I134148,I134454,);
not I_7698 (I134140,I134454);
not I_7699 (I134476,I134437);
nand I_7700 (I134125,I134476,I134315);
nor I_7701 (I134507,I682126,I682120);
not I_7702 (I134524,I134507);
nor I_7703 (I134541,I134476,I134524);
nor I_7704 (I134558,I134182,I134541);
DFFARX1 I_7705 (I134558,I3563,I134148,I134134,);
nor I_7706 (I134589,I134242,I134524);
nor I_7707 (I134122,I134437,I134589);
nor I_7708 (I134131,I134372,I134507);
nor I_7709 (I134119,I134242,I134507);
not I_7710 (I134675,I3570);
DFFARX1 I_7711 (I1395205,I3563,I134675,I134701,);
not I_7712 (I134709,I134701);
nand I_7713 (I134726,I1395199,I1395220);
and I_7714 (I134743,I134726,I1395196);
DFFARX1 I_7715 (I134743,I3563,I134675,I134769,);
DFFARX1 I_7716 (I1395217,I3563,I134675,I134786,);
and I_7717 (I134794,I134786,I1395214);
nor I_7718 (I134811,I134769,I134794);
DFFARX1 I_7719 (I134811,I3563,I134675,I134643,);
nand I_7720 (I134842,I134786,I1395214);
nand I_7721 (I134859,I134709,I134842);
not I_7722 (I134655,I134859);
DFFARX1 I_7723 (I1395202,I3563,I134675,I134899,);
DFFARX1 I_7724 (I134899,I3563,I134675,I134664,);
nand I_7725 (I134921,I1395211,I1395208);
and I_7726 (I134938,I134921,I1395193);
DFFARX1 I_7727 (I134938,I3563,I134675,I134964,);
DFFARX1 I_7728 (I134964,I3563,I134675,I134981,);
not I_7729 (I134667,I134981);
not I_7730 (I135003,I134964);
nand I_7731 (I134652,I135003,I134842);
nor I_7732 (I135034,I1395193,I1395208);
not I_7733 (I135051,I135034);
nor I_7734 (I135068,I135003,I135051);
nor I_7735 (I135085,I134709,I135068);
DFFARX1 I_7736 (I135085,I3563,I134675,I134661,);
nor I_7737 (I135116,I134769,I135051);
nor I_7738 (I134649,I134964,I135116);
nor I_7739 (I134658,I134899,I135034);
nor I_7740 (I134646,I134769,I135034);
not I_7741 (I135202,I3570);
DFFARX1 I_7742 (I1129727,I3563,I135202,I135228,);
not I_7743 (I135236,I135228);
nand I_7744 (I135253,I1129742,I1129721);
and I_7745 (I135270,I135253,I1129724);
DFFARX1 I_7746 (I135270,I3563,I135202,I135296,);
DFFARX1 I_7747 (I1129745,I3563,I135202,I135313,);
and I_7748 (I135321,I135313,I1129724);
nor I_7749 (I135338,I135296,I135321);
DFFARX1 I_7750 (I135338,I3563,I135202,I135170,);
nand I_7751 (I135369,I135313,I1129724);
nand I_7752 (I135386,I135236,I135369);
not I_7753 (I135182,I135386);
DFFARX1 I_7754 (I1129721,I3563,I135202,I135426,);
DFFARX1 I_7755 (I135426,I3563,I135202,I135191,);
nand I_7756 (I135448,I1129733,I1129730);
and I_7757 (I135465,I135448,I1129736);
DFFARX1 I_7758 (I135465,I3563,I135202,I135491,);
DFFARX1 I_7759 (I135491,I3563,I135202,I135508,);
not I_7760 (I135194,I135508);
not I_7761 (I135530,I135491);
nand I_7762 (I135179,I135530,I135369);
nor I_7763 (I135561,I1129739,I1129730);
not I_7764 (I135578,I135561);
nor I_7765 (I135595,I135530,I135578);
nor I_7766 (I135612,I135236,I135595);
DFFARX1 I_7767 (I135612,I3563,I135202,I135188,);
nor I_7768 (I135643,I135296,I135578);
nor I_7769 (I135176,I135491,I135643);
nor I_7770 (I135185,I135426,I135561);
nor I_7771 (I135173,I135296,I135561);
not I_7772 (I135729,I3570);
DFFARX1 I_7773 (I308580,I3563,I135729,I135755,);
not I_7774 (I135763,I135755);
nand I_7775 (I135780,I308562,I308577);
and I_7776 (I135797,I135780,I308553);
DFFARX1 I_7777 (I135797,I3563,I135729,I135823,);
DFFARX1 I_7778 (I308556,I3563,I135729,I135840,);
and I_7779 (I135848,I135840,I308571);
nor I_7780 (I135865,I135823,I135848);
DFFARX1 I_7781 (I135865,I3563,I135729,I135697,);
nand I_7782 (I135896,I135840,I308571);
nand I_7783 (I135913,I135763,I135896);
not I_7784 (I135709,I135913);
DFFARX1 I_7785 (I308574,I3563,I135729,I135953,);
DFFARX1 I_7786 (I135953,I3563,I135729,I135718,);
nand I_7787 (I135975,I308553,I308565);
and I_7788 (I135992,I135975,I308559);
DFFARX1 I_7789 (I135992,I3563,I135729,I136018,);
DFFARX1 I_7790 (I136018,I3563,I135729,I136035,);
not I_7791 (I135721,I136035);
not I_7792 (I136057,I136018);
nand I_7793 (I135706,I136057,I135896);
nor I_7794 (I136088,I308568,I308565);
not I_7795 (I136105,I136088);
nor I_7796 (I136122,I136057,I136105);
nor I_7797 (I136139,I135763,I136122);
DFFARX1 I_7798 (I136139,I3563,I135729,I135715,);
nor I_7799 (I136170,I135823,I136105);
nor I_7800 (I135703,I136018,I136170);
nor I_7801 (I135712,I135953,I136088);
nor I_7802 (I135700,I135823,I136088);
not I_7803 (I136256,I3570);
DFFARX1 I_7804 (I1233767,I3563,I136256,I136282,);
not I_7805 (I136290,I136282);
nand I_7806 (I136307,I1233782,I1233761);
and I_7807 (I136324,I136307,I1233764);
DFFARX1 I_7808 (I136324,I3563,I136256,I136350,);
DFFARX1 I_7809 (I1233785,I3563,I136256,I136367,);
and I_7810 (I136375,I136367,I1233764);
nor I_7811 (I136392,I136350,I136375);
DFFARX1 I_7812 (I136392,I3563,I136256,I136224,);
nand I_7813 (I136423,I136367,I1233764);
nand I_7814 (I136440,I136290,I136423);
not I_7815 (I136236,I136440);
DFFARX1 I_7816 (I1233761,I3563,I136256,I136480,);
DFFARX1 I_7817 (I136480,I3563,I136256,I136245,);
nand I_7818 (I136502,I1233773,I1233770);
and I_7819 (I136519,I136502,I1233776);
DFFARX1 I_7820 (I136519,I3563,I136256,I136545,);
DFFARX1 I_7821 (I136545,I3563,I136256,I136562,);
not I_7822 (I136248,I136562);
not I_7823 (I136584,I136545);
nand I_7824 (I136233,I136584,I136423);
nor I_7825 (I136615,I1233779,I1233770);
not I_7826 (I136632,I136615);
nor I_7827 (I136649,I136584,I136632);
nor I_7828 (I136666,I136290,I136649);
DFFARX1 I_7829 (I136666,I3563,I136256,I136242,);
nor I_7830 (I136697,I136350,I136632);
nor I_7831 (I136230,I136545,I136697);
nor I_7832 (I136239,I136480,I136615);
nor I_7833 (I136227,I136350,I136615);
not I_7834 (I136783,I3570);
DFFARX1 I_7835 (I14893,I3563,I136783,I136809,);
not I_7836 (I136817,I136809);
nand I_7837 (I136834,I14878,I14878);
and I_7838 (I136851,I136834,I14899);
DFFARX1 I_7839 (I136851,I3563,I136783,I136877,);
DFFARX1 I_7840 (I14881,I3563,I136783,I136894,);
and I_7841 (I136902,I136894,I14890);
nor I_7842 (I136919,I136877,I136902);
DFFARX1 I_7843 (I136919,I3563,I136783,I136751,);
nand I_7844 (I136950,I136894,I14890);
nand I_7845 (I136967,I136817,I136950);
not I_7846 (I136763,I136967);
DFFARX1 I_7847 (I14884,I3563,I136783,I137007,);
DFFARX1 I_7848 (I137007,I3563,I136783,I136772,);
nand I_7849 (I137029,I14887,I14896);
and I_7850 (I137046,I137029,I14881);
DFFARX1 I_7851 (I137046,I3563,I136783,I137072,);
DFFARX1 I_7852 (I137072,I3563,I136783,I137089,);
not I_7853 (I136775,I137089);
not I_7854 (I137111,I137072);
nand I_7855 (I136760,I137111,I136950);
nor I_7856 (I137142,I14884,I14896);
not I_7857 (I137159,I137142);
nor I_7858 (I137176,I137111,I137159);
nor I_7859 (I137193,I136817,I137176);
DFFARX1 I_7860 (I137193,I3563,I136783,I136769,);
nor I_7861 (I137224,I136877,I137159);
nor I_7862 (I136757,I137072,I137224);
nor I_7863 (I136766,I137007,I137142);
nor I_7864 (I136754,I136877,I137142);
not I_7865 (I137310,I3570);
DFFARX1 I_7866 (I321755,I3563,I137310,I137336,);
not I_7867 (I137344,I137336);
nand I_7868 (I137361,I321737,I321752);
and I_7869 (I137378,I137361,I321728);
DFFARX1 I_7870 (I137378,I3563,I137310,I137404,);
DFFARX1 I_7871 (I321731,I3563,I137310,I137421,);
and I_7872 (I137429,I137421,I321746);
nor I_7873 (I137446,I137404,I137429);
DFFARX1 I_7874 (I137446,I3563,I137310,I137278,);
nand I_7875 (I137477,I137421,I321746);
nand I_7876 (I137494,I137344,I137477);
not I_7877 (I137290,I137494);
DFFARX1 I_7878 (I321749,I3563,I137310,I137534,);
DFFARX1 I_7879 (I137534,I3563,I137310,I137299,);
nand I_7880 (I137556,I321728,I321740);
and I_7881 (I137573,I137556,I321734);
DFFARX1 I_7882 (I137573,I3563,I137310,I137599,);
DFFARX1 I_7883 (I137599,I3563,I137310,I137616,);
not I_7884 (I137302,I137616);
not I_7885 (I137638,I137599);
nand I_7886 (I137287,I137638,I137477);
nor I_7887 (I137669,I321743,I321740);
not I_7888 (I137686,I137669);
nor I_7889 (I137703,I137638,I137686);
nor I_7890 (I137720,I137344,I137703);
DFFARX1 I_7891 (I137720,I3563,I137310,I137296,);
nor I_7892 (I137751,I137404,I137686);
nor I_7893 (I137284,I137599,I137751);
nor I_7894 (I137293,I137534,I137669);
nor I_7895 (I137281,I137404,I137669);
not I_7896 (I137837,I3570);
DFFARX1 I_7897 (I17146,I3563,I137837,I137863,);
not I_7898 (I137871,I137863);
nand I_7899 (I137888,I17134,I17140);
and I_7900 (I137905,I137888,I17143);
DFFARX1 I_7901 (I137905,I3563,I137837,I137931,);
DFFARX1 I_7902 (I17125,I3563,I137837,I137948,);
and I_7903 (I137956,I137948,I17131);
nor I_7904 (I137973,I137931,I137956);
DFFARX1 I_7905 (I137973,I3563,I137837,I137805,);
nand I_7906 (I138004,I137948,I17131);
nand I_7907 (I138021,I137871,I138004);
not I_7908 (I137817,I138021);
DFFARX1 I_7909 (I17125,I3563,I137837,I138061,);
DFFARX1 I_7910 (I138061,I3563,I137837,I137826,);
nand I_7911 (I138083,I17128,I17122);
and I_7912 (I138100,I138083,I17137);
DFFARX1 I_7913 (I138100,I3563,I137837,I138126,);
DFFARX1 I_7914 (I138126,I3563,I137837,I138143,);
not I_7915 (I137829,I138143);
not I_7916 (I138165,I138126);
nand I_7917 (I137814,I138165,I138004);
nor I_7918 (I138196,I17122,I17122);
not I_7919 (I138213,I138196);
nor I_7920 (I138230,I138165,I138213);
nor I_7921 (I138247,I137871,I138230);
DFFARX1 I_7922 (I138247,I3563,I137837,I137823,);
nor I_7923 (I138278,I137931,I138213);
nor I_7924 (I137811,I138126,I138278);
nor I_7925 (I137820,I138061,I138196);
nor I_7926 (I137808,I137931,I138196);
not I_7927 (I138364,I3570);
DFFARX1 I_7928 (I492596,I3563,I138364,I138390,);
not I_7929 (I138398,I138390);
nand I_7930 (I138415,I492590,I492581);
and I_7931 (I138432,I138415,I492602);
DFFARX1 I_7932 (I138432,I3563,I138364,I138458,);
DFFARX1 I_7933 (I492584,I3563,I138364,I138475,);
and I_7934 (I138483,I138475,I492578);
nor I_7935 (I138500,I138458,I138483);
DFFARX1 I_7936 (I138500,I3563,I138364,I138332,);
nand I_7937 (I138531,I138475,I492578);
nand I_7938 (I138548,I138398,I138531);
not I_7939 (I138344,I138548);
DFFARX1 I_7940 (I492578,I3563,I138364,I138588,);
DFFARX1 I_7941 (I138588,I3563,I138364,I138353,);
nand I_7942 (I138610,I492605,I492587);
and I_7943 (I138627,I138610,I492593);
DFFARX1 I_7944 (I138627,I3563,I138364,I138653,);
DFFARX1 I_7945 (I138653,I3563,I138364,I138670,);
not I_7946 (I138356,I138670);
not I_7947 (I138692,I138653);
nand I_7948 (I138341,I138692,I138531);
nor I_7949 (I138723,I492599,I492587);
not I_7950 (I138740,I138723);
nor I_7951 (I138757,I138692,I138740);
nor I_7952 (I138774,I138398,I138757);
DFFARX1 I_7953 (I138774,I3563,I138364,I138350,);
nor I_7954 (I138805,I138458,I138740);
nor I_7955 (I138338,I138653,I138805);
nor I_7956 (I138347,I138588,I138723);
nor I_7957 (I138335,I138458,I138723);
not I_7958 (I138891,I3570);
DFFARX1 I_7959 (I292243,I3563,I138891,I138917,);
not I_7960 (I138925,I138917);
nand I_7961 (I138942,I292225,I292240);
and I_7962 (I138959,I138942,I292216);
DFFARX1 I_7963 (I138959,I3563,I138891,I138985,);
DFFARX1 I_7964 (I292219,I3563,I138891,I139002,);
and I_7965 (I139010,I139002,I292234);
nor I_7966 (I139027,I138985,I139010);
DFFARX1 I_7967 (I139027,I3563,I138891,I138859,);
nand I_7968 (I139058,I139002,I292234);
nand I_7969 (I139075,I138925,I139058);
not I_7970 (I138871,I139075);
DFFARX1 I_7971 (I292237,I3563,I138891,I139115,);
DFFARX1 I_7972 (I139115,I3563,I138891,I138880,);
nand I_7973 (I139137,I292216,I292228);
and I_7974 (I139154,I139137,I292222);
DFFARX1 I_7975 (I139154,I3563,I138891,I139180,);
DFFARX1 I_7976 (I139180,I3563,I138891,I139197,);
not I_7977 (I138883,I139197);
not I_7978 (I139219,I139180);
nand I_7979 (I138868,I139219,I139058);
nor I_7980 (I139250,I292231,I292228);
not I_7981 (I139267,I139250);
nor I_7982 (I139284,I139219,I139267);
nor I_7983 (I139301,I138925,I139284);
DFFARX1 I_7984 (I139301,I3563,I138891,I138877,);
nor I_7985 (I139332,I138985,I139267);
nor I_7986 (I138865,I139180,I139332);
nor I_7987 (I138874,I139115,I139250);
nor I_7988 (I138862,I138985,I139250);
not I_7989 (I139418,I3570);
DFFARX1 I_7990 (I580392,I3563,I139418,I139444,);
not I_7991 (I139452,I139444);
nand I_7992 (I139469,I580404,I580389);
and I_7993 (I139486,I139469,I580383);
DFFARX1 I_7994 (I139486,I3563,I139418,I139512,);
DFFARX1 I_7995 (I580398,I3563,I139418,I139529,);
and I_7996 (I139537,I139529,I580386);
nor I_7997 (I139554,I139512,I139537);
DFFARX1 I_7998 (I139554,I3563,I139418,I139386,);
nand I_7999 (I139585,I139529,I580386);
nand I_8000 (I139602,I139452,I139585);
not I_8001 (I139398,I139602);
DFFARX1 I_8002 (I580395,I3563,I139418,I139642,);
DFFARX1 I_8003 (I139642,I3563,I139418,I139407,);
nand I_8004 (I139664,I580401,I580407);
and I_8005 (I139681,I139664,I580383);
DFFARX1 I_8006 (I139681,I3563,I139418,I139707,);
DFFARX1 I_8007 (I139707,I3563,I139418,I139724,);
not I_8008 (I139410,I139724);
not I_8009 (I139746,I139707);
nand I_8010 (I139395,I139746,I139585);
nor I_8011 (I139777,I580386,I580407);
not I_8012 (I139794,I139777);
nor I_8013 (I139811,I139746,I139794);
nor I_8014 (I139828,I139452,I139811);
DFFARX1 I_8015 (I139828,I3563,I139418,I139404,);
nor I_8016 (I139859,I139512,I139794);
nor I_8017 (I139392,I139707,I139859);
nor I_8018 (I139401,I139642,I139777);
nor I_8019 (I139389,I139512,I139777);
not I_8020 (I139945,I3570);
DFFARX1 I_8021 (I668251,I3563,I139945,I139971,);
not I_8022 (I139979,I139971);
nand I_8023 (I139996,I668242,I668260);
and I_8024 (I140013,I139996,I668239);
DFFARX1 I_8025 (I140013,I3563,I139945,I140039,);
DFFARX1 I_8026 (I668242,I3563,I139945,I140056,);
and I_8027 (I140064,I140056,I668245);
nor I_8028 (I140081,I140039,I140064);
DFFARX1 I_8029 (I140081,I3563,I139945,I139913,);
nand I_8030 (I140112,I140056,I668245);
nand I_8031 (I140129,I139979,I140112);
not I_8032 (I139925,I140129);
DFFARX1 I_8033 (I668239,I3563,I139945,I140169,);
DFFARX1 I_8034 (I140169,I3563,I139945,I139934,);
nand I_8035 (I140191,I668257,I668248);
and I_8036 (I140208,I140191,I668263);
DFFARX1 I_8037 (I140208,I3563,I139945,I140234,);
DFFARX1 I_8038 (I140234,I3563,I139945,I140251,);
not I_8039 (I139937,I140251);
not I_8040 (I140273,I140234);
nand I_8041 (I139922,I140273,I140112);
nor I_8042 (I140304,I668254,I668248);
not I_8043 (I140321,I140304);
nor I_8044 (I140338,I140273,I140321);
nor I_8045 (I140355,I139979,I140338);
DFFARX1 I_8046 (I140355,I3563,I139945,I139931,);
nor I_8047 (I140386,I140039,I140321);
nor I_8048 (I139919,I140234,I140386);
nor I_8049 (I139928,I140169,I140304);
nor I_8050 (I139916,I140039,I140304);
not I_8051 (I140472,I3570);
DFFARX1 I_8052 (I952998,I3563,I140472,I140498,);
not I_8053 (I140506,I140498);
nand I_8054 (I140523,I953016,I953010);
and I_8055 (I140540,I140523,I952989);
DFFARX1 I_8056 (I140540,I3563,I140472,I140566,);
DFFARX1 I_8057 (I953007,I3563,I140472,I140583,);
and I_8058 (I140591,I140583,I952992);
nor I_8059 (I140608,I140566,I140591);
DFFARX1 I_8060 (I140608,I3563,I140472,I140440,);
nand I_8061 (I140639,I140583,I952992);
nand I_8062 (I140656,I140506,I140639);
not I_8063 (I140452,I140656);
DFFARX1 I_8064 (I953004,I3563,I140472,I140696,);
DFFARX1 I_8065 (I140696,I3563,I140472,I140461,);
nand I_8066 (I140718,I953013,I953001);
and I_8067 (I140735,I140718,I952995);
DFFARX1 I_8068 (I140735,I3563,I140472,I140761,);
DFFARX1 I_8069 (I140761,I3563,I140472,I140778,);
not I_8070 (I140464,I140778);
not I_8071 (I140800,I140761);
nand I_8072 (I140449,I140800,I140639);
nor I_8073 (I140831,I952989,I953001);
not I_8074 (I140848,I140831);
nor I_8075 (I140865,I140800,I140848);
nor I_8076 (I140882,I140506,I140865);
DFFARX1 I_8077 (I140882,I3563,I140472,I140458,);
nor I_8078 (I140913,I140566,I140848);
nor I_8079 (I140446,I140761,I140913);
nor I_8080 (I140455,I140696,I140831);
nor I_8081 (I140443,I140566,I140831);
not I_8082 (I140999,I3570);
DFFARX1 I_8083 (I685591,I3563,I140999,I141025,);
not I_8084 (I141033,I141025);
nand I_8085 (I141050,I685582,I685600);
and I_8086 (I141067,I141050,I685579);
DFFARX1 I_8087 (I141067,I3563,I140999,I141093,);
DFFARX1 I_8088 (I685582,I3563,I140999,I141110,);
and I_8089 (I141118,I141110,I685585);
nor I_8090 (I141135,I141093,I141118);
DFFARX1 I_8091 (I141135,I3563,I140999,I140967,);
nand I_8092 (I141166,I141110,I685585);
nand I_8093 (I141183,I141033,I141166);
not I_8094 (I140979,I141183);
DFFARX1 I_8095 (I685579,I3563,I140999,I141223,);
DFFARX1 I_8096 (I141223,I3563,I140999,I140988,);
nand I_8097 (I141245,I685597,I685588);
and I_8098 (I141262,I141245,I685603);
DFFARX1 I_8099 (I141262,I3563,I140999,I141288,);
DFFARX1 I_8100 (I141288,I3563,I140999,I141305,);
not I_8101 (I140991,I141305);
not I_8102 (I141327,I141288);
nand I_8103 (I140976,I141327,I141166);
nor I_8104 (I141358,I685594,I685588);
not I_8105 (I141375,I141358);
nor I_8106 (I141392,I141327,I141375);
nor I_8107 (I141409,I141033,I141392);
DFFARX1 I_8108 (I141409,I3563,I140999,I140985,);
nor I_8109 (I141440,I141093,I141375);
nor I_8110 (I140973,I141288,I141440);
nor I_8111 (I140982,I141223,I141358);
nor I_8112 (I140970,I141093,I141358);
not I_8113 (I141526,I3570);
DFFARX1 I_8114 (I1053955,I3563,I141526,I141552,);
not I_8115 (I141560,I141552);
nand I_8116 (I141577,I1053952,I1053958);
and I_8117 (I141594,I141577,I1053955);
DFFARX1 I_8118 (I141594,I3563,I141526,I141620,);
DFFARX1 I_8119 (I1053958,I3563,I141526,I141637,);
and I_8120 (I141645,I141637,I1053952);
nor I_8121 (I141662,I141620,I141645);
DFFARX1 I_8122 (I141662,I3563,I141526,I141494,);
nand I_8123 (I141693,I141637,I1053952);
nand I_8124 (I141710,I141560,I141693);
not I_8125 (I141506,I141710);
DFFARX1 I_8126 (I1053961,I3563,I141526,I141750,);
DFFARX1 I_8127 (I141750,I3563,I141526,I141515,);
nand I_8128 (I141772,I1053964,I1053973);
and I_8129 (I141789,I141772,I1053967);
DFFARX1 I_8130 (I141789,I3563,I141526,I141815,);
DFFARX1 I_8131 (I141815,I3563,I141526,I141832,);
not I_8132 (I141518,I141832);
not I_8133 (I141854,I141815);
nand I_8134 (I141503,I141854,I141693);
nor I_8135 (I141885,I1053970,I1053973);
not I_8136 (I141902,I141885);
nor I_8137 (I141919,I141854,I141902);
nor I_8138 (I141936,I141560,I141919);
DFFARX1 I_8139 (I141936,I3563,I141526,I141512,);
nor I_8140 (I141967,I141620,I141902);
nor I_8141 (I141500,I141815,I141967);
nor I_8142 (I141509,I141750,I141885);
nor I_8143 (I141497,I141620,I141885);
not I_8144 (I142053,I3570);
DFFARX1 I_8145 (I1070785,I3563,I142053,I142079,);
not I_8146 (I142087,I142079);
nand I_8147 (I142104,I1070782,I1070788);
and I_8148 (I142121,I142104,I1070785);
DFFARX1 I_8149 (I142121,I3563,I142053,I142147,);
DFFARX1 I_8150 (I1070788,I3563,I142053,I142164,);
and I_8151 (I142172,I142164,I1070782);
nor I_8152 (I142189,I142147,I142172);
DFFARX1 I_8153 (I142189,I3563,I142053,I142021,);
nand I_8154 (I142220,I142164,I1070782);
nand I_8155 (I142237,I142087,I142220);
not I_8156 (I142033,I142237);
DFFARX1 I_8157 (I1070791,I3563,I142053,I142277,);
DFFARX1 I_8158 (I142277,I3563,I142053,I142042,);
nand I_8159 (I142299,I1070794,I1070803);
and I_8160 (I142316,I142299,I1070797);
DFFARX1 I_8161 (I142316,I3563,I142053,I142342,);
DFFARX1 I_8162 (I142342,I3563,I142053,I142359,);
not I_8163 (I142045,I142359);
not I_8164 (I142381,I142342);
nand I_8165 (I142030,I142381,I142220);
nor I_8166 (I142412,I1070800,I1070803);
not I_8167 (I142429,I142412);
nor I_8168 (I142446,I142381,I142429);
nor I_8169 (I142463,I142087,I142446);
DFFARX1 I_8170 (I142463,I3563,I142053,I142039,);
nor I_8171 (I142494,I142147,I142429);
nor I_8172 (I142027,I142342,I142494);
nor I_8173 (I142036,I142277,I142412);
nor I_8174 (I142024,I142147,I142412);
not I_8175 (I142580,I3570);
DFFARX1 I_8176 (I605824,I3563,I142580,I142606,);
not I_8177 (I142614,I142606);
nand I_8178 (I142631,I605836,I605821);
and I_8179 (I142648,I142631,I605815);
DFFARX1 I_8180 (I142648,I3563,I142580,I142674,);
DFFARX1 I_8181 (I605830,I3563,I142580,I142691,);
and I_8182 (I142699,I142691,I605818);
nor I_8183 (I142716,I142674,I142699);
DFFARX1 I_8184 (I142716,I3563,I142580,I142548,);
nand I_8185 (I142747,I142691,I605818);
nand I_8186 (I142764,I142614,I142747);
not I_8187 (I142560,I142764);
DFFARX1 I_8188 (I605827,I3563,I142580,I142804,);
DFFARX1 I_8189 (I142804,I3563,I142580,I142569,);
nand I_8190 (I142826,I605833,I605839);
and I_8191 (I142843,I142826,I605815);
DFFARX1 I_8192 (I142843,I3563,I142580,I142869,);
DFFARX1 I_8193 (I142869,I3563,I142580,I142886,);
not I_8194 (I142572,I142886);
not I_8195 (I142908,I142869);
nand I_8196 (I142557,I142908,I142747);
nor I_8197 (I142939,I605818,I605839);
not I_8198 (I142956,I142939);
nor I_8199 (I142973,I142908,I142956);
nor I_8200 (I142990,I142614,I142973);
DFFARX1 I_8201 (I142990,I3563,I142580,I142566,);
nor I_8202 (I143021,I142674,I142956);
nor I_8203 (I142554,I142869,I143021);
nor I_8204 (I142563,I142804,I142939);
nor I_8205 (I142551,I142674,I142939);
not I_8206 (I143107,I3570);
DFFARX1 I_8207 (I1263823,I3563,I143107,I143133,);
not I_8208 (I143141,I143133);
nand I_8209 (I143158,I1263817,I1263838);
and I_8210 (I143175,I143158,I1263829);
DFFARX1 I_8211 (I143175,I3563,I143107,I143201,);
DFFARX1 I_8212 (I1263820,I3563,I143107,I143218,);
and I_8213 (I143226,I143218,I1263832);
nor I_8214 (I143243,I143201,I143226);
DFFARX1 I_8215 (I143243,I3563,I143107,I143075,);
nand I_8216 (I143274,I143218,I1263832);
nand I_8217 (I143291,I143141,I143274);
not I_8218 (I143087,I143291);
DFFARX1 I_8219 (I1263820,I3563,I143107,I143331,);
DFFARX1 I_8220 (I143331,I3563,I143107,I143096,);
nand I_8221 (I143353,I1263841,I1263826);
and I_8222 (I143370,I143353,I1263817);
DFFARX1 I_8223 (I143370,I3563,I143107,I143396,);
DFFARX1 I_8224 (I143396,I3563,I143107,I143413,);
not I_8225 (I143099,I143413);
not I_8226 (I143435,I143396);
nand I_8227 (I143084,I143435,I143274);
nor I_8228 (I143466,I1263835,I1263826);
not I_8229 (I143483,I143466);
nor I_8230 (I143500,I143435,I143483);
nor I_8231 (I143517,I143141,I143500);
DFFARX1 I_8232 (I143517,I3563,I143107,I143093,);
nor I_8233 (I143548,I143201,I143483);
nor I_8234 (I143081,I143396,I143548);
nor I_8235 (I143090,I143331,I143466);
nor I_8236 (I143078,I143201,I143466);
not I_8237 (I143634,I3570);
DFFARX1 I_8238 (I450708,I3563,I143634,I143660,);
not I_8239 (I143668,I143660);
nand I_8240 (I143685,I450702,I450693);
and I_8241 (I143702,I143685,I450714);
DFFARX1 I_8242 (I143702,I3563,I143634,I143728,);
DFFARX1 I_8243 (I450696,I3563,I143634,I143745,);
and I_8244 (I143753,I143745,I450690);
nor I_8245 (I143770,I143728,I143753);
DFFARX1 I_8246 (I143770,I3563,I143634,I143602,);
nand I_8247 (I143801,I143745,I450690);
nand I_8248 (I143818,I143668,I143801);
not I_8249 (I143614,I143818);
DFFARX1 I_8250 (I450690,I3563,I143634,I143858,);
DFFARX1 I_8251 (I143858,I3563,I143634,I143623,);
nand I_8252 (I143880,I450717,I450699);
and I_8253 (I143897,I143880,I450705);
DFFARX1 I_8254 (I143897,I3563,I143634,I143923,);
DFFARX1 I_8255 (I143923,I3563,I143634,I143940,);
not I_8256 (I143626,I143940);
not I_8257 (I143962,I143923);
nand I_8258 (I143611,I143962,I143801);
nor I_8259 (I143993,I450711,I450699);
not I_8260 (I144010,I143993);
nor I_8261 (I144027,I143962,I144010);
nor I_8262 (I144044,I143668,I144027);
DFFARX1 I_8263 (I144044,I3563,I143634,I143620,);
nor I_8264 (I144075,I143728,I144010);
nor I_8265 (I143608,I143923,I144075);
nor I_8266 (I143617,I143858,I143993);
nor I_8267 (I143605,I143728,I143993);
not I_8268 (I144161,I3570);
DFFARX1 I_8269 (I383414,I3563,I144161,I144187,);
not I_8270 (I144195,I144187);
nand I_8271 (I144212,I383396,I383411);
and I_8272 (I144229,I144212,I383387);
DFFARX1 I_8273 (I144229,I3563,I144161,I144255,);
DFFARX1 I_8274 (I383390,I3563,I144161,I144272,);
and I_8275 (I144280,I144272,I383405);
nor I_8276 (I144297,I144255,I144280);
DFFARX1 I_8277 (I144297,I3563,I144161,I144129,);
nand I_8278 (I144328,I144272,I383405);
nand I_8279 (I144345,I144195,I144328);
not I_8280 (I144141,I144345);
DFFARX1 I_8281 (I383408,I3563,I144161,I144385,);
DFFARX1 I_8282 (I144385,I3563,I144161,I144150,);
nand I_8283 (I144407,I383387,I383399);
and I_8284 (I144424,I144407,I383393);
DFFARX1 I_8285 (I144424,I3563,I144161,I144450,);
DFFARX1 I_8286 (I144450,I3563,I144161,I144467,);
not I_8287 (I144153,I144467);
not I_8288 (I144489,I144450);
nand I_8289 (I144138,I144489,I144328);
nor I_8290 (I144520,I383402,I383399);
not I_8291 (I144537,I144520);
nor I_8292 (I144554,I144489,I144537);
nor I_8293 (I144571,I144195,I144554);
DFFARX1 I_8294 (I144571,I3563,I144161,I144147,);
nor I_8295 (I144602,I144255,I144537);
nor I_8296 (I144135,I144450,I144602);
nor I_8297 (I144144,I144385,I144520);
nor I_8298 (I144132,I144255,I144520);
not I_8299 (I144688,I3570);
DFFARX1 I_8300 (I306999,I3563,I144688,I144714,);
not I_8301 (I144722,I144714);
nand I_8302 (I144739,I306981,I306996);
and I_8303 (I144756,I144739,I306972);
DFFARX1 I_8304 (I144756,I3563,I144688,I144782,);
DFFARX1 I_8305 (I306975,I3563,I144688,I144799,);
and I_8306 (I144807,I144799,I306990);
nor I_8307 (I144824,I144782,I144807);
DFFARX1 I_8308 (I144824,I3563,I144688,I144656,);
nand I_8309 (I144855,I144799,I306990);
nand I_8310 (I144872,I144722,I144855);
not I_8311 (I144668,I144872);
DFFARX1 I_8312 (I306993,I3563,I144688,I144912,);
DFFARX1 I_8313 (I144912,I3563,I144688,I144677,);
nand I_8314 (I144934,I306972,I306984);
and I_8315 (I144951,I144934,I306978);
DFFARX1 I_8316 (I144951,I3563,I144688,I144977,);
DFFARX1 I_8317 (I144977,I3563,I144688,I144994,);
not I_8318 (I144680,I144994);
not I_8319 (I145016,I144977);
nand I_8320 (I144665,I145016,I144855);
nor I_8321 (I145047,I306987,I306984);
not I_8322 (I145064,I145047);
nor I_8323 (I145081,I145016,I145064);
nor I_8324 (I145098,I144722,I145081);
DFFARX1 I_8325 (I145098,I3563,I144688,I144674,);
nor I_8326 (I145129,I144782,I145064);
nor I_8327 (I144662,I144977,I145129);
nor I_8328 (I144671,I144912,I145047);
nor I_8329 (I144659,I144782,I145047);
not I_8330 (I145215,I3570);
DFFARX1 I_8331 (I1294710,I3563,I145215,I145241,);
not I_8332 (I145249,I145241);
nand I_8333 (I145266,I1294713,I1294707);
and I_8334 (I145283,I145266,I1294704);
DFFARX1 I_8335 (I145283,I3563,I145215,I145309,);
DFFARX1 I_8336 (I1294689,I3563,I145215,I145326,);
and I_8337 (I145334,I145326,I1294698);
nor I_8338 (I145351,I145309,I145334);
DFFARX1 I_8339 (I145351,I3563,I145215,I145183,);
nand I_8340 (I145382,I145326,I1294698);
nand I_8341 (I145399,I145249,I145382);
not I_8342 (I145195,I145399);
DFFARX1 I_8343 (I1294689,I3563,I145215,I145439,);
DFFARX1 I_8344 (I145439,I3563,I145215,I145204,);
nand I_8345 (I145461,I1294692,I1294695);
and I_8346 (I145478,I145461,I1294701);
DFFARX1 I_8347 (I145478,I3563,I145215,I145504,);
DFFARX1 I_8348 (I145504,I3563,I145215,I145521,);
not I_8349 (I145207,I145521);
not I_8350 (I145543,I145504);
nand I_8351 (I145192,I145543,I145382);
nor I_8352 (I145574,I1294692,I1294695);
not I_8353 (I145591,I145574);
nor I_8354 (I145608,I145543,I145591);
nor I_8355 (I145625,I145249,I145608);
DFFARX1 I_8356 (I145625,I3563,I145215,I145201,);
nor I_8357 (I145656,I145309,I145591);
nor I_8358 (I145189,I145504,I145656);
nor I_8359 (I145198,I145439,I145574);
nor I_8360 (I145186,I145309,I145574);
not I_8361 (I145742,I3570);
DFFARX1 I_8362 (I353375,I3563,I145742,I145768,);
not I_8363 (I145776,I145768);
nand I_8364 (I145793,I353357,I353372);
and I_8365 (I145810,I145793,I353348);
DFFARX1 I_8366 (I145810,I3563,I145742,I145836,);
DFFARX1 I_8367 (I353351,I3563,I145742,I145853,);
and I_8368 (I145861,I145853,I353366);
nor I_8369 (I145878,I145836,I145861);
DFFARX1 I_8370 (I145878,I3563,I145742,I145710,);
nand I_8371 (I145909,I145853,I353366);
nand I_8372 (I145926,I145776,I145909);
not I_8373 (I145722,I145926);
DFFARX1 I_8374 (I353369,I3563,I145742,I145966,);
DFFARX1 I_8375 (I145966,I3563,I145742,I145731,);
nand I_8376 (I145988,I353348,I353360);
and I_8377 (I146005,I145988,I353354);
DFFARX1 I_8378 (I146005,I3563,I145742,I146031,);
DFFARX1 I_8379 (I146031,I3563,I145742,I146048,);
not I_8380 (I145734,I146048);
not I_8381 (I146070,I146031);
nand I_8382 (I145719,I146070,I145909);
nor I_8383 (I146101,I353363,I353360);
not I_8384 (I146118,I146101);
nor I_8385 (I146135,I146070,I146118);
nor I_8386 (I146152,I145776,I146135);
DFFARX1 I_8387 (I146152,I3563,I145742,I145728,);
nor I_8388 (I146183,I145836,I146118);
nor I_8389 (I145716,I146031,I146183);
nor I_8390 (I145725,I145966,I146101);
nor I_8391 (I145713,I145836,I146101);
not I_8392 (I146269,I3570);
DFFARX1 I_8393 (I732409,I3563,I146269,I146295,);
not I_8394 (I146303,I146295);
nand I_8395 (I146320,I732400,I732418);
and I_8396 (I146337,I146320,I732397);
DFFARX1 I_8397 (I146337,I3563,I146269,I146363,);
DFFARX1 I_8398 (I732400,I3563,I146269,I146380,);
and I_8399 (I146388,I146380,I732403);
nor I_8400 (I146405,I146363,I146388);
DFFARX1 I_8401 (I146405,I3563,I146269,I146237,);
nand I_8402 (I146436,I146380,I732403);
nand I_8403 (I146453,I146303,I146436);
not I_8404 (I146249,I146453);
DFFARX1 I_8405 (I732397,I3563,I146269,I146493,);
DFFARX1 I_8406 (I146493,I3563,I146269,I146258,);
nand I_8407 (I146515,I732415,I732406);
and I_8408 (I146532,I146515,I732421);
DFFARX1 I_8409 (I146532,I3563,I146269,I146558,);
DFFARX1 I_8410 (I146558,I3563,I146269,I146575,);
not I_8411 (I146261,I146575);
not I_8412 (I146597,I146558);
nand I_8413 (I146246,I146597,I146436);
nor I_8414 (I146628,I732412,I732406);
not I_8415 (I146645,I146628);
nor I_8416 (I146662,I146597,I146645);
nor I_8417 (I146679,I146303,I146662);
DFFARX1 I_8418 (I146679,I3563,I146269,I146255,);
nor I_8419 (I146710,I146363,I146645);
nor I_8420 (I146243,I146558,I146710);
nor I_8421 (I146252,I146493,I146628);
nor I_8422 (I146240,I146363,I146628);
not I_8423 (I146796,I3570);
DFFARX1 I_8424 (I334930,I3563,I146796,I146822,);
not I_8425 (I146830,I146822);
nand I_8426 (I146847,I334912,I334927);
and I_8427 (I146864,I146847,I334903);
DFFARX1 I_8428 (I146864,I3563,I146796,I146890,);
DFFARX1 I_8429 (I334906,I3563,I146796,I146907,);
and I_8430 (I146915,I146907,I334921);
nor I_8431 (I146932,I146890,I146915);
DFFARX1 I_8432 (I146932,I3563,I146796,I146764,);
nand I_8433 (I146963,I146907,I334921);
nand I_8434 (I146980,I146830,I146963);
not I_8435 (I146776,I146980);
DFFARX1 I_8436 (I334924,I3563,I146796,I147020,);
DFFARX1 I_8437 (I147020,I3563,I146796,I146785,);
nand I_8438 (I147042,I334903,I334915);
and I_8439 (I147059,I147042,I334909);
DFFARX1 I_8440 (I147059,I3563,I146796,I147085,);
DFFARX1 I_8441 (I147085,I3563,I146796,I147102,);
not I_8442 (I146788,I147102);
not I_8443 (I147124,I147085);
nand I_8444 (I146773,I147124,I146963);
nor I_8445 (I147155,I334918,I334915);
not I_8446 (I147172,I147155);
nor I_8447 (I147189,I147124,I147172);
nor I_8448 (I147206,I146830,I147189);
DFFARX1 I_8449 (I147206,I3563,I146796,I146782,);
nor I_8450 (I147237,I146890,I147172);
nor I_8451 (I146770,I147085,I147237);
nor I_8452 (I146779,I147020,I147155);
nor I_8453 (I146767,I146890,I147155);
not I_8454 (I147323,I3570);
DFFARX1 I_8455 (I207755,I3563,I147323,I147349,);
not I_8456 (I147357,I147349);
nand I_8457 (I147374,I207749,I207743);
and I_8458 (I147391,I147374,I207764);
DFFARX1 I_8459 (I147391,I3563,I147323,I147417,);
DFFARX1 I_8460 (I207761,I3563,I147323,I147434,);
and I_8461 (I147442,I147434,I207758);
nor I_8462 (I147459,I147417,I147442);
DFFARX1 I_8463 (I147459,I3563,I147323,I147291,);
nand I_8464 (I147490,I147434,I207758);
nand I_8465 (I147507,I147357,I147490);
not I_8466 (I147303,I147507);
DFFARX1 I_8467 (I207743,I3563,I147323,I147547,);
DFFARX1 I_8468 (I147547,I3563,I147323,I147312,);
nand I_8469 (I147569,I207746,I207746);
and I_8470 (I147586,I147569,I207767);
DFFARX1 I_8471 (I147586,I3563,I147323,I147612,);
DFFARX1 I_8472 (I147612,I3563,I147323,I147629,);
not I_8473 (I147315,I147629);
not I_8474 (I147651,I147612);
nand I_8475 (I147300,I147651,I147490);
nor I_8476 (I147682,I207752,I207746);
not I_8477 (I147699,I147682);
nor I_8478 (I147716,I147651,I147699);
nor I_8479 (I147733,I147357,I147716);
DFFARX1 I_8480 (I147733,I3563,I147323,I147309,);
nor I_8481 (I147764,I147417,I147699);
nor I_8482 (I147297,I147612,I147764);
nor I_8483 (I147306,I147547,I147682);
nor I_8484 (I147294,I147417,I147682);
not I_8485 (I147850,I3570);
DFFARX1 I_8486 (I316485,I3563,I147850,I147876,);
not I_8487 (I147884,I147876);
nand I_8488 (I147901,I316467,I316482);
and I_8489 (I147918,I147901,I316458);
DFFARX1 I_8490 (I147918,I3563,I147850,I147944,);
DFFARX1 I_8491 (I316461,I3563,I147850,I147961,);
and I_8492 (I147969,I147961,I316476);
nor I_8493 (I147986,I147944,I147969);
DFFARX1 I_8494 (I147986,I3563,I147850,I147818,);
nand I_8495 (I148017,I147961,I316476);
nand I_8496 (I148034,I147884,I148017);
not I_8497 (I147830,I148034);
DFFARX1 I_8498 (I316479,I3563,I147850,I148074,);
DFFARX1 I_8499 (I148074,I3563,I147850,I147839,);
nand I_8500 (I148096,I316458,I316470);
and I_8501 (I148113,I148096,I316464);
DFFARX1 I_8502 (I148113,I3563,I147850,I148139,);
DFFARX1 I_8503 (I148139,I3563,I147850,I148156,);
not I_8504 (I147842,I148156);
not I_8505 (I148178,I148139);
nand I_8506 (I147827,I148178,I148017);
nor I_8507 (I148209,I316473,I316470);
not I_8508 (I148226,I148209);
nor I_8509 (I148243,I148178,I148226);
nor I_8510 (I148260,I147884,I148243);
DFFARX1 I_8511 (I148260,I3563,I147850,I147836,);
nor I_8512 (I148291,I147944,I148226);
nor I_8513 (I147824,I148139,I148291);
nor I_8514 (I147833,I148074,I148209);
nor I_8515 (I147821,I147944,I148209);
not I_8516 (I148377,I3570);
DFFARX1 I_8517 (I702931,I3563,I148377,I148403,);
not I_8518 (I148411,I148403);
nand I_8519 (I148428,I702922,I702940);
and I_8520 (I148445,I148428,I702919);
DFFARX1 I_8521 (I148445,I3563,I148377,I148471,);
DFFARX1 I_8522 (I702922,I3563,I148377,I148488,);
and I_8523 (I148496,I148488,I702925);
nor I_8524 (I148513,I148471,I148496);
DFFARX1 I_8525 (I148513,I3563,I148377,I148345,);
nand I_8526 (I148544,I148488,I702925);
nand I_8527 (I148561,I148411,I148544);
not I_8528 (I148357,I148561);
DFFARX1 I_8529 (I702919,I3563,I148377,I148601,);
DFFARX1 I_8530 (I148601,I3563,I148377,I148366,);
nand I_8531 (I148623,I702937,I702928);
and I_8532 (I148640,I148623,I702943);
DFFARX1 I_8533 (I148640,I3563,I148377,I148666,);
DFFARX1 I_8534 (I148666,I3563,I148377,I148683,);
not I_8535 (I148369,I148683);
not I_8536 (I148705,I148666);
nand I_8537 (I148354,I148705,I148544);
nor I_8538 (I148736,I702934,I702928);
not I_8539 (I148753,I148736);
nor I_8540 (I148770,I148705,I148753);
nor I_8541 (I148787,I148411,I148770);
DFFARX1 I_8542 (I148787,I3563,I148377,I148363,);
nor I_8543 (I148818,I148471,I148753);
nor I_8544 (I148351,I148666,I148818);
nor I_8545 (I148360,I148601,I148736);
nor I_8546 (I148348,I148471,I148736);
not I_8547 (I148904,I3570);
DFFARX1 I_8548 (I694261,I3563,I148904,I148930,);
not I_8549 (I148938,I148930);
nand I_8550 (I148955,I694252,I694270);
and I_8551 (I148972,I148955,I694249);
DFFARX1 I_8552 (I148972,I3563,I148904,I148998,);
DFFARX1 I_8553 (I694252,I3563,I148904,I149015,);
and I_8554 (I149023,I149015,I694255);
nor I_8555 (I149040,I148998,I149023);
DFFARX1 I_8556 (I149040,I3563,I148904,I148872,);
nand I_8557 (I149071,I149015,I694255);
nand I_8558 (I149088,I148938,I149071);
not I_8559 (I148884,I149088);
DFFARX1 I_8560 (I694249,I3563,I148904,I149128,);
DFFARX1 I_8561 (I149128,I3563,I148904,I148893,);
nand I_8562 (I149150,I694267,I694258);
and I_8563 (I149167,I149150,I694273);
DFFARX1 I_8564 (I149167,I3563,I148904,I149193,);
DFFARX1 I_8565 (I149193,I3563,I148904,I149210,);
not I_8566 (I148896,I149210);
not I_8567 (I149232,I149193);
nand I_8568 (I148881,I149232,I149071);
nor I_8569 (I149263,I694264,I694258);
not I_8570 (I149280,I149263);
nor I_8571 (I149297,I149232,I149280);
nor I_8572 (I149314,I148938,I149297);
DFFARX1 I_8573 (I149314,I3563,I148904,I148890,);
nor I_8574 (I149345,I148998,I149280);
nor I_8575 (I148878,I149193,I149345);
nor I_8576 (I148887,I149128,I149263);
nor I_8577 (I148875,I148998,I149263);
not I_8578 (I149431,I3570);
DFFARX1 I_8579 (I1239547,I3563,I149431,I149457,);
not I_8580 (I149465,I149457);
nand I_8581 (I149482,I1239562,I1239541);
and I_8582 (I149499,I149482,I1239544);
DFFARX1 I_8583 (I149499,I3563,I149431,I149525,);
DFFARX1 I_8584 (I1239565,I3563,I149431,I149542,);
and I_8585 (I149550,I149542,I1239544);
nor I_8586 (I149567,I149525,I149550);
DFFARX1 I_8587 (I149567,I3563,I149431,I149399,);
nand I_8588 (I149598,I149542,I1239544);
nand I_8589 (I149615,I149465,I149598);
not I_8590 (I149411,I149615);
DFFARX1 I_8591 (I1239541,I3563,I149431,I149655,);
DFFARX1 I_8592 (I149655,I3563,I149431,I149420,);
nand I_8593 (I149677,I1239553,I1239550);
and I_8594 (I149694,I149677,I1239556);
DFFARX1 I_8595 (I149694,I3563,I149431,I149720,);
DFFARX1 I_8596 (I149720,I3563,I149431,I149737,);
not I_8597 (I149423,I149737);
not I_8598 (I149759,I149720);
nand I_8599 (I149408,I149759,I149598);
nor I_8600 (I149790,I1239559,I1239550);
not I_8601 (I149807,I149790);
nor I_8602 (I149824,I149759,I149807);
nor I_8603 (I149841,I149465,I149824);
DFFARX1 I_8604 (I149841,I3563,I149431,I149417,);
nor I_8605 (I149872,I149525,I149807);
nor I_8606 (I149405,I149720,I149872);
nor I_8607 (I149414,I149655,I149790);
nor I_8608 (I149402,I149525,I149790);
not I_8609 (I149958,I3570);
DFFARX1 I_8610 (I1057882,I3563,I149958,I149984,);
not I_8611 (I149992,I149984);
nand I_8612 (I150009,I1057879,I1057885);
and I_8613 (I150026,I150009,I1057882);
DFFARX1 I_8614 (I150026,I3563,I149958,I150052,);
DFFARX1 I_8615 (I1057885,I3563,I149958,I150069,);
and I_8616 (I150077,I150069,I1057879);
nor I_8617 (I150094,I150052,I150077);
DFFARX1 I_8618 (I150094,I3563,I149958,I149926,);
nand I_8619 (I150125,I150069,I1057879);
nand I_8620 (I150142,I149992,I150125);
not I_8621 (I149938,I150142);
DFFARX1 I_8622 (I1057888,I3563,I149958,I150182,);
DFFARX1 I_8623 (I150182,I3563,I149958,I149947,);
nand I_8624 (I150204,I1057891,I1057900);
and I_8625 (I150221,I150204,I1057894);
DFFARX1 I_8626 (I150221,I3563,I149958,I150247,);
DFFARX1 I_8627 (I150247,I3563,I149958,I150264,);
not I_8628 (I149950,I150264);
not I_8629 (I150286,I150247);
nand I_8630 (I149935,I150286,I150125);
nor I_8631 (I150317,I1057897,I1057900);
not I_8632 (I150334,I150317);
nor I_8633 (I150351,I150286,I150334);
nor I_8634 (I150368,I149992,I150351);
DFFARX1 I_8635 (I150368,I3563,I149958,I149944,);
nor I_8636 (I150399,I150052,I150334);
nor I_8637 (I149932,I150247,I150399);
nor I_8638 (I149941,I150182,I150317);
nor I_8639 (I149929,I150052,I150317);
not I_8640 (I150485,I3570);
DFFARX1 I_8641 (I843739,I3563,I150485,I150511,);
not I_8642 (I150519,I150511);
nand I_8643 (I150536,I843736,I843751);
and I_8644 (I150553,I150536,I843733);
DFFARX1 I_8645 (I150553,I3563,I150485,I150579,);
DFFARX1 I_8646 (I843730,I3563,I150485,I150596,);
and I_8647 (I150604,I150596,I843730);
nor I_8648 (I150621,I150579,I150604);
DFFARX1 I_8649 (I150621,I3563,I150485,I150453,);
nand I_8650 (I150652,I150596,I843730);
nand I_8651 (I150669,I150519,I150652);
not I_8652 (I150465,I150669);
DFFARX1 I_8653 (I843733,I3563,I150485,I150709,);
DFFARX1 I_8654 (I150709,I3563,I150485,I150474,);
nand I_8655 (I150731,I843745,I843736);
and I_8656 (I150748,I150731,I843748);
DFFARX1 I_8657 (I150748,I3563,I150485,I150774,);
DFFARX1 I_8658 (I150774,I3563,I150485,I150791,);
not I_8659 (I150477,I150791);
not I_8660 (I150813,I150774);
nand I_8661 (I150462,I150813,I150652);
nor I_8662 (I150844,I843742,I843736);
not I_8663 (I150861,I150844);
nor I_8664 (I150878,I150813,I150861);
nor I_8665 (I150895,I150519,I150878);
DFFARX1 I_8666 (I150895,I3563,I150485,I150471,);
nor I_8667 (I150926,I150579,I150861);
nor I_8668 (I150459,I150774,I150926);
nor I_8669 (I150468,I150709,I150844);
nor I_8670 (I150456,I150579,I150844);
not I_8671 (I151012,I3570);
DFFARX1 I_8672 (I381833,I3563,I151012,I151038,);
not I_8673 (I151046,I151038);
nand I_8674 (I151063,I381815,I381830);
and I_8675 (I151080,I151063,I381806);
DFFARX1 I_8676 (I151080,I3563,I151012,I151106,);
DFFARX1 I_8677 (I381809,I3563,I151012,I151123,);
and I_8678 (I151131,I151123,I381824);
nor I_8679 (I151148,I151106,I151131);
DFFARX1 I_8680 (I151148,I3563,I151012,I150980,);
nand I_8681 (I151179,I151123,I381824);
nand I_8682 (I151196,I151046,I151179);
not I_8683 (I150992,I151196);
DFFARX1 I_8684 (I381827,I3563,I151012,I151236,);
DFFARX1 I_8685 (I151236,I3563,I151012,I151001,);
nand I_8686 (I151258,I381806,I381818);
and I_8687 (I151275,I151258,I381812);
DFFARX1 I_8688 (I151275,I3563,I151012,I151301,);
DFFARX1 I_8689 (I151301,I3563,I151012,I151318,);
not I_8690 (I151004,I151318);
not I_8691 (I151340,I151301);
nand I_8692 (I150989,I151340,I151179);
nor I_8693 (I151371,I381821,I381818);
not I_8694 (I151388,I151371);
nor I_8695 (I151405,I151340,I151388);
nor I_8696 (I151422,I151046,I151405);
DFFARX1 I_8697 (I151422,I3563,I151012,I150998,);
nor I_8698 (I151453,I151106,I151388);
nor I_8699 (I150986,I151301,I151453);
nor I_8700 (I150995,I151236,I151371);
nor I_8701 (I150983,I151106,I151371);
not I_8702 (I151539,I3570);
DFFARX1 I_8703 (I1052272,I3563,I151539,I151565,);
not I_8704 (I151573,I151565);
nand I_8705 (I151590,I1052269,I1052275);
and I_8706 (I151607,I151590,I1052272);
DFFARX1 I_8707 (I151607,I3563,I151539,I151633,);
DFFARX1 I_8708 (I1052275,I3563,I151539,I151650,);
and I_8709 (I151658,I151650,I1052269);
nor I_8710 (I151675,I151633,I151658);
DFFARX1 I_8711 (I151675,I3563,I151539,I151507,);
nand I_8712 (I151706,I151650,I1052269);
nand I_8713 (I151723,I151573,I151706);
not I_8714 (I151519,I151723);
DFFARX1 I_8715 (I1052278,I3563,I151539,I151763,);
DFFARX1 I_8716 (I151763,I3563,I151539,I151528,);
nand I_8717 (I151785,I1052281,I1052290);
and I_8718 (I151802,I151785,I1052284);
DFFARX1 I_8719 (I151802,I3563,I151539,I151828,);
DFFARX1 I_8720 (I151828,I3563,I151539,I151845,);
not I_8721 (I151531,I151845);
not I_8722 (I151867,I151828);
nand I_8723 (I151516,I151867,I151706);
nor I_8724 (I151898,I1052287,I1052290);
not I_8725 (I151915,I151898);
nor I_8726 (I151932,I151867,I151915);
nor I_8727 (I151949,I151573,I151932);
DFFARX1 I_8728 (I151949,I3563,I151539,I151525,);
nor I_8729 (I151980,I151633,I151915);
nor I_8730 (I151513,I151828,I151980);
nor I_8731 (I151522,I151763,I151898);
nor I_8732 (I151510,I151633,I151898);
not I_8733 (I152066,I3570);
DFFARX1 I_8734 (I201210,I3563,I152066,I152092,);
not I_8735 (I152100,I152092);
nand I_8736 (I152117,I201204,I201198);
and I_8737 (I152134,I152117,I201219);
DFFARX1 I_8738 (I152134,I3563,I152066,I152160,);
DFFARX1 I_8739 (I201216,I3563,I152066,I152177,);
and I_8740 (I152185,I152177,I201213);
nor I_8741 (I152202,I152160,I152185);
DFFARX1 I_8742 (I152202,I3563,I152066,I152034,);
nand I_8743 (I152233,I152177,I201213);
nand I_8744 (I152250,I152100,I152233);
not I_8745 (I152046,I152250);
DFFARX1 I_8746 (I201198,I3563,I152066,I152290,);
DFFARX1 I_8747 (I152290,I3563,I152066,I152055,);
nand I_8748 (I152312,I201201,I201201);
and I_8749 (I152329,I152312,I201222);
DFFARX1 I_8750 (I152329,I3563,I152066,I152355,);
DFFARX1 I_8751 (I152355,I3563,I152066,I152372,);
not I_8752 (I152058,I152372);
not I_8753 (I152394,I152355);
nand I_8754 (I152043,I152394,I152233);
nor I_8755 (I152425,I201207,I201201);
not I_8756 (I152442,I152425);
nor I_8757 (I152459,I152394,I152442);
nor I_8758 (I152476,I152100,I152459);
DFFARX1 I_8759 (I152476,I3563,I152066,I152052,);
nor I_8760 (I152507,I152160,I152442);
nor I_8761 (I152040,I152355,I152507);
nor I_8762 (I152049,I152290,I152425);
nor I_8763 (I152037,I152160,I152425);
not I_8764 (I152593,I3570);
DFFARX1 I_8765 (I1206601,I3563,I152593,I152619,);
not I_8766 (I152627,I152619);
nand I_8767 (I152644,I1206616,I1206595);
and I_8768 (I152661,I152644,I1206598);
DFFARX1 I_8769 (I152661,I3563,I152593,I152687,);
DFFARX1 I_8770 (I1206619,I3563,I152593,I152704,);
and I_8771 (I152712,I152704,I1206598);
nor I_8772 (I152729,I152687,I152712);
DFFARX1 I_8773 (I152729,I3563,I152593,I152561,);
nand I_8774 (I152760,I152704,I1206598);
nand I_8775 (I152777,I152627,I152760);
not I_8776 (I152573,I152777);
DFFARX1 I_8777 (I1206595,I3563,I152593,I152817,);
DFFARX1 I_8778 (I152817,I3563,I152593,I152582,);
nand I_8779 (I152839,I1206607,I1206604);
and I_8780 (I152856,I152839,I1206610);
DFFARX1 I_8781 (I152856,I3563,I152593,I152882,);
DFFARX1 I_8782 (I152882,I3563,I152593,I152899,);
not I_8783 (I152585,I152899);
not I_8784 (I152921,I152882);
nand I_8785 (I152570,I152921,I152760);
nor I_8786 (I152952,I1206613,I1206604);
not I_8787 (I152969,I152952);
nor I_8788 (I152986,I152921,I152969);
nor I_8789 (I153003,I152627,I152986);
DFFARX1 I_8790 (I153003,I3563,I152593,I152579,);
nor I_8791 (I153034,I152687,I152969);
nor I_8792 (I152567,I152882,I153034);
nor I_8793 (I152576,I152817,I152952);
nor I_8794 (I152564,I152687,I152952);
not I_8795 (I153120,I3570);
DFFARX1 I_8796 (I711601,I3563,I153120,I153146,);
not I_8797 (I153154,I153146);
nand I_8798 (I153171,I711592,I711610);
and I_8799 (I153188,I153171,I711589);
DFFARX1 I_8800 (I153188,I3563,I153120,I153214,);
DFFARX1 I_8801 (I711592,I3563,I153120,I153231,);
and I_8802 (I153239,I153231,I711595);
nor I_8803 (I153256,I153214,I153239);
DFFARX1 I_8804 (I153256,I3563,I153120,I153088,);
nand I_8805 (I153287,I153231,I711595);
nand I_8806 (I153304,I153154,I153287);
not I_8807 (I153100,I153304);
DFFARX1 I_8808 (I711589,I3563,I153120,I153344,);
DFFARX1 I_8809 (I153344,I3563,I153120,I153109,);
nand I_8810 (I153366,I711607,I711598);
and I_8811 (I153383,I153366,I711613);
DFFARX1 I_8812 (I153383,I3563,I153120,I153409,);
DFFARX1 I_8813 (I153409,I3563,I153120,I153426,);
not I_8814 (I153112,I153426);
not I_8815 (I153448,I153409);
nand I_8816 (I153097,I153448,I153287);
nor I_8817 (I153479,I711604,I711598);
not I_8818 (I153496,I153479);
nor I_8819 (I153513,I153448,I153496);
nor I_8820 (I153530,I153154,I153513);
DFFARX1 I_8821 (I153530,I3563,I153120,I153106,);
nor I_8822 (I153561,I153214,I153496);
nor I_8823 (I153094,I153409,I153561);
nor I_8824 (I153103,I153344,I153479);
nor I_8825 (I153091,I153214,I153479);
not I_8826 (I153647,I3570);
DFFARX1 I_8827 (I272610,I3563,I153647,I153673,);
not I_8828 (I153681,I153673);
nand I_8829 (I153698,I272604,I272598);
and I_8830 (I153715,I153698,I272619);
DFFARX1 I_8831 (I153715,I3563,I153647,I153741,);
DFFARX1 I_8832 (I272616,I3563,I153647,I153758,);
and I_8833 (I153766,I153758,I272613);
nor I_8834 (I153783,I153741,I153766);
DFFARX1 I_8835 (I153783,I3563,I153647,I153615,);
nand I_8836 (I153814,I153758,I272613);
nand I_8837 (I153831,I153681,I153814);
not I_8838 (I153627,I153831);
DFFARX1 I_8839 (I272598,I3563,I153647,I153871,);
DFFARX1 I_8840 (I153871,I3563,I153647,I153636,);
nand I_8841 (I153893,I272601,I272601);
and I_8842 (I153910,I153893,I272622);
DFFARX1 I_8843 (I153910,I3563,I153647,I153936,);
DFFARX1 I_8844 (I153936,I3563,I153647,I153953,);
not I_8845 (I153639,I153953);
not I_8846 (I153975,I153936);
nand I_8847 (I153624,I153975,I153814);
nor I_8848 (I154006,I272607,I272601);
not I_8849 (I154023,I154006);
nor I_8850 (I154040,I153975,I154023);
nor I_8851 (I154057,I153681,I154040);
DFFARX1 I_8852 (I154057,I3563,I153647,I153633,);
nor I_8853 (I154088,I153741,I154023);
nor I_8854 (I153621,I153936,I154088);
nor I_8855 (I153630,I153871,I154006);
nor I_8856 (I153618,I153741,I154006);
not I_8857 (I154174,I3570);
DFFARX1 I_8858 (I327552,I3563,I154174,I154200,);
not I_8859 (I154208,I154200);
nand I_8860 (I154225,I327534,I327549);
and I_8861 (I154242,I154225,I327525);
DFFARX1 I_8862 (I154242,I3563,I154174,I154268,);
DFFARX1 I_8863 (I327528,I3563,I154174,I154285,);
and I_8864 (I154293,I154285,I327543);
nor I_8865 (I154310,I154268,I154293);
DFFARX1 I_8866 (I154310,I3563,I154174,I154142,);
nand I_8867 (I154341,I154285,I327543);
nand I_8868 (I154358,I154208,I154341);
not I_8869 (I154154,I154358);
DFFARX1 I_8870 (I327546,I3563,I154174,I154398,);
DFFARX1 I_8871 (I154398,I3563,I154174,I154163,);
nand I_8872 (I154420,I327525,I327537);
and I_8873 (I154437,I154420,I327531);
DFFARX1 I_8874 (I154437,I3563,I154174,I154463,);
DFFARX1 I_8875 (I154463,I3563,I154174,I154480,);
not I_8876 (I154166,I154480);
not I_8877 (I154502,I154463);
nand I_8878 (I154151,I154502,I154341);
nor I_8879 (I154533,I327540,I327537);
not I_8880 (I154550,I154533);
nor I_8881 (I154567,I154502,I154550);
nor I_8882 (I154584,I154208,I154567);
DFFARX1 I_8883 (I154584,I3563,I154174,I154160,);
nor I_8884 (I154615,I154268,I154550);
nor I_8885 (I154148,I154463,I154615);
nor I_8886 (I154157,I154398,I154533);
nor I_8887 (I154145,I154268,I154533);
not I_8888 (I154701,I3570);
DFFARX1 I_8889 (I379198,I3563,I154701,I154727,);
not I_8890 (I154735,I154727);
nand I_8891 (I154752,I379180,I379195);
and I_8892 (I154769,I154752,I379171);
DFFARX1 I_8893 (I154769,I3563,I154701,I154795,);
DFFARX1 I_8894 (I379174,I3563,I154701,I154812,);
and I_8895 (I154820,I154812,I379189);
nor I_8896 (I154837,I154795,I154820);
DFFARX1 I_8897 (I154837,I3563,I154701,I154669,);
nand I_8898 (I154868,I154812,I379189);
nand I_8899 (I154885,I154735,I154868);
not I_8900 (I154681,I154885);
DFFARX1 I_8901 (I379192,I3563,I154701,I154925,);
DFFARX1 I_8902 (I154925,I3563,I154701,I154690,);
nand I_8903 (I154947,I379171,I379183);
and I_8904 (I154964,I154947,I379177);
DFFARX1 I_8905 (I154964,I3563,I154701,I154990,);
DFFARX1 I_8906 (I154990,I3563,I154701,I155007,);
not I_8907 (I154693,I155007);
not I_8908 (I155029,I154990);
nand I_8909 (I154678,I155029,I154868);
nor I_8910 (I155060,I379186,I379183);
not I_8911 (I155077,I155060);
nor I_8912 (I155094,I155029,I155077);
nor I_8913 (I155111,I154735,I155094);
DFFARX1 I_8914 (I155111,I3563,I154701,I154687,);
nor I_8915 (I155142,I154795,I155077);
nor I_8916 (I154675,I154990,I155142);
nor I_8917 (I154684,I154925,I155060);
nor I_8918 (I154672,I154795,I155060);
not I_8919 (I155228,I3570);
DFFARX1 I_8920 (I1360100,I3563,I155228,I155254,);
not I_8921 (I155262,I155254);
nand I_8922 (I155279,I1360094,I1360115);
and I_8923 (I155296,I155279,I1360091);
DFFARX1 I_8924 (I155296,I3563,I155228,I155322,);
DFFARX1 I_8925 (I1360112,I3563,I155228,I155339,);
and I_8926 (I155347,I155339,I1360109);
nor I_8927 (I155364,I155322,I155347);
DFFARX1 I_8928 (I155364,I3563,I155228,I155196,);
nand I_8929 (I155395,I155339,I1360109);
nand I_8930 (I155412,I155262,I155395);
not I_8931 (I155208,I155412);
DFFARX1 I_8932 (I1360097,I3563,I155228,I155452,);
DFFARX1 I_8933 (I155452,I3563,I155228,I155217,);
nand I_8934 (I155474,I1360106,I1360103);
and I_8935 (I155491,I155474,I1360088);
DFFARX1 I_8936 (I155491,I3563,I155228,I155517,);
DFFARX1 I_8937 (I155517,I3563,I155228,I155534,);
not I_8938 (I155220,I155534);
not I_8939 (I155556,I155517);
nand I_8940 (I155205,I155556,I155395);
nor I_8941 (I155587,I1360088,I1360103);
not I_8942 (I155604,I155587);
nor I_8943 (I155621,I155556,I155604);
nor I_8944 (I155638,I155262,I155621);
DFFARX1 I_8945 (I155638,I3563,I155228,I155214,);
nor I_8946 (I155669,I155322,I155604);
nor I_8947 (I155202,I155517,I155669);
nor I_8948 (I155211,I155452,I155587);
nor I_8949 (I155199,I155322,I155587);
not I_8950 (I155755,I3570);
DFFARX1 I_8951 (I1130305,I3563,I155755,I155781,);
not I_8952 (I155789,I155781);
nand I_8953 (I155806,I1130320,I1130299);
and I_8954 (I155823,I155806,I1130302);
DFFARX1 I_8955 (I155823,I3563,I155755,I155849,);
DFFARX1 I_8956 (I1130323,I3563,I155755,I155866,);
and I_8957 (I155874,I155866,I1130302);
nor I_8958 (I155891,I155849,I155874);
DFFARX1 I_8959 (I155891,I3563,I155755,I155723,);
nand I_8960 (I155922,I155866,I1130302);
nand I_8961 (I155939,I155789,I155922);
not I_8962 (I155735,I155939);
DFFARX1 I_8963 (I1130299,I3563,I155755,I155979,);
DFFARX1 I_8964 (I155979,I3563,I155755,I155744,);
nand I_8965 (I156001,I1130311,I1130308);
and I_8966 (I156018,I156001,I1130314);
DFFARX1 I_8967 (I156018,I3563,I155755,I156044,);
DFFARX1 I_8968 (I156044,I3563,I155755,I156061,);
not I_8969 (I155747,I156061);
not I_8970 (I156083,I156044);
nand I_8971 (I155732,I156083,I155922);
nor I_8972 (I156114,I1130317,I1130308);
not I_8973 (I156131,I156114);
nor I_8974 (I156148,I156083,I156131);
nor I_8975 (I156165,I155789,I156148);
DFFARX1 I_8976 (I156165,I3563,I155755,I155741,);
nor I_8977 (I156196,I155849,I156131);
nor I_8978 (I155729,I156044,I156196);
nor I_8979 (I155738,I155979,I156114);
nor I_8980 (I155726,I155849,I156114);
not I_8981 (I156282,I3570);
DFFARX1 I_8982 (I985298,I3563,I156282,I156308,);
not I_8983 (I156316,I156308);
nand I_8984 (I156333,I985316,I985310);
and I_8985 (I156350,I156333,I985289);
DFFARX1 I_8986 (I156350,I3563,I156282,I156376,);
DFFARX1 I_8987 (I985307,I3563,I156282,I156393,);
and I_8988 (I156401,I156393,I985292);
nor I_8989 (I156418,I156376,I156401);
DFFARX1 I_8990 (I156418,I3563,I156282,I156250,);
nand I_8991 (I156449,I156393,I985292);
nand I_8992 (I156466,I156316,I156449);
not I_8993 (I156262,I156466);
DFFARX1 I_8994 (I985304,I3563,I156282,I156506,);
DFFARX1 I_8995 (I156506,I3563,I156282,I156271,);
nand I_8996 (I156528,I985313,I985301);
and I_8997 (I156545,I156528,I985295);
DFFARX1 I_8998 (I156545,I3563,I156282,I156571,);
DFFARX1 I_8999 (I156571,I3563,I156282,I156588,);
not I_9000 (I156274,I156588);
not I_9001 (I156610,I156571);
nand I_9002 (I156259,I156610,I156449);
nor I_9003 (I156641,I985289,I985301);
not I_9004 (I156658,I156641);
nor I_9005 (I156675,I156610,I156658);
nor I_9006 (I156692,I156316,I156675);
DFFARX1 I_9007 (I156692,I3563,I156282,I156268,);
nor I_9008 (I156723,I156376,I156658);
nor I_9009 (I156256,I156571,I156723);
nor I_9010 (I156265,I156506,I156641);
nor I_9011 (I156253,I156376,I156641);
not I_9012 (I156809,I3570);
DFFARX1 I_9013 (I1089298,I3563,I156809,I156835,);
not I_9014 (I156843,I156835);
nand I_9015 (I156860,I1089295,I1089301);
and I_9016 (I156877,I156860,I1089298);
DFFARX1 I_9017 (I156877,I3563,I156809,I156903,);
DFFARX1 I_9018 (I1089301,I3563,I156809,I156920,);
and I_9019 (I156928,I156920,I1089295);
nor I_9020 (I156945,I156903,I156928);
DFFARX1 I_9021 (I156945,I3563,I156809,I156777,);
nand I_9022 (I156976,I156920,I1089295);
nand I_9023 (I156993,I156843,I156976);
not I_9024 (I156789,I156993);
DFFARX1 I_9025 (I1089304,I3563,I156809,I157033,);
DFFARX1 I_9026 (I157033,I3563,I156809,I156798,);
nand I_9027 (I157055,I1089307,I1089316);
and I_9028 (I157072,I157055,I1089310);
DFFARX1 I_9029 (I157072,I3563,I156809,I157098,);
DFFARX1 I_9030 (I157098,I3563,I156809,I157115,);
not I_9031 (I156801,I157115);
not I_9032 (I157137,I157098);
nand I_9033 (I156786,I157137,I156976);
nor I_9034 (I157168,I1089313,I1089316);
not I_9035 (I157185,I157168);
nor I_9036 (I157202,I157137,I157185);
nor I_9037 (I157219,I156843,I157202);
DFFARX1 I_9038 (I157219,I3563,I156809,I156795,);
nor I_9039 (I157250,I156903,I157185);
nor I_9040 (I156783,I157098,I157250);
nor I_9041 (I156792,I157033,I157168);
nor I_9042 (I156780,I156903,I157168);
not I_9043 (I157336,I3570);
DFFARX1 I_9044 (I1293554,I3563,I157336,I157362,);
not I_9045 (I157370,I157362);
nand I_9046 (I157387,I1293557,I1293551);
and I_9047 (I157404,I157387,I1293548);
DFFARX1 I_9048 (I157404,I3563,I157336,I157430,);
DFFARX1 I_9049 (I1293533,I3563,I157336,I157447,);
and I_9050 (I157455,I157447,I1293542);
nor I_9051 (I157472,I157430,I157455);
DFFARX1 I_9052 (I157472,I3563,I157336,I157304,);
nand I_9053 (I157503,I157447,I1293542);
nand I_9054 (I157520,I157370,I157503);
not I_9055 (I157316,I157520);
DFFARX1 I_9056 (I1293533,I3563,I157336,I157560,);
DFFARX1 I_9057 (I157560,I3563,I157336,I157325,);
nand I_9058 (I157582,I1293536,I1293539);
and I_9059 (I157599,I157582,I1293545);
DFFARX1 I_9060 (I157599,I3563,I157336,I157625,);
DFFARX1 I_9061 (I157625,I3563,I157336,I157642,);
not I_9062 (I157328,I157642);
not I_9063 (I157664,I157625);
nand I_9064 (I157313,I157664,I157503);
nor I_9065 (I157695,I1293536,I1293539);
not I_9066 (I157712,I157695);
nor I_9067 (I157729,I157664,I157712);
nor I_9068 (I157746,I157370,I157729);
DFFARX1 I_9069 (I157746,I3563,I157336,I157322,);
nor I_9070 (I157777,I157430,I157712);
nor I_9071 (I157310,I157625,I157777);
nor I_9072 (I157319,I157560,I157695);
nor I_9073 (I157307,I157430,I157695);
not I_9074 (I157863,I3570);
DFFARX1 I_9075 (I228580,I3563,I157863,I157889,);
not I_9076 (I157897,I157889);
nand I_9077 (I157914,I228574,I228568);
and I_9078 (I157931,I157914,I228589);
DFFARX1 I_9079 (I157931,I3563,I157863,I157957,);
DFFARX1 I_9080 (I228586,I3563,I157863,I157974,);
and I_9081 (I157982,I157974,I228583);
nor I_9082 (I157999,I157957,I157982);
DFFARX1 I_9083 (I157999,I3563,I157863,I157831,);
nand I_9084 (I158030,I157974,I228583);
nand I_9085 (I158047,I157897,I158030);
not I_9086 (I157843,I158047);
DFFARX1 I_9087 (I228568,I3563,I157863,I158087,);
DFFARX1 I_9088 (I158087,I3563,I157863,I157852,);
nand I_9089 (I158109,I228571,I228571);
and I_9090 (I158126,I158109,I228592);
DFFARX1 I_9091 (I158126,I3563,I157863,I158152,);
DFFARX1 I_9092 (I158152,I3563,I157863,I158169,);
not I_9093 (I157855,I158169);
not I_9094 (I158191,I158152);
nand I_9095 (I157840,I158191,I158030);
nor I_9096 (I158222,I228577,I228571);
not I_9097 (I158239,I158222);
nor I_9098 (I158256,I158191,I158239);
nor I_9099 (I158273,I157897,I158256);
DFFARX1 I_9100 (I158273,I3563,I157863,I157849,);
nor I_9101 (I158304,I157957,I158239);
nor I_9102 (I157837,I158152,I158304);
nor I_9103 (I157846,I158087,I158222);
nor I_9104 (I157834,I157957,I158222);
not I_9105 (I158393,I3570);
DFFARX1 I_9106 (I1264364,I3563,I158393,I158419,);
not I_9107 (I158427,I158419);
DFFARX1 I_9108 (I1264376,I3563,I158393,I158453,);
not I_9109 (I158461,I1264382);
or I_9110 (I158478,I1264361,I1264382);
nor I_9111 (I158495,I158453,I1264361);
nand I_9112 (I158370,I158461,I158495);
nor I_9113 (I158526,I1264379,I1264361);
nand I_9114 (I158364,I158526,I158461);
not I_9115 (I158557,I1264364);
nand I_9116 (I158574,I158461,I158557);
nor I_9117 (I158591,I1264367,I1264361);
not I_9118 (I158608,I158591);
nor I_9119 (I158625,I158608,I158574);
nor I_9120 (I158642,I158526,I158625);
DFFARX1 I_9121 (I158642,I3563,I158393,I158379,);
nor I_9122 (I158376,I158591,I158478);
DFFARX1 I_9123 (I158591,I3563,I158393,I158382,);
nor I_9124 (I158701,I158557,I1264367);
nor I_9125 (I158718,I158701,I1264382);
nor I_9126 (I158735,I1264385,I1264373);
DFFARX1 I_9127 (I158735,I3563,I158393,I158761,);
nor I_9128 (I158361,I158761,I158718);
DFFARX1 I_9129 (I158761,I3563,I158393,I158792,);
nand I_9130 (I158800,I158792,I1264370);
nor I_9131 (I158385,I158427,I158800);
not I_9132 (I158831,I158761);
nand I_9133 (I158848,I158831,I1264370);
nor I_9134 (I158865,I158427,I158848);
nor I_9135 (I158367,I158453,I158865);
nor I_9136 (I158896,I1264385,I1264379);
nor I_9137 (I158913,I158453,I158896);
DFFARX1 I_9138 (I158913,I3563,I158393,I158358,);
and I_9139 (I158373,I158526,I1264385);
not I_9140 (I158988,I3570);
DFFARX1 I_9141 (I2532,I3563,I158988,I159014,);
not I_9142 (I159022,I159014);
DFFARX1 I_9143 (I2988,I3563,I158988,I159048,);
not I_9144 (I159056,I2652);
or I_9145 (I159073,I3556,I2652);
nor I_9146 (I159090,I159048,I3556);
nand I_9147 (I158965,I159056,I159090);
nor I_9148 (I159121,I2244,I3556);
nand I_9149 (I158959,I159121,I159056);
not I_9150 (I159152,I2284);
nand I_9151 (I159169,I159056,I159152);
nor I_9152 (I159186,I2964,I2468);
not I_9153 (I159203,I159186);
nor I_9154 (I159220,I159203,I159169);
nor I_9155 (I159237,I159121,I159220);
DFFARX1 I_9156 (I159237,I3563,I158988,I158974,);
nor I_9157 (I158971,I159186,I159073);
DFFARX1 I_9158 (I159186,I3563,I158988,I158977,);
nor I_9159 (I159296,I159152,I2964);
nor I_9160 (I159313,I159296,I2652);
nor I_9161 (I159330,I2292,I2892);
DFFARX1 I_9162 (I159330,I3563,I158988,I159356,);
nor I_9163 (I158956,I159356,I159313);
DFFARX1 I_9164 (I159356,I3563,I158988,I159387,);
nand I_9165 (I159395,I159387,I1908);
nor I_9166 (I158980,I159022,I159395);
not I_9167 (I159426,I159356);
nand I_9168 (I159443,I159426,I1908);
nor I_9169 (I159460,I159022,I159443);
nor I_9170 (I158962,I159048,I159460);
nor I_9171 (I159491,I2292,I2244);
nor I_9172 (I159508,I159048,I159491);
DFFARX1 I_9173 (I159508,I3563,I158988,I158953,);
and I_9174 (I158968,I159121,I2292);
not I_9175 (I159583,I3570);
DFFARX1 I_9176 (I394990,I3563,I159583,I159609,);
not I_9177 (I159617,I159609);
DFFARX1 I_9178 (I394987,I3563,I159583,I159643,);
not I_9179 (I159651,I394984);
or I_9180 (I159668,I394996,I394984);
nor I_9181 (I159685,I159643,I394996);
nand I_9182 (I159560,I159651,I159685);
nor I_9183 (I159716,I395005,I394996);
nand I_9184 (I159554,I159716,I159651);
not I_9185 (I159747,I395002);
nand I_9186 (I159764,I159651,I159747);
nor I_9187 (I159781,I394981,I394981);
not I_9188 (I159798,I159781);
nor I_9189 (I159815,I159798,I159764);
nor I_9190 (I159832,I159716,I159815);
DFFARX1 I_9191 (I159832,I3563,I159583,I159569,);
nor I_9192 (I159566,I159781,I159668);
DFFARX1 I_9193 (I159781,I3563,I159583,I159572,);
nor I_9194 (I159891,I159747,I394981);
nor I_9195 (I159908,I159891,I394984);
nor I_9196 (I159925,I394993,I395008);
DFFARX1 I_9197 (I159925,I3563,I159583,I159951,);
nor I_9198 (I159551,I159951,I159908);
DFFARX1 I_9199 (I159951,I3563,I159583,I159982,);
nand I_9200 (I159990,I159982,I394999);
nor I_9201 (I159575,I159617,I159990);
not I_9202 (I160021,I159951);
nand I_9203 (I160038,I160021,I394999);
nor I_9204 (I160055,I159617,I160038);
nor I_9205 (I159557,I159643,I160055);
nor I_9206 (I160086,I394993,I395005);
nor I_9207 (I160103,I159643,I160086);
DFFARX1 I_9208 (I160103,I3563,I159583,I159548,);
and I_9209 (I159563,I159716,I394993);
not I_9210 (I160178,I3570);
DFFARX1 I_9211 (I520890,I3563,I160178,I160204,);
not I_9212 (I160212,I160204);
DFFARX1 I_9213 (I520884,I3563,I160178,I160238,);
not I_9214 (I160246,I520881);
or I_9215 (I160263,I520872,I520881);
nor I_9216 (I160280,I160238,I520872);
nand I_9217 (I160155,I160246,I160280);
nor I_9218 (I160311,I520875,I520872);
nand I_9219 (I160149,I160311,I160246);
not I_9220 (I160342,I520878);
nand I_9221 (I160359,I160246,I160342);
nor I_9222 (I160376,I520866,I520893);
not I_9223 (I160393,I160376);
nor I_9224 (I160410,I160393,I160359);
nor I_9225 (I160427,I160311,I160410);
DFFARX1 I_9226 (I160427,I3563,I160178,I160164,);
nor I_9227 (I160161,I160376,I160263);
DFFARX1 I_9228 (I160376,I3563,I160178,I160167,);
nor I_9229 (I160486,I160342,I520866);
nor I_9230 (I160503,I160486,I520881);
nor I_9231 (I160520,I520869,I520866);
DFFARX1 I_9232 (I160520,I3563,I160178,I160546,);
nor I_9233 (I160146,I160546,I160503);
DFFARX1 I_9234 (I160546,I3563,I160178,I160577,);
nand I_9235 (I160585,I160577,I520887);
nor I_9236 (I160170,I160212,I160585);
not I_9237 (I160616,I160546);
nand I_9238 (I160633,I160616,I520887);
nor I_9239 (I160650,I160212,I160633);
nor I_9240 (I160152,I160238,I160650);
nor I_9241 (I160681,I520869,I520875);
nor I_9242 (I160698,I160238,I160681);
DFFARX1 I_9243 (I160698,I3563,I160178,I160143,);
and I_9244 (I160158,I160311,I520869);
not I_9245 (I160773,I3570);
DFFARX1 I_9246 (I129921,I3563,I160773,I160799,);
not I_9247 (I160807,I160799);
DFFARX1 I_9248 (I129915,I3563,I160773,I160833,);
not I_9249 (I160841,I129924);
or I_9250 (I160858,I129909,I129924);
nor I_9251 (I160875,I160833,I129909);
nand I_9252 (I160750,I160841,I160875);
nor I_9253 (I160906,I129900,I129909);
nand I_9254 (I160744,I160906,I160841);
not I_9255 (I160937,I129900);
nand I_9256 (I160954,I160841,I160937);
nor I_9257 (I160971,I129903,I129918);
not I_9258 (I160988,I160971);
nor I_9259 (I161005,I160988,I160954);
nor I_9260 (I161022,I160906,I161005);
DFFARX1 I_9261 (I161022,I3563,I160773,I160759,);
nor I_9262 (I160756,I160971,I160858);
DFFARX1 I_9263 (I160971,I3563,I160773,I160762,);
nor I_9264 (I161081,I160937,I129903);
nor I_9265 (I161098,I161081,I129924);
nor I_9266 (I161115,I129903,I129912);
DFFARX1 I_9267 (I161115,I3563,I160773,I161141,);
nor I_9268 (I160741,I161141,I161098);
DFFARX1 I_9269 (I161141,I3563,I160773,I161172,);
nand I_9270 (I161180,I161172,I129906);
nor I_9271 (I160765,I160807,I161180);
not I_9272 (I161211,I161141);
nand I_9273 (I161228,I161211,I129906);
nor I_9274 (I161245,I160807,I161228);
nor I_9275 (I160747,I160833,I161245);
nor I_9276 (I161276,I129903,I129900);
nor I_9277 (I161293,I160833,I161276);
DFFARX1 I_9278 (I161293,I3563,I160773,I160738,);
and I_9279 (I160753,I160906,I129903);
not I_9280 (I161368,I3570);
DFFARX1 I_9281 (I1277964,I3563,I161368,I161394,);
not I_9282 (I161402,I161394);
DFFARX1 I_9283 (I1277976,I3563,I161368,I161428,);
not I_9284 (I161436,I1277982);
or I_9285 (I161453,I1277961,I1277982);
nor I_9286 (I161470,I161428,I1277961);
nand I_9287 (I161345,I161436,I161470);
nor I_9288 (I161501,I1277979,I1277961);
nand I_9289 (I161339,I161501,I161436);
not I_9290 (I161532,I1277964);
nand I_9291 (I161549,I161436,I161532);
nor I_9292 (I161566,I1277967,I1277961);
not I_9293 (I161583,I161566);
nor I_9294 (I161600,I161583,I161549);
nor I_9295 (I161617,I161501,I161600);
DFFARX1 I_9296 (I161617,I3563,I161368,I161354,);
nor I_9297 (I161351,I161566,I161453);
DFFARX1 I_9298 (I161566,I3563,I161368,I161357,);
nor I_9299 (I161676,I161532,I1277967);
nor I_9300 (I161693,I161676,I1277982);
nor I_9301 (I161710,I1277985,I1277973);
DFFARX1 I_9302 (I161710,I3563,I161368,I161736,);
nor I_9303 (I161336,I161736,I161693);
DFFARX1 I_9304 (I161736,I3563,I161368,I161767,);
nand I_9305 (I161775,I161767,I1277970);
nor I_9306 (I161360,I161402,I161775);
not I_9307 (I161806,I161736);
nand I_9308 (I161823,I161806,I1277970);
nor I_9309 (I161840,I161402,I161823);
nor I_9310 (I161342,I161428,I161840);
nor I_9311 (I161871,I1277985,I1277979);
nor I_9312 (I161888,I161428,I161871);
DFFARX1 I_9313 (I161888,I3563,I161368,I161333,);
and I_9314 (I161348,I161501,I1277985);
not I_9315 (I161963,I3570);
DFFARX1 I_9316 (I350195,I3563,I161963,I161989,);
not I_9317 (I161997,I161989);
DFFARX1 I_9318 (I350192,I3563,I161963,I162023,);
not I_9319 (I162031,I350189);
or I_9320 (I162048,I350201,I350189);
nor I_9321 (I162065,I162023,I350201);
nand I_9322 (I161940,I162031,I162065);
nor I_9323 (I162096,I350210,I350201);
nand I_9324 (I161934,I162096,I162031);
not I_9325 (I162127,I350207);
nand I_9326 (I162144,I162031,I162127);
nor I_9327 (I162161,I350186,I350186);
not I_9328 (I162178,I162161);
nor I_9329 (I162195,I162178,I162144);
nor I_9330 (I162212,I162096,I162195);
DFFARX1 I_9331 (I162212,I3563,I161963,I161949,);
nor I_9332 (I161946,I162161,I162048);
DFFARX1 I_9333 (I162161,I3563,I161963,I161952,);
nor I_9334 (I162271,I162127,I350186);
nor I_9335 (I162288,I162271,I350189);
nor I_9336 (I162305,I350198,I350213);
DFFARX1 I_9337 (I162305,I3563,I161963,I162331,);
nor I_9338 (I161931,I162331,I162288);
DFFARX1 I_9339 (I162331,I3563,I161963,I162362,);
nand I_9340 (I162370,I162362,I350204);
nor I_9341 (I161955,I161997,I162370);
not I_9342 (I162401,I162331);
nand I_9343 (I162418,I162401,I350204);
nor I_9344 (I162435,I161997,I162418);
nor I_9345 (I161937,I162023,I162435);
nor I_9346 (I162466,I350198,I350210);
nor I_9347 (I162483,I162023,I162466);
DFFARX1 I_9348 (I162483,I3563,I161963,I161928,);
and I_9349 (I161943,I162096,I350198);
not I_9350 (I162558,I3570);
DFFARX1 I_9351 (I411327,I3563,I162558,I162584,);
not I_9352 (I162592,I162584);
DFFARX1 I_9353 (I411324,I3563,I162558,I162618,);
not I_9354 (I162626,I411321);
or I_9355 (I162643,I411333,I411321);
nor I_9356 (I162660,I162618,I411333);
nand I_9357 (I162535,I162626,I162660);
nor I_9358 (I162691,I411342,I411333);
nand I_9359 (I162529,I162691,I162626);
not I_9360 (I162722,I411339);
nand I_9361 (I162739,I162626,I162722);
nor I_9362 (I162756,I411318,I411318);
not I_9363 (I162773,I162756);
nor I_9364 (I162790,I162773,I162739);
nor I_9365 (I162807,I162691,I162790);
DFFARX1 I_9366 (I162807,I3563,I162558,I162544,);
nor I_9367 (I162541,I162756,I162643);
DFFARX1 I_9368 (I162756,I3563,I162558,I162547,);
nor I_9369 (I162866,I162722,I411318);
nor I_9370 (I162883,I162866,I411321);
nor I_9371 (I162900,I411330,I411345);
DFFARX1 I_9372 (I162900,I3563,I162558,I162926,);
nor I_9373 (I162526,I162926,I162883);
DFFARX1 I_9374 (I162926,I3563,I162558,I162957,);
nand I_9375 (I162965,I162957,I411336);
nor I_9376 (I162550,I162592,I162965);
not I_9377 (I162996,I162926);
nand I_9378 (I163013,I162996,I411336);
nor I_9379 (I163030,I162592,I163013);
nor I_9380 (I162532,I162618,I163030);
nor I_9381 (I163061,I411330,I411342);
nor I_9382 (I163078,I162618,I163061);
DFFARX1 I_9383 (I163078,I3563,I162558,I162523,);
and I_9384 (I162538,I162691,I411330);
not I_9385 (I163153,I3570);
DFFARX1 I_9386 (I776903,I3563,I163153,I163179,);
not I_9387 (I163187,I163179);
DFFARX1 I_9388 (I776924,I3563,I163153,I163213,);
not I_9389 (I163221,I776903);
or I_9390 (I163238,I776915,I776903);
nor I_9391 (I163255,I163213,I776915);
nand I_9392 (I163130,I163221,I163255);
nor I_9393 (I163286,I776912,I776915);
nand I_9394 (I163124,I163286,I163221);
not I_9395 (I163317,I776921);
nand I_9396 (I163334,I163221,I163317);
nor I_9397 (I163351,I776906,I776906);
not I_9398 (I163368,I163351);
nor I_9399 (I163385,I163368,I163334);
nor I_9400 (I163402,I163286,I163385);
DFFARX1 I_9401 (I163402,I3563,I163153,I163139,);
nor I_9402 (I163136,I163351,I163238);
DFFARX1 I_9403 (I163351,I3563,I163153,I163142,);
nor I_9404 (I163461,I163317,I776906);
nor I_9405 (I163478,I163461,I776903);
nor I_9406 (I163495,I776927,I776909);
DFFARX1 I_9407 (I163495,I3563,I163153,I163521,);
nor I_9408 (I163121,I163521,I163478);
DFFARX1 I_9409 (I163521,I3563,I163153,I163552,);
nand I_9410 (I163560,I163552,I776918);
nor I_9411 (I163145,I163187,I163560);
not I_9412 (I163591,I163521);
nand I_9413 (I163608,I163591,I776918);
nor I_9414 (I163625,I163187,I163608);
nor I_9415 (I163127,I163213,I163625);
nor I_9416 (I163656,I776927,I776912);
nor I_9417 (I163673,I163213,I163656);
DFFARX1 I_9418 (I163673,I3563,I163153,I163118,);
and I_9419 (I163133,I163286,I776927);
not I_9420 (I163748,I3570);
DFFARX1 I_9421 (I1130880,I3563,I163748,I163774,);
not I_9422 (I163782,I163774);
DFFARX1 I_9423 (I1130877,I3563,I163748,I163808,);
not I_9424 (I163816,I1130886);
or I_9425 (I163833,I1130877,I1130886);
nor I_9426 (I163850,I163808,I1130877);
nand I_9427 (I163725,I163816,I163850);
nor I_9428 (I163881,I1130889,I1130877);
nand I_9429 (I163719,I163881,I163816);
not I_9430 (I163912,I1130883);
nand I_9431 (I163929,I163816,I163912);
nor I_9432 (I163946,I1130880,I1130898);
not I_9433 (I163963,I163946);
nor I_9434 (I163980,I163963,I163929);
nor I_9435 (I163997,I163881,I163980);
DFFARX1 I_9436 (I163997,I3563,I163748,I163734,);
nor I_9437 (I163731,I163946,I163833);
DFFARX1 I_9438 (I163946,I3563,I163748,I163737,);
nor I_9439 (I164056,I163912,I1130880);
nor I_9440 (I164073,I164056,I1130886);
nor I_9441 (I164090,I1130901,I1130895);
DFFARX1 I_9442 (I164090,I3563,I163748,I164116,);
nor I_9443 (I163716,I164116,I164073);
DFFARX1 I_9444 (I164116,I3563,I163748,I164147,);
nand I_9445 (I164155,I164147,I1130892);
nor I_9446 (I163740,I163782,I164155);
not I_9447 (I164186,I164116);
nand I_9448 (I164203,I164186,I1130892);
nor I_9449 (I164220,I163782,I164203);
nor I_9450 (I163722,I163808,I164220);
nor I_9451 (I164251,I1130901,I1130889);
nor I_9452 (I164268,I163808,I164251);
DFFARX1 I_9453 (I164268,I3563,I163748,I163713,);
and I_9454 (I163728,I163881,I1130901);
not I_9455 (I164343,I3570);
DFFARX1 I_9456 (I724883,I3563,I164343,I164369,);
not I_9457 (I164377,I164369);
DFFARX1 I_9458 (I724904,I3563,I164343,I164403,);
not I_9459 (I164411,I724883);
or I_9460 (I164428,I724895,I724883);
nor I_9461 (I164445,I164403,I724895);
nand I_9462 (I164320,I164411,I164445);
nor I_9463 (I164476,I724892,I724895);
nand I_9464 (I164314,I164476,I164411);
not I_9465 (I164507,I724901);
nand I_9466 (I164524,I164411,I164507);
nor I_9467 (I164541,I724886,I724886);
not I_9468 (I164558,I164541);
nor I_9469 (I164575,I164558,I164524);
nor I_9470 (I164592,I164476,I164575);
DFFARX1 I_9471 (I164592,I3563,I164343,I164329,);
nor I_9472 (I164326,I164541,I164428);
DFFARX1 I_9473 (I164541,I3563,I164343,I164332,);
nor I_9474 (I164651,I164507,I724886);
nor I_9475 (I164668,I164651,I724883);
nor I_9476 (I164685,I724907,I724889);
DFFARX1 I_9477 (I164685,I3563,I164343,I164711,);
nor I_9478 (I164311,I164711,I164668);
DFFARX1 I_9479 (I164711,I3563,I164343,I164742,);
nand I_9480 (I164750,I164742,I724898);
nor I_9481 (I164335,I164377,I164750);
not I_9482 (I164781,I164711);
nand I_9483 (I164798,I164781,I724898);
nor I_9484 (I164815,I164377,I164798);
nor I_9485 (I164317,I164403,I164815);
nor I_9486 (I164846,I724907,I724892);
nor I_9487 (I164863,I164403,I164846);
DFFARX1 I_9488 (I164863,I3563,I164343,I164308,);
and I_9489 (I164323,I164476,I724907);
not I_9490 (I164938,I3570);
DFFARX1 I_9491 (I1027931,I3563,I164938,I164964,);
not I_9492 (I164972,I164964);
DFFARX1 I_9493 (I1027952,I3563,I164938,I164998,);
not I_9494 (I165006,I1027934);
or I_9495 (I165023,I1027925,I1027934);
nor I_9496 (I165040,I164998,I1027925);
nand I_9497 (I164915,I165006,I165040);
nor I_9498 (I165071,I1027937,I1027925);
nand I_9499 (I164909,I165071,I165006);
not I_9500 (I165102,I1027928);
nand I_9501 (I165119,I165006,I165102);
nor I_9502 (I165136,I1027946,I1027949);
not I_9503 (I165153,I165136);
nor I_9504 (I165170,I165153,I165119);
nor I_9505 (I165187,I165071,I165170);
DFFARX1 I_9506 (I165187,I3563,I164938,I164924,);
nor I_9507 (I164921,I165136,I165023);
DFFARX1 I_9508 (I165136,I3563,I164938,I164927,);
nor I_9509 (I165246,I165102,I1027946);
nor I_9510 (I165263,I165246,I1027934);
nor I_9511 (I165280,I1027940,I1027943);
DFFARX1 I_9512 (I165280,I3563,I164938,I165306,);
nor I_9513 (I164906,I165306,I165263);
DFFARX1 I_9514 (I165306,I3563,I164938,I165337,);
nand I_9515 (I165345,I165337,I1027925);
nor I_9516 (I164930,I164972,I165345);
not I_9517 (I165376,I165306);
nand I_9518 (I165393,I165376,I1027925);
nor I_9519 (I165410,I164972,I165393);
nor I_9520 (I164912,I164998,I165410);
nor I_9521 (I165441,I1027940,I1027937);
nor I_9522 (I165458,I164998,I165441);
DFFARX1 I_9523 (I165458,I3563,I164938,I164903,);
and I_9524 (I164918,I165071,I1027940);
not I_9525 (I165530,I3570);
DFFARX1 I_9526 (I1096775,I3563,I165530,I165556,);
DFFARX1 I_9527 (I165556,I3563,I165530,I165573,);
not I_9528 (I165522,I165573);
not I_9529 (I165595,I165556);
DFFARX1 I_9530 (I1096775,I3563,I165530,I165621,);
not I_9531 (I165629,I165621);
and I_9532 (I165646,I165595,I1096778);
not I_9533 (I165663,I1096790);
nand I_9534 (I165680,I165663,I1096778);
not I_9535 (I165697,I1096796);
nor I_9536 (I165714,I165697,I1096787);
nand I_9537 (I165731,I165714,I1096793);
nor I_9538 (I165748,I165731,I165680);
DFFARX1 I_9539 (I165748,I3563,I165530,I165498,);
not I_9540 (I165779,I165731);
not I_9541 (I165796,I1096787);
nand I_9542 (I165813,I165796,I1096778);
nor I_9543 (I165830,I1096787,I1096790);
nand I_9544 (I165510,I165646,I165830);
nand I_9545 (I165504,I165595,I1096787);
nand I_9546 (I165875,I165697,I1096784);
DFFARX1 I_9547 (I165875,I3563,I165530,I165519,);
DFFARX1 I_9548 (I165875,I3563,I165530,I165513,);
not I_9549 (I165920,I1096784);
nor I_9550 (I165937,I165920,I1096781);
and I_9551 (I165954,I165937,I1096799);
or I_9552 (I165971,I165954,I1096778);
DFFARX1 I_9553 (I165971,I3563,I165530,I165997,);
nand I_9554 (I166005,I165997,I165663);
nor I_9555 (I165507,I166005,I165813);
nor I_9556 (I165501,I165997,I165629);
DFFARX1 I_9557 (I165997,I3563,I165530,I166059,);
not I_9558 (I166067,I166059);
nor I_9559 (I165516,I166067,I165779);
not I_9560 (I166125,I3570);
DFFARX1 I_9561 (I1250235,I3563,I166125,I166151,);
DFFARX1 I_9562 (I166151,I3563,I166125,I166168,);
not I_9563 (I166117,I166168);
not I_9564 (I166190,I166151);
DFFARX1 I_9565 (I1250220,I3563,I166125,I166216,);
not I_9566 (I166224,I166216);
and I_9567 (I166241,I166190,I1250238);
not I_9568 (I166258,I1250220);
nand I_9569 (I166275,I166258,I1250238);
not I_9570 (I166292,I1250241);
nor I_9571 (I166309,I166292,I1250232);
nand I_9572 (I166326,I166309,I1250229);
nor I_9573 (I166343,I166326,I166275);
DFFARX1 I_9574 (I166343,I3563,I166125,I166093,);
not I_9575 (I166374,I166326);
not I_9576 (I166391,I1250232);
nand I_9577 (I166408,I166391,I1250238);
nor I_9578 (I166425,I1250232,I1250220);
nand I_9579 (I166105,I166241,I166425);
nand I_9580 (I166099,I166190,I1250232);
nand I_9581 (I166470,I166292,I1250226);
DFFARX1 I_9582 (I166470,I3563,I166125,I166114,);
DFFARX1 I_9583 (I166470,I3563,I166125,I166108,);
not I_9584 (I166515,I1250226);
nor I_9585 (I166532,I166515,I1250217);
and I_9586 (I166549,I166532,I1250223);
or I_9587 (I166566,I166549,I1250217);
DFFARX1 I_9588 (I166566,I3563,I166125,I166592,);
nand I_9589 (I166600,I166592,I166258);
nor I_9590 (I166102,I166600,I166408);
nor I_9591 (I166096,I166592,I166224);
DFFARX1 I_9592 (I166592,I3563,I166125,I166654,);
not I_9593 (I166662,I166654);
nor I_9594 (I166111,I166662,I166374);
not I_9595 (I166720,I3570);
DFFARX1 I_9596 (I64561,I3563,I166720,I166746,);
DFFARX1 I_9597 (I166746,I3563,I166720,I166763,);
not I_9598 (I166712,I166763);
not I_9599 (I166785,I166746);
DFFARX1 I_9600 (I64555,I3563,I166720,I166811,);
not I_9601 (I166819,I166811);
and I_9602 (I166836,I166785,I64552);
not I_9603 (I166853,I64573);
nand I_9604 (I166870,I166853,I64552);
not I_9605 (I166887,I64567);
nor I_9606 (I166904,I166887,I64558);
nand I_9607 (I166921,I166904,I64564);
nor I_9608 (I166938,I166921,I166870);
DFFARX1 I_9609 (I166938,I3563,I166720,I166688,);
not I_9610 (I166969,I166921);
not I_9611 (I166986,I64558);
nand I_9612 (I167003,I166986,I64552);
nor I_9613 (I167020,I64558,I64573);
nand I_9614 (I166700,I166836,I167020);
nand I_9615 (I166694,I166785,I64558);
nand I_9616 (I167065,I166887,I64552);
DFFARX1 I_9617 (I167065,I3563,I166720,I166709,);
DFFARX1 I_9618 (I167065,I3563,I166720,I166703,);
not I_9619 (I167110,I64552);
nor I_9620 (I167127,I167110,I64570);
and I_9621 (I167144,I167127,I64576);
or I_9622 (I167161,I167144,I64555);
DFFARX1 I_9623 (I167161,I3563,I166720,I167187,);
nand I_9624 (I167195,I167187,I166853);
nor I_9625 (I166697,I167195,I167003);
nor I_9626 (I166691,I167187,I166819);
DFFARX1 I_9627 (I167187,I3563,I166720,I167249,);
not I_9628 (I167257,I167249);
nor I_9629 (I166706,I167257,I166969);
not I_9630 (I167315,I3570);
DFFARX1 I_9631 (I1612,I3563,I167315,I167341,);
DFFARX1 I_9632 (I167341,I3563,I167315,I167358,);
not I_9633 (I167307,I167358);
not I_9634 (I167380,I167341);
DFFARX1 I_9635 (I2228,I3563,I167315,I167406,);
not I_9636 (I167414,I167406);
and I_9637 (I167431,I167380,I3116);
not I_9638 (I167448,I3092);
nand I_9639 (I167465,I167448,I3116);
not I_9640 (I167482,I1660);
nor I_9641 (I167499,I167482,I1644);
nand I_9642 (I167516,I167499,I1372);
nor I_9643 (I167533,I167516,I167465);
DFFARX1 I_9644 (I167533,I3563,I167315,I167283,);
not I_9645 (I167564,I167516);
not I_9646 (I167581,I1644);
nand I_9647 (I167598,I167581,I3116);
nor I_9648 (I167615,I1644,I3092);
nand I_9649 (I167295,I167431,I167615);
nand I_9650 (I167289,I167380,I1644);
nand I_9651 (I167660,I167482,I2572);
DFFARX1 I_9652 (I167660,I3563,I167315,I167304,);
DFFARX1 I_9653 (I167660,I3563,I167315,I167298,);
not I_9654 (I167705,I2572);
nor I_9655 (I167722,I167705,I1548);
and I_9656 (I167739,I167722,I3412);
or I_9657 (I167756,I167739,I1956);
DFFARX1 I_9658 (I167756,I3563,I167315,I167782,);
nand I_9659 (I167790,I167782,I167448);
nor I_9660 (I167292,I167790,I167598);
nor I_9661 (I167286,I167782,I167414);
DFFARX1 I_9662 (I167782,I3563,I167315,I167844,);
not I_9663 (I167852,I167844);
nor I_9664 (I167301,I167852,I167564);
not I_9665 (I167910,I3570);
DFFARX1 I_9666 (I124112,I3563,I167910,I167936,);
DFFARX1 I_9667 (I167936,I3563,I167910,I167953,);
not I_9668 (I167902,I167953);
not I_9669 (I167975,I167936);
DFFARX1 I_9670 (I124106,I3563,I167910,I168001,);
not I_9671 (I168009,I168001);
and I_9672 (I168026,I167975,I124103);
not I_9673 (I168043,I124124);
nand I_9674 (I168060,I168043,I124103);
not I_9675 (I168077,I124118);
nor I_9676 (I168094,I168077,I124109);
nand I_9677 (I168111,I168094,I124115);
nor I_9678 (I168128,I168111,I168060);
DFFARX1 I_9679 (I168128,I3563,I167910,I167878,);
not I_9680 (I168159,I168111);
not I_9681 (I168176,I124109);
nand I_9682 (I168193,I168176,I124103);
nor I_9683 (I168210,I124109,I124124);
nand I_9684 (I167890,I168026,I168210);
nand I_9685 (I167884,I167975,I124109);
nand I_9686 (I168255,I168077,I124103);
DFFARX1 I_9687 (I168255,I3563,I167910,I167899,);
DFFARX1 I_9688 (I168255,I3563,I167910,I167893,);
not I_9689 (I168300,I124103);
nor I_9690 (I168317,I168300,I124121);
and I_9691 (I168334,I168317,I124127);
or I_9692 (I168351,I168334,I124106);
DFFARX1 I_9693 (I168351,I3563,I167910,I168377,);
nand I_9694 (I168385,I168377,I168043);
nor I_9695 (I167887,I168385,I168193);
nor I_9696 (I167881,I168377,I168009);
DFFARX1 I_9697 (I168377,I3563,I167910,I168439,);
not I_9698 (I168447,I168439);
nor I_9699 (I167896,I168447,I168159);
not I_9700 (I168505,I3570);
DFFARX1 I_9701 (I1082005,I3563,I168505,I168531,);
DFFARX1 I_9702 (I168531,I3563,I168505,I168548,);
not I_9703 (I168497,I168548);
not I_9704 (I168570,I168531);
DFFARX1 I_9705 (I1082014,I3563,I168505,I168596,);
not I_9706 (I168604,I168596);
and I_9707 (I168621,I168570,I1082008);
not I_9708 (I168638,I1082002);
nand I_9709 (I168655,I168638,I1082008);
not I_9710 (I168672,I1082017);
nor I_9711 (I168689,I168672,I1082005);
nand I_9712 (I168706,I168689,I1082011);
nor I_9713 (I168723,I168706,I168655);
DFFARX1 I_9714 (I168723,I3563,I168505,I168473,);
not I_9715 (I168754,I168706);
not I_9716 (I168771,I1082005);
nand I_9717 (I168788,I168771,I1082008);
nor I_9718 (I168805,I1082005,I1082002);
nand I_9719 (I168485,I168621,I168805);
nand I_9720 (I168479,I168570,I1082005);
nand I_9721 (I168850,I168672,I1082008);
DFFARX1 I_9722 (I168850,I3563,I168505,I168494,);
DFFARX1 I_9723 (I168850,I3563,I168505,I168488,);
not I_9724 (I168895,I1082008);
nor I_9725 (I168912,I168895,I1082023);
and I_9726 (I168929,I168912,I1082020);
or I_9727 (I168946,I168929,I1082002);
DFFARX1 I_9728 (I168946,I3563,I168505,I168972,);
nand I_9729 (I168980,I168972,I168638);
nor I_9730 (I168482,I168980,I168788);
nor I_9731 (I168476,I168972,I168604);
DFFARX1 I_9732 (I168972,I3563,I168505,I169034,);
not I_9733 (I169042,I169034);
nor I_9734 (I168491,I169042,I168754);
not I_9735 (I169100,I3570);
DFFARX1 I_9736 (I1056199,I3563,I169100,I169126,);
DFFARX1 I_9737 (I169126,I3563,I169100,I169143,);
not I_9738 (I169092,I169143);
not I_9739 (I169165,I169126);
DFFARX1 I_9740 (I1056208,I3563,I169100,I169191,);
not I_9741 (I169199,I169191);
and I_9742 (I169216,I169165,I1056202);
not I_9743 (I169233,I1056196);
nand I_9744 (I169250,I169233,I1056202);
not I_9745 (I169267,I1056211);
nor I_9746 (I169284,I169267,I1056199);
nand I_9747 (I169301,I169284,I1056205);
nor I_9748 (I169318,I169301,I169250);
DFFARX1 I_9749 (I169318,I3563,I169100,I169068,);
not I_9750 (I169349,I169301);
not I_9751 (I169366,I1056199);
nand I_9752 (I169383,I169366,I1056202);
nor I_9753 (I169400,I1056199,I1056196);
nand I_9754 (I169080,I169216,I169400);
nand I_9755 (I169074,I169165,I1056199);
nand I_9756 (I169445,I169267,I1056202);
DFFARX1 I_9757 (I169445,I3563,I169100,I169089,);
DFFARX1 I_9758 (I169445,I3563,I169100,I169083,);
not I_9759 (I169490,I1056202);
nor I_9760 (I169507,I169490,I1056217);
and I_9761 (I169524,I169507,I1056214);
or I_9762 (I169541,I169524,I1056196);
DFFARX1 I_9763 (I169541,I3563,I169100,I169567,);
nand I_9764 (I169575,I169567,I169233);
nor I_9765 (I169077,I169575,I169383);
nor I_9766 (I169071,I169567,I169199);
DFFARX1 I_9767 (I169567,I3563,I169100,I169629,);
not I_9768 (I169637,I169629);
nor I_9769 (I169086,I169637,I169349);
not I_9770 (I169695,I3570);
DFFARX1 I_9771 (I782695,I3563,I169695,I169721,);
DFFARX1 I_9772 (I169721,I3563,I169695,I169738,);
not I_9773 (I169687,I169738);
not I_9774 (I169760,I169721);
DFFARX1 I_9775 (I782692,I3563,I169695,I169786,);
not I_9776 (I169794,I169786);
and I_9777 (I169811,I169760,I782698);
not I_9778 (I169828,I782683);
nand I_9779 (I169845,I169828,I782698);
not I_9780 (I169862,I782686);
nor I_9781 (I169879,I169862,I782707);
nand I_9782 (I169896,I169879,I782704);
nor I_9783 (I169913,I169896,I169845);
DFFARX1 I_9784 (I169913,I3563,I169695,I169663,);
not I_9785 (I169944,I169896);
not I_9786 (I169961,I782707);
nand I_9787 (I169978,I169961,I782698);
nor I_9788 (I169995,I782707,I782683);
nand I_9789 (I169675,I169811,I169995);
nand I_9790 (I169669,I169760,I782707);
nand I_9791 (I170040,I169862,I782683);
DFFARX1 I_9792 (I170040,I3563,I169695,I169684,);
DFFARX1 I_9793 (I170040,I3563,I169695,I169678,);
not I_9794 (I170085,I782683);
nor I_9795 (I170102,I170085,I782689);
and I_9796 (I170119,I170102,I782701);
or I_9797 (I170136,I170119,I782686);
DFFARX1 I_9798 (I170136,I3563,I169695,I170162,);
nand I_9799 (I170170,I170162,I169828);
nor I_9800 (I169672,I170170,I169978);
nor I_9801 (I169666,I170162,I169794);
DFFARX1 I_9802 (I170162,I3563,I169695,I170224,);
not I_9803 (I170232,I170224);
nor I_9804 (I169681,I170232,I169944);
not I_9805 (I170290,I3570);
DFFARX1 I_9806 (I1126831,I3563,I170290,I170316,);
DFFARX1 I_9807 (I170316,I3563,I170290,I170333,);
not I_9808 (I170282,I170333);
not I_9809 (I170355,I170316);
DFFARX1 I_9810 (I1126831,I3563,I170290,I170381,);
not I_9811 (I170389,I170381);
and I_9812 (I170406,I170355,I1126834);
not I_9813 (I170423,I1126846);
nand I_9814 (I170440,I170423,I1126834);
not I_9815 (I170457,I1126852);
nor I_9816 (I170474,I170457,I1126843);
nand I_9817 (I170491,I170474,I1126849);
nor I_9818 (I170508,I170491,I170440);
DFFARX1 I_9819 (I170508,I3563,I170290,I170258,);
not I_9820 (I170539,I170491);
not I_9821 (I170556,I1126843);
nand I_9822 (I170573,I170556,I1126834);
nor I_9823 (I170590,I1126843,I1126846);
nand I_9824 (I170270,I170406,I170590);
nand I_9825 (I170264,I170355,I1126843);
nand I_9826 (I170635,I170457,I1126840);
DFFARX1 I_9827 (I170635,I3563,I170290,I170279,);
DFFARX1 I_9828 (I170635,I3563,I170290,I170273,);
not I_9829 (I170680,I1126840);
nor I_9830 (I170697,I170680,I1126837);
and I_9831 (I170714,I170697,I1126855);
or I_9832 (I170731,I170714,I1126834);
DFFARX1 I_9833 (I170731,I3563,I170290,I170757,);
nand I_9834 (I170765,I170757,I170423);
nor I_9835 (I170267,I170765,I170573);
nor I_9836 (I170261,I170757,I170389);
DFFARX1 I_9837 (I170757,I3563,I170290,I170819,);
not I_9838 (I170827,I170819);
nor I_9839 (I170276,I170827,I170539);
not I_9840 (I170885,I3570);
DFFARX1 I_9841 (I142557,I3563,I170885,I170911,);
DFFARX1 I_9842 (I170911,I3563,I170885,I170928,);
not I_9843 (I170877,I170928);
not I_9844 (I170950,I170911);
DFFARX1 I_9845 (I142551,I3563,I170885,I170976,);
not I_9846 (I170984,I170976);
and I_9847 (I171001,I170950,I142548);
not I_9848 (I171018,I142569);
nand I_9849 (I171035,I171018,I142548);
not I_9850 (I171052,I142563);
nor I_9851 (I171069,I171052,I142554);
nand I_9852 (I171086,I171069,I142560);
nor I_9853 (I171103,I171086,I171035);
DFFARX1 I_9854 (I171103,I3563,I170885,I170853,);
not I_9855 (I171134,I171086);
not I_9856 (I171151,I142554);
nand I_9857 (I171168,I171151,I142548);
nor I_9858 (I171185,I142554,I142569);
nand I_9859 (I170865,I171001,I171185);
nand I_9860 (I170859,I170950,I142554);
nand I_9861 (I171230,I171052,I142548);
DFFARX1 I_9862 (I171230,I3563,I170885,I170874,);
DFFARX1 I_9863 (I171230,I3563,I170885,I170868,);
not I_9864 (I171275,I142548);
nor I_9865 (I171292,I171275,I142566);
and I_9866 (I171309,I171292,I142572);
or I_9867 (I171326,I171309,I142551);
DFFARX1 I_9868 (I171326,I3563,I170885,I171352,);
nand I_9869 (I171360,I171352,I171018);
nor I_9870 (I170862,I171360,I171168);
nor I_9871 (I170856,I171352,I170984);
DFFARX1 I_9872 (I171352,I3563,I170885,I171414,);
not I_9873 (I171422,I171414);
nor I_9874 (I170871,I171422,I171134);
not I_9875 (I171480,I3570);
DFFARX1 I_9876 (I1250779,I3563,I171480,I171506,);
DFFARX1 I_9877 (I171506,I3563,I171480,I171523,);
not I_9878 (I171472,I171523);
not I_9879 (I171545,I171506);
DFFARX1 I_9880 (I1250764,I3563,I171480,I171571,);
not I_9881 (I171579,I171571);
and I_9882 (I171596,I171545,I1250782);
not I_9883 (I171613,I1250764);
nand I_9884 (I171630,I171613,I1250782);
not I_9885 (I171647,I1250785);
nor I_9886 (I171664,I171647,I1250776);
nand I_9887 (I171681,I171664,I1250773);
nor I_9888 (I171698,I171681,I171630);
DFFARX1 I_9889 (I171698,I3563,I171480,I171448,);
not I_9890 (I171729,I171681);
not I_9891 (I171746,I1250776);
nand I_9892 (I171763,I171746,I1250782);
nor I_9893 (I171780,I1250776,I1250764);
nand I_9894 (I171460,I171596,I171780);
nand I_9895 (I171454,I171545,I1250776);
nand I_9896 (I171825,I171647,I1250770);
DFFARX1 I_9897 (I171825,I3563,I171480,I171469,);
DFFARX1 I_9898 (I171825,I3563,I171480,I171463,);
not I_9899 (I171870,I1250770);
nor I_9900 (I171887,I171870,I1250761);
and I_9901 (I171904,I171887,I1250767);
or I_9902 (I171921,I171904,I1250761);
DFFARX1 I_9903 (I171921,I3563,I171480,I171947,);
nand I_9904 (I171955,I171947,I171613);
nor I_9905 (I171457,I171955,I171763);
nor I_9906 (I171451,I171947,I171579);
DFFARX1 I_9907 (I171947,I3563,I171480,I172009,);
not I_9908 (I172017,I172009);
nor I_9909 (I171466,I172017,I171729);
not I_9910 (I172075,I3570);
DFFARX1 I_9911 (I1234917,I3563,I172075,I172101,);
DFFARX1 I_9912 (I172101,I3563,I172075,I172118,);
not I_9913 (I172067,I172118);
not I_9914 (I172140,I172101);
DFFARX1 I_9915 (I1234917,I3563,I172075,I172166,);
not I_9916 (I172174,I172166);
and I_9917 (I172191,I172140,I1234920);
not I_9918 (I172208,I1234932);
nand I_9919 (I172225,I172208,I1234920);
not I_9920 (I172242,I1234938);
nor I_9921 (I172259,I172242,I1234929);
nand I_9922 (I172276,I172259,I1234935);
nor I_9923 (I172293,I172276,I172225);
DFFARX1 I_9924 (I172293,I3563,I172075,I172043,);
not I_9925 (I172324,I172276);
not I_9926 (I172341,I1234929);
nand I_9927 (I172358,I172341,I1234920);
nor I_9928 (I172375,I1234929,I1234932);
nand I_9929 (I172055,I172191,I172375);
nand I_9930 (I172049,I172140,I1234929);
nand I_9931 (I172420,I172242,I1234926);
DFFARX1 I_9932 (I172420,I3563,I172075,I172064,);
DFFARX1 I_9933 (I172420,I3563,I172075,I172058,);
not I_9934 (I172465,I1234926);
nor I_9935 (I172482,I172465,I1234923);
and I_9936 (I172499,I172482,I1234941);
or I_9937 (I172516,I172499,I1234920);
DFFARX1 I_9938 (I172516,I3563,I172075,I172542,);
nand I_9939 (I172550,I172542,I172208);
nor I_9940 (I172052,I172550,I172358);
nor I_9941 (I172046,I172542,I172174);
DFFARX1 I_9942 (I172542,I3563,I172075,I172604,);
not I_9943 (I172612,I172604);
nor I_9944 (I172061,I172612,I172324);
not I_9945 (I172670,I3570);
DFFARX1 I_9946 (I1313188,I3563,I172670,I172696,);
DFFARX1 I_9947 (I172696,I3563,I172670,I172713,);
not I_9948 (I172662,I172713);
not I_9949 (I172735,I172696);
DFFARX1 I_9950 (I1313200,I3563,I172670,I172761,);
not I_9951 (I172769,I172761);
and I_9952 (I172786,I172735,I1313194);
not I_9953 (I172803,I1313206);
nand I_9954 (I172820,I172803,I1313194);
not I_9955 (I172837,I1313191);
nor I_9956 (I172854,I172837,I1313203);
nand I_9957 (I172871,I172854,I1313185);
nor I_9958 (I172888,I172871,I172820);
DFFARX1 I_9959 (I172888,I3563,I172670,I172638,);
not I_9960 (I172919,I172871);
not I_9961 (I172936,I1313203);
nand I_9962 (I172953,I172936,I1313194);
nor I_9963 (I172970,I1313203,I1313206);
nand I_9964 (I172650,I172786,I172970);
nand I_9965 (I172644,I172735,I1313203);
nand I_9966 (I173015,I172837,I1313197);
DFFARX1 I_9967 (I173015,I3563,I172670,I172659,);
DFFARX1 I_9968 (I173015,I3563,I172670,I172653,);
not I_9969 (I173060,I1313197);
nor I_9970 (I173077,I173060,I1313188);
and I_9971 (I173094,I173077,I1313185);
or I_9972 (I173111,I173094,I1313209);
DFFARX1 I_9973 (I173111,I3563,I172670,I173137,);
nand I_9974 (I173145,I173137,I172803);
nor I_9975 (I172647,I173145,I172953);
nor I_9976 (I172641,I173137,I172769);
DFFARX1 I_9977 (I173137,I3563,I172670,I173199,);
not I_9978 (I173207,I173199);
nor I_9979 (I172656,I173207,I172919);
not I_9980 (I173265,I3570);
DFFARX1 I_9981 (I477914,I3563,I173265,I173291,);
DFFARX1 I_9982 (I173291,I3563,I173265,I173308,);
not I_9983 (I173257,I173308);
not I_9984 (I173330,I173291);
DFFARX1 I_9985 (I477902,I3563,I173265,I173356,);
not I_9986 (I173364,I173356);
and I_9987 (I173381,I173330,I477911);
not I_9988 (I173398,I477908);
nand I_9989 (I173415,I173398,I477911);
not I_9990 (I173432,I477899);
nor I_9991 (I173449,I173432,I477905);
nand I_9992 (I173466,I173449,I477890);
nor I_9993 (I173483,I173466,I173415);
DFFARX1 I_9994 (I173483,I3563,I173265,I173233,);
not I_9995 (I173514,I173466);
not I_9996 (I173531,I477905);
nand I_9997 (I173548,I173531,I477911);
nor I_9998 (I173565,I477905,I477908);
nand I_9999 (I173245,I173381,I173565);
nand I_10000 (I173239,I173330,I477905);
nand I_10001 (I173610,I173432,I477890);
DFFARX1 I_10002 (I173610,I3563,I173265,I173254,);
DFFARX1 I_10003 (I173610,I3563,I173265,I173248,);
not I_10004 (I173655,I477890);
nor I_10005 (I173672,I173655,I477896);
and I_10006 (I173689,I173672,I477893);
or I_10007 (I173706,I173689,I477917);
DFFARX1 I_10008 (I173706,I3563,I173265,I173732,);
nand I_10009 (I173740,I173732,I173398);
nor I_10010 (I173242,I173740,I173548);
nor I_10011 (I173236,I173732,I173364);
DFFARX1 I_10012 (I173732,I3563,I173265,I173794,);
not I_10013 (I173802,I173794);
nor I_10014 (I173251,I173802,I173514);
not I_10015 (I173860,I3570);
DFFARX1 I_10016 (I151516,I3563,I173860,I173886,);
DFFARX1 I_10017 (I173886,I3563,I173860,I173903,);
not I_10018 (I173852,I173903);
not I_10019 (I173925,I173886);
DFFARX1 I_10020 (I151510,I3563,I173860,I173951,);
not I_10021 (I173959,I173951);
and I_10022 (I173976,I173925,I151507);
not I_10023 (I173993,I151528);
nand I_10024 (I174010,I173993,I151507);
not I_10025 (I174027,I151522);
nor I_10026 (I174044,I174027,I151513);
nand I_10027 (I174061,I174044,I151519);
nor I_10028 (I174078,I174061,I174010);
DFFARX1 I_10029 (I174078,I3563,I173860,I173828,);
not I_10030 (I174109,I174061);
not I_10031 (I174126,I151513);
nand I_10032 (I174143,I174126,I151507);
nor I_10033 (I174160,I151513,I151528);
nand I_10034 (I173840,I173976,I174160);
nand I_10035 (I173834,I173925,I151513);
nand I_10036 (I174205,I174027,I151507);
DFFARX1 I_10037 (I174205,I3563,I173860,I173849,);
DFFARX1 I_10038 (I174205,I3563,I173860,I173843,);
not I_10039 (I174250,I151507);
nor I_10040 (I174267,I174250,I151525);
and I_10041 (I174284,I174267,I151531);
or I_10042 (I174301,I174284,I151510);
DFFARX1 I_10043 (I174301,I3563,I173860,I174327,);
nand I_10044 (I174335,I174327,I173993);
nor I_10045 (I173837,I174335,I174143);
nor I_10046 (I173831,I174327,I173959);
DFFARX1 I_10047 (I174327,I3563,I173860,I174389,);
not I_10048 (I174397,I174389);
nor I_10049 (I173846,I174397,I174109);
not I_10050 (I174455,I3570);
DFFARX1 I_10051 (I370212,I3563,I174455,I174481,);
DFFARX1 I_10052 (I174481,I3563,I174455,I174498,);
not I_10053 (I174447,I174498);
not I_10054 (I174520,I174481);
DFFARX1 I_10055 (I370227,I3563,I174455,I174546,);
not I_10056 (I174554,I174546);
and I_10057 (I174571,I174520,I370224);
not I_10058 (I174588,I370212);
nand I_10059 (I174605,I174588,I370224);
not I_10060 (I174622,I370221);
nor I_10061 (I174639,I174622,I370236);
nand I_10062 (I174656,I174639,I370233);
nor I_10063 (I174673,I174656,I174605);
DFFARX1 I_10064 (I174673,I3563,I174455,I174423,);
not I_10065 (I174704,I174656);
not I_10066 (I174721,I370236);
nand I_10067 (I174738,I174721,I370224);
nor I_10068 (I174755,I370236,I370212);
nand I_10069 (I174435,I174571,I174755);
nand I_10070 (I174429,I174520,I370236);
nand I_10071 (I174800,I174622,I370230);
DFFARX1 I_10072 (I174800,I3563,I174455,I174444,);
DFFARX1 I_10073 (I174800,I3563,I174455,I174438,);
not I_10074 (I174845,I370230);
nor I_10075 (I174862,I174845,I370218);
and I_10076 (I174879,I174862,I370239);
or I_10077 (I174896,I174879,I370215);
DFFARX1 I_10078 (I174896,I3563,I174455,I174922,);
nand I_10079 (I174930,I174922,I174588);
nor I_10080 (I174432,I174930,I174738);
nor I_10081 (I174426,I174922,I174554);
DFFARX1 I_10082 (I174922,I3563,I174455,I174984,);
not I_10083 (I174992,I174984);
nor I_10084 (I174441,I174992,I174704);
not I_10085 (I175050,I3570);
DFFARX1 I_10086 (I127801,I3563,I175050,I175076,);
DFFARX1 I_10087 (I175076,I3563,I175050,I175093,);
not I_10088 (I175042,I175093);
not I_10089 (I175115,I175076);
DFFARX1 I_10090 (I127795,I3563,I175050,I175141,);
not I_10091 (I175149,I175141);
and I_10092 (I175166,I175115,I127792);
not I_10093 (I175183,I127813);
nand I_10094 (I175200,I175183,I127792);
not I_10095 (I175217,I127807);
nor I_10096 (I175234,I175217,I127798);
nand I_10097 (I175251,I175234,I127804);
nor I_10098 (I175268,I175251,I175200);
DFFARX1 I_10099 (I175268,I3563,I175050,I175018,);
not I_10100 (I175299,I175251);
not I_10101 (I175316,I127798);
nand I_10102 (I175333,I175316,I127792);
nor I_10103 (I175350,I127798,I127813);
nand I_10104 (I175030,I175166,I175350);
nand I_10105 (I175024,I175115,I127798);
nand I_10106 (I175395,I175217,I127792);
DFFARX1 I_10107 (I175395,I3563,I175050,I175039,);
DFFARX1 I_10108 (I175395,I3563,I175050,I175033,);
not I_10109 (I175440,I127792);
nor I_10110 (I175457,I175440,I127810);
and I_10111 (I175474,I175457,I127816);
or I_10112 (I175491,I175474,I127795);
DFFARX1 I_10113 (I175491,I3563,I175050,I175517,);
nand I_10114 (I175525,I175517,I175183);
nor I_10115 (I175027,I175525,I175333);
nor I_10116 (I175021,I175517,I175149);
DFFARX1 I_10117 (I175517,I3563,I175050,I175579,);
not I_10118 (I175587,I175579);
nor I_10119 (I175036,I175587,I175299);
not I_10120 (I175645,I3570);
DFFARX1 I_10121 (I951066,I3563,I175645,I175671,);
DFFARX1 I_10122 (I175671,I3563,I175645,I175688,);
not I_10123 (I175637,I175688);
not I_10124 (I175710,I175671);
DFFARX1 I_10125 (I951075,I3563,I175645,I175736,);
not I_10126 (I175744,I175736);
and I_10127 (I175761,I175710,I951063);
not I_10128 (I175778,I951054);
nand I_10129 (I175795,I175778,I951063);
not I_10130 (I175812,I951060);
nor I_10131 (I175829,I175812,I951078);
nand I_10132 (I175846,I175829,I951051);
nor I_10133 (I175863,I175846,I175795);
DFFARX1 I_10134 (I175863,I3563,I175645,I175613,);
not I_10135 (I175894,I175846);
not I_10136 (I175911,I951078);
nand I_10137 (I175928,I175911,I951063);
nor I_10138 (I175945,I951078,I951054);
nand I_10139 (I175625,I175761,I175945);
nand I_10140 (I175619,I175710,I951078);
nand I_10141 (I175990,I175812,I951057);
DFFARX1 I_10142 (I175990,I3563,I175645,I175634,);
DFFARX1 I_10143 (I175990,I3563,I175645,I175628,);
not I_10144 (I176035,I951057);
nor I_10145 (I176052,I176035,I951069);
and I_10146 (I176069,I176052,I951051);
or I_10147 (I176086,I176069,I951072);
DFFARX1 I_10148 (I176086,I3563,I175645,I176112,);
nand I_10149 (I176120,I176112,I175778);
nor I_10150 (I175622,I176120,I175928);
nor I_10151 (I175616,I176112,I175744);
DFFARX1 I_10152 (I176112,I3563,I175645,I176174,);
not I_10153 (I176182,I176174);
nor I_10154 (I175631,I176182,I175894);
not I_10155 (I176240,I3570);
DFFARX1 I_10156 (I661893,I3563,I176240,I176266,);
DFFARX1 I_10157 (I176266,I3563,I176240,I176283,);
not I_10158 (I176232,I176283);
not I_10159 (I176305,I176266);
DFFARX1 I_10160 (I661890,I3563,I176240,I176331,);
not I_10161 (I176339,I176331);
and I_10162 (I176356,I176305,I661896);
not I_10163 (I176373,I661881);
nand I_10164 (I176390,I176373,I661896);
not I_10165 (I176407,I661884);
nor I_10166 (I176424,I176407,I661905);
nand I_10167 (I176441,I176424,I661902);
nor I_10168 (I176458,I176441,I176390);
DFFARX1 I_10169 (I176458,I3563,I176240,I176208,);
not I_10170 (I176489,I176441);
not I_10171 (I176506,I661905);
nand I_10172 (I176523,I176506,I661896);
nor I_10173 (I176540,I661905,I661881);
nand I_10174 (I176220,I176356,I176540);
nand I_10175 (I176214,I176305,I661905);
nand I_10176 (I176585,I176407,I661881);
DFFARX1 I_10177 (I176585,I3563,I176240,I176229,);
DFFARX1 I_10178 (I176585,I3563,I176240,I176223,);
not I_10179 (I176630,I661881);
nor I_10180 (I176647,I176630,I661887);
and I_10181 (I176664,I176647,I661899);
or I_10182 (I176681,I176664,I661884);
DFFARX1 I_10183 (I176681,I3563,I176240,I176707,);
nand I_10184 (I176715,I176707,I176373);
nor I_10185 (I176217,I176715,I176523);
nor I_10186 (I176211,I176707,I176339);
DFFARX1 I_10187 (I176707,I3563,I176240,I176769,);
not I_10188 (I176777,I176769);
nor I_10189 (I176226,I176777,I176489);
not I_10190 (I176835,I3570);
DFFARX1 I_10191 (I1066858,I3563,I176835,I176861,);
DFFARX1 I_10192 (I176861,I3563,I176835,I176878,);
not I_10193 (I176827,I176878);
not I_10194 (I176900,I176861);
DFFARX1 I_10195 (I1066867,I3563,I176835,I176926,);
not I_10196 (I176934,I176926);
and I_10197 (I176951,I176900,I1066861);
not I_10198 (I176968,I1066855);
nand I_10199 (I176985,I176968,I1066861);
not I_10200 (I177002,I1066870);
nor I_10201 (I177019,I177002,I1066858);
nand I_10202 (I177036,I177019,I1066864);
nor I_10203 (I177053,I177036,I176985);
DFFARX1 I_10204 (I177053,I3563,I176835,I176803,);
not I_10205 (I177084,I177036);
not I_10206 (I177101,I1066858);
nand I_10207 (I177118,I177101,I1066861);
nor I_10208 (I177135,I1066858,I1066855);
nand I_10209 (I176815,I176951,I177135);
nand I_10210 (I176809,I176900,I1066858);
nand I_10211 (I177180,I177002,I1066861);
DFFARX1 I_10212 (I177180,I3563,I176835,I176824,);
DFFARX1 I_10213 (I177180,I3563,I176835,I176818,);
not I_10214 (I177225,I1066861);
nor I_10215 (I177242,I177225,I1066876);
and I_10216 (I177259,I177242,I1066873);
or I_10217 (I177276,I177259,I1066855);
DFFARX1 I_10218 (I177276,I3563,I176835,I177302,);
nand I_10219 (I177310,I177302,I176968);
nor I_10220 (I176812,I177310,I177118);
nor I_10221 (I176806,I177302,I176934);
DFFARX1 I_10222 (I177302,I3563,I176835,I177364,);
not I_10223 (I177372,I177364);
nor I_10224 (I176821,I177372,I177084);
not I_10225 (I177430,I3570);
DFFARX1 I_10226 (I896436,I3563,I177430,I177456,);
DFFARX1 I_10227 (I177456,I3563,I177430,I177473,);
not I_10228 (I177422,I177473);
not I_10229 (I177495,I177456);
DFFARX1 I_10230 (I896430,I3563,I177430,I177521,);
not I_10231 (I177529,I177521);
and I_10232 (I177546,I177495,I896448);
not I_10233 (I177563,I896436);
nand I_10234 (I177580,I177563,I896448);
not I_10235 (I177597,I896430);
nor I_10236 (I177614,I177597,I896442);
nand I_10237 (I177631,I177614,I896433);
nor I_10238 (I177648,I177631,I177580);
DFFARX1 I_10239 (I177648,I3563,I177430,I177398,);
not I_10240 (I177679,I177631);
not I_10241 (I177696,I896442);
nand I_10242 (I177713,I177696,I896448);
nor I_10243 (I177730,I896442,I896436);
nand I_10244 (I177410,I177546,I177730);
nand I_10245 (I177404,I177495,I896442);
nand I_10246 (I177775,I177597,I896445);
DFFARX1 I_10247 (I177775,I3563,I177430,I177419,);
DFFARX1 I_10248 (I177775,I3563,I177430,I177413,);
not I_10249 (I177820,I896445);
nor I_10250 (I177837,I177820,I896451);
and I_10251 (I177854,I177837,I896433);
or I_10252 (I177871,I177854,I896439);
DFFARX1 I_10253 (I177871,I3563,I177430,I177897,);
nand I_10254 (I177905,I177897,I177563);
nor I_10255 (I177407,I177905,I177713);
nor I_10256 (I177401,I177897,I177529);
DFFARX1 I_10257 (I177897,I3563,I177430,I177959,);
not I_10258 (I177967,I177959);
nor I_10259 (I177416,I177967,I177679);
not I_10260 (I178025,I3570);
DFFARX1 I_10261 (I1107757,I3563,I178025,I178051,);
DFFARX1 I_10262 (I178051,I3563,I178025,I178068,);
not I_10263 (I178017,I178068);
not I_10264 (I178090,I178051);
DFFARX1 I_10265 (I1107757,I3563,I178025,I178116,);
not I_10266 (I178124,I178116);
and I_10267 (I178141,I178090,I1107760);
not I_10268 (I178158,I1107772);
nand I_10269 (I178175,I178158,I1107760);
not I_10270 (I178192,I1107778);
nor I_10271 (I178209,I178192,I1107769);
nand I_10272 (I178226,I178209,I1107775);
nor I_10273 (I178243,I178226,I178175);
DFFARX1 I_10274 (I178243,I3563,I178025,I177993,);
not I_10275 (I178274,I178226);
not I_10276 (I178291,I1107769);
nand I_10277 (I178308,I178291,I1107760);
nor I_10278 (I178325,I1107769,I1107772);
nand I_10279 (I178005,I178141,I178325);
nand I_10280 (I177999,I178090,I1107769);
nand I_10281 (I178370,I178192,I1107766);
DFFARX1 I_10282 (I178370,I3563,I178025,I178014,);
DFFARX1 I_10283 (I178370,I3563,I178025,I178008,);
not I_10284 (I178415,I1107766);
nor I_10285 (I178432,I178415,I1107763);
and I_10286 (I178449,I178432,I1107781);
or I_10287 (I178466,I178449,I1107760);
DFFARX1 I_10288 (I178466,I3563,I178025,I178492,);
nand I_10289 (I178500,I178492,I178158);
nor I_10290 (I178002,I178500,I178308);
nor I_10291 (I177996,I178492,I178124);
DFFARX1 I_10292 (I178492,I3563,I178025,I178554,);
not I_10293 (I178562,I178554);
nor I_10294 (I178011,I178562,I178274);
not I_10295 (I178620,I3570);
DFFARX1 I_10296 (I714491,I3563,I178620,I178646,);
DFFARX1 I_10297 (I178646,I3563,I178620,I178663,);
not I_10298 (I178612,I178663);
not I_10299 (I178685,I178646);
DFFARX1 I_10300 (I714488,I3563,I178620,I178711,);
not I_10301 (I178719,I178711);
and I_10302 (I178736,I178685,I714494);
not I_10303 (I178753,I714479);
nand I_10304 (I178770,I178753,I714494);
not I_10305 (I178787,I714482);
nor I_10306 (I178804,I178787,I714503);
nand I_10307 (I178821,I178804,I714500);
nor I_10308 (I178838,I178821,I178770);
DFFARX1 I_10309 (I178838,I3563,I178620,I178588,);
not I_10310 (I178869,I178821);
not I_10311 (I178886,I714503);
nand I_10312 (I178903,I178886,I714494);
nor I_10313 (I178920,I714503,I714479);
nand I_10314 (I178600,I178736,I178920);
nand I_10315 (I178594,I178685,I714503);
nand I_10316 (I178965,I178787,I714479);
DFFARX1 I_10317 (I178965,I3563,I178620,I178609,);
DFFARX1 I_10318 (I178965,I3563,I178620,I178603,);
not I_10319 (I179010,I714479);
nor I_10320 (I179027,I179010,I714485);
and I_10321 (I179044,I179027,I714497);
or I_10322 (I179061,I179044,I714482);
DFFARX1 I_10323 (I179061,I3563,I178620,I179087,);
nand I_10324 (I179095,I179087,I178753);
nor I_10325 (I178597,I179095,I178903);
nor I_10326 (I178591,I179087,I178719);
DFFARX1 I_10327 (I179087,I3563,I178620,I179149,);
not I_10328 (I179157,I179149);
nor I_10329 (I178606,I179157,I178869);
not I_10330 (I179215,I3570);
DFFARX1 I_10331 (I414480,I3563,I179215,I179241,);
DFFARX1 I_10332 (I179241,I3563,I179215,I179258,);
not I_10333 (I179207,I179258);
not I_10334 (I179280,I179241);
DFFARX1 I_10335 (I414495,I3563,I179215,I179306,);
not I_10336 (I179314,I179306);
and I_10337 (I179331,I179280,I414492);
not I_10338 (I179348,I414480);
nand I_10339 (I179365,I179348,I414492);
not I_10340 (I179382,I414489);
nor I_10341 (I179399,I179382,I414504);
nand I_10342 (I179416,I179399,I414501);
nor I_10343 (I179433,I179416,I179365);
DFFARX1 I_10344 (I179433,I3563,I179215,I179183,);
not I_10345 (I179464,I179416);
not I_10346 (I179481,I414504);
nand I_10347 (I179498,I179481,I414492);
nor I_10348 (I179515,I414504,I414480);
nand I_10349 (I179195,I179331,I179515);
nand I_10350 (I179189,I179280,I414504);
nand I_10351 (I179560,I179382,I414498);
DFFARX1 I_10352 (I179560,I3563,I179215,I179204,);
DFFARX1 I_10353 (I179560,I3563,I179215,I179198,);
not I_10354 (I179605,I414498);
nor I_10355 (I179622,I179605,I414486);
and I_10356 (I179639,I179622,I414507);
or I_10357 (I179656,I179639,I414483);
DFFARX1 I_10358 (I179656,I3563,I179215,I179682,);
nand I_10359 (I179690,I179682,I179348);
nor I_10360 (I179192,I179690,I179498);
nor I_10361 (I179186,I179682,I179314);
DFFARX1 I_10362 (I179682,I3563,I179215,I179744,);
not I_10363 (I179752,I179744);
nor I_10364 (I179201,I179752,I179464);
not I_10365 (I179810,I3570);
DFFARX1 I_10366 (I760153,I3563,I179810,I179836,);
DFFARX1 I_10367 (I179836,I3563,I179810,I179853,);
not I_10368 (I179802,I179853);
not I_10369 (I179875,I179836);
DFFARX1 I_10370 (I760150,I3563,I179810,I179901,);
not I_10371 (I179909,I179901);
and I_10372 (I179926,I179875,I760156);
not I_10373 (I179943,I760141);
nand I_10374 (I179960,I179943,I760156);
not I_10375 (I179977,I760144);
nor I_10376 (I179994,I179977,I760165);
nand I_10377 (I180011,I179994,I760162);
nor I_10378 (I180028,I180011,I179960);
DFFARX1 I_10379 (I180028,I3563,I179810,I179778,);
not I_10380 (I180059,I180011);
not I_10381 (I180076,I760165);
nand I_10382 (I180093,I180076,I760156);
nor I_10383 (I180110,I760165,I760141);
nand I_10384 (I179790,I179926,I180110);
nand I_10385 (I179784,I179875,I760165);
nand I_10386 (I180155,I179977,I760141);
DFFARX1 I_10387 (I180155,I3563,I179810,I179799,);
DFFARX1 I_10388 (I180155,I3563,I179810,I179793,);
not I_10389 (I180200,I760141);
nor I_10390 (I180217,I180200,I760147);
and I_10391 (I180234,I180217,I760159);
or I_10392 (I180251,I180234,I760144);
DFFARX1 I_10393 (I180251,I3563,I179810,I180277,);
nand I_10394 (I180285,I180277,I179943);
nor I_10395 (I179787,I180285,I180093);
nor I_10396 (I179781,I180277,I179909);
DFFARX1 I_10397 (I180277,I3563,I179810,I180339,);
not I_10398 (I180347,I180339);
nor I_10399 (I179796,I180347,I180059);
not I_10400 (I180405,I3570);
DFFARX1 I_10401 (I116207,I3563,I180405,I180431,);
DFFARX1 I_10402 (I180431,I3563,I180405,I180448,);
not I_10403 (I180397,I180448);
not I_10404 (I180470,I180431);
DFFARX1 I_10405 (I116201,I3563,I180405,I180496,);
not I_10406 (I180504,I180496);
and I_10407 (I180521,I180470,I116198);
not I_10408 (I180538,I116219);
nand I_10409 (I180555,I180538,I116198);
not I_10410 (I180572,I116213);
nor I_10411 (I180589,I180572,I116204);
nand I_10412 (I180606,I180589,I116210);
nor I_10413 (I180623,I180606,I180555);
DFFARX1 I_10414 (I180623,I3563,I180405,I180373,);
not I_10415 (I180654,I180606);
not I_10416 (I180671,I116204);
nand I_10417 (I180688,I180671,I116198);
nor I_10418 (I180705,I116204,I116219);
nand I_10419 (I180385,I180521,I180705);
nand I_10420 (I180379,I180470,I116204);
nand I_10421 (I180750,I180572,I116198);
DFFARX1 I_10422 (I180750,I3563,I180405,I180394,);
DFFARX1 I_10423 (I180750,I3563,I180405,I180388,);
not I_10424 (I180795,I116198);
nor I_10425 (I180812,I180795,I116216);
and I_10426 (I180829,I180812,I116222);
or I_10427 (I180846,I180829,I116201);
DFFARX1 I_10428 (I180846,I3563,I180405,I180872,);
nand I_10429 (I180880,I180872,I180538);
nor I_10430 (I180382,I180880,I180688);
nor I_10431 (I180376,I180872,I180504);
DFFARX1 I_10432 (I180872,I3563,I180405,I180934,);
not I_10433 (I180942,I180934);
nor I_10434 (I180391,I180942,I180654);
not I_10435 (I181000,I3570);
DFFARX1 I_10436 (I328579,I3563,I181000,I181026,);
DFFARX1 I_10437 (I181026,I3563,I181000,I181043,);
not I_10438 (I180992,I181043);
not I_10439 (I181065,I181026);
DFFARX1 I_10440 (I328594,I3563,I181000,I181091,);
not I_10441 (I181099,I181091);
and I_10442 (I181116,I181065,I328591);
not I_10443 (I181133,I328579);
nand I_10444 (I181150,I181133,I328591);
not I_10445 (I181167,I328588);
nor I_10446 (I181184,I181167,I328603);
nand I_10447 (I181201,I181184,I328600);
nor I_10448 (I181218,I181201,I181150);
DFFARX1 I_10449 (I181218,I3563,I181000,I180968,);
not I_10450 (I181249,I181201);
not I_10451 (I181266,I328603);
nand I_10452 (I181283,I181266,I328591);
nor I_10453 (I181300,I328603,I328579);
nand I_10454 (I180980,I181116,I181300);
nand I_10455 (I180974,I181065,I328603);
nand I_10456 (I181345,I181167,I328597);
DFFARX1 I_10457 (I181345,I3563,I181000,I180989,);
DFFARX1 I_10458 (I181345,I3563,I181000,I180983,);
not I_10459 (I181390,I328597);
nor I_10460 (I181407,I181390,I328585);
and I_10461 (I181424,I181407,I328606);
or I_10462 (I181441,I181424,I328582);
DFFARX1 I_10463 (I181441,I3563,I181000,I181467,);
nand I_10464 (I181475,I181467,I181133);
nor I_10465 (I180977,I181475,I181283);
nor I_10466 (I180971,I181467,I181099);
DFFARX1 I_10467 (I181467,I3563,I181000,I181529,);
not I_10468 (I181537,I181529);
nor I_10469 (I180986,I181537,I181249);
not I_10470 (I181595,I3570);
DFFARX1 I_10471 (I735877,I3563,I181595,I181621,);
DFFARX1 I_10472 (I181621,I3563,I181595,I181638,);
not I_10473 (I181587,I181638);
not I_10474 (I181660,I181621);
DFFARX1 I_10475 (I735874,I3563,I181595,I181686,);
not I_10476 (I181694,I181686);
and I_10477 (I181711,I181660,I735880);
not I_10478 (I181728,I735865);
nand I_10479 (I181745,I181728,I735880);
not I_10480 (I181762,I735868);
nor I_10481 (I181779,I181762,I735889);
nand I_10482 (I181796,I181779,I735886);
nor I_10483 (I181813,I181796,I181745);
DFFARX1 I_10484 (I181813,I3563,I181595,I181563,);
not I_10485 (I181844,I181796);
not I_10486 (I181861,I735889);
nand I_10487 (I181878,I181861,I735880);
nor I_10488 (I181895,I735889,I735865);
nand I_10489 (I181575,I181711,I181895);
nand I_10490 (I181569,I181660,I735889);
nand I_10491 (I181940,I181762,I735865);
DFFARX1 I_10492 (I181940,I3563,I181595,I181584,);
DFFARX1 I_10493 (I181940,I3563,I181595,I181578,);
not I_10494 (I181985,I735865);
nor I_10495 (I182002,I181985,I735871);
and I_10496 (I182019,I182002,I735883);
or I_10497 (I182036,I182019,I735868);
DFFARX1 I_10498 (I182036,I3563,I181595,I182062,);
nand I_10499 (I182070,I182062,I181728);
nor I_10500 (I181572,I182070,I181878);
nor I_10501 (I181566,I182062,I181694);
DFFARX1 I_10502 (I182062,I3563,I181595,I182124,);
not I_10503 (I182132,I182124);
nor I_10504 (I181581,I182132,I181844);
not I_10505 (I182190,I3570);
DFFARX1 I_10506 (I141503,I3563,I182190,I182216,);
DFFARX1 I_10507 (I182216,I3563,I182190,I182233,);
not I_10508 (I182182,I182233);
not I_10509 (I182255,I182216);
DFFARX1 I_10510 (I141497,I3563,I182190,I182281,);
not I_10511 (I182289,I182281);
and I_10512 (I182306,I182255,I141494);
not I_10513 (I182323,I141515);
nand I_10514 (I182340,I182323,I141494);
not I_10515 (I182357,I141509);
nor I_10516 (I182374,I182357,I141500);
nand I_10517 (I182391,I182374,I141506);
nor I_10518 (I182408,I182391,I182340);
DFFARX1 I_10519 (I182408,I3563,I182190,I182158,);
not I_10520 (I182439,I182391);
not I_10521 (I182456,I141500);
nand I_10522 (I182473,I182456,I141494);
nor I_10523 (I182490,I141500,I141515);
nand I_10524 (I182170,I182306,I182490);
nand I_10525 (I182164,I182255,I141500);
nand I_10526 (I182535,I182357,I141494);
DFFARX1 I_10527 (I182535,I3563,I182190,I182179,);
DFFARX1 I_10528 (I182535,I3563,I182190,I182173,);
not I_10529 (I182580,I141494);
nor I_10530 (I182597,I182580,I141512);
and I_10531 (I182614,I182597,I141518);
or I_10532 (I182631,I182614,I141497);
DFFARX1 I_10533 (I182631,I3563,I182190,I182657,);
nand I_10534 (I182665,I182657,I182323);
nor I_10535 (I182167,I182665,I182473);
nor I_10536 (I182161,I182657,I182289);
DFFARX1 I_10537 (I182657,I3563,I182190,I182719,);
not I_10538 (I182727,I182719);
nor I_10539 (I182176,I182727,I182439);
not I_10540 (I182785,I3570);
DFFARX1 I_10541 (I1297004,I3563,I182785,I182811,);
DFFARX1 I_10542 (I182811,I3563,I182785,I182828,);
not I_10543 (I182777,I182828);
not I_10544 (I182850,I182811);
DFFARX1 I_10545 (I1297016,I3563,I182785,I182876,);
not I_10546 (I182884,I182876);
and I_10547 (I182901,I182850,I1297010);
not I_10548 (I182918,I1297022);
nand I_10549 (I182935,I182918,I1297010);
not I_10550 (I182952,I1297007);
nor I_10551 (I182969,I182952,I1297019);
nand I_10552 (I182986,I182969,I1297001);
nor I_10553 (I183003,I182986,I182935);
DFFARX1 I_10554 (I183003,I3563,I182785,I182753,);
not I_10555 (I183034,I182986);
not I_10556 (I183051,I1297019);
nand I_10557 (I183068,I183051,I1297010);
nor I_10558 (I183085,I1297019,I1297022);
nand I_10559 (I182765,I182901,I183085);
nand I_10560 (I182759,I182850,I1297019);
nand I_10561 (I183130,I182952,I1297013);
DFFARX1 I_10562 (I183130,I3563,I182785,I182774,);
DFFARX1 I_10563 (I183130,I3563,I182785,I182768,);
not I_10564 (I183175,I1297013);
nor I_10565 (I183192,I183175,I1297004);
and I_10566 (I183209,I183192,I1297001);
or I_10567 (I183226,I183209,I1297025);
DFFARX1 I_10568 (I183226,I3563,I182785,I183252,);
nand I_10569 (I183260,I183252,I182918);
nor I_10570 (I182762,I183260,I183068);
nor I_10571 (I182756,I183252,I182884);
DFFARX1 I_10572 (I183252,I3563,I182785,I183314,);
not I_10573 (I183322,I183314);
nor I_10574 (I182771,I183322,I183034);
not I_10575 (I183380,I3570);
DFFARX1 I_10576 (I690215,I3563,I183380,I183406,);
DFFARX1 I_10577 (I183406,I3563,I183380,I183423,);
not I_10578 (I183372,I183423);
not I_10579 (I183445,I183406);
DFFARX1 I_10580 (I690212,I3563,I183380,I183471,);
not I_10581 (I183479,I183471);
and I_10582 (I183496,I183445,I690218);
not I_10583 (I183513,I690203);
nand I_10584 (I183530,I183513,I690218);
not I_10585 (I183547,I690206);
nor I_10586 (I183564,I183547,I690227);
nand I_10587 (I183581,I183564,I690224);
nor I_10588 (I183598,I183581,I183530);
DFFARX1 I_10589 (I183598,I3563,I183380,I183348,);
not I_10590 (I183629,I183581);
not I_10591 (I183646,I690227);
nand I_10592 (I183663,I183646,I690218);
nor I_10593 (I183680,I690227,I690203);
nand I_10594 (I183360,I183496,I183680);
nand I_10595 (I183354,I183445,I690227);
nand I_10596 (I183725,I183547,I690203);
DFFARX1 I_10597 (I183725,I3563,I183380,I183369,);
DFFARX1 I_10598 (I183725,I3563,I183380,I183363,);
not I_10599 (I183770,I690203);
nor I_10600 (I183787,I183770,I690209);
and I_10601 (I183804,I183787,I690221);
or I_10602 (I183821,I183804,I690206);
DFFARX1 I_10603 (I183821,I3563,I183380,I183847,);
nand I_10604 (I183855,I183847,I183513);
nor I_10605 (I183357,I183855,I183663);
nor I_10606 (I183351,I183847,I183479);
DFFARX1 I_10607 (I183847,I3563,I183380,I183909,);
not I_10608 (I183917,I183909);
nor I_10609 (I183366,I183917,I183629);
not I_10610 (I183975,I3570);
DFFARX1 I_10611 (I591380,I3563,I183975,I184001,);
DFFARX1 I_10612 (I184001,I3563,I183975,I184018,);
not I_10613 (I183967,I184018);
not I_10614 (I184040,I184001);
DFFARX1 I_10615 (I591371,I3563,I183975,I184066,);
not I_10616 (I184074,I184066);
and I_10617 (I184091,I184040,I591389);
not I_10618 (I184108,I591386);
nand I_10619 (I184125,I184108,I591389);
not I_10620 (I184142,I591365);
nor I_10621 (I184159,I184142,I591368);
nand I_10622 (I184176,I184159,I591377);
nor I_10623 (I184193,I184176,I184125);
DFFARX1 I_10624 (I184193,I3563,I183975,I183943,);
not I_10625 (I184224,I184176);
not I_10626 (I184241,I591368);
nand I_10627 (I184258,I184241,I591389);
nor I_10628 (I184275,I591368,I591386);
nand I_10629 (I183955,I184091,I184275);
nand I_10630 (I183949,I184040,I591368);
nand I_10631 (I184320,I184142,I591383);
DFFARX1 I_10632 (I184320,I3563,I183975,I183964,);
DFFARX1 I_10633 (I184320,I3563,I183975,I183958,);
not I_10634 (I184365,I591383);
nor I_10635 (I184382,I184365,I591365);
and I_10636 (I184399,I184382,I591374);
or I_10637 (I184416,I184399,I591368);
DFFARX1 I_10638 (I184416,I3563,I183975,I184442,);
nand I_10639 (I184450,I184442,I184108);
nor I_10640 (I183952,I184450,I184258);
nor I_10641 (I183946,I184442,I184074);
DFFARX1 I_10642 (I184442,I3563,I183975,I184504,);
not I_10643 (I184512,I184504);
nor I_10644 (I183961,I184512,I184224);
not I_10645 (I184570,I3570);
DFFARX1 I_10646 (I614500,I3563,I184570,I184596,);
DFFARX1 I_10647 (I184596,I3563,I184570,I184613,);
not I_10648 (I184562,I184613);
not I_10649 (I184635,I184596);
DFFARX1 I_10650 (I614491,I3563,I184570,I184661,);
not I_10651 (I184669,I184661);
and I_10652 (I184686,I184635,I614509);
not I_10653 (I184703,I614506);
nand I_10654 (I184720,I184703,I614509);
not I_10655 (I184737,I614485);
nor I_10656 (I184754,I184737,I614488);
nand I_10657 (I184771,I184754,I614497);
nor I_10658 (I184788,I184771,I184720);
DFFARX1 I_10659 (I184788,I3563,I184570,I184538,);
not I_10660 (I184819,I184771);
not I_10661 (I184836,I614488);
nand I_10662 (I184853,I184836,I614509);
nor I_10663 (I184870,I614488,I614506);
nand I_10664 (I184550,I184686,I184870);
nand I_10665 (I184544,I184635,I614488);
nand I_10666 (I184915,I184737,I614503);
DFFARX1 I_10667 (I184915,I3563,I184570,I184559,);
DFFARX1 I_10668 (I184915,I3563,I184570,I184553,);
not I_10669 (I184960,I614503);
nor I_10670 (I184977,I184960,I614485);
and I_10671 (I184994,I184977,I614494);
or I_10672 (I185011,I184994,I614488);
DFFARX1 I_10673 (I185011,I3563,I184570,I185037,);
nand I_10674 (I185045,I185037,I184703);
nor I_10675 (I184547,I185045,I184853);
nor I_10676 (I184541,I185037,I184669);
DFFARX1 I_10677 (I185037,I3563,I184570,I185099,);
not I_10678 (I185107,I185099);
nor I_10679 (I184556,I185107,I184819);
not I_10680 (I185165,I3570);
DFFARX1 I_10681 (I1257851,I3563,I185165,I185191,);
DFFARX1 I_10682 (I185191,I3563,I185165,I185208,);
not I_10683 (I185157,I185208);
not I_10684 (I185230,I185191);
DFFARX1 I_10685 (I1257836,I3563,I185165,I185256,);
not I_10686 (I185264,I185256);
and I_10687 (I185281,I185230,I1257854);
not I_10688 (I185298,I1257836);
nand I_10689 (I185315,I185298,I1257854);
not I_10690 (I185332,I1257857);
nor I_10691 (I185349,I185332,I1257848);
nand I_10692 (I185366,I185349,I1257845);
nor I_10693 (I185383,I185366,I185315);
DFFARX1 I_10694 (I185383,I3563,I185165,I185133,);
not I_10695 (I185414,I185366);
not I_10696 (I185431,I1257848);
nand I_10697 (I185448,I185431,I1257854);
nor I_10698 (I185465,I1257848,I1257836);
nand I_10699 (I185145,I185281,I185465);
nand I_10700 (I185139,I185230,I1257848);
nand I_10701 (I185510,I185332,I1257842);
DFFARX1 I_10702 (I185510,I3563,I185165,I185154,);
DFFARX1 I_10703 (I185510,I3563,I185165,I185148,);
not I_10704 (I185555,I1257842);
nor I_10705 (I185572,I185555,I1257833);
and I_10706 (I185589,I185572,I1257839);
or I_10707 (I185606,I185589,I1257833);
DFFARX1 I_10708 (I185606,I3563,I185165,I185632,);
nand I_10709 (I185640,I185632,I185298);
nor I_10710 (I185142,I185640,I185448);
nor I_10711 (I185136,I185632,I185264);
DFFARX1 I_10712 (I185632,I3563,I185165,I185694,);
not I_10713 (I185702,I185694);
nor I_10714 (I185151,I185702,I185414);
not I_10715 (I185760,I3570);
DFFARX1 I_10716 (I1051150,I3563,I185760,I185786,);
DFFARX1 I_10717 (I185786,I3563,I185760,I185803,);
not I_10718 (I185752,I185803);
not I_10719 (I185825,I185786);
DFFARX1 I_10720 (I1051159,I3563,I185760,I185851,);
not I_10721 (I185859,I185851);
and I_10722 (I185876,I185825,I1051153);
not I_10723 (I185893,I1051147);
nand I_10724 (I185910,I185893,I1051153);
not I_10725 (I185927,I1051162);
nor I_10726 (I185944,I185927,I1051150);
nand I_10727 (I185961,I185944,I1051156);
nor I_10728 (I185978,I185961,I185910);
DFFARX1 I_10729 (I185978,I3563,I185760,I185728,);
not I_10730 (I186009,I185961);
not I_10731 (I186026,I1051150);
nand I_10732 (I186043,I186026,I1051153);
nor I_10733 (I186060,I1051150,I1051147);
nand I_10734 (I185740,I185876,I186060);
nand I_10735 (I185734,I185825,I1051150);
nand I_10736 (I186105,I185927,I1051153);
DFFARX1 I_10737 (I186105,I3563,I185760,I185749,);
DFFARX1 I_10738 (I186105,I3563,I185760,I185743,);
not I_10739 (I186150,I1051153);
nor I_10740 (I186167,I186150,I1051168);
and I_10741 (I186184,I186167,I1051165);
or I_10742 (I186201,I186184,I1051147);
DFFARX1 I_10743 (I186201,I3563,I185760,I186227,);
nand I_10744 (I186235,I186227,I185893);
nor I_10745 (I185737,I186235,I186043);
nor I_10746 (I185731,I186227,I185859);
DFFARX1 I_10747 (I186227,I3563,I185760,I186289,);
not I_10748 (I186297,I186289);
nor I_10749 (I185746,I186297,I186009);
not I_10750 (I186355,I3570);
DFFARX1 I_10751 (I485530,I3563,I186355,I186381,);
DFFARX1 I_10752 (I186381,I3563,I186355,I186398,);
not I_10753 (I186347,I186398);
not I_10754 (I186420,I186381);
DFFARX1 I_10755 (I485518,I3563,I186355,I186446,);
not I_10756 (I186454,I186446);
and I_10757 (I186471,I186420,I485527);
not I_10758 (I186488,I485524);
nand I_10759 (I186505,I186488,I485527);
not I_10760 (I186522,I485515);
nor I_10761 (I186539,I186522,I485521);
nand I_10762 (I186556,I186539,I485506);
nor I_10763 (I186573,I186556,I186505);
DFFARX1 I_10764 (I186573,I3563,I186355,I186323,);
not I_10765 (I186604,I186556);
not I_10766 (I186621,I485521);
nand I_10767 (I186638,I186621,I485527);
nor I_10768 (I186655,I485521,I485524);
nand I_10769 (I186335,I186471,I186655);
nand I_10770 (I186329,I186420,I485521);
nand I_10771 (I186700,I186522,I485506);
DFFARX1 I_10772 (I186700,I3563,I186355,I186344,);
DFFARX1 I_10773 (I186700,I3563,I186355,I186338,);
not I_10774 (I186745,I485506);
nor I_10775 (I186762,I186745,I485512);
and I_10776 (I186779,I186762,I485509);
or I_10777 (I186796,I186779,I485533);
DFFARX1 I_10778 (I186796,I3563,I186355,I186822,);
nand I_10779 (I186830,I186822,I186488);
nor I_10780 (I186332,I186830,I186638);
nor I_10781 (I186326,I186822,I186454);
DFFARX1 I_10782 (I186822,I3563,I186355,I186884,);
not I_10783 (I186892,I186884);
nor I_10784 (I186341,I186892,I186604);
not I_10785 (I186950,I3570);
DFFARX1 I_10786 (I593692,I3563,I186950,I186976,);
DFFARX1 I_10787 (I186976,I3563,I186950,I186993,);
not I_10788 (I186942,I186993);
not I_10789 (I187015,I186976);
DFFARX1 I_10790 (I593683,I3563,I186950,I187041,);
not I_10791 (I187049,I187041);
and I_10792 (I187066,I187015,I593701);
not I_10793 (I187083,I593698);
nand I_10794 (I187100,I187083,I593701);
not I_10795 (I187117,I593677);
nor I_10796 (I187134,I187117,I593680);
nand I_10797 (I187151,I187134,I593689);
nor I_10798 (I187168,I187151,I187100);
DFFARX1 I_10799 (I187168,I3563,I186950,I186918,);
not I_10800 (I187199,I187151);
not I_10801 (I187216,I593680);
nand I_10802 (I187233,I187216,I593701);
nor I_10803 (I187250,I593680,I593698);
nand I_10804 (I186930,I187066,I187250);
nand I_10805 (I186924,I187015,I593680);
nand I_10806 (I187295,I187117,I593695);
DFFARX1 I_10807 (I187295,I3563,I186950,I186939,);
DFFARX1 I_10808 (I187295,I3563,I186950,I186933,);
not I_10809 (I187340,I593695);
nor I_10810 (I187357,I187340,I593677);
and I_10811 (I187374,I187357,I593686);
or I_10812 (I187391,I187374,I593680);
DFFARX1 I_10813 (I187391,I3563,I186950,I187417,);
nand I_10814 (I187425,I187417,I187083);
nor I_10815 (I186927,I187425,I187233);
nor I_10816 (I186921,I187417,I187049);
DFFARX1 I_10817 (I187417,I3563,I186950,I187479,);
not I_10818 (I187487,I187479);
nor I_10819 (I186936,I187487,I187199);
not I_10820 (I187545,I3570);
DFFARX1 I_10821 (I578664,I3563,I187545,I187571,);
DFFARX1 I_10822 (I187571,I3563,I187545,I187588,);
not I_10823 (I187537,I187588);
not I_10824 (I187610,I187571);
DFFARX1 I_10825 (I578655,I3563,I187545,I187636,);
not I_10826 (I187644,I187636);
and I_10827 (I187661,I187610,I578673);
not I_10828 (I187678,I578670);
nand I_10829 (I187695,I187678,I578673);
not I_10830 (I187712,I578649);
nor I_10831 (I187729,I187712,I578652);
nand I_10832 (I187746,I187729,I578661);
nor I_10833 (I187763,I187746,I187695);
DFFARX1 I_10834 (I187763,I3563,I187545,I187513,);
not I_10835 (I187794,I187746);
not I_10836 (I187811,I578652);
nand I_10837 (I187828,I187811,I578673);
nor I_10838 (I187845,I578652,I578670);
nand I_10839 (I187525,I187661,I187845);
nand I_10840 (I187519,I187610,I578652);
nand I_10841 (I187890,I187712,I578667);
DFFARX1 I_10842 (I187890,I3563,I187545,I187534,);
DFFARX1 I_10843 (I187890,I3563,I187545,I187528,);
not I_10844 (I187935,I578667);
nor I_10845 (I187952,I187935,I578649);
and I_10846 (I187969,I187952,I578658);
or I_10847 (I187986,I187969,I578652);
DFFARX1 I_10848 (I187986,I3563,I187545,I188012,);
nand I_10849 (I188020,I188012,I187678);
nor I_10850 (I187522,I188020,I187828);
nor I_10851 (I187516,I188012,I187644);
DFFARX1 I_10852 (I188012,I3563,I187545,I188074,);
not I_10853 (I188082,I188074);
nor I_10854 (I187531,I188082,I187794);
not I_10855 (I188140,I3570);
DFFARX1 I_10856 (I1046028,I3563,I188140,I188166,);
DFFARX1 I_10857 (I188166,I3563,I188140,I188183,);
not I_10858 (I188132,I188183);
not I_10859 (I188205,I188166);
DFFARX1 I_10860 (I1046037,I3563,I188140,I188231,);
not I_10861 (I188239,I188231);
and I_10862 (I188256,I188205,I1046025);
not I_10863 (I188273,I1046016);
nand I_10864 (I188290,I188273,I1046025);
not I_10865 (I188307,I1046022);
nor I_10866 (I188324,I188307,I1046040);
nand I_10867 (I188341,I188324,I1046013);
nor I_10868 (I188358,I188341,I188290);
DFFARX1 I_10869 (I188358,I3563,I188140,I188108,);
not I_10870 (I188389,I188341);
not I_10871 (I188406,I1046040);
nand I_10872 (I188423,I188406,I1046025);
nor I_10873 (I188440,I1046040,I1046016);
nand I_10874 (I188120,I188256,I188440);
nand I_10875 (I188114,I188205,I1046040);
nand I_10876 (I188485,I188307,I1046019);
DFFARX1 I_10877 (I188485,I3563,I188140,I188129,);
DFFARX1 I_10878 (I188485,I3563,I188140,I188123,);
not I_10879 (I188530,I1046019);
nor I_10880 (I188547,I188530,I1046031);
and I_10881 (I188564,I188547,I1046013);
or I_10882 (I188581,I188564,I1046034);
DFFARX1 I_10883 (I188581,I3563,I188140,I188607,);
nand I_10884 (I188615,I188607,I188273);
nor I_10885 (I188117,I188615,I188423);
nor I_10886 (I188111,I188607,I188239);
DFFARX1 I_10887 (I188607,I3563,I188140,I188669,);
not I_10888 (I188677,I188669);
nor I_10889 (I188126,I188677,I188389);
not I_10890 (I188735,I3570);
DFFARX1 I_10891 (I767089,I3563,I188735,I188761,);
DFFARX1 I_10892 (I188761,I3563,I188735,I188778,);
not I_10893 (I188727,I188778);
not I_10894 (I188800,I188761);
DFFARX1 I_10895 (I767086,I3563,I188735,I188826,);
not I_10896 (I188834,I188826);
and I_10897 (I188851,I188800,I767092);
not I_10898 (I188868,I767077);
nand I_10899 (I188885,I188868,I767092);
not I_10900 (I188902,I767080);
nor I_10901 (I188919,I188902,I767101);
nand I_10902 (I188936,I188919,I767098);
nor I_10903 (I188953,I188936,I188885);
DFFARX1 I_10904 (I188953,I3563,I188735,I188703,);
not I_10905 (I188984,I188936);
not I_10906 (I189001,I767101);
nand I_10907 (I189018,I189001,I767092);
nor I_10908 (I189035,I767101,I767077);
nand I_10909 (I188715,I188851,I189035);
nand I_10910 (I188709,I188800,I767101);
nand I_10911 (I189080,I188902,I767077);
DFFARX1 I_10912 (I189080,I3563,I188735,I188724,);
DFFARX1 I_10913 (I189080,I3563,I188735,I188718,);
not I_10914 (I189125,I767077);
nor I_10915 (I189142,I189125,I767083);
and I_10916 (I189159,I189142,I767095);
or I_10917 (I189176,I189159,I767080);
DFFARX1 I_10918 (I189176,I3563,I188735,I189202,);
nand I_10919 (I189210,I189202,I188868);
nor I_10920 (I188712,I189210,I189018);
nor I_10921 (I188706,I189202,I188834);
DFFARX1 I_10922 (I189202,I3563,I188735,I189264,);
not I_10923 (I189272,I189264);
nor I_10924 (I188721,I189272,I188984);
not I_10925 (I189330,I3570);
DFFARX1 I_10926 (I1048345,I3563,I189330,I189356,);
DFFARX1 I_10927 (I189356,I3563,I189330,I189373,);
not I_10928 (I189322,I189373);
not I_10929 (I189395,I189356);
DFFARX1 I_10930 (I1048354,I3563,I189330,I189421,);
not I_10931 (I189429,I189421);
and I_10932 (I189446,I189395,I1048348);
not I_10933 (I189463,I1048342);
nand I_10934 (I189480,I189463,I1048348);
not I_10935 (I189497,I1048357);
nor I_10936 (I189514,I189497,I1048345);
nand I_10937 (I189531,I189514,I1048351);
nor I_10938 (I189548,I189531,I189480);
DFFARX1 I_10939 (I189548,I3563,I189330,I189298,);
not I_10940 (I189579,I189531);
not I_10941 (I189596,I1048345);
nand I_10942 (I189613,I189596,I1048348);
nor I_10943 (I189630,I1048345,I1048342);
nand I_10944 (I189310,I189446,I189630);
nand I_10945 (I189304,I189395,I1048345);
nand I_10946 (I189675,I189497,I1048348);
DFFARX1 I_10947 (I189675,I3563,I189330,I189319,);
DFFARX1 I_10948 (I189675,I3563,I189330,I189313,);
not I_10949 (I189720,I1048348);
nor I_10950 (I189737,I189720,I1048363);
and I_10951 (I189754,I189737,I1048360);
or I_10952 (I189771,I189754,I1048342);
DFFARX1 I_10953 (I189771,I3563,I189330,I189797,);
nand I_10954 (I189805,I189797,I189463);
nor I_10955 (I189307,I189805,I189613);
nor I_10956 (I189301,I189797,I189429);
DFFARX1 I_10957 (I189797,I3563,I189330,I189859,);
not I_10958 (I189867,I189859);
nor I_10959 (I189316,I189867,I189579);
not I_10960 (I189925,I3570);
DFFARX1 I_10961 (I671719,I3563,I189925,I189951,);
DFFARX1 I_10962 (I189951,I3563,I189925,I189968,);
not I_10963 (I189917,I189968);
not I_10964 (I189990,I189951);
DFFARX1 I_10965 (I671716,I3563,I189925,I190016,);
not I_10966 (I190024,I190016);
and I_10967 (I190041,I189990,I671722);
not I_10968 (I190058,I671707);
nand I_10969 (I190075,I190058,I671722);
not I_10970 (I190092,I671710);
nor I_10971 (I190109,I190092,I671731);
nand I_10972 (I190126,I190109,I671728);
nor I_10973 (I190143,I190126,I190075);
DFFARX1 I_10974 (I190143,I3563,I189925,I189893,);
not I_10975 (I190174,I190126);
not I_10976 (I190191,I671731);
nand I_10977 (I190208,I190191,I671722);
nor I_10978 (I190225,I671731,I671707);
nand I_10979 (I189905,I190041,I190225);
nand I_10980 (I189899,I189990,I671731);
nand I_10981 (I190270,I190092,I671707);
DFFARX1 I_10982 (I190270,I3563,I189925,I189914,);
DFFARX1 I_10983 (I190270,I3563,I189925,I189908,);
not I_10984 (I190315,I671707);
nor I_10985 (I190332,I190315,I671713);
and I_10986 (I190349,I190332,I671725);
or I_10987 (I190366,I190349,I671710);
DFFARX1 I_10988 (I190366,I3563,I189925,I190392,);
nand I_10989 (I190400,I190392,I190058);
nor I_10990 (I189902,I190400,I190208);
nor I_10991 (I189896,I190392,I190024);
DFFARX1 I_10992 (I190392,I3563,I189925,I190454,);
not I_10993 (I190462,I190454);
nor I_10994 (I189911,I190462,I190174);
not I_10995 (I190520,I3570);
DFFARX1 I_10996 (I634152,I3563,I190520,I190546,);
DFFARX1 I_10997 (I190546,I3563,I190520,I190563,);
not I_10998 (I190512,I190563);
not I_10999 (I190585,I190546);
DFFARX1 I_11000 (I634143,I3563,I190520,I190611,);
not I_11001 (I190619,I190611);
and I_11002 (I190636,I190585,I634161);
not I_11003 (I190653,I634158);
nand I_11004 (I190670,I190653,I634161);
not I_11005 (I190687,I634137);
nor I_11006 (I190704,I190687,I634140);
nand I_11007 (I190721,I190704,I634149);
nor I_11008 (I190738,I190721,I190670);
DFFARX1 I_11009 (I190738,I3563,I190520,I190488,);
not I_11010 (I190769,I190721);
not I_11011 (I190786,I634140);
nand I_11012 (I190803,I190786,I634161);
nor I_11013 (I190820,I634140,I634158);
nand I_11014 (I190500,I190636,I190820);
nand I_11015 (I190494,I190585,I634140);
nand I_11016 (I190865,I190687,I634155);
DFFARX1 I_11017 (I190865,I3563,I190520,I190509,);
DFFARX1 I_11018 (I190865,I3563,I190520,I190503,);
not I_11019 (I190910,I634155);
nor I_11020 (I190927,I190910,I634137);
and I_11021 (I190944,I190927,I634146);
or I_11022 (I190961,I190944,I634140);
DFFARX1 I_11023 (I190961,I3563,I190520,I190987,);
nand I_11024 (I190995,I190987,I190653);
nor I_11025 (I190497,I190995,I190803);
nor I_11026 (I190491,I190987,I190619);
DFFARX1 I_11027 (I190987,I3563,I190520,I191049,);
not I_11028 (I191057,I191049);
nor I_11029 (I190506,I191057,I190769);
not I_11030 (I191115,I3570);
DFFARX1 I_11031 (I1276347,I3563,I191115,I191141,);
DFFARX1 I_11032 (I191141,I3563,I191115,I191158,);
not I_11033 (I191107,I191158);
not I_11034 (I191180,I191141);
DFFARX1 I_11035 (I1276332,I3563,I191115,I191206,);
not I_11036 (I191214,I191206);
and I_11037 (I191231,I191180,I1276350);
not I_11038 (I191248,I1276332);
nand I_11039 (I191265,I191248,I1276350);
not I_11040 (I191282,I1276353);
nor I_11041 (I191299,I191282,I1276344);
nand I_11042 (I191316,I191299,I1276341);
nor I_11043 (I191333,I191316,I191265);
DFFARX1 I_11044 (I191333,I3563,I191115,I191083,);
not I_11045 (I191364,I191316);
not I_11046 (I191381,I1276344);
nand I_11047 (I191398,I191381,I1276350);
nor I_11048 (I191415,I1276344,I1276332);
nand I_11049 (I191095,I191231,I191415);
nand I_11050 (I191089,I191180,I1276344);
nand I_11051 (I191460,I191282,I1276338);
DFFARX1 I_11052 (I191460,I3563,I191115,I191104,);
DFFARX1 I_11053 (I191460,I3563,I191115,I191098,);
not I_11054 (I191505,I1276338);
nor I_11055 (I191522,I191505,I1276329);
and I_11056 (I191539,I191522,I1276335);
or I_11057 (I191556,I191539,I1276329);
DFFARX1 I_11058 (I191556,I3563,I191115,I191582,);
nand I_11059 (I191590,I191582,I191248);
nor I_11060 (I191092,I191590,I191398);
nor I_11061 (I191086,I191582,I191214);
DFFARX1 I_11062 (I191582,I3563,I191115,I191644,);
not I_11063 (I191652,I191644);
nor I_11064 (I191101,I191652,I191364);
not I_11065 (I191710,I3570);
DFFARX1 I_11066 (I356510,I3563,I191710,I191736,);
DFFARX1 I_11067 (I191736,I3563,I191710,I191753,);
not I_11068 (I191702,I191753);
not I_11069 (I191775,I191736);
DFFARX1 I_11070 (I356525,I3563,I191710,I191801,);
not I_11071 (I191809,I191801);
and I_11072 (I191826,I191775,I356522);
not I_11073 (I191843,I356510);
nand I_11074 (I191860,I191843,I356522);
not I_11075 (I191877,I356519);
nor I_11076 (I191894,I191877,I356534);
nand I_11077 (I191911,I191894,I356531);
nor I_11078 (I191928,I191911,I191860);
DFFARX1 I_11079 (I191928,I3563,I191710,I191678,);
not I_11080 (I191959,I191911);
not I_11081 (I191976,I356534);
nand I_11082 (I191993,I191976,I356522);
nor I_11083 (I192010,I356534,I356510);
nand I_11084 (I191690,I191826,I192010);
nand I_11085 (I191684,I191775,I356534);
nand I_11086 (I192055,I191877,I356528);
DFFARX1 I_11087 (I192055,I3563,I191710,I191699,);
DFFARX1 I_11088 (I192055,I3563,I191710,I191693,);
not I_11089 (I192100,I356528);
nor I_11090 (I192117,I192100,I356516);
and I_11091 (I192134,I192117,I356537);
or I_11092 (I192151,I192134,I356513);
DFFARX1 I_11093 (I192151,I3563,I191710,I192177,);
nand I_11094 (I192185,I192177,I191843);
nor I_11095 (I191687,I192185,I191993);
nor I_11096 (I191681,I192177,I191809);
DFFARX1 I_11097 (I192177,I3563,I191710,I192239,);
not I_11098 (I192247,I192239);
nor I_11099 (I191696,I192247,I191959);
not I_11100 (I192305,I3570);
DFFARX1 I_11101 (I649180,I3563,I192305,I192331,);
DFFARX1 I_11102 (I192331,I3563,I192305,I192348,);
not I_11103 (I192297,I192348);
not I_11104 (I192370,I192331);
DFFARX1 I_11105 (I649171,I3563,I192305,I192396,);
not I_11106 (I192404,I192396);
and I_11107 (I192421,I192370,I649189);
not I_11108 (I192438,I649186);
nand I_11109 (I192455,I192438,I649189);
not I_11110 (I192472,I649165);
nor I_11111 (I192489,I192472,I649168);
nand I_11112 (I192506,I192489,I649177);
nor I_11113 (I192523,I192506,I192455);
DFFARX1 I_11114 (I192523,I3563,I192305,I192273,);
not I_11115 (I192554,I192506);
not I_11116 (I192571,I649168);
nand I_11117 (I192588,I192571,I649189);
nor I_11118 (I192605,I649168,I649186);
nand I_11119 (I192285,I192421,I192605);
nand I_11120 (I192279,I192370,I649168);
nand I_11121 (I192650,I192472,I649183);
DFFARX1 I_11122 (I192650,I3563,I192305,I192294,);
DFFARX1 I_11123 (I192650,I3563,I192305,I192288,);
not I_11124 (I192695,I649183);
nor I_11125 (I192712,I192695,I649165);
and I_11126 (I192729,I192712,I649174);
or I_11127 (I192746,I192729,I649168);
DFFARX1 I_11128 (I192746,I3563,I192305,I192772,);
nand I_11129 (I192780,I192772,I192438);
nor I_11130 (I192282,I192780,I192588);
nor I_11131 (I192276,I192772,I192404);
DFFARX1 I_11132 (I192772,I3563,I192305,I192834,);
not I_11133 (I192842,I192834);
nor I_11134 (I192291,I192842,I192554);
not I_11135 (I192900,I3570);
DFFARX1 I_11136 (I77209,I3563,I192900,I192926,);
DFFARX1 I_11137 (I192926,I3563,I192900,I192943,);
not I_11138 (I192892,I192943);
not I_11139 (I192965,I192926);
DFFARX1 I_11140 (I77203,I3563,I192900,I192991,);
not I_11141 (I192999,I192991);
and I_11142 (I193016,I192965,I77200);
not I_11143 (I193033,I77221);
nand I_11144 (I193050,I193033,I77200);
not I_11145 (I193067,I77215);
nor I_11146 (I193084,I193067,I77206);
nand I_11147 (I193101,I193084,I77212);
nor I_11148 (I193118,I193101,I193050);
DFFARX1 I_11149 (I193118,I3563,I192900,I192868,);
not I_11150 (I193149,I193101);
not I_11151 (I193166,I77206);
nand I_11152 (I193183,I193166,I77200);
nor I_11153 (I193200,I77206,I77221);
nand I_11154 (I192880,I193016,I193200);
nand I_11155 (I192874,I192965,I77206);
nand I_11156 (I193245,I193067,I77200);
DFFARX1 I_11157 (I193245,I3563,I192900,I192889,);
DFFARX1 I_11158 (I193245,I3563,I192900,I192883,);
not I_11159 (I193290,I77200);
nor I_11160 (I193307,I193290,I77218);
and I_11161 (I193324,I193307,I77224);
or I_11162 (I193341,I193324,I77203);
DFFARX1 I_11163 (I193341,I3563,I192900,I193367,);
nand I_11164 (I193375,I193367,I193033);
nor I_11165 (I192877,I193375,I193183);
nor I_11166 (I192871,I193367,I192999);
DFFARX1 I_11167 (I193367,I3563,I192900,I193429,);
not I_11168 (I193437,I193429);
nor I_11169 (I192886,I193437,I193149);
not I_11170 (I193495,I3570);
DFFARX1 I_11171 (I113572,I3563,I193495,I193521,);
DFFARX1 I_11172 (I193521,I3563,I193495,I193538,);
not I_11173 (I193487,I193538);
not I_11174 (I193560,I193521);
DFFARX1 I_11175 (I113566,I3563,I193495,I193586,);
not I_11176 (I193594,I193586);
and I_11177 (I193611,I193560,I113563);
not I_11178 (I193628,I113584);
nand I_11179 (I193645,I193628,I113563);
not I_11180 (I193662,I113578);
nor I_11181 (I193679,I193662,I113569);
nand I_11182 (I193696,I193679,I113575);
nor I_11183 (I193713,I193696,I193645);
DFFARX1 I_11184 (I193713,I3563,I193495,I193463,);
not I_11185 (I193744,I193696);
not I_11186 (I193761,I113569);
nand I_11187 (I193778,I193761,I113563);
nor I_11188 (I193795,I113569,I113584);
nand I_11189 (I193475,I193611,I193795);
nand I_11190 (I193469,I193560,I113569);
nand I_11191 (I193840,I193662,I113563);
DFFARX1 I_11192 (I193840,I3563,I193495,I193484,);
DFFARX1 I_11193 (I193840,I3563,I193495,I193478,);
not I_11194 (I193885,I113563);
nor I_11195 (I193902,I193885,I113581);
and I_11196 (I193919,I193902,I113587);
or I_11197 (I193936,I193919,I113566);
DFFARX1 I_11198 (I193936,I3563,I193495,I193962,);
nand I_11199 (I193970,I193962,I193628);
nor I_11200 (I193472,I193970,I193778);
nor I_11201 (I193466,I193962,I193594);
DFFARX1 I_11202 (I193962,I3563,I193495,I194024,);
not I_11203 (I194032,I194024);
nor I_11204 (I193481,I194032,I193744);
not I_11205 (I194090,I3570);
DFFARX1 I_11206 (I1122785,I3563,I194090,I194116,);
DFFARX1 I_11207 (I194116,I3563,I194090,I194133,);
not I_11208 (I194082,I194133);
not I_11209 (I194155,I194116);
DFFARX1 I_11210 (I1122785,I3563,I194090,I194181,);
not I_11211 (I194189,I194181);
and I_11212 (I194206,I194155,I1122788);
not I_11213 (I194223,I1122800);
nand I_11214 (I194240,I194223,I1122788);
not I_11215 (I194257,I1122806);
nor I_11216 (I194274,I194257,I1122797);
nand I_11217 (I194291,I194274,I1122803);
nor I_11218 (I194308,I194291,I194240);
DFFARX1 I_11219 (I194308,I3563,I194090,I194058,);
not I_11220 (I194339,I194291);
not I_11221 (I194356,I1122797);
nand I_11222 (I194373,I194356,I1122788);
nor I_11223 (I194390,I1122797,I1122800);
nand I_11224 (I194070,I194206,I194390);
nand I_11225 (I194064,I194155,I1122797);
nand I_11226 (I194435,I194257,I1122794);
DFFARX1 I_11227 (I194435,I3563,I194090,I194079,);
DFFARX1 I_11228 (I194435,I3563,I194090,I194073,);
not I_11229 (I194480,I1122794);
nor I_11230 (I194497,I194480,I1122791);
and I_11231 (I194514,I194497,I1122809);
or I_11232 (I194531,I194514,I1122788);
DFFARX1 I_11233 (I194531,I3563,I194090,I194557,);
nand I_11234 (I194565,I194557,I194223);
nor I_11235 (I194067,I194565,I194373);
nor I_11236 (I194061,I194557,I194189);
DFFARX1 I_11237 (I194557,I3563,I194090,I194619,);
not I_11238 (I194627,I194619);
nor I_11239 (I194076,I194627,I194339);
not I_11240 (I194685,I3570);
DFFARX1 I_11241 (I661315,I3563,I194685,I194711,);
DFFARX1 I_11242 (I194711,I3563,I194685,I194728,);
not I_11243 (I194677,I194728);
not I_11244 (I194750,I194711);
DFFARX1 I_11245 (I661312,I3563,I194685,I194776,);
not I_11246 (I194784,I194776);
and I_11247 (I194801,I194750,I661318);
not I_11248 (I194818,I661303);
nand I_11249 (I194835,I194818,I661318);
not I_11250 (I194852,I661306);
nor I_11251 (I194869,I194852,I661327);
nand I_11252 (I194886,I194869,I661324);
nor I_11253 (I194903,I194886,I194835);
DFFARX1 I_11254 (I194903,I3563,I194685,I194653,);
not I_11255 (I194934,I194886);
not I_11256 (I194951,I661327);
nand I_11257 (I194968,I194951,I661318);
nor I_11258 (I194985,I661327,I661303);
nand I_11259 (I194665,I194801,I194985);
nand I_11260 (I194659,I194750,I661327);
nand I_11261 (I195030,I194852,I661303);
DFFARX1 I_11262 (I195030,I3563,I194685,I194674,);
DFFARX1 I_11263 (I195030,I3563,I194685,I194668,);
not I_11264 (I195075,I661303);
nor I_11265 (I195092,I195075,I661309);
and I_11266 (I195109,I195092,I661321);
or I_11267 (I195126,I195109,I661306);
DFFARX1 I_11268 (I195126,I3563,I194685,I195152,);
nand I_11269 (I195160,I195152,I194818);
nor I_11270 (I194662,I195160,I194968);
nor I_11271 (I194656,I195152,I194784);
DFFARX1 I_11272 (I195152,I3563,I194685,I195214,);
not I_11273 (I195222,I195214);
nor I_11274 (I194671,I195222,I194934);
not I_11275 (I195280,I3570);
DFFARX1 I_11276 (I675765,I3563,I195280,I195306,);
DFFARX1 I_11277 (I195306,I3563,I195280,I195323,);
not I_11278 (I195272,I195323);
not I_11279 (I195345,I195306);
DFFARX1 I_11280 (I675762,I3563,I195280,I195371,);
not I_11281 (I195379,I195371);
and I_11282 (I195396,I195345,I675768);
not I_11283 (I195413,I675753);
nand I_11284 (I195430,I195413,I675768);
not I_11285 (I195447,I675756);
nor I_11286 (I195464,I195447,I675777);
nand I_11287 (I195481,I195464,I675774);
nor I_11288 (I195498,I195481,I195430);
DFFARX1 I_11289 (I195498,I3563,I195280,I195248,);
not I_11290 (I195529,I195481);
not I_11291 (I195546,I675777);
nand I_11292 (I195563,I195546,I675768);
nor I_11293 (I195580,I675777,I675753);
nand I_11294 (I195260,I195396,I195580);
nand I_11295 (I195254,I195345,I675777);
nand I_11296 (I195625,I195447,I675753);
DFFARX1 I_11297 (I195625,I3563,I195280,I195269,);
DFFARX1 I_11298 (I195625,I3563,I195280,I195263,);
not I_11299 (I195670,I675753);
nor I_11300 (I195687,I195670,I675759);
and I_11301 (I195704,I195687,I675771);
or I_11302 (I195721,I195704,I675756);
DFFARX1 I_11303 (I195721,I3563,I195280,I195747,);
nand I_11304 (I195755,I195747,I195413);
nor I_11305 (I195257,I195755,I195563);
nor I_11306 (I195251,I195747,I195379);
DFFARX1 I_11307 (I195747,I3563,I195280,I195809,);
not I_11308 (I195817,I195809);
nor I_11309 (I195266,I195817,I195529);
not I_11310 (I195875,I3570);
DFFARX1 I_11311 (I435482,I3563,I195875,I195901,);
DFFARX1 I_11312 (I195901,I3563,I195875,I195918,);
not I_11313 (I195867,I195918);
not I_11314 (I195940,I195901);
DFFARX1 I_11315 (I435470,I3563,I195875,I195966,);
not I_11316 (I195974,I195966);
and I_11317 (I195991,I195940,I435479);
not I_11318 (I196008,I435476);
nand I_11319 (I196025,I196008,I435479);
not I_11320 (I196042,I435467);
nor I_11321 (I196059,I196042,I435473);
nand I_11322 (I196076,I196059,I435458);
nor I_11323 (I196093,I196076,I196025);
DFFARX1 I_11324 (I196093,I3563,I195875,I195843,);
not I_11325 (I196124,I196076);
not I_11326 (I196141,I435473);
nand I_11327 (I196158,I196141,I435479);
nor I_11328 (I196175,I435473,I435476);
nand I_11329 (I195855,I195991,I196175);
nand I_11330 (I195849,I195940,I435473);
nand I_11331 (I196220,I196042,I435458);
DFFARX1 I_11332 (I196220,I3563,I195875,I195864,);
DFFARX1 I_11333 (I196220,I3563,I195875,I195858,);
not I_11334 (I196265,I435458);
nor I_11335 (I196282,I196265,I435464);
and I_11336 (I196299,I196282,I435461);
or I_11337 (I196316,I196299,I435485);
DFFARX1 I_11338 (I196316,I3563,I195875,I196342,);
nand I_11339 (I196350,I196342,I196008);
nor I_11340 (I195852,I196350,I196158);
nor I_11341 (I195846,I196342,I195974);
DFFARX1 I_11342 (I196342,I3563,I195875,I196404,);
not I_11343 (I196412,I196404);
nor I_11344 (I195861,I196412,I196124);
not I_11345 (I196470,I3570);
DFFARX1 I_11346 (I865343,I3563,I196470,I196496,);
DFFARX1 I_11347 (I196496,I3563,I196470,I196513,);
not I_11348 (I196462,I196513);
not I_11349 (I196535,I196496);
DFFARX1 I_11350 (I865337,I3563,I196470,I196561,);
not I_11351 (I196569,I196561);
and I_11352 (I196586,I196535,I865355);
not I_11353 (I196603,I865343);
nand I_11354 (I196620,I196603,I865355);
not I_11355 (I196637,I865337);
nor I_11356 (I196654,I196637,I865349);
nand I_11357 (I196671,I196654,I865340);
nor I_11358 (I196688,I196671,I196620);
DFFARX1 I_11359 (I196688,I3563,I196470,I196438,);
not I_11360 (I196719,I196671);
not I_11361 (I196736,I865349);
nand I_11362 (I196753,I196736,I865355);
nor I_11363 (I196770,I865349,I865343);
nand I_11364 (I196450,I196586,I196770);
nand I_11365 (I196444,I196535,I865349);
nand I_11366 (I196815,I196637,I865352);
DFFARX1 I_11367 (I196815,I3563,I196470,I196459,);
DFFARX1 I_11368 (I196815,I3563,I196470,I196453,);
not I_11369 (I196860,I865352);
nor I_11370 (I196877,I196860,I865358);
and I_11371 (I196894,I196877,I865340);
or I_11372 (I196911,I196894,I865346);
DFFARX1 I_11373 (I196911,I3563,I196470,I196937,);
nand I_11374 (I196945,I196937,I196603);
nor I_11375 (I196447,I196945,I196753);
nor I_11376 (I196441,I196937,I196569);
DFFARX1 I_11377 (I196937,I3563,I196470,I196999,);
not I_11378 (I197007,I196999);
nor I_11379 (I196456,I197007,I196719);
not I_11380 (I197065,I3570);
DFFARX1 I_11381 (I1301050,I3563,I197065,I197091,);
DFFARX1 I_11382 (I197091,I3563,I197065,I197108,);
not I_11383 (I197057,I197108);
not I_11384 (I197130,I197091);
DFFARX1 I_11385 (I1301062,I3563,I197065,I197156,);
not I_11386 (I197164,I197156);
and I_11387 (I197181,I197130,I1301056);
not I_11388 (I197198,I1301068);
nand I_11389 (I197215,I197198,I1301056);
not I_11390 (I197232,I1301053);
nor I_11391 (I197249,I197232,I1301065);
nand I_11392 (I197266,I197249,I1301047);
nor I_11393 (I197283,I197266,I197215);
DFFARX1 I_11394 (I197283,I3563,I197065,I197033,);
not I_11395 (I197314,I197266);
not I_11396 (I197331,I1301065);
nand I_11397 (I197348,I197331,I1301056);
nor I_11398 (I197365,I1301065,I1301068);
nand I_11399 (I197045,I197181,I197365);
nand I_11400 (I197039,I197130,I1301065);
nand I_11401 (I197410,I197232,I1301059);
DFFARX1 I_11402 (I197410,I3563,I197065,I197054,);
DFFARX1 I_11403 (I197410,I3563,I197065,I197048,);
not I_11404 (I197455,I1301059);
nor I_11405 (I197472,I197455,I1301050);
and I_11406 (I197489,I197472,I1301047);
or I_11407 (I197506,I197489,I1301071);
DFFARX1 I_11408 (I197506,I3563,I197065,I197532,);
nand I_11409 (I197540,I197532,I197198);
nor I_11410 (I197042,I197540,I197348);
nor I_11411 (I197036,I197532,I197164);
DFFARX1 I_11412 (I197532,I3563,I197065,I197594,);
not I_11413 (I197602,I197594);
nor I_11414 (I197051,I197602,I197314);
not I_11415 (I197660,I3570);
DFFARX1 I_11416 (I660159,I3563,I197660,I197686,);
DFFARX1 I_11417 (I197686,I3563,I197660,I197703,);
not I_11418 (I197652,I197703);
not I_11419 (I197725,I197686);
DFFARX1 I_11420 (I660156,I3563,I197660,I197751,);
not I_11421 (I197759,I197751);
and I_11422 (I197776,I197725,I660162);
not I_11423 (I197793,I660147);
nand I_11424 (I197810,I197793,I660162);
not I_11425 (I197827,I660150);
nor I_11426 (I197844,I197827,I660171);
nand I_11427 (I197861,I197844,I660168);
nor I_11428 (I197878,I197861,I197810);
DFFARX1 I_11429 (I197878,I3563,I197660,I197628,);
not I_11430 (I197909,I197861);
not I_11431 (I197926,I660171);
nand I_11432 (I197943,I197926,I660162);
nor I_11433 (I197960,I660171,I660147);
nand I_11434 (I197640,I197776,I197960);
nand I_11435 (I197634,I197725,I660171);
nand I_11436 (I198005,I197827,I660147);
DFFARX1 I_11437 (I198005,I3563,I197660,I197649,);
DFFARX1 I_11438 (I198005,I3563,I197660,I197643,);
not I_11439 (I198050,I660147);
nor I_11440 (I198067,I198050,I660153);
and I_11441 (I198084,I198067,I660165);
or I_11442 (I198101,I198084,I660150);
DFFARX1 I_11443 (I198101,I3563,I197660,I198127,);
nand I_11444 (I198135,I198127,I197793);
nor I_11445 (I197637,I198135,I197943);
nor I_11446 (I197631,I198127,I197759);
DFFARX1 I_11447 (I198127,I3563,I197660,I198189,);
not I_11448 (I198197,I198189);
nor I_11449 (I197646,I198197,I197909);
not I_11450 (I198255,I3570);
DFFARX1 I_11451 (I1129143,I3563,I198255,I198281,);
DFFARX1 I_11452 (I198281,I3563,I198255,I198298,);
not I_11453 (I198247,I198298);
not I_11454 (I198320,I198281);
DFFARX1 I_11455 (I1129143,I3563,I198255,I198346,);
not I_11456 (I198354,I198346);
and I_11457 (I198371,I198320,I1129146);
not I_11458 (I198388,I1129158);
nand I_11459 (I198405,I198388,I1129146);
not I_11460 (I198422,I1129164);
nor I_11461 (I198439,I198422,I1129155);
nand I_11462 (I198456,I198439,I1129161);
nor I_11463 (I198473,I198456,I198405);
DFFARX1 I_11464 (I198473,I3563,I198255,I198223,);
not I_11465 (I198504,I198456);
not I_11466 (I198521,I1129155);
nand I_11467 (I198538,I198521,I1129146);
nor I_11468 (I198555,I1129155,I1129158);
nand I_11469 (I198235,I198371,I198555);
nand I_11470 (I198229,I198320,I1129155);
nand I_11471 (I198600,I198422,I1129152);
DFFARX1 I_11472 (I198600,I3563,I198255,I198244,);
DFFARX1 I_11473 (I198600,I3563,I198255,I198238,);
not I_11474 (I198645,I1129152);
nor I_11475 (I198662,I198645,I1129149);
and I_11476 (I198679,I198662,I1129167);
or I_11477 (I198696,I198679,I1129146);
DFFARX1 I_11478 (I198696,I3563,I198255,I198722,);
nand I_11479 (I198730,I198722,I198388);
nor I_11480 (I198232,I198730,I198538);
nor I_11481 (I198226,I198722,I198354);
DFFARX1 I_11482 (I198722,I3563,I198255,I198784,);
not I_11483 (I198792,I198784);
nor I_11484 (I198241,I198792,I198504);
not I_11485 (I198850,I3570);
DFFARX1 I_11486 (I1372604,I3563,I198850,I198876,);
DFFARX1 I_11487 (I198876,I3563,I198850,I198893,);
not I_11488 (I198842,I198893);
not I_11489 (I198915,I198876);
DFFARX1 I_11490 (I1372595,I3563,I198850,I198941,);
not I_11491 (I198949,I198941);
and I_11492 (I198966,I198915,I1372589);
not I_11493 (I198983,I1372583);
nand I_11494 (I199000,I198983,I1372589);
not I_11495 (I199017,I1372610);
nor I_11496 (I199034,I199017,I1372583);
nand I_11497 (I199051,I199034,I1372607);
nor I_11498 (I199068,I199051,I199000);
DFFARX1 I_11499 (I199068,I3563,I198850,I198818,);
not I_11500 (I199099,I199051);
not I_11501 (I199116,I1372583);
nand I_11502 (I199133,I199116,I1372589);
nor I_11503 (I199150,I1372583,I1372583);
nand I_11504 (I198830,I198966,I199150);
nand I_11505 (I198824,I198915,I1372583);
nand I_11506 (I199195,I199017,I1372592);
DFFARX1 I_11507 (I199195,I3563,I198850,I198839,);
DFFARX1 I_11508 (I199195,I3563,I198850,I198833,);
not I_11509 (I199240,I1372592);
nor I_11510 (I199257,I199240,I1372598);
and I_11511 (I199274,I199257,I1372601);
or I_11512 (I199291,I199274,I1372586);
DFFARX1 I_11513 (I199291,I3563,I198850,I199317,);
nand I_11514 (I199325,I199317,I198983);
nor I_11515 (I198827,I199325,I199133);
nor I_11516 (I198821,I199317,I198949);
DFFARX1 I_11517 (I199317,I3563,I198850,I199379,);
not I_11518 (I199387,I199379);
nor I_11519 (I198836,I199387,I199099);
not I_11520 (I199445,I3570);
DFFARX1 I_11521 (I551903,I3563,I199445,I199471,);
DFFARX1 I_11522 (I199471,I3563,I199445,I199488,);
not I_11523 (I199437,I199488);
not I_11524 (I199510,I199471);
DFFARX1 I_11525 (I551897,I3563,I199445,I199536,);
not I_11526 (I199544,I199536);
and I_11527 (I199561,I199510,I551912);
not I_11528 (I199578,I551909);
nand I_11529 (I199595,I199578,I551912);
not I_11530 (I199612,I551900);
nor I_11531 (I199629,I199612,I551891);
nand I_11532 (I199646,I199629,I551894);
nor I_11533 (I199663,I199646,I199595);
DFFARX1 I_11534 (I199663,I3563,I199445,I199413,);
not I_11535 (I199694,I199646);
not I_11536 (I199711,I551891);
nand I_11537 (I199728,I199711,I551912);
nor I_11538 (I199745,I551891,I551909);
nand I_11539 (I199425,I199561,I199745);
nand I_11540 (I199419,I199510,I551891);
nand I_11541 (I199790,I199612,I551915);
DFFARX1 I_11542 (I199790,I3563,I199445,I199434,);
DFFARX1 I_11543 (I199790,I3563,I199445,I199428,);
not I_11544 (I199835,I551915);
nor I_11545 (I199852,I199835,I551906);
and I_11546 (I199869,I199852,I551891);
or I_11547 (I199886,I199869,I551894);
DFFARX1 I_11548 (I199886,I3563,I199445,I199912,);
nand I_11549 (I199920,I199912,I199578);
nor I_11550 (I199422,I199920,I199728);
nor I_11551 (I199416,I199912,I199544);
DFFARX1 I_11552 (I199912,I3563,I199445,I199974,);
not I_11553 (I199982,I199974);
nor I_11554 (I199431,I199982,I199694);
not I_11555 (I200040,I3570);
DFFARX1 I_11556 (I122004,I3563,I200040,I200066,);
DFFARX1 I_11557 (I200066,I3563,I200040,I200083,);
not I_11558 (I200032,I200083);
not I_11559 (I200105,I200066);
DFFARX1 I_11560 (I121998,I3563,I200040,I200131,);
not I_11561 (I200139,I200131);
and I_11562 (I200156,I200105,I121995);
not I_11563 (I200173,I122016);
nand I_11564 (I200190,I200173,I121995);
not I_11565 (I200207,I122010);
nor I_11566 (I200224,I200207,I122001);
nand I_11567 (I200241,I200224,I122007);
nor I_11568 (I200258,I200241,I200190);
DFFARX1 I_11569 (I200258,I3563,I200040,I200008,);
not I_11570 (I200289,I200241);
not I_11571 (I200306,I122001);
nand I_11572 (I200323,I200306,I121995);
nor I_11573 (I200340,I122001,I122016);
nand I_11574 (I200020,I200156,I200340);
nand I_11575 (I200014,I200105,I122001);
nand I_11576 (I200385,I200207,I121995);
DFFARX1 I_11577 (I200385,I3563,I200040,I200029,);
DFFARX1 I_11578 (I200385,I3563,I200040,I200023,);
not I_11579 (I200430,I121995);
nor I_11580 (I200447,I200430,I122013);
and I_11581 (I200464,I200447,I122019);
or I_11582 (I200481,I200464,I121998);
DFFARX1 I_11583 (I200481,I3563,I200040,I200507,);
nand I_11584 (I200515,I200507,I200173);
nor I_11585 (I200017,I200515,I200323);
nor I_11586 (I200011,I200507,I200139);
DFFARX1 I_11587 (I200507,I3563,I200040,I200569,);
not I_11588 (I200577,I200569);
nor I_11589 (I200026,I200577,I200289);
not I_11590 (I200635,I3570);
DFFARX1 I_11591 (I125693,I3563,I200635,I200661,);
DFFARX1 I_11592 (I200661,I3563,I200635,I200678,);
not I_11593 (I200627,I200678);
not I_11594 (I200700,I200661);
DFFARX1 I_11595 (I125687,I3563,I200635,I200726,);
not I_11596 (I200734,I200726);
and I_11597 (I200751,I200700,I125684);
not I_11598 (I200768,I125705);
nand I_11599 (I200785,I200768,I125684);
not I_11600 (I200802,I125699);
nor I_11601 (I200819,I200802,I125690);
nand I_11602 (I200836,I200819,I125696);
nor I_11603 (I200853,I200836,I200785);
DFFARX1 I_11604 (I200853,I3563,I200635,I200603,);
not I_11605 (I200884,I200836);
not I_11606 (I200901,I125690);
nand I_11607 (I200918,I200901,I125684);
nor I_11608 (I200935,I125690,I125705);
nand I_11609 (I200615,I200751,I200935);
nand I_11610 (I200609,I200700,I125690);
nand I_11611 (I200980,I200802,I125684);
DFFARX1 I_11612 (I200980,I3563,I200635,I200624,);
DFFARX1 I_11613 (I200980,I3563,I200635,I200618,);
not I_11614 (I201025,I125684);
nor I_11615 (I201042,I201025,I125702);
and I_11616 (I201059,I201042,I125708);
or I_11617 (I201076,I201059,I125687);
DFFARX1 I_11618 (I201076,I3563,I200635,I201102,);
nand I_11619 (I201110,I201102,I200768);
nor I_11620 (I200612,I201110,I200918);
nor I_11621 (I200606,I201102,I200734);
DFFARX1 I_11622 (I201102,I3563,I200635,I201164,);
not I_11623 (I201172,I201164);
nor I_11624 (I200621,I201172,I200884);
not I_11625 (I201230,I3570);
DFFARX1 I_11626 (I611032,I3563,I201230,I201256,);
DFFARX1 I_11627 (I201256,I3563,I201230,I201273,);
not I_11628 (I201222,I201273);
not I_11629 (I201295,I201256);
DFFARX1 I_11630 (I611023,I3563,I201230,I201321,);
not I_11631 (I201329,I201321);
and I_11632 (I201346,I201295,I611041);
not I_11633 (I201363,I611038);
nand I_11634 (I201380,I201363,I611041);
not I_11635 (I201397,I611017);
nor I_11636 (I201414,I201397,I611020);
nand I_11637 (I201431,I201414,I611029);
nor I_11638 (I201448,I201431,I201380);
DFFARX1 I_11639 (I201448,I3563,I201230,I201198,);
not I_11640 (I201479,I201431);
not I_11641 (I201496,I611020);
nand I_11642 (I201513,I201496,I611041);
nor I_11643 (I201530,I611020,I611038);
nand I_11644 (I201210,I201346,I201530);
nand I_11645 (I201204,I201295,I611020);
nand I_11646 (I201575,I201397,I611035);
DFFARX1 I_11647 (I201575,I3563,I201230,I201219,);
DFFARX1 I_11648 (I201575,I3563,I201230,I201213,);
not I_11649 (I201620,I611035);
nor I_11650 (I201637,I201620,I611017);
and I_11651 (I201654,I201637,I611026);
or I_11652 (I201671,I201654,I611020);
DFFARX1 I_11653 (I201671,I3563,I201230,I201697,);
nand I_11654 (I201705,I201697,I201363);
nor I_11655 (I201207,I201705,I201513);
nor I_11656 (I201201,I201697,I201329);
DFFARX1 I_11657 (I201697,I3563,I201230,I201759,);
not I_11658 (I201767,I201759);
nor I_11659 (I201216,I201767,I201479);
not I_11660 (I201825,I3570);
DFFARX1 I_11661 (I1219889,I3563,I201825,I201851,);
DFFARX1 I_11662 (I201851,I3563,I201825,I201868,);
not I_11663 (I201817,I201868);
not I_11664 (I201890,I201851);
DFFARX1 I_11665 (I1219889,I3563,I201825,I201916,);
not I_11666 (I201924,I201916);
and I_11667 (I201941,I201890,I1219892);
not I_11668 (I201958,I1219904);
nand I_11669 (I201975,I201958,I1219892);
not I_11670 (I201992,I1219910);
nor I_11671 (I202009,I201992,I1219901);
nand I_11672 (I202026,I202009,I1219907);
nor I_11673 (I202043,I202026,I201975);
DFFARX1 I_11674 (I202043,I3563,I201825,I201793,);
not I_11675 (I202074,I202026);
not I_11676 (I202091,I1219901);
nand I_11677 (I202108,I202091,I1219892);
nor I_11678 (I202125,I1219901,I1219904);
nand I_11679 (I201805,I201941,I202125);
nand I_11680 (I201799,I201890,I1219901);
nand I_11681 (I202170,I201992,I1219898);
DFFARX1 I_11682 (I202170,I3563,I201825,I201814,);
DFFARX1 I_11683 (I202170,I3563,I201825,I201808,);
not I_11684 (I202215,I1219898);
nor I_11685 (I202232,I202215,I1219895);
and I_11686 (I202249,I202232,I1219913);
or I_11687 (I202266,I202249,I1219892);
DFFARX1 I_11688 (I202266,I3563,I201825,I202292,);
nand I_11689 (I202300,I202292,I201958);
nor I_11690 (I201802,I202300,I202108);
nor I_11691 (I201796,I202292,I201924);
DFFARX1 I_11692 (I202292,I3563,I201825,I202354,);
not I_11693 (I202362,I202354);
nor I_11694 (I201811,I202362,I202074);
not I_11695 (I202420,I3570);
DFFARX1 I_11696 (I642822,I3563,I202420,I202446,);
DFFARX1 I_11697 (I202446,I3563,I202420,I202463,);
not I_11698 (I202412,I202463);
not I_11699 (I202485,I202446);
DFFARX1 I_11700 (I642813,I3563,I202420,I202511,);
not I_11701 (I202519,I202511);
and I_11702 (I202536,I202485,I642831);
not I_11703 (I202553,I642828);
nand I_11704 (I202570,I202553,I642831);
not I_11705 (I202587,I642807);
nor I_11706 (I202604,I202587,I642810);
nand I_11707 (I202621,I202604,I642819);
nor I_11708 (I202638,I202621,I202570);
DFFARX1 I_11709 (I202638,I3563,I202420,I202388,);
not I_11710 (I202669,I202621);
not I_11711 (I202686,I642810);
nand I_11712 (I202703,I202686,I642831);
nor I_11713 (I202720,I642810,I642828);
nand I_11714 (I202400,I202536,I202720);
nand I_11715 (I202394,I202485,I642810);
nand I_11716 (I202765,I202587,I642825);
DFFARX1 I_11717 (I202765,I3563,I202420,I202409,);
DFFARX1 I_11718 (I202765,I3563,I202420,I202403,);
not I_11719 (I202810,I642825);
nor I_11720 (I202827,I202810,I642807);
and I_11721 (I202844,I202827,I642816);
or I_11722 (I202861,I202844,I642810);
DFFARX1 I_11723 (I202861,I3563,I202420,I202887,);
nand I_11724 (I202895,I202887,I202553);
nor I_11725 (I202397,I202895,I202703);
nor I_11726 (I202391,I202887,I202519);
DFFARX1 I_11727 (I202887,I3563,I202420,I202949,);
not I_11728 (I202957,I202949);
nor I_11729 (I202406,I202957,I202669);
not I_11730 (I203015,I3570);
DFFARX1 I_11731 (I736455,I3563,I203015,I203041,);
DFFARX1 I_11732 (I203041,I3563,I203015,I203058,);
not I_11733 (I203007,I203058);
not I_11734 (I203080,I203041);
DFFARX1 I_11735 (I736452,I3563,I203015,I203106,);
not I_11736 (I203114,I203106);
and I_11737 (I203131,I203080,I736458);
not I_11738 (I203148,I736443);
nand I_11739 (I203165,I203148,I736458);
not I_11740 (I203182,I736446);
nor I_11741 (I203199,I203182,I736467);
nand I_11742 (I203216,I203199,I736464);
nor I_11743 (I203233,I203216,I203165);
DFFARX1 I_11744 (I203233,I3563,I203015,I202983,);
not I_11745 (I203264,I203216);
not I_11746 (I203281,I736467);
nand I_11747 (I203298,I203281,I736458);
nor I_11748 (I203315,I736467,I736443);
nand I_11749 (I202995,I203131,I203315);
nand I_11750 (I202989,I203080,I736467);
nand I_11751 (I203360,I203182,I736443);
DFFARX1 I_11752 (I203360,I3563,I203015,I203004,);
DFFARX1 I_11753 (I203360,I3563,I203015,I202998,);
not I_11754 (I203405,I736443);
nor I_11755 (I203422,I203405,I736449);
and I_11756 (I203439,I203422,I736461);
or I_11757 (I203456,I203439,I736446);
DFFARX1 I_11758 (I203456,I3563,I203015,I203482,);
nand I_11759 (I203490,I203482,I203148);
nor I_11760 (I202992,I203490,I203298);
nor I_11761 (I202986,I203482,I203114);
DFFARX1 I_11762 (I203482,I3563,I203015,I203544,);
not I_11763 (I203552,I203544);
nor I_11764 (I203001,I203552,I203264);
not I_11765 (I203610,I3570);
DFFARX1 I_11766 (I1390454,I3563,I203610,I203636,);
DFFARX1 I_11767 (I203636,I3563,I203610,I203653,);
not I_11768 (I203602,I203653);
not I_11769 (I203675,I203636);
DFFARX1 I_11770 (I1390445,I3563,I203610,I203701,);
not I_11771 (I203709,I203701);
and I_11772 (I203726,I203675,I1390439);
not I_11773 (I203743,I1390433);
nand I_11774 (I203760,I203743,I1390439);
not I_11775 (I203777,I1390460);
nor I_11776 (I203794,I203777,I1390433);
nand I_11777 (I203811,I203794,I1390457);
nor I_11778 (I203828,I203811,I203760);
DFFARX1 I_11779 (I203828,I3563,I203610,I203578,);
not I_11780 (I203859,I203811);
not I_11781 (I203876,I1390433);
nand I_11782 (I203893,I203876,I1390439);
nor I_11783 (I203910,I1390433,I1390433);
nand I_11784 (I203590,I203726,I203910);
nand I_11785 (I203584,I203675,I1390433);
nand I_11786 (I203955,I203777,I1390442);
DFFARX1 I_11787 (I203955,I3563,I203610,I203599,);
DFFARX1 I_11788 (I203955,I3563,I203610,I203593,);
not I_11789 (I204000,I1390442);
nor I_11790 (I204017,I204000,I1390448);
and I_11791 (I204034,I204017,I1390451);
or I_11792 (I204051,I204034,I1390436);
DFFARX1 I_11793 (I204051,I3563,I203610,I204077,);
nand I_11794 (I204085,I204077,I203743);
nor I_11795 (I203587,I204085,I203893);
nor I_11796 (I203581,I204077,I203709);
DFFARX1 I_11797 (I204077,I3563,I203610,I204139,);
not I_11798 (I204147,I204139);
nor I_11799 (I203596,I204147,I203859);
not I_11800 (I204205,I3570);
DFFARX1 I_11801 (I1100243,I3563,I204205,I204231,);
DFFARX1 I_11802 (I204231,I3563,I204205,I204248,);
not I_11803 (I204197,I204248);
not I_11804 (I204270,I204231);
DFFARX1 I_11805 (I1100243,I3563,I204205,I204296,);
not I_11806 (I204304,I204296);
and I_11807 (I204321,I204270,I1100246);
not I_11808 (I204338,I1100258);
nand I_11809 (I204355,I204338,I1100246);
not I_11810 (I204372,I1100264);
nor I_11811 (I204389,I204372,I1100255);
nand I_11812 (I204406,I204389,I1100261);
nor I_11813 (I204423,I204406,I204355);
DFFARX1 I_11814 (I204423,I3563,I204205,I204173,);
not I_11815 (I204454,I204406);
not I_11816 (I204471,I1100255);
nand I_11817 (I204488,I204471,I1100246);
nor I_11818 (I204505,I1100255,I1100258);
nand I_11819 (I204185,I204321,I204505);
nand I_11820 (I204179,I204270,I1100255);
nand I_11821 (I204550,I204372,I1100252);
DFFARX1 I_11822 (I204550,I3563,I204205,I204194,);
DFFARX1 I_11823 (I204550,I3563,I204205,I204188,);
not I_11824 (I204595,I1100252);
nor I_11825 (I204612,I204595,I1100249);
and I_11826 (I204629,I204612,I1100267);
or I_11827 (I204646,I204629,I1100246);
DFFARX1 I_11828 (I204646,I3563,I204205,I204672,);
nand I_11829 (I204680,I204672,I204338);
nor I_11830 (I204182,I204680,I204488);
nor I_11831 (I204176,I204672,I204304);
DFFARX1 I_11832 (I204672,I3563,I204205,I204734,);
not I_11833 (I204742,I204734);
nor I_11834 (I204191,I204742,I204454);
not I_11835 (I204800,I3570);
DFFARX1 I_11836 (I132544,I3563,I204800,I204826,);
DFFARX1 I_11837 (I204826,I3563,I204800,I204843,);
not I_11838 (I204792,I204843);
not I_11839 (I204865,I204826);
DFFARX1 I_11840 (I132538,I3563,I204800,I204891,);
not I_11841 (I204899,I204891);
and I_11842 (I204916,I204865,I132535);
not I_11843 (I204933,I132556);
nand I_11844 (I204950,I204933,I132535);
not I_11845 (I204967,I132550);
nor I_11846 (I204984,I204967,I132541);
nand I_11847 (I205001,I204984,I132547);
nor I_11848 (I205018,I205001,I204950);
DFFARX1 I_11849 (I205018,I3563,I204800,I204768,);
not I_11850 (I205049,I205001);
not I_11851 (I205066,I132541);
nand I_11852 (I205083,I205066,I132535);
nor I_11853 (I205100,I132541,I132556);
nand I_11854 (I204780,I204916,I205100);
nand I_11855 (I204774,I204865,I132541);
nand I_11856 (I205145,I204967,I132535);
DFFARX1 I_11857 (I205145,I3563,I204800,I204789,);
DFFARX1 I_11858 (I205145,I3563,I204800,I204783,);
not I_11859 (I205190,I132535);
nor I_11860 (I205207,I205190,I132553);
and I_11861 (I205224,I205207,I132559);
or I_11862 (I205241,I205224,I132538);
DFFARX1 I_11863 (I205241,I3563,I204800,I205267,);
nand I_11864 (I205275,I205267,I204933);
nor I_11865 (I204777,I205275,I205083);
nor I_11866 (I204771,I205267,I204899);
DFFARX1 I_11867 (I205267,I3563,I204800,I205329,);
not I_11868 (I205337,I205329);
nor I_11869 (I204786,I205337,I205049);
not I_11870 (I205395,I3570);
DFFARX1 I_11871 (I541193,I3563,I205395,I205421,);
DFFARX1 I_11872 (I205421,I3563,I205395,I205438,);
not I_11873 (I205387,I205438);
not I_11874 (I205460,I205421);
DFFARX1 I_11875 (I541187,I3563,I205395,I205486,);
not I_11876 (I205494,I205486);
and I_11877 (I205511,I205460,I541202);
not I_11878 (I205528,I541199);
nand I_11879 (I205545,I205528,I541202);
not I_11880 (I205562,I541190);
nor I_11881 (I205579,I205562,I541181);
nand I_11882 (I205596,I205579,I541184);
nor I_11883 (I205613,I205596,I205545);
DFFARX1 I_11884 (I205613,I3563,I205395,I205363,);
not I_11885 (I205644,I205596);
not I_11886 (I205661,I541181);
nand I_11887 (I205678,I205661,I541202);
nor I_11888 (I205695,I541181,I541199);
nand I_11889 (I205375,I205511,I205695);
nand I_11890 (I205369,I205460,I541181);
nand I_11891 (I205740,I205562,I541205);
DFFARX1 I_11892 (I205740,I3563,I205395,I205384,);
DFFARX1 I_11893 (I205740,I3563,I205395,I205378,);
not I_11894 (I205785,I541205);
nor I_11895 (I205802,I205785,I541196);
and I_11896 (I205819,I205802,I541181);
or I_11897 (I205836,I205819,I541184);
DFFARX1 I_11898 (I205836,I3563,I205395,I205862,);
nand I_11899 (I205870,I205862,I205528);
nor I_11900 (I205372,I205870,I205678);
nor I_11901 (I205366,I205862,I205494);
DFFARX1 I_11902 (I205862,I3563,I205395,I205924,);
not I_11903 (I205932,I205924);
nor I_11904 (I205381,I205932,I205644);
not I_11905 (I205990,I3570);
DFFARX1 I_11906 (I337538,I3563,I205990,I206016,);
DFFARX1 I_11907 (I206016,I3563,I205990,I206033,);
not I_11908 (I205982,I206033);
not I_11909 (I206055,I206016);
DFFARX1 I_11910 (I337553,I3563,I205990,I206081,);
not I_11911 (I206089,I206081);
and I_11912 (I206106,I206055,I337550);
not I_11913 (I206123,I337538);
nand I_11914 (I206140,I206123,I337550);
not I_11915 (I206157,I337547);
nor I_11916 (I206174,I206157,I337562);
nand I_11917 (I206191,I206174,I337559);
nor I_11918 (I206208,I206191,I206140);
DFFARX1 I_11919 (I206208,I3563,I205990,I205958,);
not I_11920 (I206239,I206191);
not I_11921 (I206256,I337562);
nand I_11922 (I206273,I206256,I337550);
nor I_11923 (I206290,I337562,I337538);
nand I_11924 (I205970,I206106,I206290);
nand I_11925 (I205964,I206055,I337562);
nand I_11926 (I206335,I206157,I337556);
DFFARX1 I_11927 (I206335,I3563,I205990,I205979,);
DFFARX1 I_11928 (I206335,I3563,I205990,I205973,);
not I_11929 (I206380,I337556);
nor I_11930 (I206397,I206380,I337544);
and I_11931 (I206414,I206397,I337565);
or I_11932 (I206431,I206414,I337541);
DFFARX1 I_11933 (I206431,I3563,I205990,I206457,);
nand I_11934 (I206465,I206457,I206123);
nor I_11935 (I205967,I206465,I206273);
nor I_11936 (I205961,I206457,I206089);
DFFARX1 I_11937 (I206457,I3563,I205990,I206519,);
not I_11938 (I206527,I206519);
nor I_11939 (I205976,I206527,I206239);
not I_11940 (I206585,I3570);
DFFARX1 I_11941 (I1350589,I3563,I206585,I206611,);
DFFARX1 I_11942 (I206611,I3563,I206585,I206628,);
not I_11943 (I206577,I206628);
not I_11944 (I206650,I206611);
DFFARX1 I_11945 (I1350580,I3563,I206585,I206676,);
not I_11946 (I206684,I206676);
and I_11947 (I206701,I206650,I1350574);
not I_11948 (I206718,I1350568);
nand I_11949 (I206735,I206718,I1350574);
not I_11950 (I206752,I1350595);
nor I_11951 (I206769,I206752,I1350568);
nand I_11952 (I206786,I206769,I1350592);
nor I_11953 (I206803,I206786,I206735);
DFFARX1 I_11954 (I206803,I3563,I206585,I206553,);
not I_11955 (I206834,I206786);
not I_11956 (I206851,I1350568);
nand I_11957 (I206868,I206851,I1350574);
nor I_11958 (I206885,I1350568,I1350568);
nand I_11959 (I206565,I206701,I206885);
nand I_11960 (I206559,I206650,I1350568);
nand I_11961 (I206930,I206752,I1350577);
DFFARX1 I_11962 (I206930,I3563,I206585,I206574,);
DFFARX1 I_11963 (I206930,I3563,I206585,I206568,);
not I_11964 (I206975,I1350577);
nor I_11965 (I206992,I206975,I1350583);
and I_11966 (I207009,I206992,I1350586);
or I_11967 (I207026,I207009,I1350571);
DFFARX1 I_11968 (I207026,I3563,I206585,I207052,);
nand I_11969 (I207060,I207052,I206718);
nor I_11970 (I206562,I207060,I206868);
nor I_11971 (I206556,I207052,I206684);
DFFARX1 I_11972 (I207052,I3563,I206585,I207114,);
not I_11973 (I207122,I207114);
nor I_11974 (I206571,I207122,I206834);
not I_11975 (I207180,I3570);
DFFARX1 I_11976 (I1005976,I3563,I207180,I207206,);
DFFARX1 I_11977 (I207206,I3563,I207180,I207223,);
not I_11978 (I207172,I207223);
not I_11979 (I207245,I207206);
DFFARX1 I_11980 (I1005985,I3563,I207180,I207271,);
not I_11981 (I207279,I207271);
and I_11982 (I207296,I207245,I1005973);
not I_11983 (I207313,I1005964);
nand I_11984 (I207330,I207313,I1005973);
not I_11985 (I207347,I1005970);
nor I_11986 (I207364,I207347,I1005988);
nand I_11987 (I207381,I207364,I1005961);
nor I_11988 (I207398,I207381,I207330);
DFFARX1 I_11989 (I207398,I3563,I207180,I207148,);
not I_11990 (I207429,I207381);
not I_11991 (I207446,I1005988);
nand I_11992 (I207463,I207446,I1005973);
nor I_11993 (I207480,I1005988,I1005964);
nand I_11994 (I207160,I207296,I207480);
nand I_11995 (I207154,I207245,I1005988);
nand I_11996 (I207525,I207347,I1005967);
DFFARX1 I_11997 (I207525,I3563,I207180,I207169,);
DFFARX1 I_11998 (I207525,I3563,I207180,I207163,);
not I_11999 (I207570,I1005967);
nor I_12000 (I207587,I207570,I1005979);
and I_12001 (I207604,I207587,I1005961);
or I_12002 (I207621,I207604,I1005982);
DFFARX1 I_12003 (I207621,I3563,I207180,I207647,);
nand I_12004 (I207655,I207647,I207313);
nor I_12005 (I207157,I207655,I207463);
nor I_12006 (I207151,I207647,I207279);
DFFARX1 I_12007 (I207647,I3563,I207180,I207709,);
not I_12008 (I207717,I207709);
nor I_12009 (I207166,I207717,I207429);
not I_12010 (I207775,I3570);
DFFARX1 I_12011 (I889585,I3563,I207775,I207801,);
DFFARX1 I_12012 (I207801,I3563,I207775,I207818,);
not I_12013 (I207767,I207818);
not I_12014 (I207840,I207801);
DFFARX1 I_12015 (I889579,I3563,I207775,I207866,);
not I_12016 (I207874,I207866);
and I_12017 (I207891,I207840,I889597);
not I_12018 (I207908,I889585);
nand I_12019 (I207925,I207908,I889597);
not I_12020 (I207942,I889579);
nor I_12021 (I207959,I207942,I889591);
nand I_12022 (I207976,I207959,I889582);
nor I_12023 (I207993,I207976,I207925);
DFFARX1 I_12024 (I207993,I3563,I207775,I207743,);
not I_12025 (I208024,I207976);
not I_12026 (I208041,I889591);
nand I_12027 (I208058,I208041,I889597);
nor I_12028 (I208075,I889591,I889585);
nand I_12029 (I207755,I207891,I208075);
nand I_12030 (I207749,I207840,I889591);
nand I_12031 (I208120,I207942,I889594);
DFFARX1 I_12032 (I208120,I3563,I207775,I207764,);
DFFARX1 I_12033 (I208120,I3563,I207775,I207758,);
not I_12034 (I208165,I889594);
nor I_12035 (I208182,I208165,I889600);
and I_12036 (I208199,I208182,I889582);
or I_12037 (I208216,I208199,I889588);
DFFARX1 I_12038 (I208216,I3563,I207775,I208242,);
nand I_12039 (I208250,I208242,I207908);
nor I_12040 (I207752,I208250,I208058);
nor I_12041 (I207746,I208242,I207874);
DFFARX1 I_12042 (I208242,I3563,I207775,I208304,);
not I_12043 (I208312,I208304);
nor I_12044 (I207761,I208312,I208024);
not I_12045 (I208370,I3570);
DFFARX1 I_12046 (I967216,I3563,I208370,I208396,);
DFFARX1 I_12047 (I208396,I3563,I208370,I208413,);
not I_12048 (I208362,I208413);
not I_12049 (I208435,I208396);
DFFARX1 I_12050 (I967225,I3563,I208370,I208461,);
not I_12051 (I208469,I208461);
and I_12052 (I208486,I208435,I967213);
not I_12053 (I208503,I967204);
nand I_12054 (I208520,I208503,I967213);
not I_12055 (I208537,I967210);
nor I_12056 (I208554,I208537,I967228);
nand I_12057 (I208571,I208554,I967201);
nor I_12058 (I208588,I208571,I208520);
DFFARX1 I_12059 (I208588,I3563,I208370,I208338,);
not I_12060 (I208619,I208571);
not I_12061 (I208636,I967228);
nand I_12062 (I208653,I208636,I967213);
nor I_12063 (I208670,I967228,I967204);
nand I_12064 (I208350,I208486,I208670);
nand I_12065 (I208344,I208435,I967228);
nand I_12066 (I208715,I208537,I967207);
DFFARX1 I_12067 (I208715,I3563,I208370,I208359,);
DFFARX1 I_12068 (I208715,I3563,I208370,I208353,);
not I_12069 (I208760,I967207);
nor I_12070 (I208777,I208760,I967219);
and I_12071 (I208794,I208777,I967201);
or I_12072 (I208811,I208794,I967222);
DFFARX1 I_12073 (I208811,I3563,I208370,I208837,);
nand I_12074 (I208845,I208837,I208503);
nor I_12075 (I208347,I208845,I208653);
nor I_12076 (I208341,I208837,I208469);
DFFARX1 I_12077 (I208837,I3563,I208370,I208899,);
not I_12078 (I208907,I208899);
nor I_12079 (I208356,I208907,I208619);
not I_12080 (I208965,I3570);
DFFARX1 I_12081 (I306445,I3563,I208965,I208991,);
DFFARX1 I_12082 (I208991,I3563,I208965,I209008,);
not I_12083 (I208957,I209008);
not I_12084 (I209030,I208991);
DFFARX1 I_12085 (I306460,I3563,I208965,I209056,);
not I_12086 (I209064,I209056);
and I_12087 (I209081,I209030,I306457);
not I_12088 (I209098,I306445);
nand I_12089 (I209115,I209098,I306457);
not I_12090 (I209132,I306454);
nor I_12091 (I209149,I209132,I306469);
nand I_12092 (I209166,I209149,I306466);
nor I_12093 (I209183,I209166,I209115);
DFFARX1 I_12094 (I209183,I3563,I208965,I208933,);
not I_12095 (I209214,I209166);
not I_12096 (I209231,I306469);
nand I_12097 (I209248,I209231,I306457);
nor I_12098 (I209265,I306469,I306445);
nand I_12099 (I208945,I209081,I209265);
nand I_12100 (I208939,I209030,I306469);
nand I_12101 (I209310,I209132,I306463);
DFFARX1 I_12102 (I209310,I3563,I208965,I208954,);
DFFARX1 I_12103 (I209310,I3563,I208965,I208948,);
not I_12104 (I209355,I306463);
nor I_12105 (I209372,I209355,I306451);
and I_12106 (I209389,I209372,I306472);
or I_12107 (I209406,I209389,I306448);
DFFARX1 I_12108 (I209406,I3563,I208965,I209432,);
nand I_12109 (I209440,I209432,I209098);
nor I_12110 (I208942,I209440,I209248);
nor I_12111 (I208936,I209432,I209064);
DFFARX1 I_12112 (I209432,I3563,I208965,I209494,);
not I_12113 (I209502,I209494);
nor I_12114 (I208951,I209502,I209214);
not I_12115 (I209560,I3570);
DFFARX1 I_12116 (I107775,I3563,I209560,I209586,);
DFFARX1 I_12117 (I209586,I3563,I209560,I209603,);
not I_12118 (I209552,I209603);
not I_12119 (I209625,I209586);
DFFARX1 I_12120 (I107769,I3563,I209560,I209651,);
not I_12121 (I209659,I209651);
and I_12122 (I209676,I209625,I107766);
not I_12123 (I209693,I107787);
nand I_12124 (I209710,I209693,I107766);
not I_12125 (I209727,I107781);
nor I_12126 (I209744,I209727,I107772);
nand I_12127 (I209761,I209744,I107778);
nor I_12128 (I209778,I209761,I209710);
DFFARX1 I_12129 (I209778,I3563,I209560,I209528,);
not I_12130 (I209809,I209761);
not I_12131 (I209826,I107772);
nand I_12132 (I209843,I209826,I107766);
nor I_12133 (I209860,I107772,I107787);
nand I_12134 (I209540,I209676,I209860);
nand I_12135 (I209534,I209625,I107772);
nand I_12136 (I209905,I209727,I107766);
DFFARX1 I_12137 (I209905,I3563,I209560,I209549,);
DFFARX1 I_12138 (I209905,I3563,I209560,I209543,);
not I_12139 (I209950,I107766);
nor I_12140 (I209967,I209950,I107784);
and I_12141 (I209984,I209967,I107790);
or I_12142 (I210001,I209984,I107769);
DFFARX1 I_12143 (I210001,I3563,I209560,I210027,);
nand I_12144 (I210035,I210027,I209693);
nor I_12145 (I209537,I210035,I209843);
nor I_12146 (I209531,I210027,I209659);
DFFARX1 I_12147 (I210027,I3563,I209560,I210089,);
not I_12148 (I210097,I210089);
nor I_12149 (I209546,I210097,I209809);
not I_12150 (I210155,I3570);
DFFARX1 I_12151 (I108302,I3563,I210155,I210181,);
DFFARX1 I_12152 (I210181,I3563,I210155,I210198,);
not I_12153 (I210147,I210198);
not I_12154 (I210220,I210181);
DFFARX1 I_12155 (I108296,I3563,I210155,I210246,);
not I_12156 (I210254,I210246);
and I_12157 (I210271,I210220,I108293);
not I_12158 (I210288,I108314);
nand I_12159 (I210305,I210288,I108293);
not I_12160 (I210322,I108308);
nor I_12161 (I210339,I210322,I108299);
nand I_12162 (I210356,I210339,I108305);
nor I_12163 (I210373,I210356,I210305);
DFFARX1 I_12164 (I210373,I3563,I210155,I210123,);
not I_12165 (I210404,I210356);
not I_12166 (I210421,I108299);
nand I_12167 (I210438,I210421,I108293);
nor I_12168 (I210455,I108299,I108314);
nand I_12169 (I210135,I210271,I210455);
nand I_12170 (I210129,I210220,I108299);
nand I_12171 (I210500,I210322,I108293);
DFFARX1 I_12172 (I210500,I3563,I210155,I210144,);
DFFARX1 I_12173 (I210500,I3563,I210155,I210138,);
not I_12174 (I210545,I108293);
nor I_12175 (I210562,I210545,I108311);
and I_12176 (I210579,I210562,I108317);
or I_12177 (I210596,I210579,I108296);
DFFARX1 I_12178 (I210596,I3563,I210155,I210622,);
nand I_12179 (I210630,I210622,I210288);
nor I_12180 (I210132,I210630,I210438);
nor I_12181 (I210126,I210622,I210254);
DFFARX1 I_12182 (I210622,I3563,I210155,I210684,);
not I_12183 (I210692,I210684);
nor I_12184 (I210141,I210692,I210404);
not I_12185 (I210750,I3570);
DFFARX1 I_12186 (I1271451,I3563,I210750,I210776,);
DFFARX1 I_12187 (I210776,I3563,I210750,I210793,);
not I_12188 (I210742,I210793);
not I_12189 (I210815,I210776);
DFFARX1 I_12190 (I1271436,I3563,I210750,I210841,);
not I_12191 (I210849,I210841);
and I_12192 (I210866,I210815,I1271454);
not I_12193 (I210883,I1271436);
nand I_12194 (I210900,I210883,I1271454);
not I_12195 (I210917,I1271457);
nor I_12196 (I210934,I210917,I1271448);
nand I_12197 (I210951,I210934,I1271445);
nor I_12198 (I210968,I210951,I210900);
DFFARX1 I_12199 (I210968,I3563,I210750,I210718,);
not I_12200 (I210999,I210951);
not I_12201 (I211016,I1271448);
nand I_12202 (I211033,I211016,I1271454);
nor I_12203 (I211050,I1271448,I1271436);
nand I_12204 (I210730,I210866,I211050);
nand I_12205 (I210724,I210815,I1271448);
nand I_12206 (I211095,I210917,I1271442);
DFFARX1 I_12207 (I211095,I3563,I210750,I210739,);
DFFARX1 I_12208 (I211095,I3563,I210750,I210733,);
not I_12209 (I211140,I1271442);
nor I_12210 (I211157,I211140,I1271433);
and I_12211 (I211174,I211157,I1271439);
or I_12212 (I211191,I211174,I1271433);
DFFARX1 I_12213 (I211191,I3563,I210750,I211217,);
nand I_12214 (I211225,I211217,I210883);
nor I_12215 (I210727,I211225,I211033);
nor I_12216 (I210721,I211217,I210849);
DFFARX1 I_12217 (I211217,I3563,I210750,I211279,);
not I_12218 (I211287,I211279);
nor I_12219 (I210736,I211287,I210999);
not I_12220 (I211345,I3570);
DFFARX1 I_12221 (I1332144,I3563,I211345,I211371,);
DFFARX1 I_12222 (I211371,I3563,I211345,I211388,);
not I_12223 (I211337,I211388);
not I_12224 (I211410,I211371);
DFFARX1 I_12225 (I1332135,I3563,I211345,I211436,);
not I_12226 (I211444,I211436);
and I_12227 (I211461,I211410,I1332129);
not I_12228 (I211478,I1332123);
nand I_12229 (I211495,I211478,I1332129);
not I_12230 (I211512,I1332150);
nor I_12231 (I211529,I211512,I1332123);
nand I_12232 (I211546,I211529,I1332147);
nor I_12233 (I211563,I211546,I211495);
DFFARX1 I_12234 (I211563,I3563,I211345,I211313,);
not I_12235 (I211594,I211546);
not I_12236 (I211611,I1332123);
nand I_12237 (I211628,I211611,I1332129);
nor I_12238 (I211645,I1332123,I1332123);
nand I_12239 (I211325,I211461,I211645);
nand I_12240 (I211319,I211410,I1332123);
nand I_12241 (I211690,I211512,I1332132);
DFFARX1 I_12242 (I211690,I3563,I211345,I211334,);
DFFARX1 I_12243 (I211690,I3563,I211345,I211328,);
not I_12244 (I211735,I1332132);
nor I_12245 (I211752,I211735,I1332138);
and I_12246 (I211769,I211752,I1332141);
or I_12247 (I211786,I211769,I1332126);
DFFARX1 I_12248 (I211786,I3563,I211345,I211812,);
nand I_12249 (I211820,I211812,I211478);
nor I_12250 (I211322,I211820,I211628);
nor I_12251 (I211316,I211812,I211444);
DFFARX1 I_12252 (I211812,I3563,I211345,I211874,);
not I_12253 (I211882,I211874);
nor I_12254 (I211331,I211882,I211594);
not I_12255 (I211940,I3570);
DFFARX1 I_12256 (I313823,I3563,I211940,I211966,);
DFFARX1 I_12257 (I211966,I3563,I211940,I211983,);
not I_12258 (I211932,I211983);
not I_12259 (I212005,I211966);
DFFARX1 I_12260 (I313838,I3563,I211940,I212031,);
not I_12261 (I212039,I212031);
and I_12262 (I212056,I212005,I313835);
not I_12263 (I212073,I313823);
nand I_12264 (I212090,I212073,I313835);
not I_12265 (I212107,I313832);
nor I_12266 (I212124,I212107,I313847);
nand I_12267 (I212141,I212124,I313844);
nor I_12268 (I212158,I212141,I212090);
DFFARX1 I_12269 (I212158,I3563,I211940,I211908,);
not I_12270 (I212189,I212141);
not I_12271 (I212206,I313847);
nand I_12272 (I212223,I212206,I313835);
nor I_12273 (I212240,I313847,I313823);
nand I_12274 (I211920,I212056,I212240);
nand I_12275 (I211914,I212005,I313847);
nand I_12276 (I212285,I212107,I313841);
DFFARX1 I_12277 (I212285,I3563,I211940,I211929,);
DFFARX1 I_12278 (I212285,I3563,I211940,I211923,);
not I_12279 (I212330,I313841);
nor I_12280 (I212347,I212330,I313829);
and I_12281 (I212364,I212347,I313850);
or I_12282 (I212381,I212364,I313826);
DFFARX1 I_12283 (I212381,I3563,I211940,I212407,);
nand I_12284 (I212415,I212407,I212073);
nor I_12285 (I211917,I212415,I212223);
nor I_12286 (I211911,I212407,I212039);
DFFARX1 I_12287 (I212407,I3563,I211940,I212469,);
not I_12288 (I212477,I212469);
nor I_12289 (I211926,I212477,I212189);
not I_12290 (I212535,I3570);
DFFARX1 I_12291 (I354929,I3563,I212535,I212561,);
DFFARX1 I_12292 (I212561,I3563,I212535,I212578,);
not I_12293 (I212527,I212578);
not I_12294 (I212600,I212561);
DFFARX1 I_12295 (I354944,I3563,I212535,I212626,);
not I_12296 (I212634,I212626);
and I_12297 (I212651,I212600,I354941);
not I_12298 (I212668,I354929);
nand I_12299 (I212685,I212668,I354941);
not I_12300 (I212702,I354938);
nor I_12301 (I212719,I212702,I354953);
nand I_12302 (I212736,I212719,I354950);
nor I_12303 (I212753,I212736,I212685);
DFFARX1 I_12304 (I212753,I3563,I212535,I212503,);
not I_12305 (I212784,I212736);
not I_12306 (I212801,I354953);
nand I_12307 (I212818,I212801,I354941);
nor I_12308 (I212835,I354953,I354929);
nand I_12309 (I212515,I212651,I212835);
nand I_12310 (I212509,I212600,I354953);
nand I_12311 (I212880,I212702,I354947);
DFFARX1 I_12312 (I212880,I3563,I212535,I212524,);
DFFARX1 I_12313 (I212880,I3563,I212535,I212518,);
not I_12314 (I212925,I354947);
nor I_12315 (I212942,I212925,I354935);
and I_12316 (I212959,I212942,I354956);
or I_12317 (I212976,I212959,I354932);
DFFARX1 I_12318 (I212976,I3563,I212535,I213002,);
nand I_12319 (I213010,I213002,I212668);
nor I_12320 (I212512,I213010,I212818);
nor I_12321 (I212506,I213002,I212634);
DFFARX1 I_12322 (I213002,I3563,I212535,I213064,);
not I_12323 (I213072,I213064);
nor I_12324 (I212521,I213072,I212784);
not I_12325 (I213130,I3570);
DFFARX1 I_12326 (I331741,I3563,I213130,I213156,);
DFFARX1 I_12327 (I213156,I3563,I213130,I213173,);
not I_12328 (I213122,I213173);
not I_12329 (I213195,I213156);
DFFARX1 I_12330 (I331756,I3563,I213130,I213221,);
not I_12331 (I213229,I213221);
and I_12332 (I213246,I213195,I331753);
not I_12333 (I213263,I331741);
nand I_12334 (I213280,I213263,I331753);
not I_12335 (I213297,I331750);
nor I_12336 (I213314,I213297,I331765);
nand I_12337 (I213331,I213314,I331762);
nor I_12338 (I213348,I213331,I213280);
DFFARX1 I_12339 (I213348,I3563,I213130,I213098,);
not I_12340 (I213379,I213331);
not I_12341 (I213396,I331765);
nand I_12342 (I213413,I213396,I331753);
nor I_12343 (I213430,I331765,I331741);
nand I_12344 (I213110,I213246,I213430);
nand I_12345 (I213104,I213195,I331765);
nand I_12346 (I213475,I213297,I331759);
DFFARX1 I_12347 (I213475,I3563,I213130,I213119,);
DFFARX1 I_12348 (I213475,I3563,I213130,I213113,);
not I_12349 (I213520,I331759);
nor I_12350 (I213537,I213520,I331747);
and I_12351 (I213554,I213537,I331768);
or I_12352 (I213571,I213554,I331744);
DFFARX1 I_12353 (I213571,I3563,I213130,I213597,);
nand I_12354 (I213605,I213597,I213263);
nor I_12355 (I213107,I213605,I213413);
nor I_12356 (I213101,I213597,I213229);
DFFARX1 I_12357 (I213597,I3563,I213130,I213659,);
not I_12358 (I213667,I213659);
nor I_12359 (I213116,I213667,I213379);
not I_12360 (I213725,I3570);
DFFARX1 I_12361 (I449082,I3563,I213725,I213751,);
DFFARX1 I_12362 (I213751,I3563,I213725,I213768,);
not I_12363 (I213717,I213768);
not I_12364 (I213790,I213751);
DFFARX1 I_12365 (I449070,I3563,I213725,I213816,);
not I_12366 (I213824,I213816);
and I_12367 (I213841,I213790,I449079);
not I_12368 (I213858,I449076);
nand I_12369 (I213875,I213858,I449079);
not I_12370 (I213892,I449067);
nor I_12371 (I213909,I213892,I449073);
nand I_12372 (I213926,I213909,I449058);
nor I_12373 (I213943,I213926,I213875);
DFFARX1 I_12374 (I213943,I3563,I213725,I213693,);
not I_12375 (I213974,I213926);
not I_12376 (I213991,I449073);
nand I_12377 (I214008,I213991,I449079);
nor I_12378 (I214025,I449073,I449076);
nand I_12379 (I213705,I213841,I214025);
nand I_12380 (I213699,I213790,I449073);
nand I_12381 (I214070,I213892,I449058);
DFFARX1 I_12382 (I214070,I3563,I213725,I213714,);
DFFARX1 I_12383 (I214070,I3563,I213725,I213708,);
not I_12384 (I214115,I449058);
nor I_12385 (I214132,I214115,I449064);
and I_12386 (I214149,I214132,I449061);
or I_12387 (I214166,I214149,I449085);
DFFARX1 I_12388 (I214166,I3563,I213725,I214192,);
nand I_12389 (I214200,I214192,I213858);
nor I_12390 (I213702,I214200,I214008);
nor I_12391 (I213696,I214192,I213824);
DFFARX1 I_12392 (I214192,I3563,I213725,I214254,);
not I_12393 (I214262,I214254);
nor I_12394 (I213711,I214262,I213974);
not I_12395 (I214320,I3570);
DFFARX1 I_12396 (I1051711,I3563,I214320,I214346,);
DFFARX1 I_12397 (I214346,I3563,I214320,I214363,);
not I_12398 (I214312,I214363);
not I_12399 (I214385,I214346);
DFFARX1 I_12400 (I1051720,I3563,I214320,I214411,);
not I_12401 (I214419,I214411);
and I_12402 (I214436,I214385,I1051714);
not I_12403 (I214453,I1051708);
nand I_12404 (I214470,I214453,I1051714);
not I_12405 (I214487,I1051723);
nor I_12406 (I214504,I214487,I1051711);
nand I_12407 (I214521,I214504,I1051717);
nor I_12408 (I214538,I214521,I214470);
DFFARX1 I_12409 (I214538,I3563,I214320,I214288,);
not I_12410 (I214569,I214521);
not I_12411 (I214586,I1051711);
nand I_12412 (I214603,I214586,I1051714);
nor I_12413 (I214620,I1051711,I1051708);
nand I_12414 (I214300,I214436,I214620);
nand I_12415 (I214294,I214385,I1051711);
nand I_12416 (I214665,I214487,I1051714);
DFFARX1 I_12417 (I214665,I3563,I214320,I214309,);
DFFARX1 I_12418 (I214665,I3563,I214320,I214303,);
not I_12419 (I214710,I1051714);
nor I_12420 (I214727,I214710,I1051729);
and I_12421 (I214744,I214727,I1051726);
or I_12422 (I214761,I214744,I1051708);
DFFARX1 I_12423 (I214761,I3563,I214320,I214787,);
nand I_12424 (I214795,I214787,I214453);
nor I_12425 (I214297,I214795,I214603);
nor I_12426 (I214291,I214787,I214419);
DFFARX1 I_12427 (I214787,I3563,I214320,I214849,);
not I_12428 (I214857,I214849);
nor I_12429 (I214306,I214857,I214569);
not I_12430 (I214915,I3570);
DFFARX1 I_12431 (I860073,I3563,I214915,I214941,);
DFFARX1 I_12432 (I214941,I3563,I214915,I214958,);
not I_12433 (I214907,I214958);
not I_12434 (I214980,I214941);
DFFARX1 I_12435 (I860067,I3563,I214915,I215006,);
not I_12436 (I215014,I215006);
and I_12437 (I215031,I214980,I860085);
not I_12438 (I215048,I860073);
nand I_12439 (I215065,I215048,I860085);
not I_12440 (I215082,I860067);
nor I_12441 (I215099,I215082,I860079);
nand I_12442 (I215116,I215099,I860070);
nor I_12443 (I215133,I215116,I215065);
DFFARX1 I_12444 (I215133,I3563,I214915,I214883,);
not I_12445 (I215164,I215116);
not I_12446 (I215181,I860079);
nand I_12447 (I215198,I215181,I860085);
nor I_12448 (I215215,I860079,I860073);
nand I_12449 (I214895,I215031,I215215);
nand I_12450 (I214889,I214980,I860079);
nand I_12451 (I215260,I215082,I860082);
DFFARX1 I_12452 (I215260,I3563,I214915,I214904,);
DFFARX1 I_12453 (I215260,I3563,I214915,I214898,);
not I_12454 (I215305,I860082);
nor I_12455 (I215322,I215305,I860088);
and I_12456 (I215339,I215322,I860070);
or I_12457 (I215356,I215339,I860076);
DFFARX1 I_12458 (I215356,I3563,I214915,I215382,);
nand I_12459 (I215390,I215382,I215048);
nor I_12460 (I214892,I215390,I215198);
nor I_12461 (I214886,I215382,I215014);
DFFARX1 I_12462 (I215382,I3563,I214915,I215444,);
not I_12463 (I215452,I215444);
nor I_12464 (I214901,I215452,I215164);
not I_12465 (I215510,I3570);
DFFARX1 I_12466 (I357037,I3563,I215510,I215536,);
DFFARX1 I_12467 (I215536,I3563,I215510,I215553,);
not I_12468 (I215502,I215553);
not I_12469 (I215575,I215536);
DFFARX1 I_12470 (I357052,I3563,I215510,I215601,);
not I_12471 (I215609,I215601);
and I_12472 (I215626,I215575,I357049);
not I_12473 (I215643,I357037);
nand I_12474 (I215660,I215643,I357049);
not I_12475 (I215677,I357046);
nor I_12476 (I215694,I215677,I357061);
nand I_12477 (I215711,I215694,I357058);
nor I_12478 (I215728,I215711,I215660);
DFFARX1 I_12479 (I215728,I3563,I215510,I215478,);
not I_12480 (I215759,I215711);
not I_12481 (I215776,I357061);
nand I_12482 (I215793,I215776,I357049);
nor I_12483 (I215810,I357061,I357037);
nand I_12484 (I215490,I215626,I215810);
nand I_12485 (I215484,I215575,I357061);
nand I_12486 (I215855,I215677,I357055);
DFFARX1 I_12487 (I215855,I3563,I215510,I215499,);
DFFARX1 I_12488 (I215855,I3563,I215510,I215493,);
not I_12489 (I215900,I357055);
nor I_12490 (I215917,I215900,I357043);
and I_12491 (I215934,I215917,I357064);
or I_12492 (I215951,I215934,I357040);
DFFARX1 I_12493 (I215951,I3563,I215510,I215977,);
nand I_12494 (I215985,I215977,I215643);
nor I_12495 (I215487,I215985,I215793);
nor I_12496 (I215481,I215977,I215609);
DFFARX1 I_12497 (I215977,I3563,I215510,I216039,);
not I_12498 (I216047,I216039);
nor I_12499 (I215496,I216047,I215759);
not I_12500 (I216105,I3570);
DFFARX1 I_12501 (I120950,I3563,I216105,I216131,);
DFFARX1 I_12502 (I216131,I3563,I216105,I216148,);
not I_12503 (I216097,I216148);
not I_12504 (I216170,I216131);
DFFARX1 I_12505 (I120944,I3563,I216105,I216196,);
not I_12506 (I216204,I216196);
and I_12507 (I216221,I216170,I120941);
not I_12508 (I216238,I120962);
nand I_12509 (I216255,I216238,I120941);
not I_12510 (I216272,I120956);
nor I_12511 (I216289,I216272,I120947);
nand I_12512 (I216306,I216289,I120953);
nor I_12513 (I216323,I216306,I216255);
DFFARX1 I_12514 (I216323,I3563,I216105,I216073,);
not I_12515 (I216354,I216306);
not I_12516 (I216371,I120947);
nand I_12517 (I216388,I216371,I120941);
nor I_12518 (I216405,I120947,I120962);
nand I_12519 (I216085,I216221,I216405);
nand I_12520 (I216079,I216170,I120947);
nand I_12521 (I216450,I216272,I120941);
DFFARX1 I_12522 (I216450,I3563,I216105,I216094,);
DFFARX1 I_12523 (I216450,I3563,I216105,I216088,);
not I_12524 (I216495,I120941);
nor I_12525 (I216512,I216495,I120959);
and I_12526 (I216529,I216512,I120965);
or I_12527 (I216546,I216529,I120944);
DFFARX1 I_12528 (I216546,I3563,I216105,I216572,);
nand I_12529 (I216580,I216572,I216238);
nor I_12530 (I216082,I216580,I216388);
nor I_12531 (I216076,I216572,I216204);
DFFARX1 I_12532 (I216572,I3563,I216105,I216634,);
not I_12533 (I216642,I216634);
nor I_12534 (I216091,I216642,I216354);
not I_12535 (I216700,I3570);
DFFARX1 I_12536 (I1262747,I3563,I216700,I216726,);
DFFARX1 I_12537 (I216726,I3563,I216700,I216743,);
not I_12538 (I216692,I216743);
not I_12539 (I216765,I216726);
DFFARX1 I_12540 (I1262732,I3563,I216700,I216791,);
not I_12541 (I216799,I216791);
and I_12542 (I216816,I216765,I1262750);
not I_12543 (I216833,I1262732);
nand I_12544 (I216850,I216833,I1262750);
not I_12545 (I216867,I1262753);
nor I_12546 (I216884,I216867,I1262744);
nand I_12547 (I216901,I216884,I1262741);
nor I_12548 (I216918,I216901,I216850);
DFFARX1 I_12549 (I216918,I3563,I216700,I216668,);
not I_12550 (I216949,I216901);
not I_12551 (I216966,I1262744);
nand I_12552 (I216983,I216966,I1262750);
nor I_12553 (I217000,I1262744,I1262732);
nand I_12554 (I216680,I216816,I217000);
nand I_12555 (I216674,I216765,I1262744);
nand I_12556 (I217045,I216867,I1262738);
DFFARX1 I_12557 (I217045,I3563,I216700,I216689,);
DFFARX1 I_12558 (I217045,I3563,I216700,I216683,);
not I_12559 (I217090,I1262738);
nor I_12560 (I217107,I217090,I1262729);
and I_12561 (I217124,I217107,I1262735);
or I_12562 (I217141,I217124,I1262729);
DFFARX1 I_12563 (I217141,I3563,I216700,I217167,);
nand I_12564 (I217175,I217167,I216833);
nor I_12565 (I216677,I217175,I216983);
nor I_12566 (I216671,I217167,I216799);
DFFARX1 I_12567 (I217167,I3563,I216700,I217229,);
not I_12568 (I217237,I217229);
nor I_12569 (I216686,I217237,I216949);
not I_12570 (I217295,I3570);
DFFARX1 I_12571 (I1120473,I3563,I217295,I217321,);
DFFARX1 I_12572 (I217321,I3563,I217295,I217338,);
not I_12573 (I217287,I217338);
not I_12574 (I217360,I217321);
DFFARX1 I_12575 (I1120473,I3563,I217295,I217386,);
not I_12576 (I217394,I217386);
and I_12577 (I217411,I217360,I1120476);
not I_12578 (I217428,I1120488);
nand I_12579 (I217445,I217428,I1120476);
not I_12580 (I217462,I1120494);
nor I_12581 (I217479,I217462,I1120485);
nand I_12582 (I217496,I217479,I1120491);
nor I_12583 (I217513,I217496,I217445);
DFFARX1 I_12584 (I217513,I3563,I217295,I217263,);
not I_12585 (I217544,I217496);
not I_12586 (I217561,I1120485);
nand I_12587 (I217578,I217561,I1120476);
nor I_12588 (I217595,I1120485,I1120488);
nand I_12589 (I217275,I217411,I217595);
nand I_12590 (I217269,I217360,I1120485);
nand I_12591 (I217640,I217462,I1120482);
DFFARX1 I_12592 (I217640,I3563,I217295,I217284,);
DFFARX1 I_12593 (I217640,I3563,I217295,I217278,);
not I_12594 (I217685,I1120482);
nor I_12595 (I217702,I217685,I1120479);
and I_12596 (I217719,I217702,I1120497);
or I_12597 (I217736,I217719,I1120476);
DFFARX1 I_12598 (I217736,I3563,I217295,I217762,);
nand I_12599 (I217770,I217762,I217428);
nor I_12600 (I217272,I217770,I217578);
nor I_12601 (I217266,I217762,I217394);
DFFARX1 I_12602 (I217762,I3563,I217295,I217824,);
not I_12603 (I217832,I217824);
nor I_12604 (I217281,I217832,I217544);
not I_12605 (I217890,I3570);
DFFARX1 I_12606 (I734143,I3563,I217890,I217916,);
DFFARX1 I_12607 (I217916,I3563,I217890,I217933,);
not I_12608 (I217882,I217933);
not I_12609 (I217955,I217916);
DFFARX1 I_12610 (I734140,I3563,I217890,I217981,);
not I_12611 (I217989,I217981);
and I_12612 (I218006,I217955,I734146);
not I_12613 (I218023,I734131);
nand I_12614 (I218040,I218023,I734146);
not I_12615 (I218057,I734134);
nor I_12616 (I218074,I218057,I734155);
nand I_12617 (I218091,I218074,I734152);
nor I_12618 (I218108,I218091,I218040);
DFFARX1 I_12619 (I218108,I3563,I217890,I217858,);
not I_12620 (I218139,I218091);
not I_12621 (I218156,I734155);
nand I_12622 (I218173,I218156,I734146);
nor I_12623 (I218190,I734155,I734131);
nand I_12624 (I217870,I218006,I218190);
nand I_12625 (I217864,I217955,I734155);
nand I_12626 (I218235,I218057,I734131);
DFFARX1 I_12627 (I218235,I3563,I217890,I217879,);
DFFARX1 I_12628 (I218235,I3563,I217890,I217873,);
not I_12629 (I218280,I734131);
nor I_12630 (I218297,I218280,I734137);
and I_12631 (I218314,I218297,I734149);
or I_12632 (I218331,I218314,I734134);
DFFARX1 I_12633 (I218331,I3563,I217890,I218357,);
nand I_12634 (I218365,I218357,I218023);
nor I_12635 (I217867,I218365,I218173);
nor I_12636 (I217861,I218357,I217989);
DFFARX1 I_12637 (I218357,I3563,I217890,I218419,);
not I_12638 (I218427,I218419);
nor I_12639 (I217876,I218427,I218139);
not I_12640 (I218485,I3570);
DFFARX1 I_12641 (I844790,I3563,I218485,I218511,);
DFFARX1 I_12642 (I218511,I3563,I218485,I218528,);
not I_12643 (I218477,I218528);
not I_12644 (I218550,I218511);
DFFARX1 I_12645 (I844784,I3563,I218485,I218576,);
not I_12646 (I218584,I218576);
and I_12647 (I218601,I218550,I844802);
not I_12648 (I218618,I844790);
nand I_12649 (I218635,I218618,I844802);
not I_12650 (I218652,I844784);
nor I_12651 (I218669,I218652,I844796);
nand I_12652 (I218686,I218669,I844787);
nor I_12653 (I218703,I218686,I218635);
DFFARX1 I_12654 (I218703,I3563,I218485,I218453,);
not I_12655 (I218734,I218686);
not I_12656 (I218751,I844796);
nand I_12657 (I218768,I218751,I844802);
nor I_12658 (I218785,I844796,I844790);
nand I_12659 (I218465,I218601,I218785);
nand I_12660 (I218459,I218550,I844796);
nand I_12661 (I218830,I218652,I844799);
DFFARX1 I_12662 (I218830,I3563,I218485,I218474,);
DFFARX1 I_12663 (I218830,I3563,I218485,I218468,);
not I_12664 (I218875,I844799);
nor I_12665 (I218892,I218875,I844805);
and I_12666 (I218909,I218892,I844787);
or I_12667 (I218926,I218909,I844793);
DFFARX1 I_12668 (I218926,I3563,I218485,I218952,);
nand I_12669 (I218960,I218952,I218618);
nor I_12670 (I218462,I218960,I218768);
nor I_12671 (I218456,I218952,I218584);
DFFARX1 I_12672 (I218952,I3563,I218485,I219014,);
not I_12673 (I219022,I219014);
nor I_12674 (I218471,I219022,I218734);
not I_12675 (I219080,I3570);
DFFARX1 I_12676 (I686169,I3563,I219080,I219106,);
DFFARX1 I_12677 (I219106,I3563,I219080,I219123,);
not I_12678 (I219072,I219123);
not I_12679 (I219145,I219106);
DFFARX1 I_12680 (I686166,I3563,I219080,I219171,);
not I_12681 (I219179,I219171);
and I_12682 (I219196,I219145,I686172);
not I_12683 (I219213,I686157);
nand I_12684 (I219230,I219213,I686172);
not I_12685 (I219247,I686160);
nor I_12686 (I219264,I219247,I686181);
nand I_12687 (I219281,I219264,I686178);
nor I_12688 (I219298,I219281,I219230);
DFFARX1 I_12689 (I219298,I3563,I219080,I219048,);
not I_12690 (I219329,I219281);
not I_12691 (I219346,I686181);
nand I_12692 (I219363,I219346,I686172);
nor I_12693 (I219380,I686181,I686157);
nand I_12694 (I219060,I219196,I219380);
nand I_12695 (I219054,I219145,I686181);
nand I_12696 (I219425,I219247,I686157);
DFFARX1 I_12697 (I219425,I3563,I219080,I219069,);
DFFARX1 I_12698 (I219425,I3563,I219080,I219063,);
not I_12699 (I219470,I686157);
nor I_12700 (I219487,I219470,I686163);
and I_12701 (I219504,I219487,I686175);
or I_12702 (I219521,I219504,I686160);
DFFARX1 I_12703 (I219521,I3563,I219080,I219547,);
nand I_12704 (I219555,I219547,I219213);
nor I_12705 (I219057,I219555,I219363);
nor I_12706 (I219051,I219547,I219179);
DFFARX1 I_12707 (I219547,I3563,I219080,I219609,);
not I_12708 (I219617,I219609);
nor I_12709 (I219066,I219617,I219329);
not I_12710 (I219675,I3570);
DFFARX1 I_12711 (I152043,I3563,I219675,I219701,);
DFFARX1 I_12712 (I219701,I3563,I219675,I219718,);
not I_12713 (I219667,I219718);
not I_12714 (I219740,I219701);
DFFARX1 I_12715 (I152037,I3563,I219675,I219766,);
not I_12716 (I219774,I219766);
and I_12717 (I219791,I219740,I152034);
not I_12718 (I219808,I152055);
nand I_12719 (I219825,I219808,I152034);
not I_12720 (I219842,I152049);
nor I_12721 (I219859,I219842,I152040);
nand I_12722 (I219876,I219859,I152046);
nor I_12723 (I219893,I219876,I219825);
DFFARX1 I_12724 (I219893,I3563,I219675,I219643,);
not I_12725 (I219924,I219876);
not I_12726 (I219941,I152040);
nand I_12727 (I219958,I219941,I152034);
nor I_12728 (I219975,I152040,I152055);
nand I_12729 (I219655,I219791,I219975);
nand I_12730 (I219649,I219740,I152040);
nand I_12731 (I220020,I219842,I152034);
DFFARX1 I_12732 (I220020,I3563,I219675,I219664,);
DFFARX1 I_12733 (I220020,I3563,I219675,I219658,);
not I_12734 (I220065,I152034);
nor I_12735 (I220082,I220065,I152052);
and I_12736 (I220099,I220082,I152058);
or I_12737 (I220116,I220099,I152037);
DFFARX1 I_12738 (I220116,I3563,I219675,I220142,);
nand I_12739 (I220150,I220142,I219808);
nor I_12740 (I219652,I220150,I219958);
nor I_12741 (I219646,I220142,I219774);
DFFARX1 I_12742 (I220142,I3563,I219675,I220204,);
not I_12743 (I220212,I220204);
nor I_12744 (I219661,I220212,I219924);
not I_12745 (I220270,I3570);
DFFARX1 I_12746 (I1072468,I3563,I220270,I220296,);
DFFARX1 I_12747 (I220296,I3563,I220270,I220313,);
not I_12748 (I220262,I220313);
not I_12749 (I220335,I220296);
DFFARX1 I_12750 (I1072477,I3563,I220270,I220361,);
not I_12751 (I220369,I220361);
and I_12752 (I220386,I220335,I1072471);
not I_12753 (I220403,I1072465);
nand I_12754 (I220420,I220403,I1072471);
not I_12755 (I220437,I1072480);
nor I_12756 (I220454,I220437,I1072468);
nand I_12757 (I220471,I220454,I1072474);
nor I_12758 (I220488,I220471,I220420);
DFFARX1 I_12759 (I220488,I3563,I220270,I220238,);
not I_12760 (I220519,I220471);
not I_12761 (I220536,I1072468);
nand I_12762 (I220553,I220536,I1072471);
nor I_12763 (I220570,I1072468,I1072465);
nand I_12764 (I220250,I220386,I220570);
nand I_12765 (I220244,I220335,I1072468);
nand I_12766 (I220615,I220437,I1072471);
DFFARX1 I_12767 (I220615,I3563,I220270,I220259,);
DFFARX1 I_12768 (I220615,I3563,I220270,I220253,);
not I_12769 (I220660,I1072471);
nor I_12770 (I220677,I220660,I1072486);
and I_12771 (I220694,I220677,I1072483);
or I_12772 (I220711,I220694,I1072465);
DFFARX1 I_12773 (I220711,I3563,I220270,I220737,);
nand I_12774 (I220745,I220737,I220403);
nor I_12775 (I220247,I220745,I220553);
nor I_12776 (I220241,I220737,I220369);
DFFARX1 I_12777 (I220737,I3563,I220270,I220799,);
not I_12778 (I220807,I220799);
nor I_12779 (I220256,I220807,I220519);
not I_12780 (I220865,I3570);
DFFARX1 I_12781 (I947190,I3563,I220865,I220891,);
DFFARX1 I_12782 (I220891,I3563,I220865,I220908,);
not I_12783 (I220857,I220908);
not I_12784 (I220930,I220891);
DFFARX1 I_12785 (I947199,I3563,I220865,I220956,);
not I_12786 (I220964,I220956);
and I_12787 (I220981,I220930,I947187);
not I_12788 (I220998,I947178);
nand I_12789 (I221015,I220998,I947187);
not I_12790 (I221032,I947184);
nor I_12791 (I221049,I221032,I947202);
nand I_12792 (I221066,I221049,I947175);
nor I_12793 (I221083,I221066,I221015);
DFFARX1 I_12794 (I221083,I3563,I220865,I220833,);
not I_12795 (I221114,I221066);
not I_12796 (I221131,I947202);
nand I_12797 (I221148,I221131,I947187);
nor I_12798 (I221165,I947202,I947178);
nand I_12799 (I220845,I220981,I221165);
nand I_12800 (I220839,I220930,I947202);
nand I_12801 (I221210,I221032,I947181);
DFFARX1 I_12802 (I221210,I3563,I220865,I220854,);
DFFARX1 I_12803 (I221210,I3563,I220865,I220848,);
not I_12804 (I221255,I947181);
nor I_12805 (I221272,I221255,I947193);
and I_12806 (I221289,I221272,I947175);
or I_12807 (I221306,I221289,I947196);
DFFARX1 I_12808 (I221306,I3563,I220865,I221332,);
nand I_12809 (I221340,I221332,I220998);
nor I_12810 (I220842,I221340,I221148);
nor I_12811 (I220836,I221332,I220964);
DFFARX1 I_12812 (I221332,I3563,I220865,I221394,);
not I_12813 (I221402,I221394);
nor I_12814 (I220851,I221402,I221114);
not I_12815 (I221460,I3570);
DFFARX1 I_12816 (I992410,I3563,I221460,I221486,);
DFFARX1 I_12817 (I221486,I3563,I221460,I221503,);
not I_12818 (I221452,I221503);
not I_12819 (I221525,I221486);
DFFARX1 I_12820 (I992419,I3563,I221460,I221551,);
not I_12821 (I221559,I221551);
and I_12822 (I221576,I221525,I992407);
not I_12823 (I221593,I992398);
nand I_12824 (I221610,I221593,I992407);
not I_12825 (I221627,I992404);
nor I_12826 (I221644,I221627,I992422);
nand I_12827 (I221661,I221644,I992395);
nor I_12828 (I221678,I221661,I221610);
DFFARX1 I_12829 (I221678,I3563,I221460,I221428,);
not I_12830 (I221709,I221661);
not I_12831 (I221726,I992422);
nand I_12832 (I221743,I221726,I992407);
nor I_12833 (I221760,I992422,I992398);
nand I_12834 (I221440,I221576,I221760);
nand I_12835 (I221434,I221525,I992422);
nand I_12836 (I221805,I221627,I992401);
DFFARX1 I_12837 (I221805,I3563,I221460,I221449,);
DFFARX1 I_12838 (I221805,I3563,I221460,I221443,);
not I_12839 (I221850,I992401);
nor I_12840 (I221867,I221850,I992413);
and I_12841 (I221884,I221867,I992395);
or I_12842 (I221901,I221884,I992416);
DFFARX1 I_12843 (I221901,I3563,I221460,I221927,);
nand I_12844 (I221935,I221927,I221593);
nor I_12845 (I221437,I221935,I221743);
nor I_12846 (I221431,I221927,I221559);
DFFARX1 I_12847 (I221927,I3563,I221460,I221989,);
not I_12848 (I221997,I221989);
nor I_12849 (I221446,I221997,I221709);
not I_12850 (I222055,I3570);
DFFARX1 I_12851 (I1358919,I3563,I222055,I222081,);
DFFARX1 I_12852 (I222081,I3563,I222055,I222098,);
not I_12853 (I222047,I222098);
not I_12854 (I222120,I222081);
DFFARX1 I_12855 (I1358910,I3563,I222055,I222146,);
not I_12856 (I222154,I222146);
and I_12857 (I222171,I222120,I1358904);
not I_12858 (I222188,I1358898);
nand I_12859 (I222205,I222188,I1358904);
not I_12860 (I222222,I1358925);
nor I_12861 (I222239,I222222,I1358898);
nand I_12862 (I222256,I222239,I1358922);
nor I_12863 (I222273,I222256,I222205);
DFFARX1 I_12864 (I222273,I3563,I222055,I222023,);
not I_12865 (I222304,I222256);
not I_12866 (I222321,I1358898);
nand I_12867 (I222338,I222321,I1358904);
nor I_12868 (I222355,I1358898,I1358898);
nand I_12869 (I222035,I222171,I222355);
nand I_12870 (I222029,I222120,I1358898);
nand I_12871 (I222400,I222222,I1358907);
DFFARX1 I_12872 (I222400,I3563,I222055,I222044,);
DFFARX1 I_12873 (I222400,I3563,I222055,I222038,);
not I_12874 (I222445,I1358907);
nor I_12875 (I222462,I222445,I1358913);
and I_12876 (I222479,I222462,I1358916);
or I_12877 (I222496,I222479,I1358901);
DFFARX1 I_12878 (I222496,I3563,I222055,I222522,);
nand I_12879 (I222530,I222522,I222188);
nor I_12880 (I222032,I222530,I222338);
nor I_12881 (I222026,I222522,I222154);
DFFARX1 I_12882 (I222522,I3563,I222055,I222584,);
not I_12883 (I222592,I222584);
nor I_12884 (I222041,I222592,I222304);
not I_12885 (I222650,I3570);
DFFARX1 I_12886 (I60345,I3563,I222650,I222676,);
DFFARX1 I_12887 (I222676,I3563,I222650,I222693,);
not I_12888 (I222642,I222693);
not I_12889 (I222715,I222676);
DFFARX1 I_12890 (I60339,I3563,I222650,I222741,);
not I_12891 (I222749,I222741);
and I_12892 (I222766,I222715,I60336);
not I_12893 (I222783,I60357);
nand I_12894 (I222800,I222783,I60336);
not I_12895 (I222817,I60351);
nor I_12896 (I222834,I222817,I60342);
nand I_12897 (I222851,I222834,I60348);
nor I_12898 (I222868,I222851,I222800);
DFFARX1 I_12899 (I222868,I3563,I222650,I222618,);
not I_12900 (I222899,I222851);
not I_12901 (I222916,I60342);
nand I_12902 (I222933,I222916,I60336);
nor I_12903 (I222950,I60342,I60357);
nand I_12904 (I222630,I222766,I222950);
nand I_12905 (I222624,I222715,I60342);
nand I_12906 (I222995,I222817,I60336);
DFFARX1 I_12907 (I222995,I3563,I222650,I222639,);
DFFARX1 I_12908 (I222995,I3563,I222650,I222633,);
not I_12909 (I223040,I60336);
nor I_12910 (I223057,I223040,I60354);
and I_12911 (I223074,I223057,I60360);
or I_12912 (I223091,I223074,I60339);
DFFARX1 I_12913 (I223091,I3563,I222650,I223117,);
nand I_12914 (I223125,I223117,I222783);
nor I_12915 (I222627,I223125,I222933);
nor I_12916 (I222621,I223117,I222749);
DFFARX1 I_12917 (I223117,I3563,I222650,I223179,);
not I_12918 (I223187,I223179);
nor I_12919 (I222636,I223187,I222899);
not I_12920 (I223245,I3570);
DFFARX1 I_12921 (I1391049,I3563,I223245,I223271,);
DFFARX1 I_12922 (I223271,I3563,I223245,I223288,);
not I_12923 (I223237,I223288);
not I_12924 (I223310,I223271);
DFFARX1 I_12925 (I1391040,I3563,I223245,I223336,);
not I_12926 (I223344,I223336);
and I_12927 (I223361,I223310,I1391034);
not I_12928 (I223378,I1391028);
nand I_12929 (I223395,I223378,I1391034);
not I_12930 (I223412,I1391055);
nor I_12931 (I223429,I223412,I1391028);
nand I_12932 (I223446,I223429,I1391052);
nor I_12933 (I223463,I223446,I223395);
DFFARX1 I_12934 (I223463,I3563,I223245,I223213,);
not I_12935 (I223494,I223446);
not I_12936 (I223511,I1391028);
nand I_12937 (I223528,I223511,I1391034);
nor I_12938 (I223545,I1391028,I1391028);
nand I_12939 (I223225,I223361,I223545);
nand I_12940 (I223219,I223310,I1391028);
nand I_12941 (I223590,I223412,I1391037);
DFFARX1 I_12942 (I223590,I3563,I223245,I223234,);
DFFARX1 I_12943 (I223590,I3563,I223245,I223228,);
not I_12944 (I223635,I1391037);
nor I_12945 (I223652,I223635,I1391043);
and I_12946 (I223669,I223652,I1391046);
or I_12947 (I223686,I223669,I1391031);
DFFARX1 I_12948 (I223686,I3563,I223245,I223712,);
nand I_12949 (I223720,I223712,I223378);
nor I_12950 (I223222,I223720,I223528);
nor I_12951 (I223216,I223712,I223344);
DFFARX1 I_12952 (I223712,I3563,I223245,I223774,);
not I_12953 (I223782,I223774);
nor I_12954 (I223231,I223782,I223494);
not I_12955 (I223840,I3570);
DFFARX1 I_12956 (I75101,I3563,I223840,I223866,);
DFFARX1 I_12957 (I223866,I3563,I223840,I223883,);
not I_12958 (I223832,I223883);
not I_12959 (I223905,I223866);
DFFARX1 I_12960 (I75095,I3563,I223840,I223931,);
not I_12961 (I223939,I223931);
and I_12962 (I223956,I223905,I75092);
not I_12963 (I223973,I75113);
nand I_12964 (I223990,I223973,I75092);
not I_12965 (I224007,I75107);
nor I_12966 (I224024,I224007,I75098);
nand I_12967 (I224041,I224024,I75104);
nor I_12968 (I224058,I224041,I223990);
DFFARX1 I_12969 (I224058,I3563,I223840,I223808,);
not I_12970 (I224089,I224041);
not I_12971 (I224106,I75098);
nand I_12972 (I224123,I224106,I75092);
nor I_12973 (I224140,I75098,I75113);
nand I_12974 (I223820,I223956,I224140);
nand I_12975 (I223814,I223905,I75098);
nand I_12976 (I224185,I224007,I75092);
DFFARX1 I_12977 (I224185,I3563,I223840,I223829,);
DFFARX1 I_12978 (I224185,I3563,I223840,I223823,);
not I_12979 (I224230,I75092);
nor I_12980 (I224247,I224230,I75110);
and I_12981 (I224264,I224247,I75116);
or I_12982 (I224281,I224264,I75095);
DFFARX1 I_12983 (I224281,I3563,I223840,I224307,);
nand I_12984 (I224315,I224307,I223973);
nor I_12985 (I223817,I224315,I224123);
nor I_12986 (I223811,I224307,I223939);
DFFARX1 I_12987 (I224307,I3563,I223840,I224369,);
not I_12988 (I224377,I224369);
nor I_12989 (I223826,I224377,I224089);
not I_12990 (I224435,I3570);
DFFARX1 I_12991 (I1295848,I3563,I224435,I224461,);
DFFARX1 I_12992 (I224461,I3563,I224435,I224478,);
not I_12993 (I224427,I224478);
not I_12994 (I224500,I224461);
DFFARX1 I_12995 (I1295860,I3563,I224435,I224526,);
not I_12996 (I224534,I224526);
and I_12997 (I224551,I224500,I1295854);
not I_12998 (I224568,I1295866);
nand I_12999 (I224585,I224568,I1295854);
not I_13000 (I224602,I1295851);
nor I_13001 (I224619,I224602,I1295863);
nand I_13002 (I224636,I224619,I1295845);
nor I_13003 (I224653,I224636,I224585);
DFFARX1 I_13004 (I224653,I3563,I224435,I224403,);
not I_13005 (I224684,I224636);
not I_13006 (I224701,I1295863);
nand I_13007 (I224718,I224701,I1295854);
nor I_13008 (I224735,I1295863,I1295866);
nand I_13009 (I224415,I224551,I224735);
nand I_13010 (I224409,I224500,I1295863);
nand I_13011 (I224780,I224602,I1295857);
DFFARX1 I_13012 (I224780,I3563,I224435,I224424,);
DFFARX1 I_13013 (I224780,I3563,I224435,I224418,);
not I_13014 (I224825,I1295857);
nor I_13015 (I224842,I224825,I1295848);
and I_13016 (I224859,I224842,I1295845);
or I_13017 (I224876,I224859,I1295869);
DFFARX1 I_13018 (I224876,I3563,I224435,I224902,);
nand I_13019 (I224910,I224902,I224568);
nor I_13020 (I224412,I224910,I224718);
nor I_13021 (I224406,I224902,I224534);
DFFARX1 I_13022 (I224902,I3563,I224435,I224964,);
not I_13023 (I224972,I224964);
nor I_13024 (I224421,I224972,I224684);
not I_13025 (I225030,I3570);
DFFARX1 I_13026 (I395508,I3563,I225030,I225056,);
DFFARX1 I_13027 (I225056,I3563,I225030,I225073,);
not I_13028 (I225022,I225073);
not I_13029 (I225095,I225056);
DFFARX1 I_13030 (I395523,I3563,I225030,I225121,);
not I_13031 (I225129,I225121);
and I_13032 (I225146,I225095,I395520);
not I_13033 (I225163,I395508);
nand I_13034 (I225180,I225163,I395520);
not I_13035 (I225197,I395517);
nor I_13036 (I225214,I225197,I395532);
nand I_13037 (I225231,I225214,I395529);
nor I_13038 (I225248,I225231,I225180);
DFFARX1 I_13039 (I225248,I3563,I225030,I224998,);
not I_13040 (I225279,I225231);
not I_13041 (I225296,I395532);
nand I_13042 (I225313,I225296,I395520);
nor I_13043 (I225330,I395532,I395508);
nand I_13044 (I225010,I225146,I225330);
nand I_13045 (I225004,I225095,I395532);
nand I_13046 (I225375,I225197,I395526);
DFFARX1 I_13047 (I225375,I3563,I225030,I225019,);
DFFARX1 I_13048 (I225375,I3563,I225030,I225013,);
not I_13049 (I225420,I395526);
nor I_13050 (I225437,I225420,I395514);
and I_13051 (I225454,I225437,I395535);
or I_13052 (I225471,I225454,I395511);
DFFARX1 I_13053 (I225471,I3563,I225030,I225497,);
nand I_13054 (I225505,I225497,I225163);
nor I_13055 (I225007,I225505,I225313);
nor I_13056 (I225001,I225497,I225129);
DFFARX1 I_13057 (I225497,I3563,I225030,I225559,);
not I_13058 (I225567,I225559);
nor I_13059 (I225016,I225567,I225279);
not I_13060 (I225625,I3570);
DFFARX1 I_13061 (I326998,I3563,I225625,I225651,);
DFFARX1 I_13062 (I225651,I3563,I225625,I225668,);
not I_13063 (I225617,I225668);
not I_13064 (I225690,I225651);
DFFARX1 I_13065 (I327013,I3563,I225625,I225716,);
not I_13066 (I225724,I225716);
and I_13067 (I225741,I225690,I327010);
not I_13068 (I225758,I326998);
nand I_13069 (I225775,I225758,I327010);
not I_13070 (I225792,I327007);
nor I_13071 (I225809,I225792,I327022);
nand I_13072 (I225826,I225809,I327019);
nor I_13073 (I225843,I225826,I225775);
DFFARX1 I_13074 (I225843,I3563,I225625,I225593,);
not I_13075 (I225874,I225826);
not I_13076 (I225891,I327022);
nand I_13077 (I225908,I225891,I327010);
nor I_13078 (I225925,I327022,I326998);
nand I_13079 (I225605,I225741,I225925);
nand I_13080 (I225599,I225690,I327022);
nand I_13081 (I225970,I225792,I327016);
DFFARX1 I_13082 (I225970,I3563,I225625,I225614,);
DFFARX1 I_13083 (I225970,I3563,I225625,I225608,);
not I_13084 (I226015,I327016);
nor I_13085 (I226032,I226015,I327004);
and I_13086 (I226049,I226032,I327025);
or I_13087 (I226066,I226049,I327001);
DFFARX1 I_13088 (I226066,I3563,I225625,I226092,);
nand I_13089 (I226100,I226092,I225758);
nor I_13090 (I225602,I226100,I225908);
nor I_13091 (I225596,I226092,I225724);
DFFARX1 I_13092 (I226092,I3563,I225625,I226154,);
not I_13093 (I226162,I226154);
nor I_13094 (I225611,I226162,I225874);
not I_13095 (I226220,I3570);
DFFARX1 I_13096 (I798879,I3563,I226220,I226246,);
DFFARX1 I_13097 (I226246,I3563,I226220,I226263,);
not I_13098 (I226212,I226263);
not I_13099 (I226285,I226246);
DFFARX1 I_13100 (I798876,I3563,I226220,I226311,);
not I_13101 (I226319,I226311);
and I_13102 (I226336,I226285,I798882);
not I_13103 (I226353,I798867);
nand I_13104 (I226370,I226353,I798882);
not I_13105 (I226387,I798870);
nor I_13106 (I226404,I226387,I798891);
nand I_13107 (I226421,I226404,I798888);
nor I_13108 (I226438,I226421,I226370);
DFFARX1 I_13109 (I226438,I3563,I226220,I226188,);
not I_13110 (I226469,I226421);
not I_13111 (I226486,I798891);
nand I_13112 (I226503,I226486,I798882);
nor I_13113 (I226520,I798891,I798867);
nand I_13114 (I226200,I226336,I226520);
nand I_13115 (I226194,I226285,I798891);
nand I_13116 (I226565,I226387,I798867);
DFFARX1 I_13117 (I226565,I3563,I226220,I226209,);
DFFARX1 I_13118 (I226565,I3563,I226220,I226203,);
not I_13119 (I226610,I798867);
nor I_13120 (I226627,I226610,I798873);
and I_13121 (I226644,I226627,I798885);
or I_13122 (I226661,I226644,I798870);
DFFARX1 I_13123 (I226661,I3563,I226220,I226687,);
nand I_13124 (I226695,I226687,I226353);
nor I_13125 (I226197,I226695,I226503);
nor I_13126 (I226191,I226687,I226319);
DFFARX1 I_13127 (I226687,I3563,I226220,I226749,);
not I_13128 (I226757,I226749);
nor I_13129 (I226206,I226757,I226469);
not I_13130 (I226815,I3570);
DFFARX1 I_13131 (I1372009,I3563,I226815,I226841,);
DFFARX1 I_13132 (I226841,I3563,I226815,I226858,);
not I_13133 (I226807,I226858);
not I_13134 (I226880,I226841);
DFFARX1 I_13135 (I1372000,I3563,I226815,I226906,);
not I_13136 (I226914,I226906);
and I_13137 (I226931,I226880,I1371994);
not I_13138 (I226948,I1371988);
nand I_13139 (I226965,I226948,I1371994);
not I_13140 (I226982,I1372015);
nor I_13141 (I226999,I226982,I1371988);
nand I_13142 (I227016,I226999,I1372012);
nor I_13143 (I227033,I227016,I226965);
DFFARX1 I_13144 (I227033,I3563,I226815,I226783,);
not I_13145 (I227064,I227016);
not I_13146 (I227081,I1371988);
nand I_13147 (I227098,I227081,I1371994);
nor I_13148 (I227115,I1371988,I1371988);
nand I_13149 (I226795,I226931,I227115);
nand I_13150 (I226789,I226880,I1371988);
nand I_13151 (I227160,I226982,I1371997);
DFFARX1 I_13152 (I227160,I3563,I226815,I226804,);
DFFARX1 I_13153 (I227160,I3563,I226815,I226798,);
not I_13154 (I227205,I1371997);
nor I_13155 (I227222,I227205,I1372003);
and I_13156 (I227239,I227222,I1372006);
or I_13157 (I227256,I227239,I1371991);
DFFARX1 I_13158 (I227256,I3563,I226815,I227282,);
nand I_13159 (I227290,I227282,I226948);
nor I_13160 (I226792,I227290,I227098);
nor I_13161 (I226786,I227282,I226914);
DFFARX1 I_13162 (I227282,I3563,I226815,I227344,);
not I_13163 (I227352,I227344);
nor I_13164 (I226801,I227352,I227064);
not I_13165 (I227410,I3570);
DFFARX1 I_13166 (I934270,I3563,I227410,I227436,);
DFFARX1 I_13167 (I227436,I3563,I227410,I227453,);
not I_13168 (I227402,I227453);
not I_13169 (I227475,I227436);
DFFARX1 I_13170 (I934279,I3563,I227410,I227501,);
not I_13171 (I227509,I227501);
and I_13172 (I227526,I227475,I934267);
not I_13173 (I227543,I934258);
nand I_13174 (I227560,I227543,I934267);
not I_13175 (I227577,I934264);
nor I_13176 (I227594,I227577,I934282);
nand I_13177 (I227611,I227594,I934255);
nor I_13178 (I227628,I227611,I227560);
DFFARX1 I_13179 (I227628,I3563,I227410,I227378,);
not I_13180 (I227659,I227611);
not I_13181 (I227676,I934282);
nand I_13182 (I227693,I227676,I934267);
nor I_13183 (I227710,I934282,I934258);
nand I_13184 (I227390,I227526,I227710);
nand I_13185 (I227384,I227475,I934282);
nand I_13186 (I227755,I227577,I934261);
DFFARX1 I_13187 (I227755,I3563,I227410,I227399,);
DFFARX1 I_13188 (I227755,I3563,I227410,I227393,);
not I_13189 (I227800,I934261);
nor I_13190 (I227817,I227800,I934273);
and I_13191 (I227834,I227817,I934255);
or I_13192 (I227851,I227834,I934276);
DFFARX1 I_13193 (I227851,I3563,I227410,I227877,);
nand I_13194 (I227885,I227877,I227543);
nor I_13195 (I227387,I227885,I227693);
nor I_13196 (I227381,I227877,I227509);
DFFARX1 I_13197 (I227877,I3563,I227410,I227939,);
not I_13198 (I227947,I227939);
nor I_13199 (I227396,I227947,I227659);
not I_13200 (I228005,I3570);
DFFARX1 I_13201 (I2580,I3563,I228005,I228031,);
DFFARX1 I_13202 (I228031,I3563,I228005,I228048,);
not I_13203 (I227997,I228048);
not I_13204 (I228070,I228031);
DFFARX1 I_13205 (I1876,I3563,I228005,I228096,);
not I_13206 (I228104,I228096);
and I_13207 (I228121,I228070,I2828);
not I_13208 (I228138,I1420);
nand I_13209 (I228155,I228138,I2828);
not I_13210 (I228172,I2564);
nor I_13211 (I228189,I228172,I2300);
nand I_13212 (I228206,I228189,I2588);
nor I_13213 (I228223,I228206,I228155);
DFFARX1 I_13214 (I228223,I3563,I228005,I227973,);
not I_13215 (I228254,I228206);
not I_13216 (I228271,I2300);
nand I_13217 (I228288,I228271,I2828);
nor I_13218 (I228305,I2300,I1420);
nand I_13219 (I227985,I228121,I228305);
nand I_13220 (I227979,I228070,I2300);
nand I_13221 (I228350,I228172,I2388);
DFFARX1 I_13222 (I228350,I3563,I228005,I227994,);
DFFARX1 I_13223 (I228350,I3563,I228005,I227988,);
not I_13224 (I228395,I2388);
nor I_13225 (I228412,I228395,I3212);
and I_13226 (I228429,I228412,I2732);
or I_13227 (I228446,I228429,I1948);
DFFARX1 I_13228 (I228446,I3563,I228005,I228472,);
nand I_13229 (I228480,I228472,I228138);
nor I_13230 (I227982,I228480,I228288);
nor I_13231 (I227976,I228472,I228104);
DFFARX1 I_13232 (I228472,I3563,I228005,I228534,);
not I_13233 (I228542,I228534);
nor I_13234 (I227991,I228542,I228254);
not I_13235 (I228600,I3570);
DFFARX1 I_13236 (I497498,I3563,I228600,I228626,);
DFFARX1 I_13237 (I228626,I3563,I228600,I228643,);
not I_13238 (I228592,I228643);
not I_13239 (I228665,I228626);
DFFARX1 I_13240 (I497486,I3563,I228600,I228691,);
not I_13241 (I228699,I228691);
and I_13242 (I228716,I228665,I497495);
not I_13243 (I228733,I497492);
nand I_13244 (I228750,I228733,I497495);
not I_13245 (I228767,I497483);
nor I_13246 (I228784,I228767,I497489);
nand I_13247 (I228801,I228784,I497474);
nor I_13248 (I228818,I228801,I228750);
DFFARX1 I_13249 (I228818,I3563,I228600,I228568,);
not I_13250 (I228849,I228801);
not I_13251 (I228866,I497489);
nand I_13252 (I228883,I228866,I497495);
nor I_13253 (I228900,I497489,I497492);
nand I_13254 (I228580,I228716,I228900);
nand I_13255 (I228574,I228665,I497489);
nand I_13256 (I228945,I228767,I497474);
DFFARX1 I_13257 (I228945,I3563,I228600,I228589,);
DFFARX1 I_13258 (I228945,I3563,I228600,I228583,);
not I_13259 (I228990,I497474);
nor I_13260 (I229007,I228990,I497480);
and I_13261 (I229024,I229007,I497477);
or I_13262 (I229041,I229024,I497501);
DFFARX1 I_13263 (I229041,I3563,I228600,I229067,);
nand I_13264 (I229075,I229067,I228733);
nor I_13265 (I228577,I229075,I228883);
nor I_13266 (I228571,I229067,I228699);
DFFARX1 I_13267 (I229067,I3563,I228600,I229129,);
not I_13268 (I229137,I229129);
nor I_13269 (I228586,I229137,I228849);
not I_13270 (I229195,I3570);
DFFARX1 I_13271 (I104613,I3563,I229195,I229221,);
DFFARX1 I_13272 (I229221,I3563,I229195,I229238,);
not I_13273 (I229187,I229238);
not I_13274 (I229260,I229221);
DFFARX1 I_13275 (I104607,I3563,I229195,I229286,);
not I_13276 (I229294,I229286);
and I_13277 (I229311,I229260,I104604);
not I_13278 (I229328,I104625);
nand I_13279 (I229345,I229328,I104604);
not I_13280 (I229362,I104619);
nor I_13281 (I229379,I229362,I104610);
nand I_13282 (I229396,I229379,I104616);
nor I_13283 (I229413,I229396,I229345);
DFFARX1 I_13284 (I229413,I3563,I229195,I229163,);
not I_13285 (I229444,I229396);
not I_13286 (I229461,I104610);
nand I_13287 (I229478,I229461,I104604);
nor I_13288 (I229495,I104610,I104625);
nand I_13289 (I229175,I229311,I229495);
nand I_13290 (I229169,I229260,I104610);
nand I_13291 (I229540,I229362,I104604);
DFFARX1 I_13292 (I229540,I3563,I229195,I229184,);
DFFARX1 I_13293 (I229540,I3563,I229195,I229178,);
not I_13294 (I229585,I104604);
nor I_13295 (I229602,I229585,I104622);
and I_13296 (I229619,I229602,I104628);
or I_13297 (I229636,I229619,I104607);
DFFARX1 I_13298 (I229636,I3563,I229195,I229662,);
nand I_13299 (I229670,I229662,I229328);
nor I_13300 (I229172,I229670,I229478);
nor I_13301 (I229166,I229662,I229294);
DFFARX1 I_13302 (I229662,I3563,I229195,I229724,);
not I_13303 (I229732,I229724);
nor I_13304 (I229181,I229732,I229444);
not I_13305 (I229790,I3570);
DFFARX1 I_13306 (I647446,I3563,I229790,I229816,);
DFFARX1 I_13307 (I229816,I3563,I229790,I229833,);
not I_13308 (I229782,I229833);
not I_13309 (I229855,I229816);
DFFARX1 I_13310 (I647437,I3563,I229790,I229881,);
not I_13311 (I229889,I229881);
and I_13312 (I229906,I229855,I647455);
not I_13313 (I229923,I647452);
nand I_13314 (I229940,I229923,I647455);
not I_13315 (I229957,I647431);
nor I_13316 (I229974,I229957,I647434);
nand I_13317 (I229991,I229974,I647443);
nor I_13318 (I230008,I229991,I229940);
DFFARX1 I_13319 (I230008,I3563,I229790,I229758,);
not I_13320 (I230039,I229991);
not I_13321 (I230056,I647434);
nand I_13322 (I230073,I230056,I647455);
nor I_13323 (I230090,I647434,I647452);
nand I_13324 (I229770,I229906,I230090);
nand I_13325 (I229764,I229855,I647434);
nand I_13326 (I230135,I229957,I647449);
DFFARX1 I_13327 (I230135,I3563,I229790,I229779,);
DFFARX1 I_13328 (I230135,I3563,I229790,I229773,);
not I_13329 (I230180,I647449);
nor I_13330 (I230197,I230180,I647431);
and I_13331 (I230214,I230197,I647440);
or I_13332 (I230231,I230214,I647434);
DFFARX1 I_13333 (I230231,I3563,I229790,I230257,);
nand I_13334 (I230265,I230257,I229923);
nor I_13335 (I229767,I230265,I230073);
nor I_13336 (I229761,I230257,I229889);
DFFARX1 I_13337 (I230257,I3563,I229790,I230319,);
not I_13338 (I230327,I230319);
nor I_13339 (I229776,I230327,I230039);
not I_13340 (I230385,I3570);
DFFARX1 I_13341 (I758997,I3563,I230385,I230411,);
DFFARX1 I_13342 (I230411,I3563,I230385,I230428,);
not I_13343 (I230377,I230428);
not I_13344 (I230450,I230411);
DFFARX1 I_13345 (I758994,I3563,I230385,I230476,);
not I_13346 (I230484,I230476);
and I_13347 (I230501,I230450,I759000);
not I_13348 (I230518,I758985);
nand I_13349 (I230535,I230518,I759000);
not I_13350 (I230552,I758988);
nor I_13351 (I230569,I230552,I759009);
nand I_13352 (I230586,I230569,I759006);
nor I_13353 (I230603,I230586,I230535);
DFFARX1 I_13354 (I230603,I3563,I230385,I230353,);
not I_13355 (I230634,I230586);
not I_13356 (I230651,I759009);
nand I_13357 (I230668,I230651,I759000);
nor I_13358 (I230685,I759009,I758985);
nand I_13359 (I230365,I230501,I230685);
nand I_13360 (I230359,I230450,I759009);
nand I_13361 (I230730,I230552,I758985);
DFFARX1 I_13362 (I230730,I3563,I230385,I230374,);
DFFARX1 I_13363 (I230730,I3563,I230385,I230368,);
not I_13364 (I230775,I758985);
nor I_13365 (I230792,I230775,I758991);
and I_13366 (I230809,I230792,I759003);
or I_13367 (I230826,I230809,I758988);
DFFARX1 I_13368 (I230826,I3563,I230385,I230852,);
nand I_13369 (I230860,I230852,I230518);
nor I_13370 (I230362,I230860,I230668);
nor I_13371 (I230356,I230852,I230484);
DFFARX1 I_13372 (I230852,I3563,I230385,I230914,);
not I_13373 (I230922,I230914);
nor I_13374 (I230371,I230922,I230634);
not I_13375 (I230980,I3570);
DFFARX1 I_13376 (I1294114,I3563,I230980,I231006,);
DFFARX1 I_13377 (I231006,I3563,I230980,I231023,);
not I_13378 (I230972,I231023);
not I_13379 (I231045,I231006);
DFFARX1 I_13380 (I1294126,I3563,I230980,I231071,);
not I_13381 (I231079,I231071);
and I_13382 (I231096,I231045,I1294120);
not I_13383 (I231113,I1294132);
nand I_13384 (I231130,I231113,I1294120);
not I_13385 (I231147,I1294117);
nor I_13386 (I231164,I231147,I1294129);
nand I_13387 (I231181,I231164,I1294111);
nor I_13388 (I231198,I231181,I231130);
DFFARX1 I_13389 (I231198,I3563,I230980,I230948,);
not I_13390 (I231229,I231181);
not I_13391 (I231246,I1294129);
nand I_13392 (I231263,I231246,I1294120);
nor I_13393 (I231280,I1294129,I1294132);
nand I_13394 (I230960,I231096,I231280);
nand I_13395 (I230954,I231045,I1294129);
nand I_13396 (I231325,I231147,I1294123);
DFFARX1 I_13397 (I231325,I3563,I230980,I230969,);
DFFARX1 I_13398 (I231325,I3563,I230980,I230963,);
not I_13399 (I231370,I1294123);
nor I_13400 (I231387,I231370,I1294114);
and I_13401 (I231404,I231387,I1294111);
or I_13402 (I231421,I231404,I1294135);
DFFARX1 I_13403 (I231421,I3563,I230980,I231447,);
nand I_13404 (I231455,I231447,I231113);
nor I_13405 (I230957,I231455,I231263);
nor I_13406 (I230951,I231447,I231079);
DFFARX1 I_13407 (I231447,I3563,I230980,I231509,);
not I_13408 (I231517,I231509);
nor I_13409 (I230966,I231517,I231229);
not I_13410 (I231575,I3570);
DFFARX1 I_13411 (I553688,I3563,I231575,I231601,);
DFFARX1 I_13412 (I231601,I3563,I231575,I231618,);
not I_13413 (I231567,I231618);
not I_13414 (I231640,I231601);
DFFARX1 I_13415 (I553682,I3563,I231575,I231666,);
not I_13416 (I231674,I231666);
and I_13417 (I231691,I231640,I553697);
not I_13418 (I231708,I553694);
nand I_13419 (I231725,I231708,I553697);
not I_13420 (I231742,I553685);
nor I_13421 (I231759,I231742,I553676);
nand I_13422 (I231776,I231759,I553679);
nor I_13423 (I231793,I231776,I231725);
DFFARX1 I_13424 (I231793,I3563,I231575,I231543,);
not I_13425 (I231824,I231776);
not I_13426 (I231841,I553676);
nand I_13427 (I231858,I231841,I553697);
nor I_13428 (I231875,I553676,I553694);
nand I_13429 (I231555,I231691,I231875);
nand I_13430 (I231549,I231640,I553676);
nand I_13431 (I231920,I231742,I553700);
DFFARX1 I_13432 (I231920,I3563,I231575,I231564,);
DFFARX1 I_13433 (I231920,I3563,I231575,I231558,);
not I_13434 (I231965,I553700);
nor I_13435 (I231982,I231965,I553691);
and I_13436 (I231999,I231982,I553676);
or I_13437 (I232016,I231999,I553679);
DFFARX1 I_13438 (I232016,I3563,I231575,I232042,);
nand I_13439 (I232050,I232042,I231708);
nor I_13440 (I231552,I232050,I231858);
nor I_13441 (I231546,I232042,I231674);
DFFARX1 I_13442 (I232042,I3563,I231575,I232104,);
not I_13443 (I232112,I232104);
nor I_13444 (I231561,I232112,I231824);
not I_13445 (I232170,I3570);
DFFARX1 I_13446 (I96181,I3563,I232170,I232196,);
DFFARX1 I_13447 (I232196,I3563,I232170,I232213,);
not I_13448 (I232162,I232213);
not I_13449 (I232235,I232196);
DFFARX1 I_13450 (I96175,I3563,I232170,I232261,);
not I_13451 (I232269,I232261);
and I_13452 (I232286,I232235,I96172);
not I_13453 (I232303,I96193);
nand I_13454 (I232320,I232303,I96172);
not I_13455 (I232337,I96187);
nor I_13456 (I232354,I232337,I96178);
nand I_13457 (I232371,I232354,I96184);
nor I_13458 (I232388,I232371,I232320);
DFFARX1 I_13459 (I232388,I3563,I232170,I232138,);
not I_13460 (I232419,I232371);
not I_13461 (I232436,I96178);
nand I_13462 (I232453,I232436,I96172);
nor I_13463 (I232470,I96178,I96193);
nand I_13464 (I232150,I232286,I232470);
nand I_13465 (I232144,I232235,I96178);
nand I_13466 (I232515,I232337,I96172);
DFFARX1 I_13467 (I232515,I3563,I232170,I232159,);
DFFARX1 I_13468 (I232515,I3563,I232170,I232153,);
not I_13469 (I232560,I96172);
nor I_13470 (I232577,I232560,I96190);
and I_13471 (I232594,I232577,I96196);
or I_13472 (I232611,I232594,I96175);
DFFARX1 I_13473 (I232611,I3563,I232170,I232637,);
nand I_13474 (I232645,I232637,I232303);
nor I_13475 (I232147,I232645,I232453);
nor I_13476 (I232141,I232637,I232269);
DFFARX1 I_13477 (I232637,I3563,I232170,I232699,);
not I_13478 (I232707,I232699);
nor I_13479 (I232156,I232707,I232419);
not I_13480 (I232765,I3570);
DFFARX1 I_13481 (I833196,I3563,I232765,I232791,);
DFFARX1 I_13482 (I232791,I3563,I232765,I232808,);
not I_13483 (I232757,I232808);
not I_13484 (I232830,I232791);
DFFARX1 I_13485 (I833190,I3563,I232765,I232856,);
not I_13486 (I232864,I232856);
and I_13487 (I232881,I232830,I833208);
not I_13488 (I232898,I833196);
nand I_13489 (I232915,I232898,I833208);
not I_13490 (I232932,I833190);
nor I_13491 (I232949,I232932,I833202);
nand I_13492 (I232966,I232949,I833193);
nor I_13493 (I232983,I232966,I232915);
DFFARX1 I_13494 (I232983,I3563,I232765,I232733,);
not I_13495 (I233014,I232966);
not I_13496 (I233031,I833202);
nand I_13497 (I233048,I233031,I833208);
nor I_13498 (I233065,I833202,I833196);
nand I_13499 (I232745,I232881,I233065);
nand I_13500 (I232739,I232830,I833202);
nand I_13501 (I233110,I232932,I833205);
DFFARX1 I_13502 (I233110,I3563,I232765,I232754,);
DFFARX1 I_13503 (I233110,I3563,I232765,I232748,);
not I_13504 (I233155,I833205);
nor I_13505 (I233172,I233155,I833211);
and I_13506 (I233189,I233172,I833193);
or I_13507 (I233206,I233189,I833199);
DFFARX1 I_13508 (I233206,I3563,I232765,I233232,);
nand I_13509 (I233240,I233232,I232898);
nor I_13510 (I232742,I233240,I233048);
nor I_13511 (I232736,I233232,I232864);
DFFARX1 I_13512 (I233232,I3563,I232765,I233294,);
not I_13513 (I233302,I233294);
nor I_13514 (I232751,I233302,I233014);
not I_13515 (I233360,I3570);
DFFARX1 I_13516 (I125166,I3563,I233360,I233386,);
DFFARX1 I_13517 (I233386,I3563,I233360,I233403,);
not I_13518 (I233352,I233403);
not I_13519 (I233425,I233386);
DFFARX1 I_13520 (I125160,I3563,I233360,I233451,);
not I_13521 (I233459,I233451);
and I_13522 (I233476,I233425,I125157);
not I_13523 (I233493,I125178);
nand I_13524 (I233510,I233493,I125157);
not I_13525 (I233527,I125172);
nor I_13526 (I233544,I233527,I125163);
nand I_13527 (I233561,I233544,I125169);
nor I_13528 (I233578,I233561,I233510);
DFFARX1 I_13529 (I233578,I3563,I233360,I233328,);
not I_13530 (I233609,I233561);
not I_13531 (I233626,I125163);
nand I_13532 (I233643,I233626,I125157);
nor I_13533 (I233660,I125163,I125178);
nand I_13534 (I233340,I233476,I233660);
nand I_13535 (I233334,I233425,I125163);
nand I_13536 (I233705,I233527,I125157);
DFFARX1 I_13537 (I233705,I3563,I233360,I233349,);
DFFARX1 I_13538 (I233705,I3563,I233360,I233343,);
not I_13539 (I233750,I125157);
nor I_13540 (I233767,I233750,I125175);
and I_13541 (I233784,I233767,I125181);
or I_13542 (I233801,I233784,I125160);
DFFARX1 I_13543 (I233801,I3563,I233360,I233827,);
nand I_13544 (I233835,I233827,I233493);
nor I_13545 (I233337,I233835,I233643);
nor I_13546 (I233331,I233827,I233459);
DFFARX1 I_13547 (I233827,I3563,I233360,I233889,);
not I_13548 (I233897,I233889);
nor I_13549 (I233346,I233897,I233609);
not I_13550 (I233955,I3570);
DFFARX1 I_13551 (I1101399,I3563,I233955,I233981,);
DFFARX1 I_13552 (I233981,I3563,I233955,I233998,);
not I_13553 (I233947,I233998);
not I_13554 (I234020,I233981);
DFFARX1 I_13555 (I1101399,I3563,I233955,I234046,);
not I_13556 (I234054,I234046);
and I_13557 (I234071,I234020,I1101402);
not I_13558 (I234088,I1101414);
nand I_13559 (I234105,I234088,I1101402);
not I_13560 (I234122,I1101420);
nor I_13561 (I234139,I234122,I1101411);
nand I_13562 (I234156,I234139,I1101417);
nor I_13563 (I234173,I234156,I234105);
DFFARX1 I_13564 (I234173,I3563,I233955,I233923,);
not I_13565 (I234204,I234156);
not I_13566 (I234221,I1101411);
nand I_13567 (I234238,I234221,I1101402);
nor I_13568 (I234255,I1101411,I1101414);
nand I_13569 (I233935,I234071,I234255);
nand I_13570 (I233929,I234020,I1101411);
nand I_13571 (I234300,I234122,I1101408);
DFFARX1 I_13572 (I234300,I3563,I233955,I233944,);
DFFARX1 I_13573 (I234300,I3563,I233955,I233938,);
not I_13574 (I234345,I1101408);
nor I_13575 (I234362,I234345,I1101405);
and I_13576 (I234379,I234362,I1101423);
or I_13577 (I234396,I234379,I1101402);
DFFARX1 I_13578 (I234396,I3563,I233955,I234422,);
nand I_13579 (I234430,I234422,I234088);
nor I_13580 (I233932,I234430,I234238);
nor I_13581 (I233926,I234422,I234054);
DFFARX1 I_13582 (I234422,I3563,I233955,I234484,);
not I_13583 (I234492,I234484);
nor I_13584 (I233941,I234492,I234204);
not I_13585 (I234550,I3570);
DFFARX1 I_13586 (I907503,I3563,I234550,I234576,);
DFFARX1 I_13587 (I234576,I3563,I234550,I234593,);
not I_13588 (I234542,I234593);
not I_13589 (I234615,I234576);
DFFARX1 I_13590 (I907497,I3563,I234550,I234641,);
not I_13591 (I234649,I234641);
and I_13592 (I234666,I234615,I907515);
not I_13593 (I234683,I907503);
nand I_13594 (I234700,I234683,I907515);
not I_13595 (I234717,I907497);
nor I_13596 (I234734,I234717,I907509);
nand I_13597 (I234751,I234734,I907500);
nor I_13598 (I234768,I234751,I234700);
DFFARX1 I_13599 (I234768,I3563,I234550,I234518,);
not I_13600 (I234799,I234751);
not I_13601 (I234816,I907509);
nand I_13602 (I234833,I234816,I907515);
nor I_13603 (I234850,I907509,I907503);
nand I_13604 (I234530,I234666,I234850);
nand I_13605 (I234524,I234615,I907509);
nand I_13606 (I234895,I234717,I907512);
DFFARX1 I_13607 (I234895,I3563,I234550,I234539,);
DFFARX1 I_13608 (I234895,I3563,I234550,I234533,);
not I_13609 (I234940,I907512);
nor I_13610 (I234957,I234940,I907518);
and I_13611 (I234974,I234957,I907500);
or I_13612 (I234991,I234974,I907506);
DFFARX1 I_13613 (I234991,I3563,I234550,I235017,);
nand I_13614 (I235025,I235017,I234683);
nor I_13615 (I234527,I235025,I234833);
nor I_13616 (I234521,I235017,I234649);
DFFARX1 I_13617 (I235017,I3563,I234550,I235079,);
not I_13618 (I235087,I235079);
nor I_13619 (I234536,I235087,I234799);
not I_13620 (I235145,I3570);
DFFARX1 I_13621 (I457786,I3563,I235145,I235171,);
DFFARX1 I_13622 (I235171,I3563,I235145,I235188,);
not I_13623 (I235137,I235188);
not I_13624 (I235210,I235171);
DFFARX1 I_13625 (I457774,I3563,I235145,I235236,);
not I_13626 (I235244,I235236);
and I_13627 (I235261,I235210,I457783);
not I_13628 (I235278,I457780);
nand I_13629 (I235295,I235278,I457783);
not I_13630 (I235312,I457771);
nor I_13631 (I235329,I235312,I457777);
nand I_13632 (I235346,I235329,I457762);
nor I_13633 (I235363,I235346,I235295);
DFFARX1 I_13634 (I235363,I3563,I235145,I235113,);
not I_13635 (I235394,I235346);
not I_13636 (I235411,I457777);
nand I_13637 (I235428,I235411,I457783);
nor I_13638 (I235445,I457777,I457780);
nand I_13639 (I235125,I235261,I235445);
nand I_13640 (I235119,I235210,I457777);
nand I_13641 (I235490,I235312,I457762);
DFFARX1 I_13642 (I235490,I3563,I235145,I235134,);
DFFARX1 I_13643 (I235490,I3563,I235145,I235128,);
not I_13644 (I235535,I457762);
nor I_13645 (I235552,I235535,I457768);
and I_13646 (I235569,I235552,I457765);
or I_13647 (I235586,I235569,I457789);
DFFARX1 I_13648 (I235586,I3563,I235145,I235612,);
nand I_13649 (I235620,I235612,I235278);
nor I_13650 (I235122,I235620,I235428);
nor I_13651 (I235116,I235612,I235244);
DFFARX1 I_13652 (I235612,I3563,I235145,I235674,);
not I_13653 (I235682,I235674);
nor I_13654 (I235131,I235682,I235394);
not I_13655 (I235740,I3570);
DFFARX1 I_13656 (I503482,I3563,I235740,I235766,);
DFFARX1 I_13657 (I235766,I3563,I235740,I235783,);
not I_13658 (I235732,I235783);
not I_13659 (I235805,I235766);
DFFARX1 I_13660 (I503470,I3563,I235740,I235831,);
not I_13661 (I235839,I235831);
and I_13662 (I235856,I235805,I503479);
not I_13663 (I235873,I503476);
nand I_13664 (I235890,I235873,I503479);
not I_13665 (I235907,I503467);
nor I_13666 (I235924,I235907,I503473);
nand I_13667 (I235941,I235924,I503458);
nor I_13668 (I235958,I235941,I235890);
DFFARX1 I_13669 (I235958,I3563,I235740,I235708,);
not I_13670 (I235989,I235941);
not I_13671 (I236006,I503473);
nand I_13672 (I236023,I236006,I503479);
nor I_13673 (I236040,I503473,I503476);
nand I_13674 (I235720,I235856,I236040);
nand I_13675 (I235714,I235805,I503473);
nand I_13676 (I236085,I235907,I503458);
DFFARX1 I_13677 (I236085,I3563,I235740,I235729,);
DFFARX1 I_13678 (I236085,I3563,I235740,I235723,);
not I_13679 (I236130,I503458);
nor I_13680 (I236147,I236130,I503464);
and I_13681 (I236164,I236147,I503461);
or I_13682 (I236181,I236164,I503485);
DFFARX1 I_13683 (I236181,I3563,I235740,I236207,);
nand I_13684 (I236215,I236207,I235873);
nor I_13685 (I235717,I236215,I236023);
nor I_13686 (I235711,I236207,I235839);
DFFARX1 I_13687 (I236207,I3563,I235740,I236269,);
not I_13688 (I236277,I236269);
nor I_13689 (I235726,I236277,I235989);
not I_13690 (I236335,I3570);
DFFARX1 I_13691 (I946544,I3563,I236335,I236361,);
DFFARX1 I_13692 (I236361,I3563,I236335,I236378,);
not I_13693 (I236327,I236378);
not I_13694 (I236400,I236361);
DFFARX1 I_13695 (I946553,I3563,I236335,I236426,);
not I_13696 (I236434,I236426);
and I_13697 (I236451,I236400,I946541);
not I_13698 (I236468,I946532);
nand I_13699 (I236485,I236468,I946541);
not I_13700 (I236502,I946538);
nor I_13701 (I236519,I236502,I946556);
nand I_13702 (I236536,I236519,I946529);
nor I_13703 (I236553,I236536,I236485);
DFFARX1 I_13704 (I236553,I3563,I236335,I236303,);
not I_13705 (I236584,I236536);
not I_13706 (I236601,I946556);
nand I_13707 (I236618,I236601,I946541);
nor I_13708 (I236635,I946556,I946532);
nand I_13709 (I236315,I236451,I236635);
nand I_13710 (I236309,I236400,I946556);
nand I_13711 (I236680,I236502,I946535);
DFFARX1 I_13712 (I236680,I3563,I236335,I236324,);
DFFARX1 I_13713 (I236680,I3563,I236335,I236318,);
not I_13714 (I236725,I946535);
nor I_13715 (I236742,I236725,I946547);
and I_13716 (I236759,I236742,I946529);
or I_13717 (I236776,I236759,I946550);
DFFARX1 I_13718 (I236776,I3563,I236335,I236802,);
nand I_13719 (I236810,I236802,I236468);
nor I_13720 (I236312,I236810,I236618);
nor I_13721 (I236306,I236802,I236434);
DFFARX1 I_13722 (I236802,I3563,I236335,I236864,);
not I_13723 (I236872,I236864);
nor I_13724 (I236321,I236872,I236584);
not I_13725 (I236930,I3570);
DFFARX1 I_13726 (I1102555,I3563,I236930,I236956,);
DFFARX1 I_13727 (I236956,I3563,I236930,I236973,);
not I_13728 (I236922,I236973);
not I_13729 (I236995,I236956);
DFFARX1 I_13730 (I1102555,I3563,I236930,I237021,);
not I_13731 (I237029,I237021);
and I_13732 (I237046,I236995,I1102558);
not I_13733 (I237063,I1102570);
nand I_13734 (I237080,I237063,I1102558);
not I_13735 (I237097,I1102576);
nor I_13736 (I237114,I237097,I1102567);
nand I_13737 (I237131,I237114,I1102573);
nor I_13738 (I237148,I237131,I237080);
DFFARX1 I_13739 (I237148,I3563,I236930,I236898,);
not I_13740 (I237179,I237131);
not I_13741 (I237196,I1102567);
nand I_13742 (I237213,I237196,I1102558);
nor I_13743 (I237230,I1102567,I1102570);
nand I_13744 (I236910,I237046,I237230);
nand I_13745 (I236904,I236995,I1102567);
nand I_13746 (I237275,I237097,I1102564);
DFFARX1 I_13747 (I237275,I3563,I236930,I236919,);
DFFARX1 I_13748 (I237275,I3563,I236930,I236913,);
not I_13749 (I237320,I1102564);
nor I_13750 (I237337,I237320,I1102561);
and I_13751 (I237354,I237337,I1102579);
or I_13752 (I237371,I237354,I1102558);
DFFARX1 I_13753 (I237371,I3563,I236930,I237397,);
nand I_13754 (I237405,I237397,I237063);
nor I_13755 (I236907,I237405,I237213);
nor I_13756 (I236901,I237397,I237029);
DFFARX1 I_13757 (I237397,I3563,I236930,I237459,);
not I_13758 (I237467,I237459);
nor I_13759 (I236916,I237467,I237179);
not I_13760 (I237525,I3570);
DFFARX1 I_13761 (I737611,I3563,I237525,I237551,);
DFFARX1 I_13762 (I237551,I3563,I237525,I237568,);
not I_13763 (I237517,I237568);
not I_13764 (I237590,I237551);
DFFARX1 I_13765 (I737608,I3563,I237525,I237616,);
not I_13766 (I237624,I237616);
and I_13767 (I237641,I237590,I737614);
not I_13768 (I237658,I737599);
nand I_13769 (I237675,I237658,I737614);
not I_13770 (I237692,I737602);
nor I_13771 (I237709,I237692,I737623);
nand I_13772 (I237726,I237709,I737620);
nor I_13773 (I237743,I237726,I237675);
DFFARX1 I_13774 (I237743,I3563,I237525,I237493,);
not I_13775 (I237774,I237726);
not I_13776 (I237791,I737623);
nand I_13777 (I237808,I237791,I737614);
nor I_13778 (I237825,I737623,I737599);
nand I_13779 (I237505,I237641,I237825);
nand I_13780 (I237499,I237590,I737623);
nand I_13781 (I237870,I237692,I737599);
DFFARX1 I_13782 (I237870,I3563,I237525,I237514,);
DFFARX1 I_13783 (I237870,I3563,I237525,I237508,);
not I_13784 (I237915,I737599);
nor I_13785 (I237932,I237915,I737605);
and I_13786 (I237949,I237932,I737617);
or I_13787 (I237966,I237949,I737602);
DFFARX1 I_13788 (I237966,I3563,I237525,I237992,);
nand I_13789 (I238000,I237992,I237658);
nor I_13790 (I237502,I238000,I237808);
nor I_13791 (I237496,I237992,I237624);
DFFARX1 I_13792 (I237992,I3563,I237525,I238054,);
not I_13793 (I238062,I238054);
nor I_13794 (I237511,I238062,I237774);
not I_13795 (I238120,I3570);
DFFARX1 I_13796 (I1323592,I3563,I238120,I238146,);
DFFARX1 I_13797 (I238146,I3563,I238120,I238163,);
not I_13798 (I238112,I238163);
not I_13799 (I238185,I238146);
DFFARX1 I_13800 (I1323604,I3563,I238120,I238211,);
not I_13801 (I238219,I238211);
and I_13802 (I238236,I238185,I1323598);
not I_13803 (I238253,I1323610);
nand I_13804 (I238270,I238253,I1323598);
not I_13805 (I238287,I1323595);
nor I_13806 (I238304,I238287,I1323607);
nand I_13807 (I238321,I238304,I1323589);
nor I_13808 (I238338,I238321,I238270);
DFFARX1 I_13809 (I238338,I3563,I238120,I238088,);
not I_13810 (I238369,I238321);
not I_13811 (I238386,I1323607);
nand I_13812 (I238403,I238386,I1323598);
nor I_13813 (I238420,I1323607,I1323610);
nand I_13814 (I238100,I238236,I238420);
nand I_13815 (I238094,I238185,I1323607);
nand I_13816 (I238465,I238287,I1323601);
DFFARX1 I_13817 (I238465,I3563,I238120,I238109,);
DFFARX1 I_13818 (I238465,I3563,I238120,I238103,);
not I_13819 (I238510,I1323601);
nor I_13820 (I238527,I238510,I1323592);
and I_13821 (I238544,I238527,I1323589);
or I_13822 (I238561,I238544,I1323613);
DFFARX1 I_13823 (I238561,I3563,I238120,I238587,);
nand I_13824 (I238595,I238587,I238253);
nor I_13825 (I238097,I238595,I238403);
nor I_13826 (I238091,I238587,I238219);
DFFARX1 I_13827 (I238587,I3563,I238120,I238649,);
not I_13828 (I238657,I238649);
nor I_13829 (I238106,I238657,I238369);
not I_13830 (I238715,I3570);
DFFARX1 I_13831 (I729519,I3563,I238715,I238741,);
DFFARX1 I_13832 (I238741,I3563,I238715,I238758,);
not I_13833 (I238707,I238758);
not I_13834 (I238780,I238741);
DFFARX1 I_13835 (I729516,I3563,I238715,I238806,);
not I_13836 (I238814,I238806);
and I_13837 (I238831,I238780,I729522);
not I_13838 (I238848,I729507);
nand I_13839 (I238865,I238848,I729522);
not I_13840 (I238882,I729510);
nor I_13841 (I238899,I238882,I729531);
nand I_13842 (I238916,I238899,I729528);
nor I_13843 (I238933,I238916,I238865);
DFFARX1 I_13844 (I238933,I3563,I238715,I238683,);
not I_13845 (I238964,I238916);
not I_13846 (I238981,I729531);
nand I_13847 (I238998,I238981,I729522);
nor I_13848 (I239015,I729531,I729507);
nand I_13849 (I238695,I238831,I239015);
nand I_13850 (I238689,I238780,I729531);
nand I_13851 (I239060,I238882,I729507);
DFFARX1 I_13852 (I239060,I3563,I238715,I238704,);
DFFARX1 I_13853 (I239060,I3563,I238715,I238698,);
not I_13854 (I239105,I729507);
nor I_13855 (I239122,I239105,I729513);
and I_13856 (I239139,I239122,I729525);
or I_13857 (I239156,I239139,I729510);
DFFARX1 I_13858 (I239156,I3563,I238715,I239182,);
nand I_13859 (I239190,I239182,I238848);
nor I_13860 (I238692,I239190,I238998);
nor I_13861 (I238686,I239182,I238814);
DFFARX1 I_13862 (I239182,I3563,I238715,I239244,);
not I_13863 (I239252,I239244);
nor I_13864 (I238701,I239252,I238964);
not I_13865 (I239310,I3570);
DFFARX1 I_13866 (I641088,I3563,I239310,I239336,);
DFFARX1 I_13867 (I239336,I3563,I239310,I239353,);
not I_13868 (I239302,I239353);
not I_13869 (I239375,I239336);
DFFARX1 I_13870 (I641079,I3563,I239310,I239401,);
not I_13871 (I239409,I239401);
and I_13872 (I239426,I239375,I641097);
not I_13873 (I239443,I641094);
nand I_13874 (I239460,I239443,I641097);
not I_13875 (I239477,I641073);
nor I_13876 (I239494,I239477,I641076);
nand I_13877 (I239511,I239494,I641085);
nor I_13878 (I239528,I239511,I239460);
DFFARX1 I_13879 (I239528,I3563,I239310,I239278,);
not I_13880 (I239559,I239511);
not I_13881 (I239576,I641076);
nand I_13882 (I239593,I239576,I641097);
nor I_13883 (I239610,I641076,I641094);
nand I_13884 (I239290,I239426,I239610);
nand I_13885 (I239284,I239375,I641076);
nand I_13886 (I239655,I239477,I641091);
DFFARX1 I_13887 (I239655,I3563,I239310,I239299,);
DFFARX1 I_13888 (I239655,I3563,I239310,I239293,);
not I_13889 (I239700,I641091);
nor I_13890 (I239717,I239700,I641073);
and I_13891 (I239734,I239717,I641082);
or I_13892 (I239751,I239734,I641076);
DFFARX1 I_13893 (I239751,I3563,I239310,I239777,);
nand I_13894 (I239785,I239777,I239443);
nor I_13895 (I239287,I239785,I239593);
nor I_13896 (I239281,I239777,I239409);
DFFARX1 I_13897 (I239777,I3563,I239310,I239839,);
not I_13898 (I239847,I239839);
nor I_13899 (I239296,I239847,I239559);
not I_13900 (I239905,I3570);
DFFARX1 I_13901 (I535243,I3563,I239905,I239931,);
DFFARX1 I_13902 (I239931,I3563,I239905,I239948,);
not I_13903 (I239897,I239948);
not I_13904 (I239970,I239931);
DFFARX1 I_13905 (I535237,I3563,I239905,I239996,);
not I_13906 (I240004,I239996);
and I_13907 (I240021,I239970,I535252);
not I_13908 (I240038,I535249);
nand I_13909 (I240055,I240038,I535252);
not I_13910 (I240072,I535240);
nor I_13911 (I240089,I240072,I535231);
nand I_13912 (I240106,I240089,I535234);
nor I_13913 (I240123,I240106,I240055);
DFFARX1 I_13914 (I240123,I3563,I239905,I239873,);
not I_13915 (I240154,I240106);
not I_13916 (I240171,I535231);
nand I_13917 (I240188,I240171,I535252);
nor I_13918 (I240205,I535231,I535249);
nand I_13919 (I239885,I240021,I240205);
nand I_13920 (I239879,I239970,I535231);
nand I_13921 (I240250,I240072,I535255);
DFFARX1 I_13922 (I240250,I3563,I239905,I239894,);
DFFARX1 I_13923 (I240250,I3563,I239905,I239888,);
not I_13924 (I240295,I535255);
nor I_13925 (I240312,I240295,I535246);
and I_13926 (I240329,I240312,I535231);
or I_13927 (I240346,I240329,I535234);
DFFARX1 I_13928 (I240346,I3563,I239905,I240372,);
nand I_13929 (I240380,I240372,I240038);
nor I_13930 (I239882,I240380,I240188);
nor I_13931 (I239876,I240372,I240004);
DFFARX1 I_13932 (I240372,I3563,I239905,I240434,);
not I_13933 (I240442,I240434);
nor I_13934 (I239891,I240442,I240154);
not I_13935 (I240500,I3570);
DFFARX1 I_13936 (I586178,I3563,I240500,I240526,);
DFFARX1 I_13937 (I240526,I3563,I240500,I240543,);
not I_13938 (I240492,I240543);
not I_13939 (I240565,I240526);
DFFARX1 I_13940 (I586169,I3563,I240500,I240591,);
not I_13941 (I240599,I240591);
and I_13942 (I240616,I240565,I586187);
not I_13943 (I240633,I586184);
nand I_13944 (I240650,I240633,I586187);
not I_13945 (I240667,I586163);
nor I_13946 (I240684,I240667,I586166);
nand I_13947 (I240701,I240684,I586175);
nor I_13948 (I240718,I240701,I240650);
DFFARX1 I_13949 (I240718,I3563,I240500,I240468,);
not I_13950 (I240749,I240701);
not I_13951 (I240766,I586166);
nand I_13952 (I240783,I240766,I586187);
nor I_13953 (I240800,I586166,I586184);
nand I_13954 (I240480,I240616,I240800);
nand I_13955 (I240474,I240565,I586166);
nand I_13956 (I240845,I240667,I586181);
DFFARX1 I_13957 (I240845,I3563,I240500,I240489,);
DFFARX1 I_13958 (I240845,I3563,I240500,I240483,);
not I_13959 (I240890,I586181);
nor I_13960 (I240907,I240890,I586163);
and I_13961 (I240924,I240907,I586172);
or I_13962 (I240941,I240924,I586166);
DFFARX1 I_13963 (I240941,I3563,I240500,I240967,);
nand I_13964 (I240975,I240967,I240633);
nor I_13965 (I240477,I240975,I240783);
nor I_13966 (I240471,I240967,I240599);
DFFARX1 I_13967 (I240967,I3563,I240500,I241029,);
not I_13968 (I241037,I241029);
nor I_13969 (I240486,I241037,I240749);
not I_13970 (I241095,I3570);
DFFARX1 I_13971 (I1240697,I3563,I241095,I241121,);
DFFARX1 I_13972 (I241121,I3563,I241095,I241138,);
not I_13973 (I241087,I241138);
not I_13974 (I241160,I241121);
DFFARX1 I_13975 (I1240697,I3563,I241095,I241186,);
not I_13976 (I241194,I241186);
and I_13977 (I241211,I241160,I1240700);
not I_13978 (I241228,I1240712);
nand I_13979 (I241245,I241228,I1240700);
not I_13980 (I241262,I1240718);
nor I_13981 (I241279,I241262,I1240709);
nand I_13982 (I241296,I241279,I1240715);
nor I_13983 (I241313,I241296,I241245);
DFFARX1 I_13984 (I241313,I3563,I241095,I241063,);
not I_13985 (I241344,I241296);
not I_13986 (I241361,I1240709);
nand I_13987 (I241378,I241361,I1240700);
nor I_13988 (I241395,I1240709,I1240712);
nand I_13989 (I241075,I241211,I241395);
nand I_13990 (I241069,I241160,I1240709);
nand I_13991 (I241440,I241262,I1240706);
DFFARX1 I_13992 (I241440,I3563,I241095,I241084,);
DFFARX1 I_13993 (I241440,I3563,I241095,I241078,);
not I_13994 (I241485,I1240706);
nor I_13995 (I241502,I241485,I1240703);
and I_13996 (I241519,I241502,I1240721);
or I_13997 (I241536,I241519,I1240700);
DFFARX1 I_13998 (I241536,I3563,I241095,I241562,);
nand I_13999 (I241570,I241562,I241228);
nor I_14000 (I241072,I241570,I241378);
nor I_14001 (I241066,I241562,I241194);
DFFARX1 I_14002 (I241562,I3563,I241095,I241624,);
not I_14003 (I241632,I241624);
nor I_14004 (I241081,I241632,I241344);
not I_14005 (I241690,I3570);
DFFARX1 I_14006 (I419750,I3563,I241690,I241716,);
DFFARX1 I_14007 (I241716,I3563,I241690,I241733,);
not I_14008 (I241682,I241733);
not I_14009 (I241755,I241716);
DFFARX1 I_14010 (I419765,I3563,I241690,I241781,);
not I_14011 (I241789,I241781);
and I_14012 (I241806,I241755,I419762);
not I_14013 (I241823,I419750);
nand I_14014 (I241840,I241823,I419762);
not I_14015 (I241857,I419759);
nor I_14016 (I241874,I241857,I419774);
nand I_14017 (I241891,I241874,I419771);
nor I_14018 (I241908,I241891,I241840);
DFFARX1 I_14019 (I241908,I3563,I241690,I241658,);
not I_14020 (I241939,I241891);
not I_14021 (I241956,I419774);
nand I_14022 (I241973,I241956,I419762);
nor I_14023 (I241990,I419774,I419750);
nand I_14024 (I241670,I241806,I241990);
nand I_14025 (I241664,I241755,I419774);
nand I_14026 (I242035,I241857,I419768);
DFFARX1 I_14027 (I242035,I3563,I241690,I241679,);
DFFARX1 I_14028 (I242035,I3563,I241690,I241673,);
not I_14029 (I242080,I419768);
nor I_14030 (I242097,I242080,I419756);
and I_14031 (I242114,I242097,I419777);
or I_14032 (I242131,I242114,I419753);
DFFARX1 I_14033 (I242131,I3563,I241690,I242157,);
nand I_14034 (I242165,I242157,I241823);
nor I_14035 (I241667,I242165,I241973);
nor I_14036 (I241661,I242157,I241789);
DFFARX1 I_14037 (I242157,I3563,I241690,I242219,);
not I_14038 (I242227,I242219);
nor I_14039 (I241676,I242227,I241939);
not I_14040 (I242285,I3570);
DFFARX1 I_14041 (I51928,I3563,I242285,I242311,);
DFFARX1 I_14042 (I242311,I3563,I242285,I242328,);
not I_14043 (I242277,I242328);
not I_14044 (I242350,I242311);
DFFARX1 I_14045 (I51904,I3563,I242285,I242376,);
not I_14046 (I242384,I242376);
and I_14047 (I242401,I242350,I51919);
not I_14048 (I242418,I51907);
nand I_14049 (I242435,I242418,I51919);
not I_14050 (I242452,I51910);
nor I_14051 (I242469,I242452,I51922);
nand I_14052 (I242486,I242469,I51913);
nor I_14053 (I242503,I242486,I242435);
DFFARX1 I_14054 (I242503,I3563,I242285,I242253,);
not I_14055 (I242534,I242486);
not I_14056 (I242551,I51922);
nand I_14057 (I242568,I242551,I51919);
nor I_14058 (I242585,I51922,I51907);
nand I_14059 (I242265,I242401,I242585);
nand I_14060 (I242259,I242350,I51922);
nand I_14061 (I242630,I242452,I51916);
DFFARX1 I_14062 (I242630,I3563,I242285,I242274,);
DFFARX1 I_14063 (I242630,I3563,I242285,I242268,);
not I_14064 (I242675,I51916);
nor I_14065 (I242692,I242675,I51907);
and I_14066 (I242709,I242692,I51904);
or I_14067 (I242726,I242709,I51925);
DFFARX1 I_14068 (I242726,I3563,I242285,I242752,);
nand I_14069 (I242760,I242752,I242418);
nor I_14070 (I242262,I242760,I242568);
nor I_14071 (I242256,I242752,I242384);
DFFARX1 I_14072 (I242752,I3563,I242285,I242814,);
not I_14073 (I242822,I242814);
nor I_14074 (I242271,I242822,I242534);
not I_14075 (I242880,I3570);
DFFARX1 I_14076 (I144138,I3563,I242880,I242906,);
DFFARX1 I_14077 (I242906,I3563,I242880,I242923,);
not I_14078 (I242872,I242923);
not I_14079 (I242945,I242906);
DFFARX1 I_14080 (I144132,I3563,I242880,I242971,);
not I_14081 (I242979,I242971);
and I_14082 (I242996,I242945,I144129);
not I_14083 (I243013,I144150);
nand I_14084 (I243030,I243013,I144129);
not I_14085 (I243047,I144144);
nor I_14086 (I243064,I243047,I144135);
nand I_14087 (I243081,I243064,I144141);
nor I_14088 (I243098,I243081,I243030);
DFFARX1 I_14089 (I243098,I3563,I242880,I242848,);
not I_14090 (I243129,I243081);
not I_14091 (I243146,I144135);
nand I_14092 (I243163,I243146,I144129);
nor I_14093 (I243180,I144135,I144150);
nand I_14094 (I242860,I242996,I243180);
nand I_14095 (I242854,I242945,I144135);
nand I_14096 (I243225,I243047,I144129);
DFFARX1 I_14097 (I243225,I3563,I242880,I242869,);
DFFARX1 I_14098 (I243225,I3563,I242880,I242863,);
not I_14099 (I243270,I144129);
nor I_14100 (I243287,I243270,I144147);
and I_14101 (I243304,I243287,I144153);
or I_14102 (I243321,I243304,I144132);
DFFARX1 I_14103 (I243321,I3563,I242880,I243347,);
nand I_14104 (I243355,I243347,I243013);
nor I_14105 (I242857,I243355,I243163);
nor I_14106 (I242851,I243347,I242979);
DFFARX1 I_14107 (I243347,I3563,I242880,I243409,);
not I_14108 (I243417,I243409);
nor I_14109 (I242866,I243417,I243129);
not I_14110 (I243475,I3570);
DFFARX1 I_14111 (I872194,I3563,I243475,I243501,);
DFFARX1 I_14112 (I243501,I3563,I243475,I243518,);
not I_14113 (I243467,I243518);
not I_14114 (I243540,I243501);
DFFARX1 I_14115 (I872188,I3563,I243475,I243566,);
not I_14116 (I243574,I243566);
and I_14117 (I243591,I243540,I872206);
not I_14118 (I243608,I872194);
nand I_14119 (I243625,I243608,I872206);
not I_14120 (I243642,I872188);
nor I_14121 (I243659,I243642,I872200);
nand I_14122 (I243676,I243659,I872191);
nor I_14123 (I243693,I243676,I243625);
DFFARX1 I_14124 (I243693,I3563,I243475,I243443,);
not I_14125 (I243724,I243676);
not I_14126 (I243741,I872200);
nand I_14127 (I243758,I243741,I872206);
nor I_14128 (I243775,I872200,I872194);
nand I_14129 (I243455,I243591,I243775);
nand I_14130 (I243449,I243540,I872200);
nand I_14131 (I243820,I243642,I872203);
DFFARX1 I_14132 (I243820,I3563,I243475,I243464,);
DFFARX1 I_14133 (I243820,I3563,I243475,I243458,);
not I_14134 (I243865,I872203);
nor I_14135 (I243882,I243865,I872209);
and I_14136 (I243899,I243882,I872191);
or I_14137 (I243916,I243899,I872197);
DFFARX1 I_14138 (I243916,I3563,I243475,I243942,);
nand I_14139 (I243950,I243942,I243608);
nor I_14140 (I243452,I243950,I243758);
nor I_14141 (I243446,I243942,I243574);
DFFARX1 I_14142 (I243942,I3563,I243475,I244004,);
not I_14143 (I244012,I244004);
nor I_14144 (I243461,I244012,I243724);
not I_14145 (I244070,I3570);
DFFARX1 I_14146 (I1061809,I3563,I244070,I244096,);
DFFARX1 I_14147 (I244096,I3563,I244070,I244113,);
not I_14148 (I244062,I244113);
not I_14149 (I244135,I244096);
DFFARX1 I_14150 (I1061818,I3563,I244070,I244161,);
not I_14151 (I244169,I244161);
and I_14152 (I244186,I244135,I1061812);
not I_14153 (I244203,I1061806);
nand I_14154 (I244220,I244203,I1061812);
not I_14155 (I244237,I1061821);
nor I_14156 (I244254,I244237,I1061809);
nand I_14157 (I244271,I244254,I1061815);
nor I_14158 (I244288,I244271,I244220);
DFFARX1 I_14159 (I244288,I3563,I244070,I244038,);
not I_14160 (I244319,I244271);
not I_14161 (I244336,I1061809);
nand I_14162 (I244353,I244336,I1061812);
nor I_14163 (I244370,I1061809,I1061806);
nand I_14164 (I244050,I244186,I244370);
nand I_14165 (I244044,I244135,I1061809);
nand I_14166 (I244415,I244237,I1061812);
DFFARX1 I_14167 (I244415,I3563,I244070,I244059,);
DFFARX1 I_14168 (I244415,I3563,I244070,I244053,);
not I_14169 (I244460,I1061812);
nor I_14170 (I244477,I244460,I1061827);
and I_14171 (I244494,I244477,I1061824);
or I_14172 (I244511,I244494,I1061806);
DFFARX1 I_14173 (I244511,I3563,I244070,I244537,);
nand I_14174 (I244545,I244537,I244203);
nor I_14175 (I244047,I244545,I244353);
nor I_14176 (I244041,I244537,I244169);
DFFARX1 I_14177 (I244537,I3563,I244070,I244599,);
not I_14178 (I244607,I244599);
nor I_14179 (I244056,I244607,I244319);
not I_14180 (I244665,I3570);
DFFARX1 I_14181 (I1316656,I3563,I244665,I244691,);
DFFARX1 I_14182 (I244691,I3563,I244665,I244708,);
not I_14183 (I244657,I244708);
not I_14184 (I244730,I244691);
DFFARX1 I_14185 (I1316668,I3563,I244665,I244756,);
not I_14186 (I244764,I244756);
and I_14187 (I244781,I244730,I1316662);
not I_14188 (I244798,I1316674);
nand I_14189 (I244815,I244798,I1316662);
not I_14190 (I244832,I1316659);
nor I_14191 (I244849,I244832,I1316671);
nand I_14192 (I244866,I244849,I1316653);
nor I_14193 (I244883,I244866,I244815);
DFFARX1 I_14194 (I244883,I3563,I244665,I244633,);
not I_14195 (I244914,I244866);
not I_14196 (I244931,I1316671);
nand I_14197 (I244948,I244931,I1316662);
nor I_14198 (I244965,I1316671,I1316674);
nand I_14199 (I244645,I244781,I244965);
nand I_14200 (I244639,I244730,I1316671);
nand I_14201 (I245010,I244832,I1316665);
DFFARX1 I_14202 (I245010,I3563,I244665,I244654,);
DFFARX1 I_14203 (I245010,I3563,I244665,I244648,);
not I_14204 (I245055,I1316665);
nor I_14205 (I245072,I245055,I1316656);
and I_14206 (I245089,I245072,I1316653);
or I_14207 (I245106,I245089,I1316677);
DFFARX1 I_14208 (I245106,I3563,I244665,I245132,);
nand I_14209 (I245140,I245132,I244798);
nor I_14210 (I244642,I245140,I244948);
nor I_14211 (I244636,I245132,I244764);
DFFARX1 I_14212 (I245132,I3563,I244665,I245194,);
not I_14213 (I245202,I245194);
nor I_14214 (I244651,I245202,I244914);
not I_14215 (I245260,I3570);
DFFARX1 I_14216 (I25578,I3563,I245260,I245286,);
DFFARX1 I_14217 (I245286,I3563,I245260,I245303,);
not I_14218 (I245252,I245303);
not I_14219 (I245325,I245286);
DFFARX1 I_14220 (I25554,I3563,I245260,I245351,);
not I_14221 (I245359,I245351);
and I_14222 (I245376,I245325,I25569);
not I_14223 (I245393,I25557);
nand I_14224 (I245410,I245393,I25569);
not I_14225 (I245427,I25560);
nor I_14226 (I245444,I245427,I25572);
nand I_14227 (I245461,I245444,I25563);
nor I_14228 (I245478,I245461,I245410);
DFFARX1 I_14229 (I245478,I3563,I245260,I245228,);
not I_14230 (I245509,I245461);
not I_14231 (I245526,I25572);
nand I_14232 (I245543,I245526,I25569);
nor I_14233 (I245560,I25572,I25557);
nand I_14234 (I245240,I245376,I245560);
nand I_14235 (I245234,I245325,I25572);
nand I_14236 (I245605,I245427,I25566);
DFFARX1 I_14237 (I245605,I3563,I245260,I245249,);
DFFARX1 I_14238 (I245605,I3563,I245260,I245243,);
not I_14239 (I245650,I25566);
nor I_14240 (I245667,I245650,I25557);
and I_14241 (I245684,I245667,I25554);
or I_14242 (I245701,I245684,I25575);
DFFARX1 I_14243 (I245701,I3563,I245260,I245727,);
nand I_14244 (I245735,I245727,I245393);
nor I_14245 (I245237,I245735,I245543);
nor I_14246 (I245231,I245727,I245359);
DFFARX1 I_14247 (I245727,I3563,I245260,I245789,);
not I_14248 (I245797,I245789);
nor I_14249 (I245246,I245797,I245509);
not I_14250 (I245855,I3570);
DFFARX1 I_14251 (I294324,I3563,I245855,I245881,);
DFFARX1 I_14252 (I245881,I3563,I245855,I245898,);
not I_14253 (I245847,I245898);
not I_14254 (I245920,I245881);
DFFARX1 I_14255 (I294339,I3563,I245855,I245946,);
not I_14256 (I245954,I245946);
and I_14257 (I245971,I245920,I294336);
not I_14258 (I245988,I294324);
nand I_14259 (I246005,I245988,I294336);
not I_14260 (I246022,I294333);
nor I_14261 (I246039,I246022,I294348);
nand I_14262 (I246056,I246039,I294345);
nor I_14263 (I246073,I246056,I246005);
DFFARX1 I_14264 (I246073,I3563,I245855,I245823,);
not I_14265 (I246104,I246056);
not I_14266 (I246121,I294348);
nand I_14267 (I246138,I246121,I294336);
nor I_14268 (I246155,I294348,I294324);
nand I_14269 (I245835,I245971,I246155);
nand I_14270 (I245829,I245920,I294348);
nand I_14271 (I246200,I246022,I294342);
DFFARX1 I_14272 (I246200,I3563,I245855,I245844,);
DFFARX1 I_14273 (I246200,I3563,I245855,I245838,);
not I_14274 (I246245,I294342);
nor I_14275 (I246262,I246245,I294330);
and I_14276 (I246279,I246262,I294351);
or I_14277 (I246296,I246279,I294327);
DFFARX1 I_14278 (I246296,I3563,I245855,I246322,);
nand I_14279 (I246330,I246322,I245988);
nor I_14280 (I245832,I246330,I246138);
nor I_14281 (I245826,I246322,I245954);
DFFARX1 I_14282 (I246322,I3563,I245855,I246384,);
not I_14283 (I246392,I246384);
nor I_14284 (I245841,I246392,I246104);
not I_14285 (I246450,I3570);
DFFARX1 I_14286 (I482810,I3563,I246450,I246476,);
DFFARX1 I_14287 (I246476,I3563,I246450,I246493,);
not I_14288 (I246442,I246493);
not I_14289 (I246515,I246476);
DFFARX1 I_14290 (I482798,I3563,I246450,I246541,);
not I_14291 (I246549,I246541);
and I_14292 (I246566,I246515,I482807);
not I_14293 (I246583,I482804);
nand I_14294 (I246600,I246583,I482807);
not I_14295 (I246617,I482795);
nor I_14296 (I246634,I246617,I482801);
nand I_14297 (I246651,I246634,I482786);
nor I_14298 (I246668,I246651,I246600);
DFFARX1 I_14299 (I246668,I3563,I246450,I246418,);
not I_14300 (I246699,I246651);
not I_14301 (I246716,I482801);
nand I_14302 (I246733,I246716,I482807);
nor I_14303 (I246750,I482801,I482804);
nand I_14304 (I246430,I246566,I246750);
nand I_14305 (I246424,I246515,I482801);
nand I_14306 (I246795,I246617,I482786);
DFFARX1 I_14307 (I246795,I3563,I246450,I246439,);
DFFARX1 I_14308 (I246795,I3563,I246450,I246433,);
not I_14309 (I246840,I482786);
nor I_14310 (I246857,I246840,I482792);
and I_14311 (I246874,I246857,I482789);
or I_14312 (I246891,I246874,I482813);
DFFARX1 I_14313 (I246891,I3563,I246450,I246917,);
nand I_14314 (I246925,I246917,I246583);
nor I_14315 (I246427,I246925,I246733);
nor I_14316 (I246421,I246917,I246549);
DFFARX1 I_14317 (I246917,I3563,I246450,I246979,);
not I_14318 (I246987,I246979);
nor I_14319 (I246436,I246987,I246699);
not I_14320 (I247045,I3570);
DFFARX1 I_14321 (I965924,I3563,I247045,I247071,);
DFFARX1 I_14322 (I247071,I3563,I247045,I247088,);
not I_14323 (I247037,I247088);
not I_14324 (I247110,I247071);
DFFARX1 I_14325 (I965933,I3563,I247045,I247136,);
not I_14326 (I247144,I247136);
and I_14327 (I247161,I247110,I965921);
not I_14328 (I247178,I965912);
nand I_14329 (I247195,I247178,I965921);
not I_14330 (I247212,I965918);
nor I_14331 (I247229,I247212,I965936);
nand I_14332 (I247246,I247229,I965909);
nor I_14333 (I247263,I247246,I247195);
DFFARX1 I_14334 (I247263,I3563,I247045,I247013,);
not I_14335 (I247294,I247246);
not I_14336 (I247311,I965936);
nand I_14337 (I247328,I247311,I965921);
nor I_14338 (I247345,I965936,I965912);
nand I_14339 (I247025,I247161,I247345);
nand I_14340 (I247019,I247110,I965936);
nand I_14341 (I247390,I247212,I965915);
DFFARX1 I_14342 (I247390,I3563,I247045,I247034,);
DFFARX1 I_14343 (I247390,I3563,I247045,I247028,);
not I_14344 (I247435,I965915);
nor I_14345 (I247452,I247435,I965927);
and I_14346 (I247469,I247452,I965909);
or I_14347 (I247486,I247469,I965930);
DFFARX1 I_14348 (I247486,I3563,I247045,I247512,);
nand I_14349 (I247520,I247512,I247178);
nor I_14350 (I247022,I247520,I247328);
nor I_14351 (I247016,I247512,I247144);
DFFARX1 I_14352 (I247512,I3563,I247045,I247574,);
not I_14353 (I247582,I247574);
nor I_14354 (I247031,I247582,I247294);
not I_14355 (I247640,I3570);
DFFARX1 I_14356 (I1166135,I3563,I247640,I247666,);
DFFARX1 I_14357 (I247666,I3563,I247640,I247683,);
not I_14358 (I247632,I247683);
not I_14359 (I247705,I247666);
DFFARX1 I_14360 (I1166135,I3563,I247640,I247731,);
not I_14361 (I247739,I247731);
and I_14362 (I247756,I247705,I1166138);
not I_14363 (I247773,I1166150);
nand I_14364 (I247790,I247773,I1166138);
not I_14365 (I247807,I1166156);
nor I_14366 (I247824,I247807,I1166147);
nand I_14367 (I247841,I247824,I1166153);
nor I_14368 (I247858,I247841,I247790);
DFFARX1 I_14369 (I247858,I3563,I247640,I247608,);
not I_14370 (I247889,I247841);
not I_14371 (I247906,I1166147);
nand I_14372 (I247923,I247906,I1166138);
nor I_14373 (I247940,I1166147,I1166150);
nand I_14374 (I247620,I247756,I247940);
nand I_14375 (I247614,I247705,I1166147);
nand I_14376 (I247985,I247807,I1166144);
DFFARX1 I_14377 (I247985,I3563,I247640,I247629,);
DFFARX1 I_14378 (I247985,I3563,I247640,I247623,);
not I_14379 (I248030,I1166144);
nor I_14380 (I248047,I248030,I1166141);
and I_14381 (I248064,I248047,I1166159);
or I_14382 (I248081,I248064,I1166138);
DFFARX1 I_14383 (I248081,I3563,I247640,I248107,);
nand I_14384 (I248115,I248107,I247773);
nor I_14385 (I247617,I248115,I247923);
nor I_14386 (I247611,I248107,I247739);
DFFARX1 I_14387 (I248107,I3563,I247640,I248169,);
not I_14388 (I248177,I248169);
nor I_14389 (I247626,I248177,I247889);
not I_14390 (I248235,I3570);
DFFARX1 I_14391 (I1181163,I3563,I248235,I248261,);
DFFARX1 I_14392 (I248261,I3563,I248235,I248278,);
not I_14393 (I248227,I248278);
not I_14394 (I248300,I248261);
DFFARX1 I_14395 (I1181163,I3563,I248235,I248326,);
not I_14396 (I248334,I248326);
and I_14397 (I248351,I248300,I1181166);
not I_14398 (I248368,I1181178);
nand I_14399 (I248385,I248368,I1181166);
not I_14400 (I248402,I1181184);
nor I_14401 (I248419,I248402,I1181175);
nand I_14402 (I248436,I248419,I1181181);
nor I_14403 (I248453,I248436,I248385);
DFFARX1 I_14404 (I248453,I3563,I248235,I248203,);
not I_14405 (I248484,I248436);
not I_14406 (I248501,I1181175);
nand I_14407 (I248518,I248501,I1181166);
nor I_14408 (I248535,I1181175,I1181178);
nand I_14409 (I248215,I248351,I248535);
nand I_14410 (I248209,I248300,I1181175);
nand I_14411 (I248580,I248402,I1181172);
DFFARX1 I_14412 (I248580,I3563,I248235,I248224,);
DFFARX1 I_14413 (I248580,I3563,I248235,I248218,);
not I_14414 (I248625,I1181172);
nor I_14415 (I248642,I248625,I1181169);
and I_14416 (I248659,I248642,I1181187);
or I_14417 (I248676,I248659,I1181166);
DFFARX1 I_14418 (I248676,I3563,I248235,I248702,);
nand I_14419 (I248710,I248702,I248368);
nor I_14420 (I248212,I248710,I248518);
nor I_14421 (I248206,I248702,I248334);
DFFARX1 I_14422 (I248702,I3563,I248235,I248764,);
not I_14423 (I248772,I248764);
nor I_14424 (I248221,I248772,I248484);
not I_14425 (I248830,I3570);
DFFARX1 I_14426 (I1365464,I3563,I248830,I248856,);
DFFARX1 I_14427 (I248856,I3563,I248830,I248873,);
not I_14428 (I248822,I248873);
not I_14429 (I248895,I248856);
DFFARX1 I_14430 (I1365455,I3563,I248830,I248921,);
not I_14431 (I248929,I248921);
and I_14432 (I248946,I248895,I1365449);
not I_14433 (I248963,I1365443);
nand I_14434 (I248980,I248963,I1365449);
not I_14435 (I248997,I1365470);
nor I_14436 (I249014,I248997,I1365443);
nand I_14437 (I249031,I249014,I1365467);
nor I_14438 (I249048,I249031,I248980);
DFFARX1 I_14439 (I249048,I3563,I248830,I248798,);
not I_14440 (I249079,I249031);
not I_14441 (I249096,I1365443);
nand I_14442 (I249113,I249096,I1365449);
nor I_14443 (I249130,I1365443,I1365443);
nand I_14444 (I248810,I248946,I249130);
nand I_14445 (I248804,I248895,I1365443);
nand I_14446 (I249175,I248997,I1365452);
DFFARX1 I_14447 (I249175,I3563,I248830,I248819,);
DFFARX1 I_14448 (I249175,I3563,I248830,I248813,);
not I_14449 (I249220,I1365452);
nor I_14450 (I249237,I249220,I1365458);
and I_14451 (I249254,I249237,I1365461);
or I_14452 (I249271,I249254,I1365446);
DFFARX1 I_14453 (I249271,I3563,I248830,I249297,);
nand I_14454 (I249305,I249297,I248963);
nor I_14455 (I248807,I249305,I249113);
nor I_14456 (I248801,I249297,I248929);
DFFARX1 I_14457 (I249297,I3563,I248830,I249359,);
not I_14458 (I249367,I249359);
nor I_14459 (I248816,I249367,I249079);
not I_14460 (I249425,I3570);
DFFARX1 I_14461 (I389711,I3563,I249425,I249451,);
DFFARX1 I_14462 (I249451,I3563,I249425,I249468,);
not I_14463 (I249417,I249468);
not I_14464 (I249490,I249451);
DFFARX1 I_14465 (I389726,I3563,I249425,I249516,);
not I_14466 (I249524,I249516);
and I_14467 (I249541,I249490,I389723);
not I_14468 (I249558,I389711);
nand I_14469 (I249575,I249558,I389723);
not I_14470 (I249592,I389720);
nor I_14471 (I249609,I249592,I389735);
nand I_14472 (I249626,I249609,I389732);
nor I_14473 (I249643,I249626,I249575);
DFFARX1 I_14474 (I249643,I3563,I249425,I249393,);
not I_14475 (I249674,I249626);
not I_14476 (I249691,I389735);
nand I_14477 (I249708,I249691,I389723);
nor I_14478 (I249725,I389735,I389711);
nand I_14479 (I249405,I249541,I249725);
nand I_14480 (I249399,I249490,I389735);
nand I_14481 (I249770,I249592,I389729);
DFFARX1 I_14482 (I249770,I3563,I249425,I249414,);
DFFARX1 I_14483 (I249770,I3563,I249425,I249408,);
not I_14484 (I249815,I389729);
nor I_14485 (I249832,I249815,I389717);
and I_14486 (I249849,I249832,I389738);
or I_14487 (I249866,I249849,I389714);
DFFARX1 I_14488 (I249866,I3563,I249425,I249892,);
nand I_14489 (I249900,I249892,I249558);
nor I_14490 (I249402,I249900,I249708);
nor I_14491 (I249396,I249892,I249524);
DFFARX1 I_14492 (I249892,I3563,I249425,I249954,);
not I_14493 (I249962,I249954);
nor I_14494 (I249411,I249962,I249674);
not I_14495 (I250020,I3570);
DFFARX1 I_14496 (I718537,I3563,I250020,I250046,);
DFFARX1 I_14497 (I250046,I3563,I250020,I250063,);
not I_14498 (I250012,I250063);
not I_14499 (I250085,I250046);
DFFARX1 I_14500 (I718534,I3563,I250020,I250111,);
not I_14501 (I250119,I250111);
and I_14502 (I250136,I250085,I718540);
not I_14503 (I250153,I718525);
nand I_14504 (I250170,I250153,I718540);
not I_14505 (I250187,I718528);
nor I_14506 (I250204,I250187,I718549);
nand I_14507 (I250221,I250204,I718546);
nor I_14508 (I250238,I250221,I250170);
DFFARX1 I_14509 (I250238,I3563,I250020,I249988,);
not I_14510 (I250269,I250221);
not I_14511 (I250286,I718549);
nand I_14512 (I250303,I250286,I718540);
nor I_14513 (I250320,I718549,I718525);
nand I_14514 (I250000,I250136,I250320);
nand I_14515 (I249994,I250085,I718549);
nand I_14516 (I250365,I250187,I718525);
DFFARX1 I_14517 (I250365,I3563,I250020,I250009,);
DFFARX1 I_14518 (I250365,I3563,I250020,I250003,);
not I_14519 (I250410,I718525);
nor I_14520 (I250427,I250410,I718531);
and I_14521 (I250444,I250427,I718543);
or I_14522 (I250461,I250444,I718528);
DFFARX1 I_14523 (I250461,I3563,I250020,I250487,);
nand I_14524 (I250495,I250487,I250153);
nor I_14525 (I249997,I250495,I250303);
nor I_14526 (I249991,I250487,I250119);
DFFARX1 I_14527 (I250487,I3563,I250020,I250549,);
not I_14528 (I250557,I250549);
nor I_14529 (I250006,I250557,I250269);
not I_14530 (I250615,I3570);
DFFARX1 I_14531 (I1066297,I3563,I250615,I250641,);
DFFARX1 I_14532 (I250641,I3563,I250615,I250658,);
not I_14533 (I250607,I250658);
not I_14534 (I250680,I250641);
DFFARX1 I_14535 (I1066306,I3563,I250615,I250706,);
not I_14536 (I250714,I250706);
and I_14537 (I250731,I250680,I1066300);
not I_14538 (I250748,I1066294);
nand I_14539 (I250765,I250748,I1066300);
not I_14540 (I250782,I1066309);
nor I_14541 (I250799,I250782,I1066297);
nand I_14542 (I250816,I250799,I1066303);
nor I_14543 (I250833,I250816,I250765);
DFFARX1 I_14544 (I250833,I3563,I250615,I250583,);
not I_14545 (I250864,I250816);
not I_14546 (I250881,I1066297);
nand I_14547 (I250898,I250881,I1066300);
nor I_14548 (I250915,I1066297,I1066294);
nand I_14549 (I250595,I250731,I250915);
nand I_14550 (I250589,I250680,I1066297);
nand I_14551 (I250960,I250782,I1066300);
DFFARX1 I_14552 (I250960,I3563,I250615,I250604,);
DFFARX1 I_14553 (I250960,I3563,I250615,I250598,);
not I_14554 (I251005,I1066300);
nor I_14555 (I251022,I251005,I1066315);
and I_14556 (I251039,I251022,I1066312);
or I_14557 (I251056,I251039,I1066294);
DFFARX1 I_14558 (I251056,I3563,I250615,I251082,);
nand I_14559 (I251090,I251082,I250748);
nor I_14560 (I250592,I251090,I250898);
nor I_14561 (I250586,I251082,I250714);
DFFARX1 I_14562 (I251082,I3563,I250615,I251144,);
not I_14563 (I251152,I251144);
nor I_14564 (I250601,I251152,I250864);
not I_14565 (I251210,I3570);
DFFARX1 I_14566 (I1392239,I3563,I251210,I251236,);
DFFARX1 I_14567 (I251236,I3563,I251210,I251253,);
not I_14568 (I251202,I251253);
not I_14569 (I251275,I251236);
DFFARX1 I_14570 (I1392230,I3563,I251210,I251301,);
not I_14571 (I251309,I251301);
and I_14572 (I251326,I251275,I1392224);
not I_14573 (I251343,I1392218);
nand I_14574 (I251360,I251343,I1392224);
not I_14575 (I251377,I1392245);
nor I_14576 (I251394,I251377,I1392218);
nand I_14577 (I251411,I251394,I1392242);
nor I_14578 (I251428,I251411,I251360);
DFFARX1 I_14579 (I251428,I3563,I251210,I251178,);
not I_14580 (I251459,I251411);
not I_14581 (I251476,I1392218);
nand I_14582 (I251493,I251476,I1392224);
nor I_14583 (I251510,I1392218,I1392218);
nand I_14584 (I251190,I251326,I251510);
nand I_14585 (I251184,I251275,I1392218);
nand I_14586 (I251555,I251377,I1392227);
DFFARX1 I_14587 (I251555,I3563,I251210,I251199,);
DFFARX1 I_14588 (I251555,I3563,I251210,I251193,);
not I_14589 (I251600,I1392227);
nor I_14590 (I251617,I251600,I1392233);
and I_14591 (I251634,I251617,I1392236);
or I_14592 (I251651,I251634,I1392221);
DFFARX1 I_14593 (I251651,I3563,I251210,I251677,);
nand I_14594 (I251685,I251677,I251343);
nor I_14595 (I251187,I251685,I251493);
nor I_14596 (I251181,I251677,I251309);
DFFARX1 I_14597 (I251677,I3563,I251210,I251739,);
not I_14598 (I251747,I251739);
nor I_14599 (I251196,I251747,I251459);
not I_14600 (I251805,I3570);
DFFARX1 I_14601 (I536433,I3563,I251805,I251831,);
DFFARX1 I_14602 (I251831,I3563,I251805,I251848,);
not I_14603 (I251797,I251848);
not I_14604 (I251870,I251831);
DFFARX1 I_14605 (I536427,I3563,I251805,I251896,);
not I_14606 (I251904,I251896);
and I_14607 (I251921,I251870,I536442);
not I_14608 (I251938,I536439);
nand I_14609 (I251955,I251938,I536442);
not I_14610 (I251972,I536430);
nor I_14611 (I251989,I251972,I536421);
nand I_14612 (I252006,I251989,I536424);
nor I_14613 (I252023,I252006,I251955);
DFFARX1 I_14614 (I252023,I3563,I251805,I251773,);
not I_14615 (I252054,I252006);
not I_14616 (I252071,I536421);
nand I_14617 (I252088,I252071,I536442);
nor I_14618 (I252105,I536421,I536439);
nand I_14619 (I251785,I251921,I252105);
nand I_14620 (I251779,I251870,I536421);
nand I_14621 (I252150,I251972,I536445);
DFFARX1 I_14622 (I252150,I3563,I251805,I251794,);
DFFARX1 I_14623 (I252150,I3563,I251805,I251788,);
not I_14624 (I252195,I536445);
nor I_14625 (I252212,I252195,I536436);
and I_14626 (I252229,I252212,I536421);
or I_14627 (I252246,I252229,I536424);
DFFARX1 I_14628 (I252246,I3563,I251805,I252272,);
nand I_14629 (I252280,I252272,I251938);
nor I_14630 (I251782,I252280,I252088);
nor I_14631 (I251776,I252272,I251904);
DFFARX1 I_14632 (I252272,I3563,I251805,I252334,);
not I_14633 (I252342,I252334);
nor I_14634 (I251791,I252342,I252054);
not I_14635 (I252400,I3570);
DFFARX1 I_14636 (I490426,I3563,I252400,I252426,);
DFFARX1 I_14637 (I252426,I3563,I252400,I252443,);
not I_14638 (I252392,I252443);
not I_14639 (I252465,I252426);
DFFARX1 I_14640 (I490414,I3563,I252400,I252491,);
not I_14641 (I252499,I252491);
and I_14642 (I252516,I252465,I490423);
not I_14643 (I252533,I490420);
nand I_14644 (I252550,I252533,I490423);
not I_14645 (I252567,I490411);
nor I_14646 (I252584,I252567,I490417);
nand I_14647 (I252601,I252584,I490402);
nor I_14648 (I252618,I252601,I252550);
DFFARX1 I_14649 (I252618,I3563,I252400,I252368,);
not I_14650 (I252649,I252601);
not I_14651 (I252666,I490417);
nand I_14652 (I252683,I252666,I490423);
nor I_14653 (I252700,I490417,I490420);
nand I_14654 (I252380,I252516,I252700);
nand I_14655 (I252374,I252465,I490417);
nand I_14656 (I252745,I252567,I490402);
DFFARX1 I_14657 (I252745,I3563,I252400,I252389,);
DFFARX1 I_14658 (I252745,I3563,I252400,I252383,);
not I_14659 (I252790,I490402);
nor I_14660 (I252807,I252790,I490408);
and I_14661 (I252824,I252807,I490405);
or I_14662 (I252841,I252824,I490429);
DFFARX1 I_14663 (I252841,I3563,I252400,I252867,);
nand I_14664 (I252875,I252867,I252533);
nor I_14665 (I252377,I252875,I252683);
nor I_14666 (I252371,I252867,I252499);
DFFARX1 I_14667 (I252867,I3563,I252400,I252929,);
not I_14668 (I252937,I252929);
nor I_14669 (I252386,I252937,I252649);
not I_14670 (I252995,I3570);
DFFARX1 I_14671 (I632996,I3563,I252995,I253021,);
DFFARX1 I_14672 (I253021,I3563,I252995,I253038,);
not I_14673 (I252987,I253038);
not I_14674 (I253060,I253021);
DFFARX1 I_14675 (I632987,I3563,I252995,I253086,);
not I_14676 (I253094,I253086);
and I_14677 (I253111,I253060,I633005);
not I_14678 (I253128,I633002);
nand I_14679 (I253145,I253128,I633005);
not I_14680 (I253162,I632981);
nor I_14681 (I253179,I253162,I632984);
nand I_14682 (I253196,I253179,I632993);
nor I_14683 (I253213,I253196,I253145);
DFFARX1 I_14684 (I253213,I3563,I252995,I252963,);
not I_14685 (I253244,I253196);
not I_14686 (I253261,I632984);
nand I_14687 (I253278,I253261,I633005);
nor I_14688 (I253295,I632984,I633002);
nand I_14689 (I252975,I253111,I253295);
nand I_14690 (I252969,I253060,I632984);
nand I_14691 (I253340,I253162,I632999);
DFFARX1 I_14692 (I253340,I3563,I252995,I252984,);
DFFARX1 I_14693 (I253340,I3563,I252995,I252978,);
not I_14694 (I253385,I632999);
nor I_14695 (I253402,I253385,I632981);
and I_14696 (I253419,I253402,I632990);
or I_14697 (I253436,I253419,I632984);
DFFARX1 I_14698 (I253436,I3563,I252995,I253462,);
nand I_14699 (I253470,I253462,I253128);
nor I_14700 (I252972,I253470,I253278);
nor I_14701 (I252966,I253462,I253094);
DFFARX1 I_14702 (I253462,I3563,I252995,I253524,);
not I_14703 (I253532,I253524);
nor I_14704 (I252981,I253532,I253244);
not I_14705 (I253590,I3570);
DFFARX1 I_14706 (I59291,I3563,I253590,I253616,);
DFFARX1 I_14707 (I253616,I3563,I253590,I253633,);
not I_14708 (I253582,I253633);
not I_14709 (I253655,I253616);
DFFARX1 I_14710 (I59285,I3563,I253590,I253681,);
not I_14711 (I253689,I253681);
and I_14712 (I253706,I253655,I59282);
not I_14713 (I253723,I59303);
nand I_14714 (I253740,I253723,I59282);
not I_14715 (I253757,I59297);
nor I_14716 (I253774,I253757,I59288);
nand I_14717 (I253791,I253774,I59294);
nor I_14718 (I253808,I253791,I253740);
DFFARX1 I_14719 (I253808,I3563,I253590,I253558,);
not I_14720 (I253839,I253791);
not I_14721 (I253856,I59288);
nand I_14722 (I253873,I253856,I59282);
nor I_14723 (I253890,I59288,I59303);
nand I_14724 (I253570,I253706,I253890);
nand I_14725 (I253564,I253655,I59288);
nand I_14726 (I253935,I253757,I59282);
DFFARX1 I_14727 (I253935,I3563,I253590,I253579,);
DFFARX1 I_14728 (I253935,I3563,I253590,I253573,);
not I_14729 (I253980,I59282);
nor I_14730 (I253997,I253980,I59300);
and I_14731 (I254014,I253997,I59306);
or I_14732 (I254031,I254014,I59285);
DFFARX1 I_14733 (I254031,I3563,I253590,I254057,);
nand I_14734 (I254065,I254057,I253723);
nor I_14735 (I253567,I254065,I253873);
nor I_14736 (I253561,I254057,I253689);
DFFARX1 I_14737 (I254057,I3563,I253590,I254119,);
not I_14738 (I254127,I254119);
nor I_14739 (I253576,I254127,I253839);
not I_14740 (I254185,I3570);
DFFARX1 I_14741 (I1191567,I3563,I254185,I254211,);
DFFARX1 I_14742 (I254211,I3563,I254185,I254228,);
not I_14743 (I254177,I254228);
not I_14744 (I254250,I254211);
DFFARX1 I_14745 (I1191567,I3563,I254185,I254276,);
not I_14746 (I254284,I254276);
and I_14747 (I254301,I254250,I1191570);
not I_14748 (I254318,I1191582);
nand I_14749 (I254335,I254318,I1191570);
not I_14750 (I254352,I1191588);
nor I_14751 (I254369,I254352,I1191579);
nand I_14752 (I254386,I254369,I1191585);
nor I_14753 (I254403,I254386,I254335);
DFFARX1 I_14754 (I254403,I3563,I254185,I254153,);
not I_14755 (I254434,I254386);
not I_14756 (I254451,I1191579);
nand I_14757 (I254468,I254451,I1191570);
nor I_14758 (I254485,I1191579,I1191582);
nand I_14759 (I254165,I254301,I254485);
nand I_14760 (I254159,I254250,I1191579);
nand I_14761 (I254530,I254352,I1191576);
DFFARX1 I_14762 (I254530,I3563,I254185,I254174,);
DFFARX1 I_14763 (I254530,I3563,I254185,I254168,);
not I_14764 (I254575,I1191576);
nor I_14765 (I254592,I254575,I1191573);
and I_14766 (I254609,I254592,I1191591);
or I_14767 (I254626,I254609,I1191570);
DFFARX1 I_14768 (I254626,I3563,I254185,I254652,);
nand I_14769 (I254660,I254652,I254318);
nor I_14770 (I254162,I254660,I254468);
nor I_14771 (I254156,I254652,I254284);
DFFARX1 I_14772 (I254652,I3563,I254185,I254714,);
not I_14773 (I254722,I254714);
nor I_14774 (I254171,I254722,I254434);
not I_14775 (I254780,I3570);
DFFARX1 I_14776 (I1118161,I3563,I254780,I254806,);
DFFARX1 I_14777 (I254806,I3563,I254780,I254823,);
not I_14778 (I254772,I254823);
not I_14779 (I254845,I254806);
DFFARX1 I_14780 (I1118161,I3563,I254780,I254871,);
not I_14781 (I254879,I254871);
and I_14782 (I254896,I254845,I1118164);
not I_14783 (I254913,I1118176);
nand I_14784 (I254930,I254913,I1118164);
not I_14785 (I254947,I1118182);
nor I_14786 (I254964,I254947,I1118173);
nand I_14787 (I254981,I254964,I1118179);
nor I_14788 (I254998,I254981,I254930);
DFFARX1 I_14789 (I254998,I3563,I254780,I254748,);
not I_14790 (I255029,I254981);
not I_14791 (I255046,I1118173);
nand I_14792 (I255063,I255046,I1118164);
nor I_14793 (I255080,I1118173,I1118176);
nand I_14794 (I254760,I254896,I255080);
nand I_14795 (I254754,I254845,I1118173);
nand I_14796 (I255125,I254947,I1118170);
DFFARX1 I_14797 (I255125,I3563,I254780,I254769,);
DFFARX1 I_14798 (I255125,I3563,I254780,I254763,);
not I_14799 (I255170,I1118170);
nor I_14800 (I255187,I255170,I1118167);
and I_14801 (I255204,I255187,I1118185);
or I_14802 (I255221,I255204,I1118164);
DFFARX1 I_14803 (I255221,I3563,I254780,I255247,);
nand I_14804 (I255255,I255247,I254913);
nor I_14805 (I254757,I255255,I255063);
nor I_14806 (I254751,I255247,I254879);
DFFARX1 I_14807 (I255247,I3563,I254780,I255309,);
not I_14808 (I255317,I255309);
nor I_14809 (I254766,I255317,I255029);
not I_14810 (I255375,I3570);
DFFARX1 I_14811 (I11326,I3563,I255375,I255401,);
DFFARX1 I_14812 (I255401,I3563,I255375,I255418,);
not I_14813 (I255367,I255418);
not I_14814 (I255440,I255401);
DFFARX1 I_14815 (I11323,I3563,I255375,I255466,);
not I_14816 (I255474,I255466);
and I_14817 (I255491,I255440,I11314);
not I_14818 (I255508,I11311);
nand I_14819 (I255525,I255508,I11314);
not I_14820 (I255542,I11311);
nor I_14821 (I255559,I255542,I11308);
nand I_14822 (I255576,I255559,I11320);
nor I_14823 (I255593,I255576,I255525);
DFFARX1 I_14824 (I255593,I3563,I255375,I255343,);
not I_14825 (I255624,I255576);
not I_14826 (I255641,I11308);
nand I_14827 (I255658,I255641,I11314);
nor I_14828 (I255675,I11308,I11311);
nand I_14829 (I255355,I255491,I255675);
nand I_14830 (I255349,I255440,I11308);
nand I_14831 (I255720,I255542,I11317);
DFFARX1 I_14832 (I255720,I3563,I255375,I255364,);
DFFARX1 I_14833 (I255720,I3563,I255375,I255358,);
not I_14834 (I255765,I11317);
nor I_14835 (I255782,I255765,I11329);
and I_14836 (I255799,I255782,I11314);
or I_14837 (I255816,I255799,I11308);
DFFARX1 I_14838 (I255816,I3563,I255375,I255842,);
nand I_14839 (I255850,I255842,I255508);
nor I_14840 (I255352,I255850,I255658);
nor I_14841 (I255346,I255842,I255474);
DFFARX1 I_14842 (I255842,I3563,I255375,I255904,);
not I_14843 (I255912,I255904);
nor I_14844 (I255361,I255912,I255624);
not I_14845 (I255970,I3570);
DFFARX1 I_14846 (I1238963,I3563,I255970,I255996,);
DFFARX1 I_14847 (I255996,I3563,I255970,I256013,);
not I_14848 (I255962,I256013);
not I_14849 (I256035,I255996);
DFFARX1 I_14850 (I1238963,I3563,I255970,I256061,);
not I_14851 (I256069,I256061);
and I_14852 (I256086,I256035,I1238966);
not I_14853 (I256103,I1238978);
nand I_14854 (I256120,I256103,I1238966);
not I_14855 (I256137,I1238984);
nor I_14856 (I256154,I256137,I1238975);
nand I_14857 (I256171,I256154,I1238981);
nor I_14858 (I256188,I256171,I256120);
DFFARX1 I_14859 (I256188,I3563,I255970,I255938,);
not I_14860 (I256219,I256171);
not I_14861 (I256236,I1238975);
nand I_14862 (I256253,I256236,I1238966);
nor I_14863 (I256270,I1238975,I1238978);
nand I_14864 (I255950,I256086,I256270);
nand I_14865 (I255944,I256035,I1238975);
nand I_14866 (I256315,I256137,I1238972);
DFFARX1 I_14867 (I256315,I3563,I255970,I255959,);
DFFARX1 I_14868 (I256315,I3563,I255970,I255953,);
not I_14869 (I256360,I1238972);
nor I_14870 (I256377,I256360,I1238969);
and I_14871 (I256394,I256377,I1238987);
or I_14872 (I256411,I256394,I1238966);
DFFARX1 I_14873 (I256411,I3563,I255970,I256437,);
nand I_14874 (I256445,I256437,I256103);
nor I_14875 (I255947,I256445,I256253);
nor I_14876 (I255941,I256437,I256069);
DFFARX1 I_14877 (I256437,I3563,I255970,I256499,);
not I_14878 (I256507,I256499);
nor I_14879 (I255956,I256507,I256219);
not I_14880 (I256565,I3570);
DFFARX1 I_14881 (I418169,I3563,I256565,I256591,);
DFFARX1 I_14882 (I256591,I3563,I256565,I256608,);
not I_14883 (I256557,I256608);
not I_14884 (I256630,I256591);
DFFARX1 I_14885 (I418184,I3563,I256565,I256656,);
not I_14886 (I256664,I256656);
and I_14887 (I256681,I256630,I418181);
not I_14888 (I256698,I418169);
nand I_14889 (I256715,I256698,I418181);
not I_14890 (I256732,I418178);
nor I_14891 (I256749,I256732,I418193);
nand I_14892 (I256766,I256749,I418190);
nor I_14893 (I256783,I256766,I256715);
DFFARX1 I_14894 (I256783,I3563,I256565,I256533,);
not I_14895 (I256814,I256766);
not I_14896 (I256831,I418193);
nand I_14897 (I256848,I256831,I418181);
nor I_14898 (I256865,I418193,I418169);
nand I_14899 (I256545,I256681,I256865);
nand I_14900 (I256539,I256630,I418193);
nand I_14901 (I256910,I256732,I418187);
DFFARX1 I_14902 (I256910,I3563,I256565,I256554,);
DFFARX1 I_14903 (I256910,I3563,I256565,I256548,);
not I_14904 (I256955,I418187);
nor I_14905 (I256972,I256955,I418175);
and I_14906 (I256989,I256972,I418196);
or I_14907 (I257006,I256989,I418172);
DFFARX1 I_14908 (I257006,I3563,I256565,I257032,);
nand I_14909 (I257040,I257032,I256698);
nor I_14910 (I256542,I257040,I256848);
nor I_14911 (I256536,I257032,I256664);
DFFARX1 I_14912 (I257032,I3563,I256565,I257094,);
not I_14913 (I257102,I257094);
nor I_14914 (I256551,I257102,I256814);
not I_14915 (I257160,I3570);
DFFARX1 I_14916 (I774603,I3563,I257160,I257186,);
DFFARX1 I_14917 (I257186,I3563,I257160,I257203,);
not I_14918 (I257152,I257203);
not I_14919 (I257225,I257186);
DFFARX1 I_14920 (I774600,I3563,I257160,I257251,);
not I_14921 (I257259,I257251);
and I_14922 (I257276,I257225,I774606);
not I_14923 (I257293,I774591);
nand I_14924 (I257310,I257293,I774606);
not I_14925 (I257327,I774594);
nor I_14926 (I257344,I257327,I774615);
nand I_14927 (I257361,I257344,I774612);
nor I_14928 (I257378,I257361,I257310);
DFFARX1 I_14929 (I257378,I3563,I257160,I257128,);
not I_14930 (I257409,I257361);
not I_14931 (I257426,I774615);
nand I_14932 (I257443,I257426,I774606);
nor I_14933 (I257460,I774615,I774591);
nand I_14934 (I257140,I257276,I257460);
nand I_14935 (I257134,I257225,I774615);
nand I_14936 (I257505,I257327,I774591);
DFFARX1 I_14937 (I257505,I3563,I257160,I257149,);
DFFARX1 I_14938 (I257505,I3563,I257160,I257143,);
not I_14939 (I257550,I774591);
nor I_14940 (I257567,I257550,I774597);
and I_14941 (I257584,I257567,I774609);
or I_14942 (I257601,I257584,I774594);
DFFARX1 I_14943 (I257601,I3563,I257160,I257627,);
nand I_14944 (I257635,I257627,I257293);
nor I_14945 (I257137,I257635,I257443);
nor I_14946 (I257131,I257627,I257259);
DFFARX1 I_14947 (I257627,I3563,I257160,I257689,);
not I_14948 (I257697,I257689);
nor I_14949 (I257146,I257697,I257409);
not I_14950 (I257755,I3570);
DFFARX1 I_14951 (I44023,I3563,I257755,I257781,);
DFFARX1 I_14952 (I257781,I3563,I257755,I257798,);
not I_14953 (I257747,I257798);
not I_14954 (I257820,I257781);
DFFARX1 I_14955 (I43999,I3563,I257755,I257846,);
not I_14956 (I257854,I257846);
and I_14957 (I257871,I257820,I44014);
not I_14958 (I257888,I44002);
nand I_14959 (I257905,I257888,I44014);
not I_14960 (I257922,I44005);
nor I_14961 (I257939,I257922,I44017);
nand I_14962 (I257956,I257939,I44008);
nor I_14963 (I257973,I257956,I257905);
DFFARX1 I_14964 (I257973,I3563,I257755,I257723,);
not I_14965 (I258004,I257956);
not I_14966 (I258021,I44017);
nand I_14967 (I258038,I258021,I44014);
nor I_14968 (I258055,I44017,I44002);
nand I_14969 (I257735,I257871,I258055);
nand I_14970 (I257729,I257820,I44017);
nand I_14971 (I258100,I257922,I44011);
DFFARX1 I_14972 (I258100,I3563,I257755,I257744,);
DFFARX1 I_14973 (I258100,I3563,I257755,I257738,);
not I_14974 (I258145,I44011);
nor I_14975 (I258162,I258145,I44002);
and I_14976 (I258179,I258162,I43999);
or I_14977 (I258196,I258179,I44020);
DFFARX1 I_14978 (I258196,I3563,I257755,I258222,);
nand I_14979 (I258230,I258222,I257888);
nor I_14980 (I257732,I258230,I258038);
nor I_14981 (I257726,I258222,I257854);
DFFARX1 I_14982 (I258222,I3563,I257755,I258284,);
not I_14983 (I258292,I258284);
nor I_14984 (I257741,I258292,I258004);
not I_14985 (I258350,I3570);
DFFARX1 I_14986 (I995640,I3563,I258350,I258376,);
DFFARX1 I_14987 (I258376,I3563,I258350,I258393,);
not I_14988 (I258342,I258393);
not I_14989 (I258415,I258376);
DFFARX1 I_14990 (I995649,I3563,I258350,I258441,);
not I_14991 (I258449,I258441);
and I_14992 (I258466,I258415,I995637);
not I_14993 (I258483,I995628);
nand I_14994 (I258500,I258483,I995637);
not I_14995 (I258517,I995634);
nor I_14996 (I258534,I258517,I995652);
nand I_14997 (I258551,I258534,I995625);
nor I_14998 (I258568,I258551,I258500);
DFFARX1 I_14999 (I258568,I3563,I258350,I258318,);
not I_15000 (I258599,I258551);
not I_15001 (I258616,I995652);
nand I_15002 (I258633,I258616,I995637);
nor I_15003 (I258650,I995652,I995628);
nand I_15004 (I258330,I258466,I258650);
nand I_15005 (I258324,I258415,I995652);
nand I_15006 (I258695,I258517,I995631);
DFFARX1 I_15007 (I258695,I3563,I258350,I258339,);
DFFARX1 I_15008 (I258695,I3563,I258350,I258333,);
not I_15009 (I258740,I995631);
nor I_15010 (I258757,I258740,I995643);
and I_15011 (I258774,I258757,I995625);
or I_15012 (I258791,I258774,I995646);
DFFARX1 I_15013 (I258791,I3563,I258350,I258817,);
nand I_15014 (I258825,I258817,I258483);
nor I_15015 (I258327,I258825,I258633);
nor I_15016 (I258321,I258817,I258449);
DFFARX1 I_15017 (I258817,I3563,I258350,I258879,);
not I_15018 (I258887,I258879);
nor I_15019 (I258336,I258887,I258599);
not I_15020 (I258945,I3570);
DFFARX1 I_15021 (I763043,I3563,I258945,I258971,);
DFFARX1 I_15022 (I258971,I3563,I258945,I258988,);
not I_15023 (I258937,I258988);
not I_15024 (I259010,I258971);
DFFARX1 I_15025 (I763040,I3563,I258945,I259036,);
not I_15026 (I259044,I259036);
and I_15027 (I259061,I259010,I763046);
not I_15028 (I259078,I763031);
nand I_15029 (I259095,I259078,I763046);
not I_15030 (I259112,I763034);
nor I_15031 (I259129,I259112,I763055);
nand I_15032 (I259146,I259129,I763052);
nor I_15033 (I259163,I259146,I259095);
DFFARX1 I_15034 (I259163,I3563,I258945,I258913,);
not I_15035 (I259194,I259146);
not I_15036 (I259211,I763055);
nand I_15037 (I259228,I259211,I763046);
nor I_15038 (I259245,I763055,I763031);
nand I_15039 (I258925,I259061,I259245);
nand I_15040 (I258919,I259010,I763055);
nand I_15041 (I259290,I259112,I763031);
DFFARX1 I_15042 (I259290,I3563,I258945,I258934,);
DFFARX1 I_15043 (I259290,I3563,I258945,I258928,);
not I_15044 (I259335,I763031);
nor I_15045 (I259352,I259335,I763037);
and I_15046 (I259369,I259352,I763049);
or I_15047 (I259386,I259369,I763034);
DFFARX1 I_15048 (I259386,I3563,I258945,I259412,);
nand I_15049 (I259420,I259412,I259078);
nor I_15050 (I258922,I259420,I259228);
nor I_15051 (I258916,I259412,I259044);
DFFARX1 I_15052 (I259412,I3563,I258945,I259474,);
not I_15053 (I259482,I259474);
nor I_15054 (I258931,I259482,I259194);
not I_15055 (I259540,I3570);
DFFARX1 I_15056 (I869032,I3563,I259540,I259566,);
DFFARX1 I_15057 (I259566,I3563,I259540,I259583,);
not I_15058 (I259532,I259583);
not I_15059 (I259605,I259566);
DFFARX1 I_15060 (I869026,I3563,I259540,I259631,);
not I_15061 (I259639,I259631);
and I_15062 (I259656,I259605,I869044);
not I_15063 (I259673,I869032);
nand I_15064 (I259690,I259673,I869044);
not I_15065 (I259707,I869026);
nor I_15066 (I259724,I259707,I869038);
nand I_15067 (I259741,I259724,I869029);
nor I_15068 (I259758,I259741,I259690);
DFFARX1 I_15069 (I259758,I3563,I259540,I259508,);
not I_15070 (I259789,I259741);
not I_15071 (I259806,I869038);
nand I_15072 (I259823,I259806,I869044);
nor I_15073 (I259840,I869038,I869032);
nand I_15074 (I259520,I259656,I259840);
nand I_15075 (I259514,I259605,I869038);
nand I_15076 (I259885,I259707,I869041);
DFFARX1 I_15077 (I259885,I3563,I259540,I259529,);
DFFARX1 I_15078 (I259885,I3563,I259540,I259523,);
not I_15079 (I259930,I869041);
nor I_15080 (I259947,I259930,I869047);
and I_15081 (I259964,I259947,I869029);
or I_15082 (I259981,I259964,I869035);
DFFARX1 I_15083 (I259981,I3563,I259540,I260007,);
nand I_15084 (I260015,I260007,I259673);
nor I_15085 (I259517,I260015,I259823);
nor I_15086 (I259511,I260007,I259639);
DFFARX1 I_15087 (I260007,I3563,I259540,I260069,);
not I_15088 (I260077,I260069);
nor I_15089 (I259526,I260077,I259789);
not I_15090 (I260135,I3570);
DFFARX1 I_15091 (I301702,I3563,I260135,I260161,);
DFFARX1 I_15092 (I260161,I3563,I260135,I260178,);
not I_15093 (I260127,I260178);
not I_15094 (I260200,I260161);
DFFARX1 I_15095 (I301717,I3563,I260135,I260226,);
not I_15096 (I260234,I260226);
and I_15097 (I260251,I260200,I301714);
not I_15098 (I260268,I301702);
nand I_15099 (I260285,I260268,I301714);
not I_15100 (I260302,I301711);
nor I_15101 (I260319,I260302,I301726);
nand I_15102 (I260336,I260319,I301723);
nor I_15103 (I260353,I260336,I260285);
DFFARX1 I_15104 (I260353,I3563,I260135,I260103,);
not I_15105 (I260384,I260336);
not I_15106 (I260401,I301726);
nand I_15107 (I260418,I260401,I301714);
nor I_15108 (I260435,I301726,I301702);
nand I_15109 (I260115,I260251,I260435);
nand I_15110 (I260109,I260200,I301726);
nand I_15111 (I260480,I260302,I301720);
DFFARX1 I_15112 (I260480,I3563,I260135,I260124,);
DFFARX1 I_15113 (I260480,I3563,I260135,I260118,);
not I_15114 (I260525,I301720);
nor I_15115 (I260542,I260525,I301708);
and I_15116 (I260559,I260542,I301729);
or I_15117 (I260576,I260559,I301705);
DFFARX1 I_15118 (I260576,I3563,I260135,I260602,);
nand I_15119 (I260610,I260602,I260268);
nor I_15120 (I260112,I260610,I260418);
nor I_15121 (I260106,I260602,I260234);
DFFARX1 I_15122 (I260602,I3563,I260135,I260664,);
not I_15123 (I260672,I260664);
nor I_15124 (I260121,I260672,I260384);
not I_15125 (I260730,I3570);
DFFARX1 I_15126 (I1243587,I3563,I260730,I260756,);
DFFARX1 I_15127 (I260756,I3563,I260730,I260773,);
not I_15128 (I260722,I260773);
not I_15129 (I260795,I260756);
DFFARX1 I_15130 (I1243587,I3563,I260730,I260821,);
not I_15131 (I260829,I260821);
and I_15132 (I260846,I260795,I1243590);
not I_15133 (I260863,I1243602);
nand I_15134 (I260880,I260863,I1243590);
not I_15135 (I260897,I1243608);
nor I_15136 (I260914,I260897,I1243599);
nand I_15137 (I260931,I260914,I1243605);
nor I_15138 (I260948,I260931,I260880);
DFFARX1 I_15139 (I260948,I3563,I260730,I260698,);
not I_15140 (I260979,I260931);
not I_15141 (I260996,I1243599);
nand I_15142 (I261013,I260996,I1243590);
nor I_15143 (I261030,I1243599,I1243602);
nand I_15144 (I260710,I260846,I261030);
nand I_15145 (I260704,I260795,I1243599);
nand I_15146 (I261075,I260897,I1243596);
DFFARX1 I_15147 (I261075,I3563,I260730,I260719,);
DFFARX1 I_15148 (I261075,I3563,I260730,I260713,);
not I_15149 (I261120,I1243596);
nor I_15150 (I261137,I261120,I1243593);
and I_15151 (I261154,I261137,I1243611);
or I_15152 (I261171,I261154,I1243590);
DFFARX1 I_15153 (I261171,I3563,I260730,I261197,);
nand I_15154 (I261205,I261197,I260863);
nor I_15155 (I260707,I261205,I261013);
nor I_15156 (I260701,I261197,I260829);
DFFARX1 I_15157 (I261197,I3563,I260730,I261259,);
not I_15158 (I261267,I261259);
nor I_15159 (I260716,I261267,I260979);
not I_15160 (I261325,I3570);
DFFARX1 I_15161 (I12516,I3563,I261325,I261351,);
DFFARX1 I_15162 (I261351,I3563,I261325,I261368,);
not I_15163 (I261317,I261368);
not I_15164 (I261390,I261351);
DFFARX1 I_15165 (I12513,I3563,I261325,I261416,);
not I_15166 (I261424,I261416);
and I_15167 (I261441,I261390,I12504);
not I_15168 (I261458,I12501);
nand I_15169 (I261475,I261458,I12504);
not I_15170 (I261492,I12501);
nor I_15171 (I261509,I261492,I12498);
nand I_15172 (I261526,I261509,I12510);
nor I_15173 (I261543,I261526,I261475);
DFFARX1 I_15174 (I261543,I3563,I261325,I261293,);
not I_15175 (I261574,I261526);
not I_15176 (I261591,I12498);
nand I_15177 (I261608,I261591,I12504);
nor I_15178 (I261625,I12498,I12501);
nand I_15179 (I261305,I261441,I261625);
nand I_15180 (I261299,I261390,I12498);
nand I_15181 (I261670,I261492,I12507);
DFFARX1 I_15182 (I261670,I3563,I261325,I261314,);
DFFARX1 I_15183 (I261670,I3563,I261325,I261308,);
not I_15184 (I261715,I12507);
nor I_15185 (I261732,I261715,I12519);
and I_15186 (I261749,I261732,I12504);
or I_15187 (I261766,I261749,I12498);
DFFARX1 I_15188 (I261766,I3563,I261325,I261792,);
nand I_15189 (I261800,I261792,I261458);
nor I_15190 (I261302,I261800,I261608);
nor I_15191 (I261296,I261792,I261424);
DFFARX1 I_15192 (I261792,I3563,I261325,I261854,);
not I_15193 (I261862,I261854);
nor I_15194 (I261311,I261862,I261574);
not I_15195 (I261920,I3570);
DFFARX1 I_15196 (I956880,I3563,I261920,I261946,);
DFFARX1 I_15197 (I261946,I3563,I261920,I261963,);
not I_15198 (I261912,I261963);
not I_15199 (I261985,I261946);
DFFARX1 I_15200 (I956889,I3563,I261920,I262011,);
not I_15201 (I262019,I262011);
and I_15202 (I262036,I261985,I956877);
not I_15203 (I262053,I956868);
nand I_15204 (I262070,I262053,I956877);
not I_15205 (I262087,I956874);
nor I_15206 (I262104,I262087,I956892);
nand I_15207 (I262121,I262104,I956865);
nor I_15208 (I262138,I262121,I262070);
DFFARX1 I_15209 (I262138,I3563,I261920,I261888,);
not I_15210 (I262169,I262121);
not I_15211 (I262186,I956892);
nand I_15212 (I262203,I262186,I956877);
nor I_15213 (I262220,I956892,I956868);
nand I_15214 (I261900,I262036,I262220);
nand I_15215 (I261894,I261985,I956892);
nand I_15216 (I262265,I262087,I956871);
DFFARX1 I_15217 (I262265,I3563,I261920,I261909,);
DFFARX1 I_15218 (I262265,I3563,I261920,I261903,);
not I_15219 (I262310,I956871);
nor I_15220 (I262327,I262310,I956883);
and I_15221 (I262344,I262327,I956865);
or I_15222 (I262361,I262344,I956886);
DFFARX1 I_15223 (I262361,I3563,I261920,I262387,);
nand I_15224 (I262395,I262387,I262053);
nor I_15225 (I261897,I262395,I262203);
nor I_15226 (I261891,I262387,I262019);
DFFARX1 I_15227 (I262387,I3563,I261920,I262449,);
not I_15228 (I262457,I262449);
nor I_15229 (I261906,I262457,I262169);
not I_15230 (I262515,I3570);
DFFARX1 I_15231 (I1228559,I3563,I262515,I262541,);
DFFARX1 I_15232 (I262541,I3563,I262515,I262558,);
not I_15233 (I262507,I262558);
not I_15234 (I262580,I262541);
DFFARX1 I_15235 (I1228559,I3563,I262515,I262606,);
not I_15236 (I262614,I262606);
and I_15237 (I262631,I262580,I1228562);
not I_15238 (I262648,I1228574);
nand I_15239 (I262665,I262648,I1228562);
not I_15240 (I262682,I1228580);
nor I_15241 (I262699,I262682,I1228571);
nand I_15242 (I262716,I262699,I1228577);
nor I_15243 (I262733,I262716,I262665);
DFFARX1 I_15244 (I262733,I3563,I262515,I262483,);
not I_15245 (I262764,I262716);
not I_15246 (I262781,I1228571);
nand I_15247 (I262798,I262781,I1228562);
nor I_15248 (I262815,I1228571,I1228574);
nand I_15249 (I262495,I262631,I262815);
nand I_15250 (I262489,I262580,I1228571);
nand I_15251 (I262860,I262682,I1228568);
DFFARX1 I_15252 (I262860,I3563,I262515,I262504,);
DFFARX1 I_15253 (I262860,I3563,I262515,I262498,);
not I_15254 (I262905,I1228568);
nor I_15255 (I262922,I262905,I1228565);
and I_15256 (I262939,I262922,I1228583);
or I_15257 (I262956,I262939,I1228562);
DFFARX1 I_15258 (I262956,I3563,I262515,I262982,);
nand I_15259 (I262990,I262982,I262648);
nor I_15260 (I262492,I262990,I262798);
nor I_15261 (I262486,I262982,I262614);
DFFARX1 I_15262 (I262982,I3563,I262515,I263044,);
not I_15263 (I263052,I263044);
nor I_15264 (I262501,I263052,I262764);
not I_15265 (I263110,I3570);
DFFARX1 I_15266 (I2524,I3563,I263110,I263136,);
DFFARX1 I_15267 (I263136,I3563,I263110,I263153,);
not I_15268 (I263102,I263153);
not I_15269 (I263175,I263136);
DFFARX1 I_15270 (I3108,I3563,I263110,I263201,);
not I_15271 (I263209,I263201);
and I_15272 (I263226,I263175,I1676);
not I_15273 (I263243,I3524);
nand I_15274 (I263260,I263243,I1676);
not I_15275 (I263277,I1636);
nor I_15276 (I263294,I263277,I2132);
nand I_15277 (I263311,I263294,I3332);
nor I_15278 (I263328,I263311,I263260);
DFFARX1 I_15279 (I263328,I3563,I263110,I263078,);
not I_15280 (I263359,I263311);
not I_15281 (I263376,I2132);
nand I_15282 (I263393,I263376,I1676);
nor I_15283 (I263410,I2132,I3524);
nand I_15284 (I263090,I263226,I263410);
nand I_15285 (I263084,I263175,I2132);
nand I_15286 (I263455,I263277,I1444);
DFFARX1 I_15287 (I263455,I3563,I263110,I263099,);
DFFARX1 I_15288 (I263455,I3563,I263110,I263093,);
not I_15289 (I263500,I1444);
nor I_15290 (I263517,I263500,I3012);
and I_15291 (I263534,I263517,I1860);
or I_15292 (I263551,I263534,I2900);
DFFARX1 I_15293 (I263551,I3563,I263110,I263577,);
nand I_15294 (I263585,I263577,I263243);
nor I_15295 (I263087,I263585,I263393);
nor I_15296 (I263081,I263577,I263209);
DFFARX1 I_15297 (I263577,I3563,I263110,I263639,);
not I_15298 (I263647,I263639);
nor I_15299 (I263096,I263647,I263359);
not I_15300 (I263705,I3570);
DFFARX1 I_15301 (I681545,I3563,I263705,I263731,);
DFFARX1 I_15302 (I263731,I3563,I263705,I263748,);
not I_15303 (I263697,I263748);
not I_15304 (I263770,I263731);
DFFARX1 I_15305 (I681542,I3563,I263705,I263796,);
not I_15306 (I263804,I263796);
and I_15307 (I263821,I263770,I681548);
not I_15308 (I263838,I681533);
nand I_15309 (I263855,I263838,I681548);
not I_15310 (I263872,I681536);
nor I_15311 (I263889,I263872,I681557);
nand I_15312 (I263906,I263889,I681554);
nor I_15313 (I263923,I263906,I263855);
DFFARX1 I_15314 (I263923,I3563,I263705,I263673,);
not I_15315 (I263954,I263906);
not I_15316 (I263971,I681557);
nand I_15317 (I263988,I263971,I681548);
nor I_15318 (I264005,I681557,I681533);
nand I_15319 (I263685,I263821,I264005);
nand I_15320 (I263679,I263770,I681557);
nand I_15321 (I264050,I263872,I681533);
DFFARX1 I_15322 (I264050,I3563,I263705,I263694,);
DFFARX1 I_15323 (I264050,I3563,I263705,I263688,);
not I_15324 (I264095,I681533);
nor I_15325 (I264112,I264095,I681539);
and I_15326 (I264129,I264112,I681551);
or I_15327 (I264146,I264129,I681536);
DFFARX1 I_15328 (I264146,I3563,I263705,I264172,);
nand I_15329 (I264180,I264172,I263838);
nor I_15330 (I263682,I264180,I263988);
nor I_15331 (I263676,I264172,I263804);
DFFARX1 I_15332 (I264172,I3563,I263705,I264234,);
not I_15333 (I264242,I264234);
nor I_15334 (I263691,I264242,I263954);
not I_15335 (I264300,I3570);
DFFARX1 I_15336 (I417115,I3563,I264300,I264326,);
DFFARX1 I_15337 (I264326,I3563,I264300,I264343,);
not I_15338 (I264292,I264343);
not I_15339 (I264365,I264326);
DFFARX1 I_15340 (I417130,I3563,I264300,I264391,);
not I_15341 (I264399,I264391);
and I_15342 (I264416,I264365,I417127);
not I_15343 (I264433,I417115);
nand I_15344 (I264450,I264433,I417127);
not I_15345 (I264467,I417124);
nor I_15346 (I264484,I264467,I417139);
nand I_15347 (I264501,I264484,I417136);
nor I_15348 (I264518,I264501,I264450);
DFFARX1 I_15349 (I264518,I3563,I264300,I264268,);
not I_15350 (I264549,I264501);
not I_15351 (I264566,I417139);
nand I_15352 (I264583,I264566,I417127);
nor I_15353 (I264600,I417139,I417115);
nand I_15354 (I264280,I264416,I264600);
nand I_15355 (I264274,I264365,I417139);
nand I_15356 (I264645,I264467,I417133);
DFFARX1 I_15357 (I264645,I3563,I264300,I264289,);
DFFARX1 I_15358 (I264645,I3563,I264300,I264283,);
not I_15359 (I264690,I417133);
nor I_15360 (I264707,I264690,I417121);
and I_15361 (I264724,I264707,I417142);
or I_15362 (I264741,I264724,I417118);
DFFARX1 I_15363 (I264741,I3563,I264300,I264767,);
nand I_15364 (I264775,I264767,I264433);
nor I_15365 (I264277,I264775,I264583);
nor I_15366 (I264271,I264767,I264399);
DFFARX1 I_15367 (I264767,I3563,I264300,I264829,);
not I_15368 (I264837,I264829);
nor I_15369 (I264286,I264837,I264549);
not I_15370 (I264895,I3570);
DFFARX1 I_15371 (I931040,I3563,I264895,I264921,);
DFFARX1 I_15372 (I264921,I3563,I264895,I264938,);
not I_15373 (I264887,I264938);
not I_15374 (I264960,I264921);
DFFARX1 I_15375 (I931049,I3563,I264895,I264986,);
not I_15376 (I264994,I264986);
and I_15377 (I265011,I264960,I931037);
not I_15378 (I265028,I931028);
nand I_15379 (I265045,I265028,I931037);
not I_15380 (I265062,I931034);
nor I_15381 (I265079,I265062,I931052);
nand I_15382 (I265096,I265079,I931025);
nor I_15383 (I265113,I265096,I265045);
DFFARX1 I_15384 (I265113,I3563,I264895,I264863,);
not I_15385 (I265144,I265096);
not I_15386 (I265161,I931052);
nand I_15387 (I265178,I265161,I931037);
nor I_15388 (I265195,I931052,I931028);
nand I_15389 (I264875,I265011,I265195);
nand I_15390 (I264869,I264960,I931052);
nand I_15391 (I265240,I265062,I931031);
DFFARX1 I_15392 (I265240,I3563,I264895,I264884,);
DFFARX1 I_15393 (I265240,I3563,I264895,I264878,);
not I_15394 (I265285,I931031);
nor I_15395 (I265302,I265285,I931043);
and I_15396 (I265319,I265302,I931025);
or I_15397 (I265336,I265319,I931046);
DFFARX1 I_15398 (I265336,I3563,I264895,I265362,);
nand I_15399 (I265370,I265362,I265028);
nor I_15400 (I264872,I265370,I265178);
nor I_15401 (I264866,I265362,I264994);
DFFARX1 I_15402 (I265362,I3563,I264895,I265424,);
not I_15403 (I265432,I265424);
nor I_15404 (I264881,I265432,I265144);
not I_15405 (I265490,I3570);
DFFARX1 I_15406 (I1013728,I3563,I265490,I265516,);
DFFARX1 I_15407 (I265516,I3563,I265490,I265533,);
not I_15408 (I265482,I265533);
not I_15409 (I265555,I265516);
DFFARX1 I_15410 (I1013737,I3563,I265490,I265581,);
not I_15411 (I265589,I265581);
and I_15412 (I265606,I265555,I1013725);
not I_15413 (I265623,I1013716);
nand I_15414 (I265640,I265623,I1013725);
not I_15415 (I265657,I1013722);
nor I_15416 (I265674,I265657,I1013740);
nand I_15417 (I265691,I265674,I1013713);
nor I_15418 (I265708,I265691,I265640);
DFFARX1 I_15419 (I265708,I3563,I265490,I265458,);
not I_15420 (I265739,I265691);
not I_15421 (I265756,I1013740);
nand I_15422 (I265773,I265756,I1013725);
nor I_15423 (I265790,I1013740,I1013716);
nand I_15424 (I265470,I265606,I265790);
nand I_15425 (I265464,I265555,I1013740);
nand I_15426 (I265835,I265657,I1013719);
DFFARX1 I_15427 (I265835,I3563,I265490,I265479,);
DFFARX1 I_15428 (I265835,I3563,I265490,I265473,);
not I_15429 (I265880,I1013719);
nor I_15430 (I265897,I265880,I1013731);
and I_15431 (I265914,I265897,I1013713);
or I_15432 (I265931,I265914,I1013734);
DFFARX1 I_15433 (I265931,I3563,I265490,I265957,);
nand I_15434 (I265965,I265957,I265623);
nor I_15435 (I265467,I265965,I265773);
nor I_15436 (I265461,I265957,I265589);
DFFARX1 I_15437 (I265957,I3563,I265490,I266019,);
not I_15438 (I266027,I266019);
nor I_15439 (I265476,I266027,I265739);
not I_15440 (I266085,I3570);
DFFARX1 I_15441 (I32956,I3563,I266085,I266111,);
DFFARX1 I_15442 (I266111,I3563,I266085,I266128,);
not I_15443 (I266077,I266128);
not I_15444 (I266150,I266111);
DFFARX1 I_15445 (I32932,I3563,I266085,I266176,);
not I_15446 (I266184,I266176);
and I_15447 (I266201,I266150,I32947);
not I_15448 (I266218,I32935);
nand I_15449 (I266235,I266218,I32947);
not I_15450 (I266252,I32938);
nor I_15451 (I266269,I266252,I32950);
nand I_15452 (I266286,I266269,I32941);
nor I_15453 (I266303,I266286,I266235);
DFFARX1 I_15454 (I266303,I3563,I266085,I266053,);
not I_15455 (I266334,I266286);
not I_15456 (I266351,I32950);
nand I_15457 (I266368,I266351,I32947);
nor I_15458 (I266385,I32950,I32935);
nand I_15459 (I266065,I266201,I266385);
nand I_15460 (I266059,I266150,I32950);
nand I_15461 (I266430,I266252,I32944);
DFFARX1 I_15462 (I266430,I3563,I266085,I266074,);
DFFARX1 I_15463 (I266430,I3563,I266085,I266068,);
not I_15464 (I266475,I32944);
nor I_15465 (I266492,I266475,I32935);
and I_15466 (I266509,I266492,I32932);
or I_15467 (I266526,I266509,I32953);
DFFARX1 I_15468 (I266526,I3563,I266085,I266552,);
nand I_15469 (I266560,I266552,I266218);
nor I_15470 (I266062,I266560,I266368);
nor I_15471 (I266056,I266552,I266184);
DFFARX1 I_15472 (I266552,I3563,I266085,I266614,);
not I_15473 (I266622,I266614);
nor I_15474 (I266071,I266622,I266334);
not I_15475 (I266680,I3570);
DFFARX1 I_15476 (I1266555,I3563,I266680,I266706,);
DFFARX1 I_15477 (I266706,I3563,I266680,I266723,);
not I_15478 (I266672,I266723);
not I_15479 (I266745,I266706);
DFFARX1 I_15480 (I1266540,I3563,I266680,I266771,);
not I_15481 (I266779,I266771);
and I_15482 (I266796,I266745,I1266558);
not I_15483 (I266813,I1266540);
nand I_15484 (I266830,I266813,I1266558);
not I_15485 (I266847,I1266561);
nor I_15486 (I266864,I266847,I1266552);
nand I_15487 (I266881,I266864,I1266549);
nor I_15488 (I266898,I266881,I266830);
DFFARX1 I_15489 (I266898,I3563,I266680,I266648,);
not I_15490 (I266929,I266881);
not I_15491 (I266946,I1266552);
nand I_15492 (I266963,I266946,I1266558);
nor I_15493 (I266980,I1266552,I1266540);
nand I_15494 (I266660,I266796,I266980);
nand I_15495 (I266654,I266745,I1266552);
nand I_15496 (I267025,I266847,I1266546);
DFFARX1 I_15497 (I267025,I3563,I266680,I266669,);
DFFARX1 I_15498 (I267025,I3563,I266680,I266663,);
not I_15499 (I267070,I1266546);
nor I_15500 (I267087,I267070,I1266537);
and I_15501 (I267104,I267087,I1266543);
or I_15502 (I267121,I267104,I1266537);
DFFARX1 I_15503 (I267121,I3563,I266680,I267147,);
nand I_15504 (I267155,I267147,I266813);
nor I_15505 (I266657,I267155,I266963);
nor I_15506 (I266651,I267147,I266779);
DFFARX1 I_15507 (I267147,I3563,I266680,I267209,);
not I_15508 (I267217,I267209);
nor I_15509 (I266666,I267217,I266929);
not I_15510 (I267275,I3570);
DFFARX1 I_15511 (I836358,I3563,I267275,I267301,);
DFFARX1 I_15512 (I267301,I3563,I267275,I267318,);
not I_15513 (I267267,I267318);
not I_15514 (I267340,I267301);
DFFARX1 I_15515 (I836352,I3563,I267275,I267366,);
not I_15516 (I267374,I267366);
and I_15517 (I267391,I267340,I836370);
not I_15518 (I267408,I836358);
nand I_15519 (I267425,I267408,I836370);
not I_15520 (I267442,I836352);
nor I_15521 (I267459,I267442,I836364);
nand I_15522 (I267476,I267459,I836355);
nor I_15523 (I267493,I267476,I267425);
DFFARX1 I_15524 (I267493,I3563,I267275,I267243,);
not I_15525 (I267524,I267476);
not I_15526 (I267541,I836364);
nand I_15527 (I267558,I267541,I836370);
nor I_15528 (I267575,I836364,I836358);
nand I_15529 (I267255,I267391,I267575);
nand I_15530 (I267249,I267340,I836364);
nand I_15531 (I267620,I267442,I836367);
DFFARX1 I_15532 (I267620,I3563,I267275,I267264,);
DFFARX1 I_15533 (I267620,I3563,I267275,I267258,);
not I_15534 (I267665,I836367);
nor I_15535 (I267682,I267665,I836373);
and I_15536 (I267699,I267682,I836355);
or I_15537 (I267716,I267699,I836361);
DFFARX1 I_15538 (I267716,I3563,I267275,I267742,);
nand I_15539 (I267750,I267742,I267408);
nor I_15540 (I267252,I267750,I267558);
nor I_15541 (I267246,I267742,I267374);
DFFARX1 I_15542 (I267742,I3563,I267275,I267804,);
not I_15543 (I267812,I267804);
nor I_15544 (I267261,I267812,I267524);
not I_15545 (I267870,I3570);
DFFARX1 I_15546 (I1386289,I3563,I267870,I267896,);
DFFARX1 I_15547 (I267896,I3563,I267870,I267913,);
not I_15548 (I267862,I267913);
not I_15549 (I267935,I267896);
DFFARX1 I_15550 (I1386280,I3563,I267870,I267961,);
not I_15551 (I267969,I267961);
and I_15552 (I267986,I267935,I1386274);
not I_15553 (I268003,I1386268);
nand I_15554 (I268020,I268003,I1386274);
not I_15555 (I268037,I1386295);
nor I_15556 (I268054,I268037,I1386268);
nand I_15557 (I268071,I268054,I1386292);
nor I_15558 (I268088,I268071,I268020);
DFFARX1 I_15559 (I268088,I3563,I267870,I267838,);
not I_15560 (I268119,I268071);
not I_15561 (I268136,I1386268);
nand I_15562 (I268153,I268136,I1386274);
nor I_15563 (I268170,I1386268,I1386268);
nand I_15564 (I267850,I267986,I268170);
nand I_15565 (I267844,I267935,I1386268);
nand I_15566 (I268215,I268037,I1386277);
DFFARX1 I_15567 (I268215,I3563,I267870,I267859,);
DFFARX1 I_15568 (I268215,I3563,I267870,I267853,);
not I_15569 (I268260,I1386277);
nor I_15570 (I268277,I268260,I1386283);
and I_15571 (I268294,I268277,I1386286);
or I_15572 (I268311,I268294,I1386271);
DFFARX1 I_15573 (I268311,I3563,I267870,I268337,);
nand I_15574 (I268345,I268337,I268003);
nor I_15575 (I267847,I268345,I268153);
nor I_15576 (I267841,I268337,I267969);
DFFARX1 I_15577 (I268337,I3563,I267870,I268399,);
not I_15578 (I268407,I268399);
nor I_15579 (I267856,I268407,I268119);
not I_15580 (I268465,I3570);
DFFARX1 I_15581 (I601784,I3563,I268465,I268491,);
DFFARX1 I_15582 (I268491,I3563,I268465,I268508,);
not I_15583 (I268457,I268508);
not I_15584 (I268530,I268491);
DFFARX1 I_15585 (I601775,I3563,I268465,I268556,);
not I_15586 (I268564,I268556);
and I_15587 (I268581,I268530,I601793);
not I_15588 (I268598,I601790);
nand I_15589 (I268615,I268598,I601793);
not I_15590 (I268632,I601769);
nor I_15591 (I268649,I268632,I601772);
nand I_15592 (I268666,I268649,I601781);
nor I_15593 (I268683,I268666,I268615);
DFFARX1 I_15594 (I268683,I3563,I268465,I268433,);
not I_15595 (I268714,I268666);
not I_15596 (I268731,I601772);
nand I_15597 (I268748,I268731,I601793);
nor I_15598 (I268765,I601772,I601790);
nand I_15599 (I268445,I268581,I268765);
nand I_15600 (I268439,I268530,I601772);
nand I_15601 (I268810,I268632,I601787);
DFFARX1 I_15602 (I268810,I3563,I268465,I268454,);
DFFARX1 I_15603 (I268810,I3563,I268465,I268448,);
not I_15604 (I268855,I601787);
nor I_15605 (I268872,I268855,I601769);
and I_15606 (I268889,I268872,I601778);
or I_15607 (I268906,I268889,I601772);
DFFARX1 I_15608 (I268906,I3563,I268465,I268932,);
nand I_15609 (I268940,I268932,I268598);
nor I_15610 (I268442,I268940,I268748);
nor I_15611 (I268436,I268932,I268564);
DFFARX1 I_15612 (I268932,I3563,I268465,I268994,);
not I_15613 (I269002,I268994);
nor I_15614 (I268451,I269002,I268714);
not I_15615 (I269060,I3570);
DFFARX1 I_15616 (I673453,I3563,I269060,I269086,);
DFFARX1 I_15617 (I269086,I3563,I269060,I269103,);
not I_15618 (I269052,I269103);
not I_15619 (I269125,I269086);
DFFARX1 I_15620 (I673450,I3563,I269060,I269151,);
not I_15621 (I269159,I269151);
and I_15622 (I269176,I269125,I673456);
not I_15623 (I269193,I673441);
nand I_15624 (I269210,I269193,I673456);
not I_15625 (I269227,I673444);
nor I_15626 (I269244,I269227,I673465);
nand I_15627 (I269261,I269244,I673462);
nor I_15628 (I269278,I269261,I269210);
DFFARX1 I_15629 (I269278,I3563,I269060,I269028,);
not I_15630 (I269309,I269261);
not I_15631 (I269326,I673465);
nand I_15632 (I269343,I269326,I673456);
nor I_15633 (I269360,I673465,I673441);
nand I_15634 (I269040,I269176,I269360);
nand I_15635 (I269034,I269125,I673465);
nand I_15636 (I269405,I269227,I673441);
DFFARX1 I_15637 (I269405,I3563,I269060,I269049,);
DFFARX1 I_15638 (I269405,I3563,I269060,I269043,);
not I_15639 (I269450,I673441);
nor I_15640 (I269467,I269450,I673447);
and I_15641 (I269484,I269467,I673459);
or I_15642 (I269501,I269484,I673444);
DFFARX1 I_15643 (I269501,I3563,I269060,I269527,);
nand I_15644 (I269535,I269527,I269193);
nor I_15645 (I269037,I269535,I269343);
nor I_15646 (I269031,I269527,I269159);
DFFARX1 I_15647 (I269527,I3563,I269060,I269589,);
not I_15648 (I269597,I269589);
nor I_15649 (I269046,I269597,I269309);
not I_15650 (I269655,I3570);
DFFARX1 I_15651 (I411845,I3563,I269655,I269681,);
DFFARX1 I_15652 (I269681,I3563,I269655,I269698,);
not I_15653 (I269647,I269698);
not I_15654 (I269720,I269681);
DFFARX1 I_15655 (I411860,I3563,I269655,I269746,);
not I_15656 (I269754,I269746);
and I_15657 (I269771,I269720,I411857);
not I_15658 (I269788,I411845);
nand I_15659 (I269805,I269788,I411857);
not I_15660 (I269822,I411854);
nor I_15661 (I269839,I269822,I411869);
nand I_15662 (I269856,I269839,I411866);
nor I_15663 (I269873,I269856,I269805);
DFFARX1 I_15664 (I269873,I3563,I269655,I269623,);
not I_15665 (I269904,I269856);
not I_15666 (I269921,I411869);
nand I_15667 (I269938,I269921,I411857);
nor I_15668 (I269955,I411869,I411845);
nand I_15669 (I269635,I269771,I269955);
nand I_15670 (I269629,I269720,I411869);
nand I_15671 (I270000,I269822,I411863);
DFFARX1 I_15672 (I270000,I3563,I269655,I269644,);
DFFARX1 I_15673 (I270000,I3563,I269655,I269638,);
not I_15674 (I270045,I411863);
nor I_15675 (I270062,I270045,I411851);
and I_15676 (I270079,I270062,I411872);
or I_15677 (I270096,I270079,I411848);
DFFARX1 I_15678 (I270096,I3563,I269655,I270122,);
nand I_15679 (I270130,I270122,I269788);
nor I_15680 (I269632,I270130,I269938);
nor I_15681 (I269626,I270122,I269754);
DFFARX1 I_15682 (I270122,I3563,I269655,I270184,);
not I_15683 (I270192,I270184);
nor I_15684 (I269641,I270192,I269904);
not I_15685 (I270250,I3570);
DFFARX1 I_15686 (I140449,I3563,I270250,I270276,);
DFFARX1 I_15687 (I270276,I3563,I270250,I270293,);
not I_15688 (I270242,I270293);
not I_15689 (I270315,I270276);
DFFARX1 I_15690 (I140443,I3563,I270250,I270341,);
not I_15691 (I270349,I270341);
and I_15692 (I270366,I270315,I140440);
not I_15693 (I270383,I140461);
nand I_15694 (I270400,I270383,I140440);
not I_15695 (I270417,I140455);
nor I_15696 (I270434,I270417,I140446);
nand I_15697 (I270451,I270434,I140452);
nor I_15698 (I270468,I270451,I270400);
DFFARX1 I_15699 (I270468,I3563,I270250,I270218,);
not I_15700 (I270499,I270451);
not I_15701 (I270516,I140446);
nand I_15702 (I270533,I270516,I140440);
nor I_15703 (I270550,I140446,I140461);
nand I_15704 (I270230,I270366,I270550);
nand I_15705 (I270224,I270315,I140446);
nand I_15706 (I270595,I270417,I140440);
DFFARX1 I_15707 (I270595,I3563,I270250,I270239,);
DFFARX1 I_15708 (I270595,I3563,I270250,I270233,);
not I_15709 (I270640,I140440);
nor I_15710 (I270657,I270640,I140458);
and I_15711 (I270674,I270657,I140464);
or I_15712 (I270691,I270674,I140443);
DFFARX1 I_15713 (I270691,I3563,I270250,I270717,);
nand I_15714 (I270725,I270717,I270383);
nor I_15715 (I270227,I270725,I270533);
nor I_15716 (I270221,I270717,I270349);
DFFARX1 I_15717 (I270717,I3563,I270250,I270779,);
not I_15718 (I270787,I270779);
nor I_15719 (I270236,I270787,I270499);
not I_15720 (I270845,I3570);
DFFARX1 I_15721 (I341227,I3563,I270845,I270871,);
DFFARX1 I_15722 (I270871,I3563,I270845,I270888,);
not I_15723 (I270837,I270888);
not I_15724 (I270910,I270871);
DFFARX1 I_15725 (I341242,I3563,I270845,I270936,);
not I_15726 (I270944,I270936);
and I_15727 (I270961,I270910,I341239);
not I_15728 (I270978,I341227);
nand I_15729 (I270995,I270978,I341239);
not I_15730 (I271012,I341236);
nor I_15731 (I271029,I271012,I341251);
nand I_15732 (I271046,I271029,I341248);
nor I_15733 (I271063,I271046,I270995);
DFFARX1 I_15734 (I271063,I3563,I270845,I270813,);
not I_15735 (I271094,I271046);
not I_15736 (I271111,I341251);
nand I_15737 (I271128,I271111,I341239);
nor I_15738 (I271145,I341251,I341227);
nand I_15739 (I270825,I270961,I271145);
nand I_15740 (I270819,I270910,I341251);
nand I_15741 (I271190,I271012,I341245);
DFFARX1 I_15742 (I271190,I3563,I270845,I270834,);
DFFARX1 I_15743 (I271190,I3563,I270845,I270828,);
not I_15744 (I271235,I341245);
nor I_15745 (I271252,I271235,I341233);
and I_15746 (I271269,I271252,I341254);
or I_15747 (I271286,I271269,I341230);
DFFARX1 I_15748 (I271286,I3563,I270845,I271312,);
nand I_15749 (I271320,I271312,I270978);
nor I_15750 (I270822,I271320,I271128);
nor I_15751 (I270816,I271312,I270944);
DFFARX1 I_15752 (I271312,I3563,I270845,I271374,);
not I_15753 (I271382,I271374);
nor I_15754 (I270831,I271382,I271094);
not I_15755 (I271440,I3570);
DFFARX1 I_15756 (I1143015,I3563,I271440,I271466,);
DFFARX1 I_15757 (I271466,I3563,I271440,I271483,);
not I_15758 (I271432,I271483);
not I_15759 (I271505,I271466);
DFFARX1 I_15760 (I1143015,I3563,I271440,I271531,);
not I_15761 (I271539,I271531);
and I_15762 (I271556,I271505,I1143018);
not I_15763 (I271573,I1143030);
nand I_15764 (I271590,I271573,I1143018);
not I_15765 (I271607,I1143036);
nor I_15766 (I271624,I271607,I1143027);
nand I_15767 (I271641,I271624,I1143033);
nor I_15768 (I271658,I271641,I271590);
DFFARX1 I_15769 (I271658,I3563,I271440,I271408,);
not I_15770 (I271689,I271641);
not I_15771 (I271706,I1143027);
nand I_15772 (I271723,I271706,I1143018);
nor I_15773 (I271740,I1143027,I1143030);
nand I_15774 (I271420,I271556,I271740);
nand I_15775 (I271414,I271505,I1143027);
nand I_15776 (I271785,I271607,I1143024);
DFFARX1 I_15777 (I271785,I3563,I271440,I271429,);
DFFARX1 I_15778 (I271785,I3563,I271440,I271423,);
not I_15779 (I271830,I1143024);
nor I_15780 (I271847,I271830,I1143021);
and I_15781 (I271864,I271847,I1143039);
or I_15782 (I271881,I271864,I1143018);
DFFARX1 I_15783 (I271881,I3563,I271440,I271907,);
nand I_15784 (I271915,I271907,I271573);
nor I_15785 (I271417,I271915,I271723);
nor I_15786 (I271411,I271907,I271539);
DFFARX1 I_15787 (I271907,I3563,I271440,I271969,);
not I_15788 (I271977,I271969);
nor I_15789 (I271426,I271977,I271689);
not I_15790 (I272035,I3570);
DFFARX1 I_15791 (I741079,I3563,I272035,I272061,);
DFFARX1 I_15792 (I272061,I3563,I272035,I272078,);
not I_15793 (I272027,I272078);
not I_15794 (I272100,I272061);
DFFARX1 I_15795 (I741076,I3563,I272035,I272126,);
not I_15796 (I272134,I272126);
and I_15797 (I272151,I272100,I741082);
not I_15798 (I272168,I741067);
nand I_15799 (I272185,I272168,I741082);
not I_15800 (I272202,I741070);
nor I_15801 (I272219,I272202,I741091);
nand I_15802 (I272236,I272219,I741088);
nor I_15803 (I272253,I272236,I272185);
DFFARX1 I_15804 (I272253,I3563,I272035,I272003,);
not I_15805 (I272284,I272236);
not I_15806 (I272301,I741091);
nand I_15807 (I272318,I272301,I741082);
nor I_15808 (I272335,I741091,I741067);
nand I_15809 (I272015,I272151,I272335);
nand I_15810 (I272009,I272100,I741091);
nand I_15811 (I272380,I272202,I741067);
DFFARX1 I_15812 (I272380,I3563,I272035,I272024,);
DFFARX1 I_15813 (I272380,I3563,I272035,I272018,);
not I_15814 (I272425,I741067);
nor I_15815 (I272442,I272425,I741073);
and I_15816 (I272459,I272442,I741085);
or I_15817 (I272476,I272459,I741070);
DFFARX1 I_15818 (I272476,I3563,I272035,I272502,);
nand I_15819 (I272510,I272502,I272168);
nor I_15820 (I272012,I272510,I272318);
nor I_15821 (I272006,I272502,I272134);
DFFARX1 I_15822 (I272502,I3563,I272035,I272564,);
not I_15823 (I272572,I272564);
nor I_15824 (I272021,I272572,I272284);
not I_15825 (I272630,I3570);
DFFARX1 I_15826 (I987242,I3563,I272630,I272656,);
DFFARX1 I_15827 (I272656,I3563,I272630,I272673,);
not I_15828 (I272622,I272673);
not I_15829 (I272695,I272656);
DFFARX1 I_15830 (I987251,I3563,I272630,I272721,);
not I_15831 (I272729,I272721);
and I_15832 (I272746,I272695,I987239);
not I_15833 (I272763,I987230);
nand I_15834 (I272780,I272763,I987239);
not I_15835 (I272797,I987236);
nor I_15836 (I272814,I272797,I987254);
nand I_15837 (I272831,I272814,I987227);
nor I_15838 (I272848,I272831,I272780);
DFFARX1 I_15839 (I272848,I3563,I272630,I272598,);
not I_15840 (I272879,I272831);
not I_15841 (I272896,I987254);
nand I_15842 (I272913,I272896,I987239);
nor I_15843 (I272930,I987254,I987230);
nand I_15844 (I272610,I272746,I272930);
nand I_15845 (I272604,I272695,I987254);
nand I_15846 (I272975,I272797,I987233);
DFFARX1 I_15847 (I272975,I3563,I272630,I272619,);
DFFARX1 I_15848 (I272975,I3563,I272630,I272613,);
not I_15849 (I273020,I987233);
nor I_15850 (I273037,I273020,I987245);
and I_15851 (I273054,I273037,I987227);
or I_15852 (I273071,I273054,I987248);
DFFARX1 I_15853 (I273071,I3563,I272630,I273097,);
nand I_15854 (I273105,I273097,I272763);
nor I_15855 (I272607,I273105,I272913);
nor I_15856 (I272601,I273097,I272729);
DFFARX1 I_15857 (I273097,I3563,I272630,I273159,);
not I_15858 (I273167,I273159);
nor I_15859 (I272616,I273167,I272879);
not I_15860 (I273225,I3570);
DFFARX1 I_15861 (I455066,I3563,I273225,I273251,);
DFFARX1 I_15862 (I273251,I3563,I273225,I273268,);
not I_15863 (I273217,I273268);
not I_15864 (I273290,I273251);
DFFARX1 I_15865 (I455054,I3563,I273225,I273316,);
not I_15866 (I273324,I273316);
and I_15867 (I273341,I273290,I455063);
not I_15868 (I273358,I455060);
nand I_15869 (I273375,I273358,I455063);
not I_15870 (I273392,I455051);
nor I_15871 (I273409,I273392,I455057);
nand I_15872 (I273426,I273409,I455042);
nor I_15873 (I273443,I273426,I273375);
DFFARX1 I_15874 (I273443,I3563,I273225,I273193,);
not I_15875 (I273474,I273426);
not I_15876 (I273491,I455057);
nand I_15877 (I273508,I273491,I455063);
nor I_15878 (I273525,I455057,I455060);
nand I_15879 (I273205,I273341,I273525);
nand I_15880 (I273199,I273290,I455057);
nand I_15881 (I273570,I273392,I455042);
DFFARX1 I_15882 (I273570,I3563,I273225,I273214,);
DFFARX1 I_15883 (I273570,I3563,I273225,I273208,);
not I_15884 (I273615,I455042);
nor I_15885 (I273632,I273615,I455048);
and I_15886 (I273649,I273632,I455045);
or I_15887 (I273666,I273649,I455069);
DFFARX1 I_15888 (I273666,I3563,I273225,I273692,);
nand I_15889 (I273700,I273692,I273358);
nor I_15890 (I273202,I273700,I273508);
nor I_15891 (I273196,I273692,I273324);
DFFARX1 I_15892 (I273692,I3563,I273225,I273754,);
not I_15893 (I273762,I273754);
nor I_15894 (I273211,I273762,I273474);
not I_15895 (I273820,I3570);
DFFARX1 I_15896 (I388657,I3563,I273820,I273846,);
DFFARX1 I_15897 (I273846,I3563,I273820,I273863,);
not I_15898 (I273812,I273863);
not I_15899 (I273885,I273846);
DFFARX1 I_15900 (I388672,I3563,I273820,I273911,);
not I_15901 (I273919,I273911);
and I_15902 (I273936,I273885,I388669);
not I_15903 (I273953,I388657);
nand I_15904 (I273970,I273953,I388669);
not I_15905 (I273987,I388666);
nor I_15906 (I274004,I273987,I388681);
nand I_15907 (I274021,I274004,I388678);
nor I_15908 (I274038,I274021,I273970);
DFFARX1 I_15909 (I274038,I3563,I273820,I273788,);
not I_15910 (I274069,I274021);
not I_15911 (I274086,I388681);
nand I_15912 (I274103,I274086,I388669);
nor I_15913 (I274120,I388681,I388657);
nand I_15914 (I273800,I273936,I274120);
nand I_15915 (I273794,I273885,I388681);
nand I_15916 (I274165,I273987,I388675);
DFFARX1 I_15917 (I274165,I3563,I273820,I273809,);
DFFARX1 I_15918 (I274165,I3563,I273820,I273803,);
not I_15919 (I274210,I388675);
nor I_15920 (I274227,I274210,I388663);
and I_15921 (I274244,I274227,I388684);
or I_15922 (I274261,I274244,I388660);
DFFARX1 I_15923 (I274261,I3563,I273820,I274287,);
nand I_15924 (I274295,I274287,I273953);
nor I_15925 (I273797,I274295,I274103);
nor I_15926 (I273791,I274287,I273919);
DFFARX1 I_15927 (I274287,I3563,I273820,I274349,);
not I_15928 (I274357,I274349);
nor I_15929 (I273806,I274357,I274069);
not I_15930 (I274415,I3570);
DFFARX1 I_15931 (I1175383,I3563,I274415,I274441,);
DFFARX1 I_15932 (I274441,I3563,I274415,I274458,);
not I_15933 (I274407,I274458);
not I_15934 (I274480,I274441);
DFFARX1 I_15935 (I1175383,I3563,I274415,I274506,);
not I_15936 (I274514,I274506);
and I_15937 (I274531,I274480,I1175386);
not I_15938 (I274548,I1175398);
nand I_15939 (I274565,I274548,I1175386);
not I_15940 (I274582,I1175404);
nor I_15941 (I274599,I274582,I1175395);
nand I_15942 (I274616,I274599,I1175401);
nor I_15943 (I274633,I274616,I274565);
DFFARX1 I_15944 (I274633,I3563,I274415,I274383,);
not I_15945 (I274664,I274616);
not I_15946 (I274681,I1175395);
nand I_15947 (I274698,I274681,I1175386);
nor I_15948 (I274715,I1175395,I1175398);
nand I_15949 (I274395,I274531,I274715);
nand I_15950 (I274389,I274480,I1175395);
nand I_15951 (I274760,I274582,I1175392);
DFFARX1 I_15952 (I274760,I3563,I274415,I274404,);
DFFARX1 I_15953 (I274760,I3563,I274415,I274398,);
not I_15954 (I274805,I1175392);
nor I_15955 (I274822,I274805,I1175389);
and I_15956 (I274839,I274822,I1175407);
or I_15957 (I274856,I274839,I1175386);
DFFARX1 I_15958 (I274856,I3563,I274415,I274882,);
nand I_15959 (I274890,I274882,I274548);
nor I_15960 (I274392,I274890,I274698);
nor I_15961 (I274386,I274882,I274514);
DFFARX1 I_15962 (I274882,I3563,I274415,I274944,);
not I_15963 (I274952,I274944);
nor I_15964 (I274401,I274952,I274664);
not I_15965 (I275010,I3570);
DFFARX1 I_15966 (I3540,I3563,I275010,I275036,);
DFFARX1 I_15967 (I275036,I3563,I275010,I275053,);
not I_15968 (I275002,I275053);
not I_15969 (I275075,I275036);
DFFARX1 I_15970 (I2500,I3563,I275010,I275101,);
not I_15971 (I275109,I275101);
and I_15972 (I275126,I275075,I1732);
not I_15973 (I275143,I1404);
nand I_15974 (I275160,I275143,I1732);
not I_15975 (I275177,I2764);
nor I_15976 (I275194,I275177,I1588);
nand I_15977 (I275211,I275194,I1500);
nor I_15978 (I275228,I275211,I275160);
DFFARX1 I_15979 (I275228,I3563,I275010,I274978,);
not I_15980 (I275259,I275211);
not I_15981 (I275276,I1588);
nand I_15982 (I275293,I275276,I1732);
nor I_15983 (I275310,I1588,I1404);
nand I_15984 (I274990,I275126,I275310);
nand I_15985 (I274984,I275075,I1588);
nand I_15986 (I275355,I275177,I2804);
DFFARX1 I_15987 (I275355,I3563,I275010,I274999,);
DFFARX1 I_15988 (I275355,I3563,I275010,I274993,);
not I_15989 (I275400,I2804);
nor I_15990 (I275417,I275400,I3372);
and I_15991 (I275434,I275417,I1812);
or I_15992 (I275451,I275434,I1604);
DFFARX1 I_15993 (I275451,I3563,I275010,I275477,);
nand I_15994 (I275485,I275477,I275143);
nor I_15995 (I274987,I275485,I275293);
nor I_15996 (I274981,I275477,I275109);
DFFARX1 I_15997 (I275477,I3563,I275010,I275539,);
not I_15998 (I275547,I275539);
nor I_15999 (I274996,I275547,I275259);
not I_16000 (I275605,I3570);
DFFARX1 I_16001 (I88803,I3563,I275605,I275631,);
DFFARX1 I_16002 (I275631,I3563,I275605,I275648,);
not I_16003 (I275597,I275648);
not I_16004 (I275670,I275631);
DFFARX1 I_16005 (I88797,I3563,I275605,I275696,);
not I_16006 (I275704,I275696);
and I_16007 (I275721,I275670,I88794);
not I_16008 (I275738,I88815);
nand I_16009 (I275755,I275738,I88794);
not I_16010 (I275772,I88809);
nor I_16011 (I275789,I275772,I88800);
nand I_16012 (I275806,I275789,I88806);
nor I_16013 (I275823,I275806,I275755);
DFFARX1 I_16014 (I275823,I3563,I275605,I275573,);
not I_16015 (I275854,I275806);
not I_16016 (I275871,I88800);
nand I_16017 (I275888,I275871,I88794);
nor I_16018 (I275905,I88800,I88815);
nand I_16019 (I275585,I275721,I275905);
nand I_16020 (I275579,I275670,I88800);
nand I_16021 (I275950,I275772,I88794);
DFFARX1 I_16022 (I275950,I3563,I275605,I275594,);
DFFARX1 I_16023 (I275950,I3563,I275605,I275588,);
not I_16024 (I275995,I88794);
nor I_16025 (I276012,I275995,I88812);
and I_16026 (I276029,I276012,I88818);
or I_16027 (I276046,I276029,I88797);
DFFARX1 I_16028 (I276046,I3563,I275605,I276072,);
nand I_16029 (I276080,I276072,I275738);
nor I_16030 (I275582,I276080,I275888);
nor I_16031 (I275576,I276072,I275704);
DFFARX1 I_16032 (I276072,I3563,I275605,I276134,);
not I_16033 (I276142,I276134);
nor I_16034 (I275591,I276142,I275854);
not I_16035 (I276200,I3570);
DFFARX1 I_16036 (I629528,I3563,I276200,I276226,);
DFFARX1 I_16037 (I276226,I3563,I276200,I276243,);
not I_16038 (I276192,I276243);
not I_16039 (I276265,I276226);
DFFARX1 I_16040 (I629519,I3563,I276200,I276291,);
not I_16041 (I276299,I276291);
and I_16042 (I276316,I276265,I629537);
not I_16043 (I276333,I629534);
nand I_16044 (I276350,I276333,I629537);
not I_16045 (I276367,I629513);
nor I_16046 (I276384,I276367,I629516);
nand I_16047 (I276401,I276384,I629525);
nor I_16048 (I276418,I276401,I276350);
DFFARX1 I_16049 (I276418,I3563,I276200,I276168,);
not I_16050 (I276449,I276401);
not I_16051 (I276466,I629516);
nand I_16052 (I276483,I276466,I629537);
nor I_16053 (I276500,I629516,I629534);
nand I_16054 (I276180,I276316,I276500);
nand I_16055 (I276174,I276265,I629516);
nand I_16056 (I276545,I276367,I629531);
DFFARX1 I_16057 (I276545,I3563,I276200,I276189,);
DFFARX1 I_16058 (I276545,I3563,I276200,I276183,);
not I_16059 (I276590,I629531);
nor I_16060 (I276607,I276590,I629513);
and I_16061 (I276624,I276607,I629522);
or I_16062 (I276641,I276624,I629516);
DFFARX1 I_16063 (I276641,I3563,I276200,I276667,);
nand I_16064 (I276675,I276667,I276333);
nor I_16065 (I276177,I276675,I276483);
nor I_16066 (I276171,I276667,I276299);
DFFARX1 I_16067 (I276667,I3563,I276200,I276729,);
not I_16068 (I276737,I276729);
nor I_16069 (I276186,I276737,I276449);
not I_16070 (I276795,I3570);
DFFARX1 I_16071 (I505658,I3563,I276795,I276821,);
DFFARX1 I_16072 (I276821,I3563,I276795,I276838,);
not I_16073 (I276787,I276838);
not I_16074 (I276860,I276821);
DFFARX1 I_16075 (I505646,I3563,I276795,I276886,);
not I_16076 (I276894,I276886);
and I_16077 (I276911,I276860,I505655);
not I_16078 (I276928,I505652);
nand I_16079 (I276945,I276928,I505655);
not I_16080 (I276962,I505643);
nor I_16081 (I276979,I276962,I505649);
nand I_16082 (I276996,I276979,I505634);
nor I_16083 (I277013,I276996,I276945);
DFFARX1 I_16084 (I277013,I3563,I276795,I276763,);
not I_16085 (I277044,I276996);
not I_16086 (I277061,I505649);
nand I_16087 (I277078,I277061,I505655);
nor I_16088 (I277095,I505649,I505652);
nand I_16089 (I276775,I276911,I277095);
nand I_16090 (I276769,I276860,I505649);
nand I_16091 (I277140,I276962,I505634);
DFFARX1 I_16092 (I277140,I3563,I276795,I276784,);
DFFARX1 I_16093 (I277140,I3563,I276795,I276778,);
not I_16094 (I277185,I505634);
nor I_16095 (I277202,I277185,I505640);
and I_16096 (I277219,I277202,I505637);
or I_16097 (I277236,I277219,I505661);
DFFARX1 I_16098 (I277236,I3563,I276795,I277262,);
nand I_16099 (I277270,I277262,I276928);
nor I_16100 (I276772,I277270,I277078);
nor I_16101 (I276766,I277262,I276894);
DFFARX1 I_16102 (I277262,I3563,I276795,I277324,);
not I_16103 (I277332,I277324);
nor I_16104 (I276781,I277332,I277044);
not I_16105 (I277390,I3570);
DFFARX1 I_16106 (I1242431,I3563,I277390,I277416,);
DFFARX1 I_16107 (I277416,I3563,I277390,I277433,);
not I_16108 (I277382,I277433);
not I_16109 (I277455,I277416);
DFFARX1 I_16110 (I1242431,I3563,I277390,I277481,);
not I_16111 (I277489,I277481);
and I_16112 (I277506,I277455,I1242434);
not I_16113 (I277523,I1242446);
nand I_16114 (I277540,I277523,I1242434);
not I_16115 (I277557,I1242452);
nor I_16116 (I277574,I277557,I1242443);
nand I_16117 (I277591,I277574,I1242449);
nor I_16118 (I277608,I277591,I277540);
DFFARX1 I_16119 (I277608,I3563,I277390,I277358,);
not I_16120 (I277639,I277591);
not I_16121 (I277656,I1242443);
nand I_16122 (I277673,I277656,I1242434);
nor I_16123 (I277690,I1242443,I1242446);
nand I_16124 (I277370,I277506,I277690);
nand I_16125 (I277364,I277455,I1242443);
nand I_16126 (I277735,I277557,I1242440);
DFFARX1 I_16127 (I277735,I3563,I277390,I277379,);
DFFARX1 I_16128 (I277735,I3563,I277390,I277373,);
not I_16129 (I277780,I1242440);
nor I_16130 (I277797,I277780,I1242437);
and I_16131 (I277814,I277797,I1242455);
or I_16132 (I277831,I277814,I1242434);
DFFARX1 I_16133 (I277831,I3563,I277390,I277857,);
nand I_16134 (I277865,I277857,I277523);
nor I_16135 (I277367,I277865,I277673);
nor I_16136 (I277361,I277857,I277489);
DFFARX1 I_16137 (I277857,I3563,I277390,I277919,);
not I_16138 (I277927,I277919);
nor I_16139 (I277376,I277927,I277639);
not I_16140 (I277985,I3570);
DFFARX1 I_16141 (I587334,I3563,I277985,I278011,);
DFFARX1 I_16142 (I278011,I3563,I277985,I278028,);
not I_16143 (I277977,I278028);
not I_16144 (I278050,I278011);
DFFARX1 I_16145 (I587325,I3563,I277985,I278076,);
not I_16146 (I278084,I278076);
and I_16147 (I278101,I278050,I587343);
not I_16148 (I278118,I587340);
nand I_16149 (I278135,I278118,I587343);
not I_16150 (I278152,I587319);
nor I_16151 (I278169,I278152,I587322);
nand I_16152 (I278186,I278169,I587331);
nor I_16153 (I278203,I278186,I278135);
DFFARX1 I_16154 (I278203,I3563,I277985,I277953,);
not I_16155 (I278234,I278186);
not I_16156 (I278251,I587322);
nand I_16157 (I278268,I278251,I587343);
nor I_16158 (I278285,I587322,I587340);
nand I_16159 (I277965,I278101,I278285);
nand I_16160 (I277959,I278050,I587322);
nand I_16161 (I278330,I278152,I587337);
DFFARX1 I_16162 (I278330,I3563,I277985,I277974,);
DFFARX1 I_16163 (I278330,I3563,I277985,I277968,);
not I_16164 (I278375,I587337);
nor I_16165 (I278392,I278375,I587319);
and I_16166 (I278409,I278392,I587328);
or I_16167 (I278426,I278409,I587322);
DFFARX1 I_16168 (I278426,I3563,I277985,I278452,);
nand I_16169 (I278460,I278452,I278118);
nor I_16170 (I277962,I278460,I278268);
nor I_16171 (I277956,I278452,I278084);
DFFARX1 I_16172 (I278452,I3563,I277985,I278514,);
not I_16173 (I278522,I278514);
nor I_16174 (I277971,I278522,I278234);
not I_16175 (I278580,I3570);
DFFARX1 I_16176 (I1275803,I3563,I278580,I278606,);
DFFARX1 I_16177 (I278606,I3563,I278580,I278623,);
not I_16178 (I278572,I278623);
not I_16179 (I278645,I278606);
DFFARX1 I_16180 (I1275788,I3563,I278580,I278671,);
not I_16181 (I278679,I278671);
and I_16182 (I278696,I278645,I1275806);
not I_16183 (I278713,I1275788);
nand I_16184 (I278730,I278713,I1275806);
not I_16185 (I278747,I1275809);
nor I_16186 (I278764,I278747,I1275800);
nand I_16187 (I278781,I278764,I1275797);
nor I_16188 (I278798,I278781,I278730);
DFFARX1 I_16189 (I278798,I3563,I278580,I278548,);
not I_16190 (I278829,I278781);
not I_16191 (I278846,I1275800);
nand I_16192 (I278863,I278846,I1275806);
nor I_16193 (I278880,I1275800,I1275788);
nand I_16194 (I278560,I278696,I278880);
nand I_16195 (I278554,I278645,I1275800);
nand I_16196 (I278925,I278747,I1275794);
DFFARX1 I_16197 (I278925,I3563,I278580,I278569,);
DFFARX1 I_16198 (I278925,I3563,I278580,I278563,);
not I_16199 (I278970,I1275794);
nor I_16200 (I278987,I278970,I1275785);
and I_16201 (I279004,I278987,I1275791);
or I_16202 (I279021,I279004,I1275785);
DFFARX1 I_16203 (I279021,I3563,I278580,I279047,);
nand I_16204 (I279055,I279047,I278713);
nor I_16205 (I278557,I279055,I278863);
nor I_16206 (I278551,I279047,I278679);
DFFARX1 I_16207 (I279047,I3563,I278580,I279109,);
not I_16208 (I279117,I279109);
nor I_16209 (I278566,I279117,I278829);
not I_16210 (I279175,I3570);
DFFARX1 I_16211 (I490970,I3563,I279175,I279201,);
DFFARX1 I_16212 (I279201,I3563,I279175,I279218,);
not I_16213 (I279167,I279218);
not I_16214 (I279240,I279201);
DFFARX1 I_16215 (I490958,I3563,I279175,I279266,);
not I_16216 (I279274,I279266);
and I_16217 (I279291,I279240,I490967);
not I_16218 (I279308,I490964);
nand I_16219 (I279325,I279308,I490967);
not I_16220 (I279342,I490955);
nor I_16221 (I279359,I279342,I490961);
nand I_16222 (I279376,I279359,I490946);
nor I_16223 (I279393,I279376,I279325);
DFFARX1 I_16224 (I279393,I3563,I279175,I279143,);
not I_16225 (I279424,I279376);
not I_16226 (I279441,I490961);
nand I_16227 (I279458,I279441,I490967);
nor I_16228 (I279475,I490961,I490964);
nand I_16229 (I279155,I279291,I279475);
nand I_16230 (I279149,I279240,I490961);
nand I_16231 (I279520,I279342,I490946);
DFFARX1 I_16232 (I279520,I3563,I279175,I279164,);
DFFARX1 I_16233 (I279520,I3563,I279175,I279158,);
not I_16234 (I279565,I490946);
nor I_16235 (I279582,I279565,I490952);
and I_16236 (I279599,I279582,I490949);
or I_16237 (I279616,I279599,I490973);
DFFARX1 I_16238 (I279616,I3563,I279175,I279642,);
nand I_16239 (I279650,I279642,I279308);
nor I_16240 (I279152,I279650,I279458);
nor I_16241 (I279146,I279642,I279274);
DFFARX1 I_16242 (I279642,I3563,I279175,I279704,);
not I_16243 (I279712,I279704);
nor I_16244 (I279161,I279712,I279424);
not I_16245 (I279770,I3570);
DFFARX1 I_16246 (I620858,I3563,I279770,I279796,);
DFFARX1 I_16247 (I279796,I3563,I279770,I279813,);
not I_16248 (I279762,I279813);
not I_16249 (I279835,I279796);
DFFARX1 I_16250 (I620849,I3563,I279770,I279861,);
not I_16251 (I279869,I279861);
and I_16252 (I279886,I279835,I620867);
not I_16253 (I279903,I620864);
nand I_16254 (I279920,I279903,I620867);
not I_16255 (I279937,I620843);
nor I_16256 (I279954,I279937,I620846);
nand I_16257 (I279971,I279954,I620855);
nor I_16258 (I279988,I279971,I279920);
DFFARX1 I_16259 (I279988,I3563,I279770,I279738,);
not I_16260 (I280019,I279971);
not I_16261 (I280036,I620846);
nand I_16262 (I280053,I280036,I620867);
nor I_16263 (I280070,I620846,I620864);
nand I_16264 (I279750,I279886,I280070);
nand I_16265 (I279744,I279835,I620846);
nand I_16266 (I280115,I279937,I620861);
DFFARX1 I_16267 (I280115,I3563,I279770,I279759,);
DFFARX1 I_16268 (I280115,I3563,I279770,I279753,);
not I_16269 (I280160,I620861);
nor I_16270 (I280177,I280160,I620843);
and I_16271 (I280194,I280177,I620852);
or I_16272 (I280211,I280194,I620846);
DFFARX1 I_16273 (I280211,I3563,I279770,I280237,);
nand I_16274 (I280245,I280237,I279903);
nor I_16275 (I279747,I280245,I280053);
nor I_16276 (I279741,I280237,I279869);
DFFARX1 I_16277 (I280237,I3563,I279770,I280299,);
not I_16278 (I280307,I280299);
nor I_16279 (I279756,I280307,I280019);
not I_16280 (I280365,I3570);
DFFARX1 I_16281 (I478458,I3563,I280365,I280391,);
DFFARX1 I_16282 (I280391,I3563,I280365,I280408,);
not I_16283 (I280357,I280408);
not I_16284 (I280430,I280391);
DFFARX1 I_16285 (I478446,I3563,I280365,I280456,);
not I_16286 (I280464,I280456);
and I_16287 (I280481,I280430,I478455);
not I_16288 (I280498,I478452);
nand I_16289 (I280515,I280498,I478455);
not I_16290 (I280532,I478443);
nor I_16291 (I280549,I280532,I478449);
nand I_16292 (I280566,I280549,I478434);
nor I_16293 (I280583,I280566,I280515);
DFFARX1 I_16294 (I280583,I3563,I280365,I280333,);
not I_16295 (I280614,I280566);
not I_16296 (I280631,I478449);
nand I_16297 (I280648,I280631,I478455);
nor I_16298 (I280665,I478449,I478452);
nand I_16299 (I280345,I280481,I280665);
nand I_16300 (I280339,I280430,I478449);
nand I_16301 (I280710,I280532,I478434);
DFFARX1 I_16302 (I280710,I3563,I280365,I280354,);
DFFARX1 I_16303 (I280710,I3563,I280365,I280348,);
not I_16304 (I280755,I478434);
nor I_16305 (I280772,I280755,I478440);
and I_16306 (I280789,I280772,I478437);
or I_16307 (I280806,I280789,I478461);
DFFARX1 I_16308 (I280806,I3563,I280365,I280832,);
nand I_16309 (I280840,I280832,I280498);
nor I_16310 (I280342,I280840,I280648);
nor I_16311 (I280336,I280832,I280464);
DFFARX1 I_16312 (I280832,I3563,I280365,I280894,);
not I_16313 (I280902,I280894);
nor I_16314 (I280351,I280902,I280614);
not I_16315 (I280960,I3570);
DFFARX1 I_16316 (I513274,I3563,I280960,I280986,);
DFFARX1 I_16317 (I280986,I3563,I280960,I281003,);
not I_16318 (I280952,I281003);
not I_16319 (I281025,I280986);
DFFARX1 I_16320 (I513262,I3563,I280960,I281051,);
not I_16321 (I281059,I281051);
and I_16322 (I281076,I281025,I513271);
not I_16323 (I281093,I513268);
nand I_16324 (I281110,I281093,I513271);
not I_16325 (I281127,I513259);
nor I_16326 (I281144,I281127,I513265);
nand I_16327 (I281161,I281144,I513250);
nor I_16328 (I281178,I281161,I281110);
DFFARX1 I_16329 (I281178,I3563,I280960,I280928,);
not I_16330 (I281209,I281161);
not I_16331 (I281226,I513265);
nand I_16332 (I281243,I281226,I513271);
nor I_16333 (I281260,I513265,I513268);
nand I_16334 (I280940,I281076,I281260);
nand I_16335 (I280934,I281025,I513265);
nand I_16336 (I281305,I281127,I513250);
DFFARX1 I_16337 (I281305,I3563,I280960,I280949,);
DFFARX1 I_16338 (I281305,I3563,I280960,I280943,);
not I_16339 (I281350,I513250);
nor I_16340 (I281367,I281350,I513256);
and I_16341 (I281384,I281367,I513253);
or I_16342 (I281401,I281384,I513277);
DFFARX1 I_16343 (I281401,I3563,I280960,I281427,);
nand I_16344 (I281435,I281427,I281093);
nor I_16345 (I280937,I281435,I281243);
nor I_16346 (I280931,I281427,I281059);
DFFARX1 I_16347 (I281427,I3563,I280960,I281489,);
not I_16348 (I281497,I281489);
nor I_16349 (I280946,I281497,I281209);
not I_16350 (I281555,I3570);
DFFARX1 I_16351 (I756685,I3563,I281555,I281581,);
DFFARX1 I_16352 (I281581,I3563,I281555,I281598,);
not I_16353 (I281547,I281598);
not I_16354 (I281620,I281581);
DFFARX1 I_16355 (I756682,I3563,I281555,I281646,);
not I_16356 (I281654,I281646);
and I_16357 (I281671,I281620,I756688);
not I_16358 (I281688,I756673);
nand I_16359 (I281705,I281688,I756688);
not I_16360 (I281722,I756676);
nor I_16361 (I281739,I281722,I756697);
nand I_16362 (I281756,I281739,I756694);
nor I_16363 (I281773,I281756,I281705);
DFFARX1 I_16364 (I281773,I3563,I281555,I281523,);
not I_16365 (I281804,I281756);
not I_16366 (I281821,I756697);
nand I_16367 (I281838,I281821,I756688);
nor I_16368 (I281855,I756697,I756673);
nand I_16369 (I281535,I281671,I281855);
nand I_16370 (I281529,I281620,I756697);
nand I_16371 (I281900,I281722,I756673);
DFFARX1 I_16372 (I281900,I3563,I281555,I281544,);
DFFARX1 I_16373 (I281900,I3563,I281555,I281538,);
not I_16374 (I281945,I756673);
nor I_16375 (I281962,I281945,I756679);
and I_16376 (I281979,I281962,I756691);
or I_16377 (I281996,I281979,I756676);
DFFARX1 I_16378 (I281996,I3563,I281555,I282022,);
nand I_16379 (I282030,I282022,I281688);
nor I_16380 (I281532,I282030,I281838);
nor I_16381 (I281526,I282022,I281654);
DFFARX1 I_16382 (I282022,I3563,I281555,I282084,);
not I_16383 (I282092,I282084);
nor I_16384 (I281541,I282092,I281804);
not I_16385 (I282150,I3570);
DFFARX1 I_16386 (I1046662,I3563,I282150,I282176,);
DFFARX1 I_16387 (I282176,I3563,I282150,I282193,);
not I_16388 (I282142,I282193);
not I_16389 (I282215,I282176);
DFFARX1 I_16390 (I1046671,I3563,I282150,I282241,);
not I_16391 (I282249,I282241);
and I_16392 (I282266,I282215,I1046665);
not I_16393 (I282283,I1046659);
nand I_16394 (I282300,I282283,I1046665);
not I_16395 (I282317,I1046674);
nor I_16396 (I282334,I282317,I1046662);
nand I_16397 (I282351,I282334,I1046668);
nor I_16398 (I282368,I282351,I282300);
DFFARX1 I_16399 (I282368,I3563,I282150,I282118,);
not I_16400 (I282399,I282351);
not I_16401 (I282416,I1046662);
nand I_16402 (I282433,I282416,I1046665);
nor I_16403 (I282450,I1046662,I1046659);
nand I_16404 (I282130,I282266,I282450);
nand I_16405 (I282124,I282215,I1046662);
nand I_16406 (I282495,I282317,I1046665);
DFFARX1 I_16407 (I282495,I3563,I282150,I282139,);
DFFARX1 I_16408 (I282495,I3563,I282150,I282133,);
not I_16409 (I282540,I1046665);
nor I_16410 (I282557,I282540,I1046680);
and I_16411 (I282574,I282557,I1046677);
or I_16412 (I282591,I282574,I1046659);
DFFARX1 I_16413 (I282591,I3563,I282150,I282617,);
nand I_16414 (I282625,I282617,I282283);
nor I_16415 (I282127,I282625,I282433);
nor I_16416 (I282121,I282617,I282249);
DFFARX1 I_16417 (I282617,I3563,I282150,I282679,);
not I_16418 (I282687,I282679);
nor I_16419 (I282136,I282687,I282399);
not I_16420 (I282745,I3570);
DFFARX1 I_16421 (I121477,I3563,I282745,I282771,);
DFFARX1 I_16422 (I282771,I3563,I282745,I282788,);
not I_16423 (I282737,I282788);
not I_16424 (I282810,I282771);
DFFARX1 I_16425 (I121471,I3563,I282745,I282836,);
not I_16426 (I282844,I282836);
and I_16427 (I282861,I282810,I121468);
not I_16428 (I282878,I121489);
nand I_16429 (I282895,I282878,I121468);
not I_16430 (I282912,I121483);
nor I_16431 (I282929,I282912,I121474);
nand I_16432 (I282946,I282929,I121480);
nor I_16433 (I282963,I282946,I282895);
DFFARX1 I_16434 (I282963,I3563,I282745,I282713,);
not I_16435 (I282994,I282946);
not I_16436 (I283011,I121474);
nand I_16437 (I283028,I283011,I121468);
nor I_16438 (I283045,I121474,I121489);
nand I_16439 (I282725,I282861,I283045);
nand I_16440 (I282719,I282810,I121474);
nand I_16441 (I283090,I282912,I121468);
DFFARX1 I_16442 (I283090,I3563,I282745,I282734,);
DFFARX1 I_16443 (I283090,I3563,I282745,I282728,);
not I_16444 (I283135,I121468);
nor I_16445 (I283152,I283135,I121486);
and I_16446 (I283169,I283152,I121492);
or I_16447 (I283186,I283169,I121471);
DFFARX1 I_16448 (I283186,I3563,I282745,I283212,);
nand I_16449 (I283220,I283212,I282878);
nor I_16450 (I282722,I283220,I283028);
nor I_16451 (I282716,I283212,I282844);
DFFARX1 I_16452 (I283212,I3563,I282745,I283274,);
not I_16453 (I283282,I283274);
nor I_16454 (I282731,I283282,I282994);
not I_16455 (I283340,I3570);
DFFARX1 I_16456 (I1158043,I3563,I283340,I283366,);
DFFARX1 I_16457 (I283366,I3563,I283340,I283383,);
not I_16458 (I283332,I283383);
not I_16459 (I283405,I283366);
DFFARX1 I_16460 (I1158043,I3563,I283340,I283431,);
not I_16461 (I283439,I283431);
and I_16462 (I283456,I283405,I1158046);
not I_16463 (I283473,I1158058);
nand I_16464 (I283490,I283473,I1158046);
not I_16465 (I283507,I1158064);
nor I_16466 (I283524,I283507,I1158055);
nand I_16467 (I283541,I283524,I1158061);
nor I_16468 (I283558,I283541,I283490);
DFFARX1 I_16469 (I283558,I3563,I283340,I283308,);
not I_16470 (I283589,I283541);
not I_16471 (I283606,I1158055);
nand I_16472 (I283623,I283606,I1158046);
nor I_16473 (I283640,I1158055,I1158058);
nand I_16474 (I283320,I283456,I283640);
nand I_16475 (I283314,I283405,I1158055);
nand I_16476 (I283685,I283507,I1158052);
DFFARX1 I_16477 (I283685,I3563,I283340,I283329,);
DFFARX1 I_16478 (I283685,I3563,I283340,I283323,);
not I_16479 (I283730,I1158052);
nor I_16480 (I283747,I283730,I1158049);
and I_16481 (I283764,I283747,I1158067);
or I_16482 (I283781,I283764,I1158046);
DFFARX1 I_16483 (I283781,I3563,I283340,I283807,);
nand I_16484 (I283815,I283807,I283473);
nor I_16485 (I283317,I283815,I283623);
nor I_16486 (I283311,I283807,I283439);
DFFARX1 I_16487 (I283807,I3563,I283340,I283869,);
not I_16488 (I283877,I283869);
nor I_16489 (I283326,I283877,I283589);
not I_16490 (I283935,I3570);
DFFARX1 I_16491 (I928456,I3563,I283935,I283961,);
DFFARX1 I_16492 (I283961,I3563,I283935,I283978,);
not I_16493 (I283927,I283978);
not I_16494 (I284000,I283961);
DFFARX1 I_16495 (I928465,I3563,I283935,I284026,);
not I_16496 (I284034,I284026);
and I_16497 (I284051,I284000,I928453);
not I_16498 (I284068,I928444);
nand I_16499 (I284085,I284068,I928453);
not I_16500 (I284102,I928450);
nor I_16501 (I284119,I284102,I928468);
nand I_16502 (I284136,I284119,I928441);
nor I_16503 (I284153,I284136,I284085);
DFFARX1 I_16504 (I284153,I3563,I283935,I283903,);
not I_16505 (I284184,I284136);
not I_16506 (I284201,I928468);
nand I_16507 (I284218,I284201,I928453);
nor I_16508 (I284235,I928468,I928444);
nand I_16509 (I283915,I284051,I284235);
nand I_16510 (I283909,I284000,I928468);
nand I_16511 (I284280,I284102,I928447);
DFFARX1 I_16512 (I284280,I3563,I283935,I283924,);
DFFARX1 I_16513 (I284280,I3563,I283935,I283918,);
not I_16514 (I284325,I928447);
nor I_16515 (I284342,I284325,I928459);
and I_16516 (I284359,I284342,I928441);
or I_16517 (I284376,I284359,I928462);
DFFARX1 I_16518 (I284376,I3563,I283935,I284402,);
nand I_16519 (I284410,I284402,I284068);
nor I_16520 (I283912,I284410,I284218);
nor I_16521 (I283906,I284402,I284034);
DFFARX1 I_16522 (I284402,I3563,I283935,I284464,);
not I_16523 (I284472,I284464);
nor I_16524 (I283921,I284472,I284184);
not I_16525 (I284530,I3570);
DFFARX1 I_16526 (I921350,I3563,I284530,I284556,);
DFFARX1 I_16527 (I284556,I3563,I284530,I284573,);
not I_16528 (I284522,I284573);
not I_16529 (I284595,I284556);
DFFARX1 I_16530 (I921359,I3563,I284530,I284621,);
not I_16531 (I284629,I284621);
and I_16532 (I284646,I284595,I921347);
not I_16533 (I284663,I921338);
nand I_16534 (I284680,I284663,I921347);
not I_16535 (I284697,I921344);
nor I_16536 (I284714,I284697,I921362);
nand I_16537 (I284731,I284714,I921335);
nor I_16538 (I284748,I284731,I284680);
DFFARX1 I_16539 (I284748,I3563,I284530,I284498,);
not I_16540 (I284779,I284731);
not I_16541 (I284796,I921362);
nand I_16542 (I284813,I284796,I921347);
nor I_16543 (I284830,I921362,I921338);
nand I_16544 (I284510,I284646,I284830);
nand I_16545 (I284504,I284595,I921362);
nand I_16546 (I284875,I284697,I921341);
DFFARX1 I_16547 (I284875,I3563,I284530,I284519,);
DFFARX1 I_16548 (I284875,I3563,I284530,I284513,);
not I_16549 (I284920,I921341);
nor I_16550 (I284937,I284920,I921353);
and I_16551 (I284954,I284937,I921335);
or I_16552 (I284971,I284954,I921356);
DFFARX1 I_16553 (I284971,I3563,I284530,I284997,);
nand I_16554 (I285005,I284997,I284663);
nor I_16555 (I284507,I285005,I284813);
nor I_16556 (I284501,I284997,I284629);
DFFARX1 I_16557 (I284997,I3563,I284530,I285059,);
not I_16558 (I285067,I285059);
nor I_16559 (I284516,I285067,I284779);
not I_16560 (I285125,I3570);
DFFARX1 I_16561 (I688481,I3563,I285125,I285151,);
DFFARX1 I_16562 (I285151,I3563,I285125,I285168,);
not I_16563 (I285117,I285168);
not I_16564 (I285190,I285151);
DFFARX1 I_16565 (I688478,I3563,I285125,I285216,);
not I_16566 (I285224,I285216);
and I_16567 (I285241,I285190,I688484);
not I_16568 (I285258,I688469);
nand I_16569 (I285275,I285258,I688484);
not I_16570 (I285292,I688472);
nor I_16571 (I285309,I285292,I688493);
nand I_16572 (I285326,I285309,I688490);
nor I_16573 (I285343,I285326,I285275);
DFFARX1 I_16574 (I285343,I3563,I285125,I285093,);
not I_16575 (I285374,I285326);
not I_16576 (I285391,I688493);
nand I_16577 (I285408,I285391,I688484);
nor I_16578 (I285425,I688493,I688469);
nand I_16579 (I285105,I285241,I285425);
nand I_16580 (I285099,I285190,I688493);
nand I_16581 (I285470,I285292,I688469);
DFFARX1 I_16582 (I285470,I3563,I285125,I285114,);
DFFARX1 I_16583 (I285470,I3563,I285125,I285108,);
not I_16584 (I285515,I688469);
nor I_16585 (I285532,I285515,I688475);
and I_16586 (I285549,I285532,I688487);
or I_16587 (I285566,I285549,I688472);
DFFARX1 I_16588 (I285566,I3563,I285125,I285592,);
nand I_16589 (I285600,I285592,I285258);
nor I_16590 (I285102,I285600,I285408);
nor I_16591 (I285096,I285592,I285224);
DFFARX1 I_16592 (I285592,I3563,I285125,I285654,);
not I_16593 (I285662,I285654);
nor I_16594 (I285111,I285662,I285374);
not I_16595 (I285720,I3570);
DFFARX1 I_16596 (I913827,I3563,I285720,I285746,);
DFFARX1 I_16597 (I285746,I3563,I285720,I285763,);
not I_16598 (I285712,I285763);
not I_16599 (I285785,I285746);
DFFARX1 I_16600 (I913821,I3563,I285720,I285811,);
not I_16601 (I285819,I285811);
and I_16602 (I285836,I285785,I913839);
not I_16603 (I285853,I913827);
nand I_16604 (I285870,I285853,I913839);
not I_16605 (I285887,I913821);
nor I_16606 (I285904,I285887,I913833);
nand I_16607 (I285921,I285904,I913824);
nor I_16608 (I285938,I285921,I285870);
DFFARX1 I_16609 (I285938,I3563,I285720,I285688,);
not I_16610 (I285969,I285921);
not I_16611 (I285986,I913833);
nand I_16612 (I286003,I285986,I913839);
nor I_16613 (I286020,I913833,I913827);
nand I_16614 (I285700,I285836,I286020);
nand I_16615 (I285694,I285785,I913833);
nand I_16616 (I286065,I285887,I913836);
DFFARX1 I_16617 (I286065,I3563,I285720,I285709,);
DFFARX1 I_16618 (I286065,I3563,I285720,I285703,);
not I_16619 (I286110,I913836);
nor I_16620 (I286127,I286110,I913842);
and I_16621 (I286144,I286127,I913824);
or I_16622 (I286161,I286144,I913830);
DFFARX1 I_16623 (I286161,I3563,I285720,I286187,);
nand I_16624 (I286195,I286187,I285853);
nor I_16625 (I285697,I286195,I286003);
nor I_16626 (I285691,I286187,I285819);
DFFARX1 I_16627 (I286187,I3563,I285720,I286249,);
not I_16628 (I286257,I286249);
nor I_16629 (I285706,I286257,I285969);
not I_16630 (I286315,I3570);
DFFARX1 I_16631 (I50347,I3563,I286315,I286341,);
DFFARX1 I_16632 (I286341,I3563,I286315,I286358,);
not I_16633 (I286307,I286358);
not I_16634 (I286380,I286341);
DFFARX1 I_16635 (I50323,I3563,I286315,I286406,);
not I_16636 (I286414,I286406);
and I_16637 (I286431,I286380,I50338);
not I_16638 (I286448,I50326);
nand I_16639 (I286465,I286448,I50338);
not I_16640 (I286482,I50329);
nor I_16641 (I286499,I286482,I50341);
nand I_16642 (I286516,I286499,I50332);
nor I_16643 (I286533,I286516,I286465);
DFFARX1 I_16644 (I286533,I3563,I286315,I286283,);
not I_16645 (I286564,I286516);
not I_16646 (I286581,I50341);
nand I_16647 (I286598,I286581,I50338);
nor I_16648 (I286615,I50341,I50326);
nand I_16649 (I286295,I286431,I286615);
nand I_16650 (I286289,I286380,I50341);
nand I_16651 (I286660,I286482,I50335);
DFFARX1 I_16652 (I286660,I3563,I286315,I286304,);
DFFARX1 I_16653 (I286660,I3563,I286315,I286298,);
not I_16654 (I286705,I50335);
nor I_16655 (I286722,I286705,I50326);
and I_16656 (I286739,I286722,I50323);
or I_16657 (I286756,I286739,I50344);
DFFARX1 I_16658 (I286756,I3563,I286315,I286782,);
nand I_16659 (I286790,I286782,I286448);
nor I_16660 (I286292,I286790,I286598);
nor I_16661 (I286286,I286782,I286414);
DFFARX1 I_16662 (I286782,I3563,I286315,I286844,);
not I_16663 (I286852,I286844);
nor I_16664 (I286301,I286852,I286564);
not I_16665 (I286910,I3570);
DFFARX1 I_16666 (I1004038,I3563,I286910,I286936,);
DFFARX1 I_16667 (I286936,I3563,I286910,I286953,);
not I_16668 (I286902,I286953);
not I_16669 (I286975,I286936);
DFFARX1 I_16670 (I1004047,I3563,I286910,I287001,);
not I_16671 (I287009,I287001);
and I_16672 (I287026,I286975,I1004035);
not I_16673 (I287043,I1004026);
nand I_16674 (I287060,I287043,I1004035);
not I_16675 (I287077,I1004032);
nor I_16676 (I287094,I287077,I1004050);
nand I_16677 (I287111,I287094,I1004023);
nor I_16678 (I287128,I287111,I287060);
DFFARX1 I_16679 (I287128,I3563,I286910,I286878,);
not I_16680 (I287159,I287111);
not I_16681 (I287176,I1004050);
nand I_16682 (I287193,I287176,I1004035);
nor I_16683 (I287210,I1004050,I1004026);
nand I_16684 (I286890,I287026,I287210);
nand I_16685 (I286884,I286975,I1004050);
nand I_16686 (I287255,I287077,I1004029);
DFFARX1 I_16687 (I287255,I3563,I286910,I286899,);
DFFARX1 I_16688 (I287255,I3563,I286910,I286893,);
not I_16689 (I287300,I1004029);
nor I_16690 (I287317,I287300,I1004041);
and I_16691 (I287334,I287317,I1004023);
or I_16692 (I287351,I287334,I1004044);
DFFARX1 I_16693 (I287351,I3563,I286910,I287377,);
nand I_16694 (I287385,I287377,I287043);
nor I_16695 (I286887,I287385,I287193);
nor I_16696 (I286881,I287377,I287009);
DFFARX1 I_16697 (I287377,I3563,I286910,I287439,);
not I_16698 (I287447,I287439);
nor I_16699 (I286896,I287447,I287159);
not I_16700 (I287508,I3570);
DFFARX1 I_16701 (I541779,I3563,I287508,I287534,);
nand I_16702 (I287542,I541779,I541791);
and I_16703 (I287559,I287542,I541776);
DFFARX1 I_16704 (I287559,I3563,I287508,I287585,);
nor I_16705 (I287476,I287585,I287534);
not I_16706 (I287607,I287585);
DFFARX1 I_16707 (I541800,I3563,I287508,I287633,);
nand I_16708 (I287641,I287633,I541797);
not I_16709 (I287658,I287641);
DFFARX1 I_16710 (I287658,I3563,I287508,I287684,);
not I_16711 (I287500,I287684);
nor I_16712 (I287706,I287534,I287641);
nor I_16713 (I287482,I287585,I287706);
DFFARX1 I_16714 (I541788,I3563,I287508,I287746,);
DFFARX1 I_16715 (I287746,I3563,I287508,I287763,);
not I_16716 (I287771,I287763);
not I_16717 (I287788,I287746);
nand I_16718 (I287485,I287788,I287607);
nand I_16719 (I287819,I541776,I541785);
and I_16720 (I287836,I287819,I541794);
DFFARX1 I_16721 (I287836,I3563,I287508,I287862,);
nor I_16722 (I287870,I287862,I287534);
DFFARX1 I_16723 (I287870,I3563,I287508,I287473,);
DFFARX1 I_16724 (I287862,I3563,I287508,I287491,);
nor I_16725 (I287915,I541782,I541785);
not I_16726 (I287932,I287915);
nor I_16727 (I287494,I287771,I287932);
nand I_16728 (I287479,I287788,I287932);
nor I_16729 (I287488,I287534,I287915);
DFFARX1 I_16730 (I287915,I3563,I287508,I287497,);
not I_16731 (I288035,I3570);
DFFARX1 I_16732 (I932320,I3563,I288035,I288061,);
nand I_16733 (I288069,I932317,I932335);
and I_16734 (I288086,I288069,I932326);
DFFARX1 I_16735 (I288086,I3563,I288035,I288112,);
nor I_16736 (I288003,I288112,I288061);
not I_16737 (I288134,I288112);
DFFARX1 I_16738 (I932341,I3563,I288035,I288160,);
nand I_16739 (I288168,I288160,I932323);
not I_16740 (I288185,I288168);
DFFARX1 I_16741 (I288185,I3563,I288035,I288211,);
not I_16742 (I288027,I288211);
nor I_16743 (I288233,I288061,I288168);
nor I_16744 (I288009,I288112,I288233);
DFFARX1 I_16745 (I932329,I3563,I288035,I288273,);
DFFARX1 I_16746 (I288273,I3563,I288035,I288290,);
not I_16747 (I288298,I288290);
not I_16748 (I288315,I288273);
nand I_16749 (I288012,I288315,I288134);
nand I_16750 (I288346,I932317,I932344);
and I_16751 (I288363,I288346,I932332);
DFFARX1 I_16752 (I288363,I3563,I288035,I288389,);
nor I_16753 (I288397,I288389,I288061);
DFFARX1 I_16754 (I288397,I3563,I288035,I288000,);
DFFARX1 I_16755 (I288389,I3563,I288035,I288018,);
nor I_16756 (I288442,I932338,I932344);
not I_16757 (I288459,I288442);
nor I_16758 (I288021,I288298,I288459);
nand I_16759 (I288006,I288315,I288459);
nor I_16760 (I288015,I288061,I288442);
DFFARX1 I_16761 (I288442,I3563,I288035,I288024,);
not I_16762 (I288562,I3570);
DFFARX1 I_16763 (I1096197,I3563,I288562,I288588,);
nand I_16764 (I288596,I1096212,I1096197);
and I_16765 (I288613,I288596,I1096215);
DFFARX1 I_16766 (I288613,I3563,I288562,I288639,);
nor I_16767 (I288530,I288639,I288588);
not I_16768 (I288661,I288639);
DFFARX1 I_16769 (I1096221,I3563,I288562,I288687,);
nand I_16770 (I288695,I288687,I1096203);
not I_16771 (I288712,I288695);
DFFARX1 I_16772 (I288712,I3563,I288562,I288738,);
not I_16773 (I288554,I288738);
nor I_16774 (I288760,I288588,I288695);
nor I_16775 (I288536,I288639,I288760);
DFFARX1 I_16776 (I1096200,I3563,I288562,I288800,);
DFFARX1 I_16777 (I288800,I3563,I288562,I288817,);
not I_16778 (I288825,I288817);
not I_16779 (I288842,I288800);
nand I_16780 (I288539,I288842,I288661);
nand I_16781 (I288873,I1096200,I1096206);
and I_16782 (I288890,I288873,I1096218);
DFFARX1 I_16783 (I288890,I3563,I288562,I288916,);
nor I_16784 (I288924,I288916,I288588);
DFFARX1 I_16785 (I288924,I3563,I288562,I288527,);
DFFARX1 I_16786 (I288916,I3563,I288562,I288545,);
nor I_16787 (I288969,I1096209,I1096206);
not I_16788 (I288986,I288969);
nor I_16789 (I288548,I288825,I288986);
nand I_16790 (I288533,I288842,I288986);
nor I_16791 (I288542,I288588,I288969);
DFFARX1 I_16792 (I288969,I3563,I288562,I288551,);
not I_16793 (I289089,I3570);
DFFARX1 I_16794 (I1391644,I3563,I289089,I289115,);
nand I_16795 (I289123,I1391623,I1391623);
and I_16796 (I289140,I289123,I1391650);
DFFARX1 I_16797 (I289140,I3563,I289089,I289166,);
nor I_16798 (I289057,I289166,I289115);
not I_16799 (I289188,I289166);
DFFARX1 I_16800 (I1391638,I3563,I289089,I289214,);
nand I_16801 (I289222,I289214,I1391641);
not I_16802 (I289239,I289222);
DFFARX1 I_16803 (I289239,I3563,I289089,I289265,);
not I_16804 (I289081,I289265);
nor I_16805 (I289287,I289115,I289222);
nor I_16806 (I289063,I289166,I289287);
DFFARX1 I_16807 (I1391632,I3563,I289089,I289327,);
DFFARX1 I_16808 (I289327,I3563,I289089,I289344,);
not I_16809 (I289352,I289344);
not I_16810 (I289369,I289327);
nand I_16811 (I289066,I289369,I289188);
nand I_16812 (I289400,I1391629,I1391626);
and I_16813 (I289417,I289400,I1391647);
DFFARX1 I_16814 (I289417,I3563,I289089,I289443,);
nor I_16815 (I289451,I289443,I289115);
DFFARX1 I_16816 (I289451,I3563,I289089,I289054,);
DFFARX1 I_16817 (I289443,I3563,I289089,I289072,);
nor I_16818 (I289496,I1391635,I1391626);
not I_16819 (I289513,I289496);
nor I_16820 (I289075,I289352,I289513);
nand I_16821 (I289060,I289369,I289513);
nor I_16822 (I289069,I289115,I289496);
DFFARX1 I_16823 (I289496,I3563,I289089,I289078,);
not I_16824 (I289616,I3570);
DFFARX1 I_16825 (I1134923,I3563,I289616,I289642,);
nand I_16826 (I289650,I1134938,I1134923);
and I_16827 (I289667,I289650,I1134941);
DFFARX1 I_16828 (I289667,I3563,I289616,I289693,);
nor I_16829 (I289584,I289693,I289642);
not I_16830 (I289715,I289693);
DFFARX1 I_16831 (I1134947,I3563,I289616,I289741,);
nand I_16832 (I289749,I289741,I1134929);
not I_16833 (I289766,I289749);
DFFARX1 I_16834 (I289766,I3563,I289616,I289792,);
not I_16835 (I289608,I289792);
nor I_16836 (I289814,I289642,I289749);
nor I_16837 (I289590,I289693,I289814);
DFFARX1 I_16838 (I1134926,I3563,I289616,I289854,);
DFFARX1 I_16839 (I289854,I3563,I289616,I289871,);
not I_16840 (I289879,I289871);
not I_16841 (I289896,I289854);
nand I_16842 (I289593,I289896,I289715);
nand I_16843 (I289927,I1134926,I1134932);
and I_16844 (I289944,I289927,I1134944);
DFFARX1 I_16845 (I289944,I3563,I289616,I289970,);
nor I_16846 (I289978,I289970,I289642);
DFFARX1 I_16847 (I289978,I3563,I289616,I289581,);
DFFARX1 I_16848 (I289970,I3563,I289616,I289599,);
nor I_16849 (I290023,I1134935,I1134932);
not I_16850 (I290040,I290023);
nor I_16851 (I289602,I289879,I290040);
nand I_16852 (I289587,I289896,I290040);
nor I_16853 (I289596,I289642,I290023);
DFFARX1 I_16854 (I290023,I3563,I289616,I289605,);
not I_16855 (I290143,I3570);
DFFARX1 I_16856 (I959452,I3563,I290143,I290169,);
nand I_16857 (I290177,I959449,I959467);
and I_16858 (I290194,I290177,I959458);
DFFARX1 I_16859 (I290194,I3563,I290143,I290220,);
nor I_16860 (I290111,I290220,I290169);
not I_16861 (I290242,I290220);
DFFARX1 I_16862 (I959473,I3563,I290143,I290268,);
nand I_16863 (I290276,I290268,I959455);
not I_16864 (I290293,I290276);
DFFARX1 I_16865 (I290293,I3563,I290143,I290319,);
not I_16866 (I290135,I290319);
nor I_16867 (I290341,I290169,I290276);
nor I_16868 (I290117,I290220,I290341);
DFFARX1 I_16869 (I959461,I3563,I290143,I290381,);
DFFARX1 I_16870 (I290381,I3563,I290143,I290398,);
not I_16871 (I290406,I290398);
not I_16872 (I290423,I290381);
nand I_16873 (I290120,I290423,I290242);
nand I_16874 (I290454,I959449,I959476);
and I_16875 (I290471,I290454,I959464);
DFFARX1 I_16876 (I290471,I3563,I290143,I290497,);
nor I_16877 (I290505,I290497,I290169);
DFFARX1 I_16878 (I290505,I3563,I290143,I290108,);
DFFARX1 I_16879 (I290497,I3563,I290143,I290126,);
nor I_16880 (I290550,I959470,I959476);
not I_16881 (I290567,I290550);
nor I_16882 (I290129,I290406,I290567);
nand I_16883 (I290114,I290423,I290567);
nor I_16884 (I290123,I290169,I290550);
DFFARX1 I_16885 (I290550,I3563,I290143,I290132,);
not I_16886 (I290670,I3570);
DFFARX1 I_16887 (I150456,I3563,I290670,I290696,);
nand I_16888 (I290704,I150468,I150477);
and I_16889 (I290721,I290704,I150456);
DFFARX1 I_16890 (I290721,I3563,I290670,I290747,);
nor I_16891 (I290638,I290747,I290696);
not I_16892 (I290769,I290747);
DFFARX1 I_16893 (I150471,I3563,I290670,I290795,);
nand I_16894 (I290803,I290795,I150459);
not I_16895 (I290820,I290803);
DFFARX1 I_16896 (I290820,I3563,I290670,I290846,);
not I_16897 (I290662,I290846);
nor I_16898 (I290868,I290696,I290803);
nor I_16899 (I290644,I290747,I290868);
DFFARX1 I_16900 (I150462,I3563,I290670,I290908,);
DFFARX1 I_16901 (I290908,I3563,I290670,I290925,);
not I_16902 (I290933,I290925);
not I_16903 (I290950,I290908);
nand I_16904 (I290647,I290950,I290769);
nand I_16905 (I290981,I150453,I150453);
and I_16906 (I290998,I290981,I150465);
DFFARX1 I_16907 (I290998,I3563,I290670,I291024,);
nor I_16908 (I291032,I291024,I290696);
DFFARX1 I_16909 (I291032,I3563,I290670,I290635,);
DFFARX1 I_16910 (I291024,I3563,I290670,I290653,);
nor I_16911 (I291077,I150474,I150453);
not I_16912 (I291094,I291077);
nor I_16913 (I290656,I290933,I291094);
nand I_16914 (I290641,I290950,I291094);
nor I_16915 (I290650,I290696,I291077);
DFFARX1 I_16916 (I291077,I3563,I290670,I290659,);
not I_16917 (I291197,I3570);
DFFARX1 I_16918 (I680389,I3563,I291197,I291223,);
nand I_16919 (I291231,I680380,I680395);
and I_16920 (I291248,I291231,I680401);
DFFARX1 I_16921 (I291248,I3563,I291197,I291274,);
nor I_16922 (I291165,I291274,I291223);
not I_16923 (I291296,I291274);
DFFARX1 I_16924 (I680386,I3563,I291197,I291322,);
nand I_16925 (I291330,I291322,I680380);
not I_16926 (I291347,I291330);
DFFARX1 I_16927 (I291347,I3563,I291197,I291373,);
not I_16928 (I291189,I291373);
nor I_16929 (I291395,I291223,I291330);
nor I_16930 (I291171,I291274,I291395);
DFFARX1 I_16931 (I680383,I3563,I291197,I291435,);
DFFARX1 I_16932 (I291435,I3563,I291197,I291452,);
not I_16933 (I291460,I291452);
not I_16934 (I291477,I291435);
nand I_16935 (I291174,I291477,I291296);
nand I_16936 (I291508,I680377,I680392);
and I_16937 (I291525,I291508,I680377);
DFFARX1 I_16938 (I291525,I3563,I291197,I291551,);
nor I_16939 (I291559,I291551,I291223);
DFFARX1 I_16940 (I291559,I3563,I291197,I291162,);
DFFARX1 I_16941 (I291551,I3563,I291197,I291180,);
nor I_16942 (I291604,I680398,I680392);
not I_16943 (I291621,I291604);
nor I_16944 (I291183,I291460,I291621);
nand I_16945 (I291168,I291477,I291621);
nor I_16946 (I291177,I291223,I291604);
DFFARX1 I_16947 (I291604,I3563,I291197,I291186,);
not I_16948 (I291724,I3570);
DFFARX1 I_16949 (I646868,I3563,I291724,I291750,);
nand I_16950 (I291758,I646853,I646856);
and I_16951 (I291775,I291758,I646871);
DFFARX1 I_16952 (I291775,I3563,I291724,I291801,);
nor I_16953 (I291692,I291801,I291750);
not I_16954 (I291823,I291801);
DFFARX1 I_16955 (I646865,I3563,I291724,I291849,);
nand I_16956 (I291857,I291849,I646856);
not I_16957 (I291874,I291857);
DFFARX1 I_16958 (I291874,I3563,I291724,I291900,);
not I_16959 (I291716,I291900);
nor I_16960 (I291922,I291750,I291857);
nor I_16961 (I291698,I291801,I291922);
DFFARX1 I_16962 (I646862,I3563,I291724,I291962,);
DFFARX1 I_16963 (I291962,I3563,I291724,I291979,);
not I_16964 (I291987,I291979);
not I_16965 (I292004,I291962);
nand I_16966 (I291701,I292004,I291823);
nand I_16967 (I292035,I646877,I646853);
and I_16968 (I292052,I292035,I646874);
DFFARX1 I_16969 (I292052,I3563,I291724,I292078,);
nor I_16970 (I292086,I292078,I291750);
DFFARX1 I_16971 (I292086,I3563,I291724,I291689,);
DFFARX1 I_16972 (I292078,I3563,I291724,I291707,);
nor I_16973 (I292131,I646859,I646853);
not I_16974 (I292148,I292131);
nor I_16975 (I291710,I291987,I292148);
nand I_16976 (I291695,I292004,I292148);
nor I_16977 (I291704,I291750,I292131);
DFFARX1 I_16978 (I292131,I3563,I291724,I291713,);
not I_16979 (I292251,I3570);
DFFARX1 I_16980 (I148348,I3563,I292251,I292277,);
nand I_16981 (I292285,I148360,I148369);
and I_16982 (I292302,I292285,I148348);
DFFARX1 I_16983 (I292302,I3563,I292251,I292328,);
nor I_16984 (I292219,I292328,I292277);
not I_16985 (I292350,I292328);
DFFARX1 I_16986 (I148363,I3563,I292251,I292376,);
nand I_16987 (I292384,I292376,I148351);
not I_16988 (I292401,I292384);
DFFARX1 I_16989 (I292401,I3563,I292251,I292427,);
not I_16990 (I292243,I292427);
nor I_16991 (I292449,I292277,I292384);
nor I_16992 (I292225,I292328,I292449);
DFFARX1 I_16993 (I148354,I3563,I292251,I292489,);
DFFARX1 I_16994 (I292489,I3563,I292251,I292506,);
not I_16995 (I292514,I292506);
not I_16996 (I292531,I292489);
nand I_16997 (I292228,I292531,I292350);
nand I_16998 (I292562,I148345,I148345);
and I_16999 (I292579,I292562,I148357);
DFFARX1 I_17000 (I292579,I3563,I292251,I292605,);
nor I_17001 (I292613,I292605,I292277);
DFFARX1 I_17002 (I292613,I3563,I292251,I292216,);
DFFARX1 I_17003 (I292605,I3563,I292251,I292234,);
nor I_17004 (I292658,I148366,I148345);
not I_17005 (I292675,I292658);
nor I_17006 (I292237,I292514,I292675);
nand I_17007 (I292222,I292531,I292675);
nor I_17008 (I292231,I292277,I292658);
DFFARX1 I_17009 (I292658,I3563,I292251,I292240,);
not I_17010 (I292778,I3570);
DFFARX1 I_17011 (I1344044,I3563,I292778,I292804,);
nand I_17012 (I292812,I1344023,I1344023);
and I_17013 (I292829,I292812,I1344050);
DFFARX1 I_17014 (I292829,I3563,I292778,I292855,);
nor I_17015 (I292746,I292855,I292804);
not I_17016 (I292877,I292855);
DFFARX1 I_17017 (I1344038,I3563,I292778,I292903,);
nand I_17018 (I292911,I292903,I1344041);
not I_17019 (I292928,I292911);
DFFARX1 I_17020 (I292928,I3563,I292778,I292954,);
not I_17021 (I292770,I292954);
nor I_17022 (I292976,I292804,I292911);
nor I_17023 (I292752,I292855,I292976);
DFFARX1 I_17024 (I1344032,I3563,I292778,I293016,);
DFFARX1 I_17025 (I293016,I3563,I292778,I293033,);
not I_17026 (I293041,I293033);
not I_17027 (I293058,I293016);
nand I_17028 (I292755,I293058,I292877);
nand I_17029 (I293089,I1344029,I1344026);
and I_17030 (I293106,I293089,I1344047);
DFFARX1 I_17031 (I293106,I3563,I292778,I293132,);
nor I_17032 (I293140,I293132,I292804);
DFFARX1 I_17033 (I293140,I3563,I292778,I292743,);
DFFARX1 I_17034 (I293132,I3563,I292778,I292761,);
nor I_17035 (I293185,I1344035,I1344026);
not I_17036 (I293202,I293185);
nor I_17037 (I292764,I293041,I293202);
nand I_17038 (I292749,I293058,I293202);
nor I_17039 (I292758,I292804,I293185);
DFFARX1 I_17040 (I293185,I3563,I292778,I292767,);
not I_17041 (I293305,I3570);
DFFARX1 I_17042 (I1092151,I3563,I293305,I293331,);
nand I_17043 (I293339,I1092166,I1092151);
and I_17044 (I293356,I293339,I1092169);
DFFARX1 I_17045 (I293356,I3563,I293305,I293382,);
nor I_17046 (I293273,I293382,I293331);
not I_17047 (I293404,I293382);
DFFARX1 I_17048 (I1092175,I3563,I293305,I293430,);
nand I_17049 (I293438,I293430,I1092157);
not I_17050 (I293455,I293438);
DFFARX1 I_17051 (I293455,I3563,I293305,I293481,);
not I_17052 (I293297,I293481);
nor I_17053 (I293503,I293331,I293438);
nor I_17054 (I293279,I293382,I293503);
DFFARX1 I_17055 (I1092154,I3563,I293305,I293543,);
DFFARX1 I_17056 (I293543,I3563,I293305,I293560,);
not I_17057 (I293568,I293560);
not I_17058 (I293585,I293543);
nand I_17059 (I293282,I293585,I293404);
nand I_17060 (I293616,I1092154,I1092160);
and I_17061 (I293633,I293616,I1092172);
DFFARX1 I_17062 (I293633,I3563,I293305,I293659,);
nor I_17063 (I293667,I293659,I293331);
DFFARX1 I_17064 (I293667,I3563,I293305,I293270,);
DFFARX1 I_17065 (I293659,I3563,I293305,I293288,);
nor I_17066 (I293712,I1092163,I1092160);
not I_17067 (I293729,I293712);
nor I_17068 (I293291,I293568,I293729);
nand I_17069 (I293276,I293585,I293729);
nor I_17070 (I293285,I293331,I293712);
DFFARX1 I_17071 (I293712,I3563,I293305,I293294,);
not I_17072 (I293832,I3570);
DFFARX1 I_17073 (I749749,I3563,I293832,I293858,);
nand I_17074 (I293866,I749740,I749755);
and I_17075 (I293883,I293866,I749761);
DFFARX1 I_17076 (I293883,I3563,I293832,I293909,);
nor I_17077 (I293800,I293909,I293858);
not I_17078 (I293931,I293909);
DFFARX1 I_17079 (I749746,I3563,I293832,I293957,);
nand I_17080 (I293965,I293957,I749740);
not I_17081 (I293982,I293965);
DFFARX1 I_17082 (I293982,I3563,I293832,I294008,);
not I_17083 (I293824,I294008);
nor I_17084 (I294030,I293858,I293965);
nor I_17085 (I293806,I293909,I294030);
DFFARX1 I_17086 (I749743,I3563,I293832,I294070,);
DFFARX1 I_17087 (I294070,I3563,I293832,I294087,);
not I_17088 (I294095,I294087);
not I_17089 (I294112,I294070);
nand I_17090 (I293809,I294112,I293931);
nand I_17091 (I294143,I749737,I749752);
and I_17092 (I294160,I294143,I749737);
DFFARX1 I_17093 (I294160,I3563,I293832,I294186,);
nor I_17094 (I294194,I294186,I293858);
DFFARX1 I_17095 (I294194,I3563,I293832,I293797,);
DFFARX1 I_17096 (I294186,I3563,I293832,I293815,);
nor I_17097 (I294239,I749758,I749752);
not I_17098 (I294256,I294239);
nor I_17099 (I293818,I294095,I294256);
nand I_17100 (I293803,I294112,I294256);
nor I_17101 (I293812,I293858,I294239);
DFFARX1 I_17102 (I294239,I3563,I293832,I293821,);
not I_17103 (I294359,I3570);
DFFARX1 I_17104 (I1336309,I3563,I294359,I294385,);
nand I_17105 (I294393,I1336288,I1336288);
and I_17106 (I294410,I294393,I1336315);
DFFARX1 I_17107 (I294410,I3563,I294359,I294436,);
nor I_17108 (I294327,I294436,I294385);
not I_17109 (I294458,I294436);
DFFARX1 I_17110 (I1336303,I3563,I294359,I294484,);
nand I_17111 (I294492,I294484,I1336306);
not I_17112 (I294509,I294492);
DFFARX1 I_17113 (I294509,I3563,I294359,I294535,);
not I_17114 (I294351,I294535);
nor I_17115 (I294557,I294385,I294492);
nor I_17116 (I294333,I294436,I294557);
DFFARX1 I_17117 (I1336297,I3563,I294359,I294597,);
DFFARX1 I_17118 (I294597,I3563,I294359,I294614,);
not I_17119 (I294622,I294614);
not I_17120 (I294639,I294597);
nand I_17121 (I294336,I294639,I294458);
nand I_17122 (I294670,I1336294,I1336291);
and I_17123 (I294687,I294670,I1336312);
DFFARX1 I_17124 (I294687,I3563,I294359,I294713,);
nor I_17125 (I294721,I294713,I294385);
DFFARX1 I_17126 (I294721,I3563,I294359,I294324,);
DFFARX1 I_17127 (I294713,I3563,I294359,I294342,);
nor I_17128 (I294766,I1336300,I1336291);
not I_17129 (I294783,I294766);
nor I_17130 (I294345,I294622,I294783);
nand I_17131 (I294330,I294639,I294783);
nor I_17132 (I294339,I294385,I294766);
DFFARX1 I_17133 (I294766,I3563,I294359,I294348,);
not I_17134 (I294886,I3570);
DFFARX1 I_17135 (I1452,I3563,I294886,I294912,);
nand I_17136 (I294920,I2628,I3308);
and I_17137 (I294937,I294920,I1900);
DFFARX1 I_17138 (I294937,I3563,I294886,I294963,);
nor I_17139 (I294854,I294963,I294912);
not I_17140 (I294985,I294963);
DFFARX1 I_17141 (I2076,I3563,I294886,I295011,);
nand I_17142 (I295019,I295011,I3148);
not I_17143 (I295036,I295019);
DFFARX1 I_17144 (I295036,I3563,I294886,I295062,);
not I_17145 (I294878,I295062);
nor I_17146 (I295084,I294912,I295019);
nor I_17147 (I294860,I294963,I295084);
DFFARX1 I_17148 (I1772,I3563,I294886,I295124,);
DFFARX1 I_17149 (I295124,I3563,I294886,I295141,);
not I_17150 (I295149,I295141);
not I_17151 (I295166,I295124);
nand I_17152 (I294863,I295166,I294985);
nand I_17153 (I295197,I3244,I3428);
and I_17154 (I295214,I295197,I1428);
DFFARX1 I_17155 (I295214,I3563,I294886,I295240,);
nor I_17156 (I295248,I295240,I294912);
DFFARX1 I_17157 (I295248,I3563,I294886,I294851,);
DFFARX1 I_17158 (I295240,I3563,I294886,I294869,);
nor I_17159 (I295293,I2852,I3428);
not I_17160 (I295310,I295293);
nor I_17161 (I294872,I295149,I295310);
nand I_17162 (I294857,I295166,I295310);
nor I_17163 (I294866,I294912,I295293);
DFFARX1 I_17164 (I295293,I3563,I294886,I294875,);
not I_17165 (I295413,I3570);
DFFARX1 I_17166 (I1031804,I3563,I295413,I295439,);
nand I_17167 (I295447,I1031801,I1031819);
and I_17168 (I295464,I295447,I1031810);
DFFARX1 I_17169 (I295464,I3563,I295413,I295490,);
nor I_17170 (I295381,I295490,I295439);
not I_17171 (I295512,I295490);
DFFARX1 I_17172 (I1031825,I3563,I295413,I295538,);
nand I_17173 (I295546,I295538,I1031807);
not I_17174 (I295563,I295546);
DFFARX1 I_17175 (I295563,I3563,I295413,I295589,);
not I_17176 (I295405,I295589);
nor I_17177 (I295611,I295439,I295546);
nor I_17178 (I295387,I295490,I295611);
DFFARX1 I_17179 (I1031813,I3563,I295413,I295651,);
DFFARX1 I_17180 (I295651,I3563,I295413,I295668,);
not I_17181 (I295676,I295668);
not I_17182 (I295693,I295651);
nand I_17183 (I295390,I295693,I295512);
nand I_17184 (I295724,I1031801,I1031828);
and I_17185 (I295741,I295724,I1031816);
DFFARX1 I_17186 (I295741,I3563,I295413,I295767,);
nor I_17187 (I295775,I295767,I295439);
DFFARX1 I_17188 (I295775,I3563,I295413,I295378,);
DFFARX1 I_17189 (I295767,I3563,I295413,I295396,);
nor I_17190 (I295820,I1031822,I1031828);
not I_17191 (I295837,I295820);
nor I_17192 (I295399,I295676,I295837);
nand I_17193 (I295384,I295693,I295837);
nor I_17194 (I295393,I295439,I295820);
DFFARX1 I_17195 (I295820,I3563,I295413,I295402,);
not I_17196 (I295940,I3570);
DFFARX1 I_17197 (I1159199,I3563,I295940,I295966,);
nand I_17198 (I295974,I1159214,I1159199);
and I_17199 (I295991,I295974,I1159217);
DFFARX1 I_17200 (I295991,I3563,I295940,I296017,);
nor I_17201 (I295908,I296017,I295966);
not I_17202 (I296039,I296017);
DFFARX1 I_17203 (I1159223,I3563,I295940,I296065,);
nand I_17204 (I296073,I296065,I1159205);
not I_17205 (I296090,I296073);
DFFARX1 I_17206 (I296090,I3563,I295940,I296116,);
not I_17207 (I295932,I296116);
nor I_17208 (I296138,I295966,I296073);
nor I_17209 (I295914,I296017,I296138);
DFFARX1 I_17210 (I1159202,I3563,I295940,I296178,);
DFFARX1 I_17211 (I296178,I3563,I295940,I296195,);
not I_17212 (I296203,I296195);
not I_17213 (I296220,I296178);
nand I_17214 (I295917,I296220,I296039);
nand I_17215 (I296251,I1159202,I1159208);
and I_17216 (I296268,I296251,I1159220);
DFFARX1 I_17217 (I296268,I3563,I295940,I296294,);
nor I_17218 (I296302,I296294,I295966);
DFFARX1 I_17219 (I296302,I3563,I295940,I295905,);
DFFARX1 I_17220 (I296294,I3563,I295940,I295923,);
nor I_17221 (I296347,I1159211,I1159208);
not I_17222 (I296364,I296347);
nor I_17223 (I295926,I296203,I296364);
nand I_17224 (I295911,I296220,I296364);
nor I_17225 (I295920,I295966,I296347);
DFFARX1 I_17226 (I296347,I3563,I295940,I295929,);
not I_17227 (I296467,I3570);
DFFARX1 I_17228 (I1180007,I3563,I296467,I296493,);
nand I_17229 (I296501,I1180022,I1180007);
and I_17230 (I296518,I296501,I1180025);
DFFARX1 I_17231 (I296518,I3563,I296467,I296544,);
nor I_17232 (I296435,I296544,I296493);
not I_17233 (I296566,I296544);
DFFARX1 I_17234 (I1180031,I3563,I296467,I296592,);
nand I_17235 (I296600,I296592,I1180013);
not I_17236 (I296617,I296600);
DFFARX1 I_17237 (I296617,I3563,I296467,I296643,);
not I_17238 (I296459,I296643);
nor I_17239 (I296665,I296493,I296600);
nor I_17240 (I296441,I296544,I296665);
DFFARX1 I_17241 (I1180010,I3563,I296467,I296705,);
DFFARX1 I_17242 (I296705,I3563,I296467,I296722,);
not I_17243 (I296730,I296722);
not I_17244 (I296747,I296705);
nand I_17245 (I296444,I296747,I296566);
nand I_17246 (I296778,I1180010,I1180016);
and I_17247 (I296795,I296778,I1180028);
DFFARX1 I_17248 (I296795,I3563,I296467,I296821,);
nor I_17249 (I296829,I296821,I296493);
DFFARX1 I_17250 (I296829,I3563,I296467,I296432,);
DFFARX1 I_17251 (I296821,I3563,I296467,I296450,);
nor I_17252 (I296874,I1180019,I1180016);
not I_17253 (I296891,I296874);
nor I_17254 (I296453,I296730,I296891);
nand I_17255 (I296438,I296747,I296891);
nor I_17256 (I296447,I296493,I296874);
DFFARX1 I_17257 (I296874,I3563,I296467,I296456,);
not I_17258 (I296994,I3570);
DFFARX1 I_17259 (I1199081,I3563,I296994,I297020,);
nand I_17260 (I297028,I1199096,I1199081);
and I_17261 (I297045,I297028,I1199099);
DFFARX1 I_17262 (I297045,I3563,I296994,I297071,);
nor I_17263 (I296962,I297071,I297020);
not I_17264 (I297093,I297071);
DFFARX1 I_17265 (I1199105,I3563,I296994,I297119,);
nand I_17266 (I297127,I297119,I1199087);
not I_17267 (I297144,I297127);
DFFARX1 I_17268 (I297144,I3563,I296994,I297170,);
not I_17269 (I296986,I297170);
nor I_17270 (I297192,I297020,I297127);
nor I_17271 (I296968,I297071,I297192);
DFFARX1 I_17272 (I1199084,I3563,I296994,I297232,);
DFFARX1 I_17273 (I297232,I3563,I296994,I297249,);
not I_17274 (I297257,I297249);
not I_17275 (I297274,I297232);
nand I_17276 (I296971,I297274,I297093);
nand I_17277 (I297305,I1199084,I1199090);
and I_17278 (I297322,I297305,I1199102);
DFFARX1 I_17279 (I297322,I3563,I296994,I297348,);
nor I_17280 (I297356,I297348,I297020);
DFFARX1 I_17281 (I297356,I3563,I296994,I296959,);
DFFARX1 I_17282 (I297348,I3563,I296994,I296977,);
nor I_17283 (I297401,I1199093,I1199090);
not I_17284 (I297418,I297401);
nor I_17285 (I296980,I297257,I297418);
nand I_17286 (I296965,I297274,I297418);
nor I_17287 (I296974,I297020,I297401);
DFFARX1 I_17288 (I297401,I3563,I296994,I296983,);
not I_17289 (I297521,I3570);
DFFARX1 I_17290 (I764199,I3563,I297521,I297547,);
nand I_17291 (I297555,I764190,I764205);
and I_17292 (I297572,I297555,I764211);
DFFARX1 I_17293 (I297572,I3563,I297521,I297598,);
nor I_17294 (I297489,I297598,I297547);
not I_17295 (I297620,I297598);
DFFARX1 I_17296 (I764196,I3563,I297521,I297646,);
nand I_17297 (I297654,I297646,I764190);
not I_17298 (I297671,I297654);
DFFARX1 I_17299 (I297671,I3563,I297521,I297697,);
not I_17300 (I297513,I297697);
nor I_17301 (I297719,I297547,I297654);
nor I_17302 (I297495,I297598,I297719);
DFFARX1 I_17303 (I764193,I3563,I297521,I297759,);
DFFARX1 I_17304 (I297759,I3563,I297521,I297776,);
not I_17305 (I297784,I297776);
not I_17306 (I297801,I297759);
nand I_17307 (I297498,I297801,I297620);
nand I_17308 (I297832,I764187,I764202);
and I_17309 (I297849,I297832,I764187);
DFFARX1 I_17310 (I297849,I3563,I297521,I297875,);
nor I_17311 (I297883,I297875,I297547);
DFFARX1 I_17312 (I297883,I3563,I297521,I297486,);
DFFARX1 I_17313 (I297875,I3563,I297521,I297504,);
nor I_17314 (I297928,I764208,I764202);
not I_17315 (I297945,I297928);
nor I_17316 (I297507,I297784,I297945);
nand I_17317 (I297492,I297801,I297945);
nor I_17318 (I297501,I297547,I297928);
DFFARX1 I_17319 (I297928,I3563,I297521,I297510,);
not I_17320 (I298048,I3570);
DFFARX1 I_17321 (I1185209,I3563,I298048,I298074,);
nand I_17322 (I298082,I1185224,I1185209);
and I_17323 (I298099,I298082,I1185227);
DFFARX1 I_17324 (I298099,I3563,I298048,I298125,);
nor I_17325 (I298016,I298125,I298074);
not I_17326 (I298147,I298125);
DFFARX1 I_17327 (I1185233,I3563,I298048,I298173,);
nand I_17328 (I298181,I298173,I1185215);
not I_17329 (I298198,I298181);
DFFARX1 I_17330 (I298198,I3563,I298048,I298224,);
not I_17331 (I298040,I298224);
nor I_17332 (I298246,I298074,I298181);
nor I_17333 (I298022,I298125,I298246);
DFFARX1 I_17334 (I1185212,I3563,I298048,I298286,);
DFFARX1 I_17335 (I298286,I3563,I298048,I298303,);
not I_17336 (I298311,I298303);
not I_17337 (I298328,I298286);
nand I_17338 (I298025,I298328,I298147);
nand I_17339 (I298359,I1185212,I1185218);
and I_17340 (I298376,I298359,I1185230);
DFFARX1 I_17341 (I298376,I3563,I298048,I298402,);
nor I_17342 (I298410,I298402,I298074);
DFFARX1 I_17343 (I298410,I3563,I298048,I298013,);
DFFARX1 I_17344 (I298402,I3563,I298048,I298031,);
nor I_17345 (I298455,I1185221,I1185218);
not I_17346 (I298472,I298455);
nor I_17347 (I298034,I298311,I298472);
nand I_17348 (I298019,I298328,I298472);
nor I_17349 (I298028,I298074,I298455);
DFFARX1 I_17350 (I298455,I3563,I298048,I298037,);
not I_17351 (I298575,I3570);
DFFARX1 I_17352 (I1313778,I3563,I298575,I298601,);
nand I_17353 (I298609,I1313775,I1313766);
and I_17354 (I298626,I298609,I1313763);
DFFARX1 I_17355 (I298626,I3563,I298575,I298652,);
nor I_17356 (I298543,I298652,I298601);
not I_17357 (I298674,I298652);
DFFARX1 I_17358 (I1313772,I3563,I298575,I298700,);
nand I_17359 (I298708,I298700,I1313781);
not I_17360 (I298725,I298708);
DFFARX1 I_17361 (I298725,I3563,I298575,I298751,);
not I_17362 (I298567,I298751);
nor I_17363 (I298773,I298601,I298708);
nor I_17364 (I298549,I298652,I298773);
DFFARX1 I_17365 (I1313784,I3563,I298575,I298813,);
DFFARX1 I_17366 (I298813,I3563,I298575,I298830,);
not I_17367 (I298838,I298830);
not I_17368 (I298855,I298813);
nand I_17369 (I298552,I298855,I298674);
nand I_17370 (I298886,I1313763,I1313769);
and I_17371 (I298903,I298886,I1313787);
DFFARX1 I_17372 (I298903,I3563,I298575,I298929,);
nor I_17373 (I298937,I298929,I298601);
DFFARX1 I_17374 (I298937,I3563,I298575,I298540,);
DFFARX1 I_17375 (I298929,I3563,I298575,I298558,);
nor I_17376 (I298982,I1313766,I1313769);
not I_17377 (I298999,I298982);
nor I_17378 (I298561,I298838,I298999);
nand I_17379 (I298546,I298855,I298999);
nor I_17380 (I298555,I298601,I298982);
DFFARX1 I_17381 (I298982,I3563,I298575,I298564,);
not I_17382 (I299102,I3570);
DFFARX1 I_17383 (I430030,I3563,I299102,I299128,);
nand I_17384 (I299136,I430042,I430021);
and I_17385 (I299153,I299136,I430045);
DFFARX1 I_17386 (I299153,I3563,I299102,I299179,);
nor I_17387 (I299070,I299179,I299128);
not I_17388 (I299201,I299179);
DFFARX1 I_17389 (I430036,I3563,I299102,I299227,);
nand I_17390 (I299235,I299227,I430018);
not I_17391 (I299252,I299235);
DFFARX1 I_17392 (I299252,I3563,I299102,I299278,);
not I_17393 (I299094,I299278);
nor I_17394 (I299300,I299128,I299235);
nor I_17395 (I299076,I299179,I299300);
DFFARX1 I_17396 (I430033,I3563,I299102,I299340,);
DFFARX1 I_17397 (I299340,I3563,I299102,I299357,);
not I_17398 (I299365,I299357);
not I_17399 (I299382,I299340);
nand I_17400 (I299079,I299382,I299201);
nand I_17401 (I299413,I430018,I430024);
and I_17402 (I299430,I299413,I430027);
DFFARX1 I_17403 (I299430,I3563,I299102,I299456,);
nor I_17404 (I299464,I299456,I299128);
DFFARX1 I_17405 (I299464,I3563,I299102,I299067,);
DFFARX1 I_17406 (I299456,I3563,I299102,I299085,);
nor I_17407 (I299509,I430039,I430024);
not I_17408 (I299526,I299509);
nor I_17409 (I299088,I299365,I299526);
nand I_17410 (I299073,I299382,I299526);
nor I_17411 (I299082,I299128,I299509);
DFFARX1 I_17412 (I299509,I3563,I299102,I299091,);
not I_17413 (I299629,I3570);
DFFARX1 I_17414 (I940718,I3563,I299629,I299655,);
nand I_17415 (I299663,I940715,I940733);
and I_17416 (I299680,I299663,I940724);
DFFARX1 I_17417 (I299680,I3563,I299629,I299706,);
nor I_17418 (I299597,I299706,I299655);
not I_17419 (I299728,I299706);
DFFARX1 I_17420 (I940739,I3563,I299629,I299754,);
nand I_17421 (I299762,I299754,I940721);
not I_17422 (I299779,I299762);
DFFARX1 I_17423 (I299779,I3563,I299629,I299805,);
not I_17424 (I299621,I299805);
nor I_17425 (I299827,I299655,I299762);
nor I_17426 (I299603,I299706,I299827);
DFFARX1 I_17427 (I940727,I3563,I299629,I299867,);
DFFARX1 I_17428 (I299867,I3563,I299629,I299884,);
not I_17429 (I299892,I299884);
not I_17430 (I299909,I299867);
nand I_17431 (I299606,I299909,I299728);
nand I_17432 (I299940,I940715,I940742);
and I_17433 (I299957,I299940,I940730);
DFFARX1 I_17434 (I299957,I3563,I299629,I299983,);
nor I_17435 (I299991,I299983,I299655);
DFFARX1 I_17436 (I299991,I3563,I299629,I299594,);
DFFARX1 I_17437 (I299983,I3563,I299629,I299612,);
nor I_17438 (I300036,I940736,I940742);
not I_17439 (I300053,I300036);
nor I_17440 (I299615,I299892,I300053);
nand I_17441 (I299600,I299909,I300053);
nor I_17442 (I299609,I299655,I300036);
DFFARX1 I_17443 (I300036,I3563,I299629,I299618,);
not I_17444 (I300156,I3570);
DFFARX1 I_17445 (I888001,I3563,I300156,I300182,);
nand I_17446 (I300190,I888004,I887998);
and I_17447 (I300207,I300190,I888010);
DFFARX1 I_17448 (I300207,I3563,I300156,I300233,);
nor I_17449 (I300124,I300233,I300182);
not I_17450 (I300255,I300233);
DFFARX1 I_17451 (I888013,I3563,I300156,I300281,);
nand I_17452 (I300289,I300281,I888004);
not I_17453 (I300306,I300289);
DFFARX1 I_17454 (I300306,I3563,I300156,I300332,);
not I_17455 (I300148,I300332);
nor I_17456 (I300354,I300182,I300289);
nor I_17457 (I300130,I300233,I300354);
DFFARX1 I_17458 (I888016,I3563,I300156,I300394,);
DFFARX1 I_17459 (I300394,I3563,I300156,I300411,);
not I_17460 (I300419,I300411);
not I_17461 (I300436,I300394);
nand I_17462 (I300133,I300436,I300255);
nand I_17463 (I300467,I887998,I888007);
and I_17464 (I300484,I300467,I888001);
DFFARX1 I_17465 (I300484,I3563,I300156,I300510,);
nor I_17466 (I300518,I300510,I300182);
DFFARX1 I_17467 (I300518,I3563,I300156,I300121,);
DFFARX1 I_17468 (I300510,I3563,I300156,I300139,);
nor I_17469 (I300563,I888019,I888007);
not I_17470 (I300580,I300563);
nor I_17471 (I300142,I300419,I300580);
nand I_17472 (I300127,I300436,I300580);
nor I_17473 (I300136,I300182,I300563);
DFFARX1 I_17474 (I300563,I3563,I300156,I300145,);
not I_17475 (I300683,I3570);
DFFARX1 I_17476 (I423502,I3563,I300683,I300709,);
nand I_17477 (I300717,I423514,I423493);
and I_17478 (I300734,I300717,I423517);
DFFARX1 I_17479 (I300734,I3563,I300683,I300760,);
nor I_17480 (I300651,I300760,I300709);
not I_17481 (I300782,I300760);
DFFARX1 I_17482 (I423508,I3563,I300683,I300808,);
nand I_17483 (I300816,I300808,I423490);
not I_17484 (I300833,I300816);
DFFARX1 I_17485 (I300833,I3563,I300683,I300859,);
not I_17486 (I300675,I300859);
nor I_17487 (I300881,I300709,I300816);
nor I_17488 (I300657,I300760,I300881);
DFFARX1 I_17489 (I423505,I3563,I300683,I300921,);
DFFARX1 I_17490 (I300921,I3563,I300683,I300938,);
not I_17491 (I300946,I300938);
not I_17492 (I300963,I300921);
nand I_17493 (I300660,I300963,I300782);
nand I_17494 (I300994,I423490,I423496);
and I_17495 (I301011,I300994,I423499);
DFFARX1 I_17496 (I301011,I3563,I300683,I301037,);
nor I_17497 (I301045,I301037,I300709);
DFFARX1 I_17498 (I301045,I3563,I300683,I300648,);
DFFARX1 I_17499 (I301037,I3563,I300683,I300666,);
nor I_17500 (I301090,I423511,I423496);
not I_17501 (I301107,I301090);
nor I_17502 (I300669,I300946,I301107);
nand I_17503 (I300654,I300963,I301107);
nor I_17504 (I300663,I300709,I301090);
DFFARX1 I_17505 (I301090,I3563,I300683,I300672,);
not I_17506 (I301210,I3570);
DFFARX1 I_17507 (I1219311,I3563,I301210,I301236,);
nand I_17508 (I301244,I1219326,I1219311);
and I_17509 (I301261,I301244,I1219329);
DFFARX1 I_17510 (I301261,I3563,I301210,I301287,);
nor I_17511 (I301178,I301287,I301236);
not I_17512 (I301309,I301287);
DFFARX1 I_17513 (I1219335,I3563,I301210,I301335,);
nand I_17514 (I301343,I301335,I1219317);
not I_17515 (I301360,I301343);
DFFARX1 I_17516 (I301360,I3563,I301210,I301386,);
not I_17517 (I301202,I301386);
nor I_17518 (I301408,I301236,I301343);
nor I_17519 (I301184,I301287,I301408);
DFFARX1 I_17520 (I1219314,I3563,I301210,I301448,);
DFFARX1 I_17521 (I301448,I3563,I301210,I301465,);
not I_17522 (I301473,I301465);
not I_17523 (I301490,I301448);
nand I_17524 (I301187,I301490,I301309);
nand I_17525 (I301521,I1219314,I1219320);
and I_17526 (I301538,I301521,I1219332);
DFFARX1 I_17527 (I301538,I3563,I301210,I301564,);
nor I_17528 (I301572,I301564,I301236);
DFFARX1 I_17529 (I301572,I3563,I301210,I301175,);
DFFARX1 I_17530 (I301564,I3563,I301210,I301193,);
nor I_17531 (I301617,I1219323,I1219320);
not I_17532 (I301634,I301617);
nor I_17533 (I301196,I301473,I301634);
nand I_17534 (I301181,I301490,I301634);
nor I_17535 (I301190,I301236,I301617);
DFFARX1 I_17536 (I301617,I3563,I301210,I301199,);
not I_17537 (I301737,I3570);
DFFARX1 I_17538 (I145713,I3563,I301737,I301763,);
nand I_17539 (I301771,I145725,I145734);
and I_17540 (I301788,I301771,I145713);
DFFARX1 I_17541 (I301788,I3563,I301737,I301814,);
nor I_17542 (I301705,I301814,I301763);
not I_17543 (I301836,I301814);
DFFARX1 I_17544 (I145728,I3563,I301737,I301862,);
nand I_17545 (I301870,I301862,I145716);
not I_17546 (I301887,I301870);
DFFARX1 I_17547 (I301887,I3563,I301737,I301913,);
not I_17548 (I301729,I301913);
nor I_17549 (I301935,I301763,I301870);
nor I_17550 (I301711,I301814,I301935);
DFFARX1 I_17551 (I145719,I3563,I301737,I301975,);
DFFARX1 I_17552 (I301975,I3563,I301737,I301992,);
not I_17553 (I302000,I301992);
not I_17554 (I302017,I301975);
nand I_17555 (I301714,I302017,I301836);
nand I_17556 (I302048,I145710,I145710);
and I_17557 (I302065,I302048,I145722);
DFFARX1 I_17558 (I302065,I3563,I301737,I302091,);
nor I_17559 (I302099,I302091,I301763);
DFFARX1 I_17560 (I302099,I3563,I301737,I301702,);
DFFARX1 I_17561 (I302091,I3563,I301737,I301720,);
nor I_17562 (I302144,I145731,I145710);
not I_17563 (I302161,I302144);
nor I_17564 (I301723,I302000,I302161);
nand I_17565 (I301708,I302017,I302161);
nor I_17566 (I301717,I301763,I302144);
DFFARX1 I_17567 (I302144,I3563,I301737,I301726,);
not I_17568 (I302264,I3570);
DFFARX1 I_17569 (I1152841,I3563,I302264,I302290,);
nand I_17570 (I302298,I1152856,I1152841);
and I_17571 (I302315,I302298,I1152859);
DFFARX1 I_17572 (I302315,I3563,I302264,I302341,);
nor I_17573 (I302232,I302341,I302290);
not I_17574 (I302363,I302341);
DFFARX1 I_17575 (I1152865,I3563,I302264,I302389,);
nand I_17576 (I302397,I302389,I1152847);
not I_17577 (I302414,I302397);
DFFARX1 I_17578 (I302414,I3563,I302264,I302440,);
not I_17579 (I302256,I302440);
nor I_17580 (I302462,I302290,I302397);
nor I_17581 (I302238,I302341,I302462);
DFFARX1 I_17582 (I1152844,I3563,I302264,I302502,);
DFFARX1 I_17583 (I302502,I3563,I302264,I302519,);
not I_17584 (I302527,I302519);
not I_17585 (I302544,I302502);
nand I_17586 (I302241,I302544,I302363);
nand I_17587 (I302575,I1152844,I1152850);
and I_17588 (I302592,I302575,I1152862);
DFFARX1 I_17589 (I302592,I3563,I302264,I302618,);
nor I_17590 (I302626,I302618,I302290);
DFFARX1 I_17591 (I302626,I3563,I302264,I302229,);
DFFARX1 I_17592 (I302618,I3563,I302264,I302247,);
nor I_17593 (I302671,I1152853,I1152850);
not I_17594 (I302688,I302671);
nor I_17595 (I302250,I302527,I302688);
nand I_17596 (I302235,I302544,I302688);
nor I_17597 (I302244,I302290,I302671);
DFFARX1 I_17598 (I302671,I3563,I302264,I302253,);
not I_17599 (I302791,I3570);
DFFARX1 I_17600 (I1278523,I3563,I302791,I302817,);
nand I_17601 (I302825,I1278505,I1278529);
and I_17602 (I302842,I302825,I1278520);
DFFARX1 I_17603 (I302842,I3563,I302791,I302868,);
nor I_17604 (I302759,I302868,I302817);
not I_17605 (I302890,I302868);
DFFARX1 I_17606 (I1278526,I3563,I302791,I302916,);
nand I_17607 (I302924,I302916,I1278514);
not I_17608 (I302941,I302924);
DFFARX1 I_17609 (I302941,I3563,I302791,I302967,);
not I_17610 (I302783,I302967);
nor I_17611 (I302989,I302817,I302924);
nor I_17612 (I302765,I302868,I302989);
DFFARX1 I_17613 (I1278505,I3563,I302791,I303029,);
DFFARX1 I_17614 (I303029,I3563,I302791,I303046,);
not I_17615 (I303054,I303046);
not I_17616 (I303071,I303029);
nand I_17617 (I302768,I303071,I302890);
nand I_17618 (I303102,I1278511,I1278508);
and I_17619 (I303119,I303102,I1278517);
DFFARX1 I_17620 (I303119,I3563,I302791,I303145,);
nor I_17621 (I303153,I303145,I302817);
DFFARX1 I_17622 (I303153,I3563,I302791,I302756,);
DFFARX1 I_17623 (I303145,I3563,I302791,I302774,);
nor I_17624 (I303198,I1278508,I1278508);
not I_17625 (I303215,I303198);
nor I_17626 (I302777,I303054,I303215);
nand I_17627 (I302762,I303071,I303215);
nor I_17628 (I302771,I302817,I303198);
DFFARX1 I_17629 (I303198,I3563,I302791,I302780,);
not I_17630 (I303318,I3570);
DFFARX1 I_17631 (I938780,I3563,I303318,I303344,);
nand I_17632 (I303352,I938777,I938795);
and I_17633 (I303369,I303352,I938786);
DFFARX1 I_17634 (I303369,I3563,I303318,I303395,);
nor I_17635 (I303286,I303395,I303344);
not I_17636 (I303417,I303395);
DFFARX1 I_17637 (I938801,I3563,I303318,I303443,);
nand I_17638 (I303451,I303443,I938783);
not I_17639 (I303468,I303451);
DFFARX1 I_17640 (I303468,I3563,I303318,I303494,);
not I_17641 (I303310,I303494);
nor I_17642 (I303516,I303344,I303451);
nor I_17643 (I303292,I303395,I303516);
DFFARX1 I_17644 (I938789,I3563,I303318,I303556,);
DFFARX1 I_17645 (I303556,I3563,I303318,I303573,);
not I_17646 (I303581,I303573);
not I_17647 (I303598,I303556);
nand I_17648 (I303295,I303598,I303417);
nand I_17649 (I303629,I938777,I938804);
and I_17650 (I303646,I303629,I938792);
DFFARX1 I_17651 (I303646,I3563,I303318,I303672,);
nor I_17652 (I303680,I303672,I303344);
DFFARX1 I_17653 (I303680,I3563,I303318,I303283,);
DFFARX1 I_17654 (I303672,I3563,I303318,I303301,);
nor I_17655 (I303725,I938798,I938804);
not I_17656 (I303742,I303725);
nor I_17657 (I303304,I303581,I303742);
nand I_17658 (I303289,I303598,I303742);
nor I_17659 (I303298,I303344,I303725);
DFFARX1 I_17660 (I303725,I3563,I303318,I303307,);
not I_17661 (I303845,I3570);
DFFARX1 I_17662 (I161952,I3563,I303845,I303871,);
nand I_17663 (I303879,I161937,I161928);
and I_17664 (I303896,I303879,I161943);
DFFARX1 I_17665 (I303896,I3563,I303845,I303922,);
nor I_17666 (I303813,I303922,I303871);
not I_17667 (I303944,I303922);
DFFARX1 I_17668 (I161955,I3563,I303845,I303970,);
nand I_17669 (I303978,I303970,I161946);
not I_17670 (I303995,I303978);
DFFARX1 I_17671 (I303995,I3563,I303845,I304021,);
not I_17672 (I303837,I304021);
nor I_17673 (I304043,I303871,I303978);
nor I_17674 (I303819,I303922,I304043);
DFFARX1 I_17675 (I161934,I3563,I303845,I304083,);
DFFARX1 I_17676 (I304083,I3563,I303845,I304100,);
not I_17677 (I304108,I304100);
not I_17678 (I304125,I304083);
nand I_17679 (I303822,I304125,I303944);
nand I_17680 (I304156,I161940,I161931);
and I_17681 (I304173,I304156,I161928);
DFFARX1 I_17682 (I304173,I3563,I303845,I304199,);
nor I_17683 (I304207,I304199,I303871);
DFFARX1 I_17684 (I304207,I3563,I303845,I303810,);
DFFARX1 I_17685 (I304199,I3563,I303845,I303828,);
nor I_17686 (I304252,I161949,I161931);
not I_17687 (I304269,I304252);
nor I_17688 (I303831,I304108,I304269);
nand I_17689 (I303816,I304125,I304269);
nor I_17690 (I303825,I303871,I304252);
DFFARX1 I_17691 (I304252,I3563,I303845,I303834,);
not I_17692 (I304372,I3570);
DFFARX1 I_17693 (I498030,I3563,I304372,I304398,);
nand I_17694 (I304406,I498042,I498021);
and I_17695 (I304423,I304406,I498045);
DFFARX1 I_17696 (I304423,I3563,I304372,I304449,);
nor I_17697 (I304340,I304449,I304398);
not I_17698 (I304471,I304449);
DFFARX1 I_17699 (I498036,I3563,I304372,I304497,);
nand I_17700 (I304505,I304497,I498018);
not I_17701 (I304522,I304505);
DFFARX1 I_17702 (I304522,I3563,I304372,I304548,);
not I_17703 (I304364,I304548);
nor I_17704 (I304570,I304398,I304505);
nor I_17705 (I304346,I304449,I304570);
DFFARX1 I_17706 (I498033,I3563,I304372,I304610,);
DFFARX1 I_17707 (I304610,I3563,I304372,I304627,);
not I_17708 (I304635,I304627);
not I_17709 (I304652,I304610);
nand I_17710 (I304349,I304652,I304471);
nand I_17711 (I304683,I498018,I498024);
and I_17712 (I304700,I304683,I498027);
DFFARX1 I_17713 (I304700,I3563,I304372,I304726,);
nor I_17714 (I304734,I304726,I304398);
DFFARX1 I_17715 (I304734,I3563,I304372,I304337,);
DFFARX1 I_17716 (I304726,I3563,I304372,I304355,);
nor I_17717 (I304779,I498039,I498024);
not I_17718 (I304796,I304779);
nor I_17719 (I304358,I304635,I304796);
nand I_17720 (I304343,I304652,I304796);
nor I_17721 (I304352,I304398,I304779);
DFFARX1 I_17722 (I304779,I3563,I304372,I304361,);
not I_17723 (I304899,I3570);
DFFARX1 I_17724 (I761309,I3563,I304899,I304925,);
nand I_17725 (I304933,I761300,I761315);
and I_17726 (I304950,I304933,I761321);
DFFARX1 I_17727 (I304950,I3563,I304899,I304976,);
nor I_17728 (I304867,I304976,I304925);
not I_17729 (I304998,I304976);
DFFARX1 I_17730 (I761306,I3563,I304899,I305024,);
nand I_17731 (I305032,I305024,I761300);
not I_17732 (I305049,I305032);
DFFARX1 I_17733 (I305049,I3563,I304899,I305075,);
not I_17734 (I304891,I305075);
nor I_17735 (I305097,I304925,I305032);
nor I_17736 (I304873,I304976,I305097);
DFFARX1 I_17737 (I761303,I3563,I304899,I305137,);
DFFARX1 I_17738 (I305137,I3563,I304899,I305154,);
not I_17739 (I305162,I305154);
not I_17740 (I305179,I305137);
nand I_17741 (I304876,I305179,I304998);
nand I_17742 (I305210,I761297,I761312);
and I_17743 (I305227,I305210,I761297);
DFFARX1 I_17744 (I305227,I3563,I304899,I305253,);
nor I_17745 (I305261,I305253,I304925);
DFFARX1 I_17746 (I305261,I3563,I304899,I304864,);
DFFARX1 I_17747 (I305253,I3563,I304899,I304882,);
nor I_17748 (I305306,I761318,I761312);
not I_17749 (I305323,I305306);
nor I_17750 (I304885,I305162,I305323);
nand I_17751 (I304870,I305179,I305323);
nor I_17752 (I304879,I304925,I305306);
DFFARX1 I_17753 (I305306,I3563,I304899,I304888,);
not I_17754 (I305426,I3570);
DFFARX1 I_17755 (I72460,I3563,I305426,I305452,);
nand I_17756 (I305460,I72472,I72481);
and I_17757 (I305477,I305460,I72460);
DFFARX1 I_17758 (I305477,I3563,I305426,I305503,);
nor I_17759 (I305394,I305503,I305452);
not I_17760 (I305525,I305503);
DFFARX1 I_17761 (I72475,I3563,I305426,I305551,);
nand I_17762 (I305559,I305551,I72463);
not I_17763 (I305576,I305559);
DFFARX1 I_17764 (I305576,I3563,I305426,I305602,);
not I_17765 (I305418,I305602);
nor I_17766 (I305624,I305452,I305559);
nor I_17767 (I305400,I305503,I305624);
DFFARX1 I_17768 (I72466,I3563,I305426,I305664,);
DFFARX1 I_17769 (I305664,I3563,I305426,I305681,);
not I_17770 (I305689,I305681);
not I_17771 (I305706,I305664);
nand I_17772 (I305403,I305706,I305525);
nand I_17773 (I305737,I72457,I72457);
and I_17774 (I305754,I305737,I72469);
DFFARX1 I_17775 (I305754,I3563,I305426,I305780,);
nor I_17776 (I305788,I305780,I305452);
DFFARX1 I_17777 (I305788,I3563,I305426,I305391,);
DFFARX1 I_17778 (I305780,I3563,I305426,I305409,);
nor I_17779 (I305833,I72478,I72457);
not I_17780 (I305850,I305833);
nor I_17781 (I305412,I305689,I305850);
nand I_17782 (I305397,I305706,I305850);
nor I_17783 (I305406,I305452,I305833);
DFFARX1 I_17784 (I305833,I3563,I305426,I305415,);
not I_17785 (I305953,I3570);
DFFARX1 I_17786 (I87743,I3563,I305953,I305979,);
nand I_17787 (I305987,I87755,I87764);
and I_17788 (I306004,I305987,I87743);
DFFARX1 I_17789 (I306004,I3563,I305953,I306030,);
nor I_17790 (I305921,I306030,I305979);
not I_17791 (I306052,I306030);
DFFARX1 I_17792 (I87758,I3563,I305953,I306078,);
nand I_17793 (I306086,I306078,I87746);
not I_17794 (I306103,I306086);
DFFARX1 I_17795 (I306103,I3563,I305953,I306129,);
not I_17796 (I305945,I306129);
nor I_17797 (I306151,I305979,I306086);
nor I_17798 (I305927,I306030,I306151);
DFFARX1 I_17799 (I87749,I3563,I305953,I306191,);
DFFARX1 I_17800 (I306191,I3563,I305953,I306208,);
not I_17801 (I306216,I306208);
not I_17802 (I306233,I306191);
nand I_17803 (I305930,I306233,I306052);
nand I_17804 (I306264,I87740,I87740);
and I_17805 (I306281,I306264,I87752);
DFFARX1 I_17806 (I306281,I3563,I305953,I306307,);
nor I_17807 (I306315,I306307,I305979);
DFFARX1 I_17808 (I306315,I3563,I305953,I305918,);
DFFARX1 I_17809 (I306307,I3563,I305953,I305936,);
nor I_17810 (I306360,I87761,I87740);
not I_17811 (I306377,I306360);
nor I_17812 (I305939,I306216,I306377);
nand I_17813 (I305924,I306233,I306377);
nor I_17814 (I305933,I305979,I306360);
DFFARX1 I_17815 (I306360,I3563,I305953,I305942,);
not I_17816 (I306480,I3570);
DFFARX1 I_17817 (I685013,I3563,I306480,I306506,);
nand I_17818 (I306514,I685004,I685019);
and I_17819 (I306531,I306514,I685025);
DFFARX1 I_17820 (I306531,I3563,I306480,I306557,);
nor I_17821 (I306448,I306557,I306506);
not I_17822 (I306579,I306557);
DFFARX1 I_17823 (I685010,I3563,I306480,I306605,);
nand I_17824 (I306613,I306605,I685004);
not I_17825 (I306630,I306613);
DFFARX1 I_17826 (I306630,I3563,I306480,I306656,);
not I_17827 (I306472,I306656);
nor I_17828 (I306678,I306506,I306613);
nor I_17829 (I306454,I306557,I306678);
DFFARX1 I_17830 (I685007,I3563,I306480,I306718,);
DFFARX1 I_17831 (I306718,I3563,I306480,I306735,);
not I_17832 (I306743,I306735);
not I_17833 (I306760,I306718);
nand I_17834 (I306457,I306760,I306579);
nand I_17835 (I306791,I685001,I685016);
and I_17836 (I306808,I306791,I685001);
DFFARX1 I_17837 (I306808,I3563,I306480,I306834,);
nor I_17838 (I306842,I306834,I306506);
DFFARX1 I_17839 (I306842,I3563,I306480,I306445,);
DFFARX1 I_17840 (I306834,I3563,I306480,I306463,);
nor I_17841 (I306887,I685022,I685016);
not I_17842 (I306904,I306887);
nor I_17843 (I306466,I306743,I306904);
nand I_17844 (I306451,I306760,I306904);
nor I_17845 (I306460,I306506,I306887);
DFFARX1 I_17846 (I306887,I3563,I306480,I306469,);
not I_17847 (I307007,I3570);
DFFARX1 I_17848 (I612766,I3563,I307007,I307033,);
nand I_17849 (I307041,I612751,I612754);
and I_17850 (I307058,I307041,I612769);
DFFARX1 I_17851 (I307058,I3563,I307007,I307084,);
nor I_17852 (I306975,I307084,I307033);
not I_17853 (I307106,I307084);
DFFARX1 I_17854 (I612763,I3563,I307007,I307132,);
nand I_17855 (I307140,I307132,I612754);
not I_17856 (I307157,I307140);
DFFARX1 I_17857 (I307157,I3563,I307007,I307183,);
not I_17858 (I306999,I307183);
nor I_17859 (I307205,I307033,I307140);
nor I_17860 (I306981,I307084,I307205);
DFFARX1 I_17861 (I612760,I3563,I307007,I307245,);
DFFARX1 I_17862 (I307245,I3563,I307007,I307262,);
not I_17863 (I307270,I307262);
not I_17864 (I307287,I307245);
nand I_17865 (I306984,I307287,I307106);
nand I_17866 (I307318,I612775,I612751);
and I_17867 (I307335,I307318,I612772);
DFFARX1 I_17868 (I307335,I3563,I307007,I307361,);
nor I_17869 (I307369,I307361,I307033);
DFFARX1 I_17870 (I307369,I3563,I307007,I306972,);
DFFARX1 I_17871 (I307361,I3563,I307007,I306990,);
nor I_17872 (I307414,I612757,I612751);
not I_17873 (I307431,I307414);
nor I_17874 (I306993,I307270,I307431);
nand I_17875 (I306978,I307287,I307431);
nor I_17876 (I306987,I307033,I307414);
DFFARX1 I_17877 (I307414,I3563,I307007,I306996,);
not I_17878 (I307534,I3570);
DFFARX1 I_17879 (I2092,I3563,I307534,I307560,);
nand I_17880 (I307568,I2516,I2332);
and I_17881 (I307585,I307568,I1556);
DFFARX1 I_17882 (I307585,I3563,I307534,I307611,);
nor I_17883 (I307502,I307611,I307560);
not I_17884 (I307633,I307611);
DFFARX1 I_17885 (I3316,I3563,I307534,I307659,);
nand I_17886 (I307667,I307659,I1796);
not I_17887 (I307684,I307667);
DFFARX1 I_17888 (I307684,I3563,I307534,I307710,);
not I_17889 (I307526,I307710);
nor I_17890 (I307732,I307560,I307667);
nor I_17891 (I307508,I307611,I307732);
DFFARX1 I_17892 (I2356,I3563,I307534,I307772,);
DFFARX1 I_17893 (I307772,I3563,I307534,I307789,);
not I_17894 (I307797,I307789);
not I_17895 (I307814,I307772);
nand I_17896 (I307511,I307814,I307633);
nand I_17897 (I307845,I2148,I2452);
and I_17898 (I307862,I307845,I1804);
DFFARX1 I_17899 (I307862,I3563,I307534,I307888,);
nor I_17900 (I307896,I307888,I307560);
DFFARX1 I_17901 (I307896,I3563,I307534,I307499,);
DFFARX1 I_17902 (I307888,I3563,I307534,I307517,);
nor I_17903 (I307941,I1628,I2452);
not I_17904 (I307958,I307941);
nor I_17905 (I307520,I307797,I307958);
nand I_17906 (I307505,I307814,I307958);
nor I_17907 (I307514,I307560,I307941);
DFFARX1 I_17908 (I307941,I3563,I307534,I307523,);
not I_17909 (I308061,I3570);
DFFARX1 I_17910 (I1122207,I3563,I308061,I308087,);
nand I_17911 (I308095,I1122222,I1122207);
and I_17912 (I308112,I308095,I1122225);
DFFARX1 I_17913 (I308112,I3563,I308061,I308138,);
nor I_17914 (I308029,I308138,I308087);
not I_17915 (I308160,I308138);
DFFARX1 I_17916 (I1122231,I3563,I308061,I308186,);
nand I_17917 (I308194,I308186,I1122213);
not I_17918 (I308211,I308194);
DFFARX1 I_17919 (I308211,I3563,I308061,I308237,);
not I_17920 (I308053,I308237);
nor I_17921 (I308259,I308087,I308194);
nor I_17922 (I308035,I308138,I308259);
DFFARX1 I_17923 (I1122210,I3563,I308061,I308299,);
DFFARX1 I_17924 (I308299,I3563,I308061,I308316,);
not I_17925 (I308324,I308316);
not I_17926 (I308341,I308299);
nand I_17927 (I308038,I308341,I308160);
nand I_17928 (I308372,I1122210,I1122216);
and I_17929 (I308389,I308372,I1122228);
DFFARX1 I_17930 (I308389,I3563,I308061,I308415,);
nor I_17931 (I308423,I308415,I308087);
DFFARX1 I_17932 (I308423,I3563,I308061,I308026,);
DFFARX1 I_17933 (I308415,I3563,I308061,I308044,);
nor I_17934 (I308468,I1122219,I1122216);
not I_17935 (I308485,I308468);
nor I_17936 (I308047,I308324,I308485);
nand I_17937 (I308032,I308341,I308485);
nor I_17938 (I308041,I308087,I308468);
DFFARX1 I_17939 (I308468,I3563,I308061,I308050,);
not I_17940 (I308588,I3570);
DFFARX1 I_17941 (I527499,I3563,I308588,I308614,);
nand I_17942 (I308622,I527499,I527511);
and I_17943 (I308639,I308622,I527496);
DFFARX1 I_17944 (I308639,I3563,I308588,I308665,);
nor I_17945 (I308556,I308665,I308614);
not I_17946 (I308687,I308665);
DFFARX1 I_17947 (I527520,I3563,I308588,I308713,);
nand I_17948 (I308721,I308713,I527517);
not I_17949 (I308738,I308721);
DFFARX1 I_17950 (I308738,I3563,I308588,I308764,);
not I_17951 (I308580,I308764);
nor I_17952 (I308786,I308614,I308721);
nor I_17953 (I308562,I308665,I308786);
DFFARX1 I_17954 (I527508,I3563,I308588,I308826,);
DFFARX1 I_17955 (I308826,I3563,I308588,I308843,);
not I_17956 (I308851,I308843);
not I_17957 (I308868,I308826);
nand I_17958 (I308565,I308868,I308687);
nand I_17959 (I308899,I527496,I527505);
and I_17960 (I308916,I308899,I527514);
DFFARX1 I_17961 (I308916,I3563,I308588,I308942,);
nor I_17962 (I308950,I308942,I308614);
DFFARX1 I_17963 (I308950,I3563,I308588,I308553,);
DFFARX1 I_17964 (I308942,I3563,I308588,I308571,);
nor I_17965 (I308995,I527502,I527505);
not I_17966 (I309012,I308995);
nor I_17967 (I308574,I308851,I309012);
nand I_17968 (I308559,I308868,I309012);
nor I_17969 (I308568,I308614,I308995);
DFFARX1 I_17970 (I308995,I3563,I308588,I308577,);
not I_17971 (I309115,I3570);
DFFARX1 I_17972 (I5373,I3563,I309115,I309141,);
nand I_17973 (I309149,I5364,I5367);
and I_17974 (I309166,I309149,I5358);
DFFARX1 I_17975 (I309166,I3563,I309115,I309192,);
nor I_17976 (I309083,I309192,I309141);
not I_17977 (I309214,I309192);
DFFARX1 I_17978 (I5364,I3563,I309115,I309240,);
nand I_17979 (I309248,I309240,I5370);
not I_17980 (I309265,I309248);
DFFARX1 I_17981 (I309265,I3563,I309115,I309291,);
not I_17982 (I309107,I309291);
nor I_17983 (I309313,I309141,I309248);
nor I_17984 (I309089,I309192,I309313);
DFFARX1 I_17985 (I5361,I3563,I309115,I309353,);
DFFARX1 I_17986 (I309353,I3563,I309115,I309370,);
not I_17987 (I309378,I309370);
not I_17988 (I309395,I309353);
nand I_17989 (I309092,I309395,I309214);
nand I_17990 (I309426,I5361,I5376);
and I_17991 (I309443,I309426,I5358);
DFFARX1 I_17992 (I309443,I3563,I309115,I309469,);
nor I_17993 (I309477,I309469,I309141);
DFFARX1 I_17994 (I309477,I3563,I309115,I309080,);
DFFARX1 I_17995 (I309469,I3563,I309115,I309098,);
nor I_17996 (I309522,I5379,I5376);
not I_17997 (I309539,I309522);
nor I_17998 (I309101,I309378,I309539);
nand I_17999 (I309086,I309395,I309539);
nor I_18000 (I309095,I309141,I309522);
DFFARX1 I_18001 (I309522,I3563,I309115,I309104,);
not I_18002 (I309642,I3570);
DFFARX1 I_18003 (I1405924,I3563,I309642,I309668,);
nand I_18004 (I309676,I1405903,I1405903);
and I_18005 (I309693,I309676,I1405930);
DFFARX1 I_18006 (I309693,I3563,I309642,I309719,);
nor I_18007 (I309610,I309719,I309668);
not I_18008 (I309741,I309719);
DFFARX1 I_18009 (I1405918,I3563,I309642,I309767,);
nand I_18010 (I309775,I309767,I1405921);
not I_18011 (I309792,I309775);
DFFARX1 I_18012 (I309792,I3563,I309642,I309818,);
not I_18013 (I309634,I309818);
nor I_18014 (I309840,I309668,I309775);
nor I_18015 (I309616,I309719,I309840);
DFFARX1 I_18016 (I1405912,I3563,I309642,I309880,);
DFFARX1 I_18017 (I309880,I3563,I309642,I309897,);
not I_18018 (I309905,I309897);
not I_18019 (I309922,I309880);
nand I_18020 (I309619,I309922,I309741);
nand I_18021 (I309953,I1405909,I1405906);
and I_18022 (I309970,I309953,I1405927);
DFFARX1 I_18023 (I309970,I3563,I309642,I309996,);
nor I_18024 (I310004,I309996,I309668);
DFFARX1 I_18025 (I310004,I3563,I309642,I309607,);
DFFARX1 I_18026 (I309996,I3563,I309642,I309625,);
nor I_18027 (I310049,I1405915,I1405906);
not I_18028 (I310066,I310049);
nor I_18029 (I309628,I309905,I310066);
nand I_18030 (I309613,I309922,I310066);
nor I_18031 (I309622,I309668,I310049);
DFFARX1 I_18032 (I310049,I3563,I309642,I309631,);
not I_18033 (I310169,I3570);
DFFARX1 I_18034 (I100918,I3563,I310169,I310195,);
nand I_18035 (I310203,I100930,I100939);
and I_18036 (I310220,I310203,I100918);
DFFARX1 I_18037 (I310220,I3563,I310169,I310246,);
nor I_18038 (I310137,I310246,I310195);
not I_18039 (I310268,I310246);
DFFARX1 I_18040 (I100933,I3563,I310169,I310294,);
nand I_18041 (I310302,I310294,I100921);
not I_18042 (I310319,I310302);
DFFARX1 I_18043 (I310319,I3563,I310169,I310345,);
not I_18044 (I310161,I310345);
nor I_18045 (I310367,I310195,I310302);
nor I_18046 (I310143,I310246,I310367);
DFFARX1 I_18047 (I100924,I3563,I310169,I310407,);
DFFARX1 I_18048 (I310407,I3563,I310169,I310424,);
not I_18049 (I310432,I310424);
not I_18050 (I310449,I310407);
nand I_18051 (I310146,I310449,I310268);
nand I_18052 (I310480,I100915,I100915);
and I_18053 (I310497,I310480,I100927);
DFFARX1 I_18054 (I310497,I3563,I310169,I310523,);
nor I_18055 (I310531,I310523,I310195);
DFFARX1 I_18056 (I310531,I3563,I310169,I310134,);
DFFARX1 I_18057 (I310523,I3563,I310169,I310152,);
nor I_18058 (I310576,I100936,I100915);
not I_18059 (I310593,I310576);
nor I_18060 (I310155,I310432,I310593);
nand I_18061 (I310140,I310449,I310593);
nor I_18062 (I310149,I310195,I310576);
DFFARX1 I_18063 (I310576,I3563,I310169,I310158,);
not I_18064 (I310696,I3570);
DFFARX1 I_18065 (I659581,I3563,I310696,I310722,);
nand I_18066 (I310730,I659572,I659587);
and I_18067 (I310747,I310730,I659593);
DFFARX1 I_18068 (I310747,I3563,I310696,I310773,);
nor I_18069 (I310664,I310773,I310722);
not I_18070 (I310795,I310773);
DFFARX1 I_18071 (I659578,I3563,I310696,I310821,);
nand I_18072 (I310829,I310821,I659572);
not I_18073 (I310846,I310829);
DFFARX1 I_18074 (I310846,I3563,I310696,I310872,);
not I_18075 (I310688,I310872);
nor I_18076 (I310894,I310722,I310829);
nor I_18077 (I310670,I310773,I310894);
DFFARX1 I_18078 (I659575,I3563,I310696,I310934,);
DFFARX1 I_18079 (I310934,I3563,I310696,I310951,);
not I_18080 (I310959,I310951);
not I_18081 (I310976,I310934);
nand I_18082 (I310673,I310976,I310795);
nand I_18083 (I311007,I659569,I659584);
and I_18084 (I311024,I311007,I659569);
DFFARX1 I_18085 (I311024,I3563,I310696,I311050,);
nor I_18086 (I311058,I311050,I310722);
DFFARX1 I_18087 (I311058,I3563,I310696,I310661,);
DFFARX1 I_18088 (I311050,I3563,I310696,I310679,);
nor I_18089 (I311103,I659590,I659584);
not I_18090 (I311120,I311103);
nor I_18091 (I310682,I310959,I311120);
nand I_18092 (I310667,I310976,I311120);
nor I_18093 (I310676,I310722,I311103);
DFFARX1 I_18094 (I311103,I3563,I310696,I310685,);
not I_18095 (I311223,I3570);
DFFARX1 I_18096 (I879042,I3563,I311223,I311249,);
nand I_18097 (I311257,I879045,I879039);
and I_18098 (I311274,I311257,I879051);
DFFARX1 I_18099 (I311274,I3563,I311223,I311300,);
nor I_18100 (I311191,I311300,I311249);
not I_18101 (I311322,I311300);
DFFARX1 I_18102 (I879054,I3563,I311223,I311348,);
nand I_18103 (I311356,I311348,I879045);
not I_18104 (I311373,I311356);
DFFARX1 I_18105 (I311373,I3563,I311223,I311399,);
not I_18106 (I311215,I311399);
nor I_18107 (I311421,I311249,I311356);
nor I_18108 (I311197,I311300,I311421);
DFFARX1 I_18109 (I879057,I3563,I311223,I311461,);
DFFARX1 I_18110 (I311461,I3563,I311223,I311478,);
not I_18111 (I311486,I311478);
not I_18112 (I311503,I311461);
nand I_18113 (I311200,I311503,I311322);
nand I_18114 (I311534,I879039,I879048);
and I_18115 (I311551,I311534,I879042);
DFFARX1 I_18116 (I311551,I3563,I311223,I311577,);
nor I_18117 (I311585,I311577,I311249);
DFFARX1 I_18118 (I311585,I3563,I311223,I311188,);
DFFARX1 I_18119 (I311577,I3563,I311223,I311206,);
nor I_18120 (I311630,I879060,I879048);
not I_18121 (I311647,I311630);
nor I_18122 (I311209,I311486,I311647);
nand I_18123 (I311194,I311503,I311647);
nor I_18124 (I311203,I311249,I311630);
DFFARX1 I_18125 (I311630,I3563,I311223,I311212,);
not I_18126 (I311750,I3570);
DFFARX1 I_18127 (I1103711,I3563,I311750,I311776,);
nand I_18128 (I311784,I1103726,I1103711);
and I_18129 (I311801,I311784,I1103729);
DFFARX1 I_18130 (I311801,I3563,I311750,I311827,);
nor I_18131 (I311718,I311827,I311776);
not I_18132 (I311849,I311827);
DFFARX1 I_18133 (I1103735,I3563,I311750,I311875,);
nand I_18134 (I311883,I311875,I1103717);
not I_18135 (I311900,I311883);
DFFARX1 I_18136 (I311900,I3563,I311750,I311926,);
not I_18137 (I311742,I311926);
nor I_18138 (I311948,I311776,I311883);
nor I_18139 (I311724,I311827,I311948);
DFFARX1 I_18140 (I1103714,I3563,I311750,I311988,);
DFFARX1 I_18141 (I311988,I3563,I311750,I312005,);
not I_18142 (I312013,I312005);
not I_18143 (I312030,I311988);
nand I_18144 (I311727,I312030,I311849);
nand I_18145 (I312061,I1103714,I1103720);
and I_18146 (I312078,I312061,I1103732);
DFFARX1 I_18147 (I312078,I3563,I311750,I312104,);
nor I_18148 (I312112,I312104,I311776);
DFFARX1 I_18149 (I312112,I3563,I311750,I311715,);
DFFARX1 I_18150 (I312104,I3563,I311750,I311733,);
nor I_18151 (I312157,I1103723,I1103720);
not I_18152 (I312174,I312157);
nor I_18153 (I311736,I312013,I312174);
nand I_18154 (I311721,I312030,I312174);
nor I_18155 (I311730,I311776,I312157);
DFFARX1 I_18156 (I312157,I3563,I311750,I311739,);
not I_18157 (I312277,I3570);
DFFARX1 I_18158 (I18176,I3563,I312277,I312303,);
nand I_18159 (I312311,I18200,I18179);
and I_18160 (I312328,I312311,I18176);
DFFARX1 I_18161 (I312328,I3563,I312277,I312354,);
nor I_18162 (I312245,I312354,I312303);
not I_18163 (I312376,I312354);
DFFARX1 I_18164 (I18182,I3563,I312277,I312402,);
nand I_18165 (I312410,I312402,I18191);
not I_18166 (I312427,I312410);
DFFARX1 I_18167 (I312427,I3563,I312277,I312453,);
not I_18168 (I312269,I312453);
nor I_18169 (I312475,I312303,I312410);
nor I_18170 (I312251,I312354,I312475);
DFFARX1 I_18171 (I18185,I3563,I312277,I312515,);
DFFARX1 I_18172 (I312515,I3563,I312277,I312532,);
not I_18173 (I312540,I312532);
not I_18174 (I312557,I312515);
nand I_18175 (I312254,I312557,I312376);
nand I_18176 (I312588,I18197,I18179);
and I_18177 (I312605,I312588,I18188);
DFFARX1 I_18178 (I312605,I3563,I312277,I312631,);
nor I_18179 (I312639,I312631,I312303);
DFFARX1 I_18180 (I312639,I3563,I312277,I312242,);
DFFARX1 I_18181 (I312631,I3563,I312277,I312260,);
nor I_18182 (I312684,I18194,I18179);
not I_18183 (I312701,I312684);
nor I_18184 (I312263,I312540,I312701);
nand I_18185 (I312248,I312557,I312701);
nor I_18186 (I312257,I312303,I312684);
DFFARX1 I_18187 (I312684,I3563,I312277,I312266,);
not I_18188 (I312804,I3570);
DFFARX1 I_18189 (I637620,I3563,I312804,I312830,);
nand I_18190 (I312838,I637605,I637608);
and I_18191 (I312855,I312838,I637623);
DFFARX1 I_18192 (I312855,I3563,I312804,I312881,);
nor I_18193 (I312772,I312881,I312830);
not I_18194 (I312903,I312881);
DFFARX1 I_18195 (I637617,I3563,I312804,I312929,);
nand I_18196 (I312937,I312929,I637608);
not I_18197 (I312954,I312937);
DFFARX1 I_18198 (I312954,I3563,I312804,I312980,);
not I_18199 (I312796,I312980);
nor I_18200 (I313002,I312830,I312937);
nor I_18201 (I312778,I312881,I313002);
DFFARX1 I_18202 (I637614,I3563,I312804,I313042,);
DFFARX1 I_18203 (I313042,I3563,I312804,I313059,);
not I_18204 (I313067,I313059);
not I_18205 (I313084,I313042);
nand I_18206 (I312781,I313084,I312903);
nand I_18207 (I313115,I637629,I637605);
and I_18208 (I313132,I313115,I637626);
DFFARX1 I_18209 (I313132,I3563,I312804,I313158,);
nor I_18210 (I313166,I313158,I312830);
DFFARX1 I_18211 (I313166,I3563,I312804,I312769,);
DFFARX1 I_18212 (I313158,I3563,I312804,I312787,);
nor I_18213 (I313211,I637611,I637605);
not I_18214 (I313228,I313211);
nor I_18215 (I312790,I313067,I313228);
nand I_18216 (I312775,I313084,I313228);
nor I_18217 (I312784,I312830,I313211);
DFFARX1 I_18218 (I313211,I3563,I312804,I312793,);
not I_18219 (I313331,I3570);
DFFARX1 I_18220 (I984646,I3563,I313331,I313357,);
nand I_18221 (I313365,I984643,I984661);
and I_18222 (I313382,I313365,I984652);
DFFARX1 I_18223 (I313382,I3563,I313331,I313408,);
nor I_18224 (I313299,I313408,I313357);
not I_18225 (I313430,I313408);
DFFARX1 I_18226 (I984667,I3563,I313331,I313456,);
nand I_18227 (I313464,I313456,I984649);
not I_18228 (I313481,I313464);
DFFARX1 I_18229 (I313481,I3563,I313331,I313507,);
not I_18230 (I313323,I313507);
nor I_18231 (I313529,I313357,I313464);
nor I_18232 (I313305,I313408,I313529);
DFFARX1 I_18233 (I984655,I3563,I313331,I313569,);
DFFARX1 I_18234 (I313569,I3563,I313331,I313586,);
not I_18235 (I313594,I313586);
not I_18236 (I313611,I313569);
nand I_18237 (I313308,I313611,I313430);
nand I_18238 (I313642,I984643,I984670);
and I_18239 (I313659,I313642,I984658);
DFFARX1 I_18240 (I313659,I3563,I313331,I313685,);
nor I_18241 (I313693,I313685,I313357);
DFFARX1 I_18242 (I313693,I3563,I313331,I313296,);
DFFARX1 I_18243 (I313685,I3563,I313331,I313314,);
nor I_18244 (I313738,I984664,I984670);
not I_18245 (I313755,I313738);
nor I_18246 (I313317,I313594,I313755);
nand I_18247 (I313302,I313611,I313755);
nor I_18248 (I313311,I313357,I313738);
DFFARX1 I_18249 (I313738,I3563,I313331,I313320,);
not I_18250 (I313858,I3570);
DFFARX1 I_18251 (I279738,I3563,I313858,I313884,);
nand I_18252 (I313892,I279738,I279744);
and I_18253 (I313909,I313892,I279762);
DFFARX1 I_18254 (I313909,I3563,I313858,I313935,);
nor I_18255 (I313826,I313935,I313884);
not I_18256 (I313957,I313935);
DFFARX1 I_18257 (I279750,I3563,I313858,I313983,);
nand I_18258 (I313991,I313983,I279747);
not I_18259 (I314008,I313991);
DFFARX1 I_18260 (I314008,I3563,I313858,I314034,);
not I_18261 (I313850,I314034);
nor I_18262 (I314056,I313884,I313991);
nor I_18263 (I313832,I313935,I314056);
DFFARX1 I_18264 (I279756,I3563,I313858,I314096,);
DFFARX1 I_18265 (I314096,I3563,I313858,I314113,);
not I_18266 (I314121,I314113);
not I_18267 (I314138,I314096);
nand I_18268 (I313835,I314138,I313957);
nand I_18269 (I314169,I279741,I279741);
and I_18270 (I314186,I314169,I279753);
DFFARX1 I_18271 (I314186,I3563,I313858,I314212,);
nor I_18272 (I314220,I314212,I313884);
DFFARX1 I_18273 (I314220,I3563,I313858,I313823,);
DFFARX1 I_18274 (I314212,I3563,I313858,I313841,);
nor I_18275 (I314265,I279759,I279741);
not I_18276 (I314282,I314265);
nor I_18277 (I313844,I314121,I314282);
nand I_18278 (I313829,I314138,I314282);
nor I_18279 (I313838,I313884,I314265);
DFFARX1 I_18280 (I314265,I3563,I313858,I313847,);
not I_18281 (I314385,I3570);
DFFARX1 I_18282 (I495310,I3563,I314385,I314411,);
nand I_18283 (I314419,I495322,I495301);
and I_18284 (I314436,I314419,I495325);
DFFARX1 I_18285 (I314436,I3563,I314385,I314462,);
nor I_18286 (I314353,I314462,I314411);
not I_18287 (I314484,I314462);
DFFARX1 I_18288 (I495316,I3563,I314385,I314510,);
nand I_18289 (I314518,I314510,I495298);
not I_18290 (I314535,I314518);
DFFARX1 I_18291 (I314535,I3563,I314385,I314561,);
not I_18292 (I314377,I314561);
nor I_18293 (I314583,I314411,I314518);
nor I_18294 (I314359,I314462,I314583);
DFFARX1 I_18295 (I495313,I3563,I314385,I314623,);
DFFARX1 I_18296 (I314623,I3563,I314385,I314640,);
not I_18297 (I314648,I314640);
not I_18298 (I314665,I314623);
nand I_18299 (I314362,I314665,I314484);
nand I_18300 (I314696,I495298,I495304);
and I_18301 (I314713,I314696,I495307);
DFFARX1 I_18302 (I314713,I3563,I314385,I314739,);
nor I_18303 (I314747,I314739,I314411);
DFFARX1 I_18304 (I314747,I3563,I314385,I314350,);
DFFARX1 I_18305 (I314739,I3563,I314385,I314368,);
nor I_18306 (I314792,I495319,I495304);
not I_18307 (I314809,I314792);
nor I_18308 (I314371,I314648,I314809);
nand I_18309 (I314356,I314665,I314809);
nor I_18310 (I314365,I314411,I314792);
DFFARX1 I_18311 (I314792,I3563,I314385,I314374,);
not I_18312 (I314912,I3570);
DFFARX1 I_18313 (I1168447,I3563,I314912,I314938,);
nand I_18314 (I314946,I1168462,I1168447);
and I_18315 (I314963,I314946,I1168465);
DFFARX1 I_18316 (I314963,I3563,I314912,I314989,);
nor I_18317 (I314880,I314989,I314938);
not I_18318 (I315011,I314989);
DFFARX1 I_18319 (I1168471,I3563,I314912,I315037,);
nand I_18320 (I315045,I315037,I1168453);
not I_18321 (I315062,I315045);
DFFARX1 I_18322 (I315062,I3563,I314912,I315088,);
not I_18323 (I314904,I315088);
nor I_18324 (I315110,I314938,I315045);
nor I_18325 (I314886,I314989,I315110);
DFFARX1 I_18326 (I1168450,I3563,I314912,I315150,);
DFFARX1 I_18327 (I315150,I3563,I314912,I315167,);
not I_18328 (I315175,I315167);
not I_18329 (I315192,I315150);
nand I_18330 (I314889,I315192,I315011);
nand I_18331 (I315223,I1168450,I1168456);
and I_18332 (I315240,I315223,I1168468);
DFFARX1 I_18333 (I315240,I3563,I314912,I315266,);
nor I_18334 (I315274,I315266,I314938);
DFFARX1 I_18335 (I315274,I3563,I314912,I314877,);
DFFARX1 I_18336 (I315266,I3563,I314912,I314895,);
nor I_18337 (I315319,I1168459,I1168456);
not I_18338 (I315336,I315319);
nor I_18339 (I314898,I315175,I315336);
nand I_18340 (I314883,I315192,I315336);
nor I_18341 (I314892,I314938,I315319);
DFFARX1 I_18342 (I315319,I3563,I314912,I314901,);
not I_18343 (I315439,I3570);
DFFARX1 I_18344 (I947824,I3563,I315439,I315465,);
nand I_18345 (I315473,I947821,I947839);
and I_18346 (I315490,I315473,I947830);
DFFARX1 I_18347 (I315490,I3563,I315439,I315516,);
nor I_18348 (I315407,I315516,I315465);
not I_18349 (I315538,I315516);
DFFARX1 I_18350 (I947845,I3563,I315439,I315564,);
nand I_18351 (I315572,I315564,I947827);
not I_18352 (I315589,I315572);
DFFARX1 I_18353 (I315589,I3563,I315439,I315615,);
not I_18354 (I315431,I315615);
nor I_18355 (I315637,I315465,I315572);
nor I_18356 (I315413,I315516,I315637);
DFFARX1 I_18357 (I947833,I3563,I315439,I315677,);
DFFARX1 I_18358 (I315677,I3563,I315439,I315694,);
not I_18359 (I315702,I315694);
not I_18360 (I315719,I315677);
nand I_18361 (I315416,I315719,I315538);
nand I_18362 (I315750,I947821,I947848);
and I_18363 (I315767,I315750,I947836);
DFFARX1 I_18364 (I315767,I3563,I315439,I315793,);
nor I_18365 (I315801,I315793,I315465);
DFFARX1 I_18366 (I315801,I3563,I315439,I315404,);
DFFARX1 I_18367 (I315793,I3563,I315439,I315422,);
nor I_18368 (I315846,I947842,I947848);
not I_18369 (I315863,I315846);
nor I_18370 (I315425,I315702,I315863);
nand I_18371 (I315410,I315719,I315863);
nor I_18372 (I315419,I315465,I315846);
DFFARX1 I_18373 (I315846,I3563,I315439,I315428,);
not I_18374 (I315966,I3570);
DFFARX1 I_18375 (I847422,I3563,I315966,I315992,);
nand I_18376 (I316000,I847425,I847419);
and I_18377 (I316017,I316000,I847431);
DFFARX1 I_18378 (I316017,I3563,I315966,I316043,);
nor I_18379 (I315934,I316043,I315992);
not I_18380 (I316065,I316043);
DFFARX1 I_18381 (I847434,I3563,I315966,I316091,);
nand I_18382 (I316099,I316091,I847425);
not I_18383 (I316116,I316099);
DFFARX1 I_18384 (I316116,I3563,I315966,I316142,);
not I_18385 (I315958,I316142);
nor I_18386 (I316164,I315992,I316099);
nor I_18387 (I315940,I316043,I316164);
DFFARX1 I_18388 (I847437,I3563,I315966,I316204,);
DFFARX1 I_18389 (I316204,I3563,I315966,I316221,);
not I_18390 (I316229,I316221);
not I_18391 (I316246,I316204);
nand I_18392 (I315943,I316246,I316065);
nand I_18393 (I316277,I847419,I847428);
and I_18394 (I316294,I316277,I847422);
DFFARX1 I_18395 (I316294,I3563,I315966,I316320,);
nor I_18396 (I316328,I316320,I315992);
DFFARX1 I_18397 (I316328,I3563,I315966,I315931,);
DFFARX1 I_18398 (I316320,I3563,I315966,I315949,);
nor I_18399 (I316373,I847440,I847428);
not I_18400 (I316390,I316373);
nor I_18401 (I315952,I316229,I316390);
nand I_18402 (I315937,I316246,I316390);
nor I_18403 (I315946,I315992,I316373);
DFFARX1 I_18404 (I316373,I3563,I315966,I315955,);
not I_18405 (I316493,I3570);
DFFARX1 I_18406 (I954284,I3563,I316493,I316519,);
nand I_18407 (I316527,I954281,I954299);
and I_18408 (I316544,I316527,I954290);
DFFARX1 I_18409 (I316544,I3563,I316493,I316570,);
nor I_18410 (I316461,I316570,I316519);
not I_18411 (I316592,I316570);
DFFARX1 I_18412 (I954305,I3563,I316493,I316618,);
nand I_18413 (I316626,I316618,I954287);
not I_18414 (I316643,I316626);
DFFARX1 I_18415 (I316643,I3563,I316493,I316669,);
not I_18416 (I316485,I316669);
nor I_18417 (I316691,I316519,I316626);
nor I_18418 (I316467,I316570,I316691);
DFFARX1 I_18419 (I954293,I3563,I316493,I316731,);
DFFARX1 I_18420 (I316731,I3563,I316493,I316748,);
not I_18421 (I316756,I316748);
not I_18422 (I316773,I316731);
nand I_18423 (I316470,I316773,I316592);
nand I_18424 (I316804,I954281,I954308);
and I_18425 (I316821,I316804,I954296);
DFFARX1 I_18426 (I316821,I3563,I316493,I316847,);
nor I_18427 (I316855,I316847,I316519);
DFFARX1 I_18428 (I316855,I3563,I316493,I316458,);
DFFARX1 I_18429 (I316847,I3563,I316493,I316476,);
nor I_18430 (I316900,I954302,I954308);
not I_18431 (I316917,I316900);
nor I_18432 (I316479,I316756,I316917);
nand I_18433 (I316464,I316773,I316917);
nor I_18434 (I316473,I316519,I316900);
DFFARX1 I_18435 (I316900,I3563,I316493,I316482,);
not I_18436 (I317020,I3570);
DFFARX1 I_18437 (I875880,I3563,I317020,I317046,);
nand I_18438 (I317054,I875883,I875877);
and I_18439 (I317071,I317054,I875889);
DFFARX1 I_18440 (I317071,I3563,I317020,I317097,);
nor I_18441 (I316988,I317097,I317046);
not I_18442 (I317119,I317097);
DFFARX1 I_18443 (I875892,I3563,I317020,I317145,);
nand I_18444 (I317153,I317145,I875883);
not I_18445 (I317170,I317153);
DFFARX1 I_18446 (I317170,I3563,I317020,I317196,);
not I_18447 (I317012,I317196);
nor I_18448 (I317218,I317046,I317153);
nor I_18449 (I316994,I317097,I317218);
DFFARX1 I_18450 (I875895,I3563,I317020,I317258,);
DFFARX1 I_18451 (I317258,I3563,I317020,I317275,);
not I_18452 (I317283,I317275);
not I_18453 (I317300,I317258);
nand I_18454 (I316997,I317300,I317119);
nand I_18455 (I317331,I875877,I875886);
and I_18456 (I317348,I317331,I875880);
DFFARX1 I_18457 (I317348,I3563,I317020,I317374,);
nor I_18458 (I317382,I317374,I317046);
DFFARX1 I_18459 (I317382,I3563,I317020,I316985,);
DFFARX1 I_18460 (I317374,I3563,I317020,I317003,);
nor I_18461 (I317427,I875898,I875886);
not I_18462 (I317444,I317427);
nor I_18463 (I317006,I317283,I317444);
nand I_18464 (I316991,I317300,I317444);
nor I_18465 (I317000,I317046,I317427);
DFFARX1 I_18466 (I317427,I3563,I317020,I317009,);
not I_18467 (I317547,I3570);
DFFARX1 I_18468 (I1006610,I3563,I317547,I317573,);
nand I_18469 (I317581,I1006607,I1006625);
and I_18470 (I317598,I317581,I1006616);
DFFARX1 I_18471 (I317598,I3563,I317547,I317624,);
nor I_18472 (I317515,I317624,I317573);
not I_18473 (I317646,I317624);
DFFARX1 I_18474 (I1006631,I3563,I317547,I317672,);
nand I_18475 (I317680,I317672,I1006613);
not I_18476 (I317697,I317680);
DFFARX1 I_18477 (I317697,I3563,I317547,I317723,);
not I_18478 (I317539,I317723);
nor I_18479 (I317745,I317573,I317680);
nor I_18480 (I317521,I317624,I317745);
DFFARX1 I_18481 (I1006619,I3563,I317547,I317785,);
DFFARX1 I_18482 (I317785,I3563,I317547,I317802,);
not I_18483 (I317810,I317802);
not I_18484 (I317827,I317785);
nand I_18485 (I317524,I317827,I317646);
nand I_18486 (I317858,I1006607,I1006634);
and I_18487 (I317875,I317858,I1006622);
DFFARX1 I_18488 (I317875,I3563,I317547,I317901,);
nor I_18489 (I317909,I317901,I317573);
DFFARX1 I_18490 (I317909,I3563,I317547,I317512,);
DFFARX1 I_18491 (I317901,I3563,I317547,I317530,);
nor I_18492 (I317954,I1006628,I1006634);
not I_18493 (I317971,I317954);
nor I_18494 (I317533,I317810,I317971);
nand I_18495 (I317518,I317827,I317971);
nor I_18496 (I317527,I317573,I317954);
DFFARX1 I_18497 (I317954,I3563,I317547,I317536,);
not I_18498 (I318074,I3570);
DFFARX1 I_18499 (I23446,I3563,I318074,I318100,);
nand I_18500 (I318108,I23470,I23449);
and I_18501 (I318125,I318108,I23446);
DFFARX1 I_18502 (I318125,I3563,I318074,I318151,);
nor I_18503 (I318042,I318151,I318100);
not I_18504 (I318173,I318151);
DFFARX1 I_18505 (I23452,I3563,I318074,I318199,);
nand I_18506 (I318207,I318199,I23461);
not I_18507 (I318224,I318207);
DFFARX1 I_18508 (I318224,I3563,I318074,I318250,);
not I_18509 (I318066,I318250);
nor I_18510 (I318272,I318100,I318207);
nor I_18511 (I318048,I318151,I318272);
DFFARX1 I_18512 (I23455,I3563,I318074,I318312,);
DFFARX1 I_18513 (I318312,I3563,I318074,I318329,);
not I_18514 (I318337,I318329);
not I_18515 (I318354,I318312);
nand I_18516 (I318051,I318354,I318173);
nand I_18517 (I318385,I23467,I23449);
and I_18518 (I318402,I318385,I23458);
DFFARX1 I_18519 (I318402,I3563,I318074,I318428,);
nor I_18520 (I318436,I318428,I318100);
DFFARX1 I_18521 (I318436,I3563,I318074,I318039,);
DFFARX1 I_18522 (I318428,I3563,I318074,I318057,);
nor I_18523 (I318481,I23464,I23449);
not I_18524 (I318498,I318481);
nor I_18525 (I318060,I318337,I318498);
nand I_18526 (I318045,I318354,I318498);
nor I_18527 (I318054,I318100,I318481);
DFFARX1 I_18528 (I318481,I3563,I318074,I318063,);
not I_18529 (I318601,I3570);
DFFARX1 I_18530 (I1366654,I3563,I318601,I318627,);
nand I_18531 (I318635,I1366633,I1366633);
and I_18532 (I318652,I318635,I1366660);
DFFARX1 I_18533 (I318652,I3563,I318601,I318678,);
nor I_18534 (I318569,I318678,I318627);
not I_18535 (I318700,I318678);
DFFARX1 I_18536 (I1366648,I3563,I318601,I318726,);
nand I_18537 (I318734,I318726,I1366651);
not I_18538 (I318751,I318734);
DFFARX1 I_18539 (I318751,I3563,I318601,I318777,);
not I_18540 (I318593,I318777);
nor I_18541 (I318799,I318627,I318734);
nor I_18542 (I318575,I318678,I318799);
DFFARX1 I_18543 (I1366642,I3563,I318601,I318839,);
DFFARX1 I_18544 (I318839,I3563,I318601,I318856,);
not I_18545 (I318864,I318856);
not I_18546 (I318881,I318839);
nand I_18547 (I318578,I318881,I318700);
nand I_18548 (I318912,I1366639,I1366636);
and I_18549 (I318929,I318912,I1366657);
DFFARX1 I_18550 (I318929,I3563,I318601,I318955,);
nor I_18551 (I318963,I318955,I318627);
DFFARX1 I_18552 (I318963,I3563,I318601,I318566,);
DFFARX1 I_18553 (I318955,I3563,I318601,I318584,);
nor I_18554 (I319008,I1366645,I1366636);
not I_18555 (I319025,I319008);
nor I_18556 (I318587,I318864,I319025);
nand I_18557 (I318572,I318881,I319025);
nor I_18558 (I318581,I318627,I319008);
DFFARX1 I_18559 (I319008,I3563,I318601,I318590,);
not I_18560 (I319128,I3570);
DFFARX1 I_18561 (I14298,I3563,I319128,I319154,);
nand I_18562 (I319162,I14289,I14292);
and I_18563 (I319179,I319162,I14283);
DFFARX1 I_18564 (I319179,I3563,I319128,I319205,);
nor I_18565 (I319096,I319205,I319154);
not I_18566 (I319227,I319205);
DFFARX1 I_18567 (I14289,I3563,I319128,I319253,);
nand I_18568 (I319261,I319253,I14295);
not I_18569 (I319278,I319261);
DFFARX1 I_18570 (I319278,I3563,I319128,I319304,);
not I_18571 (I319120,I319304);
nor I_18572 (I319326,I319154,I319261);
nor I_18573 (I319102,I319205,I319326);
DFFARX1 I_18574 (I14286,I3563,I319128,I319366,);
DFFARX1 I_18575 (I319366,I3563,I319128,I319383,);
not I_18576 (I319391,I319383);
not I_18577 (I319408,I319366);
nand I_18578 (I319105,I319408,I319227);
nand I_18579 (I319439,I14286,I14301);
and I_18580 (I319456,I319439,I14283);
DFFARX1 I_18581 (I319456,I3563,I319128,I319482,);
nor I_18582 (I319490,I319482,I319154);
DFFARX1 I_18583 (I319490,I3563,I319128,I319093,);
DFFARX1 I_18584 (I319482,I3563,I319128,I319111,);
nor I_18585 (I319535,I14304,I14301);
not I_18586 (I319552,I319535);
nor I_18587 (I319114,I319391,I319552);
nand I_18588 (I319099,I319408,I319552);
nor I_18589 (I319108,I319154,I319535);
DFFARX1 I_18590 (I319535,I3563,I319128,I319117,);
not I_18591 (I319655,I3570);
DFFARX1 I_18592 (I932966,I3563,I319655,I319681,);
nand I_18593 (I319689,I932963,I932981);
and I_18594 (I319706,I319689,I932972);
DFFARX1 I_18595 (I319706,I3563,I319655,I319732,);
nor I_18596 (I319623,I319732,I319681);
not I_18597 (I319754,I319732);
DFFARX1 I_18598 (I932987,I3563,I319655,I319780,);
nand I_18599 (I319788,I319780,I932969);
not I_18600 (I319805,I319788);
DFFARX1 I_18601 (I319805,I3563,I319655,I319831,);
not I_18602 (I319647,I319831);
nor I_18603 (I319853,I319681,I319788);
nor I_18604 (I319629,I319732,I319853);
DFFARX1 I_18605 (I932975,I3563,I319655,I319893,);
DFFARX1 I_18606 (I319893,I3563,I319655,I319910,);
not I_18607 (I319918,I319910);
not I_18608 (I319935,I319893);
nand I_18609 (I319632,I319935,I319754);
nand I_18610 (I319966,I932963,I932990);
and I_18611 (I319983,I319966,I932978);
DFFARX1 I_18612 (I319983,I3563,I319655,I320009,);
nor I_18613 (I320017,I320009,I319681);
DFFARX1 I_18614 (I320017,I3563,I319655,I319620,);
DFFARX1 I_18615 (I320009,I3563,I319655,I319638,);
nor I_18616 (I320062,I932984,I932990);
not I_18617 (I320079,I320062);
nor I_18618 (I319641,I319918,I320079);
nand I_18619 (I319626,I319935,I320079);
nor I_18620 (I319635,I319681,I320062);
DFFARX1 I_18621 (I320062,I3563,I319655,I319644,);
not I_18622 (I320182,I3570);
DFFARX1 I_18623 (I258913,I3563,I320182,I320208,);
nand I_18624 (I320216,I258913,I258919);
and I_18625 (I320233,I320216,I258937);
DFFARX1 I_18626 (I320233,I3563,I320182,I320259,);
nor I_18627 (I320150,I320259,I320208);
not I_18628 (I320281,I320259);
DFFARX1 I_18629 (I258925,I3563,I320182,I320307,);
nand I_18630 (I320315,I320307,I258922);
not I_18631 (I320332,I320315);
DFFARX1 I_18632 (I320332,I3563,I320182,I320358,);
not I_18633 (I320174,I320358);
nor I_18634 (I320380,I320208,I320315);
nor I_18635 (I320156,I320259,I320380);
DFFARX1 I_18636 (I258931,I3563,I320182,I320420,);
DFFARX1 I_18637 (I320420,I3563,I320182,I320437,);
not I_18638 (I320445,I320437);
not I_18639 (I320462,I320420);
nand I_18640 (I320159,I320462,I320281);
nand I_18641 (I320493,I258916,I258916);
and I_18642 (I320510,I320493,I258928);
DFFARX1 I_18643 (I320510,I3563,I320182,I320536,);
nor I_18644 (I320544,I320536,I320208);
DFFARX1 I_18645 (I320544,I3563,I320182,I320147,);
DFFARX1 I_18646 (I320536,I3563,I320182,I320165,);
nor I_18647 (I320589,I258934,I258916);
not I_18648 (I320606,I320589);
nor I_18649 (I320168,I320445,I320606);
nand I_18650 (I320153,I320462,I320606);
nor I_18651 (I320162,I320208,I320589);
DFFARX1 I_18652 (I320589,I3563,I320182,I320171,);
not I_18653 (I320709,I3570);
DFFARX1 I_18654 (I616234,I3563,I320709,I320735,);
nand I_18655 (I320743,I616219,I616222);
and I_18656 (I320760,I320743,I616237);
DFFARX1 I_18657 (I320760,I3563,I320709,I320786,);
nor I_18658 (I320677,I320786,I320735);
not I_18659 (I320808,I320786);
DFFARX1 I_18660 (I616231,I3563,I320709,I320834,);
nand I_18661 (I320842,I320834,I616222);
not I_18662 (I320859,I320842);
DFFARX1 I_18663 (I320859,I3563,I320709,I320885,);
not I_18664 (I320701,I320885);
nor I_18665 (I320907,I320735,I320842);
nor I_18666 (I320683,I320786,I320907);
DFFARX1 I_18667 (I616228,I3563,I320709,I320947,);
DFFARX1 I_18668 (I320947,I3563,I320709,I320964,);
not I_18669 (I320972,I320964);
not I_18670 (I320989,I320947);
nand I_18671 (I320686,I320989,I320808);
nand I_18672 (I321020,I616243,I616219);
and I_18673 (I321037,I321020,I616240);
DFFARX1 I_18674 (I321037,I3563,I320709,I321063,);
nor I_18675 (I321071,I321063,I320735);
DFFARX1 I_18676 (I321071,I3563,I320709,I320674,);
DFFARX1 I_18677 (I321063,I3563,I320709,I320692,);
nor I_18678 (I321116,I616225,I616219);
not I_18679 (I321133,I321116);
nor I_18680 (I320695,I320972,I321133);
nand I_18681 (I320680,I320989,I321133);
nor I_18682 (I320689,I320735,I321116);
DFFARX1 I_18683 (I321116,I3563,I320709,I320698,);
not I_18684 (I321236,I3570);
DFFARX1 I_18685 (I576289,I3563,I321236,I321262,);
nand I_18686 (I321270,I576289,I576301);
and I_18687 (I321287,I321270,I576286);
DFFARX1 I_18688 (I321287,I3563,I321236,I321313,);
nor I_18689 (I321204,I321313,I321262);
not I_18690 (I321335,I321313);
DFFARX1 I_18691 (I576310,I3563,I321236,I321361,);
nand I_18692 (I321369,I321361,I576307);
not I_18693 (I321386,I321369);
DFFARX1 I_18694 (I321386,I3563,I321236,I321412,);
not I_18695 (I321228,I321412);
nor I_18696 (I321434,I321262,I321369);
nor I_18697 (I321210,I321313,I321434);
DFFARX1 I_18698 (I576298,I3563,I321236,I321474,);
DFFARX1 I_18699 (I321474,I3563,I321236,I321491,);
not I_18700 (I321499,I321491);
not I_18701 (I321516,I321474);
nand I_18702 (I321213,I321516,I321335);
nand I_18703 (I321547,I576286,I576295);
and I_18704 (I321564,I321547,I576304);
DFFARX1 I_18705 (I321564,I3563,I321236,I321590,);
nor I_18706 (I321598,I321590,I321262);
DFFARX1 I_18707 (I321598,I3563,I321236,I321201,);
DFFARX1 I_18708 (I321590,I3563,I321236,I321219,);
nor I_18709 (I321643,I576292,I576295);
not I_18710 (I321660,I321643);
nor I_18711 (I321222,I321499,I321660);
nand I_18712 (I321207,I321516,I321660);
nor I_18713 (I321216,I321262,I321643);
DFFARX1 I_18714 (I321643,I3563,I321236,I321225,);
not I_18715 (I321763,I3570);
DFFARX1 I_18716 (I1241275,I3563,I321763,I321789,);
nand I_18717 (I321797,I1241290,I1241275);
and I_18718 (I321814,I321797,I1241293);
DFFARX1 I_18719 (I321814,I3563,I321763,I321840,);
nor I_18720 (I321731,I321840,I321789);
not I_18721 (I321862,I321840);
DFFARX1 I_18722 (I1241299,I3563,I321763,I321888,);
nand I_18723 (I321896,I321888,I1241281);
not I_18724 (I321913,I321896);
DFFARX1 I_18725 (I321913,I3563,I321763,I321939,);
not I_18726 (I321755,I321939);
nor I_18727 (I321961,I321789,I321896);
nor I_18728 (I321737,I321840,I321961);
DFFARX1 I_18729 (I1241278,I3563,I321763,I322001,);
DFFARX1 I_18730 (I322001,I3563,I321763,I322018,);
not I_18731 (I322026,I322018);
not I_18732 (I322043,I322001);
nand I_18733 (I321740,I322043,I321862);
nand I_18734 (I322074,I1241278,I1241284);
and I_18735 (I322091,I322074,I1241296);
DFFARX1 I_18736 (I322091,I3563,I321763,I322117,);
nor I_18737 (I322125,I322117,I321789);
DFFARX1 I_18738 (I322125,I3563,I321763,I321728,);
DFFARX1 I_18739 (I322117,I3563,I321763,I321746,);
nor I_18740 (I322170,I1241287,I1241284);
not I_18741 (I322187,I322170);
nor I_18742 (I321749,I322026,I322187);
nand I_18743 (I321734,I322043,I322187);
nor I_18744 (I321743,I321789,I322170);
DFFARX1 I_18745 (I322170,I3563,I321763,I321752,);
not I_18746 (I322290,I3570);
DFFARX1 I_18747 (I207148,I3563,I322290,I322316,);
nand I_18748 (I322324,I207148,I207154);
and I_18749 (I322341,I322324,I207172);
DFFARX1 I_18750 (I322341,I3563,I322290,I322367,);
nor I_18751 (I322258,I322367,I322316);
not I_18752 (I322389,I322367);
DFFARX1 I_18753 (I207160,I3563,I322290,I322415,);
nand I_18754 (I322423,I322415,I207157);
not I_18755 (I322440,I322423);
DFFARX1 I_18756 (I322440,I3563,I322290,I322466,);
not I_18757 (I322282,I322466);
nor I_18758 (I322488,I322316,I322423);
nor I_18759 (I322264,I322367,I322488);
DFFARX1 I_18760 (I207166,I3563,I322290,I322528,);
DFFARX1 I_18761 (I322528,I3563,I322290,I322545,);
not I_18762 (I322553,I322545);
not I_18763 (I322570,I322528);
nand I_18764 (I322267,I322570,I322389);
nand I_18765 (I322601,I207151,I207151);
and I_18766 (I322618,I322601,I207163);
DFFARX1 I_18767 (I322618,I3563,I322290,I322644,);
nor I_18768 (I322652,I322644,I322316);
DFFARX1 I_18769 (I322652,I3563,I322290,I322255,);
DFFARX1 I_18770 (I322644,I3563,I322290,I322273,);
nor I_18771 (I322697,I207169,I207151);
not I_18772 (I322714,I322697);
nor I_18773 (I322276,I322553,I322714);
nand I_18774 (I322261,I322570,I322714);
nor I_18775 (I322270,I322316,I322697);
DFFARX1 I_18776 (I322697,I3563,I322290,I322279,);
not I_18777 (I322817,I3570);
DFFARX1 I_18778 (I1325850,I3563,I322817,I322843,);
nand I_18779 (I322851,I1325877,I1325853);
and I_18780 (I322868,I322851,I1325862);
DFFARX1 I_18781 (I322868,I3563,I322817,I322894,);
nor I_18782 (I322785,I322894,I322843);
not I_18783 (I322916,I322894);
DFFARX1 I_18784 (I1325850,I3563,I322817,I322942,);
nand I_18785 (I322950,I322942,I1325874);
not I_18786 (I322967,I322950);
DFFARX1 I_18787 (I322967,I3563,I322817,I322993,);
not I_18788 (I322809,I322993);
nor I_18789 (I323015,I322843,I322950);
nor I_18790 (I322791,I322894,I323015);
DFFARX1 I_18791 (I1325856,I3563,I322817,I323055,);
DFFARX1 I_18792 (I323055,I3563,I322817,I323072,);
not I_18793 (I323080,I323072);
not I_18794 (I323097,I323055);
nand I_18795 (I322794,I323097,I322916);
nand I_18796 (I323128,I1325871,I1325859);
and I_18797 (I323145,I323128,I1325865);
DFFARX1 I_18798 (I323145,I3563,I322817,I323171,);
nor I_18799 (I323179,I323171,I322843);
DFFARX1 I_18800 (I323179,I3563,I322817,I322782,);
DFFARX1 I_18801 (I323171,I3563,I322817,I322800,);
nor I_18802 (I323224,I1325868,I1325859);
not I_18803 (I323241,I323224);
nor I_18804 (I322803,I323080,I323241);
nand I_18805 (I322788,I323097,I323241);
nor I_18806 (I322797,I322843,I323224);
DFFARX1 I_18807 (I323224,I3563,I322817,I322806,);
not I_18808 (I323344,I3570);
DFFARX1 I_18809 (I899595,I3563,I323344,I323370,);
nand I_18810 (I323378,I899598,I899592);
and I_18811 (I323395,I323378,I899604);
DFFARX1 I_18812 (I323395,I3563,I323344,I323421,);
nor I_18813 (I323312,I323421,I323370);
not I_18814 (I323443,I323421);
DFFARX1 I_18815 (I899607,I3563,I323344,I323469,);
nand I_18816 (I323477,I323469,I899598);
not I_18817 (I323494,I323477);
DFFARX1 I_18818 (I323494,I3563,I323344,I323520,);
not I_18819 (I323336,I323520);
nor I_18820 (I323542,I323370,I323477);
nor I_18821 (I323318,I323421,I323542);
DFFARX1 I_18822 (I899610,I3563,I323344,I323582,);
DFFARX1 I_18823 (I323582,I3563,I323344,I323599,);
not I_18824 (I323607,I323599);
not I_18825 (I323624,I323582);
nand I_18826 (I323321,I323624,I323443);
nand I_18827 (I323655,I899592,I899601);
and I_18828 (I323672,I323655,I899595);
DFFARX1 I_18829 (I323672,I3563,I323344,I323698,);
nor I_18830 (I323706,I323698,I323370);
DFFARX1 I_18831 (I323706,I3563,I323344,I323309,);
DFFARX1 I_18832 (I323698,I3563,I323344,I323327,);
nor I_18833 (I323751,I899613,I899601);
not I_18834 (I323768,I323751);
nor I_18835 (I323330,I323607,I323768);
nand I_18836 (I323315,I323624,I323768);
nor I_18837 (I323324,I323370,I323751);
DFFARX1 I_18838 (I323751,I3563,I323344,I323333,);
not I_18839 (I323871,I3570);
DFFARX1 I_18840 (I124633,I3563,I323871,I323897,);
nand I_18841 (I323905,I124645,I124654);
and I_18842 (I323922,I323905,I124633);
DFFARX1 I_18843 (I323922,I3563,I323871,I323948,);
nor I_18844 (I323839,I323948,I323897);
not I_18845 (I323970,I323948);
DFFARX1 I_18846 (I124648,I3563,I323871,I323996,);
nand I_18847 (I324004,I323996,I124636);
not I_18848 (I324021,I324004);
DFFARX1 I_18849 (I324021,I3563,I323871,I324047,);
not I_18850 (I323863,I324047);
nor I_18851 (I324069,I323897,I324004);
nor I_18852 (I323845,I323948,I324069);
DFFARX1 I_18853 (I124639,I3563,I323871,I324109,);
DFFARX1 I_18854 (I324109,I3563,I323871,I324126,);
not I_18855 (I324134,I324126);
not I_18856 (I324151,I324109);
nand I_18857 (I323848,I324151,I323970);
nand I_18858 (I324182,I124630,I124630);
and I_18859 (I324199,I324182,I124642);
DFFARX1 I_18860 (I324199,I3563,I323871,I324225,);
nor I_18861 (I324233,I324225,I323897);
DFFARX1 I_18862 (I324233,I3563,I323871,I323836,);
DFFARX1 I_18863 (I324225,I3563,I323871,I323854,);
nor I_18864 (I324278,I124651,I124630);
not I_18865 (I324295,I324278);
nor I_18866 (I323857,I324134,I324295);
nand I_18867 (I323842,I324151,I324295);
nor I_18868 (I323851,I323897,I324278);
DFFARX1 I_18869 (I324278,I3563,I323871,I323860,);
not I_18870 (I324398,I3570);
DFFARX1 I_18871 (I257128,I3563,I324398,I324424,);
nand I_18872 (I324432,I257128,I257134);
and I_18873 (I324449,I324432,I257152);
DFFARX1 I_18874 (I324449,I3563,I324398,I324475,);
nor I_18875 (I324366,I324475,I324424);
not I_18876 (I324497,I324475);
DFFARX1 I_18877 (I257140,I3563,I324398,I324523,);
nand I_18878 (I324531,I324523,I257137);
not I_18879 (I324548,I324531);
DFFARX1 I_18880 (I324548,I3563,I324398,I324574,);
not I_18881 (I324390,I324574);
nor I_18882 (I324596,I324424,I324531);
nor I_18883 (I324372,I324475,I324596);
DFFARX1 I_18884 (I257146,I3563,I324398,I324636,);
DFFARX1 I_18885 (I324636,I3563,I324398,I324653,);
not I_18886 (I324661,I324653);
not I_18887 (I324678,I324636);
nand I_18888 (I324375,I324678,I324497);
nand I_18889 (I324709,I257131,I257131);
and I_18890 (I324726,I324709,I257143);
DFFARX1 I_18891 (I324726,I3563,I324398,I324752,);
nor I_18892 (I324760,I324752,I324424);
DFFARX1 I_18893 (I324760,I3563,I324398,I324363,);
DFFARX1 I_18894 (I324752,I3563,I324398,I324381,);
nor I_18895 (I324805,I257149,I257131);
not I_18896 (I324822,I324805);
nor I_18897 (I324384,I324661,I324822);
nand I_18898 (I324369,I324678,I324822);
nor I_18899 (I324378,I324424,I324805);
DFFARX1 I_18900 (I324805,I3563,I324398,I324387,);
not I_18901 (I324925,I3570);
DFFARX1 I_18902 (I1399974,I3563,I324925,I324951,);
nand I_18903 (I324959,I1399953,I1399953);
and I_18904 (I324976,I324959,I1399980);
DFFARX1 I_18905 (I324976,I3563,I324925,I325002,);
nor I_18906 (I324893,I325002,I324951);
not I_18907 (I325024,I325002);
DFFARX1 I_18908 (I1399968,I3563,I324925,I325050,);
nand I_18909 (I325058,I325050,I1399971);
not I_18910 (I325075,I325058);
DFFARX1 I_18911 (I325075,I3563,I324925,I325101,);
not I_18912 (I324917,I325101);
nor I_18913 (I325123,I324951,I325058);
nor I_18914 (I324899,I325002,I325123);
DFFARX1 I_18915 (I1399962,I3563,I324925,I325163,);
DFFARX1 I_18916 (I325163,I3563,I324925,I325180,);
not I_18917 (I325188,I325180);
not I_18918 (I325205,I325163);
nand I_18919 (I324902,I325205,I325024);
nand I_18920 (I325236,I1399959,I1399956);
and I_18921 (I325253,I325236,I1399977);
DFFARX1 I_18922 (I325253,I3563,I324925,I325279,);
nor I_18923 (I325287,I325279,I324951);
DFFARX1 I_18924 (I325287,I3563,I324925,I324890,);
DFFARX1 I_18925 (I325279,I3563,I324925,I324908,);
nor I_18926 (I325332,I1399965,I1399956);
not I_18927 (I325349,I325332);
nor I_18928 (I324911,I325188,I325349);
nand I_18929 (I324896,I325205,I325349);
nor I_18930 (I324905,I324951,I325332);
DFFARX1 I_18931 (I325332,I3563,I324925,I324914,);
not I_18932 (I325452,I3570);
DFFARX1 I_18933 (I565579,I3563,I325452,I325478,);
nand I_18934 (I325486,I565579,I565591);
and I_18935 (I325503,I325486,I565576);
DFFARX1 I_18936 (I325503,I3563,I325452,I325529,);
nor I_18937 (I325420,I325529,I325478);
not I_18938 (I325551,I325529);
DFFARX1 I_18939 (I565600,I3563,I325452,I325577,);
nand I_18940 (I325585,I325577,I565597);
not I_18941 (I325602,I325585);
DFFARX1 I_18942 (I325602,I3563,I325452,I325628,);
not I_18943 (I325444,I325628);
nor I_18944 (I325650,I325478,I325585);
nor I_18945 (I325426,I325529,I325650);
DFFARX1 I_18946 (I565588,I3563,I325452,I325690,);
DFFARX1 I_18947 (I325690,I3563,I325452,I325707,);
not I_18948 (I325715,I325707);
not I_18949 (I325732,I325690);
nand I_18950 (I325429,I325732,I325551);
nand I_18951 (I325763,I565576,I565585);
and I_18952 (I325780,I325763,I565594);
DFFARX1 I_18953 (I325780,I3563,I325452,I325806,);
nor I_18954 (I325814,I325806,I325478);
DFFARX1 I_18955 (I325814,I3563,I325452,I325417,);
DFFARX1 I_18956 (I325806,I3563,I325452,I325435,);
nor I_18957 (I325859,I565582,I565585);
not I_18958 (I325876,I325859);
nor I_18959 (I325438,I325715,I325876);
nand I_18960 (I325423,I325732,I325876);
nor I_18961 (I325432,I325478,I325859);
DFFARX1 I_18962 (I325859,I3563,I325452,I325441,);
not I_18963 (I325979,I3570);
DFFARX1 I_18964 (I1112381,I3563,I325979,I326005,);
nand I_18965 (I326013,I1112396,I1112381);
and I_18966 (I326030,I326013,I1112399);
DFFARX1 I_18967 (I326030,I3563,I325979,I326056,);
nor I_18968 (I325947,I326056,I326005);
not I_18969 (I326078,I326056);
DFFARX1 I_18970 (I1112405,I3563,I325979,I326104,);
nand I_18971 (I326112,I326104,I1112387);
not I_18972 (I326129,I326112);
DFFARX1 I_18973 (I326129,I3563,I325979,I326155,);
not I_18974 (I325971,I326155);
nor I_18975 (I326177,I326005,I326112);
nor I_18976 (I325953,I326056,I326177);
DFFARX1 I_18977 (I1112384,I3563,I325979,I326217,);
DFFARX1 I_18978 (I326217,I3563,I325979,I326234,);
not I_18979 (I326242,I326234);
not I_18980 (I326259,I326217);
nand I_18981 (I325956,I326259,I326078);
nand I_18982 (I326290,I1112384,I1112390);
and I_18983 (I326307,I326290,I1112402);
DFFARX1 I_18984 (I326307,I3563,I325979,I326333,);
nor I_18985 (I326341,I326333,I326005);
DFFARX1 I_18986 (I326341,I3563,I325979,I325944,);
DFFARX1 I_18987 (I326333,I3563,I325979,I325962,);
nor I_18988 (I326386,I1112393,I1112390);
not I_18989 (I326403,I326386);
nor I_18990 (I325965,I326242,I326403);
nand I_18991 (I325950,I326259,I326403);
nor I_18992 (I325959,I326005,I326386);
DFFARX1 I_18993 (I326386,I3563,I325979,I325968,);
not I_18994 (I326506,I3570);
DFFARX1 I_18995 (I488782,I3563,I326506,I326532,);
nand I_18996 (I326540,I488794,I488773);
and I_18997 (I326557,I326540,I488797);
DFFARX1 I_18998 (I326557,I3563,I326506,I326583,);
nor I_18999 (I326474,I326583,I326532);
not I_19000 (I326605,I326583);
DFFARX1 I_19001 (I488788,I3563,I326506,I326631,);
nand I_19002 (I326639,I326631,I488770);
not I_19003 (I326656,I326639);
DFFARX1 I_19004 (I326656,I3563,I326506,I326682,);
not I_19005 (I326498,I326682);
nor I_19006 (I326704,I326532,I326639);
nor I_19007 (I326480,I326583,I326704);
DFFARX1 I_19008 (I488785,I3563,I326506,I326744,);
DFFARX1 I_19009 (I326744,I3563,I326506,I326761,);
not I_19010 (I326769,I326761);
not I_19011 (I326786,I326744);
nand I_19012 (I326483,I326786,I326605);
nand I_19013 (I326817,I488770,I488776);
and I_19014 (I326834,I326817,I488779);
DFFARX1 I_19015 (I326834,I3563,I326506,I326860,);
nor I_19016 (I326868,I326860,I326532);
DFFARX1 I_19017 (I326868,I3563,I326506,I326471,);
DFFARX1 I_19018 (I326860,I3563,I326506,I326489,);
nor I_19019 (I326913,I488791,I488776);
not I_19020 (I326930,I326913);
nor I_19021 (I326492,I326769,I326930);
nand I_19022 (I326477,I326786,I326930);
nor I_19023 (I326486,I326532,I326913);
DFFARX1 I_19024 (I326913,I3563,I326506,I326495,);
not I_19025 (I327033,I3570);
DFFARX1 I_19026 (I1196769,I3563,I327033,I327059,);
nand I_19027 (I327067,I1196784,I1196769);
and I_19028 (I327084,I327067,I1196787);
DFFARX1 I_19029 (I327084,I3563,I327033,I327110,);
nor I_19030 (I327001,I327110,I327059);
not I_19031 (I327132,I327110);
DFFARX1 I_19032 (I1196793,I3563,I327033,I327158,);
nand I_19033 (I327166,I327158,I1196775);
not I_19034 (I327183,I327166);
DFFARX1 I_19035 (I327183,I3563,I327033,I327209,);
not I_19036 (I327025,I327209);
nor I_19037 (I327231,I327059,I327166);
nor I_19038 (I327007,I327110,I327231);
DFFARX1 I_19039 (I1196772,I3563,I327033,I327271,);
DFFARX1 I_19040 (I327271,I3563,I327033,I327288,);
not I_19041 (I327296,I327288);
not I_19042 (I327313,I327271);
nand I_19043 (I327010,I327313,I327132);
nand I_19044 (I327344,I1196772,I1196778);
and I_19045 (I327361,I327344,I1196790);
DFFARX1 I_19046 (I327361,I3563,I327033,I327387,);
nor I_19047 (I327395,I327387,I327059);
DFFARX1 I_19048 (I327395,I3563,I327033,I326998,);
DFFARX1 I_19049 (I327387,I3563,I327033,I327016,);
nor I_19050 (I327440,I1196781,I1196778);
not I_19051 (I327457,I327440);
nor I_19052 (I327019,I327296,I327457);
nand I_19053 (I327004,I327313,I327457);
nor I_19054 (I327013,I327059,I327440);
DFFARX1 I_19055 (I327440,I3563,I327033,I327022,);
not I_19056 (I327560,I3570);
DFFARX1 I_19057 (I1180585,I3563,I327560,I327586,);
nand I_19058 (I327594,I1180600,I1180585);
and I_19059 (I327611,I327594,I1180603);
DFFARX1 I_19060 (I327611,I3563,I327560,I327637,);
nor I_19061 (I327528,I327637,I327586);
not I_19062 (I327659,I327637);
DFFARX1 I_19063 (I1180609,I3563,I327560,I327685,);
nand I_19064 (I327693,I327685,I1180591);
not I_19065 (I327710,I327693);
DFFARX1 I_19066 (I327710,I3563,I327560,I327736,);
not I_19067 (I327552,I327736);
nor I_19068 (I327758,I327586,I327693);
nor I_19069 (I327534,I327637,I327758);
DFFARX1 I_19070 (I1180588,I3563,I327560,I327798,);
DFFARX1 I_19071 (I327798,I3563,I327560,I327815,);
not I_19072 (I327823,I327815);
not I_19073 (I327840,I327798);
nand I_19074 (I327537,I327840,I327659);
nand I_19075 (I327871,I1180588,I1180594);
and I_19076 (I327888,I327871,I1180606);
DFFARX1 I_19077 (I327888,I3563,I327560,I327914,);
nor I_19078 (I327922,I327914,I327586);
DFFARX1 I_19079 (I327922,I3563,I327560,I327525,);
DFFARX1 I_19080 (I327914,I3563,I327560,I327543,);
nor I_19081 (I327967,I1180597,I1180594);
not I_19082 (I327984,I327967);
nor I_19083 (I327546,I327823,I327984);
nand I_19084 (I327531,I327840,I327984);
nor I_19085 (I327540,I327586,I327967);
DFFARX1 I_19086 (I327967,I3563,I327560,I327549,);
not I_19087 (I328087,I3570);
DFFARX1 I_19088 (I1170181,I3563,I328087,I328113,);
nand I_19089 (I328121,I1170196,I1170181);
and I_19090 (I328138,I328121,I1170199);
DFFARX1 I_19091 (I328138,I3563,I328087,I328164,);
nor I_19092 (I328055,I328164,I328113);
not I_19093 (I328186,I328164);
DFFARX1 I_19094 (I1170205,I3563,I328087,I328212,);
nand I_19095 (I328220,I328212,I1170187);
not I_19096 (I328237,I328220);
DFFARX1 I_19097 (I328237,I3563,I328087,I328263,);
not I_19098 (I328079,I328263);
nor I_19099 (I328285,I328113,I328220);
nor I_19100 (I328061,I328164,I328285);
DFFARX1 I_19101 (I1170184,I3563,I328087,I328325,);
DFFARX1 I_19102 (I328325,I3563,I328087,I328342,);
not I_19103 (I328350,I328342);
not I_19104 (I328367,I328325);
nand I_19105 (I328064,I328367,I328186);
nand I_19106 (I328398,I1170184,I1170190);
and I_19107 (I328415,I328398,I1170202);
DFFARX1 I_19108 (I328415,I3563,I328087,I328441,);
nor I_19109 (I328449,I328441,I328113);
DFFARX1 I_19110 (I328449,I3563,I328087,I328052,);
DFFARX1 I_19111 (I328441,I3563,I328087,I328070,);
nor I_19112 (I328494,I1170193,I1170190);
not I_19113 (I328511,I328494);
nor I_19114 (I328073,I328350,I328511);
nand I_19115 (I328058,I328367,I328511);
nor I_19116 (I328067,I328113,I328494);
DFFARX1 I_19117 (I328494,I3563,I328087,I328076,);
not I_19118 (I328614,I3570);
DFFARX1 I_19119 (I473550,I3563,I328614,I328640,);
nand I_19120 (I328648,I473562,I473541);
and I_19121 (I328665,I328648,I473565);
DFFARX1 I_19122 (I328665,I3563,I328614,I328691,);
nor I_19123 (I328582,I328691,I328640);
not I_19124 (I328713,I328691);
DFFARX1 I_19125 (I473556,I3563,I328614,I328739,);
nand I_19126 (I328747,I328739,I473538);
not I_19127 (I328764,I328747);
DFFARX1 I_19128 (I328764,I3563,I328614,I328790,);
not I_19129 (I328606,I328790);
nor I_19130 (I328812,I328640,I328747);
nor I_19131 (I328588,I328691,I328812);
DFFARX1 I_19132 (I473553,I3563,I328614,I328852,);
DFFARX1 I_19133 (I328852,I3563,I328614,I328869,);
not I_19134 (I328877,I328869);
not I_19135 (I328894,I328852);
nand I_19136 (I328591,I328894,I328713);
nand I_19137 (I328925,I473538,I473544);
and I_19138 (I328942,I328925,I473547);
DFFARX1 I_19139 (I328942,I3563,I328614,I328968,);
nor I_19140 (I328976,I328968,I328640);
DFFARX1 I_19141 (I328976,I3563,I328614,I328579,);
DFFARX1 I_19142 (I328968,I3563,I328614,I328597,);
nor I_19143 (I329021,I473559,I473544);
not I_19144 (I329038,I329021);
nor I_19145 (I328600,I328877,I329038);
nand I_19146 (I328585,I328894,I329038);
nor I_19147 (I328594,I328640,I329021);
DFFARX1 I_19148 (I329021,I3563,I328614,I328603,);
not I_19149 (I329141,I3570);
DFFARX1 I_19150 (I660737,I3563,I329141,I329167,);
nand I_19151 (I329175,I660728,I660743);
and I_19152 (I329192,I329175,I660749);
DFFARX1 I_19153 (I329192,I3563,I329141,I329218,);
nor I_19154 (I329109,I329218,I329167);
not I_19155 (I329240,I329218);
DFFARX1 I_19156 (I660734,I3563,I329141,I329266,);
nand I_19157 (I329274,I329266,I660728);
not I_19158 (I329291,I329274);
DFFARX1 I_19159 (I329291,I3563,I329141,I329317,);
not I_19160 (I329133,I329317);
nor I_19161 (I329339,I329167,I329274);
nor I_19162 (I329115,I329218,I329339);
DFFARX1 I_19163 (I660731,I3563,I329141,I329379,);
DFFARX1 I_19164 (I329379,I3563,I329141,I329396,);
not I_19165 (I329404,I329396);
not I_19166 (I329421,I329379);
nand I_19167 (I329118,I329421,I329240);
nand I_19168 (I329452,I660725,I660740);
and I_19169 (I329469,I329452,I660725);
DFFARX1 I_19170 (I329469,I3563,I329141,I329495,);
nor I_19171 (I329503,I329495,I329167);
DFFARX1 I_19172 (I329503,I3563,I329141,I329106,);
DFFARX1 I_19173 (I329495,I3563,I329141,I329124,);
nor I_19174 (I329548,I660746,I660740);
not I_19175 (I329565,I329548);
nor I_19176 (I329127,I329404,I329565);
nand I_19177 (I329112,I329421,I329565);
nor I_19178 (I329121,I329167,I329548);
DFFARX1 I_19179 (I329548,I3563,I329141,I329130,);
not I_19180 (I329668,I3570);
DFFARX1 I_19181 (I173828,I3563,I329668,I329694,);
nand I_19182 (I329702,I173828,I173834);
and I_19183 (I329719,I329702,I173852);
DFFARX1 I_19184 (I329719,I3563,I329668,I329745,);
nor I_19185 (I329636,I329745,I329694);
not I_19186 (I329767,I329745);
DFFARX1 I_19187 (I173840,I3563,I329668,I329793,);
nand I_19188 (I329801,I329793,I173837);
not I_19189 (I329818,I329801);
DFFARX1 I_19190 (I329818,I3563,I329668,I329844,);
not I_19191 (I329660,I329844);
nor I_19192 (I329866,I329694,I329801);
nor I_19193 (I329642,I329745,I329866);
DFFARX1 I_19194 (I173846,I3563,I329668,I329906,);
DFFARX1 I_19195 (I329906,I3563,I329668,I329923,);
not I_19196 (I329931,I329923);
not I_19197 (I329948,I329906);
nand I_19198 (I329645,I329948,I329767);
nand I_19199 (I329979,I173831,I173831);
and I_19200 (I329996,I329979,I173843);
DFFARX1 I_19201 (I329996,I3563,I329668,I330022,);
nor I_19202 (I330030,I330022,I329694);
DFFARX1 I_19203 (I330030,I3563,I329668,I329633,);
DFFARX1 I_19204 (I330022,I3563,I329668,I329651,);
nor I_19205 (I330075,I173849,I173831);
not I_19206 (I330092,I330075);
nor I_19207 (I329654,I329931,I330092);
nand I_19208 (I329639,I329948,I330092);
nor I_19209 (I329648,I329694,I330075);
DFFARX1 I_19210 (I330075,I3563,I329668,I329657,);
not I_19211 (I330195,I3570);
DFFARX1 I_19212 (I1150529,I3563,I330195,I330221,);
nand I_19213 (I330229,I1150544,I1150529);
and I_19214 (I330246,I330229,I1150547);
DFFARX1 I_19215 (I330246,I3563,I330195,I330272,);
nor I_19216 (I330163,I330272,I330221);
not I_19217 (I330294,I330272);
DFFARX1 I_19218 (I1150553,I3563,I330195,I330320,);
nand I_19219 (I330328,I330320,I1150535);
not I_19220 (I330345,I330328);
DFFARX1 I_19221 (I330345,I3563,I330195,I330371,);
not I_19222 (I330187,I330371);
nor I_19223 (I330393,I330221,I330328);
nor I_19224 (I330169,I330272,I330393);
DFFARX1 I_19225 (I1150532,I3563,I330195,I330433,);
DFFARX1 I_19226 (I330433,I3563,I330195,I330450,);
not I_19227 (I330458,I330450);
not I_19228 (I330475,I330433);
nand I_19229 (I330172,I330475,I330294);
nand I_19230 (I330506,I1150532,I1150538);
and I_19231 (I330523,I330506,I1150550);
DFFARX1 I_19232 (I330523,I3563,I330195,I330549,);
nor I_19233 (I330557,I330549,I330221);
DFFARX1 I_19234 (I330557,I3563,I330195,I330160,);
DFFARX1 I_19235 (I330549,I3563,I330195,I330178,);
nor I_19236 (I330602,I1150541,I1150538);
not I_19237 (I330619,I330602);
nor I_19238 (I330181,I330458,I330619);
nand I_19239 (I330166,I330475,I330619);
nor I_19240 (I330175,I330221,I330602);
DFFARX1 I_19241 (I330602,I3563,I330195,I330184,);
not I_19242 (I330722,I3570);
DFFARX1 I_19243 (I170258,I3563,I330722,I330748,);
nand I_19244 (I330756,I170258,I170264);
and I_19245 (I330773,I330756,I170282);
DFFARX1 I_19246 (I330773,I3563,I330722,I330799,);
nor I_19247 (I330690,I330799,I330748);
not I_19248 (I330821,I330799);
DFFARX1 I_19249 (I170270,I3563,I330722,I330847,);
nand I_19250 (I330855,I330847,I170267);
not I_19251 (I330872,I330855);
DFFARX1 I_19252 (I330872,I3563,I330722,I330898,);
not I_19253 (I330714,I330898);
nor I_19254 (I330920,I330748,I330855);
nor I_19255 (I330696,I330799,I330920);
DFFARX1 I_19256 (I170276,I3563,I330722,I330960,);
DFFARX1 I_19257 (I330960,I3563,I330722,I330977,);
not I_19258 (I330985,I330977);
not I_19259 (I331002,I330960);
nand I_19260 (I330699,I331002,I330821);
nand I_19261 (I331033,I170261,I170261);
and I_19262 (I331050,I331033,I170273);
DFFARX1 I_19263 (I331050,I3563,I330722,I331076,);
nor I_19264 (I331084,I331076,I330748);
DFFARX1 I_19265 (I331084,I3563,I330722,I330687,);
DFFARX1 I_19266 (I331076,I3563,I330722,I330705,);
nor I_19267 (I331129,I170279,I170261);
not I_19268 (I331146,I331129);
nor I_19269 (I330708,I330985,I331146);
nand I_19270 (I330693,I331002,I331146);
nor I_19271 (I330702,I330748,I331129);
DFFARX1 I_19272 (I331129,I3563,I330722,I330711,);
not I_19273 (I331249,I3570);
DFFARX1 I_19274 (I844260,I3563,I331249,I331275,);
nand I_19275 (I331283,I844263,I844257);
and I_19276 (I331300,I331283,I844269);
DFFARX1 I_19277 (I331300,I3563,I331249,I331326,);
nor I_19278 (I331217,I331326,I331275);
not I_19279 (I331348,I331326);
DFFARX1 I_19280 (I844272,I3563,I331249,I331374,);
nand I_19281 (I331382,I331374,I844263);
not I_19282 (I331399,I331382);
DFFARX1 I_19283 (I331399,I3563,I331249,I331425,);
not I_19284 (I331241,I331425);
nor I_19285 (I331447,I331275,I331382);
nor I_19286 (I331223,I331326,I331447);
DFFARX1 I_19287 (I844275,I3563,I331249,I331487,);
DFFARX1 I_19288 (I331487,I3563,I331249,I331504,);
not I_19289 (I331512,I331504);
not I_19290 (I331529,I331487);
nand I_19291 (I331226,I331529,I331348);
nand I_19292 (I331560,I844257,I844266);
and I_19293 (I331577,I331560,I844260);
DFFARX1 I_19294 (I331577,I3563,I331249,I331603,);
nor I_19295 (I331611,I331603,I331275);
DFFARX1 I_19296 (I331611,I3563,I331249,I331214,);
DFFARX1 I_19297 (I331603,I3563,I331249,I331232,);
nor I_19298 (I331656,I844278,I844266);
not I_19299 (I331673,I331656);
nor I_19300 (I331235,I331512,I331673);
nand I_19301 (I331220,I331529,I331673);
nor I_19302 (I331229,I331275,I331656);
DFFARX1 I_19303 (I331656,I3563,I331249,I331238,);
not I_19304 (I331776,I3570);
DFFARX1 I_19305 (I851638,I3563,I331776,I331802,);
nand I_19306 (I331810,I851641,I851635);
and I_19307 (I331827,I331810,I851647);
DFFARX1 I_19308 (I331827,I3563,I331776,I331853,);
nor I_19309 (I331744,I331853,I331802);
not I_19310 (I331875,I331853);
DFFARX1 I_19311 (I851650,I3563,I331776,I331901,);
nand I_19312 (I331909,I331901,I851641);
not I_19313 (I331926,I331909);
DFFARX1 I_19314 (I331926,I3563,I331776,I331952,);
not I_19315 (I331768,I331952);
nor I_19316 (I331974,I331802,I331909);
nor I_19317 (I331750,I331853,I331974);
DFFARX1 I_19318 (I851653,I3563,I331776,I332014,);
DFFARX1 I_19319 (I332014,I3563,I331776,I332031,);
not I_19320 (I332039,I332031);
not I_19321 (I332056,I332014);
nand I_19322 (I331753,I332056,I331875);
nand I_19323 (I332087,I851635,I851644);
and I_19324 (I332104,I332087,I851638);
DFFARX1 I_19325 (I332104,I3563,I331776,I332130,);
nor I_19326 (I332138,I332130,I331802);
DFFARX1 I_19327 (I332138,I3563,I331776,I331741,);
DFFARX1 I_19328 (I332130,I3563,I331776,I331759,);
nor I_19329 (I332183,I851656,I851644);
not I_19330 (I332200,I332183);
nor I_19331 (I331762,I332039,I332200);
nand I_19332 (I331747,I332056,I332200);
nor I_19333 (I331756,I331802,I332183);
DFFARX1 I_19334 (I332183,I3563,I331776,I331765,);
not I_19335 (I332303,I3570);
DFFARX1 I_19336 (I267243,I3563,I332303,I332329,);
nand I_19337 (I332337,I267243,I267249);
and I_19338 (I332354,I332337,I267267);
DFFARX1 I_19339 (I332354,I3563,I332303,I332380,);
nor I_19340 (I332271,I332380,I332329);
not I_19341 (I332402,I332380);
DFFARX1 I_19342 (I267255,I3563,I332303,I332428,);
nand I_19343 (I332436,I332428,I267252);
not I_19344 (I332453,I332436);
DFFARX1 I_19345 (I332453,I3563,I332303,I332479,);
not I_19346 (I332295,I332479);
nor I_19347 (I332501,I332329,I332436);
nor I_19348 (I332277,I332380,I332501);
DFFARX1 I_19349 (I267261,I3563,I332303,I332541,);
DFFARX1 I_19350 (I332541,I3563,I332303,I332558,);
not I_19351 (I332566,I332558);
not I_19352 (I332583,I332541);
nand I_19353 (I332280,I332583,I332402);
nand I_19354 (I332614,I267246,I267246);
and I_19355 (I332631,I332614,I267258);
DFFARX1 I_19356 (I332631,I3563,I332303,I332657,);
nor I_19357 (I332665,I332657,I332329);
DFFARX1 I_19358 (I332665,I3563,I332303,I332268,);
DFFARX1 I_19359 (I332657,I3563,I332303,I332286,);
nor I_19360 (I332710,I267264,I267246);
not I_19361 (I332727,I332710);
nor I_19362 (I332289,I332566,I332727);
nand I_19363 (I332274,I332583,I332727);
nor I_19364 (I332283,I332329,I332710);
DFFARX1 I_19365 (I332710,I3563,I332303,I332292,);
not I_19366 (I332830,I3570);
DFFARX1 I_19367 (I909081,I3563,I332830,I332856,);
nand I_19368 (I332864,I909084,I909078);
and I_19369 (I332881,I332864,I909090);
DFFARX1 I_19370 (I332881,I3563,I332830,I332907,);
nor I_19371 (I332798,I332907,I332856);
not I_19372 (I332929,I332907);
DFFARX1 I_19373 (I909093,I3563,I332830,I332955,);
nand I_19374 (I332963,I332955,I909084);
not I_19375 (I332980,I332963);
DFFARX1 I_19376 (I332980,I3563,I332830,I333006,);
not I_19377 (I332822,I333006);
nor I_19378 (I333028,I332856,I332963);
nor I_19379 (I332804,I332907,I333028);
DFFARX1 I_19380 (I909096,I3563,I332830,I333068,);
DFFARX1 I_19381 (I333068,I3563,I332830,I333085,);
not I_19382 (I333093,I333085);
not I_19383 (I333110,I333068);
nand I_19384 (I332807,I333110,I332929);
nand I_19385 (I333141,I909078,I909087);
and I_19386 (I333158,I333141,I909081);
DFFARX1 I_19387 (I333158,I3563,I332830,I333184,);
nor I_19388 (I333192,I333184,I332856);
DFFARX1 I_19389 (I333192,I3563,I332830,I332795,);
DFFARX1 I_19390 (I333184,I3563,I332830,I332813,);
nor I_19391 (I333237,I909099,I909087);
not I_19392 (I333254,I333237);
nor I_19393 (I332816,I333093,I333254);
nand I_19394 (I332801,I333110,I333254);
nor I_19395 (I332810,I332856,I333237);
DFFARX1 I_19396 (I333237,I3563,I332830,I332819,);
not I_19397 (I333357,I3570);
DFFARX1 I_19398 (I1040202,I3563,I333357,I333383,);
nand I_19399 (I333391,I1040199,I1040217);
and I_19400 (I333408,I333391,I1040208);
DFFARX1 I_19401 (I333408,I3563,I333357,I333434,);
nor I_19402 (I333325,I333434,I333383);
not I_19403 (I333456,I333434);
DFFARX1 I_19404 (I1040223,I3563,I333357,I333482,);
nand I_19405 (I333490,I333482,I1040205);
not I_19406 (I333507,I333490);
DFFARX1 I_19407 (I333507,I3563,I333357,I333533,);
not I_19408 (I333349,I333533);
nor I_19409 (I333555,I333383,I333490);
nor I_19410 (I333331,I333434,I333555);
DFFARX1 I_19411 (I1040211,I3563,I333357,I333595,);
DFFARX1 I_19412 (I333595,I3563,I333357,I333612,);
not I_19413 (I333620,I333612);
not I_19414 (I333637,I333595);
nand I_19415 (I333334,I333637,I333456);
nand I_19416 (I333668,I1040199,I1040226);
and I_19417 (I333685,I333668,I1040214);
DFFARX1 I_19418 (I333685,I3563,I333357,I333711,);
nor I_19419 (I333719,I333711,I333383);
DFFARX1 I_19420 (I333719,I3563,I333357,I333322,);
DFFARX1 I_19421 (I333711,I3563,I333357,I333340,);
nor I_19422 (I333764,I1040220,I1040226);
not I_19423 (I333781,I333764);
nor I_19424 (I333343,I333620,I333781);
nand I_19425 (I333328,I333637,I333781);
nor I_19426 (I333337,I333383,I333764);
DFFARX1 I_19427 (I333764,I3563,I333357,I333346,);
not I_19428 (I333884,I3570);
DFFARX1 I_19429 (I2484,I3563,I333884,I333910,);
nand I_19430 (I333918,I2236,I3100);
and I_19431 (I333935,I333918,I2316);
DFFARX1 I_19432 (I333935,I3563,I333884,I333961,);
nor I_19433 (I333852,I333961,I333910);
not I_19434 (I333983,I333961);
DFFARX1 I_19435 (I2796,I3563,I333884,I334009,);
nand I_19436 (I334017,I334009,I3164);
not I_19437 (I334034,I334017);
DFFARX1 I_19438 (I334034,I3563,I333884,I334060,);
not I_19439 (I333876,I334060);
nor I_19440 (I334082,I333910,I334017);
nor I_19441 (I333858,I333961,I334082);
DFFARX1 I_19442 (I3348,I3563,I333884,I334122,);
DFFARX1 I_19443 (I334122,I3563,I333884,I334139,);
not I_19444 (I334147,I334139);
not I_19445 (I334164,I334122);
nand I_19446 (I333861,I334164,I333983);
nand I_19447 (I334195,I2844,I2212);
and I_19448 (I334212,I334195,I2780);
DFFARX1 I_19449 (I334212,I3563,I333884,I334238,);
nor I_19450 (I334246,I334238,I333910);
DFFARX1 I_19451 (I334246,I3563,I333884,I333849,);
DFFARX1 I_19452 (I334238,I3563,I333884,I333867,);
nor I_19453 (I334291,I2980,I2212);
not I_19454 (I334308,I334291);
nor I_19455 (I333870,I334147,I334308);
nand I_19456 (I333855,I334164,I334308);
nor I_19457 (I333864,I333910,I334291);
DFFARX1 I_19458 (I334291,I3563,I333884,I333873,);
not I_19459 (I334411,I3570);
DFFARX1 I_19460 (I450158,I3563,I334411,I334437,);
nand I_19461 (I334445,I450170,I450149);
and I_19462 (I334462,I334445,I450173);
DFFARX1 I_19463 (I334462,I3563,I334411,I334488,);
nor I_19464 (I334379,I334488,I334437);
not I_19465 (I334510,I334488);
DFFARX1 I_19466 (I450164,I3563,I334411,I334536,);
nand I_19467 (I334544,I334536,I450146);
not I_19468 (I334561,I334544);
DFFARX1 I_19469 (I334561,I3563,I334411,I334587,);
not I_19470 (I334403,I334587);
nor I_19471 (I334609,I334437,I334544);
nor I_19472 (I334385,I334488,I334609);
DFFARX1 I_19473 (I450161,I3563,I334411,I334649,);
DFFARX1 I_19474 (I334649,I3563,I334411,I334666,);
not I_19475 (I334674,I334666);
not I_19476 (I334691,I334649);
nand I_19477 (I334388,I334691,I334510);
nand I_19478 (I334722,I450146,I450152);
and I_19479 (I334739,I334722,I450155);
DFFARX1 I_19480 (I334739,I3563,I334411,I334765,);
nor I_19481 (I334773,I334765,I334437);
DFFARX1 I_19482 (I334773,I3563,I334411,I334376,);
DFFARX1 I_19483 (I334765,I3563,I334411,I334394,);
nor I_19484 (I334818,I450167,I450152);
not I_19485 (I334835,I334818);
nor I_19486 (I334397,I334674,I334835);
nand I_19487 (I334382,I334691,I334835);
nor I_19488 (I334391,I334437,I334818);
DFFARX1 I_19489 (I334818,I3563,I334411,I334400,);
not I_19490 (I334938,I3570);
DFFARX1 I_19491 (I1402949,I3563,I334938,I334964,);
nand I_19492 (I334972,I1402928,I1402928);
and I_19493 (I334989,I334972,I1402955);
DFFARX1 I_19494 (I334989,I3563,I334938,I335015,);
nor I_19495 (I334906,I335015,I334964);
not I_19496 (I335037,I335015);
DFFARX1 I_19497 (I1402943,I3563,I334938,I335063,);
nand I_19498 (I335071,I335063,I1402946);
not I_19499 (I335088,I335071);
DFFARX1 I_19500 (I335088,I3563,I334938,I335114,);
not I_19501 (I334930,I335114);
nor I_19502 (I335136,I334964,I335071);
nor I_19503 (I334912,I335015,I335136);
DFFARX1 I_19504 (I1402937,I3563,I334938,I335176,);
DFFARX1 I_19505 (I335176,I3563,I334938,I335193,);
not I_19506 (I335201,I335193);
not I_19507 (I335218,I335176);
nand I_19508 (I334915,I335218,I335037);
nand I_19509 (I335249,I1402934,I1402931);
and I_19510 (I335266,I335249,I1402952);
DFFARX1 I_19511 (I335266,I3563,I334938,I335292,);
nor I_19512 (I335300,I335292,I334964);
DFFARX1 I_19513 (I335300,I3563,I334938,I334903,);
DFFARX1 I_19514 (I335292,I3563,I334938,I334921,);
nor I_19515 (I335345,I1402940,I1402931);
not I_19516 (I335362,I335345);
nor I_19517 (I334924,I335201,I335362);
nand I_19518 (I334909,I335218,I335362);
nor I_19519 (I334918,I334964,I335345);
DFFARX1 I_19520 (I335345,I3563,I334938,I334927,);
not I_19521 (I335465,I3570);
DFFARX1 I_19522 (I1371414,I3563,I335465,I335491,);
nand I_19523 (I335499,I1371393,I1371393);
and I_19524 (I335516,I335499,I1371420);
DFFARX1 I_19525 (I335516,I3563,I335465,I335542,);
nor I_19526 (I335433,I335542,I335491);
not I_19527 (I335564,I335542);
DFFARX1 I_19528 (I1371408,I3563,I335465,I335590,);
nand I_19529 (I335598,I335590,I1371411);
not I_19530 (I335615,I335598);
DFFARX1 I_19531 (I335615,I3563,I335465,I335641,);
not I_19532 (I335457,I335641);
nor I_19533 (I335663,I335491,I335598);
nor I_19534 (I335439,I335542,I335663);
DFFARX1 I_19535 (I1371402,I3563,I335465,I335703,);
DFFARX1 I_19536 (I335703,I3563,I335465,I335720,);
not I_19537 (I335728,I335720);
not I_19538 (I335745,I335703);
nand I_19539 (I335442,I335745,I335564);
nand I_19540 (I335776,I1371399,I1371396);
and I_19541 (I335793,I335776,I1371417);
DFFARX1 I_19542 (I335793,I3563,I335465,I335819,);
nor I_19543 (I335827,I335819,I335491);
DFFARX1 I_19544 (I335827,I3563,I335465,I335430,);
DFFARX1 I_19545 (I335819,I3563,I335465,I335448,);
nor I_19546 (I335872,I1371405,I1371396);
not I_19547 (I335889,I335872);
nor I_19548 (I335451,I335728,I335889);
nand I_19549 (I335436,I335745,I335889);
nor I_19550 (I335445,I335491,I335872);
DFFARX1 I_19551 (I335872,I3563,I335465,I335454,);
not I_19552 (I335992,I3570);
DFFARX1 I_19553 (I193463,I3563,I335992,I336018,);
nand I_19554 (I336026,I193463,I193469);
and I_19555 (I336043,I336026,I193487);
DFFARX1 I_19556 (I336043,I3563,I335992,I336069,);
nor I_19557 (I335960,I336069,I336018);
not I_19558 (I336091,I336069);
DFFARX1 I_19559 (I193475,I3563,I335992,I336117,);
nand I_19560 (I336125,I336117,I193472);
not I_19561 (I336142,I336125);
DFFARX1 I_19562 (I336142,I3563,I335992,I336168,);
not I_19563 (I335984,I336168);
nor I_19564 (I336190,I336018,I336125);
nor I_19565 (I335966,I336069,I336190);
DFFARX1 I_19566 (I193481,I3563,I335992,I336230,);
DFFARX1 I_19567 (I336230,I3563,I335992,I336247,);
not I_19568 (I336255,I336247);
not I_19569 (I336272,I336230);
nand I_19570 (I335969,I336272,I336091);
nand I_19571 (I336303,I193466,I193466);
and I_19572 (I336320,I336303,I193478);
DFFARX1 I_19573 (I336320,I3563,I335992,I336346,);
nor I_19574 (I336354,I336346,I336018);
DFFARX1 I_19575 (I336354,I3563,I335992,I335957,);
DFFARX1 I_19576 (I336346,I3563,I335992,I335975,);
nor I_19577 (I336399,I193484,I193466);
not I_19578 (I336416,I336399);
nor I_19579 (I335978,I336255,I336416);
nand I_19580 (I335963,I336272,I336416);
nor I_19581 (I335972,I336018,I336399);
DFFARX1 I_19582 (I336399,I3563,I335992,I335981,);
not I_19583 (I336519,I3570);
DFFARX1 I_19584 (I1071346,I3563,I336519,I336545,);
nand I_19585 (I336553,I1071343,I1071346);
and I_19586 (I336570,I336553,I1071355);
DFFARX1 I_19587 (I336570,I3563,I336519,I336596,);
nor I_19588 (I336487,I336596,I336545);
not I_19589 (I336618,I336596);
DFFARX1 I_19590 (I1071343,I3563,I336519,I336644,);
nand I_19591 (I336652,I336644,I1071361);
not I_19592 (I336669,I336652);
DFFARX1 I_19593 (I336669,I3563,I336519,I336695,);
not I_19594 (I336511,I336695);
nor I_19595 (I336717,I336545,I336652);
nor I_19596 (I336493,I336596,I336717);
DFFARX1 I_19597 (I1071349,I3563,I336519,I336757,);
DFFARX1 I_19598 (I336757,I3563,I336519,I336774,);
not I_19599 (I336782,I336774);
not I_19600 (I336799,I336757);
nand I_19601 (I336496,I336799,I336618);
nand I_19602 (I336830,I1071358,I1071364);
and I_19603 (I336847,I336830,I1071349);
DFFARX1 I_19604 (I336847,I3563,I336519,I336873,);
nor I_19605 (I336881,I336873,I336545);
DFFARX1 I_19606 (I336881,I3563,I336519,I336484,);
DFFARX1 I_19607 (I336873,I3563,I336519,I336502,);
nor I_19608 (I336926,I1071352,I1071364);
not I_19609 (I336943,I336926);
nor I_19610 (I336505,I336782,I336943);
nand I_19611 (I336490,I336799,I336943);
nor I_19612 (I336499,I336545,I336926);
DFFARX1 I_19613 (I336926,I3563,I336519,I336508,);
not I_19614 (I337046,I3570);
DFFARX1 I_19615 (I806971,I3563,I337046,I337072,);
nand I_19616 (I337080,I806962,I806977);
and I_19617 (I337097,I337080,I806983);
DFFARX1 I_19618 (I337097,I3563,I337046,I337123,);
nor I_19619 (I337014,I337123,I337072);
not I_19620 (I337145,I337123);
DFFARX1 I_19621 (I806968,I3563,I337046,I337171,);
nand I_19622 (I337179,I337171,I806962);
not I_19623 (I337196,I337179);
DFFARX1 I_19624 (I337196,I3563,I337046,I337222,);
not I_19625 (I337038,I337222);
nor I_19626 (I337244,I337072,I337179);
nor I_19627 (I337020,I337123,I337244);
DFFARX1 I_19628 (I806965,I3563,I337046,I337284,);
DFFARX1 I_19629 (I337284,I3563,I337046,I337301,);
not I_19630 (I337309,I337301);
not I_19631 (I337326,I337284);
nand I_19632 (I337023,I337326,I337145);
nand I_19633 (I337357,I806959,I806974);
and I_19634 (I337374,I337357,I806959);
DFFARX1 I_19635 (I337374,I3563,I337046,I337400,);
nor I_19636 (I337408,I337400,I337072);
DFFARX1 I_19637 (I337408,I3563,I337046,I337011,);
DFFARX1 I_19638 (I337400,I3563,I337046,I337029,);
nor I_19639 (I337453,I806980,I806974);
not I_19640 (I337470,I337453);
nor I_19641 (I337032,I337309,I337470);
nand I_19642 (I337017,I337326,I337470);
nor I_19643 (I337026,I337072,I337453);
DFFARX1 I_19644 (I337453,I3563,I337046,I337035,);
not I_19645 (I337573,I3570);
DFFARX1 I_19646 (I1022760,I3563,I337573,I337599,);
nand I_19647 (I337607,I1022757,I1022775);
and I_19648 (I337624,I337607,I1022766);
DFFARX1 I_19649 (I337624,I3563,I337573,I337650,);
nor I_19650 (I337541,I337650,I337599);
not I_19651 (I337672,I337650);
DFFARX1 I_19652 (I1022781,I3563,I337573,I337698,);
nand I_19653 (I337706,I337698,I1022763);
not I_19654 (I337723,I337706);
DFFARX1 I_19655 (I337723,I3563,I337573,I337749,);
not I_19656 (I337565,I337749);
nor I_19657 (I337771,I337599,I337706);
nor I_19658 (I337547,I337650,I337771);
DFFARX1 I_19659 (I1022769,I3563,I337573,I337811,);
DFFARX1 I_19660 (I337811,I3563,I337573,I337828,);
not I_19661 (I337836,I337828);
not I_19662 (I337853,I337811);
nand I_19663 (I337550,I337853,I337672);
nand I_19664 (I337884,I1022757,I1022784);
and I_19665 (I337901,I337884,I1022772);
DFFARX1 I_19666 (I337901,I3563,I337573,I337927,);
nor I_19667 (I337935,I337927,I337599);
DFFARX1 I_19668 (I337935,I3563,I337573,I337538,);
DFFARX1 I_19669 (I337927,I3563,I337573,I337556,);
nor I_19670 (I337980,I1022778,I1022784);
not I_19671 (I337997,I337980);
nor I_19672 (I337559,I337836,I337997);
nand I_19673 (I337544,I337853,I337997);
nor I_19674 (I337553,I337599,I337980);
DFFARX1 I_19675 (I337980,I3563,I337573,I337562,);
not I_19676 (I338100,I3570);
DFFARX1 I_19677 (I624326,I3563,I338100,I338126,);
nand I_19678 (I338134,I624311,I624314);
and I_19679 (I338151,I338134,I624329);
DFFARX1 I_19680 (I338151,I3563,I338100,I338177,);
nor I_19681 (I338068,I338177,I338126);
not I_19682 (I338199,I338177);
DFFARX1 I_19683 (I624323,I3563,I338100,I338225,);
nand I_19684 (I338233,I338225,I624314);
not I_19685 (I338250,I338233);
DFFARX1 I_19686 (I338250,I3563,I338100,I338276,);
not I_19687 (I338092,I338276);
nor I_19688 (I338298,I338126,I338233);
nor I_19689 (I338074,I338177,I338298);
DFFARX1 I_19690 (I624320,I3563,I338100,I338338,);
DFFARX1 I_19691 (I338338,I3563,I338100,I338355,);
not I_19692 (I338363,I338355);
not I_19693 (I338380,I338338);
nand I_19694 (I338077,I338380,I338199);
nand I_19695 (I338411,I624335,I624311);
and I_19696 (I338428,I338411,I624332);
DFFARX1 I_19697 (I338428,I3563,I338100,I338454,);
nor I_19698 (I338462,I338454,I338126);
DFFARX1 I_19699 (I338462,I3563,I338100,I338065,);
DFFARX1 I_19700 (I338454,I3563,I338100,I338083,);
nor I_19701 (I338507,I624317,I624311);
not I_19702 (I338524,I338507);
nor I_19703 (I338086,I338363,I338524);
nand I_19704 (I338071,I338380,I338524);
nor I_19705 (I338080,I338126,I338507);
DFFARX1 I_19706 (I338507,I3563,I338100,I338089,);
not I_19707 (I338627,I3570);
DFFARX1 I_19708 (I100391,I3563,I338627,I338653,);
nand I_19709 (I338661,I100403,I100412);
and I_19710 (I338678,I338661,I100391);
DFFARX1 I_19711 (I338678,I3563,I338627,I338704,);
nor I_19712 (I338595,I338704,I338653);
not I_19713 (I338726,I338704);
DFFARX1 I_19714 (I100406,I3563,I338627,I338752,);
nand I_19715 (I338760,I338752,I100394);
not I_19716 (I338777,I338760);
DFFARX1 I_19717 (I338777,I3563,I338627,I338803,);
not I_19718 (I338619,I338803);
nor I_19719 (I338825,I338653,I338760);
nor I_19720 (I338601,I338704,I338825);
DFFARX1 I_19721 (I100397,I3563,I338627,I338865,);
DFFARX1 I_19722 (I338865,I3563,I338627,I338882,);
not I_19723 (I338890,I338882);
not I_19724 (I338907,I338865);
nand I_19725 (I338604,I338907,I338726);
nand I_19726 (I338938,I100388,I100388);
and I_19727 (I338955,I338938,I100400);
DFFARX1 I_19728 (I338955,I3563,I338627,I338981,);
nor I_19729 (I338989,I338981,I338653);
DFFARX1 I_19730 (I338989,I3563,I338627,I338592,);
DFFARX1 I_19731 (I338981,I3563,I338627,I338610,);
nor I_19732 (I339034,I100409,I100388);
not I_19733 (I339051,I339034);
nor I_19734 (I338613,I338890,I339051);
nand I_19735 (I338598,I338907,I339051);
nor I_19736 (I338607,I338653,I339034);
DFFARX1 I_19737 (I339034,I3563,I338627,I338616,);
not I_19738 (I339154,I3570);
DFFARX1 I_19739 (I768245,I3563,I339154,I339180,);
nand I_19740 (I339188,I768236,I768251);
and I_19741 (I339205,I339188,I768257);
DFFARX1 I_19742 (I339205,I3563,I339154,I339231,);
nor I_19743 (I339122,I339231,I339180);
not I_19744 (I339253,I339231);
DFFARX1 I_19745 (I768242,I3563,I339154,I339279,);
nand I_19746 (I339287,I339279,I768236);
not I_19747 (I339304,I339287);
DFFARX1 I_19748 (I339304,I3563,I339154,I339330,);
not I_19749 (I339146,I339330);
nor I_19750 (I339352,I339180,I339287);
nor I_19751 (I339128,I339231,I339352);
DFFARX1 I_19752 (I768239,I3563,I339154,I339392,);
DFFARX1 I_19753 (I339392,I3563,I339154,I339409,);
not I_19754 (I339417,I339409);
not I_19755 (I339434,I339392);
nand I_19756 (I339131,I339434,I339253);
nand I_19757 (I339465,I768233,I768248);
and I_19758 (I339482,I339465,I768233);
DFFARX1 I_19759 (I339482,I3563,I339154,I339508,);
nor I_19760 (I339516,I339508,I339180);
DFFARX1 I_19761 (I339516,I3563,I339154,I339119,);
DFFARX1 I_19762 (I339508,I3563,I339154,I339137,);
nor I_19763 (I339561,I768254,I768248);
not I_19764 (I339578,I339561);
nor I_19765 (I339140,I339417,I339578);
nand I_19766 (I339125,I339434,I339578);
nor I_19767 (I339134,I339180,I339561);
DFFARX1 I_19768 (I339561,I3563,I339154,I339143,);
not I_19769 (I339681,I3570);
DFFARX1 I_19770 (I1097353,I3563,I339681,I339707,);
nand I_19771 (I339715,I1097368,I1097353);
and I_19772 (I339732,I339715,I1097371);
DFFARX1 I_19773 (I339732,I3563,I339681,I339758,);
nor I_19774 (I339649,I339758,I339707);
not I_19775 (I339780,I339758);
DFFARX1 I_19776 (I1097377,I3563,I339681,I339806,);
nand I_19777 (I339814,I339806,I1097359);
not I_19778 (I339831,I339814);
DFFARX1 I_19779 (I339831,I3563,I339681,I339857,);
not I_19780 (I339673,I339857);
nor I_19781 (I339879,I339707,I339814);
nor I_19782 (I339655,I339758,I339879);
DFFARX1 I_19783 (I1097356,I3563,I339681,I339919,);
DFFARX1 I_19784 (I339919,I3563,I339681,I339936,);
not I_19785 (I339944,I339936);
not I_19786 (I339961,I339919);
nand I_19787 (I339658,I339961,I339780);
nand I_19788 (I339992,I1097356,I1097362);
and I_19789 (I340009,I339992,I1097374);
DFFARX1 I_19790 (I340009,I3563,I339681,I340035,);
nor I_19791 (I340043,I340035,I339707);
DFFARX1 I_19792 (I340043,I3563,I339681,I339646,);
DFFARX1 I_19793 (I340035,I3563,I339681,I339664,);
nor I_19794 (I340088,I1097365,I1097362);
not I_19795 (I340105,I340088);
nor I_19796 (I339667,I339944,I340105);
nand I_19797 (I339652,I339961,I340105);
nor I_19798 (I339661,I339707,I340088);
DFFARX1 I_19799 (I340088,I3563,I339681,I339670,);
not I_19800 (I340208,I3570);
DFFARX1 I_19801 (I199413,I3563,I340208,I340234,);
nand I_19802 (I340242,I199413,I199419);
and I_19803 (I340259,I340242,I199437);
DFFARX1 I_19804 (I340259,I3563,I340208,I340285,);
nor I_19805 (I340176,I340285,I340234);
not I_19806 (I340307,I340285);
DFFARX1 I_19807 (I199425,I3563,I340208,I340333,);
nand I_19808 (I340341,I340333,I199422);
not I_19809 (I340358,I340341);
DFFARX1 I_19810 (I340358,I3563,I340208,I340384,);
not I_19811 (I340200,I340384);
nor I_19812 (I340406,I340234,I340341);
nor I_19813 (I340182,I340285,I340406);
DFFARX1 I_19814 (I199431,I3563,I340208,I340446,);
DFFARX1 I_19815 (I340446,I3563,I340208,I340463,);
not I_19816 (I340471,I340463);
not I_19817 (I340488,I340446);
nand I_19818 (I340185,I340488,I340307);
nand I_19819 (I340519,I199416,I199416);
and I_19820 (I340536,I340519,I199428);
DFFARX1 I_19821 (I340536,I3563,I340208,I340562,);
nor I_19822 (I340570,I340562,I340234);
DFFARX1 I_19823 (I340570,I3563,I340208,I340173,);
DFFARX1 I_19824 (I340562,I3563,I340208,I340191,);
nor I_19825 (I340615,I199434,I199416);
not I_19826 (I340632,I340615);
nor I_19827 (I340194,I340471,I340632);
nand I_19828 (I340179,I340488,I340632);
nor I_19829 (I340188,I340234,I340615);
DFFARX1 I_19830 (I340615,I3563,I340208,I340197,);
not I_19831 (I340735,I3570);
DFFARX1 I_19832 (I1229715,I3563,I340735,I340761,);
nand I_19833 (I340769,I1229730,I1229715);
and I_19834 (I340786,I340769,I1229733);
DFFARX1 I_19835 (I340786,I3563,I340735,I340812,);
nor I_19836 (I340703,I340812,I340761);
not I_19837 (I340834,I340812);
DFFARX1 I_19838 (I1229739,I3563,I340735,I340860,);
nand I_19839 (I340868,I340860,I1229721);
not I_19840 (I340885,I340868);
DFFARX1 I_19841 (I340885,I3563,I340735,I340911,);
not I_19842 (I340727,I340911);
nor I_19843 (I340933,I340761,I340868);
nor I_19844 (I340709,I340812,I340933);
DFFARX1 I_19845 (I1229718,I3563,I340735,I340973,);
DFFARX1 I_19846 (I340973,I3563,I340735,I340990,);
not I_19847 (I340998,I340990);
not I_19848 (I341015,I340973);
nand I_19849 (I340712,I341015,I340834);
nand I_19850 (I341046,I1229718,I1229724);
and I_19851 (I341063,I341046,I1229736);
DFFARX1 I_19852 (I341063,I3563,I340735,I341089,);
nor I_19853 (I341097,I341089,I340761);
DFFARX1 I_19854 (I341097,I3563,I340735,I340700,);
DFFARX1 I_19855 (I341089,I3563,I340735,I340718,);
nor I_19856 (I341142,I1229727,I1229724);
not I_19857 (I341159,I341142);
nor I_19858 (I340721,I340998,I341159);
nand I_19859 (I340706,I341015,I341159);
nor I_19860 (I340715,I340761,I341142);
DFFARX1 I_19861 (I341142,I3563,I340735,I340724,);
not I_19862 (I341262,I3570);
DFFARX1 I_19863 (I1211219,I3563,I341262,I341288,);
nand I_19864 (I341296,I1211234,I1211219);
and I_19865 (I341313,I341296,I1211237);
DFFARX1 I_19866 (I341313,I3563,I341262,I341339,);
nor I_19867 (I341230,I341339,I341288);
not I_19868 (I341361,I341339);
DFFARX1 I_19869 (I1211243,I3563,I341262,I341387,);
nand I_19870 (I341395,I341387,I1211225);
not I_19871 (I341412,I341395);
DFFARX1 I_19872 (I341412,I3563,I341262,I341438,);
not I_19873 (I341254,I341438);
nor I_19874 (I341460,I341288,I341395);
nor I_19875 (I341236,I341339,I341460);
DFFARX1 I_19876 (I1211222,I3563,I341262,I341500,);
DFFARX1 I_19877 (I341500,I3563,I341262,I341517,);
not I_19878 (I341525,I341517);
not I_19879 (I341542,I341500);
nand I_19880 (I341239,I341542,I341361);
nand I_19881 (I341573,I1211222,I1211228);
and I_19882 (I341590,I341573,I1211240);
DFFARX1 I_19883 (I341590,I3563,I341262,I341616,);
nor I_19884 (I341624,I341616,I341288);
DFFARX1 I_19885 (I341624,I3563,I341262,I341227,);
DFFARX1 I_19886 (I341616,I3563,I341262,I341245,);
nor I_19887 (I341669,I1211231,I1211228);
not I_19888 (I341686,I341669);
nor I_19889 (I341248,I341525,I341686);
nand I_19890 (I341233,I341542,I341686);
nor I_19891 (I341242,I341288,I341669);
DFFARX1 I_19892 (I341669,I3563,I341262,I341251,);
not I_19893 (I341789,I3570);
DFFARX1 I_19894 (I802347,I3563,I341789,I341815,);
nand I_19895 (I341823,I802338,I802353);
and I_19896 (I341840,I341823,I802359);
DFFARX1 I_19897 (I341840,I3563,I341789,I341866,);
nor I_19898 (I341757,I341866,I341815);
not I_19899 (I341888,I341866);
DFFARX1 I_19900 (I802344,I3563,I341789,I341914,);
nand I_19901 (I341922,I341914,I802338);
not I_19902 (I341939,I341922);
DFFARX1 I_19903 (I341939,I3563,I341789,I341965,);
not I_19904 (I341781,I341965);
nor I_19905 (I341987,I341815,I341922);
nor I_19906 (I341763,I341866,I341987);
DFFARX1 I_19907 (I802341,I3563,I341789,I342027,);
DFFARX1 I_19908 (I342027,I3563,I341789,I342044,);
not I_19909 (I342052,I342044);
not I_19910 (I342069,I342027);
nand I_19911 (I341766,I342069,I341888);
nand I_19912 (I342100,I802335,I802350);
and I_19913 (I342117,I342100,I802335);
DFFARX1 I_19914 (I342117,I3563,I341789,I342143,);
nor I_19915 (I342151,I342143,I341815);
DFFARX1 I_19916 (I342151,I3563,I341789,I341754,);
DFFARX1 I_19917 (I342143,I3563,I341789,I341772,);
nor I_19918 (I342196,I802356,I802350);
not I_19919 (I342213,I342196);
nor I_19920 (I341775,I342052,I342213);
nand I_19921 (I341760,I342069,I342213);
nor I_19922 (I341769,I341815,I342196);
DFFARX1 I_19923 (I342196,I3563,I341789,I341778,);
not I_19924 (I342316,I3570);
DFFARX1 I_19925 (I146767,I3563,I342316,I342342,);
nand I_19926 (I342350,I146779,I146788);
and I_19927 (I342367,I342350,I146767);
DFFARX1 I_19928 (I342367,I3563,I342316,I342393,);
nor I_19929 (I342284,I342393,I342342);
not I_19930 (I342415,I342393);
DFFARX1 I_19931 (I146782,I3563,I342316,I342441,);
nand I_19932 (I342449,I342441,I146770);
not I_19933 (I342466,I342449);
DFFARX1 I_19934 (I342466,I3563,I342316,I342492,);
not I_19935 (I342308,I342492);
nor I_19936 (I342514,I342342,I342449);
nor I_19937 (I342290,I342393,I342514);
DFFARX1 I_19938 (I146773,I3563,I342316,I342554,);
DFFARX1 I_19939 (I342554,I3563,I342316,I342571,);
not I_19940 (I342579,I342571);
not I_19941 (I342596,I342554);
nand I_19942 (I342293,I342596,I342415);
nand I_19943 (I342627,I146764,I146764);
and I_19944 (I342644,I342627,I146776);
DFFARX1 I_19945 (I342644,I3563,I342316,I342670,);
nor I_19946 (I342678,I342670,I342342);
DFFARX1 I_19947 (I342678,I3563,I342316,I342281,);
DFFARX1 I_19948 (I342670,I3563,I342316,I342299,);
nor I_19949 (I342723,I146785,I146764);
not I_19950 (I342740,I342723);
nor I_19951 (I342302,I342579,I342740);
nand I_19952 (I342287,I342596,I342740);
nor I_19953 (I342296,I342342,I342723);
DFFARX1 I_19954 (I342723,I3563,I342316,I342305,);
not I_19955 (I342843,I3570);
DFFARX1 I_19956 (I67717,I3563,I342843,I342869,);
nand I_19957 (I342877,I67729,I67738);
and I_19958 (I342894,I342877,I67717);
DFFARX1 I_19959 (I342894,I3563,I342843,I342920,);
nor I_19960 (I342811,I342920,I342869);
not I_19961 (I342942,I342920);
DFFARX1 I_19962 (I67732,I3563,I342843,I342968,);
nand I_19963 (I342976,I342968,I67720);
not I_19964 (I342993,I342976);
DFFARX1 I_19965 (I342993,I3563,I342843,I343019,);
not I_19966 (I342835,I343019);
nor I_19967 (I343041,I342869,I342976);
nor I_19968 (I342817,I342920,I343041);
DFFARX1 I_19969 (I67723,I3563,I342843,I343081,);
DFFARX1 I_19970 (I343081,I3563,I342843,I343098,);
not I_19971 (I343106,I343098);
not I_19972 (I343123,I343081);
nand I_19973 (I342820,I343123,I342942);
nand I_19974 (I343154,I67714,I67714);
and I_19975 (I343171,I343154,I67726);
DFFARX1 I_19976 (I343171,I3563,I342843,I343197,);
nor I_19977 (I343205,I343197,I342869);
DFFARX1 I_19978 (I343205,I3563,I342843,I342808,);
DFFARX1 I_19979 (I343197,I3563,I342843,I342826,);
nor I_19980 (I343250,I67735,I67714);
not I_19981 (I343267,I343250);
nor I_19982 (I342829,I343106,I343267);
nand I_19983 (I342814,I343123,I343267);
nor I_19984 (I342823,I342869,I343250);
DFFARX1 I_19985 (I343250,I3563,I342843,I342832,);
not I_19986 (I343370,I3570);
DFFARX1 I_19987 (I582132,I3563,I343370,I343396,);
nand I_19988 (I343404,I582117,I582120);
and I_19989 (I343421,I343404,I582135);
DFFARX1 I_19990 (I343421,I3563,I343370,I343447,);
nor I_19991 (I343338,I343447,I343396);
not I_19992 (I343469,I343447);
DFFARX1 I_19993 (I582129,I3563,I343370,I343495,);
nand I_19994 (I343503,I343495,I582120);
not I_19995 (I343520,I343503);
DFFARX1 I_19996 (I343520,I3563,I343370,I343546,);
not I_19997 (I343362,I343546);
nor I_19998 (I343568,I343396,I343503);
nor I_19999 (I343344,I343447,I343568);
DFFARX1 I_20000 (I582126,I3563,I343370,I343608,);
DFFARX1 I_20001 (I343608,I3563,I343370,I343625,);
not I_20002 (I343633,I343625);
not I_20003 (I343650,I343608);
nand I_20004 (I343347,I343650,I343469);
nand I_20005 (I343681,I582141,I582117);
and I_20006 (I343698,I343681,I582138);
DFFARX1 I_20007 (I343698,I3563,I343370,I343724,);
nor I_20008 (I343732,I343724,I343396);
DFFARX1 I_20009 (I343732,I3563,I343370,I343335,);
DFFARX1 I_20010 (I343724,I3563,I343370,I343353,);
nor I_20011 (I343777,I582123,I582117);
not I_20012 (I343794,I343777);
nor I_20013 (I343356,I343633,I343794);
nand I_20014 (I343341,I343650,I343794);
nor I_20015 (I343350,I343396,I343777);
DFFARX1 I_20016 (I343777,I3563,I343370,I343359,);
not I_20017 (I343897,I3570);
DFFARX1 I_20018 (I1353564,I3563,I343897,I343923,);
nand I_20019 (I343931,I1353543,I1353543);
and I_20020 (I343948,I343931,I1353570);
DFFARX1 I_20021 (I343948,I3563,I343897,I343974,);
nor I_20022 (I343865,I343974,I343923);
not I_20023 (I343996,I343974);
DFFARX1 I_20024 (I1353558,I3563,I343897,I344022,);
nand I_20025 (I344030,I344022,I1353561);
not I_20026 (I344047,I344030);
DFFARX1 I_20027 (I344047,I3563,I343897,I344073,);
not I_20028 (I343889,I344073);
nor I_20029 (I344095,I343923,I344030);
nor I_20030 (I343871,I343974,I344095);
DFFARX1 I_20031 (I1353552,I3563,I343897,I344135,);
DFFARX1 I_20032 (I344135,I3563,I343897,I344152,);
not I_20033 (I344160,I344152);
not I_20034 (I344177,I344135);
nand I_20035 (I343874,I344177,I343996);
nand I_20036 (I344208,I1353549,I1353546);
and I_20037 (I344225,I344208,I1353567);
DFFARX1 I_20038 (I344225,I3563,I343897,I344251,);
nor I_20039 (I344259,I344251,I343923);
DFFARX1 I_20040 (I344259,I3563,I343897,I343862,);
DFFARX1 I_20041 (I344251,I3563,I343897,I343880,);
nor I_20042 (I344304,I1353555,I1353546);
not I_20043 (I344321,I344304);
nor I_20044 (I343883,I344160,I344321);
nand I_20045 (I343868,I344177,I344321);
nor I_20046 (I343877,I343923,I344304);
DFFARX1 I_20047 (I344304,I3563,I343897,I343886,);
not I_20048 (I344424,I3570);
DFFARX1 I_20049 (I171448,I3563,I344424,I344450,);
nand I_20050 (I344458,I171448,I171454);
and I_20051 (I344475,I344458,I171472);
DFFARX1 I_20052 (I344475,I3563,I344424,I344501,);
nor I_20053 (I344392,I344501,I344450);
not I_20054 (I344523,I344501);
DFFARX1 I_20055 (I171460,I3563,I344424,I344549,);
nand I_20056 (I344557,I344549,I171457);
not I_20057 (I344574,I344557);
DFFARX1 I_20058 (I344574,I3563,I344424,I344600,);
not I_20059 (I344416,I344600);
nor I_20060 (I344622,I344450,I344557);
nor I_20061 (I344398,I344501,I344622);
DFFARX1 I_20062 (I171466,I3563,I344424,I344662,);
DFFARX1 I_20063 (I344662,I3563,I344424,I344679,);
not I_20064 (I344687,I344679);
not I_20065 (I344704,I344662);
nand I_20066 (I344401,I344704,I344523);
nand I_20067 (I344735,I171451,I171451);
and I_20068 (I344752,I344735,I171463);
DFFARX1 I_20069 (I344752,I3563,I344424,I344778,);
nor I_20070 (I344786,I344778,I344450);
DFFARX1 I_20071 (I344786,I3563,I344424,I344389,);
DFFARX1 I_20072 (I344778,I3563,I344424,I344407,);
nor I_20073 (I344831,I171469,I171451);
not I_20074 (I344848,I344831);
nor I_20075 (I344410,I344687,I344848);
nand I_20076 (I344395,I344704,I344848);
nor I_20077 (I344404,I344450,I344831);
DFFARX1 I_20078 (I344831,I3563,I344424,I344413,);
not I_20079 (I344951,I3570);
DFFARX1 I_20080 (I79838,I3563,I344951,I344977,);
nand I_20081 (I344985,I79850,I79859);
and I_20082 (I345002,I344985,I79838);
DFFARX1 I_20083 (I345002,I3563,I344951,I345028,);
nor I_20084 (I344919,I345028,I344977);
not I_20085 (I345050,I345028);
DFFARX1 I_20086 (I79853,I3563,I344951,I345076,);
nand I_20087 (I345084,I345076,I79841);
not I_20088 (I345101,I345084);
DFFARX1 I_20089 (I345101,I3563,I344951,I345127,);
not I_20090 (I344943,I345127);
nor I_20091 (I345149,I344977,I345084);
nor I_20092 (I344925,I345028,I345149);
DFFARX1 I_20093 (I79844,I3563,I344951,I345189,);
DFFARX1 I_20094 (I345189,I3563,I344951,I345206,);
not I_20095 (I345214,I345206);
not I_20096 (I345231,I345189);
nand I_20097 (I344928,I345231,I345050);
nand I_20098 (I345262,I79835,I79835);
and I_20099 (I345279,I345262,I79847);
DFFARX1 I_20100 (I345279,I3563,I344951,I345305,);
nor I_20101 (I345313,I345305,I344977);
DFFARX1 I_20102 (I345313,I3563,I344951,I344916,);
DFFARX1 I_20103 (I345305,I3563,I344951,I344934,);
nor I_20104 (I345358,I79856,I79835);
not I_20105 (I345375,I345358);
nor I_20106 (I344937,I345214,I345375);
nand I_20107 (I344922,I345231,I345375);
nor I_20108 (I344931,I344977,I345358);
DFFARX1 I_20109 (I345358,I3563,I344951,I344940,);
not I_20110 (I345478,I3570);
DFFARX1 I_20111 (I1352374,I3563,I345478,I345504,);
nand I_20112 (I345512,I1352353,I1352353);
and I_20113 (I345529,I345512,I1352380);
DFFARX1 I_20114 (I345529,I3563,I345478,I345555,);
nor I_20115 (I345446,I345555,I345504);
not I_20116 (I345577,I345555);
DFFARX1 I_20117 (I1352368,I3563,I345478,I345603,);
nand I_20118 (I345611,I345603,I1352371);
not I_20119 (I345628,I345611);
DFFARX1 I_20120 (I345628,I3563,I345478,I345654,);
not I_20121 (I345470,I345654);
nor I_20122 (I345676,I345504,I345611);
nor I_20123 (I345452,I345555,I345676);
DFFARX1 I_20124 (I1352362,I3563,I345478,I345716,);
DFFARX1 I_20125 (I345716,I3563,I345478,I345733,);
not I_20126 (I345741,I345733);
not I_20127 (I345758,I345716);
nand I_20128 (I345455,I345758,I345577);
nand I_20129 (I345789,I1352359,I1352356);
and I_20130 (I345806,I345789,I1352377);
DFFARX1 I_20131 (I345806,I3563,I345478,I345832,);
nor I_20132 (I345840,I345832,I345504);
DFFARX1 I_20133 (I345840,I3563,I345478,I345443,);
DFFARX1 I_20134 (I345832,I3563,I345478,I345461,);
nor I_20135 (I345885,I1352365,I1352356);
not I_20136 (I345902,I345885);
nor I_20137 (I345464,I345741,I345902);
nand I_20138 (I345449,I345758,I345902);
nor I_20139 (I345458,I345504,I345885);
DFFARX1 I_20140 (I345885,I3563,I345478,I345467,);
not I_20141 (I346005,I3570);
DFFARX1 I_20142 (I874299,I3563,I346005,I346031,);
nand I_20143 (I346039,I874302,I874296);
and I_20144 (I346056,I346039,I874308);
DFFARX1 I_20145 (I346056,I3563,I346005,I346082,);
nor I_20146 (I345973,I346082,I346031);
not I_20147 (I346104,I346082);
DFFARX1 I_20148 (I874311,I3563,I346005,I346130,);
nand I_20149 (I346138,I346130,I874302);
not I_20150 (I346155,I346138);
DFFARX1 I_20151 (I346155,I3563,I346005,I346181,);
not I_20152 (I345997,I346181);
nor I_20153 (I346203,I346031,I346138);
nor I_20154 (I345979,I346082,I346203);
DFFARX1 I_20155 (I874314,I3563,I346005,I346243,);
DFFARX1 I_20156 (I346243,I3563,I346005,I346260,);
not I_20157 (I346268,I346260);
not I_20158 (I346285,I346243);
nand I_20159 (I345982,I346285,I346104);
nand I_20160 (I346316,I874296,I874305);
and I_20161 (I346333,I346316,I874299);
DFFARX1 I_20162 (I346333,I3563,I346005,I346359,);
nor I_20163 (I346367,I346359,I346031);
DFFARX1 I_20164 (I346367,I3563,I346005,I345970,);
DFFARX1 I_20165 (I346359,I3563,I346005,I345988,);
nor I_20166 (I346412,I874317,I874305);
not I_20167 (I346429,I346412);
nor I_20168 (I345991,I346268,I346429);
nand I_20169 (I345976,I346285,I346429);
nor I_20170 (I345985,I346031,I346412);
DFFARX1 I_20171 (I346412,I3563,I346005,I345994,);
not I_20172 (I346532,I3570);
DFFARX1 I_20173 (I980770,I3563,I346532,I346558,);
nand I_20174 (I346566,I980767,I980785);
and I_20175 (I346583,I346566,I980776);
DFFARX1 I_20176 (I346583,I3563,I346532,I346609,);
nor I_20177 (I346500,I346609,I346558);
not I_20178 (I346631,I346609);
DFFARX1 I_20179 (I980791,I3563,I346532,I346657,);
nand I_20180 (I346665,I346657,I980773);
not I_20181 (I346682,I346665);
DFFARX1 I_20182 (I346682,I3563,I346532,I346708,);
not I_20183 (I346524,I346708);
nor I_20184 (I346730,I346558,I346665);
nor I_20185 (I346506,I346609,I346730);
DFFARX1 I_20186 (I980779,I3563,I346532,I346770,);
DFFARX1 I_20187 (I346770,I3563,I346532,I346787,);
not I_20188 (I346795,I346787);
not I_20189 (I346812,I346770);
nand I_20190 (I346509,I346812,I346631);
nand I_20191 (I346843,I980767,I980794);
and I_20192 (I346860,I346843,I980782);
DFFARX1 I_20193 (I346860,I3563,I346532,I346886,);
nor I_20194 (I346894,I346886,I346558);
DFFARX1 I_20195 (I346894,I3563,I346532,I346497,);
DFFARX1 I_20196 (I346886,I3563,I346532,I346515,);
nor I_20197 (I346939,I980788,I980794);
not I_20198 (I346956,I346939);
nor I_20199 (I346518,I346795,I346956);
nand I_20200 (I346503,I346812,I346956);
nor I_20201 (I346512,I346558,I346939);
DFFARX1 I_20202 (I346939,I3563,I346532,I346521,);
not I_20203 (I347059,I3570);
DFFARX1 I_20204 (I1172493,I3563,I347059,I347085,);
nand I_20205 (I347093,I1172508,I1172493);
and I_20206 (I347110,I347093,I1172511);
DFFARX1 I_20207 (I347110,I3563,I347059,I347136,);
nor I_20208 (I347027,I347136,I347085);
not I_20209 (I347158,I347136);
DFFARX1 I_20210 (I1172517,I3563,I347059,I347184,);
nand I_20211 (I347192,I347184,I1172499);
not I_20212 (I347209,I347192);
DFFARX1 I_20213 (I347209,I3563,I347059,I347235,);
not I_20214 (I347051,I347235);
nor I_20215 (I347257,I347085,I347192);
nor I_20216 (I347033,I347136,I347257);
DFFARX1 I_20217 (I1172496,I3563,I347059,I347297,);
DFFARX1 I_20218 (I347297,I3563,I347059,I347314,);
not I_20219 (I347322,I347314);
not I_20220 (I347339,I347297);
nand I_20221 (I347036,I347339,I347158);
nand I_20222 (I347370,I1172496,I1172502);
and I_20223 (I347387,I347370,I1172514);
DFFARX1 I_20224 (I347387,I3563,I347059,I347413,);
nor I_20225 (I347421,I347413,I347085);
DFFARX1 I_20226 (I347421,I3563,I347059,I347024,);
DFFARX1 I_20227 (I347413,I3563,I347059,I347042,);
nor I_20228 (I347466,I1172505,I1172502);
not I_20229 (I347483,I347466);
nor I_20230 (I347045,I347322,I347483);
nand I_20231 (I347030,I347339,I347483);
nor I_20232 (I347039,I347085,I347466);
DFFARX1 I_20233 (I347466,I3563,I347059,I347048,);
not I_20234 (I347586,I3570);
DFFARX1 I_20235 (I103026,I3563,I347586,I347612,);
nand I_20236 (I347620,I103038,I103047);
and I_20237 (I347637,I347620,I103026);
DFFARX1 I_20238 (I347637,I3563,I347586,I347663,);
nor I_20239 (I347554,I347663,I347612);
not I_20240 (I347685,I347663);
DFFARX1 I_20241 (I103041,I3563,I347586,I347711,);
nand I_20242 (I347719,I347711,I103029);
not I_20243 (I347736,I347719);
DFFARX1 I_20244 (I347736,I3563,I347586,I347762,);
not I_20245 (I347578,I347762);
nor I_20246 (I347784,I347612,I347719);
nor I_20247 (I347560,I347663,I347784);
DFFARX1 I_20248 (I103032,I3563,I347586,I347824,);
DFFARX1 I_20249 (I347824,I3563,I347586,I347841,);
not I_20250 (I347849,I347841);
not I_20251 (I347866,I347824);
nand I_20252 (I347563,I347866,I347685);
nand I_20253 (I347897,I103023,I103023);
and I_20254 (I347914,I347897,I103035);
DFFARX1 I_20255 (I347914,I3563,I347586,I347940,);
nor I_20256 (I347948,I347940,I347612);
DFFARX1 I_20257 (I347948,I3563,I347586,I347551,);
DFFARX1 I_20258 (I347940,I3563,I347586,I347569,);
nor I_20259 (I347993,I103044,I103023);
not I_20260 (I348010,I347993);
nor I_20261 (I347572,I347849,I348010);
nand I_20262 (I347557,I347866,I348010);
nor I_20263 (I347566,I347612,I347993);
DFFARX1 I_20264 (I347993,I3563,I347586,I347575,);
not I_20265 (I348113,I3570);
DFFARX1 I_20266 (I1060687,I3563,I348113,I348139,);
nand I_20267 (I348147,I1060684,I1060687);
and I_20268 (I348164,I348147,I1060696);
DFFARX1 I_20269 (I348164,I3563,I348113,I348190,);
nor I_20270 (I348081,I348190,I348139);
not I_20271 (I348212,I348190);
DFFARX1 I_20272 (I1060684,I3563,I348113,I348238,);
nand I_20273 (I348246,I348238,I1060702);
not I_20274 (I348263,I348246);
DFFARX1 I_20275 (I348263,I3563,I348113,I348289,);
not I_20276 (I348105,I348289);
nor I_20277 (I348311,I348139,I348246);
nor I_20278 (I348087,I348190,I348311);
DFFARX1 I_20279 (I1060690,I3563,I348113,I348351,);
DFFARX1 I_20280 (I348351,I3563,I348113,I348368,);
not I_20281 (I348376,I348368);
not I_20282 (I348393,I348351);
nand I_20283 (I348090,I348393,I348212);
nand I_20284 (I348424,I1060699,I1060705);
and I_20285 (I348441,I348424,I1060690);
DFFARX1 I_20286 (I348441,I3563,I348113,I348467,);
nor I_20287 (I348475,I348467,I348139);
DFFARX1 I_20288 (I348475,I3563,I348113,I348078,);
DFFARX1 I_20289 (I348467,I3563,I348113,I348096,);
nor I_20290 (I348520,I1060693,I1060705);
not I_20291 (I348537,I348520);
nor I_20292 (I348099,I348376,I348537);
nand I_20293 (I348084,I348393,I348537);
nor I_20294 (I348093,I348139,I348520);
DFFARX1 I_20295 (I348520,I3563,I348113,I348102,);
not I_20296 (I348640,I3570);
DFFARX1 I_20297 (I1068541,I3563,I348640,I348666,);
nand I_20298 (I348674,I1068538,I1068541);
and I_20299 (I348691,I348674,I1068550);
DFFARX1 I_20300 (I348691,I3563,I348640,I348717,);
nor I_20301 (I348608,I348717,I348666);
not I_20302 (I348739,I348717);
DFFARX1 I_20303 (I1068538,I3563,I348640,I348765,);
nand I_20304 (I348773,I348765,I1068556);
not I_20305 (I348790,I348773);
DFFARX1 I_20306 (I348790,I3563,I348640,I348816,);
not I_20307 (I348632,I348816);
nor I_20308 (I348838,I348666,I348773);
nor I_20309 (I348614,I348717,I348838);
DFFARX1 I_20310 (I1068544,I3563,I348640,I348878,);
DFFARX1 I_20311 (I348878,I3563,I348640,I348895,);
not I_20312 (I348903,I348895);
not I_20313 (I348920,I348878);
nand I_20314 (I348617,I348920,I348739);
nand I_20315 (I348951,I1068553,I1068559);
and I_20316 (I348968,I348951,I1068544);
DFFARX1 I_20317 (I348968,I3563,I348640,I348994,);
nor I_20318 (I349002,I348994,I348666);
DFFARX1 I_20319 (I349002,I3563,I348640,I348605,);
DFFARX1 I_20320 (I348994,I3563,I348640,I348623,);
nor I_20321 (I349047,I1068547,I1068559);
not I_20322 (I349064,I349047);
nor I_20323 (I348626,I348903,I349064);
nand I_20324 (I348611,I348920,I349064);
nor I_20325 (I348620,I348666,I349047);
DFFARX1 I_20326 (I349047,I3563,I348640,I348629,);
not I_20327 (I349167,I3570);
DFFARX1 I_20328 (I507278,I3563,I349167,I349193,);
nand I_20329 (I349201,I507290,I507269);
and I_20330 (I349218,I349201,I507293);
DFFARX1 I_20331 (I349218,I3563,I349167,I349244,);
nor I_20332 (I349135,I349244,I349193);
not I_20333 (I349266,I349244);
DFFARX1 I_20334 (I507284,I3563,I349167,I349292,);
nand I_20335 (I349300,I349292,I507266);
not I_20336 (I349317,I349300);
DFFARX1 I_20337 (I349317,I3563,I349167,I349343,);
not I_20338 (I349159,I349343);
nor I_20339 (I349365,I349193,I349300);
nor I_20340 (I349141,I349244,I349365);
DFFARX1 I_20341 (I507281,I3563,I349167,I349405,);
DFFARX1 I_20342 (I349405,I3563,I349167,I349422,);
not I_20343 (I349430,I349422);
not I_20344 (I349447,I349405);
nand I_20345 (I349144,I349447,I349266);
nand I_20346 (I349478,I507266,I507272);
and I_20347 (I349495,I349478,I507275);
DFFARX1 I_20348 (I349495,I3563,I349167,I349521,);
nor I_20349 (I349529,I349521,I349193);
DFFARX1 I_20350 (I349529,I3563,I349167,I349132,);
DFFARX1 I_20351 (I349521,I3563,I349167,I349150,);
nor I_20352 (I349574,I507287,I507272);
not I_20353 (I349591,I349574);
nor I_20354 (I349153,I349430,I349591);
nand I_20355 (I349138,I349447,I349591);
nor I_20356 (I349147,I349193,I349574);
DFFARX1 I_20357 (I349574,I3563,I349167,I349156,);
not I_20358 (I349694,I3570);
DFFARX1 I_20359 (I864286,I3563,I349694,I349720,);
nand I_20360 (I349728,I864289,I864283);
and I_20361 (I349745,I349728,I864295);
DFFARX1 I_20362 (I349745,I3563,I349694,I349771,);
nor I_20363 (I349662,I349771,I349720);
not I_20364 (I349793,I349771);
DFFARX1 I_20365 (I864298,I3563,I349694,I349819,);
nand I_20366 (I349827,I349819,I864289);
not I_20367 (I349844,I349827);
DFFARX1 I_20368 (I349844,I3563,I349694,I349870,);
not I_20369 (I349686,I349870);
nor I_20370 (I349892,I349720,I349827);
nor I_20371 (I349668,I349771,I349892);
DFFARX1 I_20372 (I864301,I3563,I349694,I349932,);
DFFARX1 I_20373 (I349932,I3563,I349694,I349949,);
not I_20374 (I349957,I349949);
not I_20375 (I349974,I349932);
nand I_20376 (I349671,I349974,I349793);
nand I_20377 (I350005,I864283,I864292);
and I_20378 (I350022,I350005,I864286);
DFFARX1 I_20379 (I350022,I3563,I349694,I350048,);
nor I_20380 (I350056,I350048,I349720);
DFFARX1 I_20381 (I350056,I3563,I349694,I349659,);
DFFARX1 I_20382 (I350048,I3563,I349694,I349677,);
nor I_20383 (I350101,I864304,I864292);
not I_20384 (I350118,I350101);
nor I_20385 (I349680,I349957,I350118);
nand I_20386 (I349665,I349974,I350118);
nor I_20387 (I349674,I349720,I350101);
DFFARX1 I_20388 (I350101,I3563,I349694,I349683,);
not I_20389 (I350221,I3570);
DFFARX1 I_20390 (I613344,I3563,I350221,I350247,);
nand I_20391 (I350255,I613329,I613332);
and I_20392 (I350272,I350255,I613347);
DFFARX1 I_20393 (I350272,I3563,I350221,I350298,);
nor I_20394 (I350189,I350298,I350247);
not I_20395 (I350320,I350298);
DFFARX1 I_20396 (I613341,I3563,I350221,I350346,);
nand I_20397 (I350354,I350346,I613332);
not I_20398 (I350371,I350354);
DFFARX1 I_20399 (I350371,I3563,I350221,I350397,);
not I_20400 (I350213,I350397);
nor I_20401 (I350419,I350247,I350354);
nor I_20402 (I350195,I350298,I350419);
DFFARX1 I_20403 (I613338,I3563,I350221,I350459,);
DFFARX1 I_20404 (I350459,I3563,I350221,I350476,);
not I_20405 (I350484,I350476);
not I_20406 (I350501,I350459);
nand I_20407 (I350198,I350501,I350320);
nand I_20408 (I350532,I613353,I613329);
and I_20409 (I350549,I350532,I613350);
DFFARX1 I_20410 (I350549,I3563,I350221,I350575,);
nor I_20411 (I350583,I350575,I350247);
DFFARX1 I_20412 (I350583,I3563,I350221,I350186,);
DFFARX1 I_20413 (I350575,I3563,I350221,I350204,);
nor I_20414 (I350628,I613335,I613329);
not I_20415 (I350645,I350628);
nor I_20416 (I350207,I350484,I350645);
nand I_20417 (I350192,I350501,I350645);
nor I_20418 (I350201,I350247,I350628);
DFFARX1 I_20419 (I350628,I3563,I350221,I350210,);
not I_20420 (I350748,I3570);
DFFARX1 I_20421 (I1290080,I3563,I350748,I350774,);
nand I_20422 (I350782,I1290077,I1290068);
and I_20423 (I350799,I350782,I1290065);
DFFARX1 I_20424 (I350799,I3563,I350748,I350825,);
nor I_20425 (I350716,I350825,I350774);
not I_20426 (I350847,I350825);
DFFARX1 I_20427 (I1290074,I3563,I350748,I350873,);
nand I_20428 (I350881,I350873,I1290083);
not I_20429 (I350898,I350881);
DFFARX1 I_20430 (I350898,I3563,I350748,I350924,);
not I_20431 (I350740,I350924);
nor I_20432 (I350946,I350774,I350881);
nor I_20433 (I350722,I350825,I350946);
DFFARX1 I_20434 (I1290086,I3563,I350748,I350986,);
DFFARX1 I_20435 (I350986,I3563,I350748,I351003,);
not I_20436 (I351011,I351003);
not I_20437 (I351028,I350986);
nand I_20438 (I350725,I351028,I350847);
nand I_20439 (I351059,I1290065,I1290071);
and I_20440 (I351076,I351059,I1290089);
DFFARX1 I_20441 (I351076,I3563,I350748,I351102,);
nor I_20442 (I351110,I351102,I350774);
DFFARX1 I_20443 (I351110,I3563,I350748,I350713,);
DFFARX1 I_20444 (I351102,I3563,I350748,I350731,);
nor I_20445 (I351155,I1290068,I1290071);
not I_20446 (I351172,I351155);
nor I_20447 (I350734,I351011,I351172);
nand I_20448 (I350719,I351028,I351172);
nor I_20449 (I350728,I350774,I351155);
DFFARX1 I_20450 (I351155,I3563,I350748,I350737,);
not I_20451 (I351275,I3570);
DFFARX1 I_20452 (I779227,I3563,I351275,I351301,);
nand I_20453 (I351309,I779218,I779233);
and I_20454 (I351326,I351309,I779239);
DFFARX1 I_20455 (I351326,I3563,I351275,I351352,);
nor I_20456 (I351243,I351352,I351301);
not I_20457 (I351374,I351352);
DFFARX1 I_20458 (I779224,I3563,I351275,I351400,);
nand I_20459 (I351408,I351400,I779218);
not I_20460 (I351425,I351408);
DFFARX1 I_20461 (I351425,I3563,I351275,I351451,);
not I_20462 (I351267,I351451);
nor I_20463 (I351473,I351301,I351408);
nor I_20464 (I351249,I351352,I351473);
DFFARX1 I_20465 (I779221,I3563,I351275,I351513,);
DFFARX1 I_20466 (I351513,I3563,I351275,I351530,);
not I_20467 (I351538,I351530);
not I_20468 (I351555,I351513);
nand I_20469 (I351252,I351555,I351374);
nand I_20470 (I351586,I779215,I779230);
and I_20471 (I351603,I351586,I779215);
DFFARX1 I_20472 (I351603,I3563,I351275,I351629,);
nor I_20473 (I351637,I351629,I351301);
DFFARX1 I_20474 (I351637,I3563,I351275,I351240,);
DFFARX1 I_20475 (I351629,I3563,I351275,I351258,);
nor I_20476 (I351682,I779236,I779230);
not I_20477 (I351699,I351682);
nor I_20478 (I351261,I351538,I351699);
nand I_20479 (I351246,I351555,I351699);
nor I_20480 (I351255,I351301,I351682);
DFFARX1 I_20481 (I351682,I3563,I351275,I351264,);
not I_20482 (I351802,I3570);
DFFARX1 I_20483 (I618546,I3563,I351802,I351828,);
nand I_20484 (I351836,I618531,I618534);
and I_20485 (I351853,I351836,I618549);
DFFARX1 I_20486 (I351853,I3563,I351802,I351879,);
nor I_20487 (I351770,I351879,I351828);
not I_20488 (I351901,I351879);
DFFARX1 I_20489 (I618543,I3563,I351802,I351927,);
nand I_20490 (I351935,I351927,I618534);
not I_20491 (I351952,I351935);
DFFARX1 I_20492 (I351952,I3563,I351802,I351978,);
not I_20493 (I351794,I351978);
nor I_20494 (I352000,I351828,I351935);
nor I_20495 (I351776,I351879,I352000);
DFFARX1 I_20496 (I618540,I3563,I351802,I352040,);
DFFARX1 I_20497 (I352040,I3563,I351802,I352057,);
not I_20498 (I352065,I352057);
not I_20499 (I352082,I352040);
nand I_20500 (I351779,I352082,I351901);
nand I_20501 (I352113,I618555,I618531);
and I_20502 (I352130,I352113,I618552);
DFFARX1 I_20503 (I352130,I3563,I351802,I352156,);
nor I_20504 (I352164,I352156,I351828);
DFFARX1 I_20505 (I352164,I3563,I351802,I351767,);
DFFARX1 I_20506 (I352156,I3563,I351802,I351785,);
nor I_20507 (I352209,I618537,I618531);
not I_20508 (I352226,I352209);
nor I_20509 (I351788,I352065,I352226);
nand I_20510 (I351773,I352082,I352226);
nor I_20511 (I351782,I351828,I352209);
DFFARX1 I_20512 (I352209,I3563,I351802,I351791,);
not I_20513 (I352329,I3570);
DFFARX1 I_20514 (I1054516,I3563,I352329,I352355,);
nand I_20515 (I352363,I1054513,I1054516);
and I_20516 (I352380,I352363,I1054525);
DFFARX1 I_20517 (I352380,I3563,I352329,I352406,);
nor I_20518 (I352297,I352406,I352355);
not I_20519 (I352428,I352406);
DFFARX1 I_20520 (I1054513,I3563,I352329,I352454,);
nand I_20521 (I352462,I352454,I1054531);
not I_20522 (I352479,I352462);
DFFARX1 I_20523 (I352479,I3563,I352329,I352505,);
not I_20524 (I352321,I352505);
nor I_20525 (I352527,I352355,I352462);
nor I_20526 (I352303,I352406,I352527);
DFFARX1 I_20527 (I1054519,I3563,I352329,I352567,);
DFFARX1 I_20528 (I352567,I3563,I352329,I352584,);
not I_20529 (I352592,I352584);
not I_20530 (I352609,I352567);
nand I_20531 (I352306,I352609,I352428);
nand I_20532 (I352640,I1054528,I1054534);
and I_20533 (I352657,I352640,I1054519);
DFFARX1 I_20534 (I352657,I3563,I352329,I352683,);
nor I_20535 (I352691,I352683,I352355);
DFFARX1 I_20536 (I352691,I3563,I352329,I352294,);
DFFARX1 I_20537 (I352683,I3563,I352329,I352312,);
nor I_20538 (I352736,I1054522,I1054534);
not I_20539 (I352753,I352736);
nor I_20540 (I352315,I352592,I352753);
nand I_20541 (I352300,I352609,I352753);
nor I_20542 (I352309,I352355,I352736);
DFFARX1 I_20543 (I352736,I3563,I352329,I352318,);
not I_20544 (I352856,I3570);
DFFARX1 I_20545 (I1177117,I3563,I352856,I352882,);
nand I_20546 (I352890,I1177132,I1177117);
and I_20547 (I352907,I352890,I1177135);
DFFARX1 I_20548 (I352907,I3563,I352856,I352933,);
nor I_20549 (I352824,I352933,I352882);
not I_20550 (I352955,I352933);
DFFARX1 I_20551 (I1177141,I3563,I352856,I352981,);
nand I_20552 (I352989,I352981,I1177123);
not I_20553 (I353006,I352989);
DFFARX1 I_20554 (I353006,I3563,I352856,I353032,);
not I_20555 (I352848,I353032);
nor I_20556 (I353054,I352882,I352989);
nor I_20557 (I352830,I352933,I353054);
DFFARX1 I_20558 (I1177120,I3563,I352856,I353094,);
DFFARX1 I_20559 (I353094,I3563,I352856,I353111,);
not I_20560 (I353119,I353111);
not I_20561 (I353136,I353094);
nand I_20562 (I352833,I353136,I352955);
nand I_20563 (I353167,I1177120,I1177126);
and I_20564 (I353184,I353167,I1177138);
DFFARX1 I_20565 (I353184,I3563,I352856,I353210,);
nor I_20566 (I353218,I353210,I352882);
DFFARX1 I_20567 (I353218,I3563,I352856,I352821,);
DFFARX1 I_20568 (I353210,I3563,I352856,I352839,);
nor I_20569 (I353263,I1177129,I1177126);
not I_20570 (I353280,I353263);
nor I_20571 (I352842,I353119,I353280);
nand I_20572 (I352827,I353136,I353280);
nor I_20573 (I352836,I352882,I353263);
DFFARX1 I_20574 (I353263,I3563,I352856,I352845,);
not I_20575 (I353383,I3570);
DFFARX1 I_20576 (I1109491,I3563,I353383,I353409,);
nand I_20577 (I353417,I1109506,I1109491);
and I_20578 (I353434,I353417,I1109509);
DFFARX1 I_20579 (I353434,I3563,I353383,I353460,);
nor I_20580 (I353351,I353460,I353409);
not I_20581 (I353482,I353460);
DFFARX1 I_20582 (I1109515,I3563,I353383,I353508,);
nand I_20583 (I353516,I353508,I1109497);
not I_20584 (I353533,I353516);
DFFARX1 I_20585 (I353533,I3563,I353383,I353559,);
not I_20586 (I353375,I353559);
nor I_20587 (I353581,I353409,I353516);
nor I_20588 (I353357,I353460,I353581);
DFFARX1 I_20589 (I1109494,I3563,I353383,I353621,);
DFFARX1 I_20590 (I353621,I3563,I353383,I353638,);
not I_20591 (I353646,I353638);
not I_20592 (I353663,I353621);
nand I_20593 (I353360,I353663,I353482);
nand I_20594 (I353694,I1109494,I1109500);
and I_20595 (I353711,I353694,I1109512);
DFFARX1 I_20596 (I353711,I3563,I353383,I353737,);
nor I_20597 (I353745,I353737,I353409);
DFFARX1 I_20598 (I353745,I3563,I353383,I353348,);
DFFARX1 I_20599 (I353737,I3563,I353383,I353366,);
nor I_20600 (I353790,I1109503,I1109500);
not I_20601 (I353807,I353790);
nor I_20602 (I353369,I353646,I353807);
nand I_20603 (I353354,I353663,I353807);
nor I_20604 (I353363,I353409,I353790);
DFFARX1 I_20605 (I353790,I3563,I353383,I353372,);
not I_20606 (I353910,I3570);
DFFARX1 I_20607 (I596004,I3563,I353910,I353936,);
nand I_20608 (I353944,I595989,I595992);
and I_20609 (I353961,I353944,I596007);
DFFARX1 I_20610 (I353961,I3563,I353910,I353987,);
nor I_20611 (I353878,I353987,I353936);
not I_20612 (I354009,I353987);
DFFARX1 I_20613 (I596001,I3563,I353910,I354035,);
nand I_20614 (I354043,I354035,I595992);
not I_20615 (I354060,I354043);
DFFARX1 I_20616 (I354060,I3563,I353910,I354086,);
not I_20617 (I353902,I354086);
nor I_20618 (I354108,I353936,I354043);
nor I_20619 (I353884,I353987,I354108);
DFFARX1 I_20620 (I595998,I3563,I353910,I354148,);
DFFARX1 I_20621 (I354148,I3563,I353910,I354165,);
not I_20622 (I354173,I354165);
not I_20623 (I354190,I354148);
nand I_20624 (I353887,I354190,I354009);
nand I_20625 (I354221,I596013,I595989);
and I_20626 (I354238,I354221,I596010);
DFFARX1 I_20627 (I354238,I3563,I353910,I354264,);
nor I_20628 (I354272,I354264,I353936);
DFFARX1 I_20629 (I354272,I3563,I353910,I353875,);
DFFARX1 I_20630 (I354264,I3563,I353910,I353893,);
nor I_20631 (I354317,I595995,I595989);
not I_20632 (I354334,I354317);
nor I_20633 (I353896,I354173,I354334);
nand I_20634 (I353881,I354190,I354334);
nor I_20635 (I353890,I353936,I354317);
DFFARX1 I_20636 (I354317,I3563,I353910,I353899,);
not I_20637 (I354437,I3570);
DFFARX1 I_20638 (I212503,I3563,I354437,I354463,);
nand I_20639 (I354471,I212503,I212509);
and I_20640 (I354488,I354471,I212527);
DFFARX1 I_20641 (I354488,I3563,I354437,I354514,);
nor I_20642 (I354405,I354514,I354463);
not I_20643 (I354536,I354514);
DFFARX1 I_20644 (I212515,I3563,I354437,I354562,);
nand I_20645 (I354570,I354562,I212512);
not I_20646 (I354587,I354570);
DFFARX1 I_20647 (I354587,I3563,I354437,I354613,);
not I_20648 (I354429,I354613);
nor I_20649 (I354635,I354463,I354570);
nor I_20650 (I354411,I354514,I354635);
DFFARX1 I_20651 (I212521,I3563,I354437,I354675,);
DFFARX1 I_20652 (I354675,I3563,I354437,I354692,);
not I_20653 (I354700,I354692);
not I_20654 (I354717,I354675);
nand I_20655 (I354414,I354717,I354536);
nand I_20656 (I354748,I212506,I212506);
and I_20657 (I354765,I354748,I212518);
DFFARX1 I_20658 (I354765,I3563,I354437,I354791,);
nor I_20659 (I354799,I354791,I354463);
DFFARX1 I_20660 (I354799,I3563,I354437,I354402,);
DFFARX1 I_20661 (I354791,I3563,I354437,I354420,);
nor I_20662 (I354844,I212524,I212506);
not I_20663 (I354861,I354844);
nor I_20664 (I354423,I354700,I354861);
nand I_20665 (I354408,I354717,I354861);
nor I_20666 (I354417,I354463,I354844);
DFFARX1 I_20667 (I354844,I3563,I354437,I354426,);
not I_20668 (I354964,I3570);
DFFARX1 I_20669 (I259508,I3563,I354964,I354990,);
nand I_20670 (I354998,I259508,I259514);
and I_20671 (I355015,I354998,I259532);
DFFARX1 I_20672 (I355015,I3563,I354964,I355041,);
nor I_20673 (I354932,I355041,I354990);
not I_20674 (I355063,I355041);
DFFARX1 I_20675 (I259520,I3563,I354964,I355089,);
nand I_20676 (I355097,I355089,I259517);
not I_20677 (I355114,I355097);
DFFARX1 I_20678 (I355114,I3563,I354964,I355140,);
not I_20679 (I354956,I355140);
nor I_20680 (I355162,I354990,I355097);
nor I_20681 (I354938,I355041,I355162);
DFFARX1 I_20682 (I259526,I3563,I354964,I355202,);
DFFARX1 I_20683 (I355202,I3563,I354964,I355219,);
not I_20684 (I355227,I355219);
not I_20685 (I355244,I355202);
nand I_20686 (I354941,I355244,I355063);
nand I_20687 (I355275,I259511,I259511);
and I_20688 (I355292,I355275,I259523);
DFFARX1 I_20689 (I355292,I3563,I354964,I355318,);
nor I_20690 (I355326,I355318,I354990);
DFFARX1 I_20691 (I355326,I3563,I354964,I354929,);
DFFARX1 I_20692 (I355318,I3563,I354964,I354947,);
nor I_20693 (I355371,I259529,I259511);
not I_20694 (I355388,I355371);
nor I_20695 (I354950,I355227,I355388);
nand I_20696 (I354935,I355244,I355388);
nor I_20697 (I354944,I354990,I355371);
DFFARX1 I_20698 (I355371,I3563,I354964,I354953,);
not I_20699 (I355491,I3570);
DFFARX1 I_20700 (I29243,I3563,I355491,I355517,);
nand I_20701 (I355525,I29267,I29246);
and I_20702 (I355542,I355525,I29243);
DFFARX1 I_20703 (I355542,I3563,I355491,I355568,);
nor I_20704 (I355459,I355568,I355517);
not I_20705 (I355590,I355568);
DFFARX1 I_20706 (I29249,I3563,I355491,I355616,);
nand I_20707 (I355624,I355616,I29258);
not I_20708 (I355641,I355624);
DFFARX1 I_20709 (I355641,I3563,I355491,I355667,);
not I_20710 (I355483,I355667);
nor I_20711 (I355689,I355517,I355624);
nor I_20712 (I355465,I355568,I355689);
DFFARX1 I_20713 (I29252,I3563,I355491,I355729,);
DFFARX1 I_20714 (I355729,I3563,I355491,I355746,);
not I_20715 (I355754,I355746);
not I_20716 (I355771,I355729);
nand I_20717 (I355468,I355771,I355590);
nand I_20718 (I355802,I29264,I29246);
and I_20719 (I355819,I355802,I29255);
DFFARX1 I_20720 (I355819,I3563,I355491,I355845,);
nor I_20721 (I355853,I355845,I355517);
DFFARX1 I_20722 (I355853,I3563,I355491,I355456,);
DFFARX1 I_20723 (I355845,I3563,I355491,I355474,);
nor I_20724 (I355898,I29261,I29246);
not I_20725 (I355915,I355898);
nor I_20726 (I355477,I355754,I355915);
nand I_20727 (I355462,I355771,I355915);
nor I_20728 (I355471,I355517,I355898);
DFFARX1 I_20729 (I355898,I3563,I355491,I355480,);
not I_20730 (I356018,I3570);
DFFARX1 I_20731 (I774025,I3563,I356018,I356044,);
nand I_20732 (I356052,I774016,I774031);
and I_20733 (I356069,I356052,I774037);
DFFARX1 I_20734 (I356069,I3563,I356018,I356095,);
nor I_20735 (I355986,I356095,I356044);
not I_20736 (I356117,I356095);
DFFARX1 I_20737 (I774022,I3563,I356018,I356143,);
nand I_20738 (I356151,I356143,I774016);
not I_20739 (I356168,I356151);
DFFARX1 I_20740 (I356168,I3563,I356018,I356194,);
not I_20741 (I356010,I356194);
nor I_20742 (I356216,I356044,I356151);
nor I_20743 (I355992,I356095,I356216);
DFFARX1 I_20744 (I774019,I3563,I356018,I356256,);
DFFARX1 I_20745 (I356256,I3563,I356018,I356273,);
not I_20746 (I356281,I356273);
not I_20747 (I356298,I356256);
nand I_20748 (I355995,I356298,I356117);
nand I_20749 (I356329,I774013,I774028);
and I_20750 (I356346,I356329,I774013);
DFFARX1 I_20751 (I356346,I3563,I356018,I356372,);
nor I_20752 (I356380,I356372,I356044);
DFFARX1 I_20753 (I356380,I3563,I356018,I355983,);
DFFARX1 I_20754 (I356372,I3563,I356018,I356001,);
nor I_20755 (I356425,I774034,I774028);
not I_20756 (I356442,I356425);
nor I_20757 (I356004,I356281,I356442);
nand I_20758 (I355989,I356298,I356442);
nor I_20759 (I355998,I356044,I356425);
DFFARX1 I_20760 (I356425,I3563,I356018,I356007,);
not I_20761 (I356545,I3570);
DFFARX1 I_20762 (I1090995,I3563,I356545,I356571,);
nand I_20763 (I356579,I1091010,I1090995);
and I_20764 (I356596,I356579,I1091013);
DFFARX1 I_20765 (I356596,I3563,I356545,I356622,);
nor I_20766 (I356513,I356622,I356571);
not I_20767 (I356644,I356622);
DFFARX1 I_20768 (I1091019,I3563,I356545,I356670,);
nand I_20769 (I356678,I356670,I1091001);
not I_20770 (I356695,I356678);
DFFARX1 I_20771 (I356695,I3563,I356545,I356721,);
not I_20772 (I356537,I356721);
nor I_20773 (I356743,I356571,I356678);
nor I_20774 (I356519,I356622,I356743);
DFFARX1 I_20775 (I1090998,I3563,I356545,I356783,);
DFFARX1 I_20776 (I356783,I3563,I356545,I356800,);
not I_20777 (I356808,I356800);
not I_20778 (I356825,I356783);
nand I_20779 (I356522,I356825,I356644);
nand I_20780 (I356856,I1090998,I1091004);
and I_20781 (I356873,I356856,I1091016);
DFFARX1 I_20782 (I356873,I3563,I356545,I356899,);
nor I_20783 (I356907,I356899,I356571);
DFFARX1 I_20784 (I356907,I3563,I356545,I356510,);
DFFARX1 I_20785 (I356899,I3563,I356545,I356528,);
nor I_20786 (I356952,I1091007,I1091004);
not I_20787 (I356969,I356952);
nor I_20788 (I356531,I356808,I356969);
nand I_20789 (I356516,I356825,I356969);
nor I_20790 (I356525,I356571,I356952);
DFFARX1 I_20791 (I356952,I3563,I356545,I356534,);
not I_20792 (I357072,I3570);
DFFARX1 I_20793 (I787319,I3563,I357072,I357098,);
nand I_20794 (I357106,I787310,I787325);
and I_20795 (I357123,I357106,I787331);
DFFARX1 I_20796 (I357123,I3563,I357072,I357149,);
nor I_20797 (I357040,I357149,I357098);
not I_20798 (I357171,I357149);
DFFARX1 I_20799 (I787316,I3563,I357072,I357197,);
nand I_20800 (I357205,I357197,I787310);
not I_20801 (I357222,I357205);
DFFARX1 I_20802 (I357222,I3563,I357072,I357248,);
not I_20803 (I357064,I357248);
nor I_20804 (I357270,I357098,I357205);
nor I_20805 (I357046,I357149,I357270);
DFFARX1 I_20806 (I787313,I3563,I357072,I357310,);
DFFARX1 I_20807 (I357310,I3563,I357072,I357327,);
not I_20808 (I357335,I357327);
not I_20809 (I357352,I357310);
nand I_20810 (I357049,I357352,I357171);
nand I_20811 (I357383,I787307,I787322);
and I_20812 (I357400,I357383,I787307);
DFFARX1 I_20813 (I357400,I3563,I357072,I357426,);
nor I_20814 (I357434,I357426,I357098);
DFFARX1 I_20815 (I357434,I3563,I357072,I357037,);
DFFARX1 I_20816 (I357426,I3563,I357072,I357055,);
nor I_20817 (I357479,I787328,I787322);
not I_20818 (I357496,I357479);
nor I_20819 (I357058,I357335,I357496);
nand I_20820 (I357043,I357352,I357496);
nor I_20821 (I357052,I357098,I357479);
DFFARX1 I_20822 (I357479,I3563,I357072,I357061,);
not I_20823 (I357599,I3570);
DFFARX1 I_20824 (I1137813,I3563,I357599,I357625,);
nand I_20825 (I357633,I1137828,I1137813);
and I_20826 (I357650,I357633,I1137831);
DFFARX1 I_20827 (I357650,I3563,I357599,I357676,);
nor I_20828 (I357567,I357676,I357625);
not I_20829 (I357698,I357676);
DFFARX1 I_20830 (I1137837,I3563,I357599,I357724,);
nand I_20831 (I357732,I357724,I1137819);
not I_20832 (I357749,I357732);
DFFARX1 I_20833 (I357749,I3563,I357599,I357775,);
not I_20834 (I357591,I357775);
nor I_20835 (I357797,I357625,I357732);
nor I_20836 (I357573,I357676,I357797);
DFFARX1 I_20837 (I1137816,I3563,I357599,I357837,);
DFFARX1 I_20838 (I357837,I3563,I357599,I357854,);
not I_20839 (I357862,I357854);
not I_20840 (I357879,I357837);
nand I_20841 (I357576,I357879,I357698);
nand I_20842 (I357910,I1137816,I1137822);
and I_20843 (I357927,I357910,I1137834);
DFFARX1 I_20844 (I357927,I3563,I357599,I357953,);
nor I_20845 (I357961,I357953,I357625);
DFFARX1 I_20846 (I357961,I3563,I357599,I357564,);
DFFARX1 I_20847 (I357953,I3563,I357599,I357582,);
nor I_20848 (I358006,I1137825,I1137822);
not I_20849 (I358023,I358006);
nor I_20850 (I357585,I357862,I358023);
nand I_20851 (I357570,I357879,I358023);
nor I_20852 (I357579,I357625,I358006);
DFFARX1 I_20853 (I358006,I3563,I357599,I357588,);
not I_20854 (I358126,I3570);
DFFARX1 I_20855 (I1135501,I3563,I358126,I358152,);
nand I_20856 (I358160,I1135516,I1135501);
and I_20857 (I358177,I358160,I1135519);
DFFARX1 I_20858 (I358177,I3563,I358126,I358203,);
nor I_20859 (I358094,I358203,I358152);
not I_20860 (I358225,I358203);
DFFARX1 I_20861 (I1135525,I3563,I358126,I358251,);
nand I_20862 (I358259,I358251,I1135507);
not I_20863 (I358276,I358259);
DFFARX1 I_20864 (I358276,I3563,I358126,I358302,);
not I_20865 (I358118,I358302);
nor I_20866 (I358324,I358152,I358259);
nor I_20867 (I358100,I358203,I358324);
DFFARX1 I_20868 (I1135504,I3563,I358126,I358364,);
DFFARX1 I_20869 (I358364,I3563,I358126,I358381,);
not I_20870 (I358389,I358381);
not I_20871 (I358406,I358364);
nand I_20872 (I358103,I358406,I358225);
nand I_20873 (I358437,I1135504,I1135510);
and I_20874 (I358454,I358437,I1135522);
DFFARX1 I_20875 (I358454,I3563,I358126,I358480,);
nor I_20876 (I358488,I358480,I358152);
DFFARX1 I_20877 (I358488,I3563,I358126,I358091,);
DFFARX1 I_20878 (I358480,I3563,I358126,I358109,);
nor I_20879 (I358533,I1135513,I1135510);
not I_20880 (I358550,I358533);
nor I_20881 (I358112,I358389,I358550);
nand I_20882 (I358097,I358406,I358550);
nor I_20883 (I358106,I358152,I358533);
DFFARX1 I_20884 (I358533,I3563,I358126,I358115,);
not I_20885 (I358653,I3570);
DFFARX1 I_20886 (I15488,I3563,I358653,I358679,);
nand I_20887 (I358687,I15479,I15482);
and I_20888 (I358704,I358687,I15473);
DFFARX1 I_20889 (I358704,I3563,I358653,I358730,);
nor I_20890 (I358621,I358730,I358679);
not I_20891 (I358752,I358730);
DFFARX1 I_20892 (I15479,I3563,I358653,I358778,);
nand I_20893 (I358786,I358778,I15485);
not I_20894 (I358803,I358786);
DFFARX1 I_20895 (I358803,I3563,I358653,I358829,);
not I_20896 (I358645,I358829);
nor I_20897 (I358851,I358679,I358786);
nor I_20898 (I358627,I358730,I358851);
DFFARX1 I_20899 (I15476,I3563,I358653,I358891,);
DFFARX1 I_20900 (I358891,I3563,I358653,I358908,);
not I_20901 (I358916,I358908);
not I_20902 (I358933,I358891);
nand I_20903 (I358630,I358933,I358752);
nand I_20904 (I358964,I15476,I15491);
and I_20905 (I358981,I358964,I15473);
DFFARX1 I_20906 (I358981,I3563,I358653,I359007,);
nor I_20907 (I359015,I359007,I358679);
DFFARX1 I_20908 (I359015,I3563,I358653,I358618,);
DFFARX1 I_20909 (I359007,I3563,I358653,I358636,);
nor I_20910 (I359060,I15494,I15491);
not I_20911 (I359077,I359060);
nor I_20912 (I358639,I358916,I359077);
nand I_20913 (I358624,I358933,I359077);
nor I_20914 (I358633,I358679,I359060);
DFFARX1 I_20915 (I359060,I3563,I358653,I358642,);
not I_20916 (I359180,I3570);
DFFARX1 I_20917 (I543564,I3563,I359180,I359206,);
nand I_20918 (I359214,I543564,I543576);
and I_20919 (I359231,I359214,I543561);
DFFARX1 I_20920 (I359231,I3563,I359180,I359257,);
nor I_20921 (I359148,I359257,I359206);
not I_20922 (I359279,I359257);
DFFARX1 I_20923 (I543585,I3563,I359180,I359305,);
nand I_20924 (I359313,I359305,I543582);
not I_20925 (I359330,I359313);
DFFARX1 I_20926 (I359330,I3563,I359180,I359356,);
not I_20927 (I359172,I359356);
nor I_20928 (I359378,I359206,I359313);
nor I_20929 (I359154,I359257,I359378);
DFFARX1 I_20930 (I543573,I3563,I359180,I359418,);
DFFARX1 I_20931 (I359418,I3563,I359180,I359435,);
not I_20932 (I359443,I359435);
not I_20933 (I359460,I359418);
nand I_20934 (I359157,I359460,I359279);
nand I_20935 (I359491,I543561,I543570);
and I_20936 (I359508,I359491,I543579);
DFFARX1 I_20937 (I359508,I3563,I359180,I359534,);
nor I_20938 (I359542,I359534,I359206);
DFFARX1 I_20939 (I359542,I3563,I359180,I359145,);
DFFARX1 I_20940 (I359534,I3563,I359180,I359163,);
nor I_20941 (I359587,I543567,I543570);
not I_20942 (I359604,I359587);
nor I_20943 (I359166,I359443,I359604);
nand I_20944 (I359151,I359460,I359604);
nor I_20945 (I359160,I359206,I359587);
DFFARX1 I_20946 (I359587,I3563,I359180,I359169,);
not I_20947 (I359707,I3570);
DFFARX1 I_20948 (I868502,I3563,I359707,I359733,);
nand I_20949 (I359741,I868505,I868499);
and I_20950 (I359758,I359741,I868511);
DFFARX1 I_20951 (I359758,I3563,I359707,I359784,);
nor I_20952 (I359675,I359784,I359733);
not I_20953 (I359806,I359784);
DFFARX1 I_20954 (I868514,I3563,I359707,I359832,);
nand I_20955 (I359840,I359832,I868505);
not I_20956 (I359857,I359840);
DFFARX1 I_20957 (I359857,I3563,I359707,I359883,);
not I_20958 (I359699,I359883);
nor I_20959 (I359905,I359733,I359840);
nor I_20960 (I359681,I359784,I359905);
DFFARX1 I_20961 (I868517,I3563,I359707,I359945,);
DFFARX1 I_20962 (I359945,I3563,I359707,I359962,);
not I_20963 (I359970,I359962);
not I_20964 (I359987,I359945);
nand I_20965 (I359684,I359987,I359806);
nand I_20966 (I360018,I868499,I868508);
and I_20967 (I360035,I360018,I868502);
DFFARX1 I_20968 (I360035,I3563,I359707,I360061,);
nor I_20969 (I360069,I360061,I359733);
DFFARX1 I_20970 (I360069,I3563,I359707,I359672,);
DFFARX1 I_20971 (I360061,I3563,I359707,I359690,);
nor I_20972 (I360114,I868520,I868508);
not I_20973 (I360131,I360114);
nor I_20974 (I359693,I359970,I360131);
nand I_20975 (I359678,I359987,I360131);
nor I_20976 (I359687,I359733,I360114);
DFFARX1 I_20977 (I360114,I3563,I359707,I359696,);
not I_20978 (I360234,I3570);
DFFARX1 I_20979 (I1404139,I3563,I360234,I360260,);
nand I_20980 (I360268,I1404118,I1404118);
and I_20981 (I360285,I360268,I1404145);
DFFARX1 I_20982 (I360285,I3563,I360234,I360311,);
nor I_20983 (I360202,I360311,I360260);
not I_20984 (I360333,I360311);
DFFARX1 I_20985 (I1404133,I3563,I360234,I360359,);
nand I_20986 (I360367,I360359,I1404136);
not I_20987 (I360384,I360367);
DFFARX1 I_20988 (I360384,I3563,I360234,I360410,);
not I_20989 (I360226,I360410);
nor I_20990 (I360432,I360260,I360367);
nor I_20991 (I360208,I360311,I360432);
DFFARX1 I_20992 (I1404127,I3563,I360234,I360472,);
DFFARX1 I_20993 (I360472,I3563,I360234,I360489,);
not I_20994 (I360497,I360489);
not I_20995 (I360514,I360472);
nand I_20996 (I360211,I360514,I360333);
nand I_20997 (I360545,I1404124,I1404121);
and I_20998 (I360562,I360545,I1404142);
DFFARX1 I_20999 (I360562,I3563,I360234,I360588,);
nor I_21000 (I360596,I360588,I360260);
DFFARX1 I_21001 (I360596,I3563,I360234,I360199,);
DFFARX1 I_21002 (I360588,I3563,I360234,I360217,);
nor I_21003 (I360641,I1404130,I1404121);
not I_21004 (I360658,I360641);
nor I_21005 (I360220,I360497,I360658);
nand I_21006 (I360205,I360514,I360658);
nor I_21007 (I360214,I360260,I360641);
DFFARX1 I_21008 (I360641,I3563,I360234,I360223,);
not I_21009 (I360761,I3570);
DFFARX1 I_21010 (I967850,I3563,I360761,I360787,);
nand I_21011 (I360795,I967847,I967865);
and I_21012 (I360812,I360795,I967856);
DFFARX1 I_21013 (I360812,I3563,I360761,I360838,);
nor I_21014 (I360729,I360838,I360787);
not I_21015 (I360860,I360838);
DFFARX1 I_21016 (I967871,I3563,I360761,I360886,);
nand I_21017 (I360894,I360886,I967853);
not I_21018 (I360911,I360894);
DFFARX1 I_21019 (I360911,I3563,I360761,I360937,);
not I_21020 (I360753,I360937);
nor I_21021 (I360959,I360787,I360894);
nor I_21022 (I360735,I360838,I360959);
DFFARX1 I_21023 (I967859,I3563,I360761,I360999,);
DFFARX1 I_21024 (I360999,I3563,I360761,I361016,);
not I_21025 (I361024,I361016);
not I_21026 (I361041,I360999);
nand I_21027 (I360738,I361041,I360860);
nand I_21028 (I361072,I967847,I967874);
and I_21029 (I361089,I361072,I967862);
DFFARX1 I_21030 (I361089,I3563,I360761,I361115,);
nor I_21031 (I361123,I361115,I360787);
DFFARX1 I_21032 (I361123,I3563,I360761,I360726,);
DFFARX1 I_21033 (I361115,I3563,I360761,I360744,);
nor I_21034 (I361168,I967868,I967874);
not I_21035 (I361185,I361168);
nor I_21036 (I360747,I361024,I361185);
nand I_21037 (I360732,I361041,I361185);
nor I_21038 (I360741,I360787,I361168);
DFFARX1 I_21039 (I361168,I3563,I360761,I360750,);
not I_21040 (I361288,I3570);
DFFARX1 I_21041 (I1080322,I3563,I361288,I361314,);
nand I_21042 (I361322,I1080319,I1080322);
and I_21043 (I361339,I361322,I1080331);
DFFARX1 I_21044 (I361339,I3563,I361288,I361365,);
nor I_21045 (I361256,I361365,I361314);
not I_21046 (I361387,I361365);
DFFARX1 I_21047 (I1080319,I3563,I361288,I361413,);
nand I_21048 (I361421,I361413,I1080337);
not I_21049 (I361438,I361421);
DFFARX1 I_21050 (I361438,I3563,I361288,I361464,);
not I_21051 (I361280,I361464);
nor I_21052 (I361486,I361314,I361421);
nor I_21053 (I361262,I361365,I361486);
DFFARX1 I_21054 (I1080325,I3563,I361288,I361526,);
DFFARX1 I_21055 (I361526,I3563,I361288,I361543,);
not I_21056 (I361551,I361543);
not I_21057 (I361568,I361526);
nand I_21058 (I361265,I361568,I361387);
nand I_21059 (I361599,I1080334,I1080340);
and I_21060 (I361616,I361599,I1080325);
DFFARX1 I_21061 (I361616,I3563,I361288,I361642,);
nor I_21062 (I361650,I361642,I361314);
DFFARX1 I_21063 (I361650,I3563,I361288,I361253,);
DFFARX1 I_21064 (I361642,I3563,I361288,I361271,);
nor I_21065 (I361695,I1080328,I1080340);
not I_21066 (I361712,I361695);
nor I_21067 (I361274,I361551,I361712);
nand I_21068 (I361259,I361568,I361712);
nor I_21069 (I361268,I361314,I361695);
DFFARX1 I_21070 (I361695,I3563,I361288,I361277,);
not I_21071 (I361815,I3570);
DFFARX1 I_21072 (I956222,I3563,I361815,I361841,);
nand I_21073 (I361849,I956219,I956237);
and I_21074 (I361866,I361849,I956228);
DFFARX1 I_21075 (I361866,I3563,I361815,I361892,);
nor I_21076 (I361783,I361892,I361841);
not I_21077 (I361914,I361892);
DFFARX1 I_21078 (I956243,I3563,I361815,I361940,);
nand I_21079 (I361948,I361940,I956225);
not I_21080 (I361965,I361948);
DFFARX1 I_21081 (I361965,I3563,I361815,I361991,);
not I_21082 (I361807,I361991);
nor I_21083 (I362013,I361841,I361948);
nor I_21084 (I361789,I361892,I362013);
DFFARX1 I_21085 (I956231,I3563,I361815,I362053,);
DFFARX1 I_21086 (I362053,I3563,I361815,I362070,);
not I_21087 (I362078,I362070);
not I_21088 (I362095,I362053);
nand I_21089 (I361792,I362095,I361914);
nand I_21090 (I362126,I956219,I956246);
and I_21091 (I362143,I362126,I956234);
DFFARX1 I_21092 (I362143,I3563,I361815,I362169,);
nor I_21093 (I362177,I362169,I361841);
DFFARX1 I_21094 (I362177,I3563,I361815,I361780,);
DFFARX1 I_21095 (I362169,I3563,I361815,I361798,);
nor I_21096 (I362222,I956240,I956246);
not I_21097 (I362239,I362222);
nor I_21098 (I361801,I362078,I362239);
nand I_21099 (I361786,I362095,I362239);
nor I_21100 (I361795,I361841,I362222);
DFFARX1 I_21101 (I362222,I3563,I361815,I361804,);
not I_21102 (I362342,I3570);
DFFARX1 I_21103 (I115674,I3563,I362342,I362368,);
nand I_21104 (I362376,I115686,I115695);
and I_21105 (I362393,I362376,I115674);
DFFARX1 I_21106 (I362393,I3563,I362342,I362419,);
nor I_21107 (I362310,I362419,I362368);
not I_21108 (I362441,I362419);
DFFARX1 I_21109 (I115689,I3563,I362342,I362467,);
nand I_21110 (I362475,I362467,I115677);
not I_21111 (I362492,I362475);
DFFARX1 I_21112 (I362492,I3563,I362342,I362518,);
not I_21113 (I362334,I362518);
nor I_21114 (I362540,I362368,I362475);
nor I_21115 (I362316,I362419,I362540);
DFFARX1 I_21116 (I115680,I3563,I362342,I362580,);
DFFARX1 I_21117 (I362580,I3563,I362342,I362597,);
not I_21118 (I362605,I362597);
not I_21119 (I362622,I362580);
nand I_21120 (I362319,I362622,I362441);
nand I_21121 (I362653,I115671,I115671);
and I_21122 (I362670,I362653,I115683);
DFFARX1 I_21123 (I362670,I3563,I362342,I362696,);
nor I_21124 (I362704,I362696,I362368);
DFFARX1 I_21125 (I362704,I3563,I362342,I362307,);
DFFARX1 I_21126 (I362696,I3563,I362342,I362325,);
nor I_21127 (I362749,I115692,I115671);
not I_21128 (I362766,I362749);
nor I_21129 (I362328,I362605,I362766);
nand I_21130 (I362313,I362622,I362766);
nor I_21131 (I362322,I362368,I362749);
DFFARX1 I_21132 (I362749,I3563,I362342,I362331,);
not I_21133 (I362869,I3570);
DFFARX1 I_21134 (I139916,I3563,I362869,I362895,);
nand I_21135 (I362903,I139928,I139937);
and I_21136 (I362920,I362903,I139916);
DFFARX1 I_21137 (I362920,I3563,I362869,I362946,);
nor I_21138 (I362837,I362946,I362895);
not I_21139 (I362968,I362946);
DFFARX1 I_21140 (I139931,I3563,I362869,I362994,);
nand I_21141 (I363002,I362994,I139919);
not I_21142 (I363019,I363002);
DFFARX1 I_21143 (I363019,I3563,I362869,I363045,);
not I_21144 (I362861,I363045);
nor I_21145 (I363067,I362895,I363002);
nor I_21146 (I362843,I362946,I363067);
DFFARX1 I_21147 (I139922,I3563,I362869,I363107,);
DFFARX1 I_21148 (I363107,I3563,I362869,I363124,);
not I_21149 (I363132,I363124);
not I_21150 (I363149,I363107);
nand I_21151 (I362846,I363149,I362968);
nand I_21152 (I363180,I139913,I139913);
and I_21153 (I363197,I363180,I139925);
DFFARX1 I_21154 (I363197,I3563,I362869,I363223,);
nor I_21155 (I363231,I363223,I362895);
DFFARX1 I_21156 (I363231,I3563,I362869,I362834,);
DFFARX1 I_21157 (I363223,I3563,I362869,I362852,);
nor I_21158 (I363276,I139934,I139913);
not I_21159 (I363293,I363276);
nor I_21160 (I362855,I363132,I363293);
nand I_21161 (I362840,I363149,I363293);
nor I_21162 (I362849,I362895,I363276);
DFFARX1 I_21163 (I363276,I3563,I362869,I362858,);
not I_21164 (I363396,I3570);
DFFARX1 I_21165 (I1124519,I3563,I363396,I363422,);
nand I_21166 (I363430,I1124534,I1124519);
and I_21167 (I363447,I363430,I1124537);
DFFARX1 I_21168 (I363447,I3563,I363396,I363473,);
nor I_21169 (I363364,I363473,I363422);
not I_21170 (I363495,I363473);
DFFARX1 I_21171 (I1124543,I3563,I363396,I363521,);
nand I_21172 (I363529,I363521,I1124525);
not I_21173 (I363546,I363529);
DFFARX1 I_21174 (I363546,I3563,I363396,I363572,);
not I_21175 (I363388,I363572);
nor I_21176 (I363594,I363422,I363529);
nor I_21177 (I363370,I363473,I363594);
DFFARX1 I_21178 (I1124522,I3563,I363396,I363634,);
DFFARX1 I_21179 (I363634,I3563,I363396,I363651,);
not I_21180 (I363659,I363651);
not I_21181 (I363676,I363634);
nand I_21182 (I363373,I363676,I363495);
nand I_21183 (I363707,I1124522,I1124528);
and I_21184 (I363724,I363707,I1124540);
DFFARX1 I_21185 (I363724,I3563,I363396,I363750,);
nor I_21186 (I363758,I363750,I363422);
DFFARX1 I_21187 (I363758,I3563,I363396,I363361,);
DFFARX1 I_21188 (I363750,I3563,I363396,I363379,);
nor I_21189 (I363803,I1124531,I1124528);
not I_21190 (I363820,I363803);
nor I_21191 (I363382,I363659,I363820);
nand I_21192 (I363367,I363676,I363820);
nor I_21193 (I363376,I363422,I363803);
DFFARX1 I_21194 (I363803,I3563,I363396,I363385,);
not I_21195 (I363923,I3570);
DFFARX1 I_21196 (I757841,I3563,I363923,I363949,);
nand I_21197 (I363957,I757832,I757847);
and I_21198 (I363974,I363957,I757853);
DFFARX1 I_21199 (I363974,I3563,I363923,I364000,);
nor I_21200 (I363891,I364000,I363949);
not I_21201 (I364022,I364000);
DFFARX1 I_21202 (I757838,I3563,I363923,I364048,);
nand I_21203 (I364056,I364048,I757832);
not I_21204 (I364073,I364056);
DFFARX1 I_21205 (I364073,I3563,I363923,I364099,);
not I_21206 (I363915,I364099);
nor I_21207 (I364121,I363949,I364056);
nor I_21208 (I363897,I364000,I364121);
DFFARX1 I_21209 (I757835,I3563,I363923,I364161,);
DFFARX1 I_21210 (I364161,I3563,I363923,I364178,);
not I_21211 (I364186,I364178);
not I_21212 (I364203,I364161);
nand I_21213 (I363900,I364203,I364022);
nand I_21214 (I364234,I757829,I757844);
and I_21215 (I364251,I364234,I757829);
DFFARX1 I_21216 (I364251,I3563,I363923,I364277,);
nor I_21217 (I364285,I364277,I363949);
DFFARX1 I_21218 (I364285,I3563,I363923,I363888,);
DFFARX1 I_21219 (I364277,I3563,I363923,I363906,);
nor I_21220 (I364330,I757850,I757844);
not I_21221 (I364347,I364330);
nor I_21222 (I363909,I364186,I364347);
nand I_21223 (I363894,I364203,I364347);
nor I_21224 (I363903,I363949,I364330);
DFFARX1 I_21225 (I364330,I3563,I363923,I363912,);
not I_21226 (I364450,I3570);
DFFARX1 I_21227 (I981416,I3563,I364450,I364476,);
nand I_21228 (I364484,I981413,I981431);
and I_21229 (I364501,I364484,I981422);
DFFARX1 I_21230 (I364501,I3563,I364450,I364527,);
nor I_21231 (I364418,I364527,I364476);
not I_21232 (I364549,I364527);
DFFARX1 I_21233 (I981437,I3563,I364450,I364575,);
nand I_21234 (I364583,I364575,I981419);
not I_21235 (I364600,I364583);
DFFARX1 I_21236 (I364600,I3563,I364450,I364626,);
not I_21237 (I364442,I364626);
nor I_21238 (I364648,I364476,I364583);
nor I_21239 (I364424,I364527,I364648);
DFFARX1 I_21240 (I981425,I3563,I364450,I364688,);
DFFARX1 I_21241 (I364688,I3563,I364450,I364705,);
not I_21242 (I364713,I364705);
not I_21243 (I364730,I364688);
nand I_21244 (I364427,I364730,I364549);
nand I_21245 (I364761,I981413,I981440);
and I_21246 (I364778,I364761,I981428);
DFFARX1 I_21247 (I364778,I3563,I364450,I364804,);
nor I_21248 (I364812,I364804,I364476);
DFFARX1 I_21249 (I364812,I3563,I364450,I364415,);
DFFARX1 I_21250 (I364804,I3563,I364450,I364433,);
nor I_21251 (I364857,I981434,I981440);
not I_21252 (I364874,I364857);
nor I_21253 (I364436,I364713,I364874);
nand I_21254 (I364421,I364730,I364874);
nor I_21255 (I364430,I364476,I364857);
DFFARX1 I_21256 (I364857,I3563,I364450,I364439,);
not I_21257 (I364977,I3570);
DFFARX1 I_21258 (I945240,I3563,I364977,I365003,);
nand I_21259 (I365011,I945237,I945255);
and I_21260 (I365028,I365011,I945246);
DFFARX1 I_21261 (I365028,I3563,I364977,I365054,);
nor I_21262 (I364945,I365054,I365003);
not I_21263 (I365076,I365054);
DFFARX1 I_21264 (I945261,I3563,I364977,I365102,);
nand I_21265 (I365110,I365102,I945243);
not I_21266 (I365127,I365110);
DFFARX1 I_21267 (I365127,I3563,I364977,I365153,);
not I_21268 (I364969,I365153);
nor I_21269 (I365175,I365003,I365110);
nor I_21270 (I364951,I365054,I365175);
DFFARX1 I_21271 (I945249,I3563,I364977,I365215,);
DFFARX1 I_21272 (I365215,I3563,I364977,I365232,);
not I_21273 (I365240,I365232);
not I_21274 (I365257,I365215);
nand I_21275 (I364954,I365257,I365076);
nand I_21276 (I365288,I945237,I945264);
and I_21277 (I365305,I365288,I945252);
DFFARX1 I_21278 (I365305,I3563,I364977,I365331,);
nor I_21279 (I365339,I365331,I365003);
DFFARX1 I_21280 (I365339,I3563,I364977,I364942,);
DFFARX1 I_21281 (I365331,I3563,I364977,I364960,);
nor I_21282 (I365384,I945258,I945264);
not I_21283 (I365401,I365384);
nor I_21284 (I364963,I365240,I365401);
nand I_21285 (I364948,I365257,I365401);
nor I_21286 (I364957,I365003,I365384);
DFFARX1 I_21287 (I365384,I3563,I364977,I364966,);
not I_21288 (I365504,I3570);
DFFARX1 I_21289 (I37148,I3563,I365504,I365530,);
nand I_21290 (I365538,I37172,I37151);
and I_21291 (I365555,I365538,I37148);
DFFARX1 I_21292 (I365555,I3563,I365504,I365581,);
nor I_21293 (I365472,I365581,I365530);
not I_21294 (I365603,I365581);
DFFARX1 I_21295 (I37154,I3563,I365504,I365629,);
nand I_21296 (I365637,I365629,I37163);
not I_21297 (I365654,I365637);
DFFARX1 I_21298 (I365654,I3563,I365504,I365680,);
not I_21299 (I365496,I365680);
nor I_21300 (I365702,I365530,I365637);
nor I_21301 (I365478,I365581,I365702);
DFFARX1 I_21302 (I37157,I3563,I365504,I365742,);
DFFARX1 I_21303 (I365742,I3563,I365504,I365759,);
not I_21304 (I365767,I365759);
not I_21305 (I365784,I365742);
nand I_21306 (I365481,I365784,I365603);
nand I_21307 (I365815,I37169,I37151);
and I_21308 (I365832,I365815,I37160);
DFFARX1 I_21309 (I365832,I3563,I365504,I365858,);
nor I_21310 (I365866,I365858,I365530);
DFFARX1 I_21311 (I365866,I3563,I365504,I365469,);
DFFARX1 I_21312 (I365858,I3563,I365504,I365487,);
nor I_21313 (I365911,I37166,I37151);
not I_21314 (I365928,I365911);
nor I_21315 (I365490,I365767,I365928);
nand I_21316 (I365475,I365784,I365928);
nor I_21317 (I365484,I365530,I365911);
DFFARX1 I_21318 (I365911,I3563,I365504,I365493,);
not I_21319 (I366031,I3570);
DFFARX1 I_21320 (I1199659,I3563,I366031,I366057,);
nand I_21321 (I366065,I1199674,I1199659);
and I_21322 (I366082,I366065,I1199677);
DFFARX1 I_21323 (I366082,I3563,I366031,I366108,);
nor I_21324 (I365999,I366108,I366057);
not I_21325 (I366130,I366108);
DFFARX1 I_21326 (I1199683,I3563,I366031,I366156,);
nand I_21327 (I366164,I366156,I1199665);
not I_21328 (I366181,I366164);
DFFARX1 I_21329 (I366181,I3563,I366031,I366207,);
not I_21330 (I366023,I366207);
nor I_21331 (I366229,I366057,I366164);
nor I_21332 (I366005,I366108,I366229);
DFFARX1 I_21333 (I1199662,I3563,I366031,I366269,);
DFFARX1 I_21334 (I366269,I3563,I366031,I366286,);
not I_21335 (I366294,I366286);
not I_21336 (I366311,I366269);
nand I_21337 (I366008,I366311,I366130);
nand I_21338 (I366342,I1199662,I1199668);
and I_21339 (I366359,I366342,I1199680);
DFFARX1 I_21340 (I366359,I3563,I366031,I366385,);
nor I_21341 (I366393,I366385,I366057);
DFFARX1 I_21342 (I366393,I3563,I366031,I365996,);
DFFARX1 I_21343 (I366385,I3563,I366031,I366014,);
nor I_21344 (I366438,I1199671,I1199668);
not I_21345 (I366455,I366438);
nor I_21346 (I366017,I366294,I366455);
nand I_21347 (I366002,I366311,I366455);
nor I_21348 (I366011,I366057,I366438);
DFFARX1 I_21349 (I366438,I3563,I366031,I366020,);
not I_21350 (I366558,I3570);
DFFARX1 I_21351 (I1210641,I3563,I366558,I366584,);
nand I_21352 (I366592,I1210656,I1210641);
and I_21353 (I366609,I366592,I1210659);
DFFARX1 I_21354 (I366609,I3563,I366558,I366635,);
nor I_21355 (I366526,I366635,I366584);
not I_21356 (I366657,I366635);
DFFARX1 I_21357 (I1210665,I3563,I366558,I366683,);
nand I_21358 (I366691,I366683,I1210647);
not I_21359 (I366708,I366691);
DFFARX1 I_21360 (I366708,I3563,I366558,I366734,);
not I_21361 (I366550,I366734);
nor I_21362 (I366756,I366584,I366691);
nor I_21363 (I366532,I366635,I366756);
DFFARX1 I_21364 (I1210644,I3563,I366558,I366796,);
DFFARX1 I_21365 (I366796,I3563,I366558,I366813,);
not I_21366 (I366821,I366813);
not I_21367 (I366838,I366796);
nand I_21368 (I366535,I366838,I366657);
nand I_21369 (I366869,I1210644,I1210650);
and I_21370 (I366886,I366869,I1210662);
DFFARX1 I_21371 (I366886,I3563,I366558,I366912,);
nor I_21372 (I366920,I366912,I366584);
DFFARX1 I_21373 (I366920,I3563,I366558,I366523,);
DFFARX1 I_21374 (I366912,I3563,I366558,I366541,);
nor I_21375 (I366965,I1210653,I1210650);
not I_21376 (I366982,I366965);
nor I_21377 (I366544,I366821,I366982);
nand I_21378 (I366529,I366838,I366982);
nor I_21379 (I366538,I366584,I366965);
DFFARX1 I_21380 (I366965,I3563,I366558,I366547,);
not I_21381 (I367085,I3570);
DFFARX1 I_21382 (I1282331,I3563,I367085,I367111,);
nand I_21383 (I367119,I1282313,I1282337);
and I_21384 (I367136,I367119,I1282328);
DFFARX1 I_21385 (I367136,I3563,I367085,I367162,);
nor I_21386 (I367053,I367162,I367111);
not I_21387 (I367184,I367162);
DFFARX1 I_21388 (I1282334,I3563,I367085,I367210,);
nand I_21389 (I367218,I367210,I1282322);
not I_21390 (I367235,I367218);
DFFARX1 I_21391 (I367235,I3563,I367085,I367261,);
not I_21392 (I367077,I367261);
nor I_21393 (I367283,I367111,I367218);
nor I_21394 (I367059,I367162,I367283);
DFFARX1 I_21395 (I1282313,I3563,I367085,I367323,);
DFFARX1 I_21396 (I367323,I3563,I367085,I367340,);
not I_21397 (I367348,I367340);
not I_21398 (I367365,I367323);
nand I_21399 (I367062,I367365,I367184);
nand I_21400 (I367396,I1282319,I1282316);
and I_21401 (I367413,I367396,I1282325);
DFFARX1 I_21402 (I367413,I3563,I367085,I367439,);
nor I_21403 (I367447,I367439,I367111);
DFFARX1 I_21404 (I367447,I3563,I367085,I367050,);
DFFARX1 I_21405 (I367439,I3563,I367085,I367068,);
nor I_21406 (I367492,I1282316,I1282316);
not I_21407 (I367509,I367492);
nor I_21408 (I367071,I367348,I367509);
nand I_21409 (I367056,I367365,I367509);
nor I_21410 (I367065,I367111,I367492);
DFFARX1 I_21411 (I367492,I3563,I367085,I367074,);
not I_21412 (I367612,I3570);
DFFARX1 I_21413 (I679811,I3563,I367612,I367638,);
nand I_21414 (I367646,I679802,I679817);
and I_21415 (I367663,I367646,I679823);
DFFARX1 I_21416 (I367663,I3563,I367612,I367689,);
nor I_21417 (I367580,I367689,I367638);
not I_21418 (I367711,I367689);
DFFARX1 I_21419 (I679808,I3563,I367612,I367737,);
nand I_21420 (I367745,I367737,I679802);
not I_21421 (I367762,I367745);
DFFARX1 I_21422 (I367762,I3563,I367612,I367788,);
not I_21423 (I367604,I367788);
nor I_21424 (I367810,I367638,I367745);
nor I_21425 (I367586,I367689,I367810);
DFFARX1 I_21426 (I679805,I3563,I367612,I367850,);
DFFARX1 I_21427 (I367850,I3563,I367612,I367867,);
not I_21428 (I367875,I367867);
not I_21429 (I367892,I367850);
nand I_21430 (I367589,I367892,I367711);
nand I_21431 (I367923,I679799,I679814);
and I_21432 (I367940,I367923,I679799);
DFFARX1 I_21433 (I367940,I3563,I367612,I367966,);
nor I_21434 (I367974,I367966,I367638);
DFFARX1 I_21435 (I367974,I3563,I367612,I367577,);
DFFARX1 I_21436 (I367966,I3563,I367612,I367595,);
nor I_21437 (I368019,I679820,I679814);
not I_21438 (I368036,I368019);
nor I_21439 (I367598,I367875,I368036);
nand I_21440 (I367583,I367892,I368036);
nor I_21441 (I367592,I367638,I368019);
DFFARX1 I_21442 (I368019,I3563,I367612,I367601,);
not I_21443 (I368139,I3570);
DFFARX1 I_21444 (I600050,I3563,I368139,I368165,);
nand I_21445 (I368173,I600035,I600038);
and I_21446 (I368190,I368173,I600053);
DFFARX1 I_21447 (I368190,I3563,I368139,I368216,);
nor I_21448 (I368107,I368216,I368165);
not I_21449 (I368238,I368216);
DFFARX1 I_21450 (I600047,I3563,I368139,I368264,);
nand I_21451 (I368272,I368264,I600038);
not I_21452 (I368289,I368272);
DFFARX1 I_21453 (I368289,I3563,I368139,I368315,);
not I_21454 (I368131,I368315);
nor I_21455 (I368337,I368165,I368272);
nor I_21456 (I368113,I368216,I368337);
DFFARX1 I_21457 (I600044,I3563,I368139,I368377,);
DFFARX1 I_21458 (I368377,I3563,I368139,I368394,);
not I_21459 (I368402,I368394);
not I_21460 (I368419,I368377);
nand I_21461 (I368116,I368419,I368238);
nand I_21462 (I368450,I600059,I600035);
and I_21463 (I368467,I368450,I600056);
DFFARX1 I_21464 (I368467,I3563,I368139,I368493,);
nor I_21465 (I368501,I368493,I368165);
DFFARX1 I_21466 (I368501,I3563,I368139,I368104,);
DFFARX1 I_21467 (I368493,I3563,I368139,I368122,);
nor I_21468 (I368546,I600041,I600035);
not I_21469 (I368563,I368546);
nor I_21470 (I368125,I368402,I368563);
nand I_21471 (I368110,I368419,I368563);
nor I_21472 (I368119,I368165,I368546);
DFFARX1 I_21473 (I368546,I3563,I368139,I368128,);
not I_21474 (I368666,I3570);
DFFARX1 I_21475 (I1170759,I3563,I368666,I368692,);
nand I_21476 (I368700,I1170774,I1170759);
and I_21477 (I368717,I368700,I1170777);
DFFARX1 I_21478 (I368717,I3563,I368666,I368743,);
nor I_21479 (I368634,I368743,I368692);
not I_21480 (I368765,I368743);
DFFARX1 I_21481 (I1170783,I3563,I368666,I368791,);
nand I_21482 (I368799,I368791,I1170765);
not I_21483 (I368816,I368799);
DFFARX1 I_21484 (I368816,I3563,I368666,I368842,);
not I_21485 (I368658,I368842);
nor I_21486 (I368864,I368692,I368799);
nor I_21487 (I368640,I368743,I368864);
DFFARX1 I_21488 (I1170762,I3563,I368666,I368904,);
DFFARX1 I_21489 (I368904,I3563,I368666,I368921,);
not I_21490 (I368929,I368921);
not I_21491 (I368946,I368904);
nand I_21492 (I368643,I368946,I368765);
nand I_21493 (I368977,I1170762,I1170768);
and I_21494 (I368994,I368977,I1170780);
DFFARX1 I_21495 (I368994,I3563,I368666,I369020,);
nor I_21496 (I369028,I369020,I368692);
DFFARX1 I_21497 (I369028,I3563,I368666,I368631,);
DFFARX1 I_21498 (I369020,I3563,I368666,I368649,);
nor I_21499 (I369073,I1170771,I1170768);
not I_21500 (I369090,I369073);
nor I_21501 (I368652,I368929,I369090);
nand I_21502 (I368637,I368946,I369090);
nor I_21503 (I368646,I368692,I369073);
DFFARX1 I_21504 (I369073,I3563,I368666,I368655,);
not I_21505 (I369193,I3570);
DFFARX1 I_21506 (I1218733,I3563,I369193,I369219,);
nand I_21507 (I369227,I1218748,I1218733);
and I_21508 (I369244,I369227,I1218751);
DFFARX1 I_21509 (I369244,I3563,I369193,I369270,);
nor I_21510 (I369161,I369270,I369219);
not I_21511 (I369292,I369270);
DFFARX1 I_21512 (I1218757,I3563,I369193,I369318,);
nand I_21513 (I369326,I369318,I1218739);
not I_21514 (I369343,I369326);
DFFARX1 I_21515 (I369343,I3563,I369193,I369369,);
not I_21516 (I369185,I369369);
nor I_21517 (I369391,I369219,I369326);
nor I_21518 (I369167,I369270,I369391);
DFFARX1 I_21519 (I1218736,I3563,I369193,I369431,);
DFFARX1 I_21520 (I369431,I3563,I369193,I369448,);
not I_21521 (I369456,I369448);
not I_21522 (I369473,I369431);
nand I_21523 (I369170,I369473,I369292);
nand I_21524 (I369504,I1218736,I1218742);
and I_21525 (I369521,I369504,I1218754);
DFFARX1 I_21526 (I369521,I3563,I369193,I369547,);
nor I_21527 (I369555,I369547,I369219);
DFFARX1 I_21528 (I369555,I3563,I369193,I369158,);
DFFARX1 I_21529 (I369547,I3563,I369193,I369176,);
nor I_21530 (I369600,I1218745,I1218742);
not I_21531 (I369617,I369600);
nor I_21532 (I369179,I369456,I369617);
nand I_21533 (I369164,I369473,I369617);
nor I_21534 (I369173,I369219,I369600);
DFFARX1 I_21535 (I369600,I3563,I369193,I369182,);
not I_21536 (I369720,I3570);
DFFARX1 I_21537 (I713335,I3563,I369720,I369746,);
nand I_21538 (I369754,I713326,I713341);
and I_21539 (I369771,I369754,I713347);
DFFARX1 I_21540 (I369771,I3563,I369720,I369797,);
nor I_21541 (I369688,I369797,I369746);
not I_21542 (I369819,I369797);
DFFARX1 I_21543 (I713332,I3563,I369720,I369845,);
nand I_21544 (I369853,I369845,I713326);
not I_21545 (I369870,I369853);
DFFARX1 I_21546 (I369870,I3563,I369720,I369896,);
not I_21547 (I369712,I369896);
nor I_21548 (I369918,I369746,I369853);
nor I_21549 (I369694,I369797,I369918);
DFFARX1 I_21550 (I713329,I3563,I369720,I369958,);
DFFARX1 I_21551 (I369958,I3563,I369720,I369975,);
not I_21552 (I369983,I369975);
not I_21553 (I370000,I369958);
nand I_21554 (I369697,I370000,I369819);
nand I_21555 (I370031,I713323,I713338);
and I_21556 (I370048,I370031,I713323);
DFFARX1 I_21557 (I370048,I3563,I369720,I370074,);
nor I_21558 (I370082,I370074,I369746);
DFFARX1 I_21559 (I370082,I3563,I369720,I369685,);
DFFARX1 I_21560 (I370074,I3563,I369720,I369703,);
nor I_21561 (I370127,I713344,I713338);
not I_21562 (I370144,I370127);
nor I_21563 (I369706,I369983,I370144);
nand I_21564 (I369691,I370000,I370144);
nor I_21565 (I369700,I369746,I370127);
DFFARX1 I_21566 (I370127,I3563,I369720,I369709,);
not I_21567 (I370247,I3570);
DFFARX1 I_21568 (I751483,I3563,I370247,I370273,);
nand I_21569 (I370281,I751474,I751489);
and I_21570 (I370298,I370281,I751495);
DFFARX1 I_21571 (I370298,I3563,I370247,I370324,);
nor I_21572 (I370215,I370324,I370273);
not I_21573 (I370346,I370324);
DFFARX1 I_21574 (I751480,I3563,I370247,I370372,);
nand I_21575 (I370380,I370372,I751474);
not I_21576 (I370397,I370380);
DFFARX1 I_21577 (I370397,I3563,I370247,I370423,);
not I_21578 (I370239,I370423);
nor I_21579 (I370445,I370273,I370380);
nor I_21580 (I370221,I370324,I370445);
DFFARX1 I_21581 (I751477,I3563,I370247,I370485,);
DFFARX1 I_21582 (I370485,I3563,I370247,I370502,);
not I_21583 (I370510,I370502);
not I_21584 (I370527,I370485);
nand I_21585 (I370224,I370527,I370346);
nand I_21586 (I370558,I751471,I751486);
and I_21587 (I370575,I370558,I751471);
DFFARX1 I_21588 (I370575,I3563,I370247,I370601,);
nor I_21589 (I370609,I370601,I370273);
DFFARX1 I_21590 (I370609,I3563,I370247,I370212,);
DFFARX1 I_21591 (I370601,I3563,I370247,I370230,);
nor I_21592 (I370654,I751492,I751486);
not I_21593 (I370671,I370654);
nor I_21594 (I370233,I370510,I370671);
nand I_21595 (I370218,I370527,I370671);
nor I_21596 (I370227,I370273,I370654);
DFFARX1 I_21597 (I370654,I3563,I370247,I370236,);
not I_21598 (I370774,I3570);
DFFARX1 I_21599 (I149402,I3563,I370774,I370800,);
nand I_21600 (I370808,I149414,I149423);
and I_21601 (I370825,I370808,I149402);
DFFARX1 I_21602 (I370825,I3563,I370774,I370851,);
nor I_21603 (I370742,I370851,I370800);
not I_21604 (I370873,I370851);
DFFARX1 I_21605 (I149417,I3563,I370774,I370899,);
nand I_21606 (I370907,I370899,I149405);
not I_21607 (I370924,I370907);
DFFARX1 I_21608 (I370924,I3563,I370774,I370950,);
not I_21609 (I370766,I370950);
nor I_21610 (I370972,I370800,I370907);
nor I_21611 (I370748,I370851,I370972);
DFFARX1 I_21612 (I149408,I3563,I370774,I371012,);
DFFARX1 I_21613 (I371012,I3563,I370774,I371029,);
not I_21614 (I371037,I371029);
not I_21615 (I371054,I371012);
nand I_21616 (I370751,I371054,I370873);
nand I_21617 (I371085,I149399,I149399);
and I_21618 (I371102,I371085,I149411);
DFFARX1 I_21619 (I371102,I3563,I370774,I371128,);
nor I_21620 (I371136,I371128,I370800);
DFFARX1 I_21621 (I371136,I3563,I370774,I370739,);
DFFARX1 I_21622 (I371128,I3563,I370774,I370757,);
nor I_21623 (I371181,I149420,I149399);
not I_21624 (I371198,I371181);
nor I_21625 (I370760,I371037,I371198);
nand I_21626 (I370745,I371054,I371198);
nor I_21627 (I370754,I370800,I371181);
DFFARX1 I_21628 (I371181,I3563,I370774,I370763,);
not I_21629 (I371301,I3570);
DFFARX1 I_21630 (I939426,I3563,I371301,I371327,);
nand I_21631 (I371335,I939423,I939441);
and I_21632 (I371352,I371335,I939432);
DFFARX1 I_21633 (I371352,I3563,I371301,I371378,);
nor I_21634 (I371269,I371378,I371327);
not I_21635 (I371400,I371378);
DFFARX1 I_21636 (I939447,I3563,I371301,I371426,);
nand I_21637 (I371434,I371426,I939429);
not I_21638 (I371451,I371434);
DFFARX1 I_21639 (I371451,I3563,I371301,I371477,);
not I_21640 (I371293,I371477);
nor I_21641 (I371499,I371327,I371434);
nor I_21642 (I371275,I371378,I371499);
DFFARX1 I_21643 (I939435,I3563,I371301,I371539,);
DFFARX1 I_21644 (I371539,I3563,I371301,I371556,);
not I_21645 (I371564,I371556);
not I_21646 (I371581,I371539);
nand I_21647 (I371278,I371581,I371400);
nand I_21648 (I371612,I939423,I939450);
and I_21649 (I371629,I371612,I939438);
DFFARX1 I_21650 (I371629,I3563,I371301,I371655,);
nor I_21651 (I371663,I371655,I371327);
DFFARX1 I_21652 (I371663,I3563,I371301,I371266,);
DFFARX1 I_21653 (I371655,I3563,I371301,I371284,);
nor I_21654 (I371708,I939444,I939450);
not I_21655 (I371725,I371708);
nor I_21656 (I371287,I371564,I371725);
nand I_21657 (I371272,I371581,I371725);
nor I_21658 (I371281,I371327,I371708);
DFFARX1 I_21659 (I371708,I3563,I371301,I371290,);
not I_21660 (I371828,I3570);
DFFARX1 I_21661 (I735299,I3563,I371828,I371854,);
nand I_21662 (I371862,I735290,I735305);
and I_21663 (I371879,I371862,I735311);
DFFARX1 I_21664 (I371879,I3563,I371828,I371905,);
nor I_21665 (I371796,I371905,I371854);
not I_21666 (I371927,I371905);
DFFARX1 I_21667 (I735296,I3563,I371828,I371953,);
nand I_21668 (I371961,I371953,I735290);
not I_21669 (I371978,I371961);
DFFARX1 I_21670 (I371978,I3563,I371828,I372004,);
not I_21671 (I371820,I372004);
nor I_21672 (I372026,I371854,I371961);
nor I_21673 (I371802,I371905,I372026);
DFFARX1 I_21674 (I735293,I3563,I371828,I372066,);
DFFARX1 I_21675 (I372066,I3563,I371828,I372083,);
not I_21676 (I372091,I372083);
not I_21677 (I372108,I372066);
nand I_21678 (I371805,I372108,I371927);
nand I_21679 (I372139,I735287,I735302);
and I_21680 (I372156,I372139,I735287);
DFFARX1 I_21681 (I372156,I3563,I371828,I372182,);
nor I_21682 (I372190,I372182,I371854);
DFFARX1 I_21683 (I372190,I3563,I371828,I371793,);
DFFARX1 I_21684 (I372182,I3563,I371828,I371811,);
nor I_21685 (I372235,I735308,I735302);
not I_21686 (I372252,I372235);
nor I_21687 (I371814,I372091,I372252);
nand I_21688 (I371799,I372108,I372252);
nor I_21689 (I371808,I371854,I372235);
DFFARX1 I_21690 (I372235,I3563,I371828,I371817,);
not I_21691 (I372355,I3570);
DFFARX1 I_21692 (I1123941,I3563,I372355,I372381,);
nand I_21693 (I372389,I1123956,I1123941);
and I_21694 (I372406,I372389,I1123959);
DFFARX1 I_21695 (I372406,I3563,I372355,I372432,);
nor I_21696 (I372323,I372432,I372381);
not I_21697 (I372454,I372432);
DFFARX1 I_21698 (I1123965,I3563,I372355,I372480,);
nand I_21699 (I372488,I372480,I1123947);
not I_21700 (I372505,I372488);
DFFARX1 I_21701 (I372505,I3563,I372355,I372531,);
not I_21702 (I372347,I372531);
nor I_21703 (I372553,I372381,I372488);
nor I_21704 (I372329,I372432,I372553);
DFFARX1 I_21705 (I1123944,I3563,I372355,I372593,);
DFFARX1 I_21706 (I372593,I3563,I372355,I372610,);
not I_21707 (I372618,I372610);
not I_21708 (I372635,I372593);
nand I_21709 (I372332,I372635,I372454);
nand I_21710 (I372666,I1123944,I1123950);
and I_21711 (I372683,I372666,I1123962);
DFFARX1 I_21712 (I372683,I3563,I372355,I372709,);
nor I_21713 (I372717,I372709,I372381);
DFFARX1 I_21714 (I372717,I3563,I372355,I372320,);
DFFARX1 I_21715 (I372709,I3563,I372355,I372338,);
nor I_21716 (I372762,I1123953,I1123950);
not I_21717 (I372779,I372762);
nor I_21718 (I372341,I372618,I372779);
nand I_21719 (I372326,I372635,I372779);
nor I_21720 (I372335,I372381,I372762);
DFFARX1 I_21721 (I372762,I3563,I372355,I372344,);
not I_21722 (I372882,I3570);
DFFARX1 I_21723 (I163142,I3563,I372882,I372908,);
nand I_21724 (I372916,I163127,I163118);
and I_21725 (I372933,I372916,I163133);
DFFARX1 I_21726 (I372933,I3563,I372882,I372959,);
nor I_21727 (I372850,I372959,I372908);
not I_21728 (I372981,I372959);
DFFARX1 I_21729 (I163145,I3563,I372882,I373007,);
nand I_21730 (I373015,I373007,I163136);
not I_21731 (I373032,I373015);
DFFARX1 I_21732 (I373032,I3563,I372882,I373058,);
not I_21733 (I372874,I373058);
nor I_21734 (I373080,I372908,I373015);
nor I_21735 (I372856,I372959,I373080);
DFFARX1 I_21736 (I163124,I3563,I372882,I373120,);
DFFARX1 I_21737 (I373120,I3563,I372882,I373137,);
not I_21738 (I373145,I373137);
not I_21739 (I373162,I373120);
nand I_21740 (I372859,I373162,I372981);
nand I_21741 (I373193,I163130,I163121);
and I_21742 (I373210,I373193,I163118);
DFFARX1 I_21743 (I373210,I3563,I372882,I373236,);
nor I_21744 (I373244,I373236,I372908);
DFFARX1 I_21745 (I373244,I3563,I372882,I372847,);
DFFARX1 I_21746 (I373236,I3563,I372882,I372865,);
nor I_21747 (I373289,I163139,I163121);
not I_21748 (I373306,I373289);
nor I_21749 (I372868,I373145,I373306);
nand I_21750 (I372853,I373162,I373306);
nor I_21751 (I372862,I372908,I373289);
DFFARX1 I_21752 (I373289,I3563,I372882,I372871,);
not I_21753 (I373409,I3570);
DFFARX1 I_21754 (I1093307,I3563,I373409,I373435,);
nand I_21755 (I373443,I1093322,I1093307);
and I_21756 (I373460,I373443,I1093325);
DFFARX1 I_21757 (I373460,I3563,I373409,I373486,);
nor I_21758 (I373377,I373486,I373435);
not I_21759 (I373508,I373486);
DFFARX1 I_21760 (I1093331,I3563,I373409,I373534,);
nand I_21761 (I373542,I373534,I1093313);
not I_21762 (I373559,I373542);
DFFARX1 I_21763 (I373559,I3563,I373409,I373585,);
not I_21764 (I373401,I373585);
nor I_21765 (I373607,I373435,I373542);
nor I_21766 (I373383,I373486,I373607);
DFFARX1 I_21767 (I1093310,I3563,I373409,I373647,);
DFFARX1 I_21768 (I373647,I3563,I373409,I373664,);
not I_21769 (I373672,I373664);
not I_21770 (I373689,I373647);
nand I_21771 (I373386,I373689,I373508);
nand I_21772 (I373720,I1093310,I1093316);
and I_21773 (I373737,I373720,I1093328);
DFFARX1 I_21774 (I373737,I3563,I373409,I373763,);
nor I_21775 (I373771,I373763,I373435);
DFFARX1 I_21776 (I373771,I3563,I373409,I373374,);
DFFARX1 I_21777 (I373763,I3563,I373409,I373392,);
nor I_21778 (I373816,I1093319,I1093316);
not I_21779 (I373833,I373816);
nor I_21780 (I373395,I373672,I373833);
nand I_21781 (I373380,I373689,I373833);
nor I_21782 (I373389,I373435,I373816);
DFFARX1 I_21783 (I373816,I3563,I373409,I373398,);
not I_21784 (I373936,I3570);
DFFARX1 I_21785 (I1373199,I3563,I373936,I373962,);
nand I_21786 (I373970,I1373178,I1373178);
and I_21787 (I373987,I373970,I1373205);
DFFARX1 I_21788 (I373987,I3563,I373936,I374013,);
nor I_21789 (I373904,I374013,I373962);
not I_21790 (I374035,I374013);
DFFARX1 I_21791 (I1373193,I3563,I373936,I374061,);
nand I_21792 (I374069,I374061,I1373196);
not I_21793 (I374086,I374069);
DFFARX1 I_21794 (I374086,I3563,I373936,I374112,);
not I_21795 (I373928,I374112);
nor I_21796 (I374134,I373962,I374069);
nor I_21797 (I373910,I374013,I374134);
DFFARX1 I_21798 (I1373187,I3563,I373936,I374174,);
DFFARX1 I_21799 (I374174,I3563,I373936,I374191,);
not I_21800 (I374199,I374191);
not I_21801 (I374216,I374174);
nand I_21802 (I373913,I374216,I374035);
nand I_21803 (I374247,I1373184,I1373181);
and I_21804 (I374264,I374247,I1373202);
DFFARX1 I_21805 (I374264,I3563,I373936,I374290,);
nor I_21806 (I374298,I374290,I373962);
DFFARX1 I_21807 (I374298,I3563,I373936,I373901,);
DFFARX1 I_21808 (I374290,I3563,I373936,I373919,);
nor I_21809 (I374343,I1373190,I1373181);
not I_21810 (I374360,I374343);
nor I_21811 (I373922,I374199,I374360);
nand I_21812 (I373907,I374216,I374360);
nor I_21813 (I373916,I373962,I374343);
DFFARX1 I_21814 (I374343,I3563,I373936,I373925,);
not I_21815 (I374463,I3570);
DFFARX1 I_21816 (I978832,I3563,I374463,I374489,);
nand I_21817 (I374497,I978829,I978847);
and I_21818 (I374514,I374497,I978838);
DFFARX1 I_21819 (I374514,I3563,I374463,I374540,);
nor I_21820 (I374431,I374540,I374489);
not I_21821 (I374562,I374540);
DFFARX1 I_21822 (I978853,I3563,I374463,I374588,);
nand I_21823 (I374596,I374588,I978835);
not I_21824 (I374613,I374596);
DFFARX1 I_21825 (I374613,I3563,I374463,I374639,);
not I_21826 (I374455,I374639);
nor I_21827 (I374661,I374489,I374596);
nor I_21828 (I374437,I374540,I374661);
DFFARX1 I_21829 (I978841,I3563,I374463,I374701,);
DFFARX1 I_21830 (I374701,I3563,I374463,I374718,);
not I_21831 (I374726,I374718);
not I_21832 (I374743,I374701);
nand I_21833 (I374440,I374743,I374562);
nand I_21834 (I374774,I978829,I978856);
and I_21835 (I374791,I374774,I978844);
DFFARX1 I_21836 (I374791,I3563,I374463,I374817,);
nor I_21837 (I374825,I374817,I374489);
DFFARX1 I_21838 (I374825,I3563,I374463,I374428,);
DFFARX1 I_21839 (I374817,I3563,I374463,I374446,);
nor I_21840 (I374870,I978850,I978856);
not I_21841 (I374887,I374870);
nor I_21842 (I374449,I374726,I374887);
nand I_21843 (I374434,I374743,I374887);
nor I_21844 (I374443,I374489,I374870);
DFFARX1 I_21845 (I374870,I3563,I374463,I374452,);
not I_21846 (I374990,I3570);
DFFARX1 I_21847 (I1107179,I3563,I374990,I375016,);
nand I_21848 (I375024,I1107194,I1107179);
and I_21849 (I375041,I375024,I1107197);
DFFARX1 I_21850 (I375041,I3563,I374990,I375067,);
nor I_21851 (I374958,I375067,I375016);
not I_21852 (I375089,I375067);
DFFARX1 I_21853 (I1107203,I3563,I374990,I375115,);
nand I_21854 (I375123,I375115,I1107185);
not I_21855 (I375140,I375123);
DFFARX1 I_21856 (I375140,I3563,I374990,I375166,);
not I_21857 (I374982,I375166);
nor I_21858 (I375188,I375016,I375123);
nor I_21859 (I374964,I375067,I375188);
DFFARX1 I_21860 (I1107182,I3563,I374990,I375228,);
DFFARX1 I_21861 (I375228,I3563,I374990,I375245,);
not I_21862 (I375253,I375245);
not I_21863 (I375270,I375228);
nand I_21864 (I374967,I375270,I375089);
nand I_21865 (I375301,I1107182,I1107188);
and I_21866 (I375318,I375301,I1107200);
DFFARX1 I_21867 (I375318,I3563,I374990,I375344,);
nor I_21868 (I375352,I375344,I375016);
DFFARX1 I_21869 (I375352,I3563,I374990,I374955,);
DFFARX1 I_21870 (I375344,I3563,I374990,I374973,);
nor I_21871 (I375397,I1107191,I1107188);
not I_21872 (I375414,I375397);
nor I_21873 (I374976,I375253,I375414);
nand I_21874 (I374961,I375270,I375414);
nor I_21875 (I374970,I375016,I375397);
DFFARX1 I_21876 (I375397,I3563,I374990,I374979,);
not I_21877 (I375517,I3570);
DFFARX1 I_21878 (I676343,I3563,I375517,I375543,);
nand I_21879 (I375551,I676334,I676349);
and I_21880 (I375568,I375551,I676355);
DFFARX1 I_21881 (I375568,I3563,I375517,I375594,);
nor I_21882 (I375485,I375594,I375543);
not I_21883 (I375616,I375594);
DFFARX1 I_21884 (I676340,I3563,I375517,I375642,);
nand I_21885 (I375650,I375642,I676334);
not I_21886 (I375667,I375650);
DFFARX1 I_21887 (I375667,I3563,I375517,I375693,);
not I_21888 (I375509,I375693);
nor I_21889 (I375715,I375543,I375650);
nor I_21890 (I375491,I375594,I375715);
DFFARX1 I_21891 (I676337,I3563,I375517,I375755,);
DFFARX1 I_21892 (I375755,I3563,I375517,I375772,);
not I_21893 (I375780,I375772);
not I_21894 (I375797,I375755);
nand I_21895 (I375494,I375797,I375616);
nand I_21896 (I375828,I676331,I676346);
and I_21897 (I375845,I375828,I676331);
DFFARX1 I_21898 (I375845,I3563,I375517,I375871,);
nor I_21899 (I375879,I375871,I375543);
DFFARX1 I_21900 (I375879,I3563,I375517,I375482,);
DFFARX1 I_21901 (I375871,I3563,I375517,I375500,);
nor I_21902 (I375924,I676352,I676346);
not I_21903 (I375941,I375924);
nor I_21904 (I375503,I375780,I375941);
nand I_21905 (I375488,I375797,I375941);
nor I_21906 (I375497,I375543,I375924);
DFFARX1 I_21907 (I375924,I3563,I375517,I375506,);
not I_21908 (I376044,I3570);
DFFARX1 I_21909 (I678655,I3563,I376044,I376070,);
nand I_21910 (I376078,I678646,I678661);
and I_21911 (I376095,I376078,I678667);
DFFARX1 I_21912 (I376095,I3563,I376044,I376121,);
nor I_21913 (I376012,I376121,I376070);
not I_21914 (I376143,I376121);
DFFARX1 I_21915 (I678652,I3563,I376044,I376169,);
nand I_21916 (I376177,I376169,I678646);
not I_21917 (I376194,I376177);
DFFARX1 I_21918 (I376194,I3563,I376044,I376220,);
not I_21919 (I376036,I376220);
nor I_21920 (I376242,I376070,I376177);
nor I_21921 (I376018,I376121,I376242);
DFFARX1 I_21922 (I678649,I3563,I376044,I376282,);
DFFARX1 I_21923 (I376282,I3563,I376044,I376299,);
not I_21924 (I376307,I376299);
not I_21925 (I376324,I376282);
nand I_21926 (I376021,I376324,I376143);
nand I_21927 (I376355,I678643,I678658);
and I_21928 (I376372,I376355,I678643);
DFFARX1 I_21929 (I376372,I3563,I376044,I376398,);
nor I_21930 (I376406,I376398,I376070);
DFFARX1 I_21931 (I376406,I3563,I376044,I376009,);
DFFARX1 I_21932 (I376398,I3563,I376044,I376027,);
nor I_21933 (I376451,I678664,I678658);
not I_21934 (I376468,I376451);
nor I_21935 (I376030,I376307,I376468);
nand I_21936 (I376015,I376324,I376468);
nor I_21937 (I376024,I376070,I376451);
DFFARX1 I_21938 (I376451,I3563,I376044,I376033,);
not I_21939 (I376571,I3570);
DFFARX1 I_21940 (I1153997,I3563,I376571,I376597,);
nand I_21941 (I376605,I1154012,I1153997);
and I_21942 (I376622,I376605,I1154015);
DFFARX1 I_21943 (I376622,I3563,I376571,I376648,);
nor I_21944 (I376539,I376648,I376597);
not I_21945 (I376670,I376648);
DFFARX1 I_21946 (I1154021,I3563,I376571,I376696,);
nand I_21947 (I376704,I376696,I1154003);
not I_21948 (I376721,I376704);
DFFARX1 I_21949 (I376721,I3563,I376571,I376747,);
not I_21950 (I376563,I376747);
nor I_21951 (I376769,I376597,I376704);
nor I_21952 (I376545,I376648,I376769);
DFFARX1 I_21953 (I1154000,I3563,I376571,I376809,);
DFFARX1 I_21954 (I376809,I3563,I376571,I376826,);
not I_21955 (I376834,I376826);
not I_21956 (I376851,I376809);
nand I_21957 (I376548,I376851,I376670);
nand I_21958 (I376882,I1154000,I1154006);
and I_21959 (I376899,I376882,I1154018);
DFFARX1 I_21960 (I376899,I3563,I376571,I376925,);
nor I_21961 (I376933,I376925,I376597);
DFFARX1 I_21962 (I376933,I3563,I376571,I376536,);
DFFARX1 I_21963 (I376925,I3563,I376571,I376554,);
nor I_21964 (I376978,I1154009,I1154006);
not I_21965 (I376995,I376978);
nor I_21966 (I376557,I376834,I376995);
nand I_21967 (I376542,I376851,I376995);
nor I_21968 (I376551,I376597,I376978);
DFFARX1 I_21969 (I376978,I3563,I376571,I376560,);
not I_21970 (I377098,I3570);
DFFARX1 I_21971 (I502926,I3563,I377098,I377124,);
nand I_21972 (I377132,I502938,I502917);
and I_21973 (I377149,I377132,I502941);
DFFARX1 I_21974 (I377149,I3563,I377098,I377175,);
nor I_21975 (I377066,I377175,I377124);
not I_21976 (I377197,I377175);
DFFARX1 I_21977 (I502932,I3563,I377098,I377223,);
nand I_21978 (I377231,I377223,I502914);
not I_21979 (I377248,I377231);
DFFARX1 I_21980 (I377248,I3563,I377098,I377274,);
not I_21981 (I377090,I377274);
nor I_21982 (I377296,I377124,I377231);
nor I_21983 (I377072,I377175,I377296);
DFFARX1 I_21984 (I502929,I3563,I377098,I377336,);
DFFARX1 I_21985 (I377336,I3563,I377098,I377353,);
not I_21986 (I377361,I377353);
not I_21987 (I377378,I377336);
nand I_21988 (I377075,I377378,I377197);
nand I_21989 (I377409,I502914,I502920);
and I_21990 (I377426,I377409,I502923);
DFFARX1 I_21991 (I377426,I3563,I377098,I377452,);
nor I_21992 (I377460,I377452,I377124);
DFFARX1 I_21993 (I377460,I3563,I377098,I377063,);
DFFARX1 I_21994 (I377452,I3563,I377098,I377081,);
nor I_21995 (I377505,I502935,I502920);
not I_21996 (I377522,I377505);
nor I_21997 (I377084,I377361,I377522);
nand I_21998 (I377069,I377378,I377522);
nor I_21999 (I377078,I377124,I377505);
DFFARX1 I_22000 (I377505,I3563,I377098,I377087,);
not I_22001 (I377625,I3570);
DFFARX1 I_22002 (I825288,I3563,I377625,I377651,);
nand I_22003 (I377659,I825291,I825285);
and I_22004 (I377676,I377659,I825297);
DFFARX1 I_22005 (I377676,I3563,I377625,I377702,);
nor I_22006 (I377593,I377702,I377651);
not I_22007 (I377724,I377702);
DFFARX1 I_22008 (I825300,I3563,I377625,I377750,);
nand I_22009 (I377758,I377750,I825291);
not I_22010 (I377775,I377758);
DFFARX1 I_22011 (I377775,I3563,I377625,I377801,);
not I_22012 (I377617,I377801);
nor I_22013 (I377823,I377651,I377758);
nor I_22014 (I377599,I377702,I377823);
DFFARX1 I_22015 (I825303,I3563,I377625,I377863,);
DFFARX1 I_22016 (I377863,I3563,I377625,I377880,);
not I_22017 (I377888,I377880);
not I_22018 (I377905,I377863);
nand I_22019 (I377602,I377905,I377724);
nand I_22020 (I377936,I825285,I825294);
and I_22021 (I377953,I377936,I825288);
DFFARX1 I_22022 (I377953,I3563,I377625,I377979,);
nor I_22023 (I377987,I377979,I377651);
DFFARX1 I_22024 (I377987,I3563,I377625,I377590,);
DFFARX1 I_22025 (I377979,I3563,I377625,I377608,);
nor I_22026 (I378032,I825306,I825294);
not I_22027 (I378049,I378032);
nor I_22028 (I377611,I377888,I378049);
nand I_22029 (I377596,I377905,I378049);
nor I_22030 (I377605,I377651,I378032);
DFFARX1 I_22031 (I378032,I3563,I377625,I377614,);
not I_22032 (I378152,I3570);
DFFARX1 I_22033 (I945886,I3563,I378152,I378178,);
nand I_22034 (I378186,I945883,I945901);
and I_22035 (I378203,I378186,I945892);
DFFARX1 I_22036 (I378203,I3563,I378152,I378229,);
nor I_22037 (I378120,I378229,I378178);
not I_22038 (I378251,I378229);
DFFARX1 I_22039 (I945907,I3563,I378152,I378277,);
nand I_22040 (I378285,I378277,I945889);
not I_22041 (I378302,I378285);
DFFARX1 I_22042 (I378302,I3563,I378152,I378328,);
not I_22043 (I378144,I378328);
nor I_22044 (I378350,I378178,I378285);
nor I_22045 (I378126,I378229,I378350);
DFFARX1 I_22046 (I945895,I3563,I378152,I378390,);
DFFARX1 I_22047 (I378390,I3563,I378152,I378407,);
not I_22048 (I378415,I378407);
not I_22049 (I378432,I378390);
nand I_22050 (I378129,I378432,I378251);
nand I_22051 (I378463,I945883,I945910);
and I_22052 (I378480,I378463,I945898);
DFFARX1 I_22053 (I378480,I3563,I378152,I378506,);
nor I_22054 (I378514,I378506,I378178);
DFFARX1 I_22055 (I378514,I3563,I378152,I378117,);
DFFARX1 I_22056 (I378506,I3563,I378152,I378135,);
nor I_22057 (I378559,I945904,I945910);
not I_22058 (I378576,I378559);
nor I_22059 (I378138,I378415,I378576);
nand I_22060 (I378123,I378432,I378576);
nor I_22061 (I378132,I378178,I378559);
DFFARX1 I_22062 (I378559,I3563,I378152,I378141,);
not I_22063 (I378679,I3570);
DFFARX1 I_22064 (I716803,I3563,I378679,I378705,);
nand I_22065 (I378713,I716794,I716809);
and I_22066 (I378730,I378713,I716815);
DFFARX1 I_22067 (I378730,I3563,I378679,I378756,);
nor I_22068 (I378647,I378756,I378705);
not I_22069 (I378778,I378756);
DFFARX1 I_22070 (I716800,I3563,I378679,I378804,);
nand I_22071 (I378812,I378804,I716794);
not I_22072 (I378829,I378812);
DFFARX1 I_22073 (I378829,I3563,I378679,I378855,);
not I_22074 (I378671,I378855);
nor I_22075 (I378877,I378705,I378812);
nor I_22076 (I378653,I378756,I378877);
DFFARX1 I_22077 (I716797,I3563,I378679,I378917,);
DFFARX1 I_22078 (I378917,I3563,I378679,I378934,);
not I_22079 (I378942,I378934);
not I_22080 (I378959,I378917);
nand I_22081 (I378656,I378959,I378778);
nand I_22082 (I378990,I716791,I716806);
and I_22083 (I379007,I378990,I716791);
DFFARX1 I_22084 (I379007,I3563,I378679,I379033,);
nor I_22085 (I379041,I379033,I378705);
DFFARX1 I_22086 (I379041,I3563,I378679,I378644,);
DFFARX1 I_22087 (I379033,I3563,I378679,I378662,);
nor I_22088 (I379086,I716812,I716806);
not I_22089 (I379103,I379086);
nor I_22090 (I378665,I378942,I379103);
nand I_22091 (I378650,I378959,I379103);
nor I_22092 (I378659,I378705,I379086);
DFFARX1 I_22093 (I379086,I3563,I378679,I378668,);
not I_22094 (I379206,I3570);
DFFARX1 I_22095 (I461582,I3563,I379206,I379232,);
nand I_22096 (I379240,I461594,I461573);
and I_22097 (I379257,I379240,I461597);
DFFARX1 I_22098 (I379257,I3563,I379206,I379283,);
nor I_22099 (I379174,I379283,I379232);
not I_22100 (I379305,I379283);
DFFARX1 I_22101 (I461588,I3563,I379206,I379331,);
nand I_22102 (I379339,I379331,I461570);
not I_22103 (I379356,I379339);
DFFARX1 I_22104 (I379356,I3563,I379206,I379382,);
not I_22105 (I379198,I379382);
nor I_22106 (I379404,I379232,I379339);
nor I_22107 (I379180,I379283,I379404);
DFFARX1 I_22108 (I461585,I3563,I379206,I379444,);
DFFARX1 I_22109 (I379444,I3563,I379206,I379461,);
not I_22110 (I379469,I379461);
not I_22111 (I379486,I379444);
nand I_22112 (I379183,I379486,I379305);
nand I_22113 (I379517,I461570,I461576);
and I_22114 (I379534,I379517,I461579);
DFFARX1 I_22115 (I379534,I3563,I379206,I379560,);
nor I_22116 (I379568,I379560,I379232);
DFFARX1 I_22117 (I379568,I3563,I379206,I379171,);
DFFARX1 I_22118 (I379560,I3563,I379206,I379189,);
nor I_22119 (I379613,I461591,I461576);
not I_22120 (I379630,I379613);
nor I_22121 (I379192,I379469,I379630);
nand I_22122 (I379177,I379486,I379630);
nor I_22123 (I379186,I379232,I379613);
DFFARX1 I_22124 (I379613,I3563,I379206,I379195,);
not I_22125 (I379733,I3570);
DFFARX1 I_22126 (I3196,I3563,I379733,I379759,);
nand I_22127 (I379767,I3492,I3260);
and I_22128 (I379784,I379767,I2308);
DFFARX1 I_22129 (I379784,I3563,I379733,I379810,);
nor I_22130 (I379701,I379810,I379759);
not I_22131 (I379832,I379810);
DFFARX1 I_22132 (I1884,I3563,I379733,I379858,);
nand I_22133 (I379866,I379858,I2052);
not I_22134 (I379883,I379866);
DFFARX1 I_22135 (I379883,I3563,I379733,I379909,);
not I_22136 (I379725,I379909);
nor I_22137 (I379931,I379759,I379866);
nor I_22138 (I379707,I379810,I379931);
DFFARX1 I_22139 (I1844,I3563,I379733,I379971,);
DFFARX1 I_22140 (I379971,I3563,I379733,I379988,);
not I_22141 (I379996,I379988);
not I_22142 (I380013,I379971);
nand I_22143 (I379710,I380013,I379832);
nand I_22144 (I380044,I1892,I2492);
and I_22145 (I380061,I380044,I1748);
DFFARX1 I_22146 (I380061,I3563,I379733,I380087,);
nor I_22147 (I380095,I380087,I379759);
DFFARX1 I_22148 (I380095,I3563,I379733,I379698,);
DFFARX1 I_22149 (I380087,I3563,I379733,I379716,);
nor I_22150 (I380140,I2108,I2492);
not I_22151 (I380157,I380140);
nor I_22152 (I379719,I379996,I380157);
nand I_22153 (I379704,I380013,I380157);
nor I_22154 (I379713,I379759,I380140);
DFFARX1 I_22155 (I380140,I3563,I379733,I379722,);
not I_22156 (I380260,I3570);
DFFARX1 I_22157 (I1159777,I3563,I380260,I380286,);
nand I_22158 (I380294,I1159792,I1159777);
and I_22159 (I380311,I380294,I1159795);
DFFARX1 I_22160 (I380311,I3563,I380260,I380337,);
nor I_22161 (I380228,I380337,I380286);
not I_22162 (I380359,I380337);
DFFARX1 I_22163 (I1159801,I3563,I380260,I380385,);
nand I_22164 (I380393,I380385,I1159783);
not I_22165 (I380410,I380393);
DFFARX1 I_22166 (I380410,I3563,I380260,I380436,);
not I_22167 (I380252,I380436);
nor I_22168 (I380458,I380286,I380393);
nor I_22169 (I380234,I380337,I380458);
DFFARX1 I_22170 (I1159780,I3563,I380260,I380498,);
DFFARX1 I_22171 (I380498,I3563,I380260,I380515,);
not I_22172 (I380523,I380515);
not I_22173 (I380540,I380498);
nand I_22174 (I380237,I380540,I380359);
nand I_22175 (I380571,I1159780,I1159786);
and I_22176 (I380588,I380571,I1159798);
DFFARX1 I_22177 (I380588,I3563,I380260,I380614,);
nor I_22178 (I380622,I380614,I380286);
DFFARX1 I_22179 (I380622,I3563,I380260,I380225,);
DFFARX1 I_22180 (I380614,I3563,I380260,I380243,);
nor I_22181 (I380667,I1159789,I1159786);
not I_22182 (I380684,I380667);
nor I_22183 (I380246,I380523,I380684);
nand I_22184 (I380231,I380540,I380684);
nor I_22185 (I380240,I380286,I380667);
DFFARX1 I_22186 (I380667,I3563,I380260,I380249,);
not I_22187 (I380787,I3570);
DFFARX1 I_22188 (I770557,I3563,I380787,I380813,);
nand I_22189 (I380821,I770548,I770563);
and I_22190 (I380838,I380821,I770569);
DFFARX1 I_22191 (I380838,I3563,I380787,I380864,);
nor I_22192 (I380755,I380864,I380813);
not I_22193 (I380886,I380864);
DFFARX1 I_22194 (I770554,I3563,I380787,I380912,);
nand I_22195 (I380920,I380912,I770548);
not I_22196 (I380937,I380920);
DFFARX1 I_22197 (I380937,I3563,I380787,I380963,);
not I_22198 (I380779,I380963);
nor I_22199 (I380985,I380813,I380920);
nor I_22200 (I380761,I380864,I380985);
DFFARX1 I_22201 (I770551,I3563,I380787,I381025,);
DFFARX1 I_22202 (I381025,I3563,I380787,I381042,);
not I_22203 (I381050,I381042);
not I_22204 (I381067,I381025);
nand I_22205 (I380764,I381067,I380886);
nand I_22206 (I381098,I770545,I770560);
and I_22207 (I381115,I381098,I770545);
DFFARX1 I_22208 (I381115,I3563,I380787,I381141,);
nor I_22209 (I381149,I381141,I380813);
DFFARX1 I_22210 (I381149,I3563,I380787,I380752,);
DFFARX1 I_22211 (I381141,I3563,I380787,I380770,);
nor I_22212 (I381194,I770566,I770560);
not I_22213 (I381211,I381194);
nor I_22214 (I380773,I381050,I381211);
nand I_22215 (I380758,I381067,I381211);
nor I_22216 (I380767,I380813,I381194);
DFFARX1 I_22217 (I381194,I3563,I380787,I380776,);
not I_22218 (I381314,I3570);
DFFARX1 I_22219 (I644556,I3563,I381314,I381340,);
nand I_22220 (I381348,I644541,I644544);
and I_22221 (I381365,I381348,I644559);
DFFARX1 I_22222 (I381365,I3563,I381314,I381391,);
nor I_22223 (I381282,I381391,I381340);
not I_22224 (I381413,I381391);
DFFARX1 I_22225 (I644553,I3563,I381314,I381439,);
nand I_22226 (I381447,I381439,I644544);
not I_22227 (I381464,I381447);
DFFARX1 I_22228 (I381464,I3563,I381314,I381490,);
not I_22229 (I381306,I381490);
nor I_22230 (I381512,I381340,I381447);
nor I_22231 (I381288,I381391,I381512);
DFFARX1 I_22232 (I644550,I3563,I381314,I381552,);
DFFARX1 I_22233 (I381552,I3563,I381314,I381569,);
not I_22234 (I381577,I381569);
not I_22235 (I381594,I381552);
nand I_22236 (I381291,I381594,I381413);
nand I_22237 (I381625,I644565,I644541);
and I_22238 (I381642,I381625,I644562);
DFFARX1 I_22239 (I381642,I3563,I381314,I381668,);
nor I_22240 (I381676,I381668,I381340);
DFFARX1 I_22241 (I381676,I3563,I381314,I381279,);
DFFARX1 I_22242 (I381668,I3563,I381314,I381297,);
nor I_22243 (I381721,I644547,I644541);
not I_22244 (I381738,I381721);
nor I_22245 (I381300,I381577,I381738);
nand I_22246 (I381285,I381594,I381738);
nor I_22247 (I381294,I381340,I381721);
DFFARX1 I_22248 (I381721,I3563,I381314,I381303,);
not I_22249 (I381841,I3570);
DFFARX1 I_22250 (I137808,I3563,I381841,I381867,);
nand I_22251 (I381875,I137820,I137829);
and I_22252 (I381892,I381875,I137808);
DFFARX1 I_22253 (I381892,I3563,I381841,I381918,);
nor I_22254 (I381809,I381918,I381867);
not I_22255 (I381940,I381918);
DFFARX1 I_22256 (I137823,I3563,I381841,I381966,);
nand I_22257 (I381974,I381966,I137811);
not I_22258 (I381991,I381974);
DFFARX1 I_22259 (I381991,I3563,I381841,I382017,);
not I_22260 (I381833,I382017);
nor I_22261 (I382039,I381867,I381974);
nor I_22262 (I381815,I381918,I382039);
DFFARX1 I_22263 (I137814,I3563,I381841,I382079,);
DFFARX1 I_22264 (I382079,I3563,I381841,I382096,);
not I_22265 (I382104,I382096);
not I_22266 (I382121,I382079);
nand I_22267 (I381818,I382121,I381940);
nand I_22268 (I382152,I137805,I137805);
and I_22269 (I382169,I382152,I137817);
DFFARX1 I_22270 (I382169,I3563,I381841,I382195,);
nor I_22271 (I382203,I382195,I381867);
DFFARX1 I_22272 (I382203,I3563,I381841,I381806,);
DFFARX1 I_22273 (I382195,I3563,I381841,I381824,);
nor I_22274 (I382248,I137826,I137805);
not I_22275 (I382265,I382248);
nor I_22276 (I381827,I382104,I382265);
nand I_22277 (I381812,I382121,I382265);
nor I_22278 (I381821,I381867,I382248);
DFFARX1 I_22279 (I382248,I3563,I381841,I381830,);
not I_22280 (I382368,I3570);
DFFARX1 I_22281 (I493134,I3563,I382368,I382394,);
nand I_22282 (I382402,I493146,I493125);
and I_22283 (I382419,I382402,I493149);
DFFARX1 I_22284 (I382419,I3563,I382368,I382445,);
nor I_22285 (I382336,I382445,I382394);
not I_22286 (I382467,I382445);
DFFARX1 I_22287 (I493140,I3563,I382368,I382493,);
nand I_22288 (I382501,I382493,I493122);
not I_22289 (I382518,I382501);
DFFARX1 I_22290 (I382518,I3563,I382368,I382544,);
not I_22291 (I382360,I382544);
nor I_22292 (I382566,I382394,I382501);
nor I_22293 (I382342,I382445,I382566);
DFFARX1 I_22294 (I493137,I3563,I382368,I382606,);
DFFARX1 I_22295 (I382606,I3563,I382368,I382623,);
not I_22296 (I382631,I382623);
not I_22297 (I382648,I382606);
nand I_22298 (I382345,I382648,I382467);
nand I_22299 (I382679,I493122,I493128);
and I_22300 (I382696,I382679,I493131);
DFFARX1 I_22301 (I382696,I3563,I382368,I382722,);
nor I_22302 (I382730,I382722,I382394);
DFFARX1 I_22303 (I382730,I3563,I382368,I382333,);
DFFARX1 I_22304 (I382722,I3563,I382368,I382351,);
nor I_22305 (I382775,I493143,I493128);
not I_22306 (I382792,I382775);
nor I_22307 (I382354,I382631,I382792);
nand I_22308 (I382339,I382648,I382792);
nor I_22309 (I382348,I382394,I382775);
DFFARX1 I_22310 (I382775,I3563,I382368,I382357,);
not I_22311 (I382895,I3570);
DFFARX1 I_22312 (I912243,I3563,I382895,I382921,);
nand I_22313 (I382929,I912246,I912240);
and I_22314 (I382946,I382929,I912252);
DFFARX1 I_22315 (I382946,I3563,I382895,I382972,);
nor I_22316 (I382863,I382972,I382921);
not I_22317 (I382994,I382972);
DFFARX1 I_22318 (I912255,I3563,I382895,I383020,);
nand I_22319 (I383028,I383020,I912246);
not I_22320 (I383045,I383028);
DFFARX1 I_22321 (I383045,I3563,I382895,I383071,);
not I_22322 (I382887,I383071);
nor I_22323 (I383093,I382921,I383028);
nor I_22324 (I382869,I382972,I383093);
DFFARX1 I_22325 (I912258,I3563,I382895,I383133,);
DFFARX1 I_22326 (I383133,I3563,I382895,I383150,);
not I_22327 (I383158,I383150);
not I_22328 (I383175,I383133);
nand I_22329 (I382872,I383175,I382994);
nand I_22330 (I383206,I912240,I912249);
and I_22331 (I383223,I383206,I912243);
DFFARX1 I_22332 (I383223,I3563,I382895,I383249,);
nor I_22333 (I383257,I383249,I382921);
DFFARX1 I_22334 (I383257,I3563,I382895,I382860,);
DFFARX1 I_22335 (I383249,I3563,I382895,I382878,);
nor I_22336 (I383302,I912261,I912249);
not I_22337 (I383319,I383302);
nor I_22338 (I382881,I383158,I383319);
nand I_22339 (I382866,I383175,I383319);
nor I_22340 (I382875,I382921,I383302);
DFFARX1 I_22341 (I383302,I3563,I382895,I382884,);
not I_22342 (I383422,I3570);
DFFARX1 I_22343 (I801769,I3563,I383422,I383448,);
nand I_22344 (I383456,I801760,I801775);
and I_22345 (I383473,I383456,I801781);
DFFARX1 I_22346 (I383473,I3563,I383422,I383499,);
nor I_22347 (I383390,I383499,I383448);
not I_22348 (I383521,I383499);
DFFARX1 I_22349 (I801766,I3563,I383422,I383547,);
nand I_22350 (I383555,I383547,I801760);
not I_22351 (I383572,I383555);
DFFARX1 I_22352 (I383572,I3563,I383422,I383598,);
not I_22353 (I383414,I383598);
nor I_22354 (I383620,I383448,I383555);
nor I_22355 (I383396,I383499,I383620);
DFFARX1 I_22356 (I801763,I3563,I383422,I383660,);
DFFARX1 I_22357 (I383660,I3563,I383422,I383677,);
not I_22358 (I383685,I383677);
not I_22359 (I383702,I383660);
nand I_22360 (I383399,I383702,I383521);
nand I_22361 (I383733,I801757,I801772);
and I_22362 (I383750,I383733,I801757);
DFFARX1 I_22363 (I383750,I3563,I383422,I383776,);
nor I_22364 (I383784,I383776,I383448);
DFFARX1 I_22365 (I383784,I3563,I383422,I383387,);
DFFARX1 I_22366 (I383776,I3563,I383422,I383405,);
nor I_22367 (I383829,I801778,I801772);
not I_22368 (I383846,I383829);
nor I_22369 (I383408,I383685,I383846);
nand I_22370 (I383393,I383702,I383846);
nor I_22371 (I383402,I383448,I383829);
DFFARX1 I_22372 (I383829,I3563,I383422,I383411,);
not I_22373 (I383949,I3570);
DFFARX1 I_22374 (I713913,I3563,I383949,I383975,);
nand I_22375 (I383983,I713904,I713919);
and I_22376 (I384000,I383983,I713925);
DFFARX1 I_22377 (I384000,I3563,I383949,I384026,);
nor I_22378 (I383917,I384026,I383975);
not I_22379 (I384048,I384026);
DFFARX1 I_22380 (I713910,I3563,I383949,I384074,);
nand I_22381 (I384082,I384074,I713904);
not I_22382 (I384099,I384082);
DFFARX1 I_22383 (I384099,I3563,I383949,I384125,);
not I_22384 (I383941,I384125);
nor I_22385 (I384147,I383975,I384082);
nor I_22386 (I383923,I384026,I384147);
DFFARX1 I_22387 (I713907,I3563,I383949,I384187,);
DFFARX1 I_22388 (I384187,I3563,I383949,I384204,);
not I_22389 (I384212,I384204);
not I_22390 (I384229,I384187);
nand I_22391 (I383926,I384229,I384048);
nand I_22392 (I384260,I713901,I713916);
and I_22393 (I384277,I384260,I713901);
DFFARX1 I_22394 (I384277,I3563,I383949,I384303,);
nor I_22395 (I384311,I384303,I383975);
DFFARX1 I_22396 (I384311,I3563,I383949,I383914,);
DFFARX1 I_22397 (I384303,I3563,I383949,I383932,);
nor I_22398 (I384356,I713922,I713916);
not I_22399 (I384373,I384356);
nor I_22400 (I383935,I384212,I384373);
nand I_22401 (I383920,I384229,I384373);
nor I_22402 (I383929,I383975,I384356);
DFFARX1 I_22403 (I384356,I3563,I383949,I383938,);
not I_22404 (I384476,I3570);
DFFARX1 I_22405 (I695417,I3563,I384476,I384502,);
nand I_22406 (I384510,I695408,I695423);
and I_22407 (I384527,I384510,I695429);
DFFARX1 I_22408 (I384527,I3563,I384476,I384553,);
nor I_22409 (I384444,I384553,I384502);
not I_22410 (I384575,I384553);
DFFARX1 I_22411 (I695414,I3563,I384476,I384601,);
nand I_22412 (I384609,I384601,I695408);
not I_22413 (I384626,I384609);
DFFARX1 I_22414 (I384626,I3563,I384476,I384652,);
not I_22415 (I384468,I384652);
nor I_22416 (I384674,I384502,I384609);
nor I_22417 (I384450,I384553,I384674);
DFFARX1 I_22418 (I695411,I3563,I384476,I384714,);
DFFARX1 I_22419 (I384714,I3563,I384476,I384731,);
not I_22420 (I384739,I384731);
not I_22421 (I384756,I384714);
nand I_22422 (I384453,I384756,I384575);
nand I_22423 (I384787,I695405,I695420);
and I_22424 (I384804,I384787,I695405);
DFFARX1 I_22425 (I384804,I3563,I384476,I384830,);
nor I_22426 (I384838,I384830,I384502);
DFFARX1 I_22427 (I384838,I3563,I384476,I384441,);
DFFARX1 I_22428 (I384830,I3563,I384476,I384459,);
nor I_22429 (I384883,I695426,I695420);
not I_22430 (I384900,I384883);
nor I_22431 (I384462,I384739,I384900);
nand I_22432 (I384447,I384756,I384900);
nor I_22433 (I384456,I384502,I384883);
DFFARX1 I_22434 (I384883,I3563,I384476,I384465,);
not I_22435 (I385003,I3570);
DFFARX1 I_22436 (I698885,I3563,I385003,I385029,);
nand I_22437 (I385037,I698876,I698891);
and I_22438 (I385054,I385037,I698897);
DFFARX1 I_22439 (I385054,I3563,I385003,I385080,);
nor I_22440 (I384971,I385080,I385029);
not I_22441 (I385102,I385080);
DFFARX1 I_22442 (I698882,I3563,I385003,I385128,);
nand I_22443 (I385136,I385128,I698876);
not I_22444 (I385153,I385136);
DFFARX1 I_22445 (I385153,I3563,I385003,I385179,);
not I_22446 (I384995,I385179);
nor I_22447 (I385201,I385029,I385136);
nor I_22448 (I384977,I385080,I385201);
DFFARX1 I_22449 (I698879,I3563,I385003,I385241,);
DFFARX1 I_22450 (I385241,I3563,I385003,I385258,);
not I_22451 (I385266,I385258);
not I_22452 (I385283,I385241);
nand I_22453 (I384980,I385283,I385102);
nand I_22454 (I385314,I698873,I698888);
and I_22455 (I385331,I385314,I698873);
DFFARX1 I_22456 (I385331,I3563,I385003,I385357,);
nor I_22457 (I385365,I385357,I385029);
DFFARX1 I_22458 (I385365,I3563,I385003,I384968,);
DFFARX1 I_22459 (I385357,I3563,I385003,I384986,);
nor I_22460 (I385410,I698894,I698888);
not I_22461 (I385427,I385410);
nor I_22462 (I384989,I385266,I385427);
nand I_22463 (I384974,I385283,I385427);
nor I_22464 (I384983,I385029,I385410);
DFFARX1 I_22465 (I385410,I3563,I385003,I384992,);
not I_22466 (I385530,I3570);
DFFARX1 I_22467 (I663627,I3563,I385530,I385556,);
nand I_22468 (I385564,I663618,I663633);
and I_22469 (I385581,I385564,I663639);
DFFARX1 I_22470 (I385581,I3563,I385530,I385607,);
nor I_22471 (I385498,I385607,I385556);
not I_22472 (I385629,I385607);
DFFARX1 I_22473 (I663624,I3563,I385530,I385655,);
nand I_22474 (I385663,I385655,I663618);
not I_22475 (I385680,I385663);
DFFARX1 I_22476 (I385680,I3563,I385530,I385706,);
not I_22477 (I385522,I385706);
nor I_22478 (I385728,I385556,I385663);
nor I_22479 (I385504,I385607,I385728);
DFFARX1 I_22480 (I663621,I3563,I385530,I385768,);
DFFARX1 I_22481 (I385768,I3563,I385530,I385785,);
not I_22482 (I385793,I385785);
not I_22483 (I385810,I385768);
nand I_22484 (I385507,I385810,I385629);
nand I_22485 (I385841,I663615,I663630);
and I_22486 (I385858,I385841,I663615);
DFFARX1 I_22487 (I385858,I3563,I385530,I385884,);
nor I_22488 (I385892,I385884,I385556);
DFFARX1 I_22489 (I385892,I3563,I385530,I385495,);
DFFARX1 I_22490 (I385884,I3563,I385530,I385513,);
nor I_22491 (I385937,I663636,I663630);
not I_22492 (I385954,I385937);
nor I_22493 (I385516,I385793,I385954);
nand I_22494 (I385501,I385810,I385954);
nor I_22495 (I385510,I385556,I385937);
DFFARX1 I_22496 (I385937,I3563,I385530,I385519,);
not I_22497 (I386057,I3570);
DFFARX1 I_22498 (I109350,I3563,I386057,I386083,);
nand I_22499 (I386091,I109362,I109371);
and I_22500 (I386108,I386091,I109350);
DFFARX1 I_22501 (I386108,I3563,I386057,I386134,);
nor I_22502 (I386025,I386134,I386083);
not I_22503 (I386156,I386134);
DFFARX1 I_22504 (I109365,I3563,I386057,I386182,);
nand I_22505 (I386190,I386182,I109353);
not I_22506 (I386207,I386190);
DFFARX1 I_22507 (I386207,I3563,I386057,I386233,);
not I_22508 (I386049,I386233);
nor I_22509 (I386255,I386083,I386190);
nor I_22510 (I386031,I386134,I386255);
DFFARX1 I_22511 (I109356,I3563,I386057,I386295,);
DFFARX1 I_22512 (I386295,I3563,I386057,I386312,);
not I_22513 (I386320,I386312);
not I_22514 (I386337,I386295);
nand I_22515 (I386034,I386337,I386156);
nand I_22516 (I386368,I109347,I109347);
and I_22517 (I386385,I386368,I109359);
DFFARX1 I_22518 (I386385,I3563,I386057,I386411,);
nor I_22519 (I386419,I386411,I386083);
DFFARX1 I_22520 (I386419,I3563,I386057,I386022,);
DFFARX1 I_22521 (I386411,I3563,I386057,I386040,);
nor I_22522 (I386464,I109368,I109347);
not I_22523 (I386481,I386464);
nor I_22524 (I386043,I386320,I386481);
nand I_22525 (I386028,I386337,I386481);
nor I_22526 (I386037,I386083,I386464);
DFFARX1 I_22527 (I386464,I3563,I386057,I386046,);
not I_22528 (I386584,I3570);
DFFARX1 I_22529 (I892217,I3563,I386584,I386610,);
nand I_22530 (I386618,I892220,I892214);
and I_22531 (I386635,I386618,I892226);
DFFARX1 I_22532 (I386635,I3563,I386584,I386661,);
nor I_22533 (I386552,I386661,I386610);
not I_22534 (I386683,I386661);
DFFARX1 I_22535 (I892229,I3563,I386584,I386709,);
nand I_22536 (I386717,I386709,I892220);
not I_22537 (I386734,I386717);
DFFARX1 I_22538 (I386734,I3563,I386584,I386760,);
not I_22539 (I386576,I386760);
nor I_22540 (I386782,I386610,I386717);
nor I_22541 (I386558,I386661,I386782);
DFFARX1 I_22542 (I892232,I3563,I386584,I386822,);
DFFARX1 I_22543 (I386822,I3563,I386584,I386839,);
not I_22544 (I386847,I386839);
not I_22545 (I386864,I386822);
nand I_22546 (I386561,I386864,I386683);
nand I_22547 (I386895,I892214,I892223);
and I_22548 (I386912,I386895,I892217);
DFFARX1 I_22549 (I386912,I3563,I386584,I386938,);
nor I_22550 (I386946,I386938,I386610);
DFFARX1 I_22551 (I386946,I3563,I386584,I386549,);
DFFARX1 I_22552 (I386938,I3563,I386584,I386567,);
nor I_22553 (I386991,I892235,I892223);
not I_22554 (I387008,I386991);
nor I_22555 (I386570,I386847,I387008);
nand I_22556 (I386555,I386864,I387008);
nor I_22557 (I386564,I386610,I386991);
DFFARX1 I_22558 (I386991,I3563,I386584,I386573,);
not I_22559 (I387111,I3570);
DFFARX1 I_22560 (I216668,I3563,I387111,I387137,);
nand I_22561 (I387145,I216668,I216674);
and I_22562 (I387162,I387145,I216692);
DFFARX1 I_22563 (I387162,I3563,I387111,I387188,);
nor I_22564 (I387079,I387188,I387137);
not I_22565 (I387210,I387188);
DFFARX1 I_22566 (I216680,I3563,I387111,I387236,);
nand I_22567 (I387244,I387236,I216677);
not I_22568 (I387261,I387244);
DFFARX1 I_22569 (I387261,I3563,I387111,I387287,);
not I_22570 (I387103,I387287);
nor I_22571 (I387309,I387137,I387244);
nor I_22572 (I387085,I387188,I387309);
DFFARX1 I_22573 (I216686,I3563,I387111,I387349,);
DFFARX1 I_22574 (I387349,I3563,I387111,I387366,);
not I_22575 (I387374,I387366);
not I_22576 (I387391,I387349);
nand I_22577 (I387088,I387391,I387210);
nand I_22578 (I387422,I216671,I216671);
and I_22579 (I387439,I387422,I216683);
DFFARX1 I_22580 (I387439,I3563,I387111,I387465,);
nor I_22581 (I387473,I387465,I387137);
DFFARX1 I_22582 (I387473,I3563,I387111,I387076,);
DFFARX1 I_22583 (I387465,I3563,I387111,I387094,);
nor I_22584 (I387518,I216689,I216671);
not I_22585 (I387535,I387518);
nor I_22586 (I387097,I387374,I387535);
nand I_22587 (I387082,I387391,I387535);
nor I_22588 (I387091,I387137,I387518);
DFFARX1 I_22589 (I387518,I3563,I387111,I387100,);
not I_22590 (I387638,I3570);
DFFARX1 I_22591 (I759575,I3563,I387638,I387664,);
nand I_22592 (I387672,I759566,I759581);
and I_22593 (I387689,I387672,I759587);
DFFARX1 I_22594 (I387689,I3563,I387638,I387715,);
nor I_22595 (I387606,I387715,I387664);
not I_22596 (I387737,I387715);
DFFARX1 I_22597 (I759572,I3563,I387638,I387763,);
nand I_22598 (I387771,I387763,I759566);
not I_22599 (I387788,I387771);
DFFARX1 I_22600 (I387788,I3563,I387638,I387814,);
not I_22601 (I387630,I387814);
nor I_22602 (I387836,I387664,I387771);
nor I_22603 (I387612,I387715,I387836);
DFFARX1 I_22604 (I759569,I3563,I387638,I387876,);
DFFARX1 I_22605 (I387876,I3563,I387638,I387893,);
not I_22606 (I387901,I387893);
not I_22607 (I387918,I387876);
nand I_22608 (I387615,I387918,I387737);
nand I_22609 (I387949,I759563,I759578);
and I_22610 (I387966,I387949,I759563);
DFFARX1 I_22611 (I387966,I3563,I387638,I387992,);
nor I_22612 (I388000,I387992,I387664);
DFFARX1 I_22613 (I388000,I3563,I387638,I387603,);
DFFARX1 I_22614 (I387992,I3563,I387638,I387621,);
nor I_22615 (I388045,I759584,I759578);
not I_22616 (I388062,I388045);
nor I_22617 (I387624,I387901,I388062);
nand I_22618 (I387609,I387918,I388062);
nor I_22619 (I387618,I387664,I388045);
DFFARX1 I_22620 (I388045,I3563,I387638,I387627,);
not I_22621 (I388165,I3570);
DFFARX1 I_22622 (I782117,I3563,I388165,I388191,);
nand I_22623 (I388199,I782108,I782123);
and I_22624 (I388216,I388199,I782129);
DFFARX1 I_22625 (I388216,I3563,I388165,I388242,);
nor I_22626 (I388133,I388242,I388191);
not I_22627 (I388264,I388242);
DFFARX1 I_22628 (I782114,I3563,I388165,I388290,);
nand I_22629 (I388298,I388290,I782108);
not I_22630 (I388315,I388298);
DFFARX1 I_22631 (I388315,I3563,I388165,I388341,);
not I_22632 (I388157,I388341);
nor I_22633 (I388363,I388191,I388298);
nor I_22634 (I388139,I388242,I388363);
DFFARX1 I_22635 (I782111,I3563,I388165,I388403,);
DFFARX1 I_22636 (I388403,I3563,I388165,I388420,);
not I_22637 (I388428,I388420);
not I_22638 (I388445,I388403);
nand I_22639 (I388142,I388445,I388264);
nand I_22640 (I388476,I782105,I782120);
and I_22641 (I388493,I388476,I782105);
DFFARX1 I_22642 (I388493,I3563,I388165,I388519,);
nor I_22643 (I388527,I388519,I388191);
DFFARX1 I_22644 (I388527,I3563,I388165,I388130,);
DFFARX1 I_22645 (I388519,I3563,I388165,I388148,);
nor I_22646 (I388572,I782126,I782120);
not I_22647 (I388589,I388572);
nor I_22648 (I388151,I388428,I388589);
nand I_22649 (I388136,I388445,I388589);
nor I_22650 (I388145,I388191,I388572);
DFFARX1 I_22651 (I388572,I3563,I388165,I388154,);
not I_22652 (I388692,I3570);
DFFARX1 I_22653 (I1267099,I3563,I388692,I388718,);
nand I_22654 (I388726,I1267081,I1267105);
and I_22655 (I388743,I388726,I1267096);
DFFARX1 I_22656 (I388743,I3563,I388692,I388769,);
nor I_22657 (I388660,I388769,I388718);
not I_22658 (I388791,I388769);
DFFARX1 I_22659 (I1267102,I3563,I388692,I388817,);
nand I_22660 (I388825,I388817,I1267090);
not I_22661 (I388842,I388825);
DFFARX1 I_22662 (I388842,I3563,I388692,I388868,);
not I_22663 (I388684,I388868);
nor I_22664 (I388890,I388718,I388825);
nor I_22665 (I388666,I388769,I388890);
DFFARX1 I_22666 (I1267081,I3563,I388692,I388930,);
DFFARX1 I_22667 (I388930,I3563,I388692,I388947,);
not I_22668 (I388955,I388947);
not I_22669 (I388972,I388930);
nand I_22670 (I388669,I388972,I388791);
nand I_22671 (I389003,I1267087,I1267084);
and I_22672 (I389020,I389003,I1267093);
DFFARX1 I_22673 (I389020,I3563,I388692,I389046,);
nor I_22674 (I389054,I389046,I388718);
DFFARX1 I_22675 (I389054,I3563,I388692,I388657,);
DFFARX1 I_22676 (I389046,I3563,I388692,I388675,);
nor I_22677 (I389099,I1267084,I1267084);
not I_22678 (I389116,I389099);
nor I_22679 (I388678,I388955,I389116);
nand I_22680 (I388663,I388972,I389116);
nor I_22681 (I388672,I388718,I389099);
DFFARX1 I_22682 (I389099,I3563,I388692,I388681,);
not I_22683 (I389219,I3570);
DFFARX1 I_22684 (I852692,I3563,I389219,I389245,);
nand I_22685 (I389253,I852695,I852689);
and I_22686 (I389270,I389253,I852701);
DFFARX1 I_22687 (I389270,I3563,I389219,I389296,);
nor I_22688 (I389187,I389296,I389245);
not I_22689 (I389318,I389296);
DFFARX1 I_22690 (I852704,I3563,I389219,I389344,);
nand I_22691 (I389352,I389344,I852695);
not I_22692 (I389369,I389352);
DFFARX1 I_22693 (I389369,I3563,I389219,I389395,);
not I_22694 (I389211,I389395);
nor I_22695 (I389417,I389245,I389352);
nor I_22696 (I389193,I389296,I389417);
DFFARX1 I_22697 (I852707,I3563,I389219,I389457,);
DFFARX1 I_22698 (I389457,I3563,I389219,I389474,);
not I_22699 (I389482,I389474);
not I_22700 (I389499,I389457);
nand I_22701 (I389196,I389499,I389318);
nand I_22702 (I389530,I852689,I852698);
and I_22703 (I389547,I389530,I852692);
DFFARX1 I_22704 (I389547,I3563,I389219,I389573,);
nor I_22705 (I389581,I389573,I389245);
DFFARX1 I_22706 (I389581,I3563,I389219,I389184,);
DFFARX1 I_22707 (I389573,I3563,I389219,I389202,);
nor I_22708 (I389626,I852710,I852698);
not I_22709 (I389643,I389626);
nor I_22710 (I389205,I389482,I389643);
nand I_22711 (I389190,I389499,I389643);
nor I_22712 (I389199,I389245,I389626);
DFFARX1 I_22713 (I389626,I3563,I389219,I389208,);
not I_22714 (I389746,I3570);
DFFARX1 I_22715 (I204768,I3563,I389746,I389772,);
nand I_22716 (I389780,I204768,I204774);
and I_22717 (I389797,I389780,I204792);
DFFARX1 I_22718 (I389797,I3563,I389746,I389823,);
nor I_22719 (I389714,I389823,I389772);
not I_22720 (I389845,I389823);
DFFARX1 I_22721 (I204780,I3563,I389746,I389871,);
nand I_22722 (I389879,I389871,I204777);
not I_22723 (I389896,I389879);
DFFARX1 I_22724 (I389896,I3563,I389746,I389922,);
not I_22725 (I389738,I389922);
nor I_22726 (I389944,I389772,I389879);
nor I_22727 (I389720,I389823,I389944);
DFFARX1 I_22728 (I204786,I3563,I389746,I389984,);
DFFARX1 I_22729 (I389984,I3563,I389746,I390001,);
not I_22730 (I390009,I390001);
not I_22731 (I390026,I389984);
nand I_22732 (I389723,I390026,I389845);
nand I_22733 (I390057,I204771,I204771);
and I_22734 (I390074,I390057,I204783);
DFFARX1 I_22735 (I390074,I3563,I389746,I390100,);
nor I_22736 (I390108,I390100,I389772);
DFFARX1 I_22737 (I390108,I3563,I389746,I389711,);
DFFARX1 I_22738 (I390100,I3563,I389746,I389729,);
nor I_22739 (I390153,I204789,I204771);
not I_22740 (I390170,I390153);
nor I_22741 (I389732,I390009,I390170);
nand I_22742 (I389717,I390026,I390170);
nor I_22743 (I389726,I389772,I390153);
DFFARX1 I_22744 (I390153,I3563,I389746,I389735,);
not I_22745 (I390273,I3570);
DFFARX1 I_22746 (I767667,I3563,I390273,I390299,);
nand I_22747 (I390307,I767658,I767673);
and I_22748 (I390324,I390307,I767679);
DFFARX1 I_22749 (I390324,I3563,I390273,I390350,);
nor I_22750 (I390241,I390350,I390299);
not I_22751 (I390372,I390350);
DFFARX1 I_22752 (I767664,I3563,I390273,I390398,);
nand I_22753 (I390406,I390398,I767658);
not I_22754 (I390423,I390406);
DFFARX1 I_22755 (I390423,I3563,I390273,I390449,);
not I_22756 (I390265,I390449);
nor I_22757 (I390471,I390299,I390406);
nor I_22758 (I390247,I390350,I390471);
DFFARX1 I_22759 (I767661,I3563,I390273,I390511,);
DFFARX1 I_22760 (I390511,I3563,I390273,I390528,);
not I_22761 (I390536,I390528);
not I_22762 (I390553,I390511);
nand I_22763 (I390250,I390553,I390372);
nand I_22764 (I390584,I767655,I767670);
and I_22765 (I390601,I390584,I767655);
DFFARX1 I_22766 (I390601,I3563,I390273,I390627,);
nor I_22767 (I390635,I390627,I390299);
DFFARX1 I_22768 (I390635,I3563,I390273,I390238,);
DFFARX1 I_22769 (I390627,I3563,I390273,I390256,);
nor I_22770 (I390680,I767676,I767670);
not I_22771 (I390697,I390680);
nor I_22772 (I390259,I390536,I390697);
nand I_22773 (I390244,I390553,I390697);
nor I_22774 (I390253,I390299,I390680);
DFFARX1 I_22775 (I390680,I3563,I390273,I390262,);
not I_22776 (I390800,I3570);
DFFARX1 I_22777 (I268433,I3563,I390800,I390826,);
nand I_22778 (I390834,I268433,I268439);
and I_22779 (I390851,I390834,I268457);
DFFARX1 I_22780 (I390851,I3563,I390800,I390877,);
nor I_22781 (I390768,I390877,I390826);
not I_22782 (I390899,I390877);
DFFARX1 I_22783 (I268445,I3563,I390800,I390925,);
nand I_22784 (I390933,I390925,I268442);
not I_22785 (I390950,I390933);
DFFARX1 I_22786 (I390950,I3563,I390800,I390976,);
not I_22787 (I390792,I390976);
nor I_22788 (I390998,I390826,I390933);
nor I_22789 (I390774,I390877,I390998);
DFFARX1 I_22790 (I268451,I3563,I390800,I391038,);
DFFARX1 I_22791 (I391038,I3563,I390800,I391055,);
not I_22792 (I391063,I391055);
not I_22793 (I391080,I391038);
nand I_22794 (I390777,I391080,I390899);
nand I_22795 (I391111,I268436,I268436);
and I_22796 (I391128,I391111,I268448);
DFFARX1 I_22797 (I391128,I3563,I390800,I391154,);
nor I_22798 (I391162,I391154,I390826);
DFFARX1 I_22799 (I391162,I3563,I390800,I390765,);
DFFARX1 I_22800 (I391154,I3563,I390800,I390783,);
nor I_22801 (I391207,I268454,I268436);
not I_22802 (I391224,I391207);
nor I_22803 (I390786,I391063,I391224);
nand I_22804 (I390771,I391080,I391224);
nor I_22805 (I390780,I390826,I391207);
DFFARX1 I_22806 (I391207,I3563,I390800,I390789,);
not I_22807 (I391327,I3570);
DFFARX1 I_22808 (I107242,I3563,I391327,I391353,);
nand I_22809 (I391361,I107254,I107263);
and I_22810 (I391378,I391361,I107242);
DFFARX1 I_22811 (I391378,I3563,I391327,I391404,);
nor I_22812 (I391295,I391404,I391353);
not I_22813 (I391426,I391404);
DFFARX1 I_22814 (I107257,I3563,I391327,I391452,);
nand I_22815 (I391460,I391452,I107245);
not I_22816 (I391477,I391460);
DFFARX1 I_22817 (I391477,I3563,I391327,I391503,);
not I_22818 (I391319,I391503);
nor I_22819 (I391525,I391353,I391460);
nor I_22820 (I391301,I391404,I391525);
DFFARX1 I_22821 (I107248,I3563,I391327,I391565,);
DFFARX1 I_22822 (I391565,I3563,I391327,I391582,);
not I_22823 (I391590,I391582);
not I_22824 (I391607,I391565);
nand I_22825 (I391304,I391607,I391426);
nand I_22826 (I391638,I107239,I107239);
and I_22827 (I391655,I391638,I107251);
DFFARX1 I_22828 (I391655,I3563,I391327,I391681,);
nor I_22829 (I391689,I391681,I391353);
DFFARX1 I_22830 (I391689,I3563,I391327,I391292,);
DFFARX1 I_22831 (I391681,I3563,I391327,I391310,);
nor I_22832 (I391734,I107260,I107239);
not I_22833 (I391751,I391734);
nor I_22834 (I391313,I391590,I391751);
nand I_22835 (I391298,I391607,I391751);
nor I_22836 (I391307,I391353,I391734);
DFFARX1 I_22837 (I391734,I3563,I391327,I391316,);
not I_22838 (I391854,I3570);
DFFARX1 I_22839 (I1062370,I3563,I391854,I391880,);
nand I_22840 (I391888,I1062367,I1062370);
and I_22841 (I391905,I391888,I1062379);
DFFARX1 I_22842 (I391905,I3563,I391854,I391931,);
nor I_22843 (I391822,I391931,I391880);
not I_22844 (I391953,I391931);
DFFARX1 I_22845 (I1062367,I3563,I391854,I391979,);
nand I_22846 (I391987,I391979,I1062385);
not I_22847 (I392004,I391987);
DFFARX1 I_22848 (I392004,I3563,I391854,I392030,);
not I_22849 (I391846,I392030);
nor I_22850 (I392052,I391880,I391987);
nor I_22851 (I391828,I391931,I392052);
DFFARX1 I_22852 (I1062373,I3563,I391854,I392092,);
DFFARX1 I_22853 (I392092,I3563,I391854,I392109,);
not I_22854 (I392117,I392109);
not I_22855 (I392134,I392092);
nand I_22856 (I391831,I392134,I391953);
nand I_22857 (I392165,I1062382,I1062388);
and I_22858 (I392182,I392165,I1062373);
DFFARX1 I_22859 (I392182,I3563,I391854,I392208,);
nor I_22860 (I392216,I392208,I391880);
DFFARX1 I_22861 (I392216,I3563,I391854,I391819,);
DFFARX1 I_22862 (I392208,I3563,I391854,I391837,);
nor I_22863 (I392261,I1062376,I1062388);
not I_22864 (I392278,I392261);
nor I_22865 (I391840,I392117,I392278);
nand I_22866 (I391825,I392134,I392278);
nor I_22867 (I391834,I391880,I392261);
DFFARX1 I_22868 (I392261,I3563,I391854,I391843,);
not I_22869 (I392381,I3570);
DFFARX1 I_22870 (I793099,I3563,I392381,I392407,);
nand I_22871 (I392415,I793090,I793105);
and I_22872 (I392432,I392415,I793111);
DFFARX1 I_22873 (I392432,I3563,I392381,I392458,);
nor I_22874 (I392349,I392458,I392407);
not I_22875 (I392480,I392458);
DFFARX1 I_22876 (I793096,I3563,I392381,I392506,);
nand I_22877 (I392514,I392506,I793090);
not I_22878 (I392531,I392514);
DFFARX1 I_22879 (I392531,I3563,I392381,I392557,);
not I_22880 (I392373,I392557);
nor I_22881 (I392579,I392407,I392514);
nor I_22882 (I392355,I392458,I392579);
DFFARX1 I_22883 (I793093,I3563,I392381,I392619,);
DFFARX1 I_22884 (I392619,I3563,I392381,I392636,);
not I_22885 (I392644,I392636);
not I_22886 (I392661,I392619);
nand I_22887 (I392358,I392661,I392480);
nand I_22888 (I392692,I793087,I793102);
and I_22889 (I392709,I392692,I793087);
DFFARX1 I_22890 (I392709,I3563,I392381,I392735,);
nor I_22891 (I392743,I392735,I392407);
DFFARX1 I_22892 (I392743,I3563,I392381,I392346,);
DFFARX1 I_22893 (I392735,I3563,I392381,I392364,);
nor I_22894 (I392788,I793108,I793102);
not I_22895 (I392805,I392788);
nor I_22896 (I392367,I392644,I392805);
nand I_22897 (I392352,I392661,I392805);
nor I_22898 (I392361,I392407,I392788);
DFFARX1 I_22899 (I392788,I3563,I392381,I392370,);
not I_22900 (I392908,I3570);
DFFARX1 I_22901 (I1186365,I3563,I392908,I392934,);
nand I_22902 (I392942,I1186380,I1186365);
and I_22903 (I392959,I392942,I1186383);
DFFARX1 I_22904 (I392959,I3563,I392908,I392985,);
nor I_22905 (I392876,I392985,I392934);
not I_22906 (I393007,I392985);
DFFARX1 I_22907 (I1186389,I3563,I392908,I393033,);
nand I_22908 (I393041,I393033,I1186371);
not I_22909 (I393058,I393041);
DFFARX1 I_22910 (I393058,I3563,I392908,I393084,);
not I_22911 (I392900,I393084);
nor I_22912 (I393106,I392934,I393041);
nor I_22913 (I392882,I392985,I393106);
DFFARX1 I_22914 (I1186368,I3563,I392908,I393146,);
DFFARX1 I_22915 (I393146,I3563,I392908,I393163,);
not I_22916 (I393171,I393163);
not I_22917 (I393188,I393146);
nand I_22918 (I392885,I393188,I393007);
nand I_22919 (I393219,I1186368,I1186374);
and I_22920 (I393236,I393219,I1186386);
DFFARX1 I_22921 (I393236,I3563,I392908,I393262,);
nor I_22922 (I393270,I393262,I392934);
DFFARX1 I_22923 (I393270,I3563,I392908,I392873,);
DFFARX1 I_22924 (I393262,I3563,I392908,I392891,);
nor I_22925 (I393315,I1186377,I1186374);
not I_22926 (I393332,I393315);
nor I_22927 (I392894,I393171,I393332);
nand I_22928 (I392879,I393188,I393332);
nor I_22929 (I392888,I392934,I393315);
DFFARX1 I_22930 (I393315,I3563,I392908,I392897,);
not I_22931 (I393435,I3570);
DFFARX1 I_22932 (I511086,I3563,I393435,I393461,);
nand I_22933 (I393469,I511098,I511077);
and I_22934 (I393486,I393469,I511101);
DFFARX1 I_22935 (I393486,I3563,I393435,I393512,);
nor I_22936 (I393403,I393512,I393461);
not I_22937 (I393534,I393512);
DFFARX1 I_22938 (I511092,I3563,I393435,I393560,);
nand I_22939 (I393568,I393560,I511074);
not I_22940 (I393585,I393568);
DFFARX1 I_22941 (I393585,I3563,I393435,I393611,);
not I_22942 (I393427,I393611);
nor I_22943 (I393633,I393461,I393568);
nor I_22944 (I393409,I393512,I393633);
DFFARX1 I_22945 (I511089,I3563,I393435,I393673,);
DFFARX1 I_22946 (I393673,I3563,I393435,I393690,);
not I_22947 (I393698,I393690);
not I_22948 (I393715,I393673);
nand I_22949 (I393412,I393715,I393534);
nand I_22950 (I393746,I511074,I511080);
and I_22951 (I393763,I393746,I511083);
DFFARX1 I_22952 (I393763,I3563,I393435,I393789,);
nor I_22953 (I393797,I393789,I393461);
DFFARX1 I_22954 (I393797,I3563,I393435,I393400,);
DFFARX1 I_22955 (I393789,I3563,I393435,I393418,);
nor I_22956 (I393842,I511095,I511080);
not I_22957 (I393859,I393842);
nor I_22958 (I393421,I393698,I393859);
nand I_22959 (I393406,I393715,I393859);
nor I_22960 (I393415,I393461,I393842);
DFFARX1 I_22961 (I393842,I3563,I393435,I393424,);
not I_22962 (I393962,I3570);
DFFARX1 I_22963 (I853219,I3563,I393962,I393988,);
nand I_22964 (I393996,I853222,I853216);
and I_22965 (I394013,I393996,I853228);
DFFARX1 I_22966 (I394013,I3563,I393962,I394039,);
nor I_22967 (I393930,I394039,I393988);
not I_22968 (I394061,I394039);
DFFARX1 I_22969 (I853231,I3563,I393962,I394087,);
nand I_22970 (I394095,I394087,I853222);
not I_22971 (I394112,I394095);
DFFARX1 I_22972 (I394112,I3563,I393962,I394138,);
not I_22973 (I393954,I394138);
nor I_22974 (I394160,I393988,I394095);
nor I_22975 (I393936,I394039,I394160);
DFFARX1 I_22976 (I853234,I3563,I393962,I394200,);
DFFARX1 I_22977 (I394200,I3563,I393962,I394217,);
not I_22978 (I394225,I394217);
not I_22979 (I394242,I394200);
nand I_22980 (I393939,I394242,I394061);
nand I_22981 (I394273,I853216,I853225);
and I_22982 (I394290,I394273,I853219);
DFFARX1 I_22983 (I394290,I3563,I393962,I394316,);
nor I_22984 (I394324,I394316,I393988);
DFFARX1 I_22985 (I394324,I3563,I393962,I393927,);
DFFARX1 I_22986 (I394316,I3563,I393962,I393945,);
nor I_22987 (I394369,I853237,I853225);
not I_22988 (I394386,I394369);
nor I_22989 (I393948,I394225,I394386);
nand I_22990 (I393933,I394242,I394386);
nor I_22991 (I393942,I393988,I394369);
DFFARX1 I_22992 (I394369,I3563,I393962,I393951,);
not I_22993 (I394489,I3570);
DFFARX1 I_22994 (I1248059,I3563,I394489,I394515,);
nand I_22995 (I394523,I1248041,I1248065);
and I_22996 (I394540,I394523,I1248056);
DFFARX1 I_22997 (I394540,I3563,I394489,I394566,);
nor I_22998 (I394457,I394566,I394515);
not I_22999 (I394588,I394566);
DFFARX1 I_23000 (I1248062,I3563,I394489,I394614,);
nand I_23001 (I394622,I394614,I1248050);
not I_23002 (I394639,I394622);
DFFARX1 I_23003 (I394639,I3563,I394489,I394665,);
not I_23004 (I394481,I394665);
nor I_23005 (I394687,I394515,I394622);
nor I_23006 (I394463,I394566,I394687);
DFFARX1 I_23007 (I1248041,I3563,I394489,I394727,);
DFFARX1 I_23008 (I394727,I3563,I394489,I394744,);
not I_23009 (I394752,I394744);
not I_23010 (I394769,I394727);
nand I_23011 (I394466,I394769,I394588);
nand I_23012 (I394800,I1248047,I1248044);
and I_23013 (I394817,I394800,I1248053);
DFFARX1 I_23014 (I394817,I3563,I394489,I394843,);
nor I_23015 (I394851,I394843,I394515);
DFFARX1 I_23016 (I394851,I3563,I394489,I394454,);
DFFARX1 I_23017 (I394843,I3563,I394489,I394472,);
nor I_23018 (I394896,I1248044,I1248044);
not I_23019 (I394913,I394896);
nor I_23020 (I394475,I394752,I394913);
nand I_23021 (I394460,I394769,I394913);
nor I_23022 (I394469,I394515,I394896);
DFFARX1 I_23023 (I394896,I3563,I394489,I394478,);
not I_23024 (I395016,I3570);
DFFARX1 I_23025 (I1136079,I3563,I395016,I395042,);
nand I_23026 (I395050,I1136094,I1136079);
and I_23027 (I395067,I395050,I1136097);
DFFARX1 I_23028 (I395067,I3563,I395016,I395093,);
nor I_23029 (I394984,I395093,I395042);
not I_23030 (I395115,I395093);
DFFARX1 I_23031 (I1136103,I3563,I395016,I395141,);
nand I_23032 (I395149,I395141,I1136085);
not I_23033 (I395166,I395149);
DFFARX1 I_23034 (I395166,I3563,I395016,I395192,);
not I_23035 (I395008,I395192);
nor I_23036 (I395214,I395042,I395149);
nor I_23037 (I394990,I395093,I395214);
DFFARX1 I_23038 (I1136082,I3563,I395016,I395254,);
DFFARX1 I_23039 (I395254,I3563,I395016,I395271,);
not I_23040 (I395279,I395271);
not I_23041 (I395296,I395254);
nand I_23042 (I394993,I395296,I395115);
nand I_23043 (I395327,I1136082,I1136088);
and I_23044 (I395344,I395327,I1136100);
DFFARX1 I_23045 (I395344,I3563,I395016,I395370,);
nor I_23046 (I395378,I395370,I395042);
DFFARX1 I_23047 (I395378,I3563,I395016,I394981,);
DFFARX1 I_23048 (I395370,I3563,I395016,I394999,);
nor I_23049 (I395423,I1136091,I1136088);
not I_23050 (I395440,I395423);
nor I_23051 (I395002,I395279,I395440);
nand I_23052 (I394987,I395296,I395440);
nor I_23053 (I394996,I395042,I395423);
DFFARX1 I_23054 (I395423,I3563,I395016,I395005,);
not I_23055 (I395543,I3570);
DFFARX1 I_23056 (I126214,I3563,I395543,I395569,);
nand I_23057 (I395577,I126226,I126235);
and I_23058 (I395594,I395577,I126214);
DFFARX1 I_23059 (I395594,I3563,I395543,I395620,);
nor I_23060 (I395511,I395620,I395569);
not I_23061 (I395642,I395620);
DFFARX1 I_23062 (I126229,I3563,I395543,I395668,);
nand I_23063 (I395676,I395668,I126217);
not I_23064 (I395693,I395676);
DFFARX1 I_23065 (I395693,I3563,I395543,I395719,);
not I_23066 (I395535,I395719);
nor I_23067 (I395741,I395569,I395676);
nor I_23068 (I395517,I395620,I395741);
DFFARX1 I_23069 (I126220,I3563,I395543,I395781,);
DFFARX1 I_23070 (I395781,I3563,I395543,I395798,);
not I_23071 (I395806,I395798);
not I_23072 (I395823,I395781);
nand I_23073 (I395520,I395823,I395642);
nand I_23074 (I395854,I126211,I126211);
and I_23075 (I395871,I395854,I126223);
DFFARX1 I_23076 (I395871,I3563,I395543,I395897,);
nor I_23077 (I395905,I395897,I395569);
DFFARX1 I_23078 (I395905,I3563,I395543,I395508,);
DFFARX1 I_23079 (I395897,I3563,I395543,I395526,);
nor I_23080 (I395950,I126232,I126211);
not I_23081 (I395967,I395950);
nor I_23082 (I395529,I395806,I395967);
nand I_23083 (I395514,I395823,I395967);
nor I_23084 (I395523,I395569,I395950);
DFFARX1 I_23085 (I395950,I3563,I395543,I395532,);
not I_23086 (I396070,I3570);
DFFARX1 I_23087 (I1093885,I3563,I396070,I396096,);
nand I_23088 (I396104,I1093900,I1093885);
and I_23089 (I396121,I396104,I1093903);
DFFARX1 I_23090 (I396121,I3563,I396070,I396147,);
nor I_23091 (I396038,I396147,I396096);
not I_23092 (I396169,I396147);
DFFARX1 I_23093 (I1093909,I3563,I396070,I396195,);
nand I_23094 (I396203,I396195,I1093891);
not I_23095 (I396220,I396203);
DFFARX1 I_23096 (I396220,I3563,I396070,I396246,);
not I_23097 (I396062,I396246);
nor I_23098 (I396268,I396096,I396203);
nor I_23099 (I396044,I396147,I396268);
DFFARX1 I_23100 (I1093888,I3563,I396070,I396308,);
DFFARX1 I_23101 (I396308,I3563,I396070,I396325,);
not I_23102 (I396333,I396325);
not I_23103 (I396350,I396308);
nand I_23104 (I396047,I396350,I396169);
nand I_23105 (I396381,I1093888,I1093894);
and I_23106 (I396398,I396381,I1093906);
DFFARX1 I_23107 (I396398,I3563,I396070,I396424,);
nor I_23108 (I396432,I396424,I396096);
DFFARX1 I_23109 (I396432,I3563,I396070,I396035,);
DFFARX1 I_23110 (I396424,I3563,I396070,I396053,);
nor I_23111 (I396477,I1093897,I1093894);
not I_23112 (I396494,I396477);
nor I_23113 (I396056,I396333,I396494);
nand I_23114 (I396041,I396350,I396494);
nor I_23115 (I396050,I396096,I396477);
DFFARX1 I_23116 (I396477,I3563,I396070,I396059,);
not I_23117 (I396597,I3570);
DFFARX1 I_23118 (I895906,I3563,I396597,I396623,);
nand I_23119 (I396631,I895909,I895903);
and I_23120 (I396648,I396631,I895915);
DFFARX1 I_23121 (I396648,I3563,I396597,I396674,);
nor I_23122 (I396565,I396674,I396623);
not I_23123 (I396696,I396674);
DFFARX1 I_23124 (I895918,I3563,I396597,I396722,);
nand I_23125 (I396730,I396722,I895909);
not I_23126 (I396747,I396730);
DFFARX1 I_23127 (I396747,I3563,I396597,I396773,);
not I_23128 (I396589,I396773);
nor I_23129 (I396795,I396623,I396730);
nor I_23130 (I396571,I396674,I396795);
DFFARX1 I_23131 (I895921,I3563,I396597,I396835,);
DFFARX1 I_23132 (I396835,I3563,I396597,I396852,);
not I_23133 (I396860,I396852);
not I_23134 (I396877,I396835);
nand I_23135 (I396574,I396877,I396696);
nand I_23136 (I396908,I895903,I895912);
and I_23137 (I396925,I396908,I895906);
DFFARX1 I_23138 (I396925,I3563,I396597,I396951,);
nor I_23139 (I396959,I396951,I396623);
DFFARX1 I_23140 (I396959,I3563,I396597,I396562,);
DFFARX1 I_23141 (I396951,I3563,I396597,I396580,);
nor I_23142 (I397004,I895924,I895912);
not I_23143 (I397021,I397004);
nor I_23144 (I396583,I396860,I397021);
nand I_23145 (I396568,I396877,I397021);
nor I_23146 (I396577,I396623,I397004);
DFFARX1 I_23147 (I397004,I3563,I396597,I396586,);
not I_23148 (I397124,I3570);
DFFARX1 I_23149 (I814221,I3563,I397124,I397150,);
nand I_23150 (I397158,I814224,I814218);
and I_23151 (I397175,I397158,I814230);
DFFARX1 I_23152 (I397175,I3563,I397124,I397201,);
nor I_23153 (I397092,I397201,I397150);
not I_23154 (I397223,I397201);
DFFARX1 I_23155 (I814233,I3563,I397124,I397249,);
nand I_23156 (I397257,I397249,I814224);
not I_23157 (I397274,I397257);
DFFARX1 I_23158 (I397274,I3563,I397124,I397300,);
not I_23159 (I397116,I397300);
nor I_23160 (I397322,I397150,I397257);
nor I_23161 (I397098,I397201,I397322);
DFFARX1 I_23162 (I814236,I3563,I397124,I397362,);
DFFARX1 I_23163 (I397362,I3563,I397124,I397379,);
not I_23164 (I397387,I397379);
not I_23165 (I397404,I397362);
nand I_23166 (I397101,I397404,I397223);
nand I_23167 (I397435,I814218,I814227);
and I_23168 (I397452,I397435,I814221);
DFFARX1 I_23169 (I397452,I3563,I397124,I397478,);
nor I_23170 (I397486,I397478,I397150);
DFFARX1 I_23171 (I397486,I3563,I397124,I397089,);
DFFARX1 I_23172 (I397478,I3563,I397124,I397107,);
nor I_23173 (I397531,I814239,I814227);
not I_23174 (I397548,I397531);
nor I_23175 (I397110,I397387,I397548);
nand I_23176 (I397095,I397404,I397548);
nor I_23177 (I397104,I397150,I397531);
DFFARX1 I_23178 (I397531,I3563,I397124,I397113,);
not I_23179 (I397651,I3570);
DFFARX1 I_23180 (I1023406,I3563,I397651,I397677,);
nand I_23181 (I397685,I1023403,I1023421);
and I_23182 (I397702,I397685,I1023412);
DFFARX1 I_23183 (I397702,I3563,I397651,I397728,);
nor I_23184 (I397619,I397728,I397677);
not I_23185 (I397750,I397728);
DFFARX1 I_23186 (I1023427,I3563,I397651,I397776,);
nand I_23187 (I397784,I397776,I1023409);
not I_23188 (I397801,I397784);
DFFARX1 I_23189 (I397801,I3563,I397651,I397827,);
not I_23190 (I397643,I397827);
nor I_23191 (I397849,I397677,I397784);
nor I_23192 (I397625,I397728,I397849);
DFFARX1 I_23193 (I1023415,I3563,I397651,I397889,);
DFFARX1 I_23194 (I397889,I3563,I397651,I397906,);
not I_23195 (I397914,I397906);
not I_23196 (I397931,I397889);
nand I_23197 (I397628,I397931,I397750);
nand I_23198 (I397962,I1023403,I1023430);
and I_23199 (I397979,I397962,I1023418);
DFFARX1 I_23200 (I397979,I3563,I397651,I398005,);
nor I_23201 (I398013,I398005,I397677);
DFFARX1 I_23202 (I398013,I3563,I397651,I397616,);
DFFARX1 I_23203 (I398005,I3563,I397651,I397634,);
nor I_23204 (I398058,I1023424,I1023430);
not I_23205 (I398075,I398058);
nor I_23206 (I397637,I397914,I398075);
nand I_23207 (I397622,I397931,I398075);
nor I_23208 (I397631,I397677,I398058);
DFFARX1 I_23209 (I398058,I3563,I397651,I397640,);
not I_23210 (I398178,I3570);
DFFARX1 I_23211 (I198223,I3563,I398178,I398204,);
nand I_23212 (I398212,I198223,I198229);
and I_23213 (I398229,I398212,I198247);
DFFARX1 I_23214 (I398229,I3563,I398178,I398255,);
nor I_23215 (I398146,I398255,I398204);
not I_23216 (I398277,I398255);
DFFARX1 I_23217 (I198235,I3563,I398178,I398303,);
nand I_23218 (I398311,I398303,I198232);
not I_23219 (I398328,I398311);
DFFARX1 I_23220 (I398328,I3563,I398178,I398354,);
not I_23221 (I398170,I398354);
nor I_23222 (I398376,I398204,I398311);
nor I_23223 (I398152,I398255,I398376);
DFFARX1 I_23224 (I198241,I3563,I398178,I398416,);
DFFARX1 I_23225 (I398416,I3563,I398178,I398433,);
not I_23226 (I398441,I398433);
not I_23227 (I398458,I398416);
nand I_23228 (I398155,I398458,I398277);
nand I_23229 (I398489,I198226,I198226);
and I_23230 (I398506,I398489,I198238);
DFFARX1 I_23231 (I398506,I3563,I398178,I398532,);
nor I_23232 (I398540,I398532,I398204);
DFFARX1 I_23233 (I398540,I3563,I398178,I398143,);
DFFARX1 I_23234 (I398532,I3563,I398178,I398161,);
nor I_23235 (I398585,I198244,I198226);
not I_23236 (I398602,I398585);
nor I_23237 (I398164,I398441,I398602);
nand I_23238 (I398149,I398458,I398602);
nor I_23239 (I398158,I398204,I398585);
DFFARX1 I_23240 (I398585,I3563,I398178,I398167,);
not I_23241 (I398705,I3570);
DFFARX1 I_23242 (I1190989,I3563,I398705,I398731,);
nand I_23243 (I398739,I1191004,I1190989);
and I_23244 (I398756,I398739,I1191007);
DFFARX1 I_23245 (I398756,I3563,I398705,I398782,);
nor I_23246 (I398673,I398782,I398731);
not I_23247 (I398804,I398782);
DFFARX1 I_23248 (I1191013,I3563,I398705,I398830,);
nand I_23249 (I398838,I398830,I1190995);
not I_23250 (I398855,I398838);
DFFARX1 I_23251 (I398855,I3563,I398705,I398881,);
not I_23252 (I398697,I398881);
nor I_23253 (I398903,I398731,I398838);
nor I_23254 (I398679,I398782,I398903);
DFFARX1 I_23255 (I1190992,I3563,I398705,I398943,);
DFFARX1 I_23256 (I398943,I3563,I398705,I398960,);
not I_23257 (I398968,I398960);
not I_23258 (I398985,I398943);
nand I_23259 (I398682,I398985,I398804);
nand I_23260 (I399016,I1190992,I1190998);
and I_23261 (I399033,I399016,I1191010);
DFFARX1 I_23262 (I399033,I3563,I398705,I399059,);
nor I_23263 (I399067,I399059,I398731);
DFFARX1 I_23264 (I399067,I3563,I398705,I398670,);
DFFARX1 I_23265 (I399059,I3563,I398705,I398688,);
nor I_23266 (I399112,I1191001,I1190998);
not I_23267 (I399129,I399112);
nor I_23268 (I398691,I398968,I399129);
nand I_23269 (I398676,I398985,I399129);
nor I_23270 (I398685,I398731,I399112);
DFFARX1 I_23271 (I399112,I3563,I398705,I398694,);
not I_23272 (I399232,I3570);
DFFARX1 I_23273 (I16595,I3563,I399232,I399258,);
nand I_23274 (I399266,I16619,I16598);
and I_23275 (I399283,I399266,I16595);
DFFARX1 I_23276 (I399283,I3563,I399232,I399309,);
nor I_23277 (I399200,I399309,I399258);
not I_23278 (I399331,I399309);
DFFARX1 I_23279 (I16601,I3563,I399232,I399357,);
nand I_23280 (I399365,I399357,I16610);
not I_23281 (I399382,I399365);
DFFARX1 I_23282 (I399382,I3563,I399232,I399408,);
not I_23283 (I399224,I399408);
nor I_23284 (I399430,I399258,I399365);
nor I_23285 (I399206,I399309,I399430);
DFFARX1 I_23286 (I16604,I3563,I399232,I399470,);
DFFARX1 I_23287 (I399470,I3563,I399232,I399487,);
not I_23288 (I399495,I399487);
not I_23289 (I399512,I399470);
nand I_23290 (I399209,I399512,I399331);
nand I_23291 (I399543,I16616,I16598);
and I_23292 (I399560,I399543,I16607);
DFFARX1 I_23293 (I399560,I3563,I399232,I399586,);
nor I_23294 (I399594,I399586,I399258);
DFFARX1 I_23295 (I399594,I3563,I399232,I399197,);
DFFARX1 I_23296 (I399586,I3563,I399232,I399215,);
nor I_23297 (I399639,I16613,I16598);
not I_23298 (I399656,I399639);
nor I_23299 (I399218,I399495,I399656);
nand I_23300 (I399203,I399512,I399656);
nor I_23301 (I399212,I399258,I399639);
DFFARX1 I_23302 (I399639,I3563,I399232,I399221,);
not I_23303 (I399759,I3570);
DFFARX1 I_23304 (I1015008,I3563,I399759,I399785,);
nand I_23305 (I399793,I1015005,I1015023);
and I_23306 (I399810,I399793,I1015014);
DFFARX1 I_23307 (I399810,I3563,I399759,I399836,);
nor I_23308 (I399727,I399836,I399785);
not I_23309 (I399858,I399836);
DFFARX1 I_23310 (I1015029,I3563,I399759,I399884,);
nand I_23311 (I399892,I399884,I1015011);
not I_23312 (I399909,I399892);
DFFARX1 I_23313 (I399909,I3563,I399759,I399935,);
not I_23314 (I399751,I399935);
nor I_23315 (I399957,I399785,I399892);
nor I_23316 (I399733,I399836,I399957);
DFFARX1 I_23317 (I1015017,I3563,I399759,I399997,);
DFFARX1 I_23318 (I399997,I3563,I399759,I400014,);
not I_23319 (I400022,I400014);
not I_23320 (I400039,I399997);
nand I_23321 (I399736,I400039,I399858);
nand I_23322 (I400070,I1015005,I1015032);
and I_23323 (I400087,I400070,I1015020);
DFFARX1 I_23324 (I400087,I3563,I399759,I400113,);
nor I_23325 (I400121,I400113,I399785);
DFFARX1 I_23326 (I400121,I3563,I399759,I399724,);
DFFARX1 I_23327 (I400113,I3563,I399759,I399742,);
nor I_23328 (I400166,I1015026,I1015032);
not I_23329 (I400183,I400166);
nor I_23330 (I399745,I400022,I400183);
nand I_23331 (I399730,I400039,I400183);
nor I_23332 (I399739,I399785,I400166);
DFFARX1 I_23333 (I400166,I3563,I399759,I399748,);
not I_23334 (I400286,I3570);
DFFARX1 I_23335 (I936196,I3563,I400286,I400312,);
nand I_23336 (I400320,I936193,I936211);
and I_23337 (I400337,I400320,I936202);
DFFARX1 I_23338 (I400337,I3563,I400286,I400363,);
nor I_23339 (I400254,I400363,I400312);
not I_23340 (I400385,I400363);
DFFARX1 I_23341 (I936217,I3563,I400286,I400411,);
nand I_23342 (I400419,I400411,I936199);
not I_23343 (I400436,I400419);
DFFARX1 I_23344 (I400436,I3563,I400286,I400462,);
not I_23345 (I400278,I400462);
nor I_23346 (I400484,I400312,I400419);
nor I_23347 (I400260,I400363,I400484);
DFFARX1 I_23348 (I936205,I3563,I400286,I400524,);
DFFARX1 I_23349 (I400524,I3563,I400286,I400541,);
not I_23350 (I400549,I400541);
not I_23351 (I400566,I400524);
nand I_23352 (I400263,I400566,I400385);
nand I_23353 (I400597,I936193,I936220);
and I_23354 (I400614,I400597,I936208);
DFFARX1 I_23355 (I400614,I3563,I400286,I400640,);
nor I_23356 (I400648,I400640,I400312);
DFFARX1 I_23357 (I400648,I3563,I400286,I400251,);
DFFARX1 I_23358 (I400640,I3563,I400286,I400269,);
nor I_23359 (I400693,I936214,I936220);
not I_23360 (I400710,I400693);
nor I_23361 (I400272,I400549,I400710);
nand I_23362 (I400257,I400566,I400710);
nor I_23363 (I400266,I400312,I400693);
DFFARX1 I_23364 (I400693,I3563,I400286,I400275,);
not I_23365 (I400813,I3570);
DFFARX1 I_23366 (I1002734,I3563,I400813,I400839,);
nand I_23367 (I400847,I1002731,I1002749);
and I_23368 (I400864,I400847,I1002740);
DFFARX1 I_23369 (I400864,I3563,I400813,I400890,);
nor I_23370 (I400781,I400890,I400839);
not I_23371 (I400912,I400890);
DFFARX1 I_23372 (I1002755,I3563,I400813,I400938,);
nand I_23373 (I400946,I400938,I1002737);
not I_23374 (I400963,I400946);
DFFARX1 I_23375 (I400963,I3563,I400813,I400989,);
not I_23376 (I400805,I400989);
nor I_23377 (I401011,I400839,I400946);
nor I_23378 (I400787,I400890,I401011);
DFFARX1 I_23379 (I1002743,I3563,I400813,I401051,);
DFFARX1 I_23380 (I401051,I3563,I400813,I401068,);
not I_23381 (I401076,I401068);
not I_23382 (I401093,I401051);
nand I_23383 (I400790,I401093,I400912);
nand I_23384 (I401124,I1002731,I1002758);
and I_23385 (I401141,I401124,I1002746);
DFFARX1 I_23386 (I401141,I3563,I400813,I401167,);
nor I_23387 (I401175,I401167,I400839);
DFFARX1 I_23388 (I401175,I3563,I400813,I400778,);
DFFARX1 I_23389 (I401167,I3563,I400813,I400796,);
nor I_23390 (I401220,I1002752,I1002758);
not I_23391 (I401237,I401220);
nor I_23392 (I400799,I401076,I401237);
nand I_23393 (I400784,I401093,I401237);
nor I_23394 (I400793,I400839,I401220);
DFFARX1 I_23395 (I401220,I3563,I400813,I400802,);
not I_23396 (I401340,I3570);
DFFARX1 I_23397 (I36094,I3563,I401340,I401366,);
nand I_23398 (I401374,I36118,I36097);
and I_23399 (I401391,I401374,I36094);
DFFARX1 I_23400 (I401391,I3563,I401340,I401417,);
nor I_23401 (I401308,I401417,I401366);
not I_23402 (I401439,I401417);
DFFARX1 I_23403 (I36100,I3563,I401340,I401465,);
nand I_23404 (I401473,I401465,I36109);
not I_23405 (I401490,I401473);
DFFARX1 I_23406 (I401490,I3563,I401340,I401516,);
not I_23407 (I401332,I401516);
nor I_23408 (I401538,I401366,I401473);
nor I_23409 (I401314,I401417,I401538);
DFFARX1 I_23410 (I36103,I3563,I401340,I401578,);
DFFARX1 I_23411 (I401578,I3563,I401340,I401595,);
not I_23412 (I401603,I401595);
not I_23413 (I401620,I401578);
nand I_23414 (I401317,I401620,I401439);
nand I_23415 (I401651,I36115,I36097);
and I_23416 (I401668,I401651,I36106);
DFFARX1 I_23417 (I401668,I3563,I401340,I401694,);
nor I_23418 (I401702,I401694,I401366);
DFFARX1 I_23419 (I401702,I3563,I401340,I401305,);
DFFARX1 I_23420 (I401694,I3563,I401340,I401323,);
nor I_23421 (I401747,I36112,I36097);
not I_23422 (I401764,I401747);
nor I_23423 (I401326,I401603,I401764);
nand I_23424 (I401311,I401620,I401764);
nor I_23425 (I401320,I401366,I401747);
DFFARX1 I_23426 (I401747,I3563,I401340,I401329,);
not I_23427 (I401867,I3570);
DFFARX1 I_23428 (I998212,I3563,I401867,I401893,);
nand I_23429 (I401901,I998209,I998227);
and I_23430 (I401918,I401901,I998218);
DFFARX1 I_23431 (I401918,I3563,I401867,I401944,);
nor I_23432 (I401835,I401944,I401893);
not I_23433 (I401966,I401944);
DFFARX1 I_23434 (I998233,I3563,I401867,I401992,);
nand I_23435 (I402000,I401992,I998215);
not I_23436 (I402017,I402000);
DFFARX1 I_23437 (I402017,I3563,I401867,I402043,);
not I_23438 (I401859,I402043);
nor I_23439 (I402065,I401893,I402000);
nor I_23440 (I401841,I401944,I402065);
DFFARX1 I_23441 (I998221,I3563,I401867,I402105,);
DFFARX1 I_23442 (I402105,I3563,I401867,I402122,);
not I_23443 (I402130,I402122);
not I_23444 (I402147,I402105);
nand I_23445 (I401844,I402147,I401966);
nand I_23446 (I402178,I998209,I998236);
and I_23447 (I402195,I402178,I998224);
DFFARX1 I_23448 (I402195,I3563,I401867,I402221,);
nor I_23449 (I402229,I402221,I401893);
DFFARX1 I_23450 (I402229,I3563,I401867,I401832,);
DFFARX1 I_23451 (I402221,I3563,I401867,I401850,);
nor I_23452 (I402274,I998230,I998236);
not I_23453 (I402291,I402274);
nor I_23454 (I401853,I402130,I402291);
nand I_23455 (I401838,I402147,I402291);
nor I_23456 (I401847,I401893,I402274);
DFFARX1 I_23457 (I402274,I3563,I401867,I401856,);
not I_23458 (I402394,I3570);
DFFARX1 I_23459 (I22392,I3563,I402394,I402420,);
nand I_23460 (I402428,I22416,I22395);
and I_23461 (I402445,I402428,I22392);
DFFARX1 I_23462 (I402445,I3563,I402394,I402471,);
nor I_23463 (I402362,I402471,I402420);
not I_23464 (I402493,I402471);
DFFARX1 I_23465 (I22398,I3563,I402394,I402519,);
nand I_23466 (I402527,I402519,I22407);
not I_23467 (I402544,I402527);
DFFARX1 I_23468 (I402544,I3563,I402394,I402570,);
not I_23469 (I402386,I402570);
nor I_23470 (I402592,I402420,I402527);
nor I_23471 (I402368,I402471,I402592);
DFFARX1 I_23472 (I22401,I3563,I402394,I402632,);
DFFARX1 I_23473 (I402632,I3563,I402394,I402649,);
not I_23474 (I402657,I402649);
not I_23475 (I402674,I402632);
nand I_23476 (I402371,I402674,I402493);
nand I_23477 (I402705,I22413,I22395);
and I_23478 (I402722,I402705,I22404);
DFFARX1 I_23479 (I402722,I3563,I402394,I402748,);
nor I_23480 (I402756,I402748,I402420);
DFFARX1 I_23481 (I402756,I3563,I402394,I402359,);
DFFARX1 I_23482 (I402748,I3563,I402394,I402377,);
nor I_23483 (I402801,I22410,I22395);
not I_23484 (I402818,I402801);
nor I_23485 (I402380,I402657,I402818);
nand I_23486 (I402365,I402674,I402818);
nor I_23487 (I402374,I402420,I402801);
DFFARX1 I_23488 (I402801,I3563,I402394,I402383,);
not I_23489 (I402921,I3570);
DFFARX1 I_23490 (I11918,I3563,I402921,I402947,);
nand I_23491 (I402955,I11909,I11912);
and I_23492 (I402972,I402955,I11903);
DFFARX1 I_23493 (I402972,I3563,I402921,I402998,);
nor I_23494 (I402889,I402998,I402947);
not I_23495 (I403020,I402998);
DFFARX1 I_23496 (I11909,I3563,I402921,I403046,);
nand I_23497 (I403054,I403046,I11915);
not I_23498 (I403071,I403054);
DFFARX1 I_23499 (I403071,I3563,I402921,I403097,);
not I_23500 (I402913,I403097);
nor I_23501 (I403119,I402947,I403054);
nor I_23502 (I402895,I402998,I403119);
DFFARX1 I_23503 (I11906,I3563,I402921,I403159,);
DFFARX1 I_23504 (I403159,I3563,I402921,I403176,);
not I_23505 (I403184,I403176);
not I_23506 (I403201,I403159);
nand I_23507 (I402898,I403201,I403020);
nand I_23508 (I403232,I11906,I11921);
and I_23509 (I403249,I403232,I11903);
DFFARX1 I_23510 (I403249,I3563,I402921,I403275,);
nor I_23511 (I403283,I403275,I402947);
DFFARX1 I_23512 (I403283,I3563,I402921,I402886,);
DFFARX1 I_23513 (I403275,I3563,I402921,I402904,);
nor I_23514 (I403328,I11924,I11921);
not I_23515 (I403345,I403328);
nor I_23516 (I402907,I403184,I403345);
nand I_23517 (I402892,I403201,I403345);
nor I_23518 (I402901,I402947,I403328);
DFFARX1 I_23519 (I403328,I3563,I402921,I402910,);
not I_23520 (I403448,I3570);
DFFARX1 I_23521 (I711023,I3563,I403448,I403474,);
nand I_23522 (I403482,I711014,I711029);
and I_23523 (I403499,I403482,I711035);
DFFARX1 I_23524 (I403499,I3563,I403448,I403525,);
nor I_23525 (I403416,I403525,I403474);
not I_23526 (I403547,I403525);
DFFARX1 I_23527 (I711020,I3563,I403448,I403573,);
nand I_23528 (I403581,I403573,I711014);
not I_23529 (I403598,I403581);
DFFARX1 I_23530 (I403598,I3563,I403448,I403624,);
not I_23531 (I403440,I403624);
nor I_23532 (I403646,I403474,I403581);
nor I_23533 (I403422,I403525,I403646);
DFFARX1 I_23534 (I711017,I3563,I403448,I403686,);
DFFARX1 I_23535 (I403686,I3563,I403448,I403703,);
not I_23536 (I403711,I403703);
not I_23537 (I403728,I403686);
nand I_23538 (I403425,I403728,I403547);
nand I_23539 (I403759,I711011,I711026);
and I_23540 (I403776,I403759,I711011);
DFFARX1 I_23541 (I403776,I3563,I403448,I403802,);
nor I_23542 (I403810,I403802,I403474);
DFFARX1 I_23543 (I403810,I3563,I403448,I403413,);
DFFARX1 I_23544 (I403802,I3563,I403448,I403431,);
nor I_23545 (I403855,I711032,I711026);
not I_23546 (I403872,I403855);
nor I_23547 (I403434,I403711,I403872);
nand I_23548 (I403419,I403728,I403872);
nor I_23549 (I403428,I403474,I403855);
DFFARX1 I_23550 (I403855,I3563,I403448,I403437,);
not I_23551 (I403975,I3570);
DFFARX1 I_23552 (I927152,I3563,I403975,I404001,);
nand I_23553 (I404009,I927149,I927167);
and I_23554 (I404026,I404009,I927158);
DFFARX1 I_23555 (I404026,I3563,I403975,I404052,);
nor I_23556 (I403943,I404052,I404001);
not I_23557 (I404074,I404052);
DFFARX1 I_23558 (I927173,I3563,I403975,I404100,);
nand I_23559 (I404108,I404100,I927155);
not I_23560 (I404125,I404108);
DFFARX1 I_23561 (I404125,I3563,I403975,I404151,);
not I_23562 (I403967,I404151);
nor I_23563 (I404173,I404001,I404108);
nor I_23564 (I403949,I404052,I404173);
DFFARX1 I_23565 (I927161,I3563,I403975,I404213,);
DFFARX1 I_23566 (I404213,I3563,I403975,I404230,);
not I_23567 (I404238,I404230);
not I_23568 (I404255,I404213);
nand I_23569 (I403952,I404255,I404074);
nand I_23570 (I404286,I927149,I927176);
and I_23571 (I404303,I404286,I927164);
DFFARX1 I_23572 (I404303,I3563,I403975,I404329,);
nor I_23573 (I404337,I404329,I404001);
DFFARX1 I_23574 (I404337,I3563,I403975,I403940,);
DFFARX1 I_23575 (I404329,I3563,I403975,I403958,);
nor I_23576 (I404382,I927170,I927176);
not I_23577 (I404399,I404382);
nor I_23578 (I403961,I404238,I404399);
nand I_23579 (I403946,I404255,I404399);
nor I_23580 (I403955,I404001,I404382);
DFFARX1 I_23581 (I404382,I3563,I403975,I403964,);
not I_23582 (I404502,I3570);
DFFARX1 I_23583 (I695995,I3563,I404502,I404528,);
nand I_23584 (I404536,I695986,I696001);
and I_23585 (I404553,I404536,I696007);
DFFARX1 I_23586 (I404553,I3563,I404502,I404579,);
nor I_23587 (I404470,I404579,I404528);
not I_23588 (I404601,I404579);
DFFARX1 I_23589 (I695992,I3563,I404502,I404627,);
nand I_23590 (I404635,I404627,I695986);
not I_23591 (I404652,I404635);
DFFARX1 I_23592 (I404652,I3563,I404502,I404678,);
not I_23593 (I404494,I404678);
nor I_23594 (I404700,I404528,I404635);
nor I_23595 (I404476,I404579,I404700);
DFFARX1 I_23596 (I695989,I3563,I404502,I404740,);
DFFARX1 I_23597 (I404740,I3563,I404502,I404757,);
not I_23598 (I404765,I404757);
not I_23599 (I404782,I404740);
nand I_23600 (I404479,I404782,I404601);
nand I_23601 (I404813,I695983,I695998);
and I_23602 (I404830,I404813,I695983);
DFFARX1 I_23603 (I404830,I3563,I404502,I404856,);
nor I_23604 (I404864,I404856,I404528);
DFFARX1 I_23605 (I404864,I3563,I404502,I404467,);
DFFARX1 I_23606 (I404856,I3563,I404502,I404485,);
nor I_23607 (I404909,I696004,I695998);
not I_23608 (I404926,I404909);
nor I_23609 (I404488,I404765,I404926);
nand I_23610 (I404473,I404782,I404926);
nor I_23611 (I404482,I404528,I404909);
DFFARX1 I_23612 (I404909,I3563,I404502,I404491,);
not I_23613 (I405029,I3570);
DFFARX1 I_23614 (I1357134,I3563,I405029,I405055,);
nand I_23615 (I405063,I1357113,I1357113);
and I_23616 (I405080,I405063,I1357140);
DFFARX1 I_23617 (I405080,I3563,I405029,I405106,);
nor I_23618 (I404997,I405106,I405055);
not I_23619 (I405128,I405106);
DFFARX1 I_23620 (I1357128,I3563,I405029,I405154,);
nand I_23621 (I405162,I405154,I1357131);
not I_23622 (I405179,I405162);
DFFARX1 I_23623 (I405179,I3563,I405029,I405205,);
not I_23624 (I405021,I405205);
nor I_23625 (I405227,I405055,I405162);
nor I_23626 (I405003,I405106,I405227);
DFFARX1 I_23627 (I1357122,I3563,I405029,I405267,);
DFFARX1 I_23628 (I405267,I3563,I405029,I405284,);
not I_23629 (I405292,I405284);
not I_23630 (I405309,I405267);
nand I_23631 (I405006,I405309,I405128);
nand I_23632 (I405340,I1357119,I1357116);
and I_23633 (I405357,I405340,I1357137);
DFFARX1 I_23634 (I405357,I3563,I405029,I405383,);
nor I_23635 (I405391,I405383,I405055);
DFFARX1 I_23636 (I405391,I3563,I405029,I404994,);
DFFARX1 I_23637 (I405383,I3563,I405029,I405012,);
nor I_23638 (I405436,I1357125,I1357116);
not I_23639 (I405453,I405436);
nor I_23640 (I405015,I405292,I405453);
nand I_23641 (I405000,I405309,I405453);
nor I_23642 (I405009,I405055,I405436);
DFFARX1 I_23643 (I405436,I3563,I405029,I405018,);
not I_23644 (I405556,I3570);
DFFARX1 I_23645 (I1028574,I3563,I405556,I405582,);
nand I_23646 (I405590,I1028571,I1028589);
and I_23647 (I405607,I405590,I1028580);
DFFARX1 I_23648 (I405607,I3563,I405556,I405633,);
nor I_23649 (I405524,I405633,I405582);
not I_23650 (I405655,I405633);
DFFARX1 I_23651 (I1028595,I3563,I405556,I405681,);
nand I_23652 (I405689,I405681,I1028577);
not I_23653 (I405706,I405689);
DFFARX1 I_23654 (I405706,I3563,I405556,I405732,);
not I_23655 (I405548,I405732);
nor I_23656 (I405754,I405582,I405689);
nor I_23657 (I405530,I405633,I405754);
DFFARX1 I_23658 (I1028583,I3563,I405556,I405794,);
DFFARX1 I_23659 (I405794,I3563,I405556,I405811,);
not I_23660 (I405819,I405811);
not I_23661 (I405836,I405794);
nand I_23662 (I405533,I405836,I405655);
nand I_23663 (I405867,I1028571,I1028598);
and I_23664 (I405884,I405867,I1028586);
DFFARX1 I_23665 (I405884,I3563,I405556,I405910,);
nor I_23666 (I405918,I405910,I405582);
DFFARX1 I_23667 (I405918,I3563,I405556,I405521,);
DFFARX1 I_23668 (I405910,I3563,I405556,I405539,);
nor I_23669 (I405963,I1028592,I1028598);
not I_23670 (I405980,I405963);
nor I_23671 (I405542,I405819,I405980);
nand I_23672 (I405527,I405836,I405980);
nor I_23673 (I405536,I405582,I405963);
DFFARX1 I_23674 (I405963,I3563,I405556,I405545,);
not I_23675 (I406083,I3570);
DFFARX1 I_23676 (I824234,I3563,I406083,I406109,);
nand I_23677 (I406117,I824237,I824231);
and I_23678 (I406134,I406117,I824243);
DFFARX1 I_23679 (I406134,I3563,I406083,I406160,);
nor I_23680 (I406051,I406160,I406109);
not I_23681 (I406182,I406160);
DFFARX1 I_23682 (I824246,I3563,I406083,I406208,);
nand I_23683 (I406216,I406208,I824237);
not I_23684 (I406233,I406216);
DFFARX1 I_23685 (I406233,I3563,I406083,I406259,);
not I_23686 (I406075,I406259);
nor I_23687 (I406281,I406109,I406216);
nor I_23688 (I406057,I406160,I406281);
DFFARX1 I_23689 (I824249,I3563,I406083,I406321,);
DFFARX1 I_23690 (I406321,I3563,I406083,I406338,);
not I_23691 (I406346,I406338);
not I_23692 (I406363,I406321);
nand I_23693 (I406060,I406363,I406182);
nand I_23694 (I406394,I824231,I824240);
and I_23695 (I406411,I406394,I824234);
DFFARX1 I_23696 (I406411,I3563,I406083,I406437,);
nor I_23697 (I406445,I406437,I406109);
DFFARX1 I_23698 (I406445,I3563,I406083,I406048,);
DFFARX1 I_23699 (I406437,I3563,I406083,I406066,);
nor I_23700 (I406490,I824252,I824240);
not I_23701 (I406507,I406490);
nor I_23702 (I406069,I406346,I406507);
nand I_23703 (I406054,I406363,I406507);
nor I_23704 (I406063,I406109,I406490);
DFFARX1 I_23705 (I406490,I3563,I406083,I406072,);
not I_23706 (I406610,I3570);
DFFARX1 I_23707 (I2956,I3563,I406610,I406636,);
nand I_23708 (I406644,I2420,I3508);
and I_23709 (I406661,I406644,I3340);
DFFARX1 I_23710 (I406661,I3563,I406610,I406687,);
nor I_23711 (I406578,I406687,I406636);
not I_23712 (I406709,I406687);
DFFARX1 I_23713 (I2084,I3563,I406610,I406735,);
nand I_23714 (I406743,I406735,I1468);
not I_23715 (I406760,I406743);
DFFARX1 I_23716 (I406760,I3563,I406610,I406786,);
not I_23717 (I406602,I406786);
nor I_23718 (I406808,I406636,I406743);
nor I_23719 (I406584,I406687,I406808);
DFFARX1 I_23720 (I2812,I3563,I406610,I406848,);
DFFARX1 I_23721 (I406848,I3563,I406610,I406865,);
not I_23722 (I406873,I406865);
not I_23723 (I406890,I406848);
nand I_23724 (I406587,I406890,I406709);
nand I_23725 (I406921,I1524,I2548);
and I_23726 (I406938,I406921,I3516);
DFFARX1 I_23727 (I406938,I3563,I406610,I406964,);
nor I_23728 (I406972,I406964,I406636);
DFFARX1 I_23729 (I406972,I3563,I406610,I406575,);
DFFARX1 I_23730 (I406964,I3563,I406610,I406593,);
nor I_23731 (I407017,I1716,I2548);
not I_23732 (I407034,I407017);
nor I_23733 (I406596,I406873,I407034);
nand I_23734 (I406581,I406890,I407034);
nor I_23735 (I406590,I406636,I407017);
DFFARX1 I_23736 (I407017,I3563,I406610,I406599,);
not I_23737 (I407137,I3570);
DFFARX1 I_23738 (I486606,I3563,I407137,I407163,);
nand I_23739 (I407171,I486618,I486597);
and I_23740 (I407188,I407171,I486621);
DFFARX1 I_23741 (I407188,I3563,I407137,I407214,);
nor I_23742 (I407105,I407214,I407163);
not I_23743 (I407236,I407214);
DFFARX1 I_23744 (I486612,I3563,I407137,I407262,);
nand I_23745 (I407270,I407262,I486594);
not I_23746 (I407287,I407270);
DFFARX1 I_23747 (I407287,I3563,I407137,I407313,);
not I_23748 (I407129,I407313);
nor I_23749 (I407335,I407163,I407270);
nor I_23750 (I407111,I407214,I407335);
DFFARX1 I_23751 (I486609,I3563,I407137,I407375,);
DFFARX1 I_23752 (I407375,I3563,I407137,I407392,);
not I_23753 (I407400,I407392);
not I_23754 (I407417,I407375);
nand I_23755 (I407114,I407417,I407236);
nand I_23756 (I407448,I486594,I486600);
and I_23757 (I407465,I407448,I486603);
DFFARX1 I_23758 (I407465,I3563,I407137,I407491,);
nor I_23759 (I407499,I407491,I407163);
DFFARX1 I_23760 (I407499,I3563,I407137,I407102,);
DFFARX1 I_23761 (I407491,I3563,I407137,I407120,);
nor I_23762 (I407544,I486615,I486600);
not I_23763 (I407561,I407544);
nor I_23764 (I407123,I407400,I407561);
nand I_23765 (I407108,I407417,I407561);
nor I_23766 (I407117,I407163,I407544);
DFFARX1 I_23767 (I407544,I3563,I407137,I407126,);
not I_23768 (I407664,I3570);
DFFARX1 I_23769 (I181563,I3563,I407664,I407690,);
nand I_23770 (I407698,I181563,I181569);
and I_23771 (I407715,I407698,I181587);
DFFARX1 I_23772 (I407715,I3563,I407664,I407741,);
nor I_23773 (I407632,I407741,I407690);
not I_23774 (I407763,I407741);
DFFARX1 I_23775 (I181575,I3563,I407664,I407789,);
nand I_23776 (I407797,I407789,I181572);
not I_23777 (I407814,I407797);
DFFARX1 I_23778 (I407814,I3563,I407664,I407840,);
not I_23779 (I407656,I407840);
nor I_23780 (I407862,I407690,I407797);
nor I_23781 (I407638,I407741,I407862);
DFFARX1 I_23782 (I181581,I3563,I407664,I407902,);
DFFARX1 I_23783 (I407902,I3563,I407664,I407919,);
not I_23784 (I407927,I407919);
not I_23785 (I407944,I407902);
nand I_23786 (I407641,I407944,I407763);
nand I_23787 (I407975,I181566,I181566);
and I_23788 (I407992,I407975,I181578);
DFFARX1 I_23789 (I407992,I3563,I407664,I408018,);
nor I_23790 (I408026,I408018,I407690);
DFFARX1 I_23791 (I408026,I3563,I407664,I407629,);
DFFARX1 I_23792 (I408018,I3563,I407664,I407647,);
nor I_23793 (I408071,I181584,I181566);
not I_23794 (I408088,I408071);
nor I_23795 (I407650,I407927,I408088);
nand I_23796 (I407635,I407944,I408088);
nor I_23797 (I407644,I407690,I408071);
DFFARX1 I_23798 (I408071,I3563,I407664,I407653,);
not I_23799 (I408191,I3570);
DFFARX1 I_23800 (I625482,I3563,I408191,I408217,);
nand I_23801 (I408225,I625467,I625470);
and I_23802 (I408242,I408225,I625485);
DFFARX1 I_23803 (I408242,I3563,I408191,I408268,);
nor I_23804 (I408159,I408268,I408217);
not I_23805 (I408290,I408268);
DFFARX1 I_23806 (I625479,I3563,I408191,I408316,);
nand I_23807 (I408324,I408316,I625470);
not I_23808 (I408341,I408324);
DFFARX1 I_23809 (I408341,I3563,I408191,I408367,);
not I_23810 (I408183,I408367);
nor I_23811 (I408389,I408217,I408324);
nor I_23812 (I408165,I408268,I408389);
DFFARX1 I_23813 (I625476,I3563,I408191,I408429,);
DFFARX1 I_23814 (I408429,I3563,I408191,I408446,);
not I_23815 (I408454,I408446);
not I_23816 (I408471,I408429);
nand I_23817 (I408168,I408471,I408290);
nand I_23818 (I408502,I625491,I625467);
and I_23819 (I408519,I408502,I625488);
DFFARX1 I_23820 (I408519,I3563,I408191,I408545,);
nor I_23821 (I408553,I408545,I408217);
DFFARX1 I_23822 (I408553,I3563,I408191,I408156,);
DFFARX1 I_23823 (I408545,I3563,I408191,I408174,);
nor I_23824 (I408598,I625473,I625467);
not I_23825 (I408615,I408598);
nor I_23826 (I408177,I408454,I408615);
nand I_23827 (I408162,I408471,I408615);
nor I_23828 (I408171,I408217,I408598);
DFFARX1 I_23829 (I408598,I3563,I408191,I408180,);
not I_23830 (I408718,I3570);
DFFARX1 I_23831 (I1032450,I3563,I408718,I408744,);
nand I_23832 (I408752,I1032447,I1032465);
and I_23833 (I408769,I408752,I1032456);
DFFARX1 I_23834 (I408769,I3563,I408718,I408795,);
nor I_23835 (I408686,I408795,I408744);
not I_23836 (I408817,I408795);
DFFARX1 I_23837 (I1032471,I3563,I408718,I408843,);
nand I_23838 (I408851,I408843,I1032453);
not I_23839 (I408868,I408851);
DFFARX1 I_23840 (I408868,I3563,I408718,I408894,);
not I_23841 (I408710,I408894);
nor I_23842 (I408916,I408744,I408851);
nor I_23843 (I408692,I408795,I408916);
DFFARX1 I_23844 (I1032459,I3563,I408718,I408956,);
DFFARX1 I_23845 (I408956,I3563,I408718,I408973,);
not I_23846 (I408981,I408973);
not I_23847 (I408998,I408956);
nand I_23848 (I408695,I408998,I408817);
nand I_23849 (I409029,I1032447,I1032474);
and I_23850 (I409046,I409029,I1032462);
DFFARX1 I_23851 (I409046,I3563,I408718,I409072,);
nor I_23852 (I409080,I409072,I408744);
DFFARX1 I_23853 (I409080,I3563,I408718,I408683,);
DFFARX1 I_23854 (I409072,I3563,I408718,I408701,);
nor I_23855 (I409125,I1032468,I1032474);
not I_23856 (I409142,I409125);
nor I_23857 (I408704,I408981,I409142);
nand I_23858 (I408689,I408998,I409142);
nor I_23859 (I408698,I408744,I409125);
DFFARX1 I_23860 (I409125,I3563,I408718,I408707,);
not I_23861 (I409245,I3570);
DFFARX1 I_23862 (I1017592,I3563,I409245,I409271,);
nand I_23863 (I409279,I1017589,I1017607);
and I_23864 (I409296,I409279,I1017598);
DFFARX1 I_23865 (I409296,I3563,I409245,I409322,);
nor I_23866 (I409213,I409322,I409271);
not I_23867 (I409344,I409322);
DFFARX1 I_23868 (I1017613,I3563,I409245,I409370,);
nand I_23869 (I409378,I409370,I1017595);
not I_23870 (I409395,I409378);
DFFARX1 I_23871 (I409395,I3563,I409245,I409421,);
not I_23872 (I409237,I409421);
nor I_23873 (I409443,I409271,I409378);
nor I_23874 (I409219,I409322,I409443);
DFFARX1 I_23875 (I1017601,I3563,I409245,I409483,);
DFFARX1 I_23876 (I409483,I3563,I409245,I409500,);
not I_23877 (I409508,I409500);
not I_23878 (I409525,I409483);
nand I_23879 (I409222,I409525,I409344);
nand I_23880 (I409556,I1017589,I1017616);
and I_23881 (I409573,I409556,I1017604);
DFFARX1 I_23882 (I409573,I3563,I409245,I409599,);
nor I_23883 (I409607,I409599,I409271);
DFFARX1 I_23884 (I409607,I3563,I409245,I409210,);
DFFARX1 I_23885 (I409599,I3563,I409245,I409228,);
nor I_23886 (I409652,I1017610,I1017616);
not I_23887 (I409669,I409652);
nor I_23888 (I409231,I409508,I409669);
nand I_23889 (I409216,I409525,I409669);
nor I_23890 (I409225,I409271,I409652);
DFFARX1 I_23891 (I409652,I3563,I409245,I409234,);
not I_23892 (I409772,I3570);
DFFARX1 I_23893 (I904338,I3563,I409772,I409798,);
nand I_23894 (I409806,I904341,I904335);
and I_23895 (I409823,I409806,I904347);
DFFARX1 I_23896 (I409823,I3563,I409772,I409849,);
nor I_23897 (I409740,I409849,I409798);
not I_23898 (I409871,I409849);
DFFARX1 I_23899 (I904350,I3563,I409772,I409897,);
nand I_23900 (I409905,I409897,I904341);
not I_23901 (I409922,I409905);
DFFARX1 I_23902 (I409922,I3563,I409772,I409948,);
not I_23903 (I409764,I409948);
nor I_23904 (I409970,I409798,I409905);
nor I_23905 (I409746,I409849,I409970);
DFFARX1 I_23906 (I904353,I3563,I409772,I410010,);
DFFARX1 I_23907 (I410010,I3563,I409772,I410027,);
not I_23908 (I410035,I410027);
not I_23909 (I410052,I410010);
nand I_23910 (I409749,I410052,I409871);
nand I_23911 (I410083,I904335,I904344);
and I_23912 (I410100,I410083,I904338);
DFFARX1 I_23913 (I410100,I3563,I409772,I410126,);
nor I_23914 (I410134,I410126,I409798);
DFFARX1 I_23915 (I410134,I3563,I409772,I409737,);
DFFARX1 I_23916 (I410126,I3563,I409772,I409755,);
nor I_23917 (I410179,I904356,I904344);
not I_23918 (I410196,I410179);
nor I_23919 (I409758,I410035,I410196);
nand I_23920 (I409743,I410052,I410196);
nor I_23921 (I409752,I409798,I410179);
DFFARX1 I_23922 (I410179,I3563,I409772,I409761,);
not I_23923 (I410299,I3570);
DFFARX1 I_23924 (I1212375,I3563,I410299,I410325,);
nand I_23925 (I410333,I1212390,I1212375);
and I_23926 (I410350,I410333,I1212393);
DFFARX1 I_23927 (I410350,I3563,I410299,I410376,);
nor I_23928 (I410267,I410376,I410325);
not I_23929 (I410398,I410376);
DFFARX1 I_23930 (I1212399,I3563,I410299,I410424,);
nand I_23931 (I410432,I410424,I1212381);
not I_23932 (I410449,I410432);
DFFARX1 I_23933 (I410449,I3563,I410299,I410475,);
not I_23934 (I410291,I410475);
nor I_23935 (I410497,I410325,I410432);
nor I_23936 (I410273,I410376,I410497);
DFFARX1 I_23937 (I1212378,I3563,I410299,I410537,);
DFFARX1 I_23938 (I410537,I3563,I410299,I410554,);
not I_23939 (I410562,I410554);
not I_23940 (I410579,I410537);
nand I_23941 (I410276,I410579,I410398);
nand I_23942 (I410610,I1212378,I1212384);
and I_23943 (I410627,I410610,I1212396);
DFFARX1 I_23944 (I410627,I3563,I410299,I410653,);
nor I_23945 (I410661,I410653,I410325);
DFFARX1 I_23946 (I410661,I3563,I410299,I410264,);
DFFARX1 I_23947 (I410653,I3563,I410299,I410282,);
nor I_23948 (I410706,I1212387,I1212384);
not I_23949 (I410723,I410706);
nor I_23950 (I410285,I410562,I410723);
nand I_23951 (I410270,I410579,I410723);
nor I_23952 (I410279,I410325,I410706);
DFFARX1 I_23953 (I410706,I3563,I410299,I410288,);
not I_23954 (I410826,I3570);
DFFARX1 I_23955 (I697729,I3563,I410826,I410852,);
nand I_23956 (I410860,I697720,I697735);
and I_23957 (I410877,I410860,I697741);
DFFARX1 I_23958 (I410877,I3563,I410826,I410903,);
nor I_23959 (I410794,I410903,I410852);
not I_23960 (I410925,I410903);
DFFARX1 I_23961 (I697726,I3563,I410826,I410951,);
nand I_23962 (I410959,I410951,I697720);
not I_23963 (I410976,I410959);
DFFARX1 I_23964 (I410976,I3563,I410826,I411002,);
not I_23965 (I410818,I411002);
nor I_23966 (I411024,I410852,I410959);
nor I_23967 (I410800,I410903,I411024);
DFFARX1 I_23968 (I697723,I3563,I410826,I411064,);
DFFARX1 I_23969 (I411064,I3563,I410826,I411081,);
not I_23970 (I411089,I411081);
not I_23971 (I411106,I411064);
nand I_23972 (I410803,I411106,I410925);
nand I_23973 (I411137,I697717,I697732);
and I_23974 (I411154,I411137,I697717);
DFFARX1 I_23975 (I411154,I3563,I410826,I411180,);
nor I_23976 (I411188,I411180,I410852);
DFFARX1 I_23977 (I411188,I3563,I410826,I410791,);
DFFARX1 I_23978 (I411180,I3563,I410826,I410809,);
nor I_23979 (I411233,I697738,I697732);
not I_23980 (I411250,I411233);
nor I_23981 (I410812,I411089,I411250);
nand I_23982 (I410797,I411106,I411250);
nor I_23983 (I410806,I410852,I411233);
DFFARX1 I_23984 (I411233,I3563,I410826,I410815,);
not I_23985 (I411353,I3570);
DFFARX1 I_23986 (I276763,I3563,I411353,I411379,);
nand I_23987 (I411387,I276763,I276769);
and I_23988 (I411404,I411387,I276787);
DFFARX1 I_23989 (I411404,I3563,I411353,I411430,);
nor I_23990 (I411321,I411430,I411379);
not I_23991 (I411452,I411430);
DFFARX1 I_23992 (I276775,I3563,I411353,I411478,);
nand I_23993 (I411486,I411478,I276772);
not I_23994 (I411503,I411486);
DFFARX1 I_23995 (I411503,I3563,I411353,I411529,);
not I_23996 (I411345,I411529);
nor I_23997 (I411551,I411379,I411486);
nor I_23998 (I411327,I411430,I411551);
DFFARX1 I_23999 (I276781,I3563,I411353,I411591,);
DFFARX1 I_24000 (I411591,I3563,I411353,I411608,);
not I_24001 (I411616,I411608);
not I_24002 (I411633,I411591);
nand I_24003 (I411330,I411633,I411452);
nand I_24004 (I411664,I276766,I276766);
and I_24005 (I411681,I411664,I276778);
DFFARX1 I_24006 (I411681,I3563,I411353,I411707,);
nor I_24007 (I411715,I411707,I411379);
DFFARX1 I_24008 (I411715,I3563,I411353,I411318,);
DFFARX1 I_24009 (I411707,I3563,I411353,I411336,);
nor I_24010 (I411760,I276784,I276766);
not I_24011 (I411777,I411760);
nor I_24012 (I411339,I411616,I411777);
nand I_24013 (I411324,I411633,I411777);
nor I_24014 (I411333,I411379,I411760);
DFFARX1 I_24015 (I411760,I3563,I411353,I411342,);
not I_24016 (I411880,I3570);
DFFARX1 I_24017 (I1184053,I3563,I411880,I411906,);
nand I_24018 (I411914,I1184068,I1184053);
and I_24019 (I411931,I411914,I1184071);
DFFARX1 I_24020 (I411931,I3563,I411880,I411957,);
nor I_24021 (I411848,I411957,I411906);
not I_24022 (I411979,I411957);
DFFARX1 I_24023 (I1184077,I3563,I411880,I412005,);
nand I_24024 (I412013,I412005,I1184059);
not I_24025 (I412030,I412013);
DFFARX1 I_24026 (I412030,I3563,I411880,I412056,);
not I_24027 (I411872,I412056);
nor I_24028 (I412078,I411906,I412013);
nor I_24029 (I411854,I411957,I412078);
DFFARX1 I_24030 (I1184056,I3563,I411880,I412118,);
DFFARX1 I_24031 (I412118,I3563,I411880,I412135,);
not I_24032 (I412143,I412135);
not I_24033 (I412160,I412118);
nand I_24034 (I411857,I412160,I411979);
nand I_24035 (I412191,I1184056,I1184062);
and I_24036 (I412208,I412191,I1184074);
DFFARX1 I_24037 (I412208,I3563,I411880,I412234,);
nor I_24038 (I412242,I412234,I411906);
DFFARX1 I_24039 (I412242,I3563,I411880,I411845,);
DFFARX1 I_24040 (I412234,I3563,I411880,I411863,);
nor I_24041 (I412287,I1184065,I1184062);
not I_24042 (I412304,I412287);
nor I_24043 (I411866,I412143,I412304);
nand I_24044 (I411851,I412160,I412304);
nor I_24045 (I411860,I411906,I412287);
DFFARX1 I_24046 (I412287,I3563,I411880,I411869,);
not I_24047 (I412407,I3570);
DFFARX1 I_24048 (I451790,I3563,I412407,I412433,);
nand I_24049 (I412441,I451802,I451781);
and I_24050 (I412458,I412441,I451805);
DFFARX1 I_24051 (I412458,I3563,I412407,I412484,);
nor I_24052 (I412375,I412484,I412433);
not I_24053 (I412506,I412484);
DFFARX1 I_24054 (I451796,I3563,I412407,I412532,);
nand I_24055 (I412540,I412532,I451778);
not I_24056 (I412557,I412540);
DFFARX1 I_24057 (I412557,I3563,I412407,I412583,);
not I_24058 (I412399,I412583);
nor I_24059 (I412605,I412433,I412540);
nor I_24060 (I412381,I412484,I412605);
DFFARX1 I_24061 (I451793,I3563,I412407,I412645,);
DFFARX1 I_24062 (I412645,I3563,I412407,I412662,);
not I_24063 (I412670,I412662);
not I_24064 (I412687,I412645);
nand I_24065 (I412384,I412687,I412506);
nand I_24066 (I412718,I451778,I451784);
and I_24067 (I412735,I412718,I451787);
DFFARX1 I_24068 (I412735,I3563,I412407,I412761,);
nor I_24069 (I412769,I412761,I412433);
DFFARX1 I_24070 (I412769,I3563,I412407,I412372,);
DFFARX1 I_24071 (I412761,I3563,I412407,I412390,);
nor I_24072 (I412814,I451799,I451784);
not I_24073 (I412831,I412814);
nor I_24074 (I412393,I412670,I412831);
nand I_24075 (I412378,I412687,I412831);
nor I_24076 (I412387,I412433,I412814);
DFFARX1 I_24077 (I412814,I3563,I412407,I412396,);
not I_24078 (I412934,I3570);
DFFARX1 I_24079 (I1379744,I3563,I412934,I412960,);
nand I_24080 (I412968,I1379723,I1379723);
and I_24081 (I412985,I412968,I1379750);
DFFARX1 I_24082 (I412985,I3563,I412934,I413011,);
nor I_24083 (I412902,I413011,I412960);
not I_24084 (I413033,I413011);
DFFARX1 I_24085 (I1379738,I3563,I412934,I413059,);
nand I_24086 (I413067,I413059,I1379741);
not I_24087 (I413084,I413067);
DFFARX1 I_24088 (I413084,I3563,I412934,I413110,);
not I_24089 (I412926,I413110);
nor I_24090 (I413132,I412960,I413067);
nor I_24091 (I412908,I413011,I413132);
DFFARX1 I_24092 (I1379732,I3563,I412934,I413172,);
DFFARX1 I_24093 (I413172,I3563,I412934,I413189,);
not I_24094 (I413197,I413189);
not I_24095 (I413214,I413172);
nand I_24096 (I412911,I413214,I413033);
nand I_24097 (I413245,I1379729,I1379726);
and I_24098 (I413262,I413245,I1379747);
DFFARX1 I_24099 (I413262,I3563,I412934,I413288,);
nor I_24100 (I413296,I413288,I412960);
DFFARX1 I_24101 (I413296,I3563,I412934,I412899,);
DFFARX1 I_24102 (I413288,I3563,I412934,I412917,);
nor I_24103 (I413341,I1379735,I1379726);
not I_24104 (I413358,I413341);
nor I_24105 (I412920,I413197,I413358);
nand I_24106 (I412905,I413214,I413358);
nor I_24107 (I412914,I412960,I413341);
DFFARX1 I_24108 (I413341,I3563,I412934,I412923,);
not I_24109 (I413461,I3570);
DFFARX1 I_24110 (I133592,I3563,I413461,I413487,);
nand I_24111 (I413495,I133604,I133613);
and I_24112 (I413512,I413495,I133592);
DFFARX1 I_24113 (I413512,I3563,I413461,I413538,);
nor I_24114 (I413429,I413538,I413487);
not I_24115 (I413560,I413538);
DFFARX1 I_24116 (I133607,I3563,I413461,I413586,);
nand I_24117 (I413594,I413586,I133595);
not I_24118 (I413611,I413594);
DFFARX1 I_24119 (I413611,I3563,I413461,I413637,);
not I_24120 (I413453,I413637);
nor I_24121 (I413659,I413487,I413594);
nor I_24122 (I413435,I413538,I413659);
DFFARX1 I_24123 (I133598,I3563,I413461,I413699,);
DFFARX1 I_24124 (I413699,I3563,I413461,I413716,);
not I_24125 (I413724,I413716);
not I_24126 (I413741,I413699);
nand I_24127 (I413438,I413741,I413560);
nand I_24128 (I413772,I133589,I133589);
and I_24129 (I413789,I413772,I133601);
DFFARX1 I_24130 (I413789,I3563,I413461,I413815,);
nor I_24131 (I413823,I413815,I413487);
DFFARX1 I_24132 (I413823,I3563,I413461,I413426,);
DFFARX1 I_24133 (I413815,I3563,I413461,I413444,);
nor I_24134 (I413868,I133610,I133589);
not I_24135 (I413885,I413868);
nor I_24136 (I413447,I413724,I413885);
nand I_24137 (I413432,I413741,I413885);
nor I_24138 (I413441,I413487,I413868);
DFFARX1 I_24139 (I413868,I3563,I413461,I413450,);
not I_24140 (I413988,I3570);
DFFARX1 I_24141 (I241658,I3563,I413988,I414014,);
nand I_24142 (I414022,I241658,I241664);
and I_24143 (I414039,I414022,I241682);
DFFARX1 I_24144 (I414039,I3563,I413988,I414065,);
nor I_24145 (I413956,I414065,I414014);
not I_24146 (I414087,I414065);
DFFARX1 I_24147 (I241670,I3563,I413988,I414113,);
nand I_24148 (I414121,I414113,I241667);
not I_24149 (I414138,I414121);
DFFARX1 I_24150 (I414138,I3563,I413988,I414164,);
not I_24151 (I413980,I414164);
nor I_24152 (I414186,I414014,I414121);
nor I_24153 (I413962,I414065,I414186);
DFFARX1 I_24154 (I241676,I3563,I413988,I414226,);
DFFARX1 I_24155 (I414226,I3563,I413988,I414243,);
not I_24156 (I414251,I414243);
not I_24157 (I414268,I414226);
nand I_24158 (I413965,I414268,I414087);
nand I_24159 (I414299,I241661,I241661);
and I_24160 (I414316,I414299,I241673);
DFFARX1 I_24161 (I414316,I3563,I413988,I414342,);
nor I_24162 (I414350,I414342,I414014);
DFFARX1 I_24163 (I414350,I3563,I413988,I413953,);
DFFARX1 I_24164 (I414342,I3563,I413988,I413971,);
nor I_24165 (I414395,I241679,I241661);
not I_24166 (I414412,I414395);
nor I_24167 (I413974,I414251,I414412);
nand I_24168 (I413959,I414268,I414412);
nor I_24169 (I413968,I414014,I414395);
DFFARX1 I_24170 (I414395,I3563,I413988,I413977,);
not I_24171 (I414515,I3570);
DFFARX1 I_24172 (I800613,I3563,I414515,I414541,);
nand I_24173 (I414549,I800604,I800619);
and I_24174 (I414566,I414549,I800625);
DFFARX1 I_24175 (I414566,I3563,I414515,I414592,);
nor I_24176 (I414483,I414592,I414541);
not I_24177 (I414614,I414592);
DFFARX1 I_24178 (I800610,I3563,I414515,I414640,);
nand I_24179 (I414648,I414640,I800604);
not I_24180 (I414665,I414648);
DFFARX1 I_24181 (I414665,I3563,I414515,I414691,);
not I_24182 (I414507,I414691);
nor I_24183 (I414713,I414541,I414648);
nor I_24184 (I414489,I414592,I414713);
DFFARX1 I_24185 (I800607,I3563,I414515,I414753,);
DFFARX1 I_24186 (I414753,I3563,I414515,I414770,);
not I_24187 (I414778,I414770);
not I_24188 (I414795,I414753);
nand I_24189 (I414492,I414795,I414614);
nand I_24190 (I414826,I800601,I800616);
and I_24191 (I414843,I414826,I800601);
DFFARX1 I_24192 (I414843,I3563,I414515,I414869,);
nor I_24193 (I414877,I414869,I414541);
DFFARX1 I_24194 (I414877,I3563,I414515,I414480,);
DFFARX1 I_24195 (I414869,I3563,I414515,I414498,);
nor I_24196 (I414922,I800622,I800616);
not I_24197 (I414939,I414922);
nor I_24198 (I414501,I414778,I414939);
nand I_24199 (I414486,I414795,I414939);
nor I_24200 (I414495,I414541,I414922);
DFFARX1 I_24201 (I414922,I3563,I414515,I414504,);
not I_24202 (I415042,I3570);
DFFARX1 I_24203 (I1284507,I3563,I415042,I415068,);
nand I_24204 (I415076,I1284489,I1284513);
and I_24205 (I415093,I415076,I1284504);
DFFARX1 I_24206 (I415093,I3563,I415042,I415119,);
nor I_24207 (I415010,I415119,I415068);
not I_24208 (I415141,I415119);
DFFARX1 I_24209 (I1284510,I3563,I415042,I415167,);
nand I_24210 (I415175,I415167,I1284498);
not I_24211 (I415192,I415175);
DFFARX1 I_24212 (I415192,I3563,I415042,I415218,);
not I_24213 (I415034,I415218);
nor I_24214 (I415240,I415068,I415175);
nor I_24215 (I415016,I415119,I415240);
DFFARX1 I_24216 (I1284489,I3563,I415042,I415280,);
DFFARX1 I_24217 (I415280,I3563,I415042,I415297,);
not I_24218 (I415305,I415297);
not I_24219 (I415322,I415280);
nand I_24220 (I415019,I415322,I415141);
nand I_24221 (I415353,I1284495,I1284492);
and I_24222 (I415370,I415353,I1284501);
DFFARX1 I_24223 (I415370,I3563,I415042,I415396,);
nor I_24224 (I415404,I415396,I415068);
DFFARX1 I_24225 (I415404,I3563,I415042,I415007,);
DFFARX1 I_24226 (I415396,I3563,I415042,I415025,);
nor I_24227 (I415449,I1284492,I1284492);
not I_24228 (I415466,I415449);
nor I_24229 (I415028,I415305,I415466);
nand I_24230 (I415013,I415322,I415466);
nor I_24231 (I415022,I415068,I415449);
DFFARX1 I_24232 (I415449,I3563,I415042,I415031,);
not I_24233 (I415569,I3570);
DFFARX1 I_24234 (I1190411,I3563,I415569,I415595,);
nand I_24235 (I415603,I1190426,I1190411);
and I_24236 (I415620,I415603,I1190429);
DFFARX1 I_24237 (I415620,I3563,I415569,I415646,);
nor I_24238 (I415537,I415646,I415595);
not I_24239 (I415668,I415646);
DFFARX1 I_24240 (I1190435,I3563,I415569,I415694,);
nand I_24241 (I415702,I415694,I1190417);
not I_24242 (I415719,I415702);
DFFARX1 I_24243 (I415719,I3563,I415569,I415745,);
not I_24244 (I415561,I415745);
nor I_24245 (I415767,I415595,I415702);
nor I_24246 (I415543,I415646,I415767);
DFFARX1 I_24247 (I1190414,I3563,I415569,I415807,);
DFFARX1 I_24248 (I415807,I3563,I415569,I415824,);
not I_24249 (I415832,I415824);
not I_24250 (I415849,I415807);
nand I_24251 (I415546,I415849,I415668);
nand I_24252 (I415880,I1190414,I1190420);
and I_24253 (I415897,I415880,I1190432);
DFFARX1 I_24254 (I415897,I3563,I415569,I415923,);
nor I_24255 (I415931,I415923,I415595);
DFFARX1 I_24256 (I415931,I3563,I415569,I415534,);
DFFARX1 I_24257 (I415923,I3563,I415569,I415552,);
nor I_24258 (I415976,I1190423,I1190420);
not I_24259 (I415993,I415976);
nor I_24260 (I415555,I415832,I415993);
nand I_24261 (I415540,I415849,I415993);
nor I_24262 (I415549,I415595,I415976);
DFFARX1 I_24263 (I415976,I3563,I415569,I415558,);
not I_24264 (I416096,I3570);
DFFARX1 I_24265 (I905392,I3563,I416096,I416122,);
nand I_24266 (I416130,I905395,I905389);
and I_24267 (I416147,I416130,I905401);
DFFARX1 I_24268 (I416147,I3563,I416096,I416173,);
nor I_24269 (I416064,I416173,I416122);
not I_24270 (I416195,I416173);
DFFARX1 I_24271 (I905404,I3563,I416096,I416221,);
nand I_24272 (I416229,I416221,I905395);
not I_24273 (I416246,I416229);
DFFARX1 I_24274 (I416246,I3563,I416096,I416272,);
not I_24275 (I416088,I416272);
nor I_24276 (I416294,I416122,I416229);
nor I_24277 (I416070,I416173,I416294);
DFFARX1 I_24278 (I905407,I3563,I416096,I416334,);
DFFARX1 I_24279 (I416334,I3563,I416096,I416351,);
not I_24280 (I416359,I416351);
not I_24281 (I416376,I416334);
nand I_24282 (I416073,I416376,I416195);
nand I_24283 (I416407,I905389,I905398);
and I_24284 (I416424,I416407,I905392);
DFFARX1 I_24285 (I416424,I3563,I416096,I416450,);
nor I_24286 (I416458,I416450,I416122);
DFFARX1 I_24287 (I416458,I3563,I416096,I416061,);
DFFARX1 I_24288 (I416450,I3563,I416096,I416079,);
nor I_24289 (I416503,I905410,I905398);
not I_24290 (I416520,I416503);
nor I_24291 (I416082,I416359,I416520);
nand I_24292 (I416067,I416376,I416520);
nor I_24293 (I416076,I416122,I416503);
DFFARX1 I_24294 (I416503,I3563,I416096,I416085,);
not I_24295 (I416623,I3570);
DFFARX1 I_24296 (I282118,I3563,I416623,I416649,);
nand I_24297 (I416657,I282118,I282124);
and I_24298 (I416674,I416657,I282142);
DFFARX1 I_24299 (I416674,I3563,I416623,I416700,);
nor I_24300 (I416591,I416700,I416649);
not I_24301 (I416722,I416700);
DFFARX1 I_24302 (I282130,I3563,I416623,I416748,);
nand I_24303 (I416756,I416748,I282127);
not I_24304 (I416773,I416756);
DFFARX1 I_24305 (I416773,I3563,I416623,I416799,);
not I_24306 (I416615,I416799);
nor I_24307 (I416821,I416649,I416756);
nor I_24308 (I416597,I416700,I416821);
DFFARX1 I_24309 (I282136,I3563,I416623,I416861,);
DFFARX1 I_24310 (I416861,I3563,I416623,I416878,);
not I_24311 (I416886,I416878);
not I_24312 (I416903,I416861);
nand I_24313 (I416600,I416903,I416722);
nand I_24314 (I416934,I282121,I282121);
and I_24315 (I416951,I416934,I282133);
DFFARX1 I_24316 (I416951,I3563,I416623,I416977,);
nor I_24317 (I416985,I416977,I416649);
DFFARX1 I_24318 (I416985,I3563,I416623,I416588,);
DFFARX1 I_24319 (I416977,I3563,I416623,I416606,);
nor I_24320 (I417030,I282139,I282121);
not I_24321 (I417047,I417030);
nor I_24322 (I416609,I416886,I417047);
nand I_24323 (I416594,I416903,I417047);
nor I_24324 (I416603,I416649,I417030);
DFFARX1 I_24325 (I417030,I3563,I416623,I416612,);
not I_24326 (I417150,I3570);
DFFARX1 I_24327 (I1147639,I3563,I417150,I417176,);
nand I_24328 (I417184,I1147654,I1147639);
and I_24329 (I417201,I417184,I1147657);
DFFARX1 I_24330 (I417201,I3563,I417150,I417227,);
nor I_24331 (I417118,I417227,I417176);
not I_24332 (I417249,I417227);
DFFARX1 I_24333 (I1147663,I3563,I417150,I417275,);
nand I_24334 (I417283,I417275,I1147645);
not I_24335 (I417300,I417283);
DFFARX1 I_24336 (I417300,I3563,I417150,I417326,);
not I_24337 (I417142,I417326);
nor I_24338 (I417348,I417176,I417283);
nor I_24339 (I417124,I417227,I417348);
DFFARX1 I_24340 (I1147642,I3563,I417150,I417388,);
DFFARX1 I_24341 (I417388,I3563,I417150,I417405,);
not I_24342 (I417413,I417405);
not I_24343 (I417430,I417388);
nand I_24344 (I417127,I417430,I417249);
nand I_24345 (I417461,I1147642,I1147648);
and I_24346 (I417478,I417461,I1147660);
DFFARX1 I_24347 (I417478,I3563,I417150,I417504,);
nor I_24348 (I417512,I417504,I417176);
DFFARX1 I_24349 (I417512,I3563,I417150,I417115,);
DFFARX1 I_24350 (I417504,I3563,I417150,I417133,);
nor I_24351 (I417557,I1147651,I1147648);
not I_24352 (I417574,I417557);
nor I_24353 (I417136,I417413,I417574);
nand I_24354 (I417121,I417430,I417574);
nor I_24355 (I417130,I417176,I417557);
DFFARX1 I_24356 (I417557,I3563,I417150,I417139,);
not I_24357 (I417677,I3570);
DFFARX1 I_24358 (I586756,I3563,I417677,I417703,);
nand I_24359 (I417711,I586741,I586744);
and I_24360 (I417728,I417711,I586759);
DFFARX1 I_24361 (I417728,I3563,I417677,I417754,);
nor I_24362 (I417645,I417754,I417703);
not I_24363 (I417776,I417754);
DFFARX1 I_24364 (I586753,I3563,I417677,I417802,);
nand I_24365 (I417810,I417802,I586744);
not I_24366 (I417827,I417810);
DFFARX1 I_24367 (I417827,I3563,I417677,I417853,);
not I_24368 (I417669,I417853);
nor I_24369 (I417875,I417703,I417810);
nor I_24370 (I417651,I417754,I417875);
DFFARX1 I_24371 (I586750,I3563,I417677,I417915,);
DFFARX1 I_24372 (I417915,I3563,I417677,I417932,);
not I_24373 (I417940,I417932);
not I_24374 (I417957,I417915);
nand I_24375 (I417654,I417957,I417776);
nand I_24376 (I417988,I586765,I586741);
and I_24377 (I418005,I417988,I586762);
DFFARX1 I_24378 (I418005,I3563,I417677,I418031,);
nor I_24379 (I418039,I418031,I417703);
DFFARX1 I_24380 (I418039,I3563,I417677,I417642,);
DFFARX1 I_24381 (I418031,I3563,I417677,I417660,);
nor I_24382 (I418084,I586747,I586741);
not I_24383 (I418101,I418084);
nor I_24384 (I417663,I417940,I418101);
nand I_24385 (I417648,I417957,I418101);
nor I_24386 (I417657,I417703,I418084);
DFFARX1 I_24387 (I418084,I3563,I417677,I417666,);
not I_24388 (I418204,I3570);
DFFARX1 I_24389 (I1357729,I3563,I418204,I418230,);
nand I_24390 (I418238,I1357708,I1357708);
and I_24391 (I418255,I418238,I1357735);
DFFARX1 I_24392 (I418255,I3563,I418204,I418281,);
nor I_24393 (I418172,I418281,I418230);
not I_24394 (I418303,I418281);
DFFARX1 I_24395 (I1357723,I3563,I418204,I418329,);
nand I_24396 (I418337,I418329,I1357726);
not I_24397 (I418354,I418337);
DFFARX1 I_24398 (I418354,I3563,I418204,I418380,);
not I_24399 (I418196,I418380);
nor I_24400 (I418402,I418230,I418337);
nor I_24401 (I418178,I418281,I418402);
DFFARX1 I_24402 (I1357717,I3563,I418204,I418442,);
DFFARX1 I_24403 (I418442,I3563,I418204,I418459,);
not I_24404 (I418467,I418459);
not I_24405 (I418484,I418442);
nand I_24406 (I418181,I418484,I418303);
nand I_24407 (I418515,I1357714,I1357711);
and I_24408 (I418532,I418515,I1357732);
DFFARX1 I_24409 (I418532,I3563,I418204,I418558,);
nor I_24410 (I418566,I418558,I418230);
DFFARX1 I_24411 (I418566,I3563,I418204,I418169,);
DFFARX1 I_24412 (I418558,I3563,I418204,I418187,);
nor I_24413 (I418611,I1357720,I1357711);
not I_24414 (I418628,I418611);
nor I_24415 (I418190,I418467,I418628);
nand I_24416 (I418175,I418484,I418628);
nor I_24417 (I418184,I418230,I418611);
DFFARX1 I_24418 (I418611,I3563,I418204,I418193,);
not I_24419 (I418731,I3570);
DFFARX1 I_24420 (I842152,I3563,I418731,I418757,);
nand I_24421 (I418765,I842155,I842149);
and I_24422 (I418782,I418765,I842161);
DFFARX1 I_24423 (I418782,I3563,I418731,I418808,);
nor I_24424 (I418699,I418808,I418757);
not I_24425 (I418830,I418808);
DFFARX1 I_24426 (I842164,I3563,I418731,I418856,);
nand I_24427 (I418864,I418856,I842155);
not I_24428 (I418881,I418864);
DFFARX1 I_24429 (I418881,I3563,I418731,I418907,);
not I_24430 (I418723,I418907);
nor I_24431 (I418929,I418757,I418864);
nor I_24432 (I418705,I418808,I418929);
DFFARX1 I_24433 (I842167,I3563,I418731,I418969,);
DFFARX1 I_24434 (I418969,I3563,I418731,I418986,);
not I_24435 (I418994,I418986);
not I_24436 (I419011,I418969);
nand I_24437 (I418708,I419011,I418830);
nand I_24438 (I419042,I842149,I842158);
and I_24439 (I419059,I419042,I842152);
DFFARX1 I_24440 (I419059,I3563,I418731,I419085,);
nor I_24441 (I419093,I419085,I418757);
DFFARX1 I_24442 (I419093,I3563,I418731,I418696,);
DFFARX1 I_24443 (I419085,I3563,I418731,I418714,);
nor I_24444 (I419138,I842170,I842158);
not I_24445 (I419155,I419138);
nor I_24446 (I418717,I418994,I419155);
nand I_24447 (I418702,I419011,I419155);
nor I_24448 (I418711,I418757,I419138);
DFFARX1 I_24449 (I419138,I3563,I418731,I418720,);
not I_24450 (I419258,I3570);
DFFARX1 I_24451 (I1348804,I3563,I419258,I419284,);
nand I_24452 (I419292,I1348783,I1348783);
and I_24453 (I419309,I419292,I1348810);
DFFARX1 I_24454 (I419309,I3563,I419258,I419335,);
nor I_24455 (I419226,I419335,I419284);
not I_24456 (I419357,I419335);
DFFARX1 I_24457 (I1348798,I3563,I419258,I419383,);
nand I_24458 (I419391,I419383,I1348801);
not I_24459 (I419408,I419391);
DFFARX1 I_24460 (I419408,I3563,I419258,I419434,);
not I_24461 (I419250,I419434);
nor I_24462 (I419456,I419284,I419391);
nor I_24463 (I419232,I419335,I419456);
DFFARX1 I_24464 (I1348792,I3563,I419258,I419496,);
DFFARX1 I_24465 (I419496,I3563,I419258,I419513,);
not I_24466 (I419521,I419513);
not I_24467 (I419538,I419496);
nand I_24468 (I419235,I419538,I419357);
nand I_24469 (I419569,I1348789,I1348786);
and I_24470 (I419586,I419569,I1348807);
DFFARX1 I_24471 (I419586,I3563,I419258,I419612,);
nor I_24472 (I419620,I419612,I419284);
DFFARX1 I_24473 (I419620,I3563,I419258,I419223,);
DFFARX1 I_24474 (I419612,I3563,I419258,I419241,);
nor I_24475 (I419665,I1348795,I1348786);
not I_24476 (I419682,I419665);
nor I_24477 (I419244,I419521,I419682);
nand I_24478 (I419229,I419538,I419682);
nor I_24479 (I419238,I419284,I419665);
DFFARX1 I_24480 (I419665,I3563,I419258,I419247,);
not I_24481 (I419785,I3570);
DFFARX1 I_24482 (I85635,I3563,I419785,I419811,);
nand I_24483 (I419819,I85647,I85656);
and I_24484 (I419836,I419819,I85635);
DFFARX1 I_24485 (I419836,I3563,I419785,I419862,);
nor I_24486 (I419753,I419862,I419811);
not I_24487 (I419884,I419862);
DFFARX1 I_24488 (I85650,I3563,I419785,I419910,);
nand I_24489 (I419918,I419910,I85638);
not I_24490 (I419935,I419918);
DFFARX1 I_24491 (I419935,I3563,I419785,I419961,);
not I_24492 (I419777,I419961);
nor I_24493 (I419983,I419811,I419918);
nor I_24494 (I419759,I419862,I419983);
DFFARX1 I_24495 (I85641,I3563,I419785,I420023,);
DFFARX1 I_24496 (I420023,I3563,I419785,I420040,);
not I_24497 (I420048,I420040);
not I_24498 (I420065,I420023);
nand I_24499 (I419762,I420065,I419884);
nand I_24500 (I420096,I85632,I85632);
and I_24501 (I420113,I420096,I85644);
DFFARX1 I_24502 (I420113,I3563,I419785,I420139,);
nor I_24503 (I420147,I420139,I419811);
DFFARX1 I_24504 (I420147,I3563,I419785,I419750,);
DFFARX1 I_24505 (I420139,I3563,I419785,I419768,);
nor I_24506 (I420192,I85653,I85632);
not I_24507 (I420209,I420192);
nor I_24508 (I419771,I420048,I420209);
nand I_24509 (I419756,I420065,I420209);
nor I_24510 (I419765,I419811,I420192);
DFFARX1 I_24511 (I420192,I3563,I419785,I419774,);
not I_24512 (I420312,I3570);
DFFARX1 I_24513 (I78257,I3563,I420312,I420338,);
nand I_24514 (I420346,I78269,I78278);
and I_24515 (I420363,I420346,I78257);
DFFARX1 I_24516 (I420363,I3563,I420312,I420389,);
nor I_24517 (I420280,I420389,I420338);
not I_24518 (I420411,I420389);
DFFARX1 I_24519 (I78272,I3563,I420312,I420437,);
nand I_24520 (I420445,I420437,I78260);
not I_24521 (I420462,I420445);
DFFARX1 I_24522 (I420462,I3563,I420312,I420488,);
not I_24523 (I420304,I420488);
nor I_24524 (I420510,I420338,I420445);
nor I_24525 (I420286,I420389,I420510);
DFFARX1 I_24526 (I78263,I3563,I420312,I420550,);
DFFARX1 I_24527 (I420550,I3563,I420312,I420567,);
not I_24528 (I420575,I420567);
not I_24529 (I420592,I420550);
nand I_24530 (I420289,I420592,I420411);
nand I_24531 (I420623,I78254,I78254);
and I_24532 (I420640,I420623,I78266);
DFFARX1 I_24533 (I420640,I3563,I420312,I420666,);
nor I_24534 (I420674,I420666,I420338);
DFFARX1 I_24535 (I420674,I3563,I420312,I420277,);
DFFARX1 I_24536 (I420666,I3563,I420312,I420295,);
nor I_24537 (I420719,I78275,I78254);
not I_24538 (I420736,I420719);
nor I_24539 (I420298,I420575,I420736);
nand I_24540 (I420283,I420592,I420736);
nor I_24541 (I420292,I420338,I420719);
DFFARX1 I_24542 (I420719,I3563,I420312,I420301,);
not I_24543 (I420839,I3570);
DFFARX1 I_24544 (I672297,I3563,I420839,I420865,);
nand I_24545 (I420873,I672288,I672303);
and I_24546 (I420890,I420873,I672309);
DFFARX1 I_24547 (I420890,I3563,I420839,I420916,);
nor I_24548 (I420807,I420916,I420865);
not I_24549 (I420938,I420916);
DFFARX1 I_24550 (I672294,I3563,I420839,I420964,);
nand I_24551 (I420972,I420964,I672288);
not I_24552 (I420989,I420972);
DFFARX1 I_24553 (I420989,I3563,I420839,I421015,);
not I_24554 (I420831,I421015);
nor I_24555 (I421037,I420865,I420972);
nor I_24556 (I420813,I420916,I421037);
DFFARX1 I_24557 (I672291,I3563,I420839,I421077,);
DFFARX1 I_24558 (I421077,I3563,I420839,I421094,);
not I_24559 (I421102,I421094);
not I_24560 (I421119,I421077);
nand I_24561 (I420816,I421119,I420938);
nand I_24562 (I421150,I672285,I672300);
and I_24563 (I421167,I421150,I672285);
DFFARX1 I_24564 (I421167,I3563,I420839,I421193,);
nor I_24565 (I421201,I421193,I420865);
DFFARX1 I_24566 (I421201,I3563,I420839,I420804,);
DFFARX1 I_24567 (I421193,I3563,I420839,I420822,);
nor I_24568 (I421246,I672306,I672300);
not I_24569 (I421263,I421246);
nor I_24570 (I420825,I421102,I421263);
nand I_24571 (I420810,I421119,I421263);
nor I_24572 (I420819,I420865,I421246);
DFFARX1 I_24573 (I421246,I3563,I420839,I420828,);
not I_24574 (I421366,I3570);
DFFARX1 I_24575 (I260103,I3563,I421366,I421392,);
nand I_24576 (I421400,I260103,I260109);
and I_24577 (I421417,I421400,I260127);
DFFARX1 I_24578 (I421417,I3563,I421366,I421443,);
nor I_24579 (I421334,I421443,I421392);
not I_24580 (I421465,I421443);
DFFARX1 I_24581 (I260115,I3563,I421366,I421491,);
nand I_24582 (I421499,I421491,I260112);
not I_24583 (I421516,I421499);
DFFARX1 I_24584 (I421516,I3563,I421366,I421542,);
not I_24585 (I421358,I421542);
nor I_24586 (I421564,I421392,I421499);
nor I_24587 (I421340,I421443,I421564);
DFFARX1 I_24588 (I260121,I3563,I421366,I421604,);
DFFARX1 I_24589 (I421604,I3563,I421366,I421621,);
not I_24590 (I421629,I421621);
not I_24591 (I421646,I421604);
nand I_24592 (I421343,I421646,I421465);
nand I_24593 (I421677,I260106,I260106);
and I_24594 (I421694,I421677,I260118);
DFFARX1 I_24595 (I421694,I3563,I421366,I421720,);
nor I_24596 (I421728,I421720,I421392);
DFFARX1 I_24597 (I421728,I3563,I421366,I421331,);
DFFARX1 I_24598 (I421720,I3563,I421366,I421349,);
nor I_24599 (I421773,I260124,I260106);
not I_24600 (I421790,I421773);
nor I_24601 (I421352,I421629,I421790);
nand I_24602 (I421337,I421646,I421790);
nor I_24603 (I421346,I421392,I421773);
DFFARX1 I_24604 (I421773,I3563,I421366,I421355,);
not I_24605 (I421893,I3570);
DFFARX1 I_24606 (I290129,I3563,I421893,I421919,);
DFFARX1 I_24607 (I421919,I3563,I421893,I421936,);
not I_24608 (I421885,I421936);
not I_24609 (I421958,I421919);
nand I_24610 (I421975,I290108,I290132);
and I_24611 (I421992,I421975,I290135);
DFFARX1 I_24612 (I421992,I3563,I421893,I422018,);
not I_24613 (I422026,I422018);
DFFARX1 I_24614 (I290117,I3563,I421893,I422052,);
and I_24615 (I422060,I422052,I290123);
nand I_24616 (I422077,I422052,I290123);
nand I_24617 (I421864,I422026,I422077);
DFFARX1 I_24618 (I290111,I3563,I421893,I422117,);
nor I_24619 (I422125,I422117,I422060);
DFFARX1 I_24620 (I422125,I3563,I421893,I421858,);
nor I_24621 (I421873,I422117,I422018);
nand I_24622 (I422170,I290120,I290108);
and I_24623 (I422187,I422170,I290114);
DFFARX1 I_24624 (I422187,I3563,I421893,I422213,);
nor I_24625 (I421861,I422213,I422117);
not I_24626 (I422235,I422213);
nor I_24627 (I422252,I422235,I422026);
nor I_24628 (I422269,I421958,I422252);
DFFARX1 I_24629 (I422269,I3563,I421893,I421876,);
nor I_24630 (I422300,I422235,I422117);
nor I_24631 (I422317,I290126,I290108);
nor I_24632 (I421867,I422317,I422300);
not I_24633 (I422348,I422317);
nand I_24634 (I421870,I422077,I422348);
DFFARX1 I_24635 (I422317,I3563,I421893,I421882,);
DFFARX1 I_24636 (I422317,I3563,I421893,I421879,);
not I_24637 (I422437,I3570);
DFFARX1 I_24638 (I921987,I3563,I422437,I422463,);
DFFARX1 I_24639 (I422463,I3563,I422437,I422480,);
not I_24640 (I422429,I422480);
not I_24641 (I422502,I422463);
nand I_24642 (I422519,I922002,I921990);
and I_24643 (I422536,I422519,I921981);
DFFARX1 I_24644 (I422536,I3563,I422437,I422562,);
not I_24645 (I422570,I422562);
DFFARX1 I_24646 (I921993,I3563,I422437,I422596,);
and I_24647 (I422604,I422596,I921984);
nand I_24648 (I422621,I422596,I921984);
nand I_24649 (I422408,I422570,I422621);
DFFARX1 I_24650 (I921999,I3563,I422437,I422661,);
nor I_24651 (I422669,I422661,I422604);
DFFARX1 I_24652 (I422669,I3563,I422437,I422402,);
nor I_24653 (I422417,I422661,I422562);
nand I_24654 (I422714,I922008,I921996);
and I_24655 (I422731,I422714,I922005);
DFFARX1 I_24656 (I422731,I3563,I422437,I422757,);
nor I_24657 (I422405,I422757,I422661);
not I_24658 (I422779,I422757);
nor I_24659 (I422796,I422779,I422570);
nor I_24660 (I422813,I422502,I422796);
DFFARX1 I_24661 (I422813,I3563,I422437,I422420,);
nor I_24662 (I422844,I422779,I422661);
nor I_24663 (I422861,I921981,I921996);
nor I_24664 (I422411,I422861,I422844);
not I_24665 (I422892,I422861);
nand I_24666 (I422414,I422621,I422892);
DFFARX1 I_24667 (I422861,I3563,I422437,I422426,);
DFFARX1 I_24668 (I422861,I3563,I422437,I422423,);
not I_24669 (I422981,I3570);
DFFARX1 I_24670 (I728932,I3563,I422981,I423007,);
DFFARX1 I_24671 (I423007,I3563,I422981,I423024,);
not I_24672 (I422973,I423024);
not I_24673 (I423046,I423007);
nand I_24674 (I423063,I728953,I728944);
and I_24675 (I423080,I423063,I728932);
DFFARX1 I_24676 (I423080,I3563,I422981,I423106,);
not I_24677 (I423114,I423106);
DFFARX1 I_24678 (I728938,I3563,I422981,I423140,);
and I_24679 (I423148,I423140,I728935);
nand I_24680 (I423165,I423140,I728935);
nand I_24681 (I422952,I423114,I423165);
DFFARX1 I_24682 (I728929,I3563,I422981,I423205,);
nor I_24683 (I423213,I423205,I423148);
DFFARX1 I_24684 (I423213,I3563,I422981,I422946,);
nor I_24685 (I422961,I423205,I423106);
nand I_24686 (I423258,I728929,I728941);
and I_24687 (I423275,I423258,I728950);
DFFARX1 I_24688 (I423275,I3563,I422981,I423301,);
nor I_24689 (I422949,I423301,I423205);
not I_24690 (I423323,I423301);
nor I_24691 (I423340,I423323,I423114);
nor I_24692 (I423357,I423046,I423340);
DFFARX1 I_24693 (I423357,I3563,I422981,I422964,);
nor I_24694 (I423388,I423323,I423205);
nor I_24695 (I423405,I728947,I728941);
nor I_24696 (I422955,I423405,I423388);
not I_24697 (I423436,I423405);
nand I_24698 (I422958,I423165,I423436);
DFFARX1 I_24699 (I423405,I3563,I422981,I422970,);
DFFARX1 I_24700 (I423405,I3563,I422981,I422967,);
not I_24701 (I423525,I3570);
DFFARX1 I_24702 (I381300,I3563,I423525,I423551,);
DFFARX1 I_24703 (I423551,I3563,I423525,I423568,);
not I_24704 (I423517,I423568);
not I_24705 (I423590,I423551);
nand I_24706 (I423607,I381279,I381303);
and I_24707 (I423624,I423607,I381306);
DFFARX1 I_24708 (I423624,I3563,I423525,I423650,);
not I_24709 (I423658,I423650);
DFFARX1 I_24710 (I381288,I3563,I423525,I423684,);
and I_24711 (I423692,I423684,I381294);
nand I_24712 (I423709,I423684,I381294);
nand I_24713 (I423496,I423658,I423709);
DFFARX1 I_24714 (I381282,I3563,I423525,I423749,);
nor I_24715 (I423757,I423749,I423692);
DFFARX1 I_24716 (I423757,I3563,I423525,I423490,);
nor I_24717 (I423505,I423749,I423650);
nand I_24718 (I423802,I381291,I381279);
and I_24719 (I423819,I423802,I381285);
DFFARX1 I_24720 (I423819,I3563,I423525,I423845,);
nor I_24721 (I423493,I423845,I423749);
not I_24722 (I423867,I423845);
nor I_24723 (I423884,I423867,I423658);
nor I_24724 (I423901,I423590,I423884);
DFFARX1 I_24725 (I423901,I3563,I423525,I423508,);
nor I_24726 (I423932,I423867,I423749);
nor I_24727 (I423949,I381297,I381279);
nor I_24728 (I423499,I423949,I423932);
not I_24729 (I423980,I423949);
nand I_24730 (I423502,I423709,I423980);
DFFARX1 I_24731 (I423949,I3563,I423525,I423514,);
DFFARX1 I_24732 (I423949,I3563,I423525,I423511,);
not I_24733 (I424069,I3570);
DFFARX1 I_24734 (I308047,I3563,I424069,I424095,);
DFFARX1 I_24735 (I424095,I3563,I424069,I424112,);
not I_24736 (I424061,I424112);
not I_24737 (I424134,I424095);
nand I_24738 (I424151,I308026,I308050);
and I_24739 (I424168,I424151,I308053);
DFFARX1 I_24740 (I424168,I3563,I424069,I424194,);
not I_24741 (I424202,I424194);
DFFARX1 I_24742 (I308035,I3563,I424069,I424228,);
and I_24743 (I424236,I424228,I308041);
nand I_24744 (I424253,I424228,I308041);
nand I_24745 (I424040,I424202,I424253);
DFFARX1 I_24746 (I308029,I3563,I424069,I424293,);
nor I_24747 (I424301,I424293,I424236);
DFFARX1 I_24748 (I424301,I3563,I424069,I424034,);
nor I_24749 (I424049,I424293,I424194);
nand I_24750 (I424346,I308038,I308026);
and I_24751 (I424363,I424346,I308032);
DFFARX1 I_24752 (I424363,I3563,I424069,I424389,);
nor I_24753 (I424037,I424389,I424293);
not I_24754 (I424411,I424389);
nor I_24755 (I424428,I424411,I424202);
nor I_24756 (I424445,I424134,I424428);
DFFARX1 I_24757 (I424445,I3563,I424069,I424052,);
nor I_24758 (I424476,I424411,I424293);
nor I_24759 (I424493,I308044,I308026);
nor I_24760 (I424043,I424493,I424476);
not I_24761 (I424524,I424493);
nand I_24762 (I424046,I424253,I424524);
DFFARX1 I_24763 (I424493,I3563,I424069,I424058,);
DFFARX1 I_24764 (I424493,I3563,I424069,I424055,);
not I_24765 (I424613,I3570);
DFFARX1 I_24766 (I1149376,I3563,I424613,I424639,);
DFFARX1 I_24767 (I424639,I3563,I424613,I424656,);
not I_24768 (I424605,I424656);
not I_24769 (I424678,I424639);
nand I_24770 (I424695,I1149388,I1149376);
and I_24771 (I424712,I424695,I1149379);
DFFARX1 I_24772 (I424712,I3563,I424613,I424738,);
not I_24773 (I424746,I424738);
DFFARX1 I_24774 (I1149397,I3563,I424613,I424772,);
and I_24775 (I424780,I424772,I1149373);
nand I_24776 (I424797,I424772,I1149373);
nand I_24777 (I424584,I424746,I424797);
DFFARX1 I_24778 (I1149391,I3563,I424613,I424837,);
nor I_24779 (I424845,I424837,I424780);
DFFARX1 I_24780 (I424845,I3563,I424613,I424578,);
nor I_24781 (I424593,I424837,I424738);
nand I_24782 (I424890,I1149385,I1149382);
and I_24783 (I424907,I424890,I1149394);
DFFARX1 I_24784 (I424907,I3563,I424613,I424933,);
nor I_24785 (I424581,I424933,I424837);
not I_24786 (I424955,I424933);
nor I_24787 (I424972,I424955,I424746);
nor I_24788 (I424989,I424678,I424972);
DFFARX1 I_24789 (I424989,I3563,I424613,I424596,);
nor I_24790 (I425020,I424955,I424837);
nor I_24791 (I425037,I1149373,I1149382);
nor I_24792 (I424587,I425037,I425020);
not I_24793 (I425068,I425037);
nand I_24794 (I424590,I424797,I425068);
DFFARX1 I_24795 (I425037,I3563,I424613,I424602,);
DFFARX1 I_24796 (I425037,I3563,I424613,I424599,);
not I_24797 (I425157,I3570);
DFFARX1 I_24798 (I885902,I3563,I425157,I425183,);
DFFARX1 I_24799 (I425183,I3563,I425157,I425200,);
not I_24800 (I425149,I425200);
not I_24801 (I425222,I425183);
nand I_24802 (I425239,I885896,I885893);
and I_24803 (I425256,I425239,I885908);
DFFARX1 I_24804 (I425256,I3563,I425157,I425282,);
not I_24805 (I425290,I425282);
DFFARX1 I_24806 (I885896,I3563,I425157,I425316,);
and I_24807 (I425324,I425316,I885890);
nand I_24808 (I425341,I425316,I885890);
nand I_24809 (I425128,I425290,I425341);
DFFARX1 I_24810 (I885890,I3563,I425157,I425381,);
nor I_24811 (I425389,I425381,I425324);
DFFARX1 I_24812 (I425389,I3563,I425157,I425122,);
nor I_24813 (I425137,I425381,I425282);
nand I_24814 (I425434,I885905,I885899);
and I_24815 (I425451,I425434,I885893);
DFFARX1 I_24816 (I425451,I3563,I425157,I425477,);
nor I_24817 (I425125,I425477,I425381);
not I_24818 (I425499,I425477);
nor I_24819 (I425516,I425499,I425290);
nor I_24820 (I425533,I425222,I425516);
DFFARX1 I_24821 (I425533,I3563,I425157,I425140,);
nor I_24822 (I425564,I425499,I425381);
nor I_24823 (I425581,I885911,I885899);
nor I_24824 (I425131,I425581,I425564);
not I_24825 (I425612,I425581);
nand I_24826 (I425134,I425341,I425612);
DFFARX1 I_24827 (I425581,I3563,I425157,I425146,);
DFFARX1 I_24828 (I425581,I3563,I425157,I425143,);
not I_24829 (I425701,I3570);
DFFARX1 I_24830 (I153621,I3563,I425701,I425727,);
DFFARX1 I_24831 (I425727,I3563,I425701,I425744,);
not I_24832 (I425693,I425744);
not I_24833 (I425766,I425727);
nand I_24834 (I425783,I153636,I153615);
and I_24835 (I425800,I425783,I153618);
DFFARX1 I_24836 (I425800,I3563,I425701,I425826,);
not I_24837 (I425834,I425826);
DFFARX1 I_24838 (I153624,I3563,I425701,I425860,);
and I_24839 (I425868,I425860,I153618);
nand I_24840 (I425885,I425860,I153618);
nand I_24841 (I425672,I425834,I425885);
DFFARX1 I_24842 (I153633,I3563,I425701,I425925,);
nor I_24843 (I425933,I425925,I425868);
DFFARX1 I_24844 (I425933,I3563,I425701,I425666,);
nor I_24845 (I425681,I425925,I425826);
nand I_24846 (I425978,I153615,I153630);
and I_24847 (I425995,I425978,I153627);
DFFARX1 I_24848 (I425995,I3563,I425701,I426021,);
nor I_24849 (I425669,I426021,I425925);
not I_24850 (I426043,I426021);
nor I_24851 (I426060,I426043,I425834);
nor I_24852 (I426077,I425766,I426060);
DFFARX1 I_24853 (I426077,I3563,I425701,I425684,);
nor I_24854 (I426108,I426043,I425925);
nor I_24855 (I426125,I153639,I153630);
nor I_24856 (I425675,I426125,I426108);
not I_24857 (I426156,I426125);
nand I_24858 (I425678,I425885,I426156);
DFFARX1 I_24859 (I426125,I3563,I425701,I425690,);
DFFARX1 I_24860 (I426125,I3563,I425701,I425687,);
not I_24861 (I426245,I3570);
DFFARX1 I_24862 (I1382130,I3563,I426245,I426271,);
DFFARX1 I_24863 (I426271,I3563,I426245,I426288,);
not I_24864 (I426237,I426288);
not I_24865 (I426310,I426271);
nand I_24866 (I426327,I1382106,I1382127);
and I_24867 (I426344,I426327,I1382124);
DFFARX1 I_24868 (I426344,I3563,I426245,I426370,);
not I_24869 (I426378,I426370);
DFFARX1 I_24870 (I1382103,I3563,I426245,I426404,);
and I_24871 (I426412,I426404,I1382115);
nand I_24872 (I426429,I426404,I1382115);
nand I_24873 (I426216,I426378,I426429);
DFFARX1 I_24874 (I1382118,I3563,I426245,I426469,);
nor I_24875 (I426477,I426469,I426412);
DFFARX1 I_24876 (I426477,I3563,I426245,I426210,);
nor I_24877 (I426225,I426469,I426370);
nand I_24878 (I426522,I1382121,I1382109);
and I_24879 (I426539,I426522,I1382112);
DFFARX1 I_24880 (I426539,I3563,I426245,I426565,);
nor I_24881 (I426213,I426565,I426469);
not I_24882 (I426587,I426565);
nor I_24883 (I426604,I426587,I426378);
nor I_24884 (I426621,I426310,I426604);
DFFARX1 I_24885 (I426621,I3563,I426245,I426228,);
nor I_24886 (I426652,I426587,I426469);
nor I_24887 (I426669,I1382103,I1382109);
nor I_24888 (I426219,I426669,I426652);
not I_24889 (I426700,I426669);
nand I_24890 (I426222,I426429,I426700);
DFFARX1 I_24891 (I426669,I3563,I426245,I426234,);
DFFARX1 I_24892 (I426669,I3563,I426245,I426231,);
not I_24893 (I426789,I3570);
DFFARX1 I_24894 (I820027,I3563,I426789,I426815,);
DFFARX1 I_24895 (I426815,I3563,I426789,I426832,);
not I_24896 (I426781,I426832);
not I_24897 (I426854,I426815);
nand I_24898 (I426871,I820021,I820018);
and I_24899 (I426888,I426871,I820033);
DFFARX1 I_24900 (I426888,I3563,I426789,I426914,);
not I_24901 (I426922,I426914);
DFFARX1 I_24902 (I820021,I3563,I426789,I426948,);
and I_24903 (I426956,I426948,I820015);
nand I_24904 (I426973,I426948,I820015);
nand I_24905 (I426760,I426922,I426973);
DFFARX1 I_24906 (I820015,I3563,I426789,I427013,);
nor I_24907 (I427021,I427013,I426956);
DFFARX1 I_24908 (I427021,I3563,I426789,I426754,);
nor I_24909 (I426769,I427013,I426914);
nand I_24910 (I427066,I820030,I820024);
and I_24911 (I427083,I427066,I820018);
DFFARX1 I_24912 (I427083,I3563,I426789,I427109,);
nor I_24913 (I426757,I427109,I427013);
not I_24914 (I427131,I427109);
nor I_24915 (I427148,I427131,I426922);
nor I_24916 (I427165,I426854,I427148);
DFFARX1 I_24917 (I427165,I3563,I426789,I426772,);
nor I_24918 (I427196,I427131,I427013);
nor I_24919 (I427213,I820036,I820024);
nor I_24920 (I426763,I427213,I427196);
not I_24921 (I427244,I427213);
nand I_24922 (I426766,I426973,I427244);
DFFARX1 I_24923 (I427213,I3563,I426789,I426778,);
DFFARX1 I_24924 (I427213,I3563,I426789,I426775,);
not I_24925 (I427333,I3570);
DFFARX1 I_24926 (I752052,I3563,I427333,I427359,);
DFFARX1 I_24927 (I427359,I3563,I427333,I427376,);
not I_24928 (I427325,I427376);
not I_24929 (I427398,I427359);
nand I_24930 (I427415,I752073,I752064);
and I_24931 (I427432,I427415,I752052);
DFFARX1 I_24932 (I427432,I3563,I427333,I427458,);
not I_24933 (I427466,I427458);
DFFARX1 I_24934 (I752058,I3563,I427333,I427492,);
and I_24935 (I427500,I427492,I752055);
nand I_24936 (I427517,I427492,I752055);
nand I_24937 (I427304,I427466,I427517);
DFFARX1 I_24938 (I752049,I3563,I427333,I427557,);
nor I_24939 (I427565,I427557,I427500);
DFFARX1 I_24940 (I427565,I3563,I427333,I427298,);
nor I_24941 (I427313,I427557,I427458);
nand I_24942 (I427610,I752049,I752061);
and I_24943 (I427627,I427610,I752070);
DFFARX1 I_24944 (I427627,I3563,I427333,I427653,);
nor I_24945 (I427301,I427653,I427557);
not I_24946 (I427675,I427653);
nor I_24947 (I427692,I427675,I427466);
nor I_24948 (I427709,I427398,I427692);
DFFARX1 I_24949 (I427709,I3563,I427333,I427316,);
nor I_24950 (I427740,I427675,I427557);
nor I_24951 (I427757,I752067,I752061);
nor I_24952 (I427307,I427757,I427740);
not I_24953 (I427788,I427757);
nand I_24954 (I427310,I427517,I427788);
DFFARX1 I_24955 (I427757,I3563,I427333,I427322,);
DFFARX1 I_24956 (I427757,I3563,I427333,I427319,);
not I_24957 (I427877,I3570);
DFFARX1 I_24958 (I1095044,I3563,I427877,I427903,);
DFFARX1 I_24959 (I427903,I3563,I427877,I427920,);
not I_24960 (I427869,I427920);
not I_24961 (I427942,I427903);
nand I_24962 (I427959,I1095056,I1095044);
and I_24963 (I427976,I427959,I1095047);
DFFARX1 I_24964 (I427976,I3563,I427877,I428002,);
not I_24965 (I428010,I428002);
DFFARX1 I_24966 (I1095065,I3563,I427877,I428036,);
and I_24967 (I428044,I428036,I1095041);
nand I_24968 (I428061,I428036,I1095041);
nand I_24969 (I427848,I428010,I428061);
DFFARX1 I_24970 (I1095059,I3563,I427877,I428101,);
nor I_24971 (I428109,I428101,I428044);
DFFARX1 I_24972 (I428109,I3563,I427877,I427842,);
nor I_24973 (I427857,I428101,I428002);
nand I_24974 (I428154,I1095053,I1095050);
and I_24975 (I428171,I428154,I1095062);
DFFARX1 I_24976 (I428171,I3563,I427877,I428197,);
nor I_24977 (I427845,I428197,I428101);
not I_24978 (I428219,I428197);
nor I_24979 (I428236,I428219,I428010);
nor I_24980 (I428253,I427942,I428236);
DFFARX1 I_24981 (I428253,I3563,I427877,I427860,);
nor I_24982 (I428284,I428219,I428101);
nor I_24983 (I428301,I1095041,I1095050);
nor I_24984 (I427851,I428301,I428284);
not I_24985 (I428332,I428301);
nand I_24986 (I427854,I428061,I428332);
DFFARX1 I_24987 (I428301,I3563,I427877,I427866,);
DFFARX1 I_24988 (I428301,I3563,I427877,I427863,);
not I_24989 (I428421,I3570);
DFFARX1 I_24990 (I283912,I3563,I428421,I428447,);
DFFARX1 I_24991 (I428447,I3563,I428421,I428464,);
not I_24992 (I428413,I428464);
not I_24993 (I428486,I428447);
nand I_24994 (I428503,I283924,I283903);
and I_24995 (I428520,I428503,I283906);
DFFARX1 I_24996 (I428520,I3563,I428421,I428546,);
not I_24997 (I428554,I428546);
DFFARX1 I_24998 (I283915,I3563,I428421,I428580,);
and I_24999 (I428588,I428580,I283927);
nand I_25000 (I428605,I428580,I283927);
nand I_25001 (I428392,I428554,I428605);
DFFARX1 I_25002 (I283921,I3563,I428421,I428645,);
nor I_25003 (I428653,I428645,I428588);
DFFARX1 I_25004 (I428653,I3563,I428421,I428386,);
nor I_25005 (I428401,I428645,I428546);
nand I_25006 (I428698,I283909,I283906);
and I_25007 (I428715,I428698,I283918);
DFFARX1 I_25008 (I428715,I3563,I428421,I428741,);
nor I_25009 (I428389,I428741,I428645);
not I_25010 (I428763,I428741);
nor I_25011 (I428780,I428763,I428554);
nor I_25012 (I428797,I428486,I428780);
DFFARX1 I_25013 (I428797,I3563,I428421,I428404,);
nor I_25014 (I428828,I428763,I428645);
nor I_25015 (I428845,I283903,I283906);
nor I_25016 (I428395,I428845,I428828);
not I_25017 (I428876,I428845);
nand I_25018 (I428398,I428605,I428876);
DFFARX1 I_25019 (I428845,I3563,I428421,I428410,);
DFFARX1 I_25020 (I428845,I3563,I428421,I428407,);
not I_25021 (I428965,I3570);
DFFARX1 I_25022 (I3484,I3563,I428965,I428991,);
DFFARX1 I_25023 (I428991,I3563,I428965,I429008,);
not I_25024 (I428957,I429008);
not I_25025 (I429030,I428991);
nand I_25026 (I429047,I3180,I2372);
and I_25027 (I429064,I429047,I1516);
DFFARX1 I_25028 (I429064,I3563,I428965,I429090,);
not I_25029 (I429098,I429090);
DFFARX1 I_25030 (I3468,I3563,I428965,I429124,);
and I_25031 (I429132,I429124,I3548);
nand I_25032 (I429149,I429124,I3548);
nand I_25033 (I428936,I429098,I429149);
DFFARX1 I_25034 (I2684,I3563,I428965,I429189,);
nor I_25035 (I429197,I429189,I429132);
DFFARX1 I_25036 (I429197,I3563,I428965,I428930,);
nor I_25037 (I428945,I429189,I429090);
nand I_25038 (I429242,I2908,I2140);
and I_25039 (I429259,I429242,I3236);
DFFARX1 I_25040 (I429259,I3563,I428965,I429285,);
nor I_25041 (I428933,I429285,I429189);
not I_25042 (I429307,I429285);
nor I_25043 (I429324,I429307,I429098);
nor I_25044 (I429341,I429030,I429324);
DFFARX1 I_25045 (I429341,I3563,I428965,I428948,);
nor I_25046 (I429372,I429307,I429189);
nor I_25047 (I429389,I1868,I2140);
nor I_25048 (I428939,I429389,I429372);
not I_25049 (I429420,I429389);
nand I_25050 (I428942,I429149,I429420);
DFFARX1 I_25051 (I429389,I3563,I428965,I428954,);
DFFARX1 I_25052 (I429389,I3563,I428965,I428951,);
not I_25053 (I429509,I3570);
DFFARX1 I_25054 (I818973,I3563,I429509,I429535,);
DFFARX1 I_25055 (I429535,I3563,I429509,I429552,);
not I_25056 (I429501,I429552);
not I_25057 (I429574,I429535);
nand I_25058 (I429591,I818967,I818964);
and I_25059 (I429608,I429591,I818979);
DFFARX1 I_25060 (I429608,I3563,I429509,I429634,);
not I_25061 (I429642,I429634);
DFFARX1 I_25062 (I818967,I3563,I429509,I429668,);
and I_25063 (I429676,I429668,I818961);
nand I_25064 (I429693,I429668,I818961);
nand I_25065 (I429480,I429642,I429693);
DFFARX1 I_25066 (I818961,I3563,I429509,I429733,);
nor I_25067 (I429741,I429733,I429676);
DFFARX1 I_25068 (I429741,I3563,I429509,I429474,);
nor I_25069 (I429489,I429733,I429634);
nand I_25070 (I429786,I818976,I818970);
and I_25071 (I429803,I429786,I818964);
DFFARX1 I_25072 (I429803,I3563,I429509,I429829,);
nor I_25073 (I429477,I429829,I429733);
not I_25074 (I429851,I429829);
nor I_25075 (I429868,I429851,I429642);
nor I_25076 (I429885,I429574,I429868);
DFFARX1 I_25077 (I429885,I3563,I429509,I429492,);
nor I_25078 (I429916,I429851,I429733);
nor I_25079 (I429933,I818982,I818970);
nor I_25080 (I429483,I429933,I429916);
not I_25081 (I429964,I429933);
nand I_25082 (I429486,I429693,I429964);
DFFARX1 I_25083 (I429933,I3563,I429509,I429498,);
DFFARX1 I_25084 (I429933,I3563,I429509,I429495,);
not I_25085 (I430053,I3570);
DFFARX1 I_25086 (I220247,I3563,I430053,I430079,);
DFFARX1 I_25087 (I430079,I3563,I430053,I430096,);
not I_25088 (I430045,I430096);
not I_25089 (I430118,I430079);
nand I_25090 (I430135,I220259,I220238);
and I_25091 (I430152,I430135,I220241);
DFFARX1 I_25092 (I430152,I3563,I430053,I430178,);
not I_25093 (I430186,I430178);
DFFARX1 I_25094 (I220250,I3563,I430053,I430212,);
and I_25095 (I430220,I430212,I220262);
nand I_25096 (I430237,I430212,I220262);
nand I_25097 (I430024,I430186,I430237);
DFFARX1 I_25098 (I220256,I3563,I430053,I430277,);
nor I_25099 (I430285,I430277,I430220);
DFFARX1 I_25100 (I430285,I3563,I430053,I430018,);
nor I_25101 (I430033,I430277,I430178);
nand I_25102 (I430330,I220244,I220241);
and I_25103 (I430347,I430330,I220253);
DFFARX1 I_25104 (I430347,I3563,I430053,I430373,);
nor I_25105 (I430021,I430373,I430277);
not I_25106 (I430395,I430373);
nor I_25107 (I430412,I430395,I430186);
nor I_25108 (I430429,I430118,I430412);
DFFARX1 I_25109 (I430429,I3563,I430053,I430036,);
nor I_25110 (I430460,I430395,I430277);
nor I_25111 (I430477,I220238,I220241);
nor I_25112 (I430027,I430477,I430460);
not I_25113 (I430508,I430477);
nand I_25114 (I430030,I430237,I430508);
DFFARX1 I_25115 (I430477,I3563,I430053,I430042,);
DFFARX1 I_25116 (I430477,I3563,I430053,I430039,);
not I_25117 (I430597,I3570);
DFFARX1 I_25118 (I1087051,I3563,I430597,I430623,);
DFFARX1 I_25119 (I430623,I3563,I430597,I430640,);
not I_25120 (I430589,I430640);
not I_25121 (I430662,I430623);
nand I_25122 (I430679,I1087051,I1087069);
and I_25123 (I430696,I430679,I1087063);
DFFARX1 I_25124 (I430696,I3563,I430597,I430722,);
not I_25125 (I430730,I430722);
DFFARX1 I_25126 (I1087057,I3563,I430597,I430756,);
and I_25127 (I430764,I430756,I1087066);
nand I_25128 (I430781,I430756,I1087066);
nand I_25129 (I430568,I430730,I430781);
DFFARX1 I_25130 (I1087054,I3563,I430597,I430821,);
nor I_25131 (I430829,I430821,I430764);
DFFARX1 I_25132 (I430829,I3563,I430597,I430562,);
nor I_25133 (I430577,I430821,I430722);
nand I_25134 (I430874,I1087054,I1087072);
and I_25135 (I430891,I430874,I1087057);
DFFARX1 I_25136 (I430891,I3563,I430597,I430917,);
nor I_25137 (I430565,I430917,I430821);
not I_25138 (I430939,I430917);
nor I_25139 (I430956,I430939,I430730);
nor I_25140 (I430973,I430662,I430956);
DFFARX1 I_25141 (I430973,I3563,I430597,I430580,);
nor I_25142 (I431004,I430939,I430821);
nor I_25143 (I431021,I1087060,I1087072);
nor I_25144 (I430571,I431021,I431004);
not I_25145 (I431052,I431021);
nand I_25146 (I430574,I430781,I431052);
DFFARX1 I_25147 (I431021,I3563,I430597,I430586,);
DFFARX1 I_25148 (I431021,I3563,I430597,I430583,);
not I_25149 (I431141,I3570);
DFFARX1 I_25150 (I66666,I3563,I431141,I431167,);
DFFARX1 I_25151 (I431167,I3563,I431141,I431184,);
not I_25152 (I431133,I431184);
not I_25153 (I431206,I431167);
nand I_25154 (I431223,I66681,I66660);
and I_25155 (I431240,I431223,I66663);
DFFARX1 I_25156 (I431240,I3563,I431141,I431266,);
not I_25157 (I431274,I431266);
DFFARX1 I_25158 (I66669,I3563,I431141,I431300,);
and I_25159 (I431308,I431300,I66663);
nand I_25160 (I431325,I431300,I66663);
nand I_25161 (I431112,I431274,I431325);
DFFARX1 I_25162 (I66678,I3563,I431141,I431365,);
nor I_25163 (I431373,I431365,I431308);
DFFARX1 I_25164 (I431373,I3563,I431141,I431106,);
nor I_25165 (I431121,I431365,I431266);
nand I_25166 (I431418,I66660,I66675);
and I_25167 (I431435,I431418,I66672);
DFFARX1 I_25168 (I431435,I3563,I431141,I431461,);
nor I_25169 (I431109,I431461,I431365);
not I_25170 (I431483,I431461);
nor I_25171 (I431500,I431483,I431274);
nor I_25172 (I431517,I431206,I431500);
DFFARX1 I_25173 (I431517,I3563,I431141,I431124,);
nor I_25174 (I431548,I431483,I431365);
nor I_25175 (I431565,I66684,I66675);
nor I_25176 (I431115,I431565,I431548);
not I_25177 (I431596,I431565);
nand I_25178 (I431118,I431325,I431596);
DFFARX1 I_25179 (I431565,I3563,I431141,I431130,);
DFFARX1 I_25180 (I431565,I3563,I431141,I431127,);
not I_25181 (I431685,I3570);
DFFARX1 I_25182 (I165507,I3563,I431685,I431711,);
DFFARX1 I_25183 (I431711,I3563,I431685,I431728,);
not I_25184 (I431677,I431728);
not I_25185 (I431750,I431711);
nand I_25186 (I431767,I165519,I165498);
and I_25187 (I431784,I431767,I165501);
DFFARX1 I_25188 (I431784,I3563,I431685,I431810,);
not I_25189 (I431818,I431810);
DFFARX1 I_25190 (I165510,I3563,I431685,I431844,);
and I_25191 (I431852,I431844,I165522);
nand I_25192 (I431869,I431844,I165522);
nand I_25193 (I431656,I431818,I431869);
DFFARX1 I_25194 (I165516,I3563,I431685,I431909,);
nor I_25195 (I431917,I431909,I431852);
DFFARX1 I_25196 (I431917,I3563,I431685,I431650,);
nor I_25197 (I431665,I431909,I431810);
nand I_25198 (I431962,I165504,I165501);
and I_25199 (I431979,I431962,I165513);
DFFARX1 I_25200 (I431979,I3563,I431685,I432005,);
nor I_25201 (I431653,I432005,I431909);
not I_25202 (I432027,I432005);
nor I_25203 (I432044,I432027,I431818);
nor I_25204 (I432061,I431750,I432044);
DFFARX1 I_25205 (I432061,I3563,I431685,I431668,);
nor I_25206 (I432092,I432027,I431909);
nor I_25207 (I432109,I165498,I165501);
nor I_25208 (I431659,I432109,I432092);
not I_25209 (I432140,I432109);
nand I_25210 (I431662,I431869,I432140);
DFFARX1 I_25211 (I432109,I3563,I431685,I431674,);
DFFARX1 I_25212 (I432109,I3563,I431685,I431671,);
not I_25213 (I432229,I3570);
DFFARX1 I_25214 (I1059001,I3563,I432229,I432255,);
DFFARX1 I_25215 (I432255,I3563,I432229,I432272,);
not I_25216 (I432221,I432272);
not I_25217 (I432294,I432255);
nand I_25218 (I432311,I1059001,I1059019);
and I_25219 (I432328,I432311,I1059013);
DFFARX1 I_25220 (I432328,I3563,I432229,I432354,);
not I_25221 (I432362,I432354);
DFFARX1 I_25222 (I1059007,I3563,I432229,I432388,);
and I_25223 (I432396,I432388,I1059016);
nand I_25224 (I432413,I432388,I1059016);
nand I_25225 (I432200,I432362,I432413);
DFFARX1 I_25226 (I1059004,I3563,I432229,I432453,);
nor I_25227 (I432461,I432453,I432396);
DFFARX1 I_25228 (I432461,I3563,I432229,I432194,);
nor I_25229 (I432209,I432453,I432354);
nand I_25230 (I432506,I1059004,I1059022);
and I_25231 (I432523,I432506,I1059007);
DFFARX1 I_25232 (I432523,I3563,I432229,I432549,);
nor I_25233 (I432197,I432549,I432453);
not I_25234 (I432571,I432549);
nor I_25235 (I432588,I432571,I432362);
nor I_25236 (I432605,I432294,I432588);
DFFARX1 I_25237 (I432605,I3563,I432229,I432212,);
nor I_25238 (I432636,I432571,I432453);
nor I_25239 (I432653,I1059010,I1059022);
nor I_25240 (I432203,I432653,I432636);
not I_25241 (I432684,I432653);
nand I_25242 (I432206,I432413,I432684);
DFFARX1 I_25243 (I432653,I3563,I432229,I432218,);
DFFARX1 I_25244 (I432653,I3563,I432229,I432215,);
not I_25245 (I432773,I3570);
DFFARX1 I_25246 (I358112,I3563,I432773,I432799,);
DFFARX1 I_25247 (I432799,I3563,I432773,I432816,);
not I_25248 (I432765,I432816);
not I_25249 (I432838,I432799);
nand I_25250 (I432855,I358091,I358115);
and I_25251 (I432872,I432855,I358118);
DFFARX1 I_25252 (I432872,I3563,I432773,I432898,);
not I_25253 (I432906,I432898);
DFFARX1 I_25254 (I358100,I3563,I432773,I432932,);
and I_25255 (I432940,I432932,I358106);
nand I_25256 (I432957,I432932,I358106);
nand I_25257 (I432744,I432906,I432957);
DFFARX1 I_25258 (I358094,I3563,I432773,I432997,);
nor I_25259 (I433005,I432997,I432940);
DFFARX1 I_25260 (I433005,I3563,I432773,I432738,);
nor I_25261 (I432753,I432997,I432898);
nand I_25262 (I433050,I358103,I358091);
and I_25263 (I433067,I433050,I358097);
DFFARX1 I_25264 (I433067,I3563,I432773,I433093,);
nor I_25265 (I432741,I433093,I432997);
not I_25266 (I433115,I433093);
nor I_25267 (I433132,I433115,I432906);
nor I_25268 (I433149,I432838,I433132);
DFFARX1 I_25269 (I433149,I3563,I432773,I432756,);
nor I_25270 (I433180,I433115,I432997);
nor I_25271 (I433197,I358109,I358091);
nor I_25272 (I432747,I433197,I433180);
not I_25273 (I433228,I433197);
nand I_25274 (I432750,I432957,I433228);
DFFARX1 I_25275 (I433197,I3563,I432773,I432762,);
DFFARX1 I_25276 (I433197,I3563,I432773,I432759,);
not I_25277 (I433317,I3570);
DFFARX1 I_25278 (I756098,I3563,I433317,I433343,);
DFFARX1 I_25279 (I433343,I3563,I433317,I433360,);
not I_25280 (I433309,I433360);
not I_25281 (I433382,I433343);
nand I_25282 (I433399,I756119,I756110);
and I_25283 (I433416,I433399,I756098);
DFFARX1 I_25284 (I433416,I3563,I433317,I433442,);
not I_25285 (I433450,I433442);
DFFARX1 I_25286 (I756104,I3563,I433317,I433476,);
and I_25287 (I433484,I433476,I756101);
nand I_25288 (I433501,I433476,I756101);
nand I_25289 (I433288,I433450,I433501);
DFFARX1 I_25290 (I756095,I3563,I433317,I433541,);
nor I_25291 (I433549,I433541,I433484);
DFFARX1 I_25292 (I433549,I3563,I433317,I433282,);
nor I_25293 (I433297,I433541,I433442);
nand I_25294 (I433594,I756095,I756107);
and I_25295 (I433611,I433594,I756116);
DFFARX1 I_25296 (I433611,I3563,I433317,I433637,);
nor I_25297 (I433285,I433637,I433541);
not I_25298 (I433659,I433637);
nor I_25299 (I433676,I433659,I433450);
nor I_25300 (I433693,I433382,I433676);
DFFARX1 I_25301 (I433693,I3563,I433317,I433300,);
nor I_25302 (I433724,I433659,I433541);
nor I_25303 (I433741,I756113,I756107);
nor I_25304 (I433291,I433741,I433724);
not I_25305 (I433772,I433741);
nand I_25306 (I433294,I433501,I433772);
DFFARX1 I_25307 (I433741,I3563,I433317,I433306,);
DFFARX1 I_25308 (I433741,I3563,I433317,I433303,);
not I_25309 (I433861,I3570);
DFFARX1 I_25310 (I1194460,I3563,I433861,I433887,);
DFFARX1 I_25311 (I433887,I3563,I433861,I433904,);
not I_25312 (I433853,I433904);
not I_25313 (I433926,I433887);
nand I_25314 (I433943,I1194472,I1194460);
and I_25315 (I433960,I433943,I1194463);
DFFARX1 I_25316 (I433960,I3563,I433861,I433986,);
not I_25317 (I433994,I433986);
DFFARX1 I_25318 (I1194481,I3563,I433861,I434020,);
and I_25319 (I434028,I434020,I1194457);
nand I_25320 (I434045,I434020,I1194457);
nand I_25321 (I433832,I433994,I434045);
DFFARX1 I_25322 (I1194475,I3563,I433861,I434085,);
nor I_25323 (I434093,I434085,I434028);
DFFARX1 I_25324 (I434093,I3563,I433861,I433826,);
nor I_25325 (I433841,I434085,I433986);
nand I_25326 (I434138,I1194469,I1194466);
and I_25327 (I434155,I434138,I1194478);
DFFARX1 I_25328 (I434155,I3563,I433861,I434181,);
nor I_25329 (I433829,I434181,I434085);
not I_25330 (I434203,I434181);
nor I_25331 (I434220,I434203,I433994);
nor I_25332 (I434237,I433926,I434220);
DFFARX1 I_25333 (I434237,I3563,I433861,I433844,);
nor I_25334 (I434268,I434203,I434085);
nor I_25335 (I434285,I1194457,I1194466);
nor I_25336 (I433835,I434285,I434268);
not I_25337 (I434316,I434285);
nand I_25338 (I433838,I434045,I434316);
DFFARX1 I_25339 (I434285,I3563,I433861,I433850,);
DFFARX1 I_25340 (I434285,I3563,I433861,I433847,);
not I_25341 (I434405,I3570);
DFFARX1 I_25342 (I1069660,I3563,I434405,I434431,);
DFFARX1 I_25343 (I434431,I3563,I434405,I434448,);
not I_25344 (I434397,I434448);
not I_25345 (I434470,I434431);
nand I_25346 (I434487,I1069660,I1069678);
and I_25347 (I434504,I434487,I1069672);
DFFARX1 I_25348 (I434504,I3563,I434405,I434530,);
not I_25349 (I434538,I434530);
DFFARX1 I_25350 (I1069666,I3563,I434405,I434564,);
and I_25351 (I434572,I434564,I1069675);
nand I_25352 (I434589,I434564,I1069675);
nand I_25353 (I434376,I434538,I434589);
DFFARX1 I_25354 (I1069663,I3563,I434405,I434629,);
nor I_25355 (I434637,I434629,I434572);
DFFARX1 I_25356 (I434637,I3563,I434405,I434370,);
nor I_25357 (I434385,I434629,I434530);
nand I_25358 (I434682,I1069663,I1069681);
and I_25359 (I434699,I434682,I1069666);
DFFARX1 I_25360 (I434699,I3563,I434405,I434725,);
nor I_25361 (I434373,I434725,I434629);
not I_25362 (I434747,I434725);
nor I_25363 (I434764,I434747,I434538);
nor I_25364 (I434781,I434470,I434764);
DFFARX1 I_25365 (I434781,I3563,I434405,I434388,);
nor I_25366 (I434812,I434747,I434629);
nor I_25367 (I434829,I1069669,I1069681);
nor I_25368 (I434379,I434829,I434812);
not I_25369 (I434860,I434829);
nand I_25370 (I434382,I434589,I434860);
DFFARX1 I_25371 (I434829,I3563,I434405,I434394,);
DFFARX1 I_25372 (I434829,I3563,I434405,I434391,);
not I_25373 (I434949,I3570);
DFFARX1 I_25374 (I776328,I3563,I434949,I434975,);
DFFARX1 I_25375 (I434975,I3563,I434949,I434992,);
not I_25376 (I434941,I434992);
not I_25377 (I435014,I434975);
nand I_25378 (I435031,I776349,I776340);
and I_25379 (I435048,I435031,I776328);
DFFARX1 I_25380 (I435048,I3563,I434949,I435074,);
not I_25381 (I435082,I435074);
DFFARX1 I_25382 (I776334,I3563,I434949,I435108,);
and I_25383 (I435116,I435108,I776331);
nand I_25384 (I435133,I435108,I776331);
nand I_25385 (I434920,I435082,I435133);
DFFARX1 I_25386 (I776325,I3563,I434949,I435173,);
nor I_25387 (I435181,I435173,I435116);
DFFARX1 I_25388 (I435181,I3563,I434949,I434914,);
nor I_25389 (I434929,I435173,I435074);
nand I_25390 (I435226,I776325,I776337);
and I_25391 (I435243,I435226,I776346);
DFFARX1 I_25392 (I435243,I3563,I434949,I435269,);
nor I_25393 (I434917,I435269,I435173);
not I_25394 (I435291,I435269);
nor I_25395 (I435308,I435291,I435082);
nor I_25396 (I435325,I435014,I435308);
DFFARX1 I_25397 (I435325,I3563,I434949,I434932,);
nor I_25398 (I435356,I435291,I435173);
nor I_25399 (I435373,I776343,I776337);
nor I_25400 (I434923,I435373,I435356);
not I_25401 (I435404,I435373);
nand I_25402 (I434926,I435133,I435404);
DFFARX1 I_25403 (I435373,I3563,I434949,I434938,);
DFFARX1 I_25404 (I435373,I3563,I434949,I434935,);
not I_25405 (I435493,I3570);
DFFARX1 I_25406 (I244047,I3563,I435493,I435519,);
DFFARX1 I_25407 (I435519,I3563,I435493,I435536,);
not I_25408 (I435485,I435536);
not I_25409 (I435558,I435519);
nand I_25410 (I435575,I244059,I244038);
and I_25411 (I435592,I435575,I244041);
DFFARX1 I_25412 (I435592,I3563,I435493,I435618,);
not I_25413 (I435626,I435618);
DFFARX1 I_25414 (I244050,I3563,I435493,I435652,);
and I_25415 (I435660,I435652,I244062);
nand I_25416 (I435677,I435652,I244062);
nand I_25417 (I435464,I435626,I435677);
DFFARX1 I_25418 (I244056,I3563,I435493,I435717,);
nor I_25419 (I435725,I435717,I435660);
DFFARX1 I_25420 (I435725,I3563,I435493,I435458,);
nor I_25421 (I435473,I435717,I435618);
nand I_25422 (I435770,I244044,I244041);
and I_25423 (I435787,I435770,I244053);
DFFARX1 I_25424 (I435787,I3563,I435493,I435813,);
nor I_25425 (I435461,I435813,I435717);
not I_25426 (I435835,I435813);
nor I_25427 (I435852,I435835,I435626);
nor I_25428 (I435869,I435558,I435852);
DFFARX1 I_25429 (I435869,I3563,I435493,I435476,);
nor I_25430 (I435900,I435835,I435717);
nor I_25431 (I435917,I244038,I244041);
nor I_25432 (I435467,I435917,I435900);
not I_25433 (I435948,I435917);
nand I_25434 (I435470,I435677,I435948);
DFFARX1 I_25435 (I435917,I3563,I435493,I435482,);
DFFARX1 I_25436 (I435917,I3563,I435493,I435479,);
not I_25437 (I436037,I3570);
DFFARX1 I_25438 (I183952,I3563,I436037,I436063,);
DFFARX1 I_25439 (I436063,I3563,I436037,I436080,);
not I_25440 (I436029,I436080);
not I_25441 (I436102,I436063);
nand I_25442 (I436119,I183964,I183943);
and I_25443 (I436136,I436119,I183946);
DFFARX1 I_25444 (I436136,I3563,I436037,I436162,);
not I_25445 (I436170,I436162);
DFFARX1 I_25446 (I183955,I3563,I436037,I436196,);
and I_25447 (I436204,I436196,I183967);
nand I_25448 (I436221,I436196,I183967);
nand I_25449 (I436008,I436170,I436221);
DFFARX1 I_25450 (I183961,I3563,I436037,I436261,);
nor I_25451 (I436269,I436261,I436204);
DFFARX1 I_25452 (I436269,I3563,I436037,I436002,);
nor I_25453 (I436017,I436261,I436162);
nand I_25454 (I436314,I183949,I183946);
and I_25455 (I436331,I436314,I183958);
DFFARX1 I_25456 (I436331,I3563,I436037,I436357,);
nor I_25457 (I436005,I436357,I436261);
not I_25458 (I436379,I436357);
nor I_25459 (I436396,I436379,I436170);
nor I_25460 (I436413,I436102,I436396);
DFFARX1 I_25461 (I436413,I3563,I436037,I436020,);
nor I_25462 (I436444,I436379,I436261);
nor I_25463 (I436461,I183943,I183946);
nor I_25464 (I436011,I436461,I436444);
not I_25465 (I436492,I436461);
nand I_25466 (I436014,I436221,I436492);
DFFARX1 I_25467 (I436461,I3563,I436037,I436026,);
DFFARX1 I_25468 (I436461,I3563,I436037,I436023,);
not I_25469 (I436581,I3570);
DFFARX1 I_25470 (I1267628,I3563,I436581,I436607,);
DFFARX1 I_25471 (I436607,I3563,I436581,I436624,);
not I_25472 (I436573,I436624);
not I_25473 (I436646,I436607);
nand I_25474 (I436663,I1267640,I1267643);
and I_25475 (I436680,I436663,I1267646);
DFFARX1 I_25476 (I436680,I3563,I436581,I436706,);
not I_25477 (I436714,I436706);
DFFARX1 I_25478 (I1267631,I3563,I436581,I436740,);
and I_25479 (I436748,I436740,I1267637);
nand I_25480 (I436765,I436740,I1267637);
nand I_25481 (I436552,I436714,I436765);
DFFARX1 I_25482 (I1267625,I3563,I436581,I436805,);
nor I_25483 (I436813,I436805,I436748);
DFFARX1 I_25484 (I436813,I3563,I436581,I436546,);
nor I_25485 (I436561,I436805,I436706);
nand I_25486 (I436858,I1267628,I1267649);
and I_25487 (I436875,I436858,I1267634);
DFFARX1 I_25488 (I436875,I3563,I436581,I436901,);
nor I_25489 (I436549,I436901,I436805);
not I_25490 (I436923,I436901);
nor I_25491 (I436940,I436923,I436714);
nor I_25492 (I436957,I436646,I436940);
DFFARX1 I_25493 (I436957,I3563,I436581,I436564,);
nor I_25494 (I436988,I436923,I436805);
nor I_25495 (I437005,I1267625,I1267649);
nor I_25496 (I436555,I437005,I436988);
not I_25497 (I437036,I437005);
nand I_25498 (I436558,I436765,I437036);
DFFARX1 I_25499 (I437005,I3563,I436581,I436570,);
DFFARX1 I_25500 (I437005,I3563,I436581,I436567,);
not I_25501 (I437125,I3570);
DFFARX1 I_25502 (I93543,I3563,I437125,I437151,);
DFFARX1 I_25503 (I437151,I3563,I437125,I437168,);
not I_25504 (I437117,I437168);
not I_25505 (I437190,I437151);
nand I_25506 (I437207,I93558,I93537);
and I_25507 (I437224,I437207,I93540);
DFFARX1 I_25508 (I437224,I3563,I437125,I437250,);
not I_25509 (I437258,I437250);
DFFARX1 I_25510 (I93546,I3563,I437125,I437284,);
and I_25511 (I437292,I437284,I93540);
nand I_25512 (I437309,I437284,I93540);
nand I_25513 (I437096,I437258,I437309);
DFFARX1 I_25514 (I93555,I3563,I437125,I437349,);
nor I_25515 (I437357,I437349,I437292);
DFFARX1 I_25516 (I437357,I3563,I437125,I437090,);
nor I_25517 (I437105,I437349,I437250);
nand I_25518 (I437402,I93537,I93552);
and I_25519 (I437419,I437402,I93549);
DFFARX1 I_25520 (I437419,I3563,I437125,I437445,);
nor I_25521 (I437093,I437445,I437349);
not I_25522 (I437467,I437445);
nor I_25523 (I437484,I437467,I437258);
nor I_25524 (I437501,I437190,I437484);
DFFARX1 I_25525 (I437501,I3563,I437125,I437108,);
nor I_25526 (I437532,I437467,I437349);
nor I_25527 (I437549,I93561,I93552);
nor I_25528 (I437099,I437549,I437532);
not I_25529 (I437580,I437549);
nand I_25530 (I437102,I437309,I437580);
DFFARX1 I_25531 (I437549,I3563,I437125,I437114,);
DFFARX1 I_25532 (I437549,I3563,I437125,I437111,);
not I_25533 (I437669,I3570);
DFFARX1 I_25534 (I969791,I3563,I437669,I437695,);
DFFARX1 I_25535 (I437695,I3563,I437669,I437712,);
not I_25536 (I437661,I437712);
not I_25537 (I437734,I437695);
nand I_25538 (I437751,I969806,I969794);
and I_25539 (I437768,I437751,I969785);
DFFARX1 I_25540 (I437768,I3563,I437669,I437794,);
not I_25541 (I437802,I437794);
DFFARX1 I_25542 (I969797,I3563,I437669,I437828,);
and I_25543 (I437836,I437828,I969788);
nand I_25544 (I437853,I437828,I969788);
nand I_25545 (I437640,I437802,I437853);
DFFARX1 I_25546 (I969803,I3563,I437669,I437893,);
nor I_25547 (I437901,I437893,I437836);
DFFARX1 I_25548 (I437901,I3563,I437669,I437634,);
nor I_25549 (I437649,I437893,I437794);
nand I_25550 (I437946,I969812,I969800);
and I_25551 (I437963,I437946,I969809);
DFFARX1 I_25552 (I437963,I3563,I437669,I437989,);
nor I_25553 (I437637,I437989,I437893);
not I_25554 (I438011,I437989);
nor I_25555 (I438028,I438011,I437802);
nor I_25556 (I438045,I437734,I438028);
DFFARX1 I_25557 (I438045,I3563,I437669,I437652,);
nor I_25558 (I438076,I438011,I437893);
nor I_25559 (I438093,I969785,I969800);
nor I_25560 (I437643,I438093,I438076);
not I_25561 (I438124,I438093);
nand I_25562 (I437646,I437853,I438124);
DFFARX1 I_25563 (I438093,I3563,I437669,I437658,);
DFFARX1 I_25564 (I438093,I3563,I437669,I437655,);
not I_25565 (I438213,I3570);
DFFARX1 I_25566 (I1175964,I3563,I438213,I438239,);
DFFARX1 I_25567 (I438239,I3563,I438213,I438256,);
not I_25568 (I438205,I438256);
not I_25569 (I438278,I438239);
nand I_25570 (I438295,I1175976,I1175964);
and I_25571 (I438312,I438295,I1175967);
DFFARX1 I_25572 (I438312,I3563,I438213,I438338,);
not I_25573 (I438346,I438338);
DFFARX1 I_25574 (I1175985,I3563,I438213,I438372,);
and I_25575 (I438380,I438372,I1175961);
nand I_25576 (I438397,I438372,I1175961);
nand I_25577 (I438184,I438346,I438397);
DFFARX1 I_25578 (I1175979,I3563,I438213,I438437,);
nor I_25579 (I438445,I438437,I438380);
DFFARX1 I_25580 (I438445,I3563,I438213,I438178,);
nor I_25581 (I438193,I438437,I438338);
nand I_25582 (I438490,I1175973,I1175970);
and I_25583 (I438507,I438490,I1175982);
DFFARX1 I_25584 (I438507,I3563,I438213,I438533,);
nor I_25585 (I438181,I438533,I438437);
not I_25586 (I438555,I438533);
nor I_25587 (I438572,I438555,I438346);
nor I_25588 (I438589,I438278,I438572);
DFFARX1 I_25589 (I438589,I3563,I438213,I438196,);
nor I_25590 (I438620,I438555,I438437);
nor I_25591 (I438637,I1175961,I1175970);
nor I_25592 (I438187,I438637,I438620);
not I_25593 (I438668,I438637);
nand I_25594 (I438190,I438397,I438668);
DFFARX1 I_25595 (I438637,I3563,I438213,I438202,);
DFFARX1 I_25596 (I438637,I3563,I438213,I438199,);
not I_25597 (I438757,I3570);
DFFARX1 I_25598 (I564984,I3563,I438757,I438783,);
DFFARX1 I_25599 (I438783,I3563,I438757,I438800,);
not I_25600 (I438749,I438800);
not I_25601 (I438822,I438783);
nand I_25602 (I438839,I564987,I565005);
and I_25603 (I438856,I438839,I564993);
DFFARX1 I_25604 (I438856,I3563,I438757,I438882,);
not I_25605 (I438890,I438882);
DFFARX1 I_25606 (I564984,I3563,I438757,I438916,);
and I_25607 (I438924,I438916,I565002);
nand I_25608 (I438941,I438916,I565002);
nand I_25609 (I438728,I438890,I438941);
DFFARX1 I_25610 (I564996,I3563,I438757,I438981,);
nor I_25611 (I438989,I438981,I438924);
DFFARX1 I_25612 (I438989,I3563,I438757,I438722,);
nor I_25613 (I438737,I438981,I438882);
nand I_25614 (I439034,I564999,I564981);
and I_25615 (I439051,I439034,I564990);
DFFARX1 I_25616 (I439051,I3563,I438757,I439077,);
nor I_25617 (I438725,I439077,I438981);
not I_25618 (I439099,I439077);
nor I_25619 (I439116,I439099,I438890);
nor I_25620 (I439133,I438822,I439116);
DFFARX1 I_25621 (I439133,I3563,I438757,I438740,);
nor I_25622 (I439164,I439099,I438981);
nor I_25623 (I439181,I564981,I564981);
nor I_25624 (I438731,I439181,I439164);
not I_25625 (I439212,I439181);
nand I_25626 (I438734,I438941,I439212);
DFFARX1 I_25627 (I439181,I3563,I438757,I438746,);
DFFARX1 I_25628 (I439181,I3563,I438757,I438743,);
not I_25629 (I439301,I3570);
DFFARX1 I_25630 (I30309,I3563,I439301,I439327,);
DFFARX1 I_25631 (I439327,I3563,I439301,I439344,);
not I_25632 (I439293,I439344);
not I_25633 (I439366,I439327);
nand I_25634 (I439383,I30297,I30312);
and I_25635 (I439400,I439383,I30300);
DFFARX1 I_25636 (I439400,I3563,I439301,I439426,);
not I_25637 (I439434,I439426);
DFFARX1 I_25638 (I30321,I3563,I439301,I439460,);
and I_25639 (I439468,I439460,I30315);
nand I_25640 (I439485,I439460,I30315);
nand I_25641 (I439272,I439434,I439485);
DFFARX1 I_25642 (I30318,I3563,I439301,I439525,);
nor I_25643 (I439533,I439525,I439468);
DFFARX1 I_25644 (I439533,I3563,I439301,I439266,);
nor I_25645 (I439281,I439525,I439426);
nand I_25646 (I439578,I30297,I30300);
and I_25647 (I439595,I439578,I30303);
DFFARX1 I_25648 (I439595,I3563,I439301,I439621,);
nor I_25649 (I439269,I439621,I439525);
not I_25650 (I439643,I439621);
nor I_25651 (I439660,I439643,I439434);
nor I_25652 (I439677,I439366,I439660);
DFFARX1 I_25653 (I439677,I3563,I439301,I439284,);
nor I_25654 (I439708,I439643,I439525);
nor I_25655 (I439725,I30306,I30300);
nor I_25656 (I439275,I439725,I439708);
not I_25657 (I439756,I439725);
nand I_25658 (I439278,I439485,I439756);
DFFARX1 I_25659 (I439725,I3563,I439301,I439290,);
DFFARX1 I_25660 (I439725,I3563,I439301,I439287,);
not I_25661 (I439845,I3570);
DFFARX1 I_25662 (I241072,I3563,I439845,I439871,);
DFFARX1 I_25663 (I439871,I3563,I439845,I439888,);
not I_25664 (I439837,I439888);
not I_25665 (I439910,I439871);
nand I_25666 (I439927,I241084,I241063);
and I_25667 (I439944,I439927,I241066);
DFFARX1 I_25668 (I439944,I3563,I439845,I439970,);
not I_25669 (I439978,I439970);
DFFARX1 I_25670 (I241075,I3563,I439845,I440004,);
and I_25671 (I440012,I440004,I241087);
nand I_25672 (I440029,I440004,I241087);
nand I_25673 (I439816,I439978,I440029);
DFFARX1 I_25674 (I241081,I3563,I439845,I440069,);
nor I_25675 (I440077,I440069,I440012);
DFFARX1 I_25676 (I440077,I3563,I439845,I439810,);
nor I_25677 (I439825,I440069,I439970);
nand I_25678 (I440122,I241069,I241066);
and I_25679 (I440139,I440122,I241078);
DFFARX1 I_25680 (I440139,I3563,I439845,I440165,);
nor I_25681 (I439813,I440165,I440069);
not I_25682 (I440187,I440165);
nor I_25683 (I440204,I440187,I439978);
nor I_25684 (I440221,I439910,I440204);
DFFARX1 I_25685 (I440221,I3563,I439845,I439828,);
nor I_25686 (I440252,I440187,I440069);
nor I_25687 (I440269,I241063,I241066);
nor I_25688 (I439819,I440269,I440252);
not I_25689 (I440300,I440269);
nand I_25690 (I439822,I440029,I440300);
DFFARX1 I_25691 (I440269,I3563,I439845,I439834,);
DFFARX1 I_25692 (I440269,I3563,I439845,I439831,);
not I_25693 (I440389,I3570);
DFFARX1 I_25694 (I183357,I3563,I440389,I440415,);
DFFARX1 I_25695 (I440415,I3563,I440389,I440432,);
not I_25696 (I440381,I440432);
not I_25697 (I440454,I440415);
nand I_25698 (I440471,I183369,I183348);
and I_25699 (I440488,I440471,I183351);
DFFARX1 I_25700 (I440488,I3563,I440389,I440514,);
not I_25701 (I440522,I440514);
DFFARX1 I_25702 (I183360,I3563,I440389,I440548,);
and I_25703 (I440556,I440548,I183372);
nand I_25704 (I440573,I440548,I183372);
nand I_25705 (I440360,I440522,I440573);
DFFARX1 I_25706 (I183366,I3563,I440389,I440613,);
nor I_25707 (I440621,I440613,I440556);
DFFARX1 I_25708 (I440621,I3563,I440389,I440354,);
nor I_25709 (I440369,I440613,I440514);
nand I_25710 (I440666,I183354,I183351);
and I_25711 (I440683,I440666,I183363);
DFFARX1 I_25712 (I440683,I3563,I440389,I440709,);
nor I_25713 (I440357,I440709,I440613);
not I_25714 (I440731,I440709);
nor I_25715 (I440748,I440731,I440522);
nor I_25716 (I440765,I440454,I440748);
DFFARX1 I_25717 (I440765,I3563,I440389,I440372,);
nor I_25718 (I440796,I440731,I440613);
nor I_25719 (I440813,I183348,I183351);
nor I_25720 (I440363,I440813,I440796);
not I_25721 (I440844,I440813);
nand I_25722 (I440366,I440573,I440844);
DFFARX1 I_25723 (I440813,I3563,I440389,I440378,);
DFFARX1 I_25724 (I440813,I3563,I440389,I440375,);
not I_25725 (I440933,I3570);
DFFARX1 I_25726 (I279152,I3563,I440933,I440959,);
DFFARX1 I_25727 (I440959,I3563,I440933,I440976,);
not I_25728 (I440925,I440976);
not I_25729 (I440998,I440959);
nand I_25730 (I441015,I279164,I279143);
and I_25731 (I441032,I441015,I279146);
DFFARX1 I_25732 (I441032,I3563,I440933,I441058,);
not I_25733 (I441066,I441058);
DFFARX1 I_25734 (I279155,I3563,I440933,I441092,);
and I_25735 (I441100,I441092,I279167);
nand I_25736 (I441117,I441092,I279167);
nand I_25737 (I440904,I441066,I441117);
DFFARX1 I_25738 (I279161,I3563,I440933,I441157,);
nor I_25739 (I441165,I441157,I441100);
DFFARX1 I_25740 (I441165,I3563,I440933,I440898,);
nor I_25741 (I440913,I441157,I441058);
nand I_25742 (I441210,I279149,I279146);
and I_25743 (I441227,I441210,I279158);
DFFARX1 I_25744 (I441227,I3563,I440933,I441253,);
nor I_25745 (I440901,I441253,I441157);
not I_25746 (I441275,I441253);
nor I_25747 (I441292,I441275,I441066);
nor I_25748 (I441309,I440998,I441292);
DFFARX1 I_25749 (I441309,I3563,I440933,I440916,);
nor I_25750 (I441340,I441275,I441157);
nor I_25751 (I441357,I279143,I279146);
nor I_25752 (I440907,I441357,I441340);
not I_25753 (I441388,I441357);
nand I_25754 (I440910,I441117,I441388);
DFFARX1 I_25755 (I441357,I3563,I440933,I440922,);
DFFARX1 I_25756 (I441357,I3563,I440933,I440919,);
not I_25757 (I441477,I3570);
DFFARX1 I_25758 (I1198506,I3563,I441477,I441503,);
DFFARX1 I_25759 (I441503,I3563,I441477,I441520,);
not I_25760 (I441469,I441520);
not I_25761 (I441542,I441503);
nand I_25762 (I441559,I1198518,I1198506);
and I_25763 (I441576,I441559,I1198509);
DFFARX1 I_25764 (I441576,I3563,I441477,I441602,);
not I_25765 (I441610,I441602);
DFFARX1 I_25766 (I1198527,I3563,I441477,I441636,);
and I_25767 (I441644,I441636,I1198503);
nand I_25768 (I441661,I441636,I1198503);
nand I_25769 (I441448,I441610,I441661);
DFFARX1 I_25770 (I1198521,I3563,I441477,I441701,);
nor I_25771 (I441709,I441701,I441644);
DFFARX1 I_25772 (I441709,I3563,I441477,I441442,);
nor I_25773 (I441457,I441701,I441602);
nand I_25774 (I441754,I1198515,I1198512);
and I_25775 (I441771,I441754,I1198524);
DFFARX1 I_25776 (I441771,I3563,I441477,I441797,);
nor I_25777 (I441445,I441797,I441701);
not I_25778 (I441819,I441797);
nor I_25779 (I441836,I441819,I441610);
nor I_25780 (I441853,I441542,I441836);
DFFARX1 I_25781 (I441853,I3563,I441477,I441460,);
nor I_25782 (I441884,I441819,I441701);
nor I_25783 (I441901,I1198503,I1198512);
nor I_25784 (I441451,I441901,I441884);
not I_25785 (I441932,I441901);
nand I_25786 (I441454,I441661,I441932);
DFFARX1 I_25787 (I441901,I3563,I441477,I441466,);
DFFARX1 I_25788 (I441901,I3563,I441477,I441463,);
not I_25789 (I442021,I3570);
DFFARX1 I_25790 (I351261,I3563,I442021,I442047,);
DFFARX1 I_25791 (I442047,I3563,I442021,I442064,);
not I_25792 (I442013,I442064);
not I_25793 (I442086,I442047);
nand I_25794 (I442103,I351240,I351264);
and I_25795 (I442120,I442103,I351267);
DFFARX1 I_25796 (I442120,I3563,I442021,I442146,);
not I_25797 (I442154,I442146);
DFFARX1 I_25798 (I351249,I3563,I442021,I442180,);
and I_25799 (I442188,I442180,I351255);
nand I_25800 (I442205,I442180,I351255);
nand I_25801 (I441992,I442154,I442205);
DFFARX1 I_25802 (I351243,I3563,I442021,I442245,);
nor I_25803 (I442253,I442245,I442188);
DFFARX1 I_25804 (I442253,I3563,I442021,I441986,);
nor I_25805 (I442001,I442245,I442146);
nand I_25806 (I442298,I351252,I351240);
and I_25807 (I442315,I442298,I351246);
DFFARX1 I_25808 (I442315,I3563,I442021,I442341,);
nor I_25809 (I441989,I442341,I442245);
not I_25810 (I442363,I442341);
nor I_25811 (I442380,I442363,I442154);
nor I_25812 (I442397,I442086,I442380);
DFFARX1 I_25813 (I442397,I3563,I442021,I442004,);
nor I_25814 (I442428,I442363,I442245);
nor I_25815 (I442445,I351258,I351240);
nor I_25816 (I441995,I442445,I442428);
not I_25817 (I442476,I442445);
nand I_25818 (I441998,I442205,I442476);
DFFARX1 I_25819 (I442445,I3563,I442021,I442010,);
DFFARX1 I_25820 (I442445,I3563,I442021,I442007,);
not I_25821 (I442565,I3570);
DFFARX1 I_25822 (I1152266,I3563,I442565,I442591,);
DFFARX1 I_25823 (I442591,I3563,I442565,I442608,);
not I_25824 (I442557,I442608);
not I_25825 (I442630,I442591);
nand I_25826 (I442647,I1152278,I1152266);
and I_25827 (I442664,I442647,I1152269);
DFFARX1 I_25828 (I442664,I3563,I442565,I442690,);
not I_25829 (I442698,I442690);
DFFARX1 I_25830 (I1152287,I3563,I442565,I442724,);
and I_25831 (I442732,I442724,I1152263);
nand I_25832 (I442749,I442724,I1152263);
nand I_25833 (I442536,I442698,I442749);
DFFARX1 I_25834 (I1152281,I3563,I442565,I442789,);
nor I_25835 (I442797,I442789,I442732);
DFFARX1 I_25836 (I442797,I3563,I442565,I442530,);
nor I_25837 (I442545,I442789,I442690);
nand I_25838 (I442842,I1152275,I1152272);
and I_25839 (I442859,I442842,I1152284);
DFFARX1 I_25840 (I442859,I3563,I442565,I442885,);
nor I_25841 (I442533,I442885,I442789);
not I_25842 (I442907,I442885);
nor I_25843 (I442924,I442907,I442698);
nor I_25844 (I442941,I442630,I442924);
DFFARX1 I_25845 (I442941,I3563,I442565,I442548,);
nor I_25846 (I442972,I442907,I442789);
nor I_25847 (I442989,I1152263,I1152272);
nor I_25848 (I442539,I442989,I442972);
not I_25849 (I443020,I442989);
nand I_25850 (I442542,I442749,I443020);
DFFARX1 I_25851 (I442989,I3563,I442565,I442554,);
DFFARX1 I_25852 (I442989,I3563,I442565,I442551,);
not I_25853 (I443109,I3570);
DFFARX1 I_25854 (I748584,I3563,I443109,I443135,);
DFFARX1 I_25855 (I443135,I3563,I443109,I443152,);
not I_25856 (I443101,I443152);
not I_25857 (I443174,I443135);
nand I_25858 (I443191,I748605,I748596);
and I_25859 (I443208,I443191,I748584);
DFFARX1 I_25860 (I443208,I3563,I443109,I443234,);
not I_25861 (I443242,I443234);
DFFARX1 I_25862 (I748590,I3563,I443109,I443268,);
and I_25863 (I443276,I443268,I748587);
nand I_25864 (I443293,I443268,I748587);
nand I_25865 (I443080,I443242,I443293);
DFFARX1 I_25866 (I748581,I3563,I443109,I443333,);
nor I_25867 (I443341,I443333,I443276);
DFFARX1 I_25868 (I443341,I3563,I443109,I443074,);
nor I_25869 (I443089,I443333,I443234);
nand I_25870 (I443386,I748581,I748593);
and I_25871 (I443403,I443386,I748602);
DFFARX1 I_25872 (I443403,I3563,I443109,I443429,);
nor I_25873 (I443077,I443429,I443333);
not I_25874 (I443451,I443429);
nor I_25875 (I443468,I443451,I443242);
nor I_25876 (I443485,I443174,I443468);
DFFARX1 I_25877 (I443485,I3563,I443109,I443092,);
nor I_25878 (I443516,I443451,I443333);
nor I_25879 (I443533,I748599,I748593);
nor I_25880 (I443083,I443533,I443516);
not I_25881 (I443564,I443533);
nand I_25882 (I443086,I443293,I443564);
DFFARX1 I_25883 (I443533,I3563,I443109,I443098,);
DFFARX1 I_25884 (I443533,I3563,I443109,I443095,);
not I_25885 (I443653,I3570);
DFFARX1 I_25886 (I933615,I3563,I443653,I443679,);
DFFARX1 I_25887 (I443679,I3563,I443653,I443696,);
not I_25888 (I443645,I443696);
not I_25889 (I443718,I443679);
nand I_25890 (I443735,I933630,I933618);
and I_25891 (I443752,I443735,I933609);
DFFARX1 I_25892 (I443752,I3563,I443653,I443778,);
not I_25893 (I443786,I443778);
DFFARX1 I_25894 (I933621,I3563,I443653,I443812,);
and I_25895 (I443820,I443812,I933612);
nand I_25896 (I443837,I443812,I933612);
nand I_25897 (I443624,I443786,I443837);
DFFARX1 I_25898 (I933627,I3563,I443653,I443877,);
nor I_25899 (I443885,I443877,I443820);
DFFARX1 I_25900 (I443885,I3563,I443653,I443618,);
nor I_25901 (I443633,I443877,I443778);
nand I_25902 (I443930,I933636,I933624);
and I_25903 (I443947,I443930,I933633);
DFFARX1 I_25904 (I443947,I3563,I443653,I443973,);
nor I_25905 (I443621,I443973,I443877);
not I_25906 (I443995,I443973);
nor I_25907 (I444012,I443995,I443786);
nor I_25908 (I444029,I443718,I444012);
DFFARX1 I_25909 (I444029,I3563,I443653,I443636,);
nor I_25910 (I444060,I443995,I443877);
nor I_25911 (I444077,I933609,I933624);
nor I_25912 (I443627,I444077,I444060);
not I_25913 (I444108,I444077);
nand I_25914 (I443630,I443837,I444108);
DFFARX1 I_25915 (I444077,I3563,I443653,I443642,);
DFFARX1 I_25916 (I444077,I3563,I443653,I443639,);
not I_25917 (I444197,I3570);
DFFARX1 I_25918 (I1306845,I3563,I444197,I444223,);
DFFARX1 I_25919 (I444223,I3563,I444197,I444240,);
not I_25920 (I444189,I444240);
not I_25921 (I444262,I444223);
nand I_25922 (I444279,I1306842,I1306839);
and I_25923 (I444296,I444279,I1306827);
DFFARX1 I_25924 (I444296,I3563,I444197,I444322,);
not I_25925 (I444330,I444322);
DFFARX1 I_25926 (I1306851,I3563,I444197,I444356,);
and I_25927 (I444364,I444356,I1306836);
nand I_25928 (I444381,I444356,I1306836);
nand I_25929 (I444168,I444330,I444381);
DFFARX1 I_25930 (I1306830,I3563,I444197,I444421,);
nor I_25931 (I444429,I444421,I444364);
DFFARX1 I_25932 (I444429,I3563,I444197,I444162,);
nor I_25933 (I444177,I444421,I444322);
nand I_25934 (I444474,I1306827,I1306833);
and I_25935 (I444491,I444474,I1306848);
DFFARX1 I_25936 (I444491,I3563,I444197,I444517,);
nor I_25937 (I444165,I444517,I444421);
not I_25938 (I444539,I444517);
nor I_25939 (I444556,I444539,I444330);
nor I_25940 (I444573,I444262,I444556);
DFFARX1 I_25941 (I444573,I3563,I444197,I444180,);
nor I_25942 (I444604,I444539,I444421);
nor I_25943 (I444621,I1306830,I1306833);
nor I_25944 (I444171,I444621,I444604);
not I_25945 (I444652,I444621);
nand I_25946 (I444174,I444381,I444652);
DFFARX1 I_25947 (I444621,I3563,I444197,I444186,);
DFFARX1 I_25948 (I444621,I3563,I444197,I444183,);
not I_25949 (I444741,I3570);
DFFARX1 I_25950 (I989171,I3563,I444741,I444767,);
DFFARX1 I_25951 (I444767,I3563,I444741,I444784,);
not I_25952 (I444733,I444784);
not I_25953 (I444806,I444767);
nand I_25954 (I444823,I989186,I989174);
and I_25955 (I444840,I444823,I989165);
DFFARX1 I_25956 (I444840,I3563,I444741,I444866,);
not I_25957 (I444874,I444866);
DFFARX1 I_25958 (I989177,I3563,I444741,I444900,);
and I_25959 (I444908,I444900,I989168);
nand I_25960 (I444925,I444900,I989168);
nand I_25961 (I444712,I444874,I444925);
DFFARX1 I_25962 (I989183,I3563,I444741,I444965,);
nor I_25963 (I444973,I444965,I444908);
DFFARX1 I_25964 (I444973,I3563,I444741,I444706,);
nor I_25965 (I444721,I444965,I444866);
nand I_25966 (I445018,I989192,I989180);
and I_25967 (I445035,I445018,I989189);
DFFARX1 I_25968 (I445035,I3563,I444741,I445061,);
nor I_25969 (I444709,I445061,I444965);
not I_25970 (I445083,I445061);
nor I_25971 (I445100,I445083,I444874);
nor I_25972 (I445117,I444806,I445100);
DFFARX1 I_25973 (I445117,I3563,I444741,I444724,);
nor I_25974 (I445148,I445083,I444965);
nor I_25975 (I445165,I989165,I989180);
nor I_25976 (I444715,I445165,I445148);
not I_25977 (I445196,I445165);
nand I_25978 (I444718,I444925,I445196);
DFFARX1 I_25979 (I445165,I3563,I444741,I444730,);
DFFARX1 I_25980 (I445165,I3563,I444741,I444727,);
not I_25981 (I445285,I3570);
DFFARX1 I_25982 (I137284,I3563,I445285,I445311,);
DFFARX1 I_25983 (I445311,I3563,I445285,I445328,);
not I_25984 (I445277,I445328);
not I_25985 (I445350,I445311);
nand I_25986 (I445367,I137299,I137278);
and I_25987 (I445384,I445367,I137281);
DFFARX1 I_25988 (I445384,I3563,I445285,I445410,);
not I_25989 (I445418,I445410);
DFFARX1 I_25990 (I137287,I3563,I445285,I445444,);
and I_25991 (I445452,I445444,I137281);
nand I_25992 (I445469,I445444,I137281);
nand I_25993 (I445256,I445418,I445469);
DFFARX1 I_25994 (I137296,I3563,I445285,I445509,);
nor I_25995 (I445517,I445509,I445452);
DFFARX1 I_25996 (I445517,I3563,I445285,I445250,);
nor I_25997 (I445265,I445509,I445410);
nand I_25998 (I445562,I137278,I137293);
and I_25999 (I445579,I445562,I137290);
DFFARX1 I_26000 (I445579,I3563,I445285,I445605,);
nor I_26001 (I445253,I445605,I445509);
not I_26002 (I445627,I445605);
nor I_26003 (I445644,I445627,I445418);
nor I_26004 (I445661,I445350,I445644);
DFFARX1 I_26005 (I445661,I3563,I445285,I445268,);
nor I_26006 (I445692,I445627,I445509);
nor I_26007 (I445709,I137302,I137293);
nor I_26008 (I445259,I445709,I445692);
not I_26009 (I445740,I445709);
nand I_26010 (I445262,I445469,I445740);
DFFARX1 I_26011 (I445709,I3563,I445285,I445274,);
DFFARX1 I_26012 (I445709,I3563,I445285,I445271,);
not I_26013 (I445829,I3570);
DFFARX1 I_26014 (I114623,I3563,I445829,I445855,);
DFFARX1 I_26015 (I445855,I3563,I445829,I445872,);
not I_26016 (I445821,I445872);
not I_26017 (I445894,I445855);
nand I_26018 (I445911,I114638,I114617);
and I_26019 (I445928,I445911,I114620);
DFFARX1 I_26020 (I445928,I3563,I445829,I445954,);
not I_26021 (I445962,I445954);
DFFARX1 I_26022 (I114626,I3563,I445829,I445988,);
and I_26023 (I445996,I445988,I114620);
nand I_26024 (I446013,I445988,I114620);
nand I_26025 (I445800,I445962,I446013);
DFFARX1 I_26026 (I114635,I3563,I445829,I446053,);
nor I_26027 (I446061,I446053,I445996);
DFFARX1 I_26028 (I446061,I3563,I445829,I445794,);
nor I_26029 (I445809,I446053,I445954);
nand I_26030 (I446106,I114617,I114632);
and I_26031 (I446123,I446106,I114629);
DFFARX1 I_26032 (I446123,I3563,I445829,I446149,);
nor I_26033 (I445797,I446149,I446053);
not I_26034 (I446171,I446149);
nor I_26035 (I446188,I446171,I445962);
nor I_26036 (I446205,I445894,I446188);
DFFARX1 I_26037 (I446205,I3563,I445829,I445812,);
nor I_26038 (I446236,I446171,I446053);
nor I_26039 (I446253,I114641,I114632);
nor I_26040 (I445803,I446253,I446236);
not I_26041 (I446284,I446253);
nand I_26042 (I445806,I446013,I446284);
DFFARX1 I_26043 (I446253,I3563,I445829,I445818,);
DFFARX1 I_26044 (I446253,I3563,I445829,I445815,);
not I_26045 (I446373,I3570);
DFFARX1 I_26046 (I1171918,I3563,I446373,I446399,);
DFFARX1 I_26047 (I446399,I3563,I446373,I446416,);
not I_26048 (I446365,I446416);
not I_26049 (I446438,I446399);
nand I_26050 (I446455,I1171930,I1171918);
and I_26051 (I446472,I446455,I1171921);
DFFARX1 I_26052 (I446472,I3563,I446373,I446498,);
not I_26053 (I446506,I446498);
DFFARX1 I_26054 (I1171939,I3563,I446373,I446532,);
and I_26055 (I446540,I446532,I1171915);
nand I_26056 (I446557,I446532,I1171915);
nand I_26057 (I446344,I446506,I446557);
DFFARX1 I_26058 (I1171933,I3563,I446373,I446597,);
nor I_26059 (I446605,I446597,I446540);
DFFARX1 I_26060 (I446605,I3563,I446373,I446338,);
nor I_26061 (I446353,I446597,I446498);
nand I_26062 (I446650,I1171927,I1171924);
and I_26063 (I446667,I446650,I1171936);
DFFARX1 I_26064 (I446667,I3563,I446373,I446693,);
nor I_26065 (I446341,I446693,I446597);
not I_26066 (I446715,I446693);
nor I_26067 (I446732,I446715,I446506);
nor I_26068 (I446749,I446438,I446732);
DFFARX1 I_26069 (I446749,I3563,I446373,I446356,);
nor I_26070 (I446780,I446715,I446597);
nor I_26071 (I446797,I1171915,I1171924);
nor I_26072 (I446347,I446797,I446780);
not I_26073 (I446828,I446797);
nand I_26074 (I446350,I446557,I446828);
DFFARX1 I_26075 (I446797,I3563,I446373,I446362,);
DFFARX1 I_26076 (I446797,I3563,I446373,I446359,);
not I_26077 (I446917,I3570);
DFFARX1 I_26078 (I883267,I3563,I446917,I446943,);
DFFARX1 I_26079 (I446943,I3563,I446917,I446960,);
not I_26080 (I446909,I446960);
not I_26081 (I446982,I446943);
nand I_26082 (I446999,I883261,I883258);
and I_26083 (I447016,I446999,I883273);
DFFARX1 I_26084 (I447016,I3563,I446917,I447042,);
not I_26085 (I447050,I447042);
DFFARX1 I_26086 (I883261,I3563,I446917,I447076,);
and I_26087 (I447084,I447076,I883255);
nand I_26088 (I447101,I447076,I883255);
nand I_26089 (I446888,I447050,I447101);
DFFARX1 I_26090 (I883255,I3563,I446917,I447141,);
nor I_26091 (I447149,I447141,I447084);
DFFARX1 I_26092 (I447149,I3563,I446917,I446882,);
nor I_26093 (I446897,I447141,I447042);
nand I_26094 (I447194,I883270,I883264);
and I_26095 (I447211,I447194,I883258);
DFFARX1 I_26096 (I447211,I3563,I446917,I447237,);
nor I_26097 (I446885,I447237,I447141);
not I_26098 (I447259,I447237);
nor I_26099 (I447276,I447259,I447050);
nor I_26100 (I447293,I446982,I447276);
DFFARX1 I_26101 (I447293,I3563,I446917,I446900,);
nor I_26102 (I447324,I447259,I447141);
nor I_26103 (I447341,I883276,I883264);
nor I_26104 (I446891,I447341,I447324);
not I_26105 (I447372,I447341);
nand I_26106 (I446894,I447101,I447372);
DFFARX1 I_26107 (I447341,I3563,I446917,I446906,);
DFFARX1 I_26108 (I447341,I3563,I446917,I446903,);
not I_26109 (I447461,I3570);
DFFARX1 I_26110 (I1055635,I3563,I447461,I447487,);
DFFARX1 I_26111 (I447487,I3563,I447461,I447504,);
not I_26112 (I447453,I447504);
not I_26113 (I447526,I447487);
nand I_26114 (I447543,I1055635,I1055653);
and I_26115 (I447560,I447543,I1055647);
DFFARX1 I_26116 (I447560,I3563,I447461,I447586,);
not I_26117 (I447594,I447586);
DFFARX1 I_26118 (I1055641,I3563,I447461,I447620,);
and I_26119 (I447628,I447620,I1055650);
nand I_26120 (I447645,I447620,I1055650);
nand I_26121 (I447432,I447594,I447645);
DFFARX1 I_26122 (I1055638,I3563,I447461,I447685,);
nor I_26123 (I447693,I447685,I447628);
DFFARX1 I_26124 (I447693,I3563,I447461,I447426,);
nor I_26125 (I447441,I447685,I447586);
nand I_26126 (I447738,I1055638,I1055656);
and I_26127 (I447755,I447738,I1055641);
DFFARX1 I_26128 (I447755,I3563,I447461,I447781,);
nor I_26129 (I447429,I447781,I447685);
not I_26130 (I447803,I447781);
nor I_26131 (I447820,I447803,I447594);
nor I_26132 (I447837,I447526,I447820);
DFFARX1 I_26133 (I447837,I3563,I447461,I447444,);
nor I_26134 (I447868,I447803,I447685);
nor I_26135 (I447885,I1055644,I1055656);
nor I_26136 (I447435,I447885,I447868);
not I_26137 (I447916,I447885);
nand I_26138 (I447438,I447645,I447916);
DFFARX1 I_26139 (I447885,I3563,I447461,I447450,);
DFFARX1 I_26140 (I447885,I3563,I447461,I447447,);
not I_26141 (I448005,I3570);
DFFARX1 I_26142 (I1200818,I3563,I448005,I448031,);
DFFARX1 I_26143 (I448031,I3563,I448005,I448048,);
not I_26144 (I447997,I448048);
not I_26145 (I448070,I448031);
nand I_26146 (I448087,I1200830,I1200818);
and I_26147 (I448104,I448087,I1200821);
DFFARX1 I_26148 (I448104,I3563,I448005,I448130,);
not I_26149 (I448138,I448130);
DFFARX1 I_26150 (I1200839,I3563,I448005,I448164,);
and I_26151 (I448172,I448164,I1200815);
nand I_26152 (I448189,I448164,I1200815);
nand I_26153 (I447976,I448138,I448189);
DFFARX1 I_26154 (I1200833,I3563,I448005,I448229,);
nor I_26155 (I448237,I448229,I448172);
DFFARX1 I_26156 (I448237,I3563,I448005,I447970,);
nor I_26157 (I447985,I448229,I448130);
nand I_26158 (I448282,I1200827,I1200824);
and I_26159 (I448299,I448282,I1200836);
DFFARX1 I_26160 (I448299,I3563,I448005,I448325,);
nor I_26161 (I447973,I448325,I448229);
not I_26162 (I448347,I448325);
nor I_26163 (I448364,I448347,I448138);
nor I_26164 (I448381,I448070,I448364);
DFFARX1 I_26165 (I448381,I3563,I448005,I447988,);
nor I_26166 (I448412,I448347,I448229);
nor I_26167 (I448429,I1200815,I1200824);
nor I_26168 (I447979,I448429,I448412);
not I_26169 (I448460,I448429);
nand I_26170 (I447982,I448189,I448460);
DFFARX1 I_26171 (I448429,I3563,I448005,I447994,);
DFFARX1 I_26172 (I448429,I3563,I448005,I447991,);
not I_26173 (I448549,I3570);
DFFARX1 I_26174 (I1364280,I3563,I448549,I448575,);
DFFARX1 I_26175 (I448575,I3563,I448549,I448592,);
not I_26176 (I448541,I448592);
not I_26177 (I448614,I448575);
nand I_26178 (I448631,I1364256,I1364277);
and I_26179 (I448648,I448631,I1364274);
DFFARX1 I_26180 (I448648,I3563,I448549,I448674,);
not I_26181 (I448682,I448674);
DFFARX1 I_26182 (I1364253,I3563,I448549,I448708,);
and I_26183 (I448716,I448708,I1364265);
nand I_26184 (I448733,I448708,I1364265);
nand I_26185 (I448520,I448682,I448733);
DFFARX1 I_26186 (I1364268,I3563,I448549,I448773,);
nor I_26187 (I448781,I448773,I448716);
DFFARX1 I_26188 (I448781,I3563,I448549,I448514,);
nor I_26189 (I448529,I448773,I448674);
nand I_26190 (I448826,I1364271,I1364259);
and I_26191 (I448843,I448826,I1364262);
DFFARX1 I_26192 (I448843,I3563,I448549,I448869,);
nor I_26193 (I448517,I448869,I448773);
not I_26194 (I448891,I448869);
nor I_26195 (I448908,I448891,I448682);
nor I_26196 (I448925,I448614,I448908);
DFFARX1 I_26197 (I448925,I3563,I448549,I448532,);
nor I_26198 (I448956,I448891,I448773);
nor I_26199 (I448973,I1364253,I1364259);
nor I_26200 (I448523,I448973,I448956);
not I_26201 (I449004,I448973);
nand I_26202 (I448526,I448733,I449004);
DFFARX1 I_26203 (I448973,I3563,I448549,I448538,);
DFFARX1 I_26204 (I448973,I3563,I448549,I448535,);
not I_26205 (I449093,I3570);
DFFARX1 I_26206 (I832675,I3563,I449093,I449119,);
DFFARX1 I_26207 (I449119,I3563,I449093,I449136,);
not I_26208 (I449085,I449136);
not I_26209 (I449158,I449119);
nand I_26210 (I449175,I832669,I832666);
and I_26211 (I449192,I449175,I832681);
DFFARX1 I_26212 (I449192,I3563,I449093,I449218,);
not I_26213 (I449226,I449218);
DFFARX1 I_26214 (I832669,I3563,I449093,I449252,);
and I_26215 (I449260,I449252,I832663);
nand I_26216 (I449277,I449252,I832663);
nand I_26217 (I449064,I449226,I449277);
DFFARX1 I_26218 (I832663,I3563,I449093,I449317,);
nor I_26219 (I449325,I449317,I449260);
DFFARX1 I_26220 (I449325,I3563,I449093,I449058,);
nor I_26221 (I449073,I449317,I449218);
nand I_26222 (I449370,I832678,I832672);
and I_26223 (I449387,I449370,I832666);
DFFARX1 I_26224 (I449387,I3563,I449093,I449413,);
nor I_26225 (I449061,I449413,I449317);
not I_26226 (I449435,I449413);
nor I_26227 (I449452,I449435,I449226);
nor I_26228 (I449469,I449158,I449452);
DFFARX1 I_26229 (I449469,I3563,I449093,I449076,);
nor I_26230 (I449500,I449435,I449317);
nor I_26231 (I449517,I832684,I832672);
nor I_26232 (I449067,I449517,I449500);
not I_26233 (I449548,I449517);
nand I_26234 (I449070,I449277,I449548);
DFFARX1 I_26235 (I449517,I3563,I449093,I449082,);
DFFARX1 I_26236 (I449517,I3563,I449093,I449079,);
not I_26237 (I449637,I3570);
DFFARX1 I_26238 (I1385105,I3563,I449637,I449663,);
DFFARX1 I_26239 (I449663,I3563,I449637,I449680,);
not I_26240 (I449629,I449680);
not I_26241 (I449702,I449663);
nand I_26242 (I449719,I1385081,I1385102);
and I_26243 (I449736,I449719,I1385099);
DFFARX1 I_26244 (I449736,I3563,I449637,I449762,);
not I_26245 (I449770,I449762);
DFFARX1 I_26246 (I1385078,I3563,I449637,I449796,);
and I_26247 (I449804,I449796,I1385090);
nand I_26248 (I449821,I449796,I1385090);
nand I_26249 (I449608,I449770,I449821);
DFFARX1 I_26250 (I1385093,I3563,I449637,I449861,);
nor I_26251 (I449869,I449861,I449804);
DFFARX1 I_26252 (I449869,I3563,I449637,I449602,);
nor I_26253 (I449617,I449861,I449762);
nand I_26254 (I449914,I1385096,I1385084);
and I_26255 (I449931,I449914,I1385087);
DFFARX1 I_26256 (I449931,I3563,I449637,I449957,);
nor I_26257 (I449605,I449957,I449861);
not I_26258 (I449979,I449957);
nor I_26259 (I449996,I449979,I449770);
nor I_26260 (I450013,I449702,I449996);
DFFARX1 I_26261 (I450013,I3563,I449637,I449620,);
nor I_26262 (I450044,I449979,I449861);
nor I_26263 (I450061,I1385078,I1385084);
nor I_26264 (I449611,I450061,I450044);
not I_26265 (I450092,I450061);
nand I_26266 (I449614,I449821,I450092);
DFFARX1 I_26267 (I450061,I3563,I449637,I449626,);
DFFARX1 I_26268 (I450061,I3563,I449637,I449623,);
not I_26269 (I450181,I3570);
DFFARX1 I_26270 (I689050,I3563,I450181,I450207,);
DFFARX1 I_26271 (I450207,I3563,I450181,I450224,);
not I_26272 (I450173,I450224);
not I_26273 (I450246,I450207);
nand I_26274 (I450263,I689071,I689062);
and I_26275 (I450280,I450263,I689050);
DFFARX1 I_26276 (I450280,I3563,I450181,I450306,);
not I_26277 (I450314,I450306);
DFFARX1 I_26278 (I689056,I3563,I450181,I450340,);
and I_26279 (I450348,I450340,I689053);
nand I_26280 (I450365,I450340,I689053);
nand I_26281 (I450152,I450314,I450365);
DFFARX1 I_26282 (I689047,I3563,I450181,I450405,);
nor I_26283 (I450413,I450405,I450348);
DFFARX1 I_26284 (I450413,I3563,I450181,I450146,);
nor I_26285 (I450161,I450405,I450306);
nand I_26286 (I450458,I689047,I689059);
and I_26287 (I450475,I450458,I689068);
DFFARX1 I_26288 (I450475,I3563,I450181,I450501,);
nor I_26289 (I450149,I450501,I450405);
not I_26290 (I450523,I450501);
nor I_26291 (I450540,I450523,I450314);
nor I_26292 (I450557,I450246,I450540);
DFFARX1 I_26293 (I450557,I3563,I450181,I450164,);
nor I_26294 (I450588,I450523,I450405);
nor I_26295 (I450605,I689065,I689059);
nor I_26296 (I450155,I450605,I450588);
not I_26297 (I450636,I450605);
nand I_26298 (I450158,I450365,I450636);
DFFARX1 I_26299 (I450605,I3563,I450181,I450170,);
DFFARX1 I_26300 (I450605,I3563,I450181,I450167,);
not I_26301 (I450725,I3570);
DFFARX1 I_26302 (I1162092,I3563,I450725,I450751,);
DFFARX1 I_26303 (I450751,I3563,I450725,I450768,);
not I_26304 (I450717,I450768);
not I_26305 (I450790,I450751);
nand I_26306 (I450807,I1162104,I1162092);
and I_26307 (I450824,I450807,I1162095);
DFFARX1 I_26308 (I450824,I3563,I450725,I450850,);
not I_26309 (I450858,I450850);
DFFARX1 I_26310 (I1162113,I3563,I450725,I450884,);
and I_26311 (I450892,I450884,I1162089);
nand I_26312 (I450909,I450884,I1162089);
nand I_26313 (I450696,I450858,I450909);
DFFARX1 I_26314 (I1162107,I3563,I450725,I450949,);
nor I_26315 (I450957,I450949,I450892);
DFFARX1 I_26316 (I450957,I3563,I450725,I450690,);
nor I_26317 (I450705,I450949,I450850);
nand I_26318 (I451002,I1162101,I1162098);
and I_26319 (I451019,I451002,I1162110);
DFFARX1 I_26320 (I451019,I3563,I450725,I451045,);
nor I_26321 (I450693,I451045,I450949);
not I_26322 (I451067,I451045);
nor I_26323 (I451084,I451067,I450858);
nor I_26324 (I451101,I450790,I451084);
DFFARX1 I_26325 (I451101,I3563,I450725,I450708,);
nor I_26326 (I451132,I451067,I450949);
nor I_26327 (I451149,I1162089,I1162098);
nor I_26328 (I450699,I451149,I451132);
not I_26329 (I451180,I451149);
nand I_26330 (I450702,I450909,I451180);
DFFARX1 I_26331 (I451149,I3563,I450725,I450714,);
DFFARX1 I_26332 (I451149,I3563,I450725,I450711,);
not I_26333 (I451269,I3570);
DFFARX1 I_26334 (I113042,I3563,I451269,I451295,);
DFFARX1 I_26335 (I451295,I3563,I451269,I451312,);
not I_26336 (I451261,I451312);
not I_26337 (I451334,I451295);
nand I_26338 (I451351,I113057,I113036);
and I_26339 (I451368,I451351,I113039);
DFFARX1 I_26340 (I451368,I3563,I451269,I451394,);
not I_26341 (I451402,I451394);
DFFARX1 I_26342 (I113045,I3563,I451269,I451428,);
and I_26343 (I451436,I451428,I113039);
nand I_26344 (I451453,I451428,I113039);
nand I_26345 (I451240,I451402,I451453);
DFFARX1 I_26346 (I113054,I3563,I451269,I451493,);
nor I_26347 (I451501,I451493,I451436);
DFFARX1 I_26348 (I451501,I3563,I451269,I451234,);
nor I_26349 (I451249,I451493,I451394);
nand I_26350 (I451546,I113036,I113051);
and I_26351 (I451563,I451546,I113048);
DFFARX1 I_26352 (I451563,I3563,I451269,I451589,);
nor I_26353 (I451237,I451589,I451493);
not I_26354 (I451611,I451589);
nor I_26355 (I451628,I451611,I451402);
nor I_26356 (I451645,I451334,I451628);
DFFARX1 I_26357 (I451645,I3563,I451269,I451252,);
nor I_26358 (I451676,I451611,I451493);
nor I_26359 (I451693,I113060,I113051);
nor I_26360 (I451243,I451693,I451676);
not I_26361 (I451724,I451693);
nand I_26362 (I451246,I451453,I451724);
DFFARX1 I_26363 (I451693,I3563,I451269,I451258,);
DFFARX1 I_26364 (I451693,I3563,I451269,I451255,);
not I_26365 (I451813,I3570);
DFFARX1 I_26366 (I906982,I3563,I451813,I451839,);
DFFARX1 I_26367 (I451839,I3563,I451813,I451856,);
not I_26368 (I451805,I451856);
not I_26369 (I451878,I451839);
nand I_26370 (I451895,I906976,I906973);
and I_26371 (I451912,I451895,I906988);
DFFARX1 I_26372 (I451912,I3563,I451813,I451938,);
not I_26373 (I451946,I451938);
DFFARX1 I_26374 (I906976,I3563,I451813,I451972,);
and I_26375 (I451980,I451972,I906970);
nand I_26376 (I451997,I451972,I906970);
nand I_26377 (I451784,I451946,I451997);
DFFARX1 I_26378 (I906970,I3563,I451813,I452037,);
nor I_26379 (I452045,I452037,I451980);
DFFARX1 I_26380 (I452045,I3563,I451813,I451778,);
nor I_26381 (I451793,I452037,I451938);
nand I_26382 (I452090,I906985,I906979);
and I_26383 (I452107,I452090,I906973);
DFFARX1 I_26384 (I452107,I3563,I451813,I452133,);
nor I_26385 (I451781,I452133,I452037);
not I_26386 (I452155,I452133);
nor I_26387 (I452172,I452155,I451946);
nor I_26388 (I452189,I451878,I452172);
DFFARX1 I_26389 (I452189,I3563,I451813,I451796,);
nor I_26390 (I452220,I452155,I452037);
nor I_26391 (I452237,I906991,I906979);
nor I_26392 (I451787,I452237,I452220);
not I_26393 (I452268,I452237);
nand I_26394 (I451790,I451997,I452268);
DFFARX1 I_26395 (I452237,I3563,I451813,I451802,);
DFFARX1 I_26396 (I452237,I3563,I451813,I451799,);
not I_26397 (I452357,I3570);
DFFARX1 I_26398 (I811008,I3563,I452357,I452383,);
DFFARX1 I_26399 (I452383,I3563,I452357,I452400,);
not I_26400 (I452349,I452400);
not I_26401 (I452422,I452383);
nand I_26402 (I452439,I811029,I811020);
and I_26403 (I452456,I452439,I811008);
DFFARX1 I_26404 (I452456,I3563,I452357,I452482,);
not I_26405 (I452490,I452482);
DFFARX1 I_26406 (I811014,I3563,I452357,I452516,);
and I_26407 (I452524,I452516,I811011);
nand I_26408 (I452541,I452516,I811011);
nand I_26409 (I452328,I452490,I452541);
DFFARX1 I_26410 (I811005,I3563,I452357,I452581,);
nor I_26411 (I452589,I452581,I452524);
DFFARX1 I_26412 (I452589,I3563,I452357,I452322,);
nor I_26413 (I452337,I452581,I452482);
nand I_26414 (I452634,I811005,I811017);
and I_26415 (I452651,I452634,I811026);
DFFARX1 I_26416 (I452651,I3563,I452357,I452677,);
nor I_26417 (I452325,I452677,I452581);
not I_26418 (I452699,I452677);
nor I_26419 (I452716,I452699,I452490);
nor I_26420 (I452733,I452422,I452716);
DFFARX1 I_26421 (I452733,I3563,I452357,I452340,);
nor I_26422 (I452764,I452699,I452581);
nor I_26423 (I452781,I811023,I811017);
nor I_26424 (I452331,I452781,I452764);
not I_26425 (I452812,I452781);
nand I_26426 (I452334,I452541,I452812);
DFFARX1 I_26427 (I452781,I3563,I452357,I452346,);
DFFARX1 I_26428 (I452781,I3563,I452357,I452343,);
not I_26429 (I452901,I3570);
DFFARX1 I_26430 (I69301,I3563,I452901,I452927,);
DFFARX1 I_26431 (I452927,I3563,I452901,I452944,);
not I_26432 (I452893,I452944);
not I_26433 (I452966,I452927);
nand I_26434 (I452983,I69316,I69295);
and I_26435 (I453000,I452983,I69298);
DFFARX1 I_26436 (I453000,I3563,I452901,I453026,);
not I_26437 (I453034,I453026);
DFFARX1 I_26438 (I69304,I3563,I452901,I453060,);
and I_26439 (I453068,I453060,I69298);
nand I_26440 (I453085,I453060,I69298);
nand I_26441 (I452872,I453034,I453085);
DFFARX1 I_26442 (I69313,I3563,I452901,I453125,);
nor I_26443 (I453133,I453125,I453068);
DFFARX1 I_26444 (I453133,I3563,I452901,I452866,);
nor I_26445 (I452881,I453125,I453026);
nand I_26446 (I453178,I69295,I69310);
and I_26447 (I453195,I453178,I69307);
DFFARX1 I_26448 (I453195,I3563,I452901,I453221,);
nor I_26449 (I452869,I453221,I453125);
not I_26450 (I453243,I453221);
nor I_26451 (I453260,I453243,I453034);
nor I_26452 (I453277,I452966,I453260);
DFFARX1 I_26453 (I453277,I3563,I452901,I452884,);
nor I_26454 (I453308,I453243,I453125);
nor I_26455 (I453325,I69319,I69310);
nor I_26456 (I452875,I453325,I453308);
not I_26457 (I453356,I453325);
nand I_26458 (I452878,I453085,I453356);
DFFARX1 I_26459 (I453325,I3563,I452901,I452890,);
DFFARX1 I_26460 (I453325,I3563,I452901,I452887,);
not I_26461 (I453445,I3570);
DFFARX1 I_26462 (I539994,I3563,I453445,I453471,);
DFFARX1 I_26463 (I453471,I3563,I453445,I453488,);
not I_26464 (I453437,I453488);
not I_26465 (I453510,I453471);
nand I_26466 (I453527,I539997,I540015);
and I_26467 (I453544,I453527,I540003);
DFFARX1 I_26468 (I453544,I3563,I453445,I453570,);
not I_26469 (I453578,I453570);
DFFARX1 I_26470 (I539994,I3563,I453445,I453604,);
and I_26471 (I453612,I453604,I540012);
nand I_26472 (I453629,I453604,I540012);
nand I_26473 (I453416,I453578,I453629);
DFFARX1 I_26474 (I540006,I3563,I453445,I453669,);
nor I_26475 (I453677,I453669,I453612);
DFFARX1 I_26476 (I453677,I3563,I453445,I453410,);
nor I_26477 (I453425,I453669,I453570);
nand I_26478 (I453722,I540009,I539991);
and I_26479 (I453739,I453722,I540000);
DFFARX1 I_26480 (I453739,I3563,I453445,I453765,);
nor I_26481 (I453413,I453765,I453669);
not I_26482 (I453787,I453765);
nor I_26483 (I453804,I453787,I453578);
nor I_26484 (I453821,I453510,I453804);
DFFARX1 I_26485 (I453821,I3563,I453445,I453428,);
nor I_26486 (I453852,I453787,I453669);
nor I_26487 (I453869,I539991,I539991);
nor I_26488 (I453419,I453869,I453852);
not I_26489 (I453900,I453869);
nand I_26490 (I453422,I453629,I453900);
DFFARX1 I_26491 (I453869,I3563,I453445,I453434,);
DFFARX1 I_26492 (I453869,I3563,I453445,I453431,);
not I_26493 (I453989,I3570);
DFFARX1 I_26494 (I810430,I3563,I453989,I454015,);
DFFARX1 I_26495 (I454015,I3563,I453989,I454032,);
not I_26496 (I453981,I454032);
not I_26497 (I454054,I454015);
nand I_26498 (I454071,I810451,I810442);
and I_26499 (I454088,I454071,I810430);
DFFARX1 I_26500 (I454088,I3563,I453989,I454114,);
not I_26501 (I454122,I454114);
DFFARX1 I_26502 (I810436,I3563,I453989,I454148,);
and I_26503 (I454156,I454148,I810433);
nand I_26504 (I454173,I454148,I810433);
nand I_26505 (I453960,I454122,I454173);
DFFARX1 I_26506 (I810427,I3563,I453989,I454213,);
nor I_26507 (I454221,I454213,I454156);
DFFARX1 I_26508 (I454221,I3563,I453989,I453954,);
nor I_26509 (I453969,I454213,I454114);
nand I_26510 (I454266,I810427,I810439);
and I_26511 (I454283,I454266,I810448);
DFFARX1 I_26512 (I454283,I3563,I453989,I454309,);
nor I_26513 (I453957,I454309,I454213);
not I_26514 (I454331,I454309);
nor I_26515 (I454348,I454331,I454122);
nor I_26516 (I454365,I454054,I454348);
DFFARX1 I_26517 (I454365,I3563,I453989,I453972,);
nor I_26518 (I454396,I454331,I454213);
nor I_26519 (I454413,I810445,I810439);
nor I_26520 (I453963,I454413,I454396);
not I_26521 (I454444,I454413);
nand I_26522 (I453966,I454173,I454444);
DFFARX1 I_26523 (I454413,I3563,I453989,I453978,);
DFFARX1 I_26524 (I454413,I3563,I453989,I453975,);
not I_26525 (I454533,I3570);
DFFARX1 I_26526 (I834256,I3563,I454533,I454559,);
DFFARX1 I_26527 (I454559,I3563,I454533,I454576,);
not I_26528 (I454525,I454576);
not I_26529 (I454598,I454559);
nand I_26530 (I454615,I834250,I834247);
and I_26531 (I454632,I454615,I834262);
DFFARX1 I_26532 (I454632,I3563,I454533,I454658,);
not I_26533 (I454666,I454658);
DFFARX1 I_26534 (I834250,I3563,I454533,I454692,);
and I_26535 (I454700,I454692,I834244);
nand I_26536 (I454717,I454692,I834244);
nand I_26537 (I454504,I454666,I454717);
DFFARX1 I_26538 (I834244,I3563,I454533,I454757,);
nor I_26539 (I454765,I454757,I454700);
DFFARX1 I_26540 (I454765,I3563,I454533,I454498,);
nor I_26541 (I454513,I454757,I454658);
nand I_26542 (I454810,I834259,I834253);
and I_26543 (I454827,I454810,I834247);
DFFARX1 I_26544 (I454827,I3563,I454533,I454853,);
nor I_26545 (I454501,I454853,I454757);
not I_26546 (I454875,I454853);
nor I_26547 (I454892,I454875,I454666);
nor I_26548 (I454909,I454598,I454892);
DFFARX1 I_26549 (I454909,I3563,I454533,I454516,);
nor I_26550 (I454940,I454875,I454757);
nor I_26551 (I454957,I834265,I834253);
nor I_26552 (I454507,I454957,I454940);
not I_26553 (I454988,I454957);
nand I_26554 (I454510,I454717,I454988);
DFFARX1 I_26555 (I454957,I3563,I454533,I454522,);
DFFARX1 I_26556 (I454957,I3563,I454533,I454519,);
not I_26557 (I455077,I3570);
DFFARX1 I_26558 (I195257,I3563,I455077,I455103,);
DFFARX1 I_26559 (I455103,I3563,I455077,I455120,);
not I_26560 (I455069,I455120);
not I_26561 (I455142,I455103);
nand I_26562 (I455159,I195269,I195248);
and I_26563 (I455176,I455159,I195251);
DFFARX1 I_26564 (I455176,I3563,I455077,I455202,);
not I_26565 (I455210,I455202);
DFFARX1 I_26566 (I195260,I3563,I455077,I455236,);
and I_26567 (I455244,I455236,I195272);
nand I_26568 (I455261,I455236,I195272);
nand I_26569 (I455048,I455210,I455261);
DFFARX1 I_26570 (I195266,I3563,I455077,I455301,);
nor I_26571 (I455309,I455301,I455244);
DFFARX1 I_26572 (I455309,I3563,I455077,I455042,);
nor I_26573 (I455057,I455301,I455202);
nand I_26574 (I455354,I195254,I195251);
and I_26575 (I455371,I455354,I195263);
DFFARX1 I_26576 (I455371,I3563,I455077,I455397,);
nor I_26577 (I455045,I455397,I455301);
not I_26578 (I455419,I455397);
nor I_26579 (I455436,I455419,I455210);
nor I_26580 (I455453,I455142,I455436);
DFFARX1 I_26581 (I455453,I3563,I455077,I455060,);
nor I_26582 (I455484,I455419,I455301);
nor I_26583 (I455501,I195248,I195251);
nor I_26584 (I455051,I455501,I455484);
not I_26585 (I455532,I455501);
nand I_26586 (I455054,I455261,I455532);
DFFARX1 I_26587 (I455501,I3563,I455077,I455066,);
DFFARX1 I_26588 (I455501,I3563,I455077,I455063,);
not I_26589 (I455621,I3570);
DFFARX1 I_26590 (I1011135,I3563,I455621,I455647,);
DFFARX1 I_26591 (I455647,I3563,I455621,I455664,);
not I_26592 (I455613,I455664);
not I_26593 (I455686,I455647);
nand I_26594 (I455703,I1011150,I1011138);
and I_26595 (I455720,I455703,I1011129);
DFFARX1 I_26596 (I455720,I3563,I455621,I455746,);
not I_26597 (I455754,I455746);
DFFARX1 I_26598 (I1011141,I3563,I455621,I455780,);
and I_26599 (I455788,I455780,I1011132);
nand I_26600 (I455805,I455780,I1011132);
nand I_26601 (I455592,I455754,I455805);
DFFARX1 I_26602 (I1011147,I3563,I455621,I455845,);
nor I_26603 (I455853,I455845,I455788);
DFFARX1 I_26604 (I455853,I3563,I455621,I455586,);
nor I_26605 (I455601,I455845,I455746);
nand I_26606 (I455898,I1011156,I1011144);
and I_26607 (I455915,I455898,I1011153);
DFFARX1 I_26608 (I455915,I3563,I455621,I455941,);
nor I_26609 (I455589,I455941,I455845);
not I_26610 (I455963,I455941);
nor I_26611 (I455980,I455963,I455754);
nor I_26612 (I455997,I455686,I455980);
DFFARX1 I_26613 (I455997,I3563,I455621,I455604,);
nor I_26614 (I456028,I455963,I455845);
nor I_26615 (I456045,I1011129,I1011144);
nor I_26616 (I455595,I456045,I456028);
not I_26617 (I456076,I456045);
nand I_26618 (I455598,I455805,I456076);
DFFARX1 I_26619 (I456045,I3563,I455621,I455610,);
DFFARX1 I_26620 (I456045,I3563,I455621,I455607,);
not I_26621 (I456165,I3570);
DFFARX1 I_26622 (I41903,I3563,I456165,I456191,);
DFFARX1 I_26623 (I456191,I3563,I456165,I456208,);
not I_26624 (I456157,I456208);
not I_26625 (I456230,I456191);
nand I_26626 (I456247,I41891,I41906);
and I_26627 (I456264,I456247,I41894);
DFFARX1 I_26628 (I456264,I3563,I456165,I456290,);
not I_26629 (I456298,I456290);
DFFARX1 I_26630 (I41915,I3563,I456165,I456324,);
and I_26631 (I456332,I456324,I41909);
nand I_26632 (I456349,I456324,I41909);
nand I_26633 (I456136,I456298,I456349);
DFFARX1 I_26634 (I41912,I3563,I456165,I456389,);
nor I_26635 (I456397,I456389,I456332);
DFFARX1 I_26636 (I456397,I3563,I456165,I456130,);
nor I_26637 (I456145,I456389,I456290);
nand I_26638 (I456442,I41891,I41894);
and I_26639 (I456459,I456442,I41897);
DFFARX1 I_26640 (I456459,I3563,I456165,I456485,);
nor I_26641 (I456133,I456485,I456389);
not I_26642 (I456507,I456485);
nor I_26643 (I456524,I456507,I456298);
nor I_26644 (I456541,I456230,I456524);
DFFARX1 I_26645 (I456541,I3563,I456165,I456148,);
nor I_26646 (I456572,I456507,I456389);
nor I_26647 (I456589,I41900,I41894);
nor I_26648 (I456139,I456589,I456572);
not I_26649 (I456620,I456589);
nand I_26650 (I456142,I456349,I456620);
DFFARX1 I_26651 (I456589,I3563,I456165,I456154,);
DFFARX1 I_26652 (I456589,I3563,I456165,I456151,);
not I_26653 (I456709,I3570);
DFFARX1 I_26654 (I969145,I3563,I456709,I456735,);
DFFARX1 I_26655 (I456735,I3563,I456709,I456752,);
not I_26656 (I456701,I456752);
not I_26657 (I456774,I456735);
nand I_26658 (I456791,I969160,I969148);
and I_26659 (I456808,I456791,I969139);
DFFARX1 I_26660 (I456808,I3563,I456709,I456834,);
not I_26661 (I456842,I456834);
DFFARX1 I_26662 (I969151,I3563,I456709,I456868,);
and I_26663 (I456876,I456868,I969142);
nand I_26664 (I456893,I456868,I969142);
nand I_26665 (I456680,I456842,I456893);
DFFARX1 I_26666 (I969157,I3563,I456709,I456933,);
nor I_26667 (I456941,I456933,I456876);
DFFARX1 I_26668 (I456941,I3563,I456709,I456674,);
nor I_26669 (I456689,I456933,I456834);
nand I_26670 (I456986,I969166,I969154);
and I_26671 (I457003,I456986,I969163);
DFFARX1 I_26672 (I457003,I3563,I456709,I457029,);
nor I_26673 (I456677,I457029,I456933);
not I_26674 (I457051,I457029);
nor I_26675 (I457068,I457051,I456842);
nor I_26676 (I457085,I456774,I457068);
DFFARX1 I_26677 (I457085,I3563,I456709,I456692,);
nor I_26678 (I457116,I457051,I456933);
nor I_26679 (I457133,I969139,I969154);
nor I_26680 (I456683,I457133,I457116);
not I_26681 (I457164,I457133);
nand I_26682 (I456686,I456893,I457164);
DFFARX1 I_26683 (I457133,I3563,I456709,I456698,);
DFFARX1 I_26684 (I457133,I3563,I456709,I456695,);
not I_26685 (I457253,I3570);
DFFARX1 I_26686 (I982711,I3563,I457253,I457279,);
DFFARX1 I_26687 (I457279,I3563,I457253,I457296,);
not I_26688 (I457245,I457296);
not I_26689 (I457318,I457279);
nand I_26690 (I457335,I982726,I982714);
and I_26691 (I457352,I457335,I982705);
DFFARX1 I_26692 (I457352,I3563,I457253,I457378,);
not I_26693 (I457386,I457378);
DFFARX1 I_26694 (I982717,I3563,I457253,I457412,);
and I_26695 (I457420,I457412,I982708);
nand I_26696 (I457437,I457412,I982708);
nand I_26697 (I457224,I457386,I457437);
DFFARX1 I_26698 (I982723,I3563,I457253,I457477,);
nor I_26699 (I457485,I457477,I457420);
DFFARX1 I_26700 (I457485,I3563,I457253,I457218,);
nor I_26701 (I457233,I457477,I457378);
nand I_26702 (I457530,I982732,I982720);
and I_26703 (I457547,I457530,I982729);
DFFARX1 I_26704 (I457547,I3563,I457253,I457573,);
nor I_26705 (I457221,I457573,I457477);
not I_26706 (I457595,I457573);
nor I_26707 (I457612,I457595,I457386);
nor I_26708 (I457629,I457318,I457612);
DFFARX1 I_26709 (I457629,I3563,I457253,I457236,);
nor I_26710 (I457660,I457595,I457477);
nor I_26711 (I457677,I982705,I982720);
nor I_26712 (I457227,I457677,I457660);
not I_26713 (I457708,I457677);
nand I_26714 (I457230,I457437,I457708);
DFFARX1 I_26715 (I457677,I3563,I457253,I457242,);
DFFARX1 I_26716 (I457677,I3563,I457253,I457239,);
not I_26717 (I457797,I3570);
DFFARX1 I_26718 (I1022117,I3563,I457797,I457823,);
DFFARX1 I_26719 (I457823,I3563,I457797,I457840,);
not I_26720 (I457789,I457840);
not I_26721 (I457862,I457823);
nand I_26722 (I457879,I1022132,I1022120);
and I_26723 (I457896,I457879,I1022111);
DFFARX1 I_26724 (I457896,I3563,I457797,I457922,);
not I_26725 (I457930,I457922);
DFFARX1 I_26726 (I1022123,I3563,I457797,I457956,);
and I_26727 (I457964,I457956,I1022114);
nand I_26728 (I457981,I457956,I1022114);
nand I_26729 (I457768,I457930,I457981);
DFFARX1 I_26730 (I1022129,I3563,I457797,I458021,);
nor I_26731 (I458029,I458021,I457964);
DFFARX1 I_26732 (I458029,I3563,I457797,I457762,);
nor I_26733 (I457777,I458021,I457922);
nand I_26734 (I458074,I1022138,I1022126);
and I_26735 (I458091,I458074,I1022135);
DFFARX1 I_26736 (I458091,I3563,I457797,I458117,);
nor I_26737 (I457765,I458117,I458021);
not I_26738 (I458139,I458117);
nor I_26739 (I458156,I458139,I457930);
nor I_26740 (I458173,I457862,I458156);
DFFARX1 I_26741 (I458173,I3563,I457797,I457780,);
nor I_26742 (I458204,I458139,I458021);
nor I_26743 (I458221,I1022111,I1022126);
nor I_26744 (I457771,I458221,I458204);
not I_26745 (I458252,I458221);
nand I_26746 (I457774,I457981,I458252);
DFFARX1 I_26747 (I458221,I3563,I457797,I457786,);
DFFARX1 I_26748 (I458221,I3563,I457797,I457783,);
not I_26749 (I458341,I3570);
DFFARX1 I_26750 (I1153422,I3563,I458341,I458367,);
DFFARX1 I_26751 (I458367,I3563,I458341,I458384,);
not I_26752 (I458333,I458384);
not I_26753 (I458406,I458367);
nand I_26754 (I458423,I1153434,I1153422);
and I_26755 (I458440,I458423,I1153425);
DFFARX1 I_26756 (I458440,I3563,I458341,I458466,);
not I_26757 (I458474,I458466);
DFFARX1 I_26758 (I1153443,I3563,I458341,I458500,);
and I_26759 (I458508,I458500,I1153419);
nand I_26760 (I458525,I458500,I1153419);
nand I_26761 (I458312,I458474,I458525);
DFFARX1 I_26762 (I1153437,I3563,I458341,I458565,);
nor I_26763 (I458573,I458565,I458508);
DFFARX1 I_26764 (I458573,I3563,I458341,I458306,);
nor I_26765 (I458321,I458565,I458466);
nand I_26766 (I458618,I1153431,I1153428);
and I_26767 (I458635,I458618,I1153440);
DFFARX1 I_26768 (I458635,I3563,I458341,I458661,);
nor I_26769 (I458309,I458661,I458565);
not I_26770 (I458683,I458661);
nor I_26771 (I458700,I458683,I458474);
nor I_26772 (I458717,I458406,I458700);
DFFARX1 I_26773 (I458717,I3563,I458341,I458324,);
nor I_26774 (I458748,I458683,I458565);
nor I_26775 (I458765,I1153419,I1153428);
nor I_26776 (I458315,I458765,I458748);
not I_26777 (I458796,I458765);
nand I_26778 (I458318,I458525,I458796);
DFFARX1 I_26779 (I458765,I3563,I458341,I458330,);
DFFARX1 I_26780 (I458765,I3563,I458341,I458327,);
not I_26781 (I458885,I3570);
DFFARX1 I_26782 (I304358,I3563,I458885,I458911,);
DFFARX1 I_26783 (I458911,I3563,I458885,I458928,);
not I_26784 (I458877,I458928);
not I_26785 (I458950,I458911);
nand I_26786 (I458967,I304337,I304361);
and I_26787 (I458984,I458967,I304364);
DFFARX1 I_26788 (I458984,I3563,I458885,I459010,);
not I_26789 (I459018,I459010);
DFFARX1 I_26790 (I304346,I3563,I458885,I459044,);
and I_26791 (I459052,I459044,I304352);
nand I_26792 (I459069,I459044,I304352);
nand I_26793 (I458856,I459018,I459069);
DFFARX1 I_26794 (I304340,I3563,I458885,I459109,);
nor I_26795 (I459117,I459109,I459052);
DFFARX1 I_26796 (I459117,I3563,I458885,I458850,);
nor I_26797 (I458865,I459109,I459010);
nand I_26798 (I459162,I304349,I304337);
and I_26799 (I459179,I459162,I304343);
DFFARX1 I_26800 (I459179,I3563,I458885,I459205,);
nor I_26801 (I458853,I459205,I459109);
not I_26802 (I459227,I459205);
nor I_26803 (I459244,I459227,I459018);
nor I_26804 (I459261,I458950,I459244);
DFFARX1 I_26805 (I459261,I3563,I458885,I458868,);
nor I_26806 (I459292,I459227,I459109);
nor I_26807 (I459309,I304355,I304337);
nor I_26808 (I458859,I459309,I459292);
not I_26809 (I459340,I459309);
nand I_26810 (I458862,I459069,I459340);
DFFARX1 I_26811 (I459309,I3563,I458885,I458874,);
DFFARX1 I_26812 (I459309,I3563,I458885,I458871,);
not I_26813 (I459429,I3570);
DFFARX1 I_26814 (I1397005,I3563,I459429,I459455,);
DFFARX1 I_26815 (I459455,I3563,I459429,I459472,);
not I_26816 (I459421,I459472);
not I_26817 (I459494,I459455);
nand I_26818 (I459511,I1396981,I1397002);
and I_26819 (I459528,I459511,I1396999);
DFFARX1 I_26820 (I459528,I3563,I459429,I459554,);
not I_26821 (I459562,I459554);
DFFARX1 I_26822 (I1396978,I3563,I459429,I459588,);
and I_26823 (I459596,I459588,I1396990);
nand I_26824 (I459613,I459588,I1396990);
nand I_26825 (I459400,I459562,I459613);
DFFARX1 I_26826 (I1396993,I3563,I459429,I459653,);
nor I_26827 (I459661,I459653,I459596);
DFFARX1 I_26828 (I459661,I3563,I459429,I459394,);
nor I_26829 (I459409,I459653,I459554);
nand I_26830 (I459706,I1396996,I1396984);
and I_26831 (I459723,I459706,I1396987);
DFFARX1 I_26832 (I459723,I3563,I459429,I459749,);
nor I_26833 (I459397,I459749,I459653);
not I_26834 (I459771,I459749);
nor I_26835 (I459788,I459771,I459562);
nor I_26836 (I459805,I459494,I459788);
DFFARX1 I_26837 (I459805,I3563,I459429,I459412,);
nor I_26838 (I459836,I459771,I459653);
nor I_26839 (I459853,I1396978,I1396984);
nor I_26840 (I459403,I459853,I459836);
not I_26841 (I459884,I459853);
nand I_26842 (I459406,I459613,I459884);
DFFARX1 I_26843 (I459853,I3563,I459429,I459418,);
DFFARX1 I_26844 (I459853,I3563,I459429,I459415,);
not I_26845 (I459973,I3570);
DFFARX1 I_26846 (I845323,I3563,I459973,I459999,);
DFFARX1 I_26847 (I459999,I3563,I459973,I460016,);
not I_26848 (I459965,I460016);
not I_26849 (I460038,I459999);
nand I_26850 (I460055,I845317,I845314);
and I_26851 (I460072,I460055,I845329);
DFFARX1 I_26852 (I460072,I3563,I459973,I460098,);
not I_26853 (I460106,I460098);
DFFARX1 I_26854 (I845317,I3563,I459973,I460132,);
and I_26855 (I460140,I460132,I845311);
nand I_26856 (I460157,I460132,I845311);
nand I_26857 (I459944,I460106,I460157);
DFFARX1 I_26858 (I845311,I3563,I459973,I460197,);
nor I_26859 (I460205,I460197,I460140);
DFFARX1 I_26860 (I460205,I3563,I459973,I459938,);
nor I_26861 (I459953,I460197,I460098);
nand I_26862 (I460250,I845326,I845320);
and I_26863 (I460267,I460250,I845314);
DFFARX1 I_26864 (I460267,I3563,I459973,I460293,);
nor I_26865 (I459941,I460293,I460197);
not I_26866 (I460315,I460293);
nor I_26867 (I460332,I460315,I460106);
nor I_26868 (I460349,I460038,I460332);
DFFARX1 I_26869 (I460349,I3563,I459973,I459956,);
nor I_26870 (I460380,I460315,I460197);
nor I_26871 (I460397,I845332,I845320);
nor I_26872 (I459947,I460397,I460380);
not I_26873 (I460428,I460397);
nand I_26874 (I459950,I460157,I460428);
DFFARX1 I_26875 (I460397,I3563,I459973,I459962,);
DFFARX1 I_26876 (I460397,I3563,I459973,I459959,);
not I_26877 (I460517,I3570);
DFFARX1 I_26878 (I1079197,I3563,I460517,I460543,);
DFFARX1 I_26879 (I460543,I3563,I460517,I460560,);
not I_26880 (I460509,I460560);
not I_26881 (I460582,I460543);
nand I_26882 (I460599,I1079197,I1079215);
and I_26883 (I460616,I460599,I1079209);
DFFARX1 I_26884 (I460616,I3563,I460517,I460642,);
not I_26885 (I460650,I460642);
DFFARX1 I_26886 (I1079203,I3563,I460517,I460676,);
and I_26887 (I460684,I460676,I1079212);
nand I_26888 (I460701,I460676,I1079212);
nand I_26889 (I460488,I460650,I460701);
DFFARX1 I_26890 (I1079200,I3563,I460517,I460741,);
nor I_26891 (I460749,I460741,I460684);
DFFARX1 I_26892 (I460749,I3563,I460517,I460482,);
nor I_26893 (I460497,I460741,I460642);
nand I_26894 (I460794,I1079200,I1079218);
and I_26895 (I460811,I460794,I1079203);
DFFARX1 I_26896 (I460811,I3563,I460517,I460837,);
nor I_26897 (I460485,I460837,I460741);
not I_26898 (I460859,I460837);
nor I_26899 (I460876,I460859,I460650);
nor I_26900 (I460893,I460582,I460876);
DFFARX1 I_26901 (I460893,I3563,I460517,I460500,);
nor I_26902 (I460924,I460859,I460741);
nor I_26903 (I460941,I1079206,I1079218);
nor I_26904 (I460491,I460941,I460924);
not I_26905 (I460972,I460941);
nand I_26906 (I460494,I460701,I460972);
DFFARX1 I_26907 (I460941,I3563,I460517,I460506,);
DFFARX1 I_26908 (I460941,I3563,I460517,I460503,);
not I_26909 (I461061,I3570);
DFFARX1 I_26910 (I819500,I3563,I461061,I461087,);
DFFARX1 I_26911 (I461087,I3563,I461061,I461104,);
not I_26912 (I461053,I461104);
not I_26913 (I461126,I461087);
nand I_26914 (I461143,I819494,I819491);
and I_26915 (I461160,I461143,I819506);
DFFARX1 I_26916 (I461160,I3563,I461061,I461186,);
not I_26917 (I461194,I461186);
DFFARX1 I_26918 (I819494,I3563,I461061,I461220,);
and I_26919 (I461228,I461220,I819488);
nand I_26920 (I461245,I461220,I819488);
nand I_26921 (I461032,I461194,I461245);
DFFARX1 I_26922 (I819488,I3563,I461061,I461285,);
nor I_26923 (I461293,I461285,I461228);
DFFARX1 I_26924 (I461293,I3563,I461061,I461026,);
nor I_26925 (I461041,I461285,I461186);
nand I_26926 (I461338,I819503,I819497);
and I_26927 (I461355,I461338,I819491);
DFFARX1 I_26928 (I461355,I3563,I461061,I461381,);
nor I_26929 (I461029,I461381,I461285);
not I_26930 (I461403,I461381);
nor I_26931 (I461420,I461403,I461194);
nor I_26932 (I461437,I461126,I461420);
DFFARX1 I_26933 (I461437,I3563,I461061,I461044,);
nor I_26934 (I461468,I461403,I461285);
nor I_26935 (I461485,I819509,I819497);
nor I_26936 (I461035,I461485,I461468);
not I_26937 (I461516,I461485);
nand I_26938 (I461038,I461245,I461516);
DFFARX1 I_26939 (I461485,I3563,I461061,I461050,);
DFFARX1 I_26940 (I461485,I3563,I461061,I461047,);
not I_26941 (I461605,I3570);
DFFARX1 I_26942 (I856390,I3563,I461605,I461631,);
DFFARX1 I_26943 (I461631,I3563,I461605,I461648,);
not I_26944 (I461597,I461648);
not I_26945 (I461670,I461631);
nand I_26946 (I461687,I856384,I856381);
and I_26947 (I461704,I461687,I856396);
DFFARX1 I_26948 (I461704,I3563,I461605,I461730,);
not I_26949 (I461738,I461730);
DFFARX1 I_26950 (I856384,I3563,I461605,I461764,);
and I_26951 (I461772,I461764,I856378);
nand I_26952 (I461789,I461764,I856378);
nand I_26953 (I461576,I461738,I461789);
DFFARX1 I_26954 (I856378,I3563,I461605,I461829,);
nor I_26955 (I461837,I461829,I461772);
DFFARX1 I_26956 (I461837,I3563,I461605,I461570,);
nor I_26957 (I461585,I461829,I461730);
nand I_26958 (I461882,I856393,I856387);
and I_26959 (I461899,I461882,I856381);
DFFARX1 I_26960 (I461899,I3563,I461605,I461925,);
nor I_26961 (I461573,I461925,I461829);
not I_26962 (I461947,I461925);
nor I_26963 (I461964,I461947,I461738);
nor I_26964 (I461981,I461670,I461964);
DFFARX1 I_26965 (I461981,I3563,I461605,I461588,);
nor I_26966 (I462012,I461947,I461829);
nor I_26967 (I462029,I856399,I856387);
nor I_26968 (I461579,I462029,I462012);
not I_26969 (I462060,I462029);
nand I_26970 (I461582,I461789,I462060);
DFFARX1 I_26971 (I462029,I3563,I461605,I461594,);
DFFARX1 I_26972 (I462029,I3563,I461605,I461591,);
not I_26973 (I462149,I3570);
DFFARX1 I_26974 (I1128568,I3563,I462149,I462175,);
DFFARX1 I_26975 (I462175,I3563,I462149,I462192,);
not I_26976 (I462141,I462192);
not I_26977 (I462214,I462175);
nand I_26978 (I462231,I1128580,I1128568);
and I_26979 (I462248,I462231,I1128571);
DFFARX1 I_26980 (I462248,I3563,I462149,I462274,);
not I_26981 (I462282,I462274);
DFFARX1 I_26982 (I1128589,I3563,I462149,I462308,);
and I_26983 (I462316,I462308,I1128565);
nand I_26984 (I462333,I462308,I1128565);
nand I_26985 (I462120,I462282,I462333);
DFFARX1 I_26986 (I1128583,I3563,I462149,I462373,);
nor I_26987 (I462381,I462373,I462316);
DFFARX1 I_26988 (I462381,I3563,I462149,I462114,);
nor I_26989 (I462129,I462373,I462274);
nand I_26990 (I462426,I1128577,I1128574);
and I_26991 (I462443,I462426,I1128586);
DFFARX1 I_26992 (I462443,I3563,I462149,I462469,);
nor I_26993 (I462117,I462469,I462373);
not I_26994 (I462491,I462469);
nor I_26995 (I462508,I462491,I462282);
nor I_26996 (I462525,I462214,I462508);
DFFARX1 I_26997 (I462525,I3563,I462149,I462132,);
nor I_26998 (I462556,I462491,I462373);
nor I_26999 (I462573,I1128565,I1128574);
nor I_27000 (I462123,I462573,I462556);
not I_27001 (I462604,I462573);
nand I_27002 (I462126,I462333,I462604);
DFFARX1 I_27003 (I462573,I3563,I462149,I462138,);
DFFARX1 I_27004 (I462573,I3563,I462149,I462135,);
not I_27005 (I462693,I3570);
DFFARX1 I_27006 (I1260556,I3563,I462693,I462719,);
DFFARX1 I_27007 (I462719,I3563,I462693,I462736,);
not I_27008 (I462685,I462736);
not I_27009 (I462758,I462719);
nand I_27010 (I462775,I1260568,I1260571);
and I_27011 (I462792,I462775,I1260574);
DFFARX1 I_27012 (I462792,I3563,I462693,I462818,);
not I_27013 (I462826,I462818);
DFFARX1 I_27014 (I1260559,I3563,I462693,I462852,);
and I_27015 (I462860,I462852,I1260565);
nand I_27016 (I462877,I462852,I1260565);
nand I_27017 (I462664,I462826,I462877);
DFFARX1 I_27018 (I1260553,I3563,I462693,I462917,);
nor I_27019 (I462925,I462917,I462860);
DFFARX1 I_27020 (I462925,I3563,I462693,I462658,);
nor I_27021 (I462673,I462917,I462818);
nand I_27022 (I462970,I1260556,I1260577);
and I_27023 (I462987,I462970,I1260562);
DFFARX1 I_27024 (I462987,I3563,I462693,I463013,);
nor I_27025 (I462661,I463013,I462917);
not I_27026 (I463035,I463013);
nor I_27027 (I463052,I463035,I462826);
nor I_27028 (I463069,I462758,I463052);
DFFARX1 I_27029 (I463069,I3563,I462693,I462676,);
nor I_27030 (I463100,I463035,I462917);
nor I_27031 (I463117,I1260553,I1260577);
nor I_27032 (I462667,I463117,I463100);
not I_27033 (I463148,I463117);
nand I_27034 (I462670,I462877,I463148);
DFFARX1 I_27035 (I463117,I3563,I462693,I462682,);
DFFARX1 I_27036 (I463117,I3563,I462693,I462679,);
not I_27037 (I463237,I3570);
DFFARX1 I_27038 (I1377370,I3563,I463237,I463263,);
DFFARX1 I_27039 (I463263,I3563,I463237,I463280,);
not I_27040 (I463229,I463280);
not I_27041 (I463302,I463263);
nand I_27042 (I463319,I1377346,I1377367);
and I_27043 (I463336,I463319,I1377364);
DFFARX1 I_27044 (I463336,I3563,I463237,I463362,);
not I_27045 (I463370,I463362);
DFFARX1 I_27046 (I1377343,I3563,I463237,I463396,);
and I_27047 (I463404,I463396,I1377355);
nand I_27048 (I463421,I463396,I1377355);
nand I_27049 (I463208,I463370,I463421);
DFFARX1 I_27050 (I1377358,I3563,I463237,I463461,);
nor I_27051 (I463469,I463461,I463404);
DFFARX1 I_27052 (I463469,I3563,I463237,I463202,);
nor I_27053 (I463217,I463461,I463362);
nand I_27054 (I463514,I1377361,I1377349);
and I_27055 (I463531,I463514,I1377352);
DFFARX1 I_27056 (I463531,I3563,I463237,I463557,);
nor I_27057 (I463205,I463557,I463461);
not I_27058 (I463579,I463557);
nor I_27059 (I463596,I463579,I463370);
nor I_27060 (I463613,I463302,I463596);
DFFARX1 I_27061 (I463613,I3563,I463237,I463220,);
nor I_27062 (I463644,I463579,I463461);
nor I_27063 (I463661,I1377343,I1377349);
nor I_27064 (I463211,I463661,I463644);
not I_27065 (I463692,I463661);
nand I_27066 (I463214,I463421,I463692);
DFFARX1 I_27067 (I463661,I3563,I463237,I463226,);
DFFARX1 I_27068 (I463661,I3563,I463237,I463223,);
not I_27069 (I463781,I3570);
DFFARX1 I_27070 (I1374990,I3563,I463781,I463807,);
DFFARX1 I_27071 (I463807,I3563,I463781,I463824,);
not I_27072 (I463773,I463824);
not I_27073 (I463846,I463807);
nand I_27074 (I463863,I1374966,I1374987);
and I_27075 (I463880,I463863,I1374984);
DFFARX1 I_27076 (I463880,I3563,I463781,I463906,);
not I_27077 (I463914,I463906);
DFFARX1 I_27078 (I1374963,I3563,I463781,I463940,);
and I_27079 (I463948,I463940,I1374975);
nand I_27080 (I463965,I463940,I1374975);
nand I_27081 (I463752,I463914,I463965);
DFFARX1 I_27082 (I1374978,I3563,I463781,I464005,);
nor I_27083 (I464013,I464005,I463948);
DFFARX1 I_27084 (I464013,I3563,I463781,I463746,);
nor I_27085 (I463761,I464005,I463906);
nand I_27086 (I464058,I1374981,I1374969);
and I_27087 (I464075,I464058,I1374972);
DFFARX1 I_27088 (I464075,I3563,I463781,I464101,);
nor I_27089 (I463749,I464101,I464005);
not I_27090 (I464123,I464101);
nor I_27091 (I464140,I464123,I463914);
nor I_27092 (I464157,I463846,I464140);
DFFARX1 I_27093 (I464157,I3563,I463781,I463764,);
nor I_27094 (I464188,I464123,I464005);
nor I_27095 (I464205,I1374963,I1374969);
nor I_27096 (I463755,I464205,I464188);
not I_27097 (I464236,I464205);
nand I_27098 (I463758,I463965,I464236);
DFFARX1 I_27099 (I464205,I3563,I463781,I463770,);
DFFARX1 I_27100 (I464205,I3563,I463781,I463767,);
not I_27101 (I464325,I3570);
DFFARX1 I_27102 (I1307423,I3563,I464325,I464351,);
DFFARX1 I_27103 (I464351,I3563,I464325,I464368,);
not I_27104 (I464317,I464368);
not I_27105 (I464390,I464351);
nand I_27106 (I464407,I1307420,I1307417);
and I_27107 (I464424,I464407,I1307405);
DFFARX1 I_27108 (I464424,I3563,I464325,I464450,);
not I_27109 (I464458,I464450);
DFFARX1 I_27110 (I1307429,I3563,I464325,I464484,);
and I_27111 (I464492,I464484,I1307414);
nand I_27112 (I464509,I464484,I1307414);
nand I_27113 (I464296,I464458,I464509);
DFFARX1 I_27114 (I1307408,I3563,I464325,I464549,);
nor I_27115 (I464557,I464549,I464492);
DFFARX1 I_27116 (I464557,I3563,I464325,I464290,);
nor I_27117 (I464305,I464549,I464450);
nand I_27118 (I464602,I1307405,I1307411);
and I_27119 (I464619,I464602,I1307426);
DFFARX1 I_27120 (I464619,I3563,I464325,I464645,);
nor I_27121 (I464293,I464645,I464549);
not I_27122 (I464667,I464645);
nor I_27123 (I464684,I464667,I464458);
nor I_27124 (I464701,I464390,I464684);
DFFARX1 I_27125 (I464701,I3563,I464325,I464308,);
nor I_27126 (I464732,I464667,I464549);
nor I_27127 (I464749,I1307408,I1307411);
nor I_27128 (I464299,I464749,I464732);
not I_27129 (I464780,I464749);
nand I_27130 (I464302,I464509,I464780);
DFFARX1 I_27131 (I464749,I3563,I464325,I464314,);
DFFARX1 I_27132 (I464749,I3563,I464325,I464311,);
not I_27133 (I464869,I3570);
DFFARX1 I_27134 (I298561,I3563,I464869,I464895,);
DFFARX1 I_27135 (I464895,I3563,I464869,I464912,);
not I_27136 (I464861,I464912);
not I_27137 (I464934,I464895);
nand I_27138 (I464951,I298540,I298564);
and I_27139 (I464968,I464951,I298567);
DFFARX1 I_27140 (I464968,I3563,I464869,I464994,);
not I_27141 (I465002,I464994);
DFFARX1 I_27142 (I298549,I3563,I464869,I465028,);
and I_27143 (I465036,I465028,I298555);
nand I_27144 (I465053,I465028,I298555);
nand I_27145 (I464840,I465002,I465053);
DFFARX1 I_27146 (I298543,I3563,I464869,I465093,);
nor I_27147 (I465101,I465093,I465036);
DFFARX1 I_27148 (I465101,I3563,I464869,I464834,);
nor I_27149 (I464849,I465093,I464994);
nand I_27150 (I465146,I298552,I298540);
and I_27151 (I465163,I465146,I298546);
DFFARX1 I_27152 (I465163,I3563,I464869,I465189,);
nor I_27153 (I464837,I465189,I465093);
not I_27154 (I465211,I465189);
nor I_27155 (I465228,I465211,I465002);
nor I_27156 (I465245,I464934,I465228);
DFFARX1 I_27157 (I465245,I3563,I464869,I464852,);
nor I_27158 (I465276,I465211,I465093);
nor I_27159 (I465293,I298558,I298540);
nor I_27160 (I464843,I465293,I465276);
not I_27161 (I465324,I465293);
nand I_27162 (I464846,I465053,I465324);
DFFARX1 I_27163 (I465293,I3563,I464869,I464858,);
DFFARX1 I_27164 (I465293,I3563,I464869,I464855,);
not I_27165 (I465413,I3570);
DFFARX1 I_27166 (I1036975,I3563,I465413,I465439,);
DFFARX1 I_27167 (I465439,I3563,I465413,I465456,);
not I_27168 (I465405,I465456);
not I_27169 (I465478,I465439);
nand I_27170 (I465495,I1036990,I1036978);
and I_27171 (I465512,I465495,I1036969);
DFFARX1 I_27172 (I465512,I3563,I465413,I465538,);
not I_27173 (I465546,I465538);
DFFARX1 I_27174 (I1036981,I3563,I465413,I465572,);
and I_27175 (I465580,I465572,I1036972);
nand I_27176 (I465597,I465572,I1036972);
nand I_27177 (I465384,I465546,I465597);
DFFARX1 I_27178 (I1036987,I3563,I465413,I465637,);
nor I_27179 (I465645,I465637,I465580);
DFFARX1 I_27180 (I465645,I3563,I465413,I465378,);
nor I_27181 (I465393,I465637,I465538);
nand I_27182 (I465690,I1036996,I1036984);
and I_27183 (I465707,I465690,I1036993);
DFFARX1 I_27184 (I465707,I3563,I465413,I465733,);
nor I_27185 (I465381,I465733,I465637);
not I_27186 (I465755,I465733);
nor I_27187 (I465772,I465755,I465546);
nor I_27188 (I465789,I465478,I465772);
DFFARX1 I_27189 (I465789,I3563,I465413,I465396,);
nor I_27190 (I465820,I465755,I465637);
nor I_27191 (I465837,I1036969,I1036984);
nor I_27192 (I465387,I465837,I465820);
not I_27193 (I465868,I465837);
nand I_27194 (I465390,I465597,I465868);
DFFARX1 I_27195 (I465837,I3563,I465413,I465402,);
DFFARX1 I_27196 (I465837,I3563,I465413,I465399,);
not I_27197 (I465957,I3570);
DFFARX1 I_27198 (I962685,I3563,I465957,I465983,);
DFFARX1 I_27199 (I465983,I3563,I465957,I466000,);
not I_27200 (I465949,I466000);
not I_27201 (I466022,I465983);
nand I_27202 (I466039,I962700,I962688);
and I_27203 (I466056,I466039,I962679);
DFFARX1 I_27204 (I466056,I3563,I465957,I466082,);
not I_27205 (I466090,I466082);
DFFARX1 I_27206 (I962691,I3563,I465957,I466116,);
and I_27207 (I466124,I466116,I962682);
nand I_27208 (I466141,I466116,I962682);
nand I_27209 (I465928,I466090,I466141);
DFFARX1 I_27210 (I962697,I3563,I465957,I466181,);
nor I_27211 (I466189,I466181,I466124);
DFFARX1 I_27212 (I466189,I3563,I465957,I465922,);
nor I_27213 (I465937,I466181,I466082);
nand I_27214 (I466234,I962706,I962694);
and I_27215 (I466251,I466234,I962703);
DFFARX1 I_27216 (I466251,I3563,I465957,I466277,);
nor I_27217 (I465925,I466277,I466181);
not I_27218 (I466299,I466277);
nor I_27219 (I466316,I466299,I466090);
nor I_27220 (I466333,I466022,I466316);
DFFARX1 I_27221 (I466333,I3563,I465957,I465940,);
nor I_27222 (I466364,I466299,I466181);
nor I_27223 (I466381,I962679,I962694);
nor I_27224 (I465931,I466381,I466364);
not I_27225 (I466412,I466381);
nand I_27226 (I465934,I466141,I466412);
DFFARX1 I_27227 (I466381,I3563,I465957,I465946,);
DFFARX1 I_27228 (I466381,I3563,I465957,I465943,);
not I_27229 (I466501,I3570);
DFFARX1 I_27230 (I643388,I3563,I466501,I466527,);
DFFARX1 I_27231 (I466527,I3563,I466501,I466544,);
not I_27232 (I466493,I466544);
not I_27233 (I466566,I466527);
nand I_27234 (I466583,I643385,I643406);
and I_27235 (I466600,I466583,I643409);
DFFARX1 I_27236 (I466600,I3563,I466501,I466626,);
not I_27237 (I466634,I466626);
DFFARX1 I_27238 (I643394,I3563,I466501,I466660,);
and I_27239 (I466668,I466660,I643397);
nand I_27240 (I466685,I466660,I643397);
nand I_27241 (I466472,I466634,I466685);
DFFARX1 I_27242 (I643400,I3563,I466501,I466725,);
nor I_27243 (I466733,I466725,I466668);
DFFARX1 I_27244 (I466733,I3563,I466501,I466466,);
nor I_27245 (I466481,I466725,I466626);
nand I_27246 (I466778,I643385,I643391);
and I_27247 (I466795,I466778,I643403);
DFFARX1 I_27248 (I466795,I3563,I466501,I466821,);
nor I_27249 (I466469,I466821,I466725);
not I_27250 (I466843,I466821);
nor I_27251 (I466860,I466843,I466634);
nor I_27252 (I466877,I466566,I466860);
DFFARX1 I_27253 (I466877,I3563,I466501,I466484,);
nor I_27254 (I466908,I466843,I466725);
nor I_27255 (I466925,I643388,I643391);
nor I_27256 (I466475,I466925,I466908);
not I_27257 (I466956,I466925);
nand I_27258 (I466478,I466685,I466956);
DFFARX1 I_27259 (I466925,I3563,I466501,I466490,);
DFFARX1 I_27260 (I466925,I3563,I466501,I466487,);
not I_27261 (I467045,I3570);
DFFARX1 I_27262 (I391840,I3563,I467045,I467071,);
DFFARX1 I_27263 (I467071,I3563,I467045,I467088,);
not I_27264 (I467037,I467088);
not I_27265 (I467110,I467071);
nand I_27266 (I467127,I391819,I391843);
and I_27267 (I467144,I467127,I391846);
DFFARX1 I_27268 (I467144,I3563,I467045,I467170,);
not I_27269 (I467178,I467170);
DFFARX1 I_27270 (I391828,I3563,I467045,I467204,);
and I_27271 (I467212,I467204,I391834);
nand I_27272 (I467229,I467204,I391834);
nand I_27273 (I467016,I467178,I467229);
DFFARX1 I_27274 (I391822,I3563,I467045,I467269,);
nor I_27275 (I467277,I467269,I467212);
DFFARX1 I_27276 (I467277,I3563,I467045,I467010,);
nor I_27277 (I467025,I467269,I467170);
nand I_27278 (I467322,I391831,I391819);
and I_27279 (I467339,I467322,I391825);
DFFARX1 I_27280 (I467339,I3563,I467045,I467365,);
nor I_27281 (I467013,I467365,I467269);
not I_27282 (I467387,I467365);
nor I_27283 (I467404,I467387,I467178);
nor I_27284 (I467421,I467110,I467404);
DFFARX1 I_27285 (I467421,I3563,I467045,I467028,);
nor I_27286 (I467452,I467387,I467269);
nor I_27287 (I467469,I391837,I391819);
nor I_27288 (I467019,I467469,I467452);
not I_27289 (I467500,I467469);
nand I_27290 (I467022,I467229,I467500);
DFFARX1 I_27291 (I467469,I3563,I467045,I467034,);
DFFARX1 I_27292 (I467469,I3563,I467045,I467031,);
not I_27293 (I467589,I3570);
DFFARX1 I_27294 (I248807,I3563,I467589,I467615,);
DFFARX1 I_27295 (I467615,I3563,I467589,I467632,);
not I_27296 (I467581,I467632);
not I_27297 (I467654,I467615);
nand I_27298 (I467671,I248819,I248798);
and I_27299 (I467688,I467671,I248801);
DFFARX1 I_27300 (I467688,I3563,I467589,I467714,);
not I_27301 (I467722,I467714);
DFFARX1 I_27302 (I248810,I3563,I467589,I467748,);
and I_27303 (I467756,I467748,I248822);
nand I_27304 (I467773,I467748,I248822);
nand I_27305 (I467560,I467722,I467773);
DFFARX1 I_27306 (I248816,I3563,I467589,I467813,);
nor I_27307 (I467821,I467813,I467756);
DFFARX1 I_27308 (I467821,I3563,I467589,I467554,);
nor I_27309 (I467569,I467813,I467714);
nand I_27310 (I467866,I248804,I248801);
and I_27311 (I467883,I467866,I248813);
DFFARX1 I_27312 (I467883,I3563,I467589,I467909,);
nor I_27313 (I467557,I467909,I467813);
not I_27314 (I467931,I467909);
nor I_27315 (I467948,I467931,I467722);
nor I_27316 (I467965,I467654,I467948);
DFFARX1 I_27317 (I467965,I3563,I467589,I467572,);
nor I_27318 (I467996,I467931,I467813);
nor I_27319 (I468013,I248798,I248801);
nor I_27320 (I467563,I468013,I467996);
not I_27321 (I468044,I468013);
nand I_27322 (I467566,I467773,I468044);
DFFARX1 I_27323 (I468013,I3563,I467589,I467578,);
DFFARX1 I_27324 (I468013,I3563,I467589,I467575,);
not I_27325 (I468133,I3570);
DFFARX1 I_27326 (I1311469,I3563,I468133,I468159,);
DFFARX1 I_27327 (I468159,I3563,I468133,I468176,);
not I_27328 (I468125,I468176);
not I_27329 (I468198,I468159);
nand I_27330 (I468215,I1311466,I1311463);
and I_27331 (I468232,I468215,I1311451);
DFFARX1 I_27332 (I468232,I3563,I468133,I468258,);
not I_27333 (I468266,I468258);
DFFARX1 I_27334 (I1311475,I3563,I468133,I468292,);
and I_27335 (I468300,I468292,I1311460);
nand I_27336 (I468317,I468292,I1311460);
nand I_27337 (I468104,I468266,I468317);
DFFARX1 I_27338 (I1311454,I3563,I468133,I468357,);
nor I_27339 (I468365,I468357,I468300);
DFFARX1 I_27340 (I468365,I3563,I468133,I468098,);
nor I_27341 (I468113,I468357,I468258);
nand I_27342 (I468410,I1311451,I1311457);
and I_27343 (I468427,I468410,I1311472);
DFFARX1 I_27344 (I468427,I3563,I468133,I468453,);
nor I_27345 (I468101,I468453,I468357);
not I_27346 (I468475,I468453);
nor I_27347 (I468492,I468475,I468266);
nor I_27348 (I468509,I468198,I468492);
DFFARX1 I_27349 (I468509,I3563,I468133,I468116,);
nor I_27350 (I468540,I468475,I468357);
nor I_27351 (I468557,I1311454,I1311457);
nor I_27352 (I468107,I468557,I468540);
not I_27353 (I468588,I468557);
nand I_27354 (I468110,I468317,I468588);
DFFARX1 I_27355 (I468557,I3563,I468133,I468122,);
DFFARX1 I_27356 (I468557,I3563,I468133,I468119,);
not I_27357 (I468677,I3570);
DFFARX1 I_27358 (I409231,I3563,I468677,I468703,);
DFFARX1 I_27359 (I468703,I3563,I468677,I468720,);
not I_27360 (I468669,I468720);
not I_27361 (I468742,I468703);
nand I_27362 (I468759,I409210,I409234);
and I_27363 (I468776,I468759,I409237);
DFFARX1 I_27364 (I468776,I3563,I468677,I468802,);
not I_27365 (I468810,I468802);
DFFARX1 I_27366 (I409219,I3563,I468677,I468836,);
and I_27367 (I468844,I468836,I409225);
nand I_27368 (I468861,I468836,I409225);
nand I_27369 (I468648,I468810,I468861);
DFFARX1 I_27370 (I409213,I3563,I468677,I468901,);
nor I_27371 (I468909,I468901,I468844);
DFFARX1 I_27372 (I468909,I3563,I468677,I468642,);
nor I_27373 (I468657,I468901,I468802);
nand I_27374 (I468954,I409222,I409210);
and I_27375 (I468971,I468954,I409216);
DFFARX1 I_27376 (I468971,I3563,I468677,I468997,);
nor I_27377 (I468645,I468997,I468901);
not I_27378 (I469019,I468997);
nor I_27379 (I469036,I469019,I468810);
nor I_27380 (I469053,I468742,I469036);
DFFARX1 I_27381 (I469053,I3563,I468677,I468660,);
nor I_27382 (I469084,I469019,I468901);
nor I_27383 (I469101,I409228,I409210);
nor I_27384 (I468651,I469101,I469084);
not I_27385 (I469132,I469101);
nand I_27386 (I468654,I468861,I469132);
DFFARX1 I_27387 (I469101,I3563,I468677,I468666,);
DFFARX1 I_27388 (I469101,I3563,I468677,I468663,);
not I_27389 (I469221,I3570);
DFFARX1 I_27390 (I917465,I3563,I469221,I469247,);
DFFARX1 I_27391 (I469247,I3563,I469221,I469264,);
not I_27392 (I469213,I469264);
not I_27393 (I469286,I469247);
nand I_27394 (I469303,I917480,I917468);
and I_27395 (I469320,I469303,I917459);
DFFARX1 I_27396 (I469320,I3563,I469221,I469346,);
not I_27397 (I469354,I469346);
DFFARX1 I_27398 (I917471,I3563,I469221,I469380,);
and I_27399 (I469388,I469380,I917462);
nand I_27400 (I469405,I469380,I917462);
nand I_27401 (I469192,I469354,I469405);
DFFARX1 I_27402 (I917477,I3563,I469221,I469445,);
nor I_27403 (I469453,I469445,I469388);
DFFARX1 I_27404 (I469453,I3563,I469221,I469186,);
nor I_27405 (I469201,I469445,I469346);
nand I_27406 (I469498,I917486,I917474);
and I_27407 (I469515,I469498,I917483);
DFFARX1 I_27408 (I469515,I3563,I469221,I469541,);
nor I_27409 (I469189,I469541,I469445);
not I_27410 (I469563,I469541);
nor I_27411 (I469580,I469563,I469354);
nor I_27412 (I469597,I469286,I469580);
DFFARX1 I_27413 (I469597,I3563,I469221,I469204,);
nor I_27414 (I469628,I469563,I469445);
nor I_27415 (I469645,I917459,I917474);
nor I_27416 (I469195,I469645,I469628);
not I_27417 (I469676,I469645);
nand I_27418 (I469198,I469405,I469676);
DFFARX1 I_27419 (I469645,I3563,I469221,I469210,);
DFFARX1 I_27420 (I469645,I3563,I469221,I469207,);
not I_27421 (I469765,I3570);
DFFARX1 I_27422 (I608130,I3563,I469765,I469791,);
DFFARX1 I_27423 (I469791,I3563,I469765,I469808,);
not I_27424 (I469757,I469808);
not I_27425 (I469830,I469791);
nand I_27426 (I469847,I608127,I608148);
and I_27427 (I469864,I469847,I608151);
DFFARX1 I_27428 (I469864,I3563,I469765,I469890,);
not I_27429 (I469898,I469890);
DFFARX1 I_27430 (I608136,I3563,I469765,I469924,);
and I_27431 (I469932,I469924,I608139);
nand I_27432 (I469949,I469924,I608139);
nand I_27433 (I469736,I469898,I469949);
DFFARX1 I_27434 (I608142,I3563,I469765,I469989,);
nor I_27435 (I469997,I469989,I469932);
DFFARX1 I_27436 (I469997,I3563,I469765,I469730,);
nor I_27437 (I469745,I469989,I469890);
nand I_27438 (I470042,I608127,I608133);
and I_27439 (I470059,I470042,I608145);
DFFARX1 I_27440 (I470059,I3563,I469765,I470085,);
nor I_27441 (I469733,I470085,I469989);
not I_27442 (I470107,I470085);
nor I_27443 (I470124,I470107,I469898);
nor I_27444 (I470141,I469830,I470124);
DFFARX1 I_27445 (I470141,I3563,I469765,I469748,);
nor I_27446 (I470172,I470107,I469989);
nor I_27447 (I470189,I608130,I608133);
nor I_27448 (I469739,I470189,I470172);
not I_27449 (I470220,I470189);
nand I_27450 (I469742,I469949,I470220);
DFFARX1 I_27451 (I470189,I3563,I469765,I469754,);
DFFARX1 I_27452 (I470189,I3563,I469765,I469751,);
not I_27453 (I470309,I3570);
DFFARX1 I_27454 (I8351,I3563,I470309,I470335,);
DFFARX1 I_27455 (I470335,I3563,I470309,I470352,);
not I_27456 (I470301,I470352);
not I_27457 (I470374,I470335);
nand I_27458 (I470391,I8354,I8342);
and I_27459 (I470408,I470391,I8348);
DFFARX1 I_27460 (I470408,I3563,I470309,I470434,);
not I_27461 (I470442,I470434);
DFFARX1 I_27462 (I8336,I3563,I470309,I470468,);
and I_27463 (I470476,I470468,I8333);
nand I_27464 (I470493,I470468,I8333);
nand I_27465 (I470280,I470442,I470493);
DFFARX1 I_27466 (I8339,I3563,I470309,I470533,);
nor I_27467 (I470541,I470533,I470476);
DFFARX1 I_27468 (I470541,I3563,I470309,I470274,);
nor I_27469 (I470289,I470533,I470434);
nand I_27470 (I470586,I8339,I8336);
and I_27471 (I470603,I470586,I8333);
DFFARX1 I_27472 (I470603,I3563,I470309,I470629,);
nor I_27473 (I470277,I470629,I470533);
not I_27474 (I470651,I470629);
nor I_27475 (I470668,I470651,I470442);
nor I_27476 (I470685,I470374,I470668);
DFFARX1 I_27477 (I470685,I3563,I470309,I470292,);
nor I_27478 (I470716,I470651,I470533);
nor I_27479 (I470733,I8345,I8336);
nor I_27480 (I470283,I470733,I470716);
not I_27481 (I470764,I470733);
nand I_27482 (I470286,I470493,I470764);
DFFARX1 I_27483 (I470733,I3563,I470309,I470298,);
DFFARX1 I_27484 (I470733,I3563,I470309,I470295,);
not I_27485 (I470853,I3570);
DFFARX1 I_27486 (I200612,I3563,I470853,I470879,);
DFFARX1 I_27487 (I470879,I3563,I470853,I470896,);
not I_27488 (I470845,I470896);
not I_27489 (I470918,I470879);
nand I_27490 (I470935,I200624,I200603);
and I_27491 (I470952,I470935,I200606);
DFFARX1 I_27492 (I470952,I3563,I470853,I470978,);
not I_27493 (I470986,I470978);
DFFARX1 I_27494 (I200615,I3563,I470853,I471012,);
and I_27495 (I471020,I471012,I200627);
nand I_27496 (I471037,I471012,I200627);
nand I_27497 (I470824,I470986,I471037);
DFFARX1 I_27498 (I200621,I3563,I470853,I471077,);
nor I_27499 (I471085,I471077,I471020);
DFFARX1 I_27500 (I471085,I3563,I470853,I470818,);
nor I_27501 (I470833,I471077,I470978);
nand I_27502 (I471130,I200609,I200606);
and I_27503 (I471147,I471130,I200618);
DFFARX1 I_27504 (I471147,I3563,I470853,I471173,);
nor I_27505 (I470821,I471173,I471077);
not I_27506 (I471195,I471173);
nor I_27507 (I471212,I471195,I470986);
nor I_27508 (I471229,I470918,I471212);
DFFARX1 I_27509 (I471229,I3563,I470853,I470836,);
nor I_27510 (I471260,I471195,I471077);
nor I_27511 (I471277,I200603,I200606);
nor I_27512 (I470827,I471277,I471260);
not I_27513 (I471308,I471277);
nand I_27514 (I470830,I471037,I471308);
DFFARX1 I_27515 (I471277,I3563,I470853,I470842,);
DFFARX1 I_27516 (I471277,I3563,I470853,I470839,);
not I_27517 (I471397,I3570);
DFFARX1 I_27518 (I1363685,I3563,I471397,I471423,);
DFFARX1 I_27519 (I471423,I3563,I471397,I471440,);
not I_27520 (I471389,I471440);
not I_27521 (I471462,I471423);
nand I_27522 (I471479,I1363661,I1363682);
and I_27523 (I471496,I471479,I1363679);
DFFARX1 I_27524 (I471496,I3563,I471397,I471522,);
not I_27525 (I471530,I471522);
DFFARX1 I_27526 (I1363658,I3563,I471397,I471556,);
and I_27527 (I471564,I471556,I1363670);
nand I_27528 (I471581,I471556,I1363670);
nand I_27529 (I471368,I471530,I471581);
DFFARX1 I_27530 (I1363673,I3563,I471397,I471621,);
nor I_27531 (I471629,I471621,I471564);
DFFARX1 I_27532 (I471629,I3563,I471397,I471362,);
nor I_27533 (I471377,I471621,I471522);
nand I_27534 (I471674,I1363676,I1363664);
and I_27535 (I471691,I471674,I1363667);
DFFARX1 I_27536 (I471691,I3563,I471397,I471717,);
nor I_27537 (I471365,I471717,I471621);
not I_27538 (I471739,I471717);
nor I_27539 (I471756,I471739,I471530);
nor I_27540 (I471773,I471462,I471756);
DFFARX1 I_27541 (I471773,I3563,I471397,I471380,);
nor I_27542 (I471804,I471739,I471621);
nor I_27543 (I471821,I1363658,I1363664);
nor I_27544 (I471371,I471821,I471804);
not I_27545 (I471852,I471821);
nand I_27546 (I471374,I471581,I471852);
DFFARX1 I_27547 (I471821,I3563,I471397,I471386,);
DFFARX1 I_27548 (I471821,I3563,I471397,I471383,);
not I_27549 (I471941,I3570);
DFFARX1 I_27550 (I1323029,I3563,I471941,I471967,);
DFFARX1 I_27551 (I471967,I3563,I471941,I471984,);
not I_27552 (I471933,I471984);
not I_27553 (I472006,I471967);
nand I_27554 (I472023,I1323026,I1323023);
and I_27555 (I472040,I472023,I1323011);
DFFARX1 I_27556 (I472040,I3563,I471941,I472066,);
not I_27557 (I472074,I472066);
DFFARX1 I_27558 (I1323035,I3563,I471941,I472100,);
and I_27559 (I472108,I472100,I1323020);
nand I_27560 (I472125,I472100,I1323020);
nand I_27561 (I471912,I472074,I472125);
DFFARX1 I_27562 (I1323014,I3563,I471941,I472165,);
nor I_27563 (I472173,I472165,I472108);
DFFARX1 I_27564 (I472173,I3563,I471941,I471906,);
nor I_27565 (I471921,I472165,I472066);
nand I_27566 (I472218,I1323011,I1323017);
and I_27567 (I472235,I472218,I1323032);
DFFARX1 I_27568 (I472235,I3563,I471941,I472261,);
nor I_27569 (I471909,I472261,I472165);
not I_27570 (I472283,I472261);
nor I_27571 (I472300,I472283,I472074);
nor I_27572 (I472317,I472006,I472300);
DFFARX1 I_27573 (I472317,I3563,I471941,I471924,);
nor I_27574 (I472348,I472283,I472165);
nor I_27575 (I472365,I1323014,I1323017);
nor I_27576 (I471915,I472365,I472348);
not I_27577 (I472396,I472365);
nand I_27578 (I471918,I472125,I472396);
DFFARX1 I_27579 (I472365,I3563,I471941,I471930,);
DFFARX1 I_27580 (I472365,I3563,I471941,I471927,);
not I_27581 (I472485,I3570);
DFFARX1 I_27582 (I698298,I3563,I472485,I472511,);
DFFARX1 I_27583 (I472511,I3563,I472485,I472528,);
not I_27584 (I472477,I472528);
not I_27585 (I472550,I472511);
nand I_27586 (I472567,I698319,I698310);
and I_27587 (I472584,I472567,I698298);
DFFARX1 I_27588 (I472584,I3563,I472485,I472610,);
not I_27589 (I472618,I472610);
DFFARX1 I_27590 (I698304,I3563,I472485,I472644,);
and I_27591 (I472652,I472644,I698301);
nand I_27592 (I472669,I472644,I698301);
nand I_27593 (I472456,I472618,I472669);
DFFARX1 I_27594 (I698295,I3563,I472485,I472709,);
nor I_27595 (I472717,I472709,I472652);
DFFARX1 I_27596 (I472717,I3563,I472485,I472450,);
nor I_27597 (I472465,I472709,I472610);
nand I_27598 (I472762,I698295,I698307);
and I_27599 (I472779,I472762,I698316);
DFFARX1 I_27600 (I472779,I3563,I472485,I472805,);
nor I_27601 (I472453,I472805,I472709);
not I_27602 (I472827,I472805);
nor I_27603 (I472844,I472827,I472618);
nor I_27604 (I472861,I472550,I472844);
DFFARX1 I_27605 (I472861,I3563,I472485,I472468,);
nor I_27606 (I472892,I472827,I472709);
nor I_27607 (I472909,I698313,I698307);
nor I_27608 (I472459,I472909,I472892);
not I_27609 (I472940,I472909);
nand I_27610 (I472462,I472669,I472940);
DFFARX1 I_27611 (I472909,I3563,I472485,I472474,);
DFFARX1 I_27612 (I472909,I3563,I472485,I472471,);
not I_27613 (I473029,I3570);
DFFARX1 I_27614 (I1350000,I3563,I473029,I473055,);
DFFARX1 I_27615 (I473055,I3563,I473029,I473072,);
not I_27616 (I473021,I473072);
not I_27617 (I473094,I473055);
nand I_27618 (I473111,I1349976,I1349997);
and I_27619 (I473128,I473111,I1349994);
DFFARX1 I_27620 (I473128,I3563,I473029,I473154,);
not I_27621 (I473162,I473154);
DFFARX1 I_27622 (I1349973,I3563,I473029,I473188,);
and I_27623 (I473196,I473188,I1349985);
nand I_27624 (I473213,I473188,I1349985);
nand I_27625 (I473000,I473162,I473213);
DFFARX1 I_27626 (I1349988,I3563,I473029,I473253,);
nor I_27627 (I473261,I473253,I473196);
DFFARX1 I_27628 (I473261,I3563,I473029,I472994,);
nor I_27629 (I473009,I473253,I473154);
nand I_27630 (I473306,I1349991,I1349979);
and I_27631 (I473323,I473306,I1349982);
DFFARX1 I_27632 (I473323,I3563,I473029,I473349,);
nor I_27633 (I472997,I473349,I473253);
not I_27634 (I473371,I473349);
nor I_27635 (I473388,I473371,I473162);
nor I_27636 (I473405,I473094,I473388);
DFFARX1 I_27637 (I473405,I3563,I473029,I473012,);
nor I_27638 (I473436,I473371,I473253);
nor I_27639 (I473453,I1349973,I1349979);
nor I_27640 (I473003,I473453,I473436);
not I_27641 (I473484,I473453);
nand I_27642 (I473006,I473213,I473484);
DFFARX1 I_27643 (I473453,I3563,I473029,I473018,);
DFFARX1 I_27644 (I473453,I3563,I473029,I473015,);
not I_27645 (I473573,I3570);
DFFARX1 I_27646 (I408177,I3563,I473573,I473599,);
DFFARX1 I_27647 (I473599,I3563,I473573,I473616,);
not I_27648 (I473565,I473616);
not I_27649 (I473638,I473599);
nand I_27650 (I473655,I408156,I408180);
and I_27651 (I473672,I473655,I408183);
DFFARX1 I_27652 (I473672,I3563,I473573,I473698,);
not I_27653 (I473706,I473698);
DFFARX1 I_27654 (I408165,I3563,I473573,I473732,);
and I_27655 (I473740,I473732,I408171);
nand I_27656 (I473757,I473732,I408171);
nand I_27657 (I473544,I473706,I473757);
DFFARX1 I_27658 (I408159,I3563,I473573,I473797,);
nor I_27659 (I473805,I473797,I473740);
DFFARX1 I_27660 (I473805,I3563,I473573,I473538,);
nor I_27661 (I473553,I473797,I473698);
nand I_27662 (I473850,I408168,I408156);
and I_27663 (I473867,I473850,I408162);
DFFARX1 I_27664 (I473867,I3563,I473573,I473893,);
nor I_27665 (I473541,I473893,I473797);
not I_27666 (I473915,I473893);
nor I_27667 (I473932,I473915,I473706);
nor I_27668 (I473949,I473638,I473932);
DFFARX1 I_27669 (I473949,I3563,I473573,I473556,);
nor I_27670 (I473980,I473915,I473797);
nor I_27671 (I473997,I408174,I408156);
nor I_27672 (I473547,I473997,I473980);
not I_27673 (I474028,I473997);
nand I_27674 (I473550,I473757,I474028);
DFFARX1 I_27675 (I473997,I3563,I473573,I473562,);
DFFARX1 I_27676 (I473997,I3563,I473573,I473559,);
not I_27677 (I474117,I3570);
DFFARX1 I_27678 (I356004,I3563,I474117,I474143,);
DFFARX1 I_27679 (I474143,I3563,I474117,I474160,);
not I_27680 (I474109,I474160);
not I_27681 (I474182,I474143);
nand I_27682 (I474199,I355983,I356007);
and I_27683 (I474216,I474199,I356010);
DFFARX1 I_27684 (I474216,I3563,I474117,I474242,);
not I_27685 (I474250,I474242);
DFFARX1 I_27686 (I355992,I3563,I474117,I474276,);
and I_27687 (I474284,I474276,I355998);
nand I_27688 (I474301,I474276,I355998);
nand I_27689 (I474088,I474250,I474301);
DFFARX1 I_27690 (I355986,I3563,I474117,I474341,);
nor I_27691 (I474349,I474341,I474284);
DFFARX1 I_27692 (I474349,I3563,I474117,I474082,);
nor I_27693 (I474097,I474341,I474242);
nand I_27694 (I474394,I355995,I355983);
and I_27695 (I474411,I474394,I355989);
DFFARX1 I_27696 (I474411,I3563,I474117,I474437,);
nor I_27697 (I474085,I474437,I474341);
not I_27698 (I474459,I474437);
nor I_27699 (I474476,I474459,I474250);
nor I_27700 (I474493,I474182,I474476);
DFFARX1 I_27701 (I474493,I3563,I474117,I474100,);
nor I_27702 (I474524,I474459,I474341);
nor I_27703 (I474541,I356001,I355983);
nor I_27704 (I474091,I474541,I474524);
not I_27705 (I474572,I474541);
nand I_27706 (I474094,I474301,I474572);
DFFARX1 I_27707 (I474541,I3563,I474117,I474106,);
DFFARX1 I_27708 (I474541,I3563,I474117,I474103,);
not I_27709 (I474661,I3570);
DFFARX1 I_27710 (I147824,I3563,I474661,I474687,);
DFFARX1 I_27711 (I474687,I3563,I474661,I474704,);
not I_27712 (I474653,I474704);
not I_27713 (I474726,I474687);
nand I_27714 (I474743,I147839,I147818);
and I_27715 (I474760,I474743,I147821);
DFFARX1 I_27716 (I474760,I3563,I474661,I474786,);
not I_27717 (I474794,I474786);
DFFARX1 I_27718 (I147827,I3563,I474661,I474820,);
and I_27719 (I474828,I474820,I147821);
nand I_27720 (I474845,I474820,I147821);
nand I_27721 (I474632,I474794,I474845);
DFFARX1 I_27722 (I147836,I3563,I474661,I474885,);
nor I_27723 (I474893,I474885,I474828);
DFFARX1 I_27724 (I474893,I3563,I474661,I474626,);
nor I_27725 (I474641,I474885,I474786);
nand I_27726 (I474938,I147818,I147833);
and I_27727 (I474955,I474938,I147830);
DFFARX1 I_27728 (I474955,I3563,I474661,I474981,);
nor I_27729 (I474629,I474981,I474885);
not I_27730 (I475003,I474981);
nor I_27731 (I475020,I475003,I474794);
nor I_27732 (I475037,I474726,I475020);
DFFARX1 I_27733 (I475037,I3563,I474661,I474644,);
nor I_27734 (I475068,I475003,I474885);
nor I_27735 (I475085,I147842,I147833);
nor I_27736 (I474635,I475085,I475068);
not I_27737 (I475116,I475085);
nand I_27738 (I474638,I474845,I475116);
DFFARX1 I_27739 (I475085,I3563,I474661,I474650,);
DFFARX1 I_27740 (I475085,I3563,I474661,I474647,);
not I_27741 (I475205,I3570);
DFFARX1 I_27742 (I994339,I3563,I475205,I475231,);
DFFARX1 I_27743 (I475231,I3563,I475205,I475248,);
not I_27744 (I475197,I475248);
not I_27745 (I475270,I475231);
nand I_27746 (I475287,I994354,I994342);
and I_27747 (I475304,I475287,I994333);
DFFARX1 I_27748 (I475304,I3563,I475205,I475330,);
not I_27749 (I475338,I475330);
DFFARX1 I_27750 (I994345,I3563,I475205,I475364,);
and I_27751 (I475372,I475364,I994336);
nand I_27752 (I475389,I475364,I994336);
nand I_27753 (I475176,I475338,I475389);
DFFARX1 I_27754 (I994351,I3563,I475205,I475429,);
nor I_27755 (I475437,I475429,I475372);
DFFARX1 I_27756 (I475437,I3563,I475205,I475170,);
nor I_27757 (I475185,I475429,I475330);
nand I_27758 (I475482,I994360,I994348);
and I_27759 (I475499,I475482,I994357);
DFFARX1 I_27760 (I475499,I3563,I475205,I475525,);
nor I_27761 (I475173,I475525,I475429);
not I_27762 (I475547,I475525);
nor I_27763 (I475564,I475547,I475338);
nor I_27764 (I475581,I475270,I475564);
DFFARX1 I_27765 (I475581,I3563,I475205,I475188,);
nor I_27766 (I475612,I475547,I475429);
nor I_27767 (I475629,I994333,I994348);
nor I_27768 (I475179,I475629,I475612);
not I_27769 (I475660,I475629);
nand I_27770 (I475182,I475389,I475660);
DFFARX1 I_27771 (I475629,I3563,I475205,I475194,);
DFFARX1 I_27772 (I475629,I3563,I475205,I475191,);
not I_27773 (I475749,I3570);
DFFARX1 I_27774 (I1002091,I3563,I475749,I475775,);
DFFARX1 I_27775 (I475775,I3563,I475749,I475792,);
not I_27776 (I475741,I475792);
not I_27777 (I475814,I475775);
nand I_27778 (I475831,I1002106,I1002094);
and I_27779 (I475848,I475831,I1002085);
DFFARX1 I_27780 (I475848,I3563,I475749,I475874,);
not I_27781 (I475882,I475874);
DFFARX1 I_27782 (I1002097,I3563,I475749,I475908,);
and I_27783 (I475916,I475908,I1002088);
nand I_27784 (I475933,I475908,I1002088);
nand I_27785 (I475720,I475882,I475933);
DFFARX1 I_27786 (I1002103,I3563,I475749,I475973,);
nor I_27787 (I475981,I475973,I475916);
DFFARX1 I_27788 (I475981,I3563,I475749,I475714,);
nor I_27789 (I475729,I475973,I475874);
nand I_27790 (I476026,I1002112,I1002100);
and I_27791 (I476043,I476026,I1002109);
DFFARX1 I_27792 (I476043,I3563,I475749,I476069,);
nor I_27793 (I475717,I476069,I475973);
not I_27794 (I476091,I476069);
nor I_27795 (I476108,I476091,I475882);
nor I_27796 (I476125,I475814,I476108);
DFFARX1 I_27797 (I476125,I3563,I475749,I475732,);
nor I_27798 (I476156,I476091,I475973);
nor I_27799 (I476173,I1002085,I1002100);
nor I_27800 (I475723,I476173,I476156);
not I_27801 (I476204,I476173);
nand I_27802 (I475726,I475933,I476204);
DFFARX1 I_27803 (I476173,I3563,I475749,I475738,);
DFFARX1 I_27804 (I476173,I3563,I475749,I475735,);
not I_27805 (I476293,I3570);
DFFARX1 I_27806 (I883794,I3563,I476293,I476319,);
DFFARX1 I_27807 (I476319,I3563,I476293,I476336,);
not I_27808 (I476285,I476336);
not I_27809 (I476358,I476319);
nand I_27810 (I476375,I883788,I883785);
and I_27811 (I476392,I476375,I883800);
DFFARX1 I_27812 (I476392,I3563,I476293,I476418,);
not I_27813 (I476426,I476418);
DFFARX1 I_27814 (I883788,I3563,I476293,I476452,);
and I_27815 (I476460,I476452,I883782);
nand I_27816 (I476477,I476452,I883782);
nand I_27817 (I476264,I476426,I476477);
DFFARX1 I_27818 (I883782,I3563,I476293,I476517,);
nor I_27819 (I476525,I476517,I476460);
DFFARX1 I_27820 (I476525,I3563,I476293,I476258,);
nor I_27821 (I476273,I476517,I476418);
nand I_27822 (I476570,I883797,I883791);
and I_27823 (I476587,I476570,I883785);
DFFARX1 I_27824 (I476587,I3563,I476293,I476613,);
nor I_27825 (I476261,I476613,I476517);
not I_27826 (I476635,I476613);
nor I_27827 (I476652,I476635,I476426);
nor I_27828 (I476669,I476358,I476652);
DFFARX1 I_27829 (I476669,I3563,I476293,I476276,);
nor I_27830 (I476700,I476635,I476517);
nor I_27831 (I476717,I883803,I883791);
nor I_27832 (I476267,I476717,I476700);
not I_27833 (I476748,I476717);
nand I_27834 (I476270,I476477,I476748);
DFFARX1 I_27835 (I476717,I3563,I476293,I476282,);
DFFARX1 I_27836 (I476717,I3563,I476293,I476279,);
not I_27837 (I476837,I3570);
DFFARX1 I_27838 (I1262188,I3563,I476837,I476863,);
DFFARX1 I_27839 (I476863,I3563,I476837,I476880,);
not I_27840 (I476829,I476880);
not I_27841 (I476902,I476863);
nand I_27842 (I476919,I1262200,I1262203);
and I_27843 (I476936,I476919,I1262206);
DFFARX1 I_27844 (I476936,I3563,I476837,I476962,);
not I_27845 (I476970,I476962);
DFFARX1 I_27846 (I1262191,I3563,I476837,I476996,);
and I_27847 (I477004,I476996,I1262197);
nand I_27848 (I477021,I476996,I1262197);
nand I_27849 (I476808,I476970,I477021);
DFFARX1 I_27850 (I1262185,I3563,I476837,I477061,);
nor I_27851 (I477069,I477061,I477004);
DFFARX1 I_27852 (I477069,I3563,I476837,I476802,);
nor I_27853 (I476817,I477061,I476962);
nand I_27854 (I477114,I1262188,I1262209);
and I_27855 (I477131,I477114,I1262194);
DFFARX1 I_27856 (I477131,I3563,I476837,I477157,);
nor I_27857 (I476805,I477157,I477061);
not I_27858 (I477179,I477157);
nor I_27859 (I477196,I477179,I476970);
nor I_27860 (I477213,I476902,I477196);
DFFARX1 I_27861 (I477213,I3563,I476837,I476820,);
nor I_27862 (I477244,I477179,I477061);
nor I_27863 (I477261,I1262185,I1262209);
nor I_27864 (I476811,I477261,I477244);
not I_27865 (I477292,I477261);
nand I_27866 (I476814,I477021,I477292);
DFFARX1 I_27867 (I477261,I3563,I476837,I476826,);
DFFARX1 I_27868 (I477261,I3563,I476837,I476823,);
not I_27869 (I477381,I3570);
DFFARX1 I_27870 (I57186,I3563,I477381,I477407,);
DFFARX1 I_27871 (I477407,I3563,I477381,I477424,);
not I_27872 (I477373,I477424);
not I_27873 (I477446,I477407);
nand I_27874 (I477463,I57174,I57189);
and I_27875 (I477480,I477463,I57177);
DFFARX1 I_27876 (I477480,I3563,I477381,I477506,);
not I_27877 (I477514,I477506);
DFFARX1 I_27878 (I57198,I3563,I477381,I477540,);
and I_27879 (I477548,I477540,I57192);
nand I_27880 (I477565,I477540,I57192);
nand I_27881 (I477352,I477514,I477565);
DFFARX1 I_27882 (I57195,I3563,I477381,I477605,);
nor I_27883 (I477613,I477605,I477548);
DFFARX1 I_27884 (I477613,I3563,I477381,I477346,);
nor I_27885 (I477361,I477605,I477506);
nand I_27886 (I477658,I57174,I57177);
and I_27887 (I477675,I477658,I57180);
DFFARX1 I_27888 (I477675,I3563,I477381,I477701,);
nor I_27889 (I477349,I477701,I477605);
not I_27890 (I477723,I477701);
nor I_27891 (I477740,I477723,I477514);
nor I_27892 (I477757,I477446,I477740);
DFFARX1 I_27893 (I477757,I3563,I477381,I477364,);
nor I_27894 (I477788,I477723,I477605);
nor I_27895 (I477805,I57183,I57177);
nor I_27896 (I477355,I477805,I477788);
not I_27897 (I477836,I477805);
nand I_27898 (I477358,I477565,I477836);
DFFARX1 I_27899 (I477805,I3563,I477381,I477370,);
DFFARX1 I_27900 (I477805,I3563,I477381,I477367,);
not I_27901 (I477925,I3570);
DFFARX1 I_27902 (I862187,I3563,I477925,I477951,);
DFFARX1 I_27903 (I477951,I3563,I477925,I477968,);
not I_27904 (I477917,I477968);
not I_27905 (I477990,I477951);
nand I_27906 (I478007,I862181,I862178);
and I_27907 (I478024,I478007,I862193);
DFFARX1 I_27908 (I478024,I3563,I477925,I478050,);
not I_27909 (I478058,I478050);
DFFARX1 I_27910 (I862181,I3563,I477925,I478084,);
and I_27911 (I478092,I478084,I862175);
nand I_27912 (I478109,I478084,I862175);
nand I_27913 (I477896,I478058,I478109);
DFFARX1 I_27914 (I862175,I3563,I477925,I478149,);
nor I_27915 (I478157,I478149,I478092);
DFFARX1 I_27916 (I478157,I3563,I477925,I477890,);
nor I_27917 (I477905,I478149,I478050);
nand I_27918 (I478202,I862190,I862184);
and I_27919 (I478219,I478202,I862178);
DFFARX1 I_27920 (I478219,I3563,I477925,I478245,);
nor I_27921 (I477893,I478245,I478149);
not I_27922 (I478267,I478245);
nor I_27923 (I478284,I478267,I478058);
nor I_27924 (I478301,I477990,I478284);
DFFARX1 I_27925 (I478301,I3563,I477925,I477908,);
nor I_27926 (I478332,I478267,I478149);
nor I_27927 (I478349,I862196,I862184);
nor I_27928 (I477899,I478349,I478332);
not I_27929 (I478380,I478349);
nand I_27930 (I477902,I478109,I478380);
DFFARX1 I_27931 (I478349,I3563,I477925,I477914,);
DFFARX1 I_27932 (I478349,I3563,I477925,I477911,);
not I_27933 (I478469,I3570);
DFFARX1 I_27934 (I1248588,I3563,I478469,I478495,);
DFFARX1 I_27935 (I478495,I3563,I478469,I478512,);
not I_27936 (I478461,I478512);
not I_27937 (I478534,I478495);
nand I_27938 (I478551,I1248600,I1248603);
and I_27939 (I478568,I478551,I1248606);
DFFARX1 I_27940 (I478568,I3563,I478469,I478594,);
not I_27941 (I478602,I478594);
DFFARX1 I_27942 (I1248591,I3563,I478469,I478628,);
and I_27943 (I478636,I478628,I1248597);
nand I_27944 (I478653,I478628,I1248597);
nand I_27945 (I478440,I478602,I478653);
DFFARX1 I_27946 (I1248585,I3563,I478469,I478693,);
nor I_27947 (I478701,I478693,I478636);
DFFARX1 I_27948 (I478701,I3563,I478469,I478434,);
nor I_27949 (I478449,I478693,I478594);
nand I_27950 (I478746,I1248588,I1248609);
and I_27951 (I478763,I478746,I1248594);
DFFARX1 I_27952 (I478763,I3563,I478469,I478789,);
nor I_27953 (I478437,I478789,I478693);
not I_27954 (I478811,I478789);
nor I_27955 (I478828,I478811,I478602);
nor I_27956 (I478845,I478534,I478828);
DFFARX1 I_27957 (I478845,I3563,I478469,I478452,);
nor I_27958 (I478876,I478811,I478693);
nor I_27959 (I478893,I1248585,I1248609);
nor I_27960 (I478443,I478893,I478876);
not I_27961 (I478924,I478893);
nand I_27962 (I478446,I478653,I478924);
DFFARX1 I_27963 (I478893,I3563,I478469,I478458,);
DFFARX1 I_27964 (I478893,I3563,I478469,I478455,);
not I_27965 (I479013,I3570);
DFFARX1 I_27966 (I1125100,I3563,I479013,I479039,);
DFFARX1 I_27967 (I479039,I3563,I479013,I479056,);
not I_27968 (I479005,I479056);
not I_27969 (I479078,I479039);
nand I_27970 (I479095,I1125112,I1125100);
and I_27971 (I479112,I479095,I1125103);
DFFARX1 I_27972 (I479112,I3563,I479013,I479138,);
not I_27973 (I479146,I479138);
DFFARX1 I_27974 (I1125121,I3563,I479013,I479172,);
and I_27975 (I479180,I479172,I1125097);
nand I_27976 (I479197,I479172,I1125097);
nand I_27977 (I478984,I479146,I479197);
DFFARX1 I_27978 (I1125115,I3563,I479013,I479237,);
nor I_27979 (I479245,I479237,I479180);
DFFARX1 I_27980 (I479245,I3563,I479013,I478978,);
nor I_27981 (I478993,I479237,I479138);
nand I_27982 (I479290,I1125109,I1125106);
and I_27983 (I479307,I479290,I1125118);
DFFARX1 I_27984 (I479307,I3563,I479013,I479333,);
nor I_27985 (I478981,I479333,I479237);
not I_27986 (I479355,I479333);
nor I_27987 (I479372,I479355,I479146);
nor I_27988 (I479389,I479078,I479372);
DFFARX1 I_27989 (I479389,I3563,I479013,I478996,);
nor I_27990 (I479420,I479355,I479237);
nor I_27991 (I479437,I1125097,I1125106);
nor I_27992 (I478987,I479437,I479420);
not I_27993 (I479468,I479437);
nand I_27994 (I478990,I479197,I479468);
DFFARX1 I_27995 (I479437,I3563,I479013,I479002,);
DFFARX1 I_27996 (I479437,I3563,I479013,I478999,);
not I_27997 (I479557,I3570);
DFFARX1 I_27998 (I720262,I3563,I479557,I479583,);
DFFARX1 I_27999 (I479583,I3563,I479557,I479600,);
not I_28000 (I479549,I479600);
not I_28001 (I479622,I479583);
nand I_28002 (I479639,I720283,I720274);
and I_28003 (I479656,I479639,I720262);
DFFARX1 I_28004 (I479656,I3563,I479557,I479682,);
not I_28005 (I479690,I479682);
DFFARX1 I_28006 (I720268,I3563,I479557,I479716,);
and I_28007 (I479724,I479716,I720265);
nand I_28008 (I479741,I479716,I720265);
nand I_28009 (I479528,I479690,I479741);
DFFARX1 I_28010 (I720259,I3563,I479557,I479781,);
nor I_28011 (I479789,I479781,I479724);
DFFARX1 I_28012 (I479789,I3563,I479557,I479522,);
nor I_28013 (I479537,I479781,I479682);
nand I_28014 (I479834,I720259,I720271);
and I_28015 (I479851,I479834,I720280);
DFFARX1 I_28016 (I479851,I3563,I479557,I479877,);
nor I_28017 (I479525,I479877,I479781);
not I_28018 (I479899,I479877);
nor I_28019 (I479916,I479899,I479690);
nor I_28020 (I479933,I479622,I479916);
DFFARX1 I_28021 (I479933,I3563,I479557,I479540,);
nor I_28022 (I479964,I479899,I479781);
nor I_28023 (I479981,I720277,I720271);
nor I_28024 (I479531,I479981,I479964);
not I_28025 (I480012,I479981);
nand I_28026 (I479534,I479741,I480012);
DFFARX1 I_28027 (I479981,I3563,I479557,I479546,);
DFFARX1 I_28028 (I479981,I3563,I479557,I479543,);
not I_28029 (I480101,I3570);
DFFARX1 I_28030 (I1173652,I3563,I480101,I480127,);
DFFARX1 I_28031 (I480127,I3563,I480101,I480144,);
not I_28032 (I480093,I480144);
not I_28033 (I480166,I480127);
nand I_28034 (I480183,I1173664,I1173652);
and I_28035 (I480200,I480183,I1173655);
DFFARX1 I_28036 (I480200,I3563,I480101,I480226,);
not I_28037 (I480234,I480226);
DFFARX1 I_28038 (I1173673,I3563,I480101,I480260,);
and I_28039 (I480268,I480260,I1173649);
nand I_28040 (I480285,I480260,I1173649);
nand I_28041 (I480072,I480234,I480285);
DFFARX1 I_28042 (I1173667,I3563,I480101,I480325,);
nor I_28043 (I480333,I480325,I480268);
DFFARX1 I_28044 (I480333,I3563,I480101,I480066,);
nor I_28045 (I480081,I480325,I480226);
nand I_28046 (I480378,I1173661,I1173658);
and I_28047 (I480395,I480378,I1173670);
DFFARX1 I_28048 (I480395,I3563,I480101,I480421,);
nor I_28049 (I480069,I480421,I480325);
not I_28050 (I480443,I480421);
nor I_28051 (I480460,I480443,I480234);
nor I_28052 (I480477,I480166,I480460);
DFFARX1 I_28053 (I480477,I3563,I480101,I480084,);
nor I_28054 (I480508,I480443,I480325);
nor I_28055 (I480525,I1173649,I1173658);
nor I_28056 (I480075,I480525,I480508);
not I_28057 (I480556,I480525);
nand I_28058 (I480078,I480285,I480556);
DFFARX1 I_28059 (I480525,I3563,I480101,I480090,);
DFFARX1 I_28060 (I480525,I3563,I480101,I480087,);
not I_28061 (I480645,I3570);
DFFARX1 I_28062 (I562009,I3563,I480645,I480671,);
DFFARX1 I_28063 (I480671,I3563,I480645,I480688,);
not I_28064 (I480637,I480688);
not I_28065 (I480710,I480671);
nand I_28066 (I480727,I562012,I562030);
and I_28067 (I480744,I480727,I562018);
DFFARX1 I_28068 (I480744,I3563,I480645,I480770,);
not I_28069 (I480778,I480770);
DFFARX1 I_28070 (I562009,I3563,I480645,I480804,);
and I_28071 (I480812,I480804,I562027);
nand I_28072 (I480829,I480804,I562027);
nand I_28073 (I480616,I480778,I480829);
DFFARX1 I_28074 (I562021,I3563,I480645,I480869,);
nor I_28075 (I480877,I480869,I480812);
DFFARX1 I_28076 (I480877,I3563,I480645,I480610,);
nor I_28077 (I480625,I480869,I480770);
nand I_28078 (I480922,I562024,I562006);
and I_28079 (I480939,I480922,I562015);
DFFARX1 I_28080 (I480939,I3563,I480645,I480965,);
nor I_28081 (I480613,I480965,I480869);
not I_28082 (I480987,I480965);
nor I_28083 (I481004,I480987,I480778);
nor I_28084 (I481021,I480710,I481004);
DFFARX1 I_28085 (I481021,I3563,I480645,I480628,);
nor I_28086 (I481052,I480987,I480869);
nor I_28087 (I481069,I562006,I562006);
nor I_28088 (I480619,I481069,I481052);
not I_28089 (I481100,I481069);
nand I_28090 (I480622,I480829,I481100);
DFFARX1 I_28091 (I481069,I3563,I480645,I480634,);
DFFARX1 I_28092 (I481069,I3563,I480645,I480631,);
not I_28093 (I481189,I3570);
DFFARX1 I_28094 (I986587,I3563,I481189,I481215,);
DFFARX1 I_28095 (I481215,I3563,I481189,I481232,);
not I_28096 (I481181,I481232);
not I_28097 (I481254,I481215);
nand I_28098 (I481271,I986602,I986590);
and I_28099 (I481288,I481271,I986581);
DFFARX1 I_28100 (I481288,I3563,I481189,I481314,);
not I_28101 (I481322,I481314);
DFFARX1 I_28102 (I986593,I3563,I481189,I481348,);
and I_28103 (I481356,I481348,I986584);
nand I_28104 (I481373,I481348,I986584);
nand I_28105 (I481160,I481322,I481373);
DFFARX1 I_28106 (I986599,I3563,I481189,I481413,);
nor I_28107 (I481421,I481413,I481356);
DFFARX1 I_28108 (I481421,I3563,I481189,I481154,);
nor I_28109 (I481169,I481413,I481314);
nand I_28110 (I481466,I986608,I986596);
and I_28111 (I481483,I481466,I986605);
DFFARX1 I_28112 (I481483,I3563,I481189,I481509,);
nor I_28113 (I481157,I481509,I481413);
not I_28114 (I481531,I481509);
nor I_28115 (I481548,I481531,I481322);
nor I_28116 (I481565,I481254,I481548);
DFFARX1 I_28117 (I481565,I3563,I481189,I481172,);
nor I_28118 (I481596,I481531,I481413);
nor I_28119 (I481613,I986581,I986596);
nor I_28120 (I481163,I481613,I481596);
not I_28121 (I481644,I481613);
nand I_28122 (I481166,I481373,I481644);
DFFARX1 I_28123 (I481613,I3563,I481189,I481178,);
DFFARX1 I_28124 (I481613,I3563,I481189,I481175,);
not I_28125 (I481733,I3570);
DFFARX1 I_28126 (I914881,I3563,I481733,I481759,);
DFFARX1 I_28127 (I481759,I3563,I481733,I481776,);
not I_28128 (I481725,I481776);
not I_28129 (I481798,I481759);
nand I_28130 (I481815,I914896,I914884);
and I_28131 (I481832,I481815,I914875);
DFFARX1 I_28132 (I481832,I3563,I481733,I481858,);
not I_28133 (I481866,I481858);
DFFARX1 I_28134 (I914887,I3563,I481733,I481892,);
and I_28135 (I481900,I481892,I914878);
nand I_28136 (I481917,I481892,I914878);
nand I_28137 (I481704,I481866,I481917);
DFFARX1 I_28138 (I914893,I3563,I481733,I481957,);
nor I_28139 (I481965,I481957,I481900);
DFFARX1 I_28140 (I481965,I3563,I481733,I481698,);
nor I_28141 (I481713,I481957,I481858);
nand I_28142 (I482010,I914902,I914890);
and I_28143 (I482027,I482010,I914899);
DFFARX1 I_28144 (I482027,I3563,I481733,I482053,);
nor I_28145 (I481701,I482053,I481957);
not I_28146 (I482075,I482053);
nor I_28147 (I482092,I482075,I481866);
nor I_28148 (I482109,I481798,I482092);
DFFARX1 I_28149 (I482109,I3563,I481733,I481716,);
nor I_28150 (I482140,I482075,I481957);
nor I_28151 (I482157,I914875,I914890);
nor I_28152 (I481707,I482157,I482140);
not I_28153 (I482188,I482157);
nand I_28154 (I481710,I481917,I482188);
DFFARX1 I_28155 (I482157,I3563,I481733,I481722,);
DFFARX1 I_28156 (I482157,I3563,I481733,I481719,);
not I_28157 (I482277,I3570);
DFFARX1 I_28158 (I383935,I3563,I482277,I482303,);
DFFARX1 I_28159 (I482303,I3563,I482277,I482320,);
not I_28160 (I482269,I482320);
not I_28161 (I482342,I482303);
nand I_28162 (I482359,I383914,I383938);
and I_28163 (I482376,I482359,I383941);
DFFARX1 I_28164 (I482376,I3563,I482277,I482402,);
not I_28165 (I482410,I482402);
DFFARX1 I_28166 (I383923,I3563,I482277,I482436,);
and I_28167 (I482444,I482436,I383929);
nand I_28168 (I482461,I482436,I383929);
nand I_28169 (I482248,I482410,I482461);
DFFARX1 I_28170 (I383917,I3563,I482277,I482501,);
nor I_28171 (I482509,I482501,I482444);
DFFARX1 I_28172 (I482509,I3563,I482277,I482242,);
nor I_28173 (I482257,I482501,I482402);
nand I_28174 (I482554,I383926,I383914);
and I_28175 (I482571,I482554,I383920);
DFFARX1 I_28176 (I482571,I3563,I482277,I482597,);
nor I_28177 (I482245,I482597,I482501);
not I_28178 (I482619,I482597);
nor I_28179 (I482636,I482619,I482410);
nor I_28180 (I482653,I482342,I482636);
DFFARX1 I_28181 (I482653,I3563,I482277,I482260,);
nor I_28182 (I482684,I482619,I482501);
nor I_28183 (I482701,I383932,I383914);
nor I_28184 (I482251,I482701,I482684);
not I_28185 (I482732,I482701);
nand I_28186 (I482254,I482461,I482732);
DFFARX1 I_28187 (I482701,I3563,I482277,I482266,);
DFFARX1 I_28188 (I482701,I3563,I482277,I482263,);
not I_28189 (I482821,I3570);
DFFARX1 I_28190 (I1236076,I3563,I482821,I482847,);
DFFARX1 I_28191 (I482847,I3563,I482821,I482864,);
not I_28192 (I482813,I482864);
not I_28193 (I482886,I482847);
nand I_28194 (I482903,I1236088,I1236076);
and I_28195 (I482920,I482903,I1236079);
DFFARX1 I_28196 (I482920,I3563,I482821,I482946,);
not I_28197 (I482954,I482946);
DFFARX1 I_28198 (I1236097,I3563,I482821,I482980,);
and I_28199 (I482988,I482980,I1236073);
nand I_28200 (I483005,I482980,I1236073);
nand I_28201 (I482792,I482954,I483005);
DFFARX1 I_28202 (I1236091,I3563,I482821,I483045,);
nor I_28203 (I483053,I483045,I482988);
DFFARX1 I_28204 (I483053,I3563,I482821,I482786,);
nor I_28205 (I482801,I483045,I482946);
nand I_28206 (I483098,I1236085,I1236082);
and I_28207 (I483115,I483098,I1236094);
DFFARX1 I_28208 (I483115,I3563,I482821,I483141,);
nor I_28209 (I482789,I483141,I483045);
not I_28210 (I483163,I483141);
nor I_28211 (I483180,I483163,I482954);
nor I_28212 (I483197,I482886,I483180);
DFFARX1 I_28213 (I483197,I3563,I482821,I482804,);
nor I_28214 (I483228,I483163,I483045);
nor I_28215 (I483245,I1236073,I1236082);
nor I_28216 (I482795,I483245,I483228);
not I_28217 (I483276,I483245);
nand I_28218 (I482798,I483005,I483276);
DFFARX1 I_28219 (I483245,I3563,I482821,I482810,);
DFFARX1 I_28220 (I483245,I3563,I482821,I482807,);
not I_28221 (I483365,I3570);
DFFARX1 I_28222 (I797136,I3563,I483365,I483391,);
DFFARX1 I_28223 (I483391,I3563,I483365,I483408,);
not I_28224 (I483357,I483408);
not I_28225 (I483430,I483391);
nand I_28226 (I483447,I797157,I797148);
and I_28227 (I483464,I483447,I797136);
DFFARX1 I_28228 (I483464,I3563,I483365,I483490,);
not I_28229 (I483498,I483490);
DFFARX1 I_28230 (I797142,I3563,I483365,I483524,);
and I_28231 (I483532,I483524,I797139);
nand I_28232 (I483549,I483524,I797139);
nand I_28233 (I483336,I483498,I483549);
DFFARX1 I_28234 (I797133,I3563,I483365,I483589,);
nor I_28235 (I483597,I483589,I483532);
DFFARX1 I_28236 (I483597,I3563,I483365,I483330,);
nor I_28237 (I483345,I483589,I483490);
nand I_28238 (I483642,I797133,I797145);
and I_28239 (I483659,I483642,I797154);
DFFARX1 I_28240 (I483659,I3563,I483365,I483685,);
nor I_28241 (I483333,I483685,I483589);
not I_28242 (I483707,I483685);
nor I_28243 (I483724,I483707,I483498);
nor I_28244 (I483741,I483430,I483724);
DFFARX1 I_28245 (I483741,I3563,I483365,I483348,);
nor I_28246 (I483772,I483707,I483589);
nor I_28247 (I483789,I797151,I797145);
nor I_28248 (I483339,I483789,I483772);
not I_28249 (I483820,I483789);
nand I_28250 (I483342,I483549,I483820);
DFFARX1 I_28251 (I483789,I3563,I483365,I483354,);
DFFARX1 I_28252 (I483789,I3563,I483365,I483351,);
not I_28253 (I483909,I3570);
DFFARX1 I_28254 (I1306267,I3563,I483909,I483935,);
DFFARX1 I_28255 (I483935,I3563,I483909,I483952,);
not I_28256 (I483901,I483952);
not I_28257 (I483974,I483935);
nand I_28258 (I483991,I1306264,I1306261);
and I_28259 (I484008,I483991,I1306249);
DFFARX1 I_28260 (I484008,I3563,I483909,I484034,);
not I_28261 (I484042,I484034);
DFFARX1 I_28262 (I1306273,I3563,I483909,I484068,);
and I_28263 (I484076,I484068,I1306258);
nand I_28264 (I484093,I484068,I1306258);
nand I_28265 (I483880,I484042,I484093);
DFFARX1 I_28266 (I1306252,I3563,I483909,I484133,);
nor I_28267 (I484141,I484133,I484076);
DFFARX1 I_28268 (I484141,I3563,I483909,I483874,);
nor I_28269 (I483889,I484133,I484034);
nand I_28270 (I484186,I1306249,I1306255);
and I_28271 (I484203,I484186,I1306270);
DFFARX1 I_28272 (I484203,I3563,I483909,I484229,);
nor I_28273 (I483877,I484229,I484133);
not I_28274 (I484251,I484229);
nor I_28275 (I484268,I484251,I484042);
nor I_28276 (I484285,I483974,I484268);
DFFARX1 I_28277 (I484285,I3563,I483909,I483892,);
nor I_28278 (I484316,I484251,I484133);
nor I_28279 (I484333,I1306252,I1306255);
nor I_28280 (I483883,I484333,I484316);
not I_28281 (I484364,I484333);
nand I_28282 (I483886,I484093,I484364);
DFFARX1 I_28283 (I484333,I3563,I483909,I483898,);
DFFARX1 I_28284 (I484333,I3563,I483909,I483895,);
not I_28285 (I484453,I3570);
DFFARX1 I_28286 (I656682,I3563,I484453,I484479,);
DFFARX1 I_28287 (I484479,I3563,I484453,I484496,);
not I_28288 (I484445,I484496);
not I_28289 (I484518,I484479);
nand I_28290 (I484535,I656679,I656700);
and I_28291 (I484552,I484535,I656703);
DFFARX1 I_28292 (I484552,I3563,I484453,I484578,);
not I_28293 (I484586,I484578);
DFFARX1 I_28294 (I656688,I3563,I484453,I484612,);
and I_28295 (I484620,I484612,I656691);
nand I_28296 (I484637,I484612,I656691);
nand I_28297 (I484424,I484586,I484637);
DFFARX1 I_28298 (I656694,I3563,I484453,I484677,);
nor I_28299 (I484685,I484677,I484620);
DFFARX1 I_28300 (I484685,I3563,I484453,I484418,);
nor I_28301 (I484433,I484677,I484578);
nand I_28302 (I484730,I656679,I656685);
and I_28303 (I484747,I484730,I656697);
DFFARX1 I_28304 (I484747,I3563,I484453,I484773,);
nor I_28305 (I484421,I484773,I484677);
not I_28306 (I484795,I484773);
nor I_28307 (I484812,I484795,I484586);
nor I_28308 (I484829,I484518,I484812);
DFFARX1 I_28309 (I484829,I3563,I484453,I484436,);
nor I_28310 (I484860,I484795,I484677);
nor I_28311 (I484877,I656682,I656685);
nor I_28312 (I484427,I484877,I484860);
not I_28313 (I484908,I484877);
nand I_28314 (I484430,I484637,I484908);
DFFARX1 I_28315 (I484877,I3563,I484453,I484442,);
DFFARX1 I_28316 (I484877,I3563,I484453,I484439,);
not I_28317 (I484997,I3570);
DFFARX1 I_28318 (I653792,I3563,I484997,I485023,);
DFFARX1 I_28319 (I485023,I3563,I484997,I485040,);
not I_28320 (I484989,I485040);
not I_28321 (I485062,I485023);
nand I_28322 (I485079,I653789,I653810);
and I_28323 (I485096,I485079,I653813);
DFFARX1 I_28324 (I485096,I3563,I484997,I485122,);
not I_28325 (I485130,I485122);
DFFARX1 I_28326 (I653798,I3563,I484997,I485156,);
and I_28327 (I485164,I485156,I653801);
nand I_28328 (I485181,I485156,I653801);
nand I_28329 (I484968,I485130,I485181);
DFFARX1 I_28330 (I653804,I3563,I484997,I485221,);
nor I_28331 (I485229,I485221,I485164);
DFFARX1 I_28332 (I485229,I3563,I484997,I484962,);
nor I_28333 (I484977,I485221,I485122);
nand I_28334 (I485274,I653789,I653795);
and I_28335 (I485291,I485274,I653807);
DFFARX1 I_28336 (I485291,I3563,I484997,I485317,);
nor I_28337 (I484965,I485317,I485221);
not I_28338 (I485339,I485317);
nor I_28339 (I485356,I485339,I485130);
nor I_28340 (I485373,I485062,I485356);
DFFARX1 I_28341 (I485373,I3563,I484997,I484980,);
nor I_28342 (I485404,I485339,I485221);
nor I_28343 (I485421,I653792,I653795);
nor I_28344 (I484971,I485421,I485404);
not I_28345 (I485452,I485421);
nand I_28346 (I484974,I485181,I485452);
DFFARX1 I_28347 (I485421,I3563,I484997,I484986,);
DFFARX1 I_28348 (I485421,I3563,I484997,I484983,);
not I_28349 (I485541,I3570);
DFFARX1 I_28350 (I764768,I3563,I485541,I485567,);
DFFARX1 I_28351 (I485567,I3563,I485541,I485584,);
not I_28352 (I485533,I485584);
not I_28353 (I485606,I485567);
nand I_28354 (I485623,I764789,I764780);
and I_28355 (I485640,I485623,I764768);
DFFARX1 I_28356 (I485640,I3563,I485541,I485666,);
not I_28357 (I485674,I485666);
DFFARX1 I_28358 (I764774,I3563,I485541,I485700,);
and I_28359 (I485708,I485700,I764771);
nand I_28360 (I485725,I485700,I764771);
nand I_28361 (I485512,I485674,I485725);
DFFARX1 I_28362 (I764765,I3563,I485541,I485765,);
nor I_28363 (I485773,I485765,I485708);
DFFARX1 I_28364 (I485773,I3563,I485541,I485506,);
nor I_28365 (I485521,I485765,I485666);
nand I_28366 (I485818,I764765,I764777);
and I_28367 (I485835,I485818,I764786);
DFFARX1 I_28368 (I485835,I3563,I485541,I485861,);
nor I_28369 (I485509,I485861,I485765);
not I_28370 (I485883,I485861);
nor I_28371 (I485900,I485883,I485674);
nor I_28372 (I485917,I485606,I485900);
DFFARX1 I_28373 (I485917,I3563,I485541,I485524,);
nor I_28374 (I485948,I485883,I485765);
nor I_28375 (I485965,I764783,I764777);
nor I_28376 (I485515,I485965,I485948);
not I_28377 (I485996,I485965);
nand I_28378 (I485518,I485725,I485996);
DFFARX1 I_28379 (I485965,I3563,I485541,I485530,);
DFFARX1 I_28380 (I485965,I3563,I485541,I485527,);
not I_28381 (I486085,I3570);
DFFARX1 I_28382 (I746850,I3563,I486085,I486111,);
DFFARX1 I_28383 (I486111,I3563,I486085,I486128,);
not I_28384 (I486077,I486128);
not I_28385 (I486150,I486111);
nand I_28386 (I486167,I746871,I746862);
and I_28387 (I486184,I486167,I746850);
DFFARX1 I_28388 (I486184,I3563,I486085,I486210,);
not I_28389 (I486218,I486210);
DFFARX1 I_28390 (I746856,I3563,I486085,I486244,);
and I_28391 (I486252,I486244,I746853);
nand I_28392 (I486269,I486244,I746853);
nand I_28393 (I486056,I486218,I486269);
DFFARX1 I_28394 (I746847,I3563,I486085,I486309,);
nor I_28395 (I486317,I486309,I486252);
DFFARX1 I_28396 (I486317,I3563,I486085,I486050,);
nor I_28397 (I486065,I486309,I486210);
nand I_28398 (I486362,I746847,I746859);
and I_28399 (I486379,I486362,I746868);
DFFARX1 I_28400 (I486379,I3563,I486085,I486405,);
nor I_28401 (I486053,I486405,I486309);
not I_28402 (I486427,I486405);
nor I_28403 (I486444,I486427,I486218);
nor I_28404 (I486461,I486150,I486444);
DFFARX1 I_28405 (I486461,I3563,I486085,I486068,);
nor I_28406 (I486492,I486427,I486309);
nor I_28407 (I486509,I746865,I746859);
nor I_28408 (I486059,I486509,I486492);
not I_28409 (I486540,I486509);
nand I_28410 (I486062,I486269,I486540);
DFFARX1 I_28411 (I486509,I3563,I486085,I486074,);
DFFARX1 I_28412 (I486509,I3563,I486085,I486071,);
not I_28413 (I486629,I3570);
DFFARX1 I_28414 (I348099,I3563,I486629,I486655,);
DFFARX1 I_28415 (I486655,I3563,I486629,I486672,);
not I_28416 (I486621,I486672);
not I_28417 (I486694,I486655);
nand I_28418 (I486711,I348078,I348102);
and I_28419 (I486728,I486711,I348105);
DFFARX1 I_28420 (I486728,I3563,I486629,I486754,);
not I_28421 (I486762,I486754);
DFFARX1 I_28422 (I348087,I3563,I486629,I486788,);
and I_28423 (I486796,I486788,I348093);
nand I_28424 (I486813,I486788,I348093);
nand I_28425 (I486600,I486762,I486813);
DFFARX1 I_28426 (I348081,I3563,I486629,I486853,);
nor I_28427 (I486861,I486853,I486796);
DFFARX1 I_28428 (I486861,I3563,I486629,I486594,);
nor I_28429 (I486609,I486853,I486754);
nand I_28430 (I486906,I348090,I348078);
and I_28431 (I486923,I486906,I348084);
DFFARX1 I_28432 (I486923,I3563,I486629,I486949,);
nor I_28433 (I486597,I486949,I486853);
not I_28434 (I486971,I486949);
nor I_28435 (I486988,I486971,I486762);
nor I_28436 (I487005,I486694,I486988);
DFFARX1 I_28437 (I487005,I3563,I486629,I486612,);
nor I_28438 (I487036,I486971,I486853);
nor I_28439 (I487053,I348096,I348078);
nor I_28440 (I486603,I487053,I487036);
not I_28441 (I487084,I487053);
nand I_28442 (I486606,I486813,I487084);
DFFARX1 I_28443 (I487053,I3563,I486629,I486618,);
DFFARX1 I_28444 (I487053,I3563,I486629,I486615,);
not I_28445 (I487173,I3570);
DFFARX1 I_28446 (I261302,I3563,I487173,I487199,);
DFFARX1 I_28447 (I487199,I3563,I487173,I487216,);
not I_28448 (I487165,I487216);
not I_28449 (I487238,I487199);
nand I_28450 (I487255,I261314,I261293);
and I_28451 (I487272,I487255,I261296);
DFFARX1 I_28452 (I487272,I3563,I487173,I487298,);
not I_28453 (I487306,I487298);
DFFARX1 I_28454 (I261305,I3563,I487173,I487332,);
and I_28455 (I487340,I487332,I261317);
nand I_28456 (I487357,I487332,I261317);
nand I_28457 (I487144,I487306,I487357);
DFFARX1 I_28458 (I261311,I3563,I487173,I487397,);
nor I_28459 (I487405,I487397,I487340);
DFFARX1 I_28460 (I487405,I3563,I487173,I487138,);
nor I_28461 (I487153,I487397,I487298);
nand I_28462 (I487450,I261299,I261296);
and I_28463 (I487467,I487450,I261308);
DFFARX1 I_28464 (I487467,I3563,I487173,I487493,);
nor I_28465 (I487141,I487493,I487397);
not I_28466 (I487515,I487493);
nor I_28467 (I487532,I487515,I487306);
nor I_28468 (I487549,I487238,I487532);
DFFARX1 I_28469 (I487549,I3563,I487173,I487156,);
nor I_28470 (I487580,I487515,I487397);
nor I_28471 (I487597,I261293,I261296);
nor I_28472 (I487147,I487597,I487580);
not I_28473 (I487628,I487597);
nand I_28474 (I487150,I487357,I487628);
DFFARX1 I_28475 (I487597,I3563,I487173,I487162,);
DFFARX1 I_28476 (I487597,I3563,I487173,I487159,);
not I_28477 (I487717,I3570);
DFFARX1 I_28478 (I419244,I3563,I487717,I487743,);
DFFARX1 I_28479 (I487743,I3563,I487717,I487760,);
not I_28480 (I487709,I487760);
not I_28481 (I487782,I487743);
nand I_28482 (I487799,I419223,I419247);
and I_28483 (I487816,I487799,I419250);
DFFARX1 I_28484 (I487816,I3563,I487717,I487842,);
not I_28485 (I487850,I487842);
DFFARX1 I_28486 (I419232,I3563,I487717,I487876,);
and I_28487 (I487884,I487876,I419238);
nand I_28488 (I487901,I487876,I419238);
nand I_28489 (I487688,I487850,I487901);
DFFARX1 I_28490 (I419226,I3563,I487717,I487941,);
nor I_28491 (I487949,I487941,I487884);
DFFARX1 I_28492 (I487949,I3563,I487717,I487682,);
nor I_28493 (I487697,I487941,I487842);
nand I_28494 (I487994,I419235,I419223);
and I_28495 (I488011,I487994,I419229);
DFFARX1 I_28496 (I488011,I3563,I487717,I488037,);
nor I_28497 (I487685,I488037,I487941);
not I_28498 (I488059,I488037);
nor I_28499 (I488076,I488059,I487850);
nor I_28500 (I488093,I487782,I488076);
DFFARX1 I_28501 (I488093,I3563,I487717,I487700,);
nor I_28502 (I488124,I488059,I487941);
nor I_28503 (I488141,I419241,I419223);
nor I_28504 (I487691,I488141,I488124);
not I_28505 (I488172,I488141);
nand I_28506 (I487694,I487901,I488172);
DFFARX1 I_28507 (I488141,I3563,I487717,I487706,);
DFFARX1 I_28508 (I488141,I3563,I487717,I487703,);
not I_28509 (I488261,I3570);
DFFARX1 I_28510 (I547134,I3563,I488261,I488287,);
DFFARX1 I_28511 (I488287,I3563,I488261,I488304,);
not I_28512 (I488253,I488304);
not I_28513 (I488326,I488287);
nand I_28514 (I488343,I547137,I547155);
and I_28515 (I488360,I488343,I547143);
DFFARX1 I_28516 (I488360,I3563,I488261,I488386,);
not I_28517 (I488394,I488386);
DFFARX1 I_28518 (I547134,I3563,I488261,I488420,);
and I_28519 (I488428,I488420,I547152);
nand I_28520 (I488445,I488420,I547152);
nand I_28521 (I488232,I488394,I488445);
DFFARX1 I_28522 (I547146,I3563,I488261,I488485,);
nor I_28523 (I488493,I488485,I488428);
DFFARX1 I_28524 (I488493,I3563,I488261,I488226,);
nor I_28525 (I488241,I488485,I488386);
nand I_28526 (I488538,I547149,I547131);
and I_28527 (I488555,I488538,I547140);
DFFARX1 I_28528 (I488555,I3563,I488261,I488581,);
nor I_28529 (I488229,I488581,I488485);
not I_28530 (I488603,I488581);
nor I_28531 (I488620,I488603,I488394);
nor I_28532 (I488637,I488326,I488620);
DFFARX1 I_28533 (I488637,I3563,I488261,I488244,);
nor I_28534 (I488668,I488603,I488485);
nor I_28535 (I488685,I547131,I547131);
nor I_28536 (I488235,I488685,I488668);
not I_28537 (I488716,I488685);
nand I_28538 (I488238,I488445,I488716);
DFFARX1 I_28539 (I488685,I3563,I488261,I488250,);
DFFARX1 I_28540 (I488685,I3563,I488261,I488247,);
not I_28541 (I488805,I3570);
DFFARX1 I_28542 (I889064,I3563,I488805,I488831,);
DFFARX1 I_28543 (I488831,I3563,I488805,I488848,);
not I_28544 (I488797,I488848);
not I_28545 (I488870,I488831);
nand I_28546 (I488887,I889058,I889055);
and I_28547 (I488904,I488887,I889070);
DFFARX1 I_28548 (I488904,I3563,I488805,I488930,);
not I_28549 (I488938,I488930);
DFFARX1 I_28550 (I889058,I3563,I488805,I488964,);
and I_28551 (I488972,I488964,I889052);
nand I_28552 (I488989,I488964,I889052);
nand I_28553 (I488776,I488938,I488989);
DFFARX1 I_28554 (I889052,I3563,I488805,I489029,);
nor I_28555 (I489037,I489029,I488972);
DFFARX1 I_28556 (I489037,I3563,I488805,I488770,);
nor I_28557 (I488785,I489029,I488930);
nand I_28558 (I489082,I889067,I889061);
and I_28559 (I489099,I489082,I889055);
DFFARX1 I_28560 (I489099,I3563,I488805,I489125,);
nor I_28561 (I488773,I489125,I489029);
not I_28562 (I489147,I489125);
nor I_28563 (I489164,I489147,I488938);
nor I_28564 (I489181,I488870,I489164);
DFFARX1 I_28565 (I489181,I3563,I488805,I488788,);
nor I_28566 (I489212,I489147,I489029);
nor I_28567 (I489229,I889073,I889061);
nor I_28568 (I488779,I489229,I489212);
not I_28569 (I489260,I489229);
nand I_28570 (I488782,I488989,I489260);
DFFARX1 I_28571 (I489229,I3563,I488805,I488794,);
DFFARX1 I_28572 (I489229,I3563,I488805,I488791,);
not I_28573 (I489349,I3570);
DFFARX1 I_28574 (I813176,I3563,I489349,I489375,);
DFFARX1 I_28575 (I489375,I3563,I489349,I489392,);
not I_28576 (I489341,I489392);
not I_28577 (I489414,I489375);
nand I_28578 (I489431,I813170,I813167);
and I_28579 (I489448,I489431,I813182);
DFFARX1 I_28580 (I489448,I3563,I489349,I489474,);
not I_28581 (I489482,I489474);
DFFARX1 I_28582 (I813170,I3563,I489349,I489508,);
and I_28583 (I489516,I489508,I813164);
nand I_28584 (I489533,I489508,I813164);
nand I_28585 (I489320,I489482,I489533);
DFFARX1 I_28586 (I813164,I3563,I489349,I489573,);
nor I_28587 (I489581,I489573,I489516);
DFFARX1 I_28588 (I489581,I3563,I489349,I489314,);
nor I_28589 (I489329,I489573,I489474);
nand I_28590 (I489626,I813179,I813173);
and I_28591 (I489643,I489626,I813167);
DFFARX1 I_28592 (I489643,I3563,I489349,I489669,);
nor I_28593 (I489317,I489669,I489573);
not I_28594 (I489691,I489669);
nor I_28595 (I489708,I489691,I489482);
nor I_28596 (I489725,I489414,I489708);
DFFARX1 I_28597 (I489725,I3563,I489349,I489332,);
nor I_28598 (I489756,I489691,I489573);
nor I_28599 (I489773,I813185,I813173);
nor I_28600 (I489323,I489773,I489756);
not I_28601 (I489804,I489773);
nand I_28602 (I489326,I489533,I489804);
DFFARX1 I_28603 (I489773,I3563,I489349,I489338,);
DFFARX1 I_28604 (I489773,I3563,I489349,I489335,);
not I_28605 (I489893,I3570);
DFFARX1 I_28606 (I684426,I3563,I489893,I489919,);
DFFARX1 I_28607 (I489919,I3563,I489893,I489936,);
not I_28608 (I489885,I489936);
not I_28609 (I489958,I489919);
nand I_28610 (I489975,I684447,I684438);
and I_28611 (I489992,I489975,I684426);
DFFARX1 I_28612 (I489992,I3563,I489893,I490018,);
not I_28613 (I490026,I490018);
DFFARX1 I_28614 (I684432,I3563,I489893,I490052,);
and I_28615 (I490060,I490052,I684429);
nand I_28616 (I490077,I490052,I684429);
nand I_28617 (I489864,I490026,I490077);
DFFARX1 I_28618 (I684423,I3563,I489893,I490117,);
nor I_28619 (I490125,I490117,I490060);
DFFARX1 I_28620 (I490125,I3563,I489893,I489858,);
nor I_28621 (I489873,I490117,I490018);
nand I_28622 (I490170,I684423,I684435);
and I_28623 (I490187,I490170,I684444);
DFFARX1 I_28624 (I490187,I3563,I489893,I490213,);
nor I_28625 (I489861,I490213,I490117);
not I_28626 (I490235,I490213);
nor I_28627 (I490252,I490235,I490026);
nor I_28628 (I490269,I489958,I490252);
DFFARX1 I_28629 (I490269,I3563,I489893,I489876,);
nor I_28630 (I490300,I490235,I490117);
nor I_28631 (I490317,I684441,I684435);
nor I_28632 (I489867,I490317,I490300);
not I_28633 (I490348,I490317);
nand I_28634 (I489870,I490077,I490348);
DFFARX1 I_28635 (I490317,I3563,I489893,I489882,);
DFFARX1 I_28636 (I490317,I3563,I489893,I489879,);
not I_28637 (I490437,I3570);
DFFARX1 I_28638 (I1091576,I3563,I490437,I490463,);
DFFARX1 I_28639 (I490463,I3563,I490437,I490480,);
not I_28640 (I490429,I490480);
not I_28641 (I490502,I490463);
nand I_28642 (I490519,I1091588,I1091576);
and I_28643 (I490536,I490519,I1091579);
DFFARX1 I_28644 (I490536,I3563,I490437,I490562,);
not I_28645 (I490570,I490562);
DFFARX1 I_28646 (I1091597,I3563,I490437,I490596,);
and I_28647 (I490604,I490596,I1091573);
nand I_28648 (I490621,I490596,I1091573);
nand I_28649 (I490408,I490570,I490621);
DFFARX1 I_28650 (I1091591,I3563,I490437,I490661,);
nor I_28651 (I490669,I490661,I490604);
DFFARX1 I_28652 (I490669,I3563,I490437,I490402,);
nor I_28653 (I490417,I490661,I490562);
nand I_28654 (I490714,I1091585,I1091582);
and I_28655 (I490731,I490714,I1091594);
DFFARX1 I_28656 (I490731,I3563,I490437,I490757,);
nor I_28657 (I490405,I490757,I490661);
not I_28658 (I490779,I490757);
nor I_28659 (I490796,I490779,I490570);
nor I_28660 (I490813,I490502,I490796);
DFFARX1 I_28661 (I490813,I3563,I490437,I490420,);
nor I_28662 (I490844,I490779,I490661);
nor I_28663 (I490861,I1091573,I1091582);
nor I_28664 (I490411,I490861,I490844);
not I_28665 (I490892,I490861);
nand I_28666 (I490414,I490621,I490892);
DFFARX1 I_28667 (I490861,I3563,I490437,I490426,);
DFFARX1 I_28668 (I490861,I3563,I490437,I490423,);
not I_28669 (I490981,I3570);
DFFARX1 I_28670 (I3591,I3563,I490981,I491007,);
DFFARX1 I_28671 (I491007,I3563,I490981,I491024,);
not I_28672 (I490973,I491024);
not I_28673 (I491046,I491007);
nand I_28674 (I491063,I3594,I3582);
and I_28675 (I491080,I491063,I3588);
DFFARX1 I_28676 (I491080,I3563,I490981,I491106,);
not I_28677 (I491114,I491106);
DFFARX1 I_28678 (I3576,I3563,I490981,I491140,);
and I_28679 (I491148,I491140,I3573);
nand I_28680 (I491165,I491140,I3573);
nand I_28681 (I490952,I491114,I491165);
DFFARX1 I_28682 (I3579,I3563,I490981,I491205,);
nor I_28683 (I491213,I491205,I491148);
DFFARX1 I_28684 (I491213,I3563,I490981,I490946,);
nor I_28685 (I490961,I491205,I491106);
nand I_28686 (I491258,I3579,I3576);
and I_28687 (I491275,I491258,I3573);
DFFARX1 I_28688 (I491275,I3563,I490981,I491301,);
nor I_28689 (I490949,I491301,I491205);
not I_28690 (I491323,I491301);
nor I_28691 (I491340,I491323,I491114);
nor I_28692 (I491357,I491046,I491340);
DFFARX1 I_28693 (I491357,I3563,I490981,I490964,);
nor I_28694 (I491388,I491323,I491205);
nor I_28695 (I491405,I3585,I3576);
nor I_28696 (I490955,I491405,I491388);
not I_28697 (I491436,I491405);
nand I_28698 (I490958,I491165,I491436);
DFFARX1 I_28699 (I491405,I3563,I490981,I490970,);
DFFARX1 I_28700 (I491405,I3563,I490981,I490967,);
not I_28701 (I491525,I3570);
DFFARX1 I_28702 (I1298175,I3563,I491525,I491551,);
DFFARX1 I_28703 (I491551,I3563,I491525,I491568,);
not I_28704 (I491517,I491568);
not I_28705 (I491590,I491551);
nand I_28706 (I491607,I1298172,I1298169);
and I_28707 (I491624,I491607,I1298157);
DFFARX1 I_28708 (I491624,I3563,I491525,I491650,);
not I_28709 (I491658,I491650);
DFFARX1 I_28710 (I1298181,I3563,I491525,I491684,);
and I_28711 (I491692,I491684,I1298166);
nand I_28712 (I491709,I491684,I1298166);
nand I_28713 (I491496,I491658,I491709);
DFFARX1 I_28714 (I1298160,I3563,I491525,I491749,);
nor I_28715 (I491757,I491749,I491692);
DFFARX1 I_28716 (I491757,I3563,I491525,I491490,);
nor I_28717 (I491505,I491749,I491650);
nand I_28718 (I491802,I1298157,I1298163);
and I_28719 (I491819,I491802,I1298178);
DFFARX1 I_28720 (I491819,I3563,I491525,I491845,);
nor I_28721 (I491493,I491845,I491749);
not I_28722 (I491867,I491845);
nor I_28723 (I491884,I491867,I491658);
nor I_28724 (I491901,I491590,I491884);
DFFARX1 I_28725 (I491901,I3563,I491525,I491508,);
nor I_28726 (I491932,I491867,I491749);
nor I_28727 (I491949,I1298160,I1298163);
nor I_28728 (I491499,I491949,I491932);
not I_28729 (I491980,I491949);
nand I_28730 (I491502,I491709,I491980);
DFFARX1 I_28731 (I491949,I3563,I491525,I491514,);
DFFARX1 I_28732 (I491949,I3563,I491525,I491511,);
not I_28733 (I492069,I3570);
DFFARX1 I_28734 (I1352975,I3563,I492069,I492095,);
DFFARX1 I_28735 (I492095,I3563,I492069,I492112,);
not I_28736 (I492061,I492112);
not I_28737 (I492134,I492095);
nand I_28738 (I492151,I1352951,I1352972);
and I_28739 (I492168,I492151,I1352969);
DFFARX1 I_28740 (I492168,I3563,I492069,I492194,);
not I_28741 (I492202,I492194);
DFFARX1 I_28742 (I1352948,I3563,I492069,I492228,);
and I_28743 (I492236,I492228,I1352960);
nand I_28744 (I492253,I492228,I1352960);
nand I_28745 (I492040,I492202,I492253);
DFFARX1 I_28746 (I1352963,I3563,I492069,I492293,);
nor I_28747 (I492301,I492293,I492236);
DFFARX1 I_28748 (I492301,I3563,I492069,I492034,);
nor I_28749 (I492049,I492293,I492194);
nand I_28750 (I492346,I1352966,I1352954);
and I_28751 (I492363,I492346,I1352957);
DFFARX1 I_28752 (I492363,I3563,I492069,I492389,);
nor I_28753 (I492037,I492389,I492293);
not I_28754 (I492411,I492389);
nor I_28755 (I492428,I492411,I492202);
nor I_28756 (I492445,I492134,I492428);
DFFARX1 I_28757 (I492445,I3563,I492069,I492052,);
nor I_28758 (I492476,I492411,I492293);
nor I_28759 (I492493,I1352948,I1352954);
nor I_28760 (I492043,I492493,I492476);
not I_28761 (I492524,I492493);
nand I_28762 (I492046,I492253,I492524);
DFFARX1 I_28763 (I492493,I3563,I492069,I492058,);
DFFARX1 I_28764 (I492493,I3563,I492069,I492055,);
not I_28765 (I492613,I3570);
DFFARX1 I_28766 (I1237810,I3563,I492613,I492639,);
DFFARX1 I_28767 (I492639,I3563,I492613,I492656,);
not I_28768 (I492605,I492656);
not I_28769 (I492678,I492639);
nand I_28770 (I492695,I1237822,I1237810);
and I_28771 (I492712,I492695,I1237813);
DFFARX1 I_28772 (I492712,I3563,I492613,I492738,);
not I_28773 (I492746,I492738);
DFFARX1 I_28774 (I1237831,I3563,I492613,I492772,);
and I_28775 (I492780,I492772,I1237807);
nand I_28776 (I492797,I492772,I1237807);
nand I_28777 (I492584,I492746,I492797);
DFFARX1 I_28778 (I1237825,I3563,I492613,I492837,);
nor I_28779 (I492845,I492837,I492780);
DFFARX1 I_28780 (I492845,I3563,I492613,I492578,);
nor I_28781 (I492593,I492837,I492738);
nand I_28782 (I492890,I1237819,I1237816);
and I_28783 (I492907,I492890,I1237828);
DFFARX1 I_28784 (I492907,I3563,I492613,I492933,);
nor I_28785 (I492581,I492933,I492837);
not I_28786 (I492955,I492933);
nor I_28787 (I492972,I492955,I492746);
nor I_28788 (I492989,I492678,I492972);
DFFARX1 I_28789 (I492989,I3563,I492613,I492596,);
nor I_28790 (I493020,I492955,I492837);
nor I_28791 (I493037,I1237807,I1237816);
nor I_28792 (I492587,I493037,I493020);
not I_28793 (I493068,I493037);
nand I_28794 (I492590,I492797,I493068);
DFFARX1 I_28795 (I493037,I3563,I492613,I492602,);
DFFARX1 I_28796 (I493037,I3563,I492613,I492599,);
not I_28797 (I493157,I3570);
DFFARX1 I_28798 (I304885,I3563,I493157,I493183,);
DFFARX1 I_28799 (I493183,I3563,I493157,I493200,);
not I_28800 (I493149,I493200);
not I_28801 (I493222,I493183);
nand I_28802 (I493239,I304864,I304888);
and I_28803 (I493256,I493239,I304891);
DFFARX1 I_28804 (I493256,I3563,I493157,I493282,);
not I_28805 (I493290,I493282);
DFFARX1 I_28806 (I304873,I3563,I493157,I493316,);
and I_28807 (I493324,I493316,I304879);
nand I_28808 (I493341,I493316,I304879);
nand I_28809 (I493128,I493290,I493341);
DFFARX1 I_28810 (I304867,I3563,I493157,I493381,);
nor I_28811 (I493389,I493381,I493324);
DFFARX1 I_28812 (I493389,I3563,I493157,I493122,);
nor I_28813 (I493137,I493381,I493282);
nand I_28814 (I493434,I304876,I304864);
and I_28815 (I493451,I493434,I304870);
DFFARX1 I_28816 (I493451,I3563,I493157,I493477,);
nor I_28817 (I493125,I493477,I493381);
not I_28818 (I493499,I493477);
nor I_28819 (I493516,I493499,I493290);
nor I_28820 (I493533,I493222,I493516);
DFFARX1 I_28821 (I493533,I3563,I493157,I493140,);
nor I_28822 (I493564,I493499,I493381);
nor I_28823 (I493581,I304882,I304864);
nor I_28824 (I493131,I493581,I493564);
not I_28825 (I493612,I493581);
nand I_28826 (I493134,I493341,I493612);
DFFARX1 I_28827 (I493581,I3563,I493157,I493146,);
DFFARX1 I_28828 (I493581,I3563,I493157,I493143,);
not I_28829 (I493701,I3570);
DFFARX1 I_28830 (I704656,I3563,I493701,I493727,);
DFFARX1 I_28831 (I493727,I3563,I493701,I493744,);
not I_28832 (I493693,I493744);
not I_28833 (I493766,I493727);
nand I_28834 (I493783,I704677,I704668);
and I_28835 (I493800,I493783,I704656);
DFFARX1 I_28836 (I493800,I3563,I493701,I493826,);
not I_28837 (I493834,I493826);
DFFARX1 I_28838 (I704662,I3563,I493701,I493860,);
and I_28839 (I493868,I493860,I704659);
nand I_28840 (I493885,I493860,I704659);
nand I_28841 (I493672,I493834,I493885);
DFFARX1 I_28842 (I704653,I3563,I493701,I493925,);
nor I_28843 (I493933,I493925,I493868);
DFFARX1 I_28844 (I493933,I3563,I493701,I493666,);
nor I_28845 (I493681,I493925,I493826);
nand I_28846 (I493978,I704653,I704665);
and I_28847 (I493995,I493978,I704674);
DFFARX1 I_28848 (I493995,I3563,I493701,I494021,);
nor I_28849 (I493669,I494021,I493925);
not I_28850 (I494043,I494021);
nor I_28851 (I494060,I494043,I493834);
nor I_28852 (I494077,I493766,I494060);
DFFARX1 I_28853 (I494077,I3563,I493701,I493684,);
nor I_28854 (I494108,I494043,I493925);
nor I_28855 (I494125,I704671,I704665);
nor I_28856 (I493675,I494125,I494108);
not I_28857 (I494156,I494125);
nand I_28858 (I493678,I493885,I494156);
DFFARX1 I_28859 (I494125,I3563,I493701,I493690,);
DFFARX1 I_28860 (I494125,I3563,I493701,I493687,);
not I_28861 (I494245,I3570);
DFFARX1 I_28862 (I652636,I3563,I494245,I494271,);
DFFARX1 I_28863 (I494271,I3563,I494245,I494288,);
not I_28864 (I494237,I494288);
not I_28865 (I494310,I494271);
nand I_28866 (I494327,I652633,I652654);
and I_28867 (I494344,I494327,I652657);
DFFARX1 I_28868 (I494344,I3563,I494245,I494370,);
not I_28869 (I494378,I494370);
DFFARX1 I_28870 (I652642,I3563,I494245,I494404,);
and I_28871 (I494412,I494404,I652645);
nand I_28872 (I494429,I494404,I652645);
nand I_28873 (I494216,I494378,I494429);
DFFARX1 I_28874 (I652648,I3563,I494245,I494469,);
nor I_28875 (I494477,I494469,I494412);
DFFARX1 I_28876 (I494477,I3563,I494245,I494210,);
nor I_28877 (I494225,I494469,I494370);
nand I_28878 (I494522,I652633,I652639);
and I_28879 (I494539,I494522,I652651);
DFFARX1 I_28880 (I494539,I3563,I494245,I494565,);
nor I_28881 (I494213,I494565,I494469);
not I_28882 (I494587,I494565);
nor I_28883 (I494604,I494587,I494378);
nor I_28884 (I494621,I494310,I494604);
DFFARX1 I_28885 (I494621,I3563,I494245,I494228,);
nor I_28886 (I494652,I494587,I494469);
nor I_28887 (I494669,I652636,I652639);
nor I_28888 (I494219,I494669,I494652);
not I_28889 (I494700,I494669);
nand I_28890 (I494222,I494429,I494700);
DFFARX1 I_28891 (I494669,I3563,I494245,I494234,);
DFFARX1 I_28892 (I494669,I3563,I494245,I494231,);
not I_28893 (I494789,I3570);
DFFARX1 I_28894 (I1025347,I3563,I494789,I494815,);
DFFARX1 I_28895 (I494815,I3563,I494789,I494832,);
not I_28896 (I494781,I494832);
not I_28897 (I494854,I494815);
nand I_28898 (I494871,I1025362,I1025350);
and I_28899 (I494888,I494871,I1025341);
DFFARX1 I_28900 (I494888,I3563,I494789,I494914,);
not I_28901 (I494922,I494914);
DFFARX1 I_28902 (I1025353,I3563,I494789,I494948,);
and I_28903 (I494956,I494948,I1025344);
nand I_28904 (I494973,I494948,I1025344);
nand I_28905 (I494760,I494922,I494973);
DFFARX1 I_28906 (I1025359,I3563,I494789,I495013,);
nor I_28907 (I495021,I495013,I494956);
DFFARX1 I_28908 (I495021,I3563,I494789,I494754,);
nor I_28909 (I494769,I495013,I494914);
nand I_28910 (I495066,I1025368,I1025356);
and I_28911 (I495083,I495066,I1025365);
DFFARX1 I_28912 (I495083,I3563,I494789,I495109,);
nor I_28913 (I494757,I495109,I495013);
not I_28914 (I495131,I495109);
nor I_28915 (I495148,I495131,I494922);
nor I_28916 (I495165,I494854,I495148);
DFFARX1 I_28917 (I495165,I3563,I494789,I494772,);
nor I_28918 (I495196,I495131,I495013);
nor I_28919 (I495213,I1025341,I1025356);
nor I_28920 (I494763,I495213,I495196);
not I_28921 (I495244,I495213);
nand I_28922 (I494766,I494973,I495244);
DFFARX1 I_28923 (I495213,I3563,I494789,I494778,);
DFFARX1 I_28924 (I495213,I3563,I494789,I494775,);
not I_28925 (I495333,I3570);
DFFARX1 I_28926 (I47173,I3563,I495333,I495359,);
DFFARX1 I_28927 (I495359,I3563,I495333,I495376,);
not I_28928 (I495325,I495376);
not I_28929 (I495398,I495359);
nand I_28930 (I495415,I47161,I47176);
and I_28931 (I495432,I495415,I47164);
DFFARX1 I_28932 (I495432,I3563,I495333,I495458,);
not I_28933 (I495466,I495458);
DFFARX1 I_28934 (I47185,I3563,I495333,I495492,);
and I_28935 (I495500,I495492,I47179);
nand I_28936 (I495517,I495492,I47179);
nand I_28937 (I495304,I495466,I495517);
DFFARX1 I_28938 (I47182,I3563,I495333,I495557,);
nor I_28939 (I495565,I495557,I495500);
DFFARX1 I_28940 (I495565,I3563,I495333,I495298,);
nor I_28941 (I495313,I495557,I495458);
nand I_28942 (I495610,I47161,I47164);
and I_28943 (I495627,I495610,I47167);
DFFARX1 I_28944 (I495627,I3563,I495333,I495653,);
nor I_28945 (I495301,I495653,I495557);
not I_28946 (I495675,I495653);
nor I_28947 (I495692,I495675,I495466);
nor I_28948 (I495709,I495398,I495692);
DFFARX1 I_28949 (I495709,I3563,I495333,I495316,);
nor I_28950 (I495740,I495675,I495557);
nor I_28951 (I495757,I47170,I47164);
nor I_28952 (I495307,I495757,I495740);
not I_28953 (I495788,I495757);
nand I_28954 (I495310,I495517,I495788);
DFFARX1 I_28955 (I495757,I3563,I495333,I495322,);
DFFARX1 I_28956 (I495757,I3563,I495333,I495319,);
not I_28957 (I495877,I3570);
DFFARX1 I_28958 (I164320,I3563,I495877,I495903,);
DFFARX1 I_28959 (I495903,I3563,I495877,I495920,);
not I_28960 (I495869,I495920);
not I_28961 (I495942,I495903);
nand I_28962 (I495959,I164329,I164332);
and I_28963 (I495976,I495959,I164311);
DFFARX1 I_28964 (I495976,I3563,I495877,I496002,);
not I_28965 (I496010,I496002);
DFFARX1 I_28966 (I164326,I3563,I495877,I496036,);
and I_28967 (I496044,I496036,I164314);
nand I_28968 (I496061,I496036,I164314);
nand I_28969 (I495848,I496010,I496061);
DFFARX1 I_28970 (I164308,I3563,I495877,I496101,);
nor I_28971 (I496109,I496101,I496044);
DFFARX1 I_28972 (I496109,I3563,I495877,I495842,);
nor I_28973 (I495857,I496101,I496002);
nand I_28974 (I496154,I164323,I164317);
and I_28975 (I496171,I496154,I164308);
DFFARX1 I_28976 (I496171,I3563,I495877,I496197,);
nor I_28977 (I495845,I496197,I496101);
not I_28978 (I496219,I496197);
nor I_28979 (I496236,I496219,I496010);
nor I_28980 (I496253,I495942,I496236);
DFFARX1 I_28981 (I496253,I3563,I495877,I495860,);
nor I_28982 (I496284,I496219,I496101);
nor I_28983 (I496301,I164335,I164317);
nor I_28984 (I495851,I496301,I496284);
not I_28985 (I496332,I496301);
nand I_28986 (I495854,I496061,I496332);
DFFARX1 I_28987 (I496301,I3563,I495877,I495866,);
DFFARX1 I_28988 (I496301,I3563,I495877,I495863,);
not I_28989 (I496421,I3570);
DFFARX1 I_28990 (I886956,I3563,I496421,I496447,);
DFFARX1 I_28991 (I496447,I3563,I496421,I496464,);
not I_28992 (I496413,I496464);
not I_28993 (I496486,I496447);
nand I_28994 (I496503,I886950,I886947);
and I_28995 (I496520,I496503,I886962);
DFFARX1 I_28996 (I496520,I3563,I496421,I496546,);
not I_28997 (I496554,I496546);
DFFARX1 I_28998 (I886950,I3563,I496421,I496580,);
and I_28999 (I496588,I496580,I886944);
nand I_29000 (I496605,I496580,I886944);
nand I_29001 (I496392,I496554,I496605);
DFFARX1 I_29002 (I886944,I3563,I496421,I496645,);
nor I_29003 (I496653,I496645,I496588);
DFFARX1 I_29004 (I496653,I3563,I496421,I496386,);
nor I_29005 (I496401,I496645,I496546);
nand I_29006 (I496698,I886959,I886953);
and I_29007 (I496715,I496698,I886947);
DFFARX1 I_29008 (I496715,I3563,I496421,I496741,);
nor I_29009 (I496389,I496741,I496645);
not I_29010 (I496763,I496741);
nor I_29011 (I496780,I496763,I496554);
nor I_29012 (I496797,I496486,I496780);
DFFARX1 I_29013 (I496797,I3563,I496421,I496404,);
nor I_29014 (I496828,I496763,I496645);
nor I_29015 (I496845,I886965,I886953);
nor I_29016 (I496395,I496845,I496828);
not I_29017 (I496876,I496845);
nand I_29018 (I496398,I496605,I496876);
DFFARX1 I_29019 (I496845,I3563,I496421,I496410,);
DFFARX1 I_29020 (I496845,I3563,I496421,I496407,);
not I_29021 (I496965,I3570);
DFFARX1 I_29022 (I1078075,I3563,I496965,I496991,);
DFFARX1 I_29023 (I496991,I3563,I496965,I497008,);
not I_29024 (I496957,I497008);
not I_29025 (I497030,I496991);
nand I_29026 (I497047,I1078075,I1078093);
and I_29027 (I497064,I497047,I1078087);
DFFARX1 I_29028 (I497064,I3563,I496965,I497090,);
not I_29029 (I497098,I497090);
DFFARX1 I_29030 (I1078081,I3563,I496965,I497124,);
and I_29031 (I497132,I497124,I1078090);
nand I_29032 (I497149,I497124,I1078090);
nand I_29033 (I496936,I497098,I497149);
DFFARX1 I_29034 (I1078078,I3563,I496965,I497189,);
nor I_29035 (I497197,I497189,I497132);
DFFARX1 I_29036 (I497197,I3563,I496965,I496930,);
nor I_29037 (I496945,I497189,I497090);
nand I_29038 (I497242,I1078078,I1078096);
and I_29039 (I497259,I497242,I1078081);
DFFARX1 I_29040 (I497259,I3563,I496965,I497285,);
nor I_29041 (I496933,I497285,I497189);
not I_29042 (I497307,I497285);
nor I_29043 (I497324,I497307,I497098);
nor I_29044 (I497341,I497030,I497324);
DFFARX1 I_29045 (I497341,I3563,I496965,I496948,);
nor I_29046 (I497372,I497307,I497189);
nor I_29047 (I497389,I1078084,I1078096);
nor I_29048 (I496939,I497389,I497372);
not I_29049 (I497420,I497389);
nand I_29050 (I496942,I497149,I497420);
DFFARX1 I_29051 (I497389,I3563,I496965,I496954,);
DFFARX1 I_29052 (I497389,I3563,I496965,I496951,);
not I_29053 (I497509,I3570);
DFFARX1 I_29054 (I1333935,I3563,I497509,I497535,);
DFFARX1 I_29055 (I497535,I3563,I497509,I497552,);
not I_29056 (I497501,I497552);
not I_29057 (I497574,I497535);
nand I_29058 (I497591,I1333911,I1333932);
and I_29059 (I497608,I497591,I1333929);
DFFARX1 I_29060 (I497608,I3563,I497509,I497634,);
not I_29061 (I497642,I497634);
DFFARX1 I_29062 (I1333908,I3563,I497509,I497668,);
and I_29063 (I497676,I497668,I1333920);
nand I_29064 (I497693,I497668,I1333920);
nand I_29065 (I497480,I497642,I497693);
DFFARX1 I_29066 (I1333923,I3563,I497509,I497733,);
nor I_29067 (I497741,I497733,I497676);
DFFARX1 I_29068 (I497741,I3563,I497509,I497474,);
nor I_29069 (I497489,I497733,I497634);
nand I_29070 (I497786,I1333926,I1333914);
and I_29071 (I497803,I497786,I1333917);
DFFARX1 I_29072 (I497803,I3563,I497509,I497829,);
nor I_29073 (I497477,I497829,I497733);
not I_29074 (I497851,I497829);
nor I_29075 (I497868,I497851,I497642);
nor I_29076 (I497885,I497574,I497868);
DFFARX1 I_29077 (I497885,I3563,I497509,I497492,);
nor I_29078 (I497916,I497851,I497733);
nor I_29079 (I497933,I1333908,I1333914);
nor I_29080 (I497483,I497933,I497916);
not I_29081 (I497964,I497933);
nand I_29082 (I497486,I497693,I497964);
DFFARX1 I_29083 (I497933,I3563,I497509,I497498,);
DFFARX1 I_29084 (I497933,I3563,I497509,I497495,);
not I_29085 (I498053,I3570);
DFFARX1 I_29086 (I57713,I3563,I498053,I498079,);
DFFARX1 I_29087 (I498079,I3563,I498053,I498096,);
not I_29088 (I498045,I498096);
not I_29089 (I498118,I498079);
nand I_29090 (I498135,I57701,I57716);
and I_29091 (I498152,I498135,I57704);
DFFARX1 I_29092 (I498152,I3563,I498053,I498178,);
not I_29093 (I498186,I498178);
DFFARX1 I_29094 (I57725,I3563,I498053,I498212,);
and I_29095 (I498220,I498212,I57719);
nand I_29096 (I498237,I498212,I57719);
nand I_29097 (I498024,I498186,I498237);
DFFARX1 I_29098 (I57722,I3563,I498053,I498277,);
nor I_29099 (I498285,I498277,I498220);
DFFARX1 I_29100 (I498285,I3563,I498053,I498018,);
nor I_29101 (I498033,I498277,I498178);
nand I_29102 (I498330,I57701,I57704);
and I_29103 (I498347,I498330,I57707);
DFFARX1 I_29104 (I498347,I3563,I498053,I498373,);
nor I_29105 (I498021,I498373,I498277);
not I_29106 (I498395,I498373);
nor I_29107 (I498412,I498395,I498186);
nor I_29108 (I498429,I498118,I498412);
DFFARX1 I_29109 (I498429,I3563,I498053,I498036,);
nor I_29110 (I498460,I498395,I498277);
nor I_29111 (I498477,I57710,I57704);
nor I_29112 (I498027,I498477,I498460);
not I_29113 (I498508,I498477);
nand I_29114 (I498030,I498237,I498508);
DFFARX1 I_29115 (I498477,I3563,I498053,I498042,);
DFFARX1 I_29116 (I498477,I3563,I498053,I498039,);
not I_29117 (I498597,I3570);
DFFARX1 I_29118 (I323857,I3563,I498597,I498623,);
DFFARX1 I_29119 (I498623,I3563,I498597,I498640,);
not I_29120 (I498589,I498640);
not I_29121 (I498662,I498623);
nand I_29122 (I498679,I323836,I323860);
and I_29123 (I498696,I498679,I323863);
DFFARX1 I_29124 (I498696,I3563,I498597,I498722,);
not I_29125 (I498730,I498722);
DFFARX1 I_29126 (I323845,I3563,I498597,I498756,);
and I_29127 (I498764,I498756,I323851);
nand I_29128 (I498781,I498756,I323851);
nand I_29129 (I498568,I498730,I498781);
DFFARX1 I_29130 (I323839,I3563,I498597,I498821,);
nor I_29131 (I498829,I498821,I498764);
DFFARX1 I_29132 (I498829,I3563,I498597,I498562,);
nor I_29133 (I498577,I498821,I498722);
nand I_29134 (I498874,I323848,I323836);
and I_29135 (I498891,I498874,I323842);
DFFARX1 I_29136 (I498891,I3563,I498597,I498917,);
nor I_29137 (I498565,I498917,I498821);
not I_29138 (I498939,I498917);
nor I_29139 (I498956,I498939,I498730);
nor I_29140 (I498973,I498662,I498956);
DFFARX1 I_29141 (I498973,I3563,I498597,I498580,);
nor I_29142 (I499004,I498939,I498821);
nor I_29143 (I499021,I323854,I323836);
nor I_29144 (I498571,I499021,I499004);
not I_29145 (I499052,I499021);
nand I_29146 (I498574,I498781,I499052);
DFFARX1 I_29147 (I499021,I3563,I498597,I498586,);
DFFARX1 I_29148 (I499021,I3563,I498597,I498583,);
not I_29149 (I499141,I3570);
DFFARX1 I_29150 (I926509,I3563,I499141,I499167,);
DFFARX1 I_29151 (I499167,I3563,I499141,I499184,);
not I_29152 (I499133,I499184);
not I_29153 (I499206,I499167);
nand I_29154 (I499223,I926524,I926512);
and I_29155 (I499240,I499223,I926503);
DFFARX1 I_29156 (I499240,I3563,I499141,I499266,);
not I_29157 (I499274,I499266);
DFFARX1 I_29158 (I926515,I3563,I499141,I499300,);
and I_29159 (I499308,I499300,I926506);
nand I_29160 (I499325,I499300,I926506);
nand I_29161 (I499112,I499274,I499325);
DFFARX1 I_29162 (I926521,I3563,I499141,I499365,);
nor I_29163 (I499373,I499365,I499308);
DFFARX1 I_29164 (I499373,I3563,I499141,I499106,);
nor I_29165 (I499121,I499365,I499266);
nand I_29166 (I499418,I926530,I926518);
and I_29167 (I499435,I499418,I926527);
DFFARX1 I_29168 (I499435,I3563,I499141,I499461,);
nor I_29169 (I499109,I499461,I499365);
not I_29170 (I499483,I499461);
nor I_29171 (I499500,I499483,I499274);
nor I_29172 (I499517,I499206,I499500);
DFFARX1 I_29173 (I499517,I3563,I499141,I499124,);
nor I_29174 (I499548,I499483,I499365);
nor I_29175 (I499565,I926503,I926518);
nor I_29176 (I499115,I499565,I499548);
not I_29177 (I499596,I499565);
nand I_29178 (I499118,I499325,I499596);
DFFARX1 I_29179 (I499565,I3563,I499141,I499130,);
DFFARX1 I_29180 (I499565,I3563,I499141,I499127,);
not I_29181 (I499685,I3570);
DFFARX1 I_29182 (I550109,I3563,I499685,I499711,);
DFFARX1 I_29183 (I499711,I3563,I499685,I499728,);
not I_29184 (I499677,I499728);
not I_29185 (I499750,I499711);
nand I_29186 (I499767,I550112,I550130);
and I_29187 (I499784,I499767,I550118);
DFFARX1 I_29188 (I499784,I3563,I499685,I499810,);
not I_29189 (I499818,I499810);
DFFARX1 I_29190 (I550109,I3563,I499685,I499844,);
and I_29191 (I499852,I499844,I550127);
nand I_29192 (I499869,I499844,I550127);
nand I_29193 (I499656,I499818,I499869);
DFFARX1 I_29194 (I550121,I3563,I499685,I499909,);
nor I_29195 (I499917,I499909,I499852);
DFFARX1 I_29196 (I499917,I3563,I499685,I499650,);
nor I_29197 (I499665,I499909,I499810);
nand I_29198 (I499962,I550124,I550106);
and I_29199 (I499979,I499962,I550115);
DFFARX1 I_29200 (I499979,I3563,I499685,I500005,);
nor I_29201 (I499653,I500005,I499909);
not I_29202 (I500027,I500005);
nor I_29203 (I500044,I500027,I499818);
nor I_29204 (I500061,I499750,I500044);
DFFARX1 I_29205 (I500061,I3563,I499685,I499668,);
nor I_29206 (I500092,I500027,I499909);
nor I_29207 (I500109,I550106,I550106);
nor I_29208 (I499659,I500109,I500092);
not I_29209 (I500140,I500109);
nand I_29210 (I499662,I499869,I500140);
DFFARX1 I_29211 (I500109,I3563,I499685,I499674,);
DFFARX1 I_29212 (I500109,I3563,I499685,I499671,);
not I_29213 (I500229,I3570);
DFFARX1 I_29214 (I143081,I3563,I500229,I500255,);
DFFARX1 I_29215 (I500255,I3563,I500229,I500272,);
not I_29216 (I500221,I500272);
not I_29217 (I500294,I500255);
nand I_29218 (I500311,I143096,I143075);
and I_29219 (I500328,I500311,I143078);
DFFARX1 I_29220 (I500328,I3563,I500229,I500354,);
not I_29221 (I500362,I500354);
DFFARX1 I_29222 (I143084,I3563,I500229,I500388,);
and I_29223 (I500396,I500388,I143078);
nand I_29224 (I500413,I500388,I143078);
nand I_29225 (I500200,I500362,I500413);
DFFARX1 I_29226 (I143093,I3563,I500229,I500453,);
nor I_29227 (I500461,I500453,I500396);
DFFARX1 I_29228 (I500461,I3563,I500229,I500194,);
nor I_29229 (I500209,I500453,I500354);
nand I_29230 (I500506,I143075,I143090);
and I_29231 (I500523,I500506,I143087);
DFFARX1 I_29232 (I500523,I3563,I500229,I500549,);
nor I_29233 (I500197,I500549,I500453);
not I_29234 (I500571,I500549);
nor I_29235 (I500588,I500571,I500362);
nor I_29236 (I500605,I500294,I500588);
DFFARX1 I_29237 (I500605,I3563,I500229,I500212,);
nor I_29238 (I500636,I500571,I500453);
nor I_29239 (I500653,I143099,I143090);
nor I_29240 (I500203,I500653,I500636);
not I_29241 (I500684,I500653);
nand I_29242 (I500206,I500413,I500684);
DFFARX1 I_29243 (I500653,I3563,I500229,I500218,);
DFFARX1 I_29244 (I500653,I3563,I500229,I500215,);
not I_29245 (I500773,I3570);
DFFARX1 I_29246 (I81949,I3563,I500773,I500799,);
DFFARX1 I_29247 (I500799,I3563,I500773,I500816,);
not I_29248 (I500765,I500816);
not I_29249 (I500838,I500799);
nand I_29250 (I500855,I81964,I81943);
and I_29251 (I500872,I500855,I81946);
DFFARX1 I_29252 (I500872,I3563,I500773,I500898,);
not I_29253 (I500906,I500898);
DFFARX1 I_29254 (I81952,I3563,I500773,I500932,);
and I_29255 (I500940,I500932,I81946);
nand I_29256 (I500957,I500932,I81946);
nand I_29257 (I500744,I500906,I500957);
DFFARX1 I_29258 (I81961,I3563,I500773,I500997,);
nor I_29259 (I501005,I500997,I500940);
DFFARX1 I_29260 (I501005,I3563,I500773,I500738,);
nor I_29261 (I500753,I500997,I500898);
nand I_29262 (I501050,I81943,I81958);
and I_29263 (I501067,I501050,I81955);
DFFARX1 I_29264 (I501067,I3563,I500773,I501093,);
nor I_29265 (I500741,I501093,I500997);
not I_29266 (I501115,I501093);
nor I_29267 (I501132,I501115,I500906);
nor I_29268 (I501149,I500838,I501132);
DFFARX1 I_29269 (I501149,I3563,I500773,I500756,);
nor I_29270 (I501180,I501115,I500997);
nor I_29271 (I501197,I81967,I81958);
nor I_29272 (I500747,I501197,I501180);
not I_29273 (I501228,I501197);
nand I_29274 (I500750,I500957,I501228);
DFFARX1 I_29275 (I501197,I3563,I500773,I500762,);
DFFARX1 I_29276 (I501197,I3563,I500773,I500759,);
not I_29277 (I501317,I3570);
DFFARX1 I_29278 (I1158624,I3563,I501317,I501343,);
DFFARX1 I_29279 (I501343,I3563,I501317,I501360,);
not I_29280 (I501309,I501360);
not I_29281 (I501382,I501343);
nand I_29282 (I501399,I1158636,I1158624);
and I_29283 (I501416,I501399,I1158627);
DFFARX1 I_29284 (I501416,I3563,I501317,I501442,);
not I_29285 (I501450,I501442);
DFFARX1 I_29286 (I1158645,I3563,I501317,I501476,);
and I_29287 (I501484,I501476,I1158621);
nand I_29288 (I501501,I501476,I1158621);
nand I_29289 (I501288,I501450,I501501);
DFFARX1 I_29290 (I1158639,I3563,I501317,I501541,);
nor I_29291 (I501549,I501541,I501484);
DFFARX1 I_29292 (I501549,I3563,I501317,I501282,);
nor I_29293 (I501297,I501541,I501442);
nand I_29294 (I501594,I1158633,I1158630);
and I_29295 (I501611,I501594,I1158642);
DFFARX1 I_29296 (I501611,I3563,I501317,I501637,);
nor I_29297 (I501285,I501637,I501541);
not I_29298 (I501659,I501637);
nor I_29299 (I501676,I501659,I501450);
nor I_29300 (I501693,I501382,I501676);
DFFARX1 I_29301 (I501693,I3563,I501317,I501300,);
nor I_29302 (I501724,I501659,I501541);
nor I_29303 (I501741,I1158621,I1158630);
nor I_29304 (I501291,I501741,I501724);
not I_29305 (I501772,I501741);
nand I_29306 (I501294,I501501,I501772);
DFFARX1 I_29307 (I501741,I3563,I501317,I501306,);
DFFARX1 I_29308 (I501741,I3563,I501317,I501303,);
not I_29309 (I501861,I3570);
DFFARX1 I_29310 (I814757,I3563,I501861,I501887,);
DFFARX1 I_29311 (I501887,I3563,I501861,I501904,);
not I_29312 (I501853,I501904);
not I_29313 (I501926,I501887);
nand I_29314 (I501943,I814751,I814748);
and I_29315 (I501960,I501943,I814763);
DFFARX1 I_29316 (I501960,I3563,I501861,I501986,);
not I_29317 (I501994,I501986);
DFFARX1 I_29318 (I814751,I3563,I501861,I502020,);
and I_29319 (I502028,I502020,I814745);
nand I_29320 (I502045,I502020,I814745);
nand I_29321 (I501832,I501994,I502045);
DFFARX1 I_29322 (I814745,I3563,I501861,I502085,);
nor I_29323 (I502093,I502085,I502028);
DFFARX1 I_29324 (I502093,I3563,I501861,I501826,);
nor I_29325 (I501841,I502085,I501986);
nand I_29326 (I502138,I814760,I814754);
and I_29327 (I502155,I502138,I814748);
DFFARX1 I_29328 (I502155,I3563,I501861,I502181,);
nor I_29329 (I501829,I502181,I502085);
not I_29330 (I502203,I502181);
nor I_29331 (I502220,I502203,I501994);
nor I_29332 (I502237,I501926,I502220);
DFFARX1 I_29333 (I502237,I3563,I501861,I501844,);
nor I_29334 (I502268,I502203,I502085);
nor I_29335 (I502285,I814766,I814754);
nor I_29336 (I501835,I502285,I502268);
not I_29337 (I502316,I502285);
nand I_29338 (I501838,I502045,I502316);
DFFARX1 I_29339 (I502285,I3563,I501861,I501850,);
DFFARX1 I_29340 (I502285,I3563,I501861,I501847,);
not I_29341 (I502405,I3570);
DFFARX1 I_29342 (I1289505,I3563,I502405,I502431,);
DFFARX1 I_29343 (I502431,I3563,I502405,I502448,);
not I_29344 (I502397,I502448);
not I_29345 (I502470,I502431);
nand I_29346 (I502487,I1289502,I1289499);
and I_29347 (I502504,I502487,I1289487);
DFFARX1 I_29348 (I502504,I3563,I502405,I502530,);
not I_29349 (I502538,I502530);
DFFARX1 I_29350 (I1289511,I3563,I502405,I502564,);
and I_29351 (I502572,I502564,I1289496);
nand I_29352 (I502589,I502564,I1289496);
nand I_29353 (I502376,I502538,I502589);
DFFARX1 I_29354 (I1289490,I3563,I502405,I502629,);
nor I_29355 (I502637,I502629,I502572);
DFFARX1 I_29356 (I502637,I3563,I502405,I502370,);
nor I_29357 (I502385,I502629,I502530);
nand I_29358 (I502682,I1289487,I1289493);
and I_29359 (I502699,I502682,I1289508);
DFFARX1 I_29360 (I502699,I3563,I502405,I502725,);
nor I_29361 (I502373,I502725,I502629);
not I_29362 (I502747,I502725);
nor I_29363 (I502764,I502747,I502538);
nor I_29364 (I502781,I502470,I502764);
DFFARX1 I_29365 (I502781,I3563,I502405,I502388,);
nor I_29366 (I502812,I502747,I502629);
nor I_29367 (I502829,I1289490,I1289493);
nor I_29368 (I502379,I502829,I502812);
not I_29369 (I502860,I502829);
nand I_29370 (I502382,I502589,I502860);
DFFARX1 I_29371 (I502829,I3563,I502405,I502394,);
DFFARX1 I_29372 (I502829,I3563,I502405,I502391,);
not I_29373 (I502949,I3570);
DFFARX1 I_29374 (I873781,I3563,I502949,I502975,);
DFFARX1 I_29375 (I502975,I3563,I502949,I502992,);
not I_29376 (I502941,I502992);
not I_29377 (I503014,I502975);
nand I_29378 (I503031,I873775,I873772);
and I_29379 (I503048,I503031,I873787);
DFFARX1 I_29380 (I503048,I3563,I502949,I503074,);
not I_29381 (I503082,I503074);
DFFARX1 I_29382 (I873775,I3563,I502949,I503108,);
and I_29383 (I503116,I503108,I873769);
nand I_29384 (I503133,I503108,I873769);
nand I_29385 (I502920,I503082,I503133);
DFFARX1 I_29386 (I873769,I3563,I502949,I503173,);
nor I_29387 (I503181,I503173,I503116);
DFFARX1 I_29388 (I503181,I3563,I502949,I502914,);
nor I_29389 (I502929,I503173,I503074);
nand I_29390 (I503226,I873784,I873778);
and I_29391 (I503243,I503226,I873772);
DFFARX1 I_29392 (I503243,I3563,I502949,I503269,);
nor I_29393 (I502917,I503269,I503173);
not I_29394 (I503291,I503269);
nor I_29395 (I503308,I503291,I503082);
nor I_29396 (I503325,I503014,I503308);
DFFARX1 I_29397 (I503325,I3563,I502949,I502932,);
nor I_29398 (I503356,I503291,I503173);
nor I_29399 (I503373,I873790,I873778);
nor I_29400 (I502923,I503373,I503356);
not I_29401 (I503404,I503373);
nand I_29402 (I502926,I503133,I503404);
DFFARX1 I_29403 (I503373,I3563,I502949,I502938,);
DFFARX1 I_29404 (I503373,I3563,I502949,I502935,);
not I_29405 (I503493,I3570);
DFFARX1 I_29406 (I897496,I3563,I503493,I503519,);
DFFARX1 I_29407 (I503519,I3563,I503493,I503536,);
not I_29408 (I503485,I503536);
not I_29409 (I503558,I503519);
nand I_29410 (I503575,I897490,I897487);
and I_29411 (I503592,I503575,I897502);
DFFARX1 I_29412 (I503592,I3563,I503493,I503618,);
not I_29413 (I503626,I503618);
DFFARX1 I_29414 (I897490,I3563,I503493,I503652,);
and I_29415 (I503660,I503652,I897484);
nand I_29416 (I503677,I503652,I897484);
nand I_29417 (I503464,I503626,I503677);
DFFARX1 I_29418 (I897484,I3563,I503493,I503717,);
nor I_29419 (I503725,I503717,I503660);
DFFARX1 I_29420 (I503725,I3563,I503493,I503458,);
nor I_29421 (I503473,I503717,I503618);
nand I_29422 (I503770,I897499,I897493);
and I_29423 (I503787,I503770,I897487);
DFFARX1 I_29424 (I503787,I3563,I503493,I503813,);
nor I_29425 (I503461,I503813,I503717);
not I_29426 (I503835,I503813);
nor I_29427 (I503852,I503835,I503626);
nor I_29428 (I503869,I503558,I503852);
DFFARX1 I_29429 (I503869,I3563,I503493,I503476,);
nor I_29430 (I503900,I503835,I503717);
nor I_29431 (I503917,I897505,I897493);
nor I_29432 (I503467,I503917,I503900);
not I_29433 (I503948,I503917);
nand I_29434 (I503470,I503677,I503948);
DFFARX1 I_29435 (I503917,I3563,I503493,I503482,);
DFFARX1 I_29436 (I503917,I3563,I503493,I503479,);
not I_29437 (I504037,I3570);
DFFARX1 I_29438 (I1253484,I3563,I504037,I504063,);
DFFARX1 I_29439 (I504063,I3563,I504037,I504080,);
not I_29440 (I504029,I504080);
not I_29441 (I504102,I504063);
nand I_29442 (I504119,I1253496,I1253499);
and I_29443 (I504136,I504119,I1253502);
DFFARX1 I_29444 (I504136,I3563,I504037,I504162,);
not I_29445 (I504170,I504162);
DFFARX1 I_29446 (I1253487,I3563,I504037,I504196,);
and I_29447 (I504204,I504196,I1253493);
nand I_29448 (I504221,I504196,I1253493);
nand I_29449 (I504008,I504170,I504221);
DFFARX1 I_29450 (I1253481,I3563,I504037,I504261,);
nor I_29451 (I504269,I504261,I504204);
DFFARX1 I_29452 (I504269,I3563,I504037,I504002,);
nor I_29453 (I504017,I504261,I504162);
nand I_29454 (I504314,I1253484,I1253505);
and I_29455 (I504331,I504314,I1253490);
DFFARX1 I_29456 (I504331,I3563,I504037,I504357,);
nor I_29457 (I504005,I504357,I504261);
not I_29458 (I504379,I504357);
nor I_29459 (I504396,I504379,I504170);
nor I_29460 (I504413,I504102,I504396);
DFFARX1 I_29461 (I504413,I3563,I504037,I504020,);
nor I_29462 (I504444,I504379,I504261);
nor I_29463 (I504461,I1253481,I1253505);
nor I_29464 (I504011,I504461,I504444);
not I_29465 (I504492,I504461);
nand I_29466 (I504014,I504221,I504492);
DFFARX1 I_29467 (I504461,I3563,I504037,I504026,);
DFFARX1 I_29468 (I504461,I3563,I504037,I504023,);
not I_29469 (I504581,I3570);
DFFARX1 I_29470 (I1086490,I3563,I504581,I504607,);
DFFARX1 I_29471 (I504607,I3563,I504581,I504624,);
not I_29472 (I504573,I504624);
not I_29473 (I504646,I504607);
nand I_29474 (I504663,I1086490,I1086508);
and I_29475 (I504680,I504663,I1086502);
DFFARX1 I_29476 (I504680,I3563,I504581,I504706,);
not I_29477 (I504714,I504706);
DFFARX1 I_29478 (I1086496,I3563,I504581,I504740,);
and I_29479 (I504748,I504740,I1086505);
nand I_29480 (I504765,I504740,I1086505);
nand I_29481 (I504552,I504714,I504765);
DFFARX1 I_29482 (I1086493,I3563,I504581,I504805,);
nor I_29483 (I504813,I504805,I504748);
DFFARX1 I_29484 (I504813,I3563,I504581,I504546,);
nor I_29485 (I504561,I504805,I504706);
nand I_29486 (I504858,I1086493,I1086511);
and I_29487 (I504875,I504858,I1086496);
DFFARX1 I_29488 (I504875,I3563,I504581,I504901,);
nor I_29489 (I504549,I504901,I504805);
not I_29490 (I504923,I504901);
nor I_29491 (I504940,I504923,I504714);
nor I_29492 (I504957,I504646,I504940);
DFFARX1 I_29493 (I504957,I3563,I504581,I504564,);
nor I_29494 (I504988,I504923,I504805);
nor I_29495 (I505005,I1086499,I1086511);
nor I_29496 (I504555,I505005,I504988);
not I_29497 (I505036,I505005);
nand I_29498 (I504558,I504765,I505036);
DFFARX1 I_29499 (I505005,I3563,I504581,I504570,);
DFFARX1 I_29500 (I505005,I3563,I504581,I504567,);
not I_29501 (I505125,I3570);
DFFARX1 I_29502 (I570934,I3563,I505125,I505151,);
DFFARX1 I_29503 (I505151,I3563,I505125,I505168,);
not I_29504 (I505117,I505168);
not I_29505 (I505190,I505151);
nand I_29506 (I505207,I570937,I570955);
and I_29507 (I505224,I505207,I570943);
DFFARX1 I_29508 (I505224,I3563,I505125,I505250,);
not I_29509 (I505258,I505250);
DFFARX1 I_29510 (I570934,I3563,I505125,I505284,);
and I_29511 (I505292,I505284,I570952);
nand I_29512 (I505309,I505284,I570952);
nand I_29513 (I505096,I505258,I505309);
DFFARX1 I_29514 (I570946,I3563,I505125,I505349,);
nor I_29515 (I505357,I505349,I505292);
DFFARX1 I_29516 (I505357,I3563,I505125,I505090,);
nor I_29517 (I505105,I505349,I505250);
nand I_29518 (I505402,I570949,I570931);
and I_29519 (I505419,I505402,I570940);
DFFARX1 I_29520 (I505419,I3563,I505125,I505445,);
nor I_29521 (I505093,I505445,I505349);
not I_29522 (I505467,I505445);
nor I_29523 (I505484,I505467,I505258);
nor I_29524 (I505501,I505190,I505484);
DFFARX1 I_29525 (I505501,I3563,I505125,I505108,);
nor I_29526 (I505532,I505467,I505349);
nor I_29527 (I505549,I570931,I570931);
nor I_29528 (I505099,I505549,I505532);
not I_29529 (I505580,I505549);
nand I_29530 (I505102,I505309,I505580);
DFFARX1 I_29531 (I505549,I3563,I505125,I505114,);
DFFARX1 I_29532 (I505549,I3563,I505125,I505111,);
not I_29533 (I505669,I3570);
DFFARX1 I_29534 (I45065,I3563,I505669,I505695,);
DFFARX1 I_29535 (I505695,I3563,I505669,I505712,);
not I_29536 (I505661,I505712);
not I_29537 (I505734,I505695);
nand I_29538 (I505751,I45053,I45068);
and I_29539 (I505768,I505751,I45056);
DFFARX1 I_29540 (I505768,I3563,I505669,I505794,);
not I_29541 (I505802,I505794);
DFFARX1 I_29542 (I45077,I3563,I505669,I505828,);
and I_29543 (I505836,I505828,I45071);
nand I_29544 (I505853,I505828,I45071);
nand I_29545 (I505640,I505802,I505853);
DFFARX1 I_29546 (I45074,I3563,I505669,I505893,);
nor I_29547 (I505901,I505893,I505836);
DFFARX1 I_29548 (I505901,I3563,I505669,I505634,);
nor I_29549 (I505649,I505893,I505794);
nand I_29550 (I505946,I45053,I45056);
and I_29551 (I505963,I505946,I45059);
DFFARX1 I_29552 (I505963,I3563,I505669,I505989,);
nor I_29553 (I505637,I505989,I505893);
not I_29554 (I506011,I505989);
nor I_29555 (I506028,I506011,I505802);
nor I_29556 (I506045,I505734,I506028);
DFFARX1 I_29557 (I506045,I3563,I505669,I505652,);
nor I_29558 (I506076,I506011,I505893);
nor I_29559 (I506093,I45062,I45056);
nor I_29560 (I505643,I506093,I506076);
not I_29561 (I506124,I506093);
nand I_29562 (I505646,I505853,I506124);
DFFARX1 I_29563 (I506093,I3563,I505669,I505658,);
DFFARX1 I_29564 (I506093,I3563,I505669,I505655,);
not I_29565 (I506213,I3570);
DFFARX1 I_29566 (I390786,I3563,I506213,I506239,);
DFFARX1 I_29567 (I506239,I3563,I506213,I506256,);
not I_29568 (I506205,I506256);
not I_29569 (I506278,I506239);
nand I_29570 (I506295,I390765,I390789);
and I_29571 (I506312,I506295,I390792);
DFFARX1 I_29572 (I506312,I3563,I506213,I506338,);
not I_29573 (I506346,I506338);
DFFARX1 I_29574 (I390774,I3563,I506213,I506372,);
and I_29575 (I506380,I506372,I390780);
nand I_29576 (I506397,I506372,I390780);
nand I_29577 (I506184,I506346,I506397);
DFFARX1 I_29578 (I390768,I3563,I506213,I506437,);
nor I_29579 (I506445,I506437,I506380);
DFFARX1 I_29580 (I506445,I3563,I506213,I506178,);
nor I_29581 (I506193,I506437,I506338);
nand I_29582 (I506490,I390777,I390765);
and I_29583 (I506507,I506490,I390771);
DFFARX1 I_29584 (I506507,I3563,I506213,I506533,);
nor I_29585 (I506181,I506533,I506437);
not I_29586 (I506555,I506533);
nor I_29587 (I506572,I506555,I506346);
nor I_29588 (I506589,I506278,I506572);
DFFARX1 I_29589 (I506589,I3563,I506213,I506196,);
nor I_29590 (I506620,I506555,I506437);
nor I_29591 (I506637,I390783,I390765);
nor I_29592 (I506187,I506637,I506620);
not I_29593 (I506668,I506637);
nand I_29594 (I506190,I506397,I506668);
DFFARX1 I_29595 (I506637,I3563,I506213,I506202,);
DFFARX1 I_29596 (I506637,I3563,I506213,I506199,);
not I_29597 (I506757,I3570);
DFFARX1 I_29598 (I61923,I3563,I506757,I506783,);
DFFARX1 I_29599 (I506783,I3563,I506757,I506800,);
not I_29600 (I506749,I506800);
not I_29601 (I506822,I506783);
nand I_29602 (I506839,I61938,I61917);
and I_29603 (I506856,I506839,I61920);
DFFARX1 I_29604 (I506856,I3563,I506757,I506882,);
not I_29605 (I506890,I506882);
DFFARX1 I_29606 (I61926,I3563,I506757,I506916,);
and I_29607 (I506924,I506916,I61920);
nand I_29608 (I506941,I506916,I61920);
nand I_29609 (I506728,I506890,I506941);
DFFARX1 I_29610 (I61935,I3563,I506757,I506981,);
nor I_29611 (I506989,I506981,I506924);
DFFARX1 I_29612 (I506989,I3563,I506757,I506722,);
nor I_29613 (I506737,I506981,I506882);
nand I_29614 (I507034,I61917,I61932);
and I_29615 (I507051,I507034,I61929);
DFFARX1 I_29616 (I507051,I3563,I506757,I507077,);
nor I_29617 (I506725,I507077,I506981);
not I_29618 (I507099,I507077);
nor I_29619 (I507116,I507099,I506890);
nor I_29620 (I507133,I506822,I507116);
DFFARX1 I_29621 (I507133,I3563,I506757,I506740,);
nor I_29622 (I507164,I507099,I506981);
nor I_29623 (I507181,I61941,I61932);
nor I_29624 (I506731,I507181,I507164);
not I_29625 (I507212,I507181);
nand I_29626 (I506734,I506941,I507212);
DFFARX1 I_29627 (I507181,I3563,I506757,I506746,);
DFFARX1 I_29628 (I507181,I3563,I506757,I506743,);
not I_29629 (I507301,I3570);
DFFARX1 I_29630 (I98286,I3563,I507301,I507327,);
DFFARX1 I_29631 (I507327,I3563,I507301,I507344,);
not I_29632 (I507293,I507344);
not I_29633 (I507366,I507327);
nand I_29634 (I507383,I98301,I98280);
and I_29635 (I507400,I507383,I98283);
DFFARX1 I_29636 (I507400,I3563,I507301,I507426,);
not I_29637 (I507434,I507426);
DFFARX1 I_29638 (I98289,I3563,I507301,I507460,);
and I_29639 (I507468,I507460,I98283);
nand I_29640 (I507485,I507460,I98283);
nand I_29641 (I507272,I507434,I507485);
DFFARX1 I_29642 (I98298,I3563,I507301,I507525,);
nor I_29643 (I507533,I507525,I507468);
DFFARX1 I_29644 (I507533,I3563,I507301,I507266,);
nor I_29645 (I507281,I507525,I507426);
nand I_29646 (I507578,I98280,I98295);
and I_29647 (I507595,I507578,I98292);
DFFARX1 I_29648 (I507595,I3563,I507301,I507621,);
nor I_29649 (I507269,I507621,I507525);
not I_29650 (I507643,I507621);
nor I_29651 (I507660,I507643,I507434);
nor I_29652 (I507677,I507366,I507660);
DFFARX1 I_29653 (I507677,I3563,I507301,I507284,);
nor I_29654 (I507708,I507643,I507525);
nor I_29655 (I507725,I98304,I98295);
nor I_29656 (I507275,I507725,I507708);
not I_29657 (I507756,I507725);
nand I_29658 (I507278,I507485,I507756);
DFFARX1 I_29659 (I507725,I3563,I507301,I507290,);
DFFARX1 I_29660 (I507725,I3563,I507301,I507287,);
not I_29661 (I507845,I3570);
DFFARX1 I_29662 (I305412,I3563,I507845,I507871,);
DFFARX1 I_29663 (I507871,I3563,I507845,I507888,);
not I_29664 (I507837,I507888);
not I_29665 (I507910,I507871);
nand I_29666 (I507927,I305391,I305415);
and I_29667 (I507944,I507927,I305418);
DFFARX1 I_29668 (I507944,I3563,I507845,I507970,);
not I_29669 (I507978,I507970);
DFFARX1 I_29670 (I305400,I3563,I507845,I508004,);
and I_29671 (I508012,I508004,I305406);
nand I_29672 (I508029,I508004,I305406);
nand I_29673 (I507816,I507978,I508029);
DFFARX1 I_29674 (I305394,I3563,I507845,I508069,);
nor I_29675 (I508077,I508069,I508012);
DFFARX1 I_29676 (I508077,I3563,I507845,I507810,);
nor I_29677 (I507825,I508069,I507970);
nand I_29678 (I508122,I305403,I305391);
and I_29679 (I508139,I508122,I305397);
DFFARX1 I_29680 (I508139,I3563,I507845,I508165,);
nor I_29681 (I507813,I508165,I508069);
not I_29682 (I508187,I508165);
nor I_29683 (I508204,I508187,I507978);
nor I_29684 (I508221,I507910,I508204);
DFFARX1 I_29685 (I508221,I3563,I507845,I507828,);
nor I_29686 (I508252,I508187,I508069);
nor I_29687 (I508269,I305409,I305391);
nor I_29688 (I507819,I508269,I508252);
not I_29689 (I508300,I508269);
nand I_29690 (I507822,I508029,I508300);
DFFARX1 I_29691 (I508269,I3563,I507845,I507834,);
DFFARX1 I_29692 (I508269,I3563,I507845,I507831,);
not I_29693 (I508389,I3570);
DFFARX1 I_29694 (I1279052,I3563,I508389,I508415,);
DFFARX1 I_29695 (I508415,I3563,I508389,I508432,);
not I_29696 (I508381,I508432);
not I_29697 (I508454,I508415);
nand I_29698 (I508471,I1279064,I1279067);
and I_29699 (I508488,I508471,I1279070);
DFFARX1 I_29700 (I508488,I3563,I508389,I508514,);
not I_29701 (I508522,I508514);
DFFARX1 I_29702 (I1279055,I3563,I508389,I508548,);
and I_29703 (I508556,I508548,I1279061);
nand I_29704 (I508573,I508548,I1279061);
nand I_29705 (I508360,I508522,I508573);
DFFARX1 I_29706 (I1279049,I3563,I508389,I508613,);
nor I_29707 (I508621,I508613,I508556);
DFFARX1 I_29708 (I508621,I3563,I508389,I508354,);
nor I_29709 (I508369,I508613,I508514);
nand I_29710 (I508666,I1279052,I1279073);
and I_29711 (I508683,I508666,I1279058);
DFFARX1 I_29712 (I508683,I3563,I508389,I508709,);
nor I_29713 (I508357,I508709,I508613);
not I_29714 (I508731,I508709);
nor I_29715 (I508748,I508731,I508522);
nor I_29716 (I508765,I508454,I508748);
DFFARX1 I_29717 (I508765,I3563,I508389,I508372,);
nor I_29718 (I508796,I508731,I508613);
nor I_29719 (I508813,I1279049,I1279073);
nor I_29720 (I508363,I508813,I508796);
not I_29721 (I508844,I508813);
nand I_29722 (I508366,I508573,I508844);
DFFARX1 I_29723 (I508813,I3563,I508389,I508378,);
DFFARX1 I_29724 (I508813,I3563,I508389,I508375,);
not I_29725 (I508933,I3570);
DFFARX1 I_29726 (I1339290,I3563,I508933,I508959,);
DFFARX1 I_29727 (I508959,I3563,I508933,I508976,);
not I_29728 (I508925,I508976);
not I_29729 (I508998,I508959);
nand I_29730 (I509015,I1339266,I1339287);
and I_29731 (I509032,I509015,I1339284);
DFFARX1 I_29732 (I509032,I3563,I508933,I509058,);
not I_29733 (I509066,I509058);
DFFARX1 I_29734 (I1339263,I3563,I508933,I509092,);
and I_29735 (I509100,I509092,I1339275);
nand I_29736 (I509117,I509092,I1339275);
nand I_29737 (I508904,I509066,I509117);
DFFARX1 I_29738 (I1339278,I3563,I508933,I509157,);
nor I_29739 (I509165,I509157,I509100);
DFFARX1 I_29740 (I509165,I3563,I508933,I508898,);
nor I_29741 (I508913,I509157,I509058);
nand I_29742 (I509210,I1339281,I1339269);
and I_29743 (I509227,I509210,I1339272);
DFFARX1 I_29744 (I509227,I3563,I508933,I509253,);
nor I_29745 (I508901,I509253,I509157);
not I_29746 (I509275,I509253);
nor I_29747 (I509292,I509275,I509066);
nor I_29748 (I509309,I508998,I509292);
DFFARX1 I_29749 (I509309,I3563,I508933,I508916,);
nor I_29750 (I509340,I509275,I509157);
nor I_29751 (I509357,I1339263,I1339269);
nor I_29752 (I508907,I509357,I509340);
not I_29753 (I509388,I509357);
nand I_29754 (I508910,I509117,I509388);
DFFARX1 I_29755 (I509357,I3563,I508933,I508922,);
DFFARX1 I_29756 (I509357,I3563,I508933,I508919,);
not I_29757 (I509477,I3570);
DFFARX1 I_29758 (I17661,I3563,I509477,I509503,);
DFFARX1 I_29759 (I509503,I3563,I509477,I509520,);
not I_29760 (I509469,I509520);
not I_29761 (I509542,I509503);
nand I_29762 (I509559,I17649,I17664);
and I_29763 (I509576,I509559,I17652);
DFFARX1 I_29764 (I509576,I3563,I509477,I509602,);
not I_29765 (I509610,I509602);
DFFARX1 I_29766 (I17673,I3563,I509477,I509636,);
and I_29767 (I509644,I509636,I17667);
nand I_29768 (I509661,I509636,I17667);
nand I_29769 (I509448,I509610,I509661);
DFFARX1 I_29770 (I17670,I3563,I509477,I509701,);
nor I_29771 (I509709,I509701,I509644);
DFFARX1 I_29772 (I509709,I3563,I509477,I509442,);
nor I_29773 (I509457,I509701,I509602);
nand I_29774 (I509754,I17649,I17652);
and I_29775 (I509771,I509754,I17655);
DFFARX1 I_29776 (I509771,I3563,I509477,I509797,);
nor I_29777 (I509445,I509797,I509701);
not I_29778 (I509819,I509797);
nor I_29779 (I509836,I509819,I509610);
nor I_29780 (I509853,I509542,I509836);
DFFARX1 I_29781 (I509853,I3563,I509477,I509460,);
nor I_29782 (I509884,I509819,I509701);
nor I_29783 (I509901,I17658,I17652);
nor I_29784 (I509451,I509901,I509884);
not I_29785 (I509932,I509901);
nand I_29786 (I509454,I509661,I509932);
DFFARX1 I_29787 (I509901,I3563,I509477,I509466,);
DFFARX1 I_29788 (I509901,I3563,I509477,I509463,);
not I_29789 (I510021,I3570);
DFFARX1 I_29790 (I325438,I3563,I510021,I510047,);
DFFARX1 I_29791 (I510047,I3563,I510021,I510064,);
not I_29792 (I510013,I510064);
not I_29793 (I510086,I510047);
nand I_29794 (I510103,I325417,I325441);
and I_29795 (I510120,I510103,I325444);
DFFARX1 I_29796 (I510120,I3563,I510021,I510146,);
not I_29797 (I510154,I510146);
DFFARX1 I_29798 (I325426,I3563,I510021,I510180,);
and I_29799 (I510188,I510180,I325432);
nand I_29800 (I510205,I510180,I325432);
nand I_29801 (I509992,I510154,I510205);
DFFARX1 I_29802 (I325420,I3563,I510021,I510245,);
nor I_29803 (I510253,I510245,I510188);
DFFARX1 I_29804 (I510253,I3563,I510021,I509986,);
nor I_29805 (I510001,I510245,I510146);
nand I_29806 (I510298,I325429,I325417);
and I_29807 (I510315,I510298,I325423);
DFFARX1 I_29808 (I510315,I3563,I510021,I510341,);
nor I_29809 (I509989,I510341,I510245);
not I_29810 (I510363,I510341);
nor I_29811 (I510380,I510363,I510154);
nor I_29812 (I510397,I510086,I510380);
DFFARX1 I_29813 (I510397,I3563,I510021,I510004,);
nor I_29814 (I510428,I510363,I510245);
nor I_29815 (I510445,I325435,I325417);
nor I_29816 (I509995,I510445,I510428);
not I_29817 (I510476,I510445);
nand I_29818 (I509998,I510205,I510476);
DFFARX1 I_29819 (I510445,I3563,I510021,I510010,);
DFFARX1 I_29820 (I510445,I3563,I510021,I510007,);
not I_29821 (I510565,I3570);
DFFARX1 I_29822 (I559034,I3563,I510565,I510591,);
DFFARX1 I_29823 (I510591,I3563,I510565,I510608,);
not I_29824 (I510557,I510608);
not I_29825 (I510630,I510591);
nand I_29826 (I510647,I559037,I559055);
and I_29827 (I510664,I510647,I559043);
DFFARX1 I_29828 (I510664,I3563,I510565,I510690,);
not I_29829 (I510698,I510690);
DFFARX1 I_29830 (I559034,I3563,I510565,I510724,);
and I_29831 (I510732,I510724,I559052);
nand I_29832 (I510749,I510724,I559052);
nand I_29833 (I510536,I510698,I510749);
DFFARX1 I_29834 (I559046,I3563,I510565,I510789,);
nor I_29835 (I510797,I510789,I510732);
DFFARX1 I_29836 (I510797,I3563,I510565,I510530,);
nor I_29837 (I510545,I510789,I510690);
nand I_29838 (I510842,I559049,I559031);
and I_29839 (I510859,I510842,I559040);
DFFARX1 I_29840 (I510859,I3563,I510565,I510885,);
nor I_29841 (I510533,I510885,I510789);
not I_29842 (I510907,I510885);
nor I_29843 (I510924,I510907,I510698);
nor I_29844 (I510941,I510630,I510924);
DFFARX1 I_29845 (I510941,I3563,I510565,I510548,);
nor I_29846 (I510972,I510907,I510789);
nor I_29847 (I510989,I559031,I559031);
nor I_29848 (I510539,I510989,I510972);
not I_29849 (I511020,I510989);
nand I_29850 (I510542,I510749,I511020);
DFFARX1 I_29851 (I510989,I3563,I510565,I510554,);
DFFARX1 I_29852 (I510989,I3563,I510565,I510551,);
not I_29853 (I511109,I3570);
DFFARX1 I_29854 (I952349,I3563,I511109,I511135,);
DFFARX1 I_29855 (I511135,I3563,I511109,I511152,);
not I_29856 (I511101,I511152);
not I_29857 (I511174,I511135);
nand I_29858 (I511191,I952364,I952352);
and I_29859 (I511208,I511191,I952343);
DFFARX1 I_29860 (I511208,I3563,I511109,I511234,);
not I_29861 (I511242,I511234);
DFFARX1 I_29862 (I952355,I3563,I511109,I511268,);
and I_29863 (I511276,I511268,I952346);
nand I_29864 (I511293,I511268,I952346);
nand I_29865 (I511080,I511242,I511293);
DFFARX1 I_29866 (I952361,I3563,I511109,I511333,);
nor I_29867 (I511341,I511333,I511276);
DFFARX1 I_29868 (I511341,I3563,I511109,I511074,);
nor I_29869 (I511089,I511333,I511234);
nand I_29870 (I511386,I952370,I952358);
and I_29871 (I511403,I511386,I952367);
DFFARX1 I_29872 (I511403,I3563,I511109,I511429,);
nor I_29873 (I511077,I511429,I511333);
not I_29874 (I511451,I511429);
nor I_29875 (I511468,I511451,I511242);
nor I_29876 (I511485,I511174,I511468);
DFFARX1 I_29877 (I511485,I3563,I511109,I511092,);
nor I_29878 (I511516,I511451,I511333);
nor I_29879 (I511533,I952343,I952358);
nor I_29880 (I511083,I511533,I511516);
not I_29881 (I511564,I511533);
nand I_29882 (I511086,I511293,I511564);
DFFARX1 I_29883 (I511533,I3563,I511109,I511098,);
DFFARX1 I_29884 (I511533,I3563,I511109,I511095,);
not I_29885 (I511653,I3570);
DFFARX1 I_29886 (I403961,I3563,I511653,I511679,);
DFFARX1 I_29887 (I511679,I3563,I511653,I511696,);
not I_29888 (I511645,I511696);
not I_29889 (I511718,I511679);
nand I_29890 (I511735,I403940,I403964);
and I_29891 (I511752,I511735,I403967);
DFFARX1 I_29892 (I511752,I3563,I511653,I511778,);
not I_29893 (I511786,I511778);
DFFARX1 I_29894 (I403949,I3563,I511653,I511812,);
and I_29895 (I511820,I511812,I403955);
nand I_29896 (I511837,I511812,I403955);
nand I_29897 (I511624,I511786,I511837);
DFFARX1 I_29898 (I403943,I3563,I511653,I511877,);
nor I_29899 (I511885,I511877,I511820);
DFFARX1 I_29900 (I511885,I3563,I511653,I511618,);
nor I_29901 (I511633,I511877,I511778);
nand I_29902 (I511930,I403952,I403940);
and I_29903 (I511947,I511930,I403946);
DFFARX1 I_29904 (I511947,I3563,I511653,I511973,);
nor I_29905 (I511621,I511973,I511877);
not I_29906 (I511995,I511973);
nor I_29907 (I512012,I511995,I511786);
nor I_29908 (I512029,I511718,I512012);
DFFARX1 I_29909 (I512029,I3563,I511653,I511636,);
nor I_29910 (I512060,I511995,I511877);
nor I_29911 (I512077,I403958,I403940);
nor I_29912 (I511627,I512077,I512060);
not I_29913 (I512108,I512077);
nand I_29914 (I511630,I511837,I512108);
DFFARX1 I_29915 (I512077,I3563,I511653,I511642,);
DFFARX1 I_29916 (I512077,I3563,I511653,I511639,);
not I_29917 (I512197,I3570);
DFFARX1 I_29918 (I1216424,I3563,I512197,I512223,);
DFFARX1 I_29919 (I512223,I3563,I512197,I512240,);
not I_29920 (I512189,I512240);
not I_29921 (I512262,I512223);
nand I_29922 (I512279,I1216436,I1216424);
and I_29923 (I512296,I512279,I1216427);
DFFARX1 I_29924 (I512296,I3563,I512197,I512322,);
not I_29925 (I512330,I512322);
DFFARX1 I_29926 (I1216445,I3563,I512197,I512356,);
and I_29927 (I512364,I512356,I1216421);
nand I_29928 (I512381,I512356,I1216421);
nand I_29929 (I512168,I512330,I512381);
DFFARX1 I_29930 (I1216439,I3563,I512197,I512421,);
nor I_29931 (I512429,I512421,I512364);
DFFARX1 I_29932 (I512429,I3563,I512197,I512162,);
nor I_29933 (I512177,I512421,I512322);
nand I_29934 (I512474,I1216433,I1216430);
and I_29935 (I512491,I512474,I1216442);
DFFARX1 I_29936 (I512491,I3563,I512197,I512517,);
nor I_29937 (I512165,I512517,I512421);
not I_29938 (I512539,I512517);
nor I_29939 (I512556,I512539,I512330);
nor I_29940 (I512573,I512262,I512556);
DFFARX1 I_29941 (I512573,I3563,I512197,I512180,);
nor I_29942 (I512604,I512539,I512421);
nor I_29943 (I512621,I1216421,I1216430);
nor I_29944 (I512171,I512621,I512604);
not I_29945 (I512652,I512621);
nand I_29946 (I512174,I512381,I512652);
DFFARX1 I_29947 (I512621,I3563,I512197,I512186,);
DFFARX1 I_29948 (I512621,I3563,I512197,I512183,);
not I_29949 (I512741,I3570);
DFFARX1 I_29950 (I211322,I3563,I512741,I512767,);
DFFARX1 I_29951 (I512767,I3563,I512741,I512784,);
not I_29952 (I512733,I512784);
not I_29953 (I512806,I512767);
nand I_29954 (I512823,I211334,I211313);
and I_29955 (I512840,I512823,I211316);
DFFARX1 I_29956 (I512840,I3563,I512741,I512866,);
not I_29957 (I512874,I512866);
DFFARX1 I_29958 (I211325,I3563,I512741,I512900,);
and I_29959 (I512908,I512900,I211337);
nand I_29960 (I512925,I512900,I211337);
nand I_29961 (I512712,I512874,I512925);
DFFARX1 I_29962 (I211331,I3563,I512741,I512965,);
nor I_29963 (I512973,I512965,I512908);
DFFARX1 I_29964 (I512973,I3563,I512741,I512706,);
nor I_29965 (I512721,I512965,I512866);
nand I_29966 (I513018,I211319,I211316);
and I_29967 (I513035,I513018,I211328);
DFFARX1 I_29968 (I513035,I3563,I512741,I513061,);
nor I_29969 (I512709,I513061,I512965);
not I_29970 (I513083,I513061);
nor I_29971 (I513100,I513083,I512874);
nor I_29972 (I513117,I512806,I513100);
DFFARX1 I_29973 (I513117,I3563,I512741,I512724,);
nor I_29974 (I513148,I513083,I512965);
nor I_29975 (I513165,I211313,I211316);
nor I_29976 (I512715,I513165,I513148);
not I_29977 (I513196,I513165);
nand I_29978 (I512718,I512925,I513196);
DFFARX1 I_29979 (I513165,I3563,I512741,I512730,);
DFFARX1 I_29980 (I513165,I3563,I512741,I512727,);
not I_29981 (I513285,I3570);
DFFARX1 I_29982 (I200017,I3563,I513285,I513311,);
DFFARX1 I_29983 (I513311,I3563,I513285,I513328,);
not I_29984 (I513277,I513328);
not I_29985 (I513350,I513311);
nand I_29986 (I513367,I200029,I200008);
and I_29987 (I513384,I513367,I200011);
DFFARX1 I_29988 (I513384,I3563,I513285,I513410,);
not I_29989 (I513418,I513410);
DFFARX1 I_29990 (I200020,I3563,I513285,I513444,);
and I_29991 (I513452,I513444,I200032);
nand I_29992 (I513469,I513444,I200032);
nand I_29993 (I513256,I513418,I513469);
DFFARX1 I_29994 (I200026,I3563,I513285,I513509,);
nor I_29995 (I513517,I513509,I513452);
DFFARX1 I_29996 (I513517,I3563,I513285,I513250,);
nor I_29997 (I513265,I513509,I513410);
nand I_29998 (I513562,I200014,I200011);
and I_29999 (I513579,I513562,I200023);
DFFARX1 I_30000 (I513579,I3563,I513285,I513605,);
nor I_30001 (I513253,I513605,I513509);
not I_30002 (I513627,I513605);
nor I_30003 (I513644,I513627,I513418);
nor I_30004 (I513661,I513350,I513644);
DFFARX1 I_30005 (I513661,I3563,I513285,I513268,);
nor I_30006 (I513692,I513627,I513509);
nor I_30007 (I513709,I200008,I200011);
nor I_30008 (I513259,I513709,I513692);
not I_30009 (I513740,I513709);
nand I_30010 (I513262,I513469,I513740);
DFFARX1 I_30011 (I513709,I3563,I513285,I513274,);
DFFARX1 I_30012 (I513709,I3563,I513285,I513271,);
not I_30013 (I513829,I3570);
DFFARX1 I_30014 (I1380345,I3563,I513829,I513855,);
DFFARX1 I_30015 (I513855,I3563,I513829,I513872,);
not I_30016 (I513821,I513872);
not I_30017 (I513894,I513855);
nand I_30018 (I513911,I1380321,I1380342);
and I_30019 (I513928,I513911,I1380339);
DFFARX1 I_30020 (I513928,I3563,I513829,I513954,);
not I_30021 (I513962,I513954);
DFFARX1 I_30022 (I1380318,I3563,I513829,I513988,);
and I_30023 (I513996,I513988,I1380330);
nand I_30024 (I514013,I513988,I1380330);
nand I_30025 (I513800,I513962,I514013);
DFFARX1 I_30026 (I1380333,I3563,I513829,I514053,);
nor I_30027 (I514061,I514053,I513996);
DFFARX1 I_30028 (I514061,I3563,I513829,I513794,);
nor I_30029 (I513809,I514053,I513954);
nand I_30030 (I514106,I1380336,I1380324);
and I_30031 (I514123,I514106,I1380327);
DFFARX1 I_30032 (I514123,I3563,I513829,I514149,);
nor I_30033 (I513797,I514149,I514053);
not I_30034 (I514171,I514149);
nor I_30035 (I514188,I514171,I513962);
nor I_30036 (I514205,I513894,I514188);
DFFARX1 I_30037 (I514205,I3563,I513829,I513812,);
nor I_30038 (I514236,I514171,I514053);
nor I_30039 (I514253,I1380318,I1380324);
nor I_30040 (I513803,I514253,I514236);
not I_30041 (I514284,I514253);
nand I_30042 (I513806,I514013,I514284);
DFFARX1 I_30043 (I514253,I3563,I513829,I513818,);
DFFARX1 I_30044 (I514253,I3563,I513829,I513815,);
not I_30045 (I514373,I3570);
DFFARX1 I_30046 (I1361305,I3563,I514373,I514399,);
DFFARX1 I_30047 (I514399,I3563,I514373,I514416,);
not I_30048 (I514365,I514416);
not I_30049 (I514438,I514399);
nand I_30050 (I514455,I1361281,I1361302);
and I_30051 (I514472,I514455,I1361299);
DFFARX1 I_30052 (I514472,I3563,I514373,I514498,);
not I_30053 (I514506,I514498);
DFFARX1 I_30054 (I1361278,I3563,I514373,I514532,);
and I_30055 (I514540,I514532,I1361290);
nand I_30056 (I514557,I514532,I1361290);
nand I_30057 (I514344,I514506,I514557);
DFFARX1 I_30058 (I1361293,I3563,I514373,I514597,);
nor I_30059 (I514605,I514597,I514540);
DFFARX1 I_30060 (I514605,I3563,I514373,I514338,);
nor I_30061 (I514353,I514597,I514498);
nand I_30062 (I514650,I1361296,I1361284);
and I_30063 (I514667,I514650,I1361287);
DFFARX1 I_30064 (I514667,I3563,I514373,I514693,);
nor I_30065 (I514341,I514693,I514597);
not I_30066 (I514715,I514693);
nor I_30067 (I514732,I514715,I514506);
nor I_30068 (I514749,I514438,I514732);
DFFARX1 I_30069 (I514749,I3563,I514373,I514356,);
nor I_30070 (I514780,I514715,I514597);
nor I_30071 (I514797,I1361278,I1361284);
nor I_30072 (I514347,I514797,I514780);
not I_30073 (I514828,I514797);
nand I_30074 (I514350,I514557,I514828);
DFFARX1 I_30075 (I514797,I3563,I514373,I514362,);
DFFARX1 I_30076 (I514797,I3563,I514373,I514359,);
not I_30077 (I514917,I3570);
DFFARX1 I_30078 (I854282,I3563,I514917,I514943,);
DFFARX1 I_30079 (I514943,I3563,I514917,I514960,);
not I_30080 (I514909,I514960);
not I_30081 (I514982,I514943);
nand I_30082 (I514999,I854276,I854273);
and I_30083 (I515016,I514999,I854288);
DFFARX1 I_30084 (I515016,I3563,I514917,I515042,);
not I_30085 (I515050,I515042);
DFFARX1 I_30086 (I854276,I3563,I514917,I515076,);
and I_30087 (I515084,I515076,I854270);
nand I_30088 (I515101,I515076,I854270);
nand I_30089 (I514888,I515050,I515101);
DFFARX1 I_30090 (I854270,I3563,I514917,I515141,);
nor I_30091 (I515149,I515141,I515084);
DFFARX1 I_30092 (I515149,I3563,I514917,I514882,);
nor I_30093 (I514897,I515141,I515042);
nand I_30094 (I515194,I854285,I854279);
and I_30095 (I515211,I515194,I854273);
DFFARX1 I_30096 (I515211,I3563,I514917,I515237,);
nor I_30097 (I514885,I515237,I515141);
not I_30098 (I515259,I515237);
nor I_30099 (I515276,I515259,I515050);
nor I_30100 (I515293,I514982,I515276);
DFFARX1 I_30101 (I515293,I3563,I514917,I514900,);
nor I_30102 (I515324,I515259,I515141);
nor I_30103 (I515341,I854291,I854279);
nor I_30104 (I514891,I515341,I515324);
not I_30105 (I515372,I515341);
nand I_30106 (I514894,I515101,I515372);
DFFARX1 I_30107 (I515341,I3563,I514917,I514906,);
DFFARX1 I_30108 (I515341,I3563,I514917,I514903,);
not I_30109 (I515461,I3570);
DFFARX1 I_30110 (I1310891,I3563,I515461,I515487,);
DFFARX1 I_30111 (I515487,I3563,I515461,I515504,);
not I_30112 (I515453,I515504);
not I_30113 (I515526,I515487);
nand I_30114 (I515543,I1310888,I1310885);
and I_30115 (I515560,I515543,I1310873);
DFFARX1 I_30116 (I515560,I3563,I515461,I515586,);
not I_30117 (I515594,I515586);
DFFARX1 I_30118 (I1310897,I3563,I515461,I515620,);
and I_30119 (I515628,I515620,I1310882);
nand I_30120 (I515645,I515620,I1310882);
nand I_30121 (I515432,I515594,I515645);
DFFARX1 I_30122 (I1310876,I3563,I515461,I515685,);
nor I_30123 (I515693,I515685,I515628);
DFFARX1 I_30124 (I515693,I3563,I515461,I515426,);
nor I_30125 (I515441,I515685,I515586);
nand I_30126 (I515738,I1310873,I1310879);
and I_30127 (I515755,I515738,I1310894);
DFFARX1 I_30128 (I515755,I3563,I515461,I515781,);
nor I_30129 (I515429,I515781,I515685);
not I_30130 (I515803,I515781);
nor I_30131 (I515820,I515803,I515594);
nor I_30132 (I515837,I515526,I515820);
DFFARX1 I_30133 (I515837,I3563,I515461,I515444,);
nor I_30134 (I515868,I515803,I515685);
nor I_30135 (I515885,I1310876,I1310879);
nor I_30136 (I515435,I515885,I515868);
not I_30137 (I515916,I515885);
nand I_30138 (I515438,I515645,I515916);
DFFARX1 I_30139 (I515885,I3563,I515461,I515450,);
DFFARX1 I_30140 (I515885,I3563,I515461,I515447,);
not I_30141 (I516005,I3570);
DFFARX1 I_30142 (I738180,I3563,I516005,I516031,);
DFFARX1 I_30143 (I516031,I3563,I516005,I516048,);
not I_30144 (I515997,I516048);
not I_30145 (I516070,I516031);
nand I_30146 (I516087,I738201,I738192);
and I_30147 (I516104,I516087,I738180);
DFFARX1 I_30148 (I516104,I3563,I516005,I516130,);
not I_30149 (I516138,I516130);
DFFARX1 I_30150 (I738186,I3563,I516005,I516164,);
and I_30151 (I516172,I516164,I738183);
nand I_30152 (I516189,I516164,I738183);
nand I_30153 (I515976,I516138,I516189);
DFFARX1 I_30154 (I738177,I3563,I516005,I516229,);
nor I_30155 (I516237,I516229,I516172);
DFFARX1 I_30156 (I516237,I3563,I516005,I515970,);
nor I_30157 (I515985,I516229,I516130);
nand I_30158 (I516282,I738177,I738189);
and I_30159 (I516299,I516282,I738198);
DFFARX1 I_30160 (I516299,I3563,I516005,I516325,);
nor I_30161 (I515973,I516325,I516229);
not I_30162 (I516347,I516325);
nor I_30163 (I516364,I516347,I516138);
nor I_30164 (I516381,I516070,I516364);
DFFARX1 I_30165 (I516381,I3563,I516005,I515988,);
nor I_30166 (I516412,I516347,I516229);
nor I_30167 (I516429,I738195,I738189);
nor I_30168 (I515979,I516429,I516412);
not I_30169 (I516460,I516429);
nand I_30170 (I515982,I516189,I516460);
DFFARX1 I_30171 (I516429,I3563,I516005,I515994,);
DFFARX1 I_30172 (I516429,I3563,I516005,I515991,);
not I_30173 (I516549,I3570);
DFFARX1 I_30174 (I1144752,I3563,I516549,I516575,);
DFFARX1 I_30175 (I516575,I3563,I516549,I516592,);
not I_30176 (I516541,I516592);
not I_30177 (I516614,I516575);
nand I_30178 (I516631,I1144764,I1144752);
and I_30179 (I516648,I516631,I1144755);
DFFARX1 I_30180 (I516648,I3563,I516549,I516674,);
not I_30181 (I516682,I516674);
DFFARX1 I_30182 (I1144773,I3563,I516549,I516708,);
and I_30183 (I516716,I516708,I1144749);
nand I_30184 (I516733,I516708,I1144749);
nand I_30185 (I516520,I516682,I516733);
DFFARX1 I_30186 (I1144767,I3563,I516549,I516773,);
nor I_30187 (I516781,I516773,I516716);
DFFARX1 I_30188 (I516781,I3563,I516549,I516514,);
nor I_30189 (I516529,I516773,I516674);
nand I_30190 (I516826,I1144761,I1144758);
and I_30191 (I516843,I516826,I1144770);
DFFARX1 I_30192 (I516843,I3563,I516549,I516869,);
nor I_30193 (I516517,I516869,I516773);
not I_30194 (I516891,I516869);
nor I_30195 (I516908,I516891,I516682);
nor I_30196 (I516925,I516614,I516908);
DFFARX1 I_30197 (I516925,I3563,I516549,I516532,);
nor I_30198 (I516956,I516891,I516773);
nor I_30199 (I516973,I1144749,I1144758);
nor I_30200 (I516523,I516973,I516956);
not I_30201 (I517004,I516973);
nand I_30202 (I516526,I516733,I517004);
DFFARX1 I_30203 (I516973,I3563,I516549,I516538,);
DFFARX1 I_30204 (I516973,I3563,I516549,I516535,);
not I_30205 (I517093,I3570);
DFFARX1 I_30206 (I1007259,I3563,I517093,I517119,);
DFFARX1 I_30207 (I517119,I3563,I517093,I517136,);
not I_30208 (I517085,I517136);
not I_30209 (I517158,I517119);
nand I_30210 (I517175,I1007274,I1007262);
and I_30211 (I517192,I517175,I1007253);
DFFARX1 I_30212 (I517192,I3563,I517093,I517218,);
not I_30213 (I517226,I517218);
DFFARX1 I_30214 (I1007265,I3563,I517093,I517252,);
and I_30215 (I517260,I517252,I1007256);
nand I_30216 (I517277,I517252,I1007256);
nand I_30217 (I517064,I517226,I517277);
DFFARX1 I_30218 (I1007271,I3563,I517093,I517317,);
nor I_30219 (I517325,I517317,I517260);
DFFARX1 I_30220 (I517325,I3563,I517093,I517058,);
nor I_30221 (I517073,I517317,I517218);
nand I_30222 (I517370,I1007280,I1007268);
and I_30223 (I517387,I517370,I1007277);
DFFARX1 I_30224 (I517387,I3563,I517093,I517413,);
nor I_30225 (I517061,I517413,I517317);
not I_30226 (I517435,I517413);
nor I_30227 (I517452,I517435,I517226);
nor I_30228 (I517469,I517158,I517452);
DFFARX1 I_30229 (I517469,I3563,I517093,I517076,);
nor I_30230 (I517500,I517435,I517317);
nor I_30231 (I517517,I1007253,I1007268);
nor I_30232 (I517067,I517517,I517500);
not I_30233 (I517548,I517517);
nand I_30234 (I517070,I517277,I517548);
DFFARX1 I_30235 (I517517,I3563,I517093,I517082,);
DFFARX1 I_30236 (I517517,I3563,I517093,I517079,);
not I_30237 (I517637,I3570);
DFFARX1 I_30238 (I542374,I3563,I517637,I517663,);
DFFARX1 I_30239 (I517663,I3563,I517637,I517680,);
not I_30240 (I517629,I517680);
not I_30241 (I517702,I517663);
nand I_30242 (I517719,I542377,I542395);
and I_30243 (I517736,I517719,I542383);
DFFARX1 I_30244 (I517736,I3563,I517637,I517762,);
not I_30245 (I517770,I517762);
DFFARX1 I_30246 (I542374,I3563,I517637,I517796,);
and I_30247 (I517804,I517796,I542392);
nand I_30248 (I517821,I517796,I542392);
nand I_30249 (I517608,I517770,I517821);
DFFARX1 I_30250 (I542386,I3563,I517637,I517861,);
nor I_30251 (I517869,I517861,I517804);
DFFARX1 I_30252 (I517869,I3563,I517637,I517602,);
nor I_30253 (I517617,I517861,I517762);
nand I_30254 (I517914,I542389,I542371);
and I_30255 (I517931,I517914,I542380);
DFFARX1 I_30256 (I517931,I3563,I517637,I517957,);
nor I_30257 (I517605,I517957,I517861);
not I_30258 (I517979,I517957);
nor I_30259 (I517996,I517979,I517770);
nor I_30260 (I518013,I517702,I517996);
DFFARX1 I_30261 (I518013,I3563,I517637,I517620,);
nor I_30262 (I518044,I517979,I517861);
nor I_30263 (I518061,I542371,I542371);
nor I_30264 (I517611,I518061,I518044);
not I_30265 (I518092,I518061);
nand I_30266 (I517614,I517821,I518092);
DFFARX1 I_30267 (I518061,I3563,I517637,I517626,);
DFFARX1 I_30268 (I518061,I3563,I517637,I517623,);
not I_30269 (I518181,I3570);
DFFARX1 I_30270 (I43484,I3563,I518181,I518207,);
DFFARX1 I_30271 (I518207,I3563,I518181,I518224,);
not I_30272 (I518173,I518224);
not I_30273 (I518246,I518207);
nand I_30274 (I518263,I43472,I43487);
and I_30275 (I518280,I518263,I43475);
DFFARX1 I_30276 (I518280,I3563,I518181,I518306,);
not I_30277 (I518314,I518306);
DFFARX1 I_30278 (I43496,I3563,I518181,I518340,);
and I_30279 (I518348,I518340,I43490);
nand I_30280 (I518365,I518340,I43490);
nand I_30281 (I518152,I518314,I518365);
DFFARX1 I_30282 (I43493,I3563,I518181,I518405,);
nor I_30283 (I518413,I518405,I518348);
DFFARX1 I_30284 (I518413,I3563,I518181,I518146,);
nor I_30285 (I518161,I518405,I518306);
nand I_30286 (I518458,I43472,I43475);
and I_30287 (I518475,I518458,I43478);
DFFARX1 I_30288 (I518475,I3563,I518181,I518501,);
nor I_30289 (I518149,I518501,I518405);
not I_30290 (I518523,I518501);
nor I_30291 (I518540,I518523,I518314);
nor I_30292 (I518557,I518246,I518540);
DFFARX1 I_30293 (I518557,I3563,I518181,I518164,);
nor I_30294 (I518588,I518523,I518405);
nor I_30295 (I518605,I43481,I43475);
nor I_30296 (I518155,I518605,I518588);
not I_30297 (I518636,I518605);
nand I_30298 (I518158,I518365,I518636);
DFFARX1 I_30299 (I518605,I3563,I518181,I518170,);
DFFARX1 I_30300 (I518605,I3563,I518181,I518167,);
not I_30301 (I518725,I3570);
DFFARX1 I_30302 (I937491,I3563,I518725,I518751,);
DFFARX1 I_30303 (I518751,I3563,I518725,I518768,);
not I_30304 (I518717,I518768);
not I_30305 (I518790,I518751);
nand I_30306 (I518807,I937506,I937494);
and I_30307 (I518824,I518807,I937485);
DFFARX1 I_30308 (I518824,I3563,I518725,I518850,);
not I_30309 (I518858,I518850);
DFFARX1 I_30310 (I937497,I3563,I518725,I518884,);
and I_30311 (I518892,I518884,I937488);
nand I_30312 (I518909,I518884,I937488);
nand I_30313 (I518696,I518858,I518909);
DFFARX1 I_30314 (I937503,I3563,I518725,I518949,);
nor I_30315 (I518957,I518949,I518892);
DFFARX1 I_30316 (I518957,I3563,I518725,I518690,);
nor I_30317 (I518705,I518949,I518850);
nand I_30318 (I519002,I937512,I937500);
and I_30319 (I519019,I519002,I937509);
DFFARX1 I_30320 (I519019,I3563,I518725,I519045,);
nor I_30321 (I518693,I519045,I518949);
not I_30322 (I519067,I519045);
nor I_30323 (I519084,I519067,I518858);
nor I_30324 (I519101,I518790,I519084);
DFFARX1 I_30325 (I519101,I3563,I518725,I518708,);
nor I_30326 (I519132,I519067,I518949);
nor I_30327 (I519149,I937485,I937500);
nor I_30328 (I518699,I519149,I519132);
not I_30329 (I519180,I519149);
nand I_30330 (I518702,I518909,I519180);
DFFARX1 I_30331 (I519149,I3563,I518725,I518714,);
DFFARX1 I_30332 (I519149,I3563,I518725,I518711,);
not I_30333 (I519269,I3570);
DFFARX1 I_30334 (I160155,I3563,I519269,I519295,);
DFFARX1 I_30335 (I519295,I3563,I519269,I519312,);
not I_30336 (I519261,I519312);
not I_30337 (I519334,I519295);
nand I_30338 (I519351,I160164,I160167);
and I_30339 (I519368,I519351,I160146);
DFFARX1 I_30340 (I519368,I3563,I519269,I519394,);
not I_30341 (I519402,I519394);
DFFARX1 I_30342 (I160161,I3563,I519269,I519428,);
and I_30343 (I519436,I519428,I160149);
nand I_30344 (I519453,I519428,I160149);
nand I_30345 (I519240,I519402,I519453);
DFFARX1 I_30346 (I160143,I3563,I519269,I519493,);
nor I_30347 (I519501,I519493,I519436);
DFFARX1 I_30348 (I519501,I3563,I519269,I519234,);
nor I_30349 (I519249,I519493,I519394);
nand I_30350 (I519546,I160158,I160152);
and I_30351 (I519563,I519546,I160143);
DFFARX1 I_30352 (I519563,I3563,I519269,I519589,);
nor I_30353 (I519237,I519589,I519493);
not I_30354 (I519611,I519589);
nor I_30355 (I519628,I519611,I519402);
nor I_30356 (I519645,I519334,I519628);
DFFARX1 I_30357 (I519645,I3563,I519269,I519252,);
nor I_30358 (I519676,I519611,I519493);
nor I_30359 (I519693,I160170,I160152);
nor I_30360 (I519243,I519693,I519676);
not I_30361 (I519724,I519693);
nand I_30362 (I519246,I519453,I519724);
DFFARX1 I_30363 (I519693,I3563,I519269,I519258,);
DFFARX1 I_30364 (I519693,I3563,I519269,I519255,);
not I_30365 (I519813,I3570);
DFFARX1 I_30366 (I805806,I3563,I519813,I519839,);
DFFARX1 I_30367 (I519839,I3563,I519813,I519856,);
not I_30368 (I519805,I519856);
not I_30369 (I519878,I519839);
nand I_30370 (I519895,I805827,I805818);
and I_30371 (I519912,I519895,I805806);
DFFARX1 I_30372 (I519912,I3563,I519813,I519938,);
not I_30373 (I519946,I519938);
DFFARX1 I_30374 (I805812,I3563,I519813,I519972,);
and I_30375 (I519980,I519972,I805809);
nand I_30376 (I519997,I519972,I805809);
nand I_30377 (I519784,I519946,I519997);
DFFARX1 I_30378 (I805803,I3563,I519813,I520037,);
nor I_30379 (I520045,I520037,I519980);
DFFARX1 I_30380 (I520045,I3563,I519813,I519778,);
nor I_30381 (I519793,I520037,I519938);
nand I_30382 (I520090,I805803,I805815);
and I_30383 (I520107,I520090,I805824);
DFFARX1 I_30384 (I520107,I3563,I519813,I520133,);
nor I_30385 (I519781,I520133,I520037);
not I_30386 (I520155,I520133);
nor I_30387 (I520172,I520155,I519946);
nor I_30388 (I520189,I519878,I520172);
DFFARX1 I_30389 (I520189,I3563,I519813,I519796,);
nor I_30390 (I520220,I520155,I520037);
nor I_30391 (I520237,I805821,I805815);
nor I_30392 (I519787,I520237,I520220);
not I_30393 (I520268,I520237);
nand I_30394 (I519790,I519997,I520268);
DFFARX1 I_30395 (I520237,I3563,I519813,I519802,);
DFFARX1 I_30396 (I520237,I3563,I519813,I519799,);
not I_30397 (I520357,I3570);
DFFARX1 I_30398 (I778640,I3563,I520357,I520383,);
DFFARX1 I_30399 (I520383,I3563,I520357,I520400,);
not I_30400 (I520349,I520400);
not I_30401 (I520422,I520383);
nand I_30402 (I520439,I778661,I778652);
and I_30403 (I520456,I520439,I778640);
DFFARX1 I_30404 (I520456,I3563,I520357,I520482,);
not I_30405 (I520490,I520482);
DFFARX1 I_30406 (I778646,I3563,I520357,I520516,);
and I_30407 (I520524,I520516,I778643);
nand I_30408 (I520541,I520516,I778643);
nand I_30409 (I520328,I520490,I520541);
DFFARX1 I_30410 (I778637,I3563,I520357,I520581,);
nor I_30411 (I520589,I520581,I520524);
DFFARX1 I_30412 (I520589,I3563,I520357,I520322,);
nor I_30413 (I520337,I520581,I520482);
nand I_30414 (I520634,I778637,I778649);
and I_30415 (I520651,I520634,I778658);
DFFARX1 I_30416 (I520651,I3563,I520357,I520677,);
nor I_30417 (I520325,I520677,I520581);
not I_30418 (I520699,I520677);
nor I_30419 (I520716,I520699,I520490);
nor I_30420 (I520733,I520422,I520716);
DFFARX1 I_30421 (I520733,I3563,I520357,I520340,);
nor I_30422 (I520764,I520699,I520581);
nor I_30423 (I520781,I778655,I778649);
nor I_30424 (I520331,I520781,I520764);
not I_30425 (I520812,I520781);
nand I_30426 (I520334,I520541,I520812);
DFFARX1 I_30427 (I520781,I3563,I520357,I520346,);
DFFARX1 I_30428 (I520781,I3563,I520357,I520343,);
not I_30429 (I520901,I3570);
DFFARX1 I_30430 (I765346,I3563,I520901,I520927,);
DFFARX1 I_30431 (I520927,I3563,I520901,I520944,);
not I_30432 (I520893,I520944);
not I_30433 (I520966,I520927);
nand I_30434 (I520983,I765367,I765358);
and I_30435 (I521000,I520983,I765346);
DFFARX1 I_30436 (I521000,I3563,I520901,I521026,);
not I_30437 (I521034,I521026);
DFFARX1 I_30438 (I765352,I3563,I520901,I521060,);
and I_30439 (I521068,I521060,I765349);
nand I_30440 (I521085,I521060,I765349);
nand I_30441 (I520872,I521034,I521085);
DFFARX1 I_30442 (I765343,I3563,I520901,I521125,);
nor I_30443 (I521133,I521125,I521068);
DFFARX1 I_30444 (I521133,I3563,I520901,I520866,);
nor I_30445 (I520881,I521125,I521026);
nand I_30446 (I521178,I765343,I765355);
and I_30447 (I521195,I521178,I765364);
DFFARX1 I_30448 (I521195,I3563,I520901,I521221,);
nor I_30449 (I520869,I521221,I521125);
not I_30450 (I521243,I521221);
nor I_30451 (I521260,I521243,I521034);
nor I_30452 (I521277,I520966,I521260);
DFFARX1 I_30453 (I521277,I3563,I520901,I520884,);
nor I_30454 (I521308,I521243,I521125);
nor I_30455 (I521325,I765361,I765355);
nor I_30456 (I520875,I521325,I521308);
not I_30457 (I521356,I521325);
nand I_30458 (I520878,I521085,I521356);
DFFARX1 I_30459 (I521325,I3563,I520901,I520890,);
DFFARX1 I_30460 (I521325,I3563,I520901,I520887,);
not I_30461 (I521445,I3570);
DFFARX1 I_30462 (I31363,I3563,I521445,I521471,);
DFFARX1 I_30463 (I521471,I3563,I521445,I521488,);
not I_30464 (I521437,I521488);
not I_30465 (I521510,I521471);
nand I_30466 (I521527,I31351,I31366);
and I_30467 (I521544,I521527,I31354);
DFFARX1 I_30468 (I521544,I3563,I521445,I521570,);
not I_30469 (I521578,I521570);
DFFARX1 I_30470 (I31375,I3563,I521445,I521604,);
and I_30471 (I521612,I521604,I31369);
nand I_30472 (I521629,I521604,I31369);
nand I_30473 (I521416,I521578,I521629);
DFFARX1 I_30474 (I31372,I3563,I521445,I521669,);
nor I_30475 (I521677,I521669,I521612);
DFFARX1 I_30476 (I521677,I3563,I521445,I521410,);
nor I_30477 (I521425,I521669,I521570);
nand I_30478 (I521722,I31351,I31354);
and I_30479 (I521739,I521722,I31357);
DFFARX1 I_30480 (I521739,I3563,I521445,I521765,);
nor I_30481 (I521413,I521765,I521669);
not I_30482 (I521787,I521765);
nor I_30483 (I521804,I521787,I521578);
nor I_30484 (I521821,I521510,I521804);
DFFARX1 I_30485 (I521821,I3563,I521445,I521428,);
nor I_30486 (I521852,I521787,I521669);
nor I_30487 (I521869,I31360,I31354);
nor I_30488 (I521419,I521869,I521852);
not I_30489 (I521900,I521869);
nand I_30490 (I521422,I521629,I521900);
DFFARX1 I_30491 (I521869,I3563,I521445,I521434,);
DFFARX1 I_30492 (I521869,I3563,I521445,I521431,);
not I_30493 (I521989,I3570);
DFFARX1 I_30494 (I1316093,I3563,I521989,I522015,);
DFFARX1 I_30495 (I522015,I3563,I521989,I522032,);
not I_30496 (I521981,I522032);
not I_30497 (I522054,I522015);
nand I_30498 (I522071,I1316090,I1316087);
and I_30499 (I522088,I522071,I1316075);
DFFARX1 I_30500 (I522088,I3563,I521989,I522114,);
not I_30501 (I522122,I522114);
DFFARX1 I_30502 (I1316099,I3563,I521989,I522148,);
and I_30503 (I522156,I522148,I1316084);
nand I_30504 (I522173,I522148,I1316084);
nand I_30505 (I521960,I522122,I522173);
DFFARX1 I_30506 (I1316078,I3563,I521989,I522213,);
nor I_30507 (I522221,I522213,I522156);
DFFARX1 I_30508 (I522221,I3563,I521989,I521954,);
nor I_30509 (I521969,I522213,I522114);
nand I_30510 (I522266,I1316075,I1316081);
and I_30511 (I522283,I522266,I1316096);
DFFARX1 I_30512 (I522283,I3563,I521989,I522309,);
nor I_30513 (I521957,I522309,I522213);
not I_30514 (I522331,I522309);
nor I_30515 (I522348,I522331,I522122);
nor I_30516 (I522365,I522054,I522348);
DFFARX1 I_30517 (I522365,I3563,I521989,I521972,);
nor I_30518 (I522396,I522331,I522213);
nor I_30519 (I522413,I1316078,I1316081);
nor I_30520 (I521963,I522413,I522396);
not I_30521 (I522444,I522413);
nand I_30522 (I521966,I522173,I522444);
DFFARX1 I_30523 (I522413,I3563,I521989,I521978,);
DFFARX1 I_30524 (I522413,I3563,I521989,I521975,);
not I_30525 (I522533,I3570);
DFFARX1 I_30526 (I135176,I3563,I522533,I522559,);
DFFARX1 I_30527 (I522559,I3563,I522533,I522576,);
not I_30528 (I522525,I522576);
not I_30529 (I522598,I522559);
nand I_30530 (I522615,I135191,I135170);
and I_30531 (I522632,I522615,I135173);
DFFARX1 I_30532 (I522632,I3563,I522533,I522658,);
not I_30533 (I522666,I522658);
DFFARX1 I_30534 (I135179,I3563,I522533,I522692,);
and I_30535 (I522700,I522692,I135173);
nand I_30536 (I522717,I522692,I135173);
nand I_30537 (I522504,I522666,I522717);
DFFARX1 I_30538 (I135188,I3563,I522533,I522757,);
nor I_30539 (I522765,I522757,I522700);
DFFARX1 I_30540 (I522765,I3563,I522533,I522498,);
nor I_30541 (I522513,I522757,I522658);
nand I_30542 (I522810,I135170,I135185);
and I_30543 (I522827,I522810,I135182);
DFFARX1 I_30544 (I522827,I3563,I522533,I522853,);
nor I_30545 (I522501,I522853,I522757);
not I_30546 (I522875,I522853);
nor I_30547 (I522892,I522875,I522666);
nor I_30548 (I522909,I522598,I522892);
DFFARX1 I_30549 (I522909,I3563,I522533,I522516,);
nor I_30550 (I522940,I522875,I522757);
nor I_30551 (I522957,I135194,I135185);
nor I_30552 (I522507,I522957,I522940);
not I_30553 (I522988,I522957);
nand I_30554 (I522510,I522717,I522988);
DFFARX1 I_30555 (I522957,I3563,I522533,I522522,);
DFFARX1 I_30556 (I522957,I3563,I522533,I522519,);
not I_30557 (I523077,I3570);
DFFARX1 I_30558 (I971729,I3563,I523077,I523103,);
DFFARX1 I_30559 (I523103,I3563,I523077,I523120,);
not I_30560 (I523069,I523120);
not I_30561 (I523142,I523103);
nand I_30562 (I523159,I971744,I971732);
and I_30563 (I523176,I523159,I971723);
DFFARX1 I_30564 (I523176,I3563,I523077,I523202,);
not I_30565 (I523210,I523202);
DFFARX1 I_30566 (I971735,I3563,I523077,I523236,);
and I_30567 (I523244,I523236,I971726);
nand I_30568 (I523261,I523236,I971726);
nand I_30569 (I523048,I523210,I523261);
DFFARX1 I_30570 (I971741,I3563,I523077,I523301,);
nor I_30571 (I523309,I523301,I523244);
DFFARX1 I_30572 (I523309,I3563,I523077,I523042,);
nor I_30573 (I523057,I523301,I523202);
nand I_30574 (I523354,I971750,I971738);
and I_30575 (I523371,I523354,I971747);
DFFARX1 I_30576 (I523371,I3563,I523077,I523397,);
nor I_30577 (I523045,I523397,I523301);
not I_30578 (I523419,I523397);
nor I_30579 (I523436,I523419,I523210);
nor I_30580 (I523453,I523142,I523436);
DFFARX1 I_30581 (I523453,I3563,I523077,I523060,);
nor I_30582 (I523484,I523419,I523301);
nor I_30583 (I523501,I971723,I971738);
nor I_30584 (I523051,I523501,I523484);
not I_30585 (I523532,I523501);
nand I_30586 (I523054,I523261,I523532);
DFFARX1 I_30587 (I523501,I3563,I523077,I523066,);
DFFARX1 I_30588 (I523501,I3563,I523077,I523063,);
not I_30589 (I523621,I3570);
DFFARX1 I_30590 (I789622,I3563,I523621,I523647,);
DFFARX1 I_30591 (I523647,I3563,I523621,I523664,);
not I_30592 (I523613,I523664);
not I_30593 (I523686,I523647);
nand I_30594 (I523703,I789643,I789634);
and I_30595 (I523720,I523703,I789622);
DFFARX1 I_30596 (I523720,I3563,I523621,I523746,);
not I_30597 (I523754,I523746);
DFFARX1 I_30598 (I789628,I3563,I523621,I523780,);
and I_30599 (I523788,I523780,I789625);
nand I_30600 (I523805,I523780,I789625);
nand I_30601 (I523592,I523754,I523805);
DFFARX1 I_30602 (I789619,I3563,I523621,I523845,);
nor I_30603 (I523853,I523845,I523788);
DFFARX1 I_30604 (I523853,I3563,I523621,I523586,);
nor I_30605 (I523601,I523845,I523746);
nand I_30606 (I523898,I789619,I789631);
and I_30607 (I523915,I523898,I789640);
DFFARX1 I_30608 (I523915,I3563,I523621,I523941,);
nor I_30609 (I523589,I523941,I523845);
not I_30610 (I523963,I523941);
nor I_30611 (I523980,I523963,I523754);
nor I_30612 (I523997,I523686,I523980);
DFFARX1 I_30613 (I523997,I3563,I523621,I523604,);
nor I_30614 (I524028,I523963,I523845);
nor I_30615 (I524045,I789637,I789631);
nor I_30616 (I523595,I524045,I524028);
not I_30617 (I524076,I524045);
nand I_30618 (I523598,I523805,I524076);
DFFARX1 I_30619 (I524045,I3563,I523621,I523610,);
DFFARX1 I_30620 (I524045,I3563,I523621,I523607,);
not I_30621 (I524165,I3570);
DFFARX1 I_30622 (I1013073,I3563,I524165,I524191,);
DFFARX1 I_30623 (I524191,I3563,I524165,I524208,);
not I_30624 (I524157,I524208);
not I_30625 (I524230,I524191);
nand I_30626 (I524247,I1013088,I1013076);
and I_30627 (I524264,I524247,I1013067);
DFFARX1 I_30628 (I524264,I3563,I524165,I524290,);
not I_30629 (I524298,I524290);
DFFARX1 I_30630 (I1013079,I3563,I524165,I524324,);
and I_30631 (I524332,I524324,I1013070);
nand I_30632 (I524349,I524324,I1013070);
nand I_30633 (I524136,I524298,I524349);
DFFARX1 I_30634 (I1013085,I3563,I524165,I524389,);
nor I_30635 (I524397,I524389,I524332);
DFFARX1 I_30636 (I524397,I3563,I524165,I524130,);
nor I_30637 (I524145,I524389,I524290);
nand I_30638 (I524442,I1013094,I1013082);
and I_30639 (I524459,I524442,I1013091);
DFFARX1 I_30640 (I524459,I3563,I524165,I524485,);
nor I_30641 (I524133,I524485,I524389);
not I_30642 (I524507,I524485);
nor I_30643 (I524524,I524507,I524298);
nor I_30644 (I524541,I524230,I524524);
DFFARX1 I_30645 (I524541,I3563,I524165,I524148,);
nor I_30646 (I524572,I524507,I524389);
nor I_30647 (I524589,I1013067,I1013082);
nor I_30648 (I524139,I524589,I524572);
not I_30649 (I524620,I524589);
nand I_30650 (I524142,I524349,I524620);
DFFARX1 I_30651 (I524589,I3563,I524165,I524154,);
DFFARX1 I_30652 (I524589,I3563,I524165,I524151,);
not I_30653 (I524709,I3570);
DFFARX1 I_30654 (I189307,I3563,I524709,I524735,);
DFFARX1 I_30655 (I524735,I3563,I524709,I524752,);
not I_30656 (I524701,I524752);
not I_30657 (I524774,I524735);
nand I_30658 (I524791,I189319,I189298);
and I_30659 (I524808,I524791,I189301);
DFFARX1 I_30660 (I524808,I3563,I524709,I524834,);
not I_30661 (I524842,I524834);
DFFARX1 I_30662 (I189310,I3563,I524709,I524868,);
and I_30663 (I524876,I524868,I189322);
nand I_30664 (I524893,I524868,I189322);
nand I_30665 (I524680,I524842,I524893);
DFFARX1 I_30666 (I189316,I3563,I524709,I524933,);
nor I_30667 (I524941,I524933,I524876);
DFFARX1 I_30668 (I524941,I3563,I524709,I524674,);
nor I_30669 (I524689,I524933,I524834);
nand I_30670 (I524986,I189304,I189301);
and I_30671 (I525003,I524986,I189313);
DFFARX1 I_30672 (I525003,I3563,I524709,I525029,);
nor I_30673 (I524677,I525029,I524933);
not I_30674 (I525051,I525029);
nor I_30675 (I525068,I525051,I524842);
nor I_30676 (I525085,I524774,I525068);
DFFARX1 I_30677 (I525085,I3563,I524709,I524692,);
nor I_30678 (I525116,I525051,I524933);
nor I_30679 (I525133,I189298,I189301);
nor I_30680 (I524683,I525133,I525116);
not I_30681 (I525164,I525133);
nand I_30682 (I524686,I524893,I525164);
DFFARX1 I_30683 (I525133,I3563,I524709,I524698,);
DFFARX1 I_30684 (I525133,I3563,I524709,I524695,);
not I_30685 (I525253,I3570);
DFFARX1 I_30686 (I837945,I3563,I525253,I525279,);
DFFARX1 I_30687 (I525279,I3563,I525253,I525296,);
not I_30688 (I525245,I525296);
not I_30689 (I525318,I525279);
nand I_30690 (I525335,I837939,I837936);
and I_30691 (I525352,I525335,I837951);
DFFARX1 I_30692 (I525352,I3563,I525253,I525378,);
not I_30693 (I525386,I525378);
DFFARX1 I_30694 (I837939,I3563,I525253,I525412,);
and I_30695 (I525420,I525412,I837933);
nand I_30696 (I525437,I525412,I837933);
nand I_30697 (I525224,I525386,I525437);
DFFARX1 I_30698 (I837933,I3563,I525253,I525477,);
nor I_30699 (I525485,I525477,I525420);
DFFARX1 I_30700 (I525485,I3563,I525253,I525218,);
nor I_30701 (I525233,I525477,I525378);
nand I_30702 (I525530,I837948,I837942);
and I_30703 (I525547,I525530,I837936);
DFFARX1 I_30704 (I525547,I3563,I525253,I525573,);
nor I_30705 (I525221,I525573,I525477);
not I_30706 (I525595,I525573);
nor I_30707 (I525612,I525595,I525386);
nor I_30708 (I525629,I525318,I525612);
DFFARX1 I_30709 (I525629,I3563,I525253,I525236,);
nor I_30710 (I525660,I525595,I525477);
nor I_30711 (I525677,I837954,I837942);
nor I_30712 (I525227,I525677,I525660);
not I_30713 (I525708,I525677);
nand I_30714 (I525230,I525437,I525708);
DFFARX1 I_30715 (I525677,I3563,I525253,I525242,);
DFFARX1 I_30716 (I525677,I3563,I525253,I525239,);
not I_30717 (I525797,I3570);
DFFARX1 I_30718 (I881686,I3563,I525797,I525823,);
DFFARX1 I_30719 (I525823,I3563,I525797,I525840,);
not I_30720 (I525789,I525840);
not I_30721 (I525862,I525823);
nand I_30722 (I525879,I881680,I881677);
and I_30723 (I525896,I525879,I881692);
DFFARX1 I_30724 (I525896,I3563,I525797,I525922,);
not I_30725 (I525930,I525922);
DFFARX1 I_30726 (I881680,I3563,I525797,I525956,);
and I_30727 (I525964,I525956,I881674);
nand I_30728 (I525981,I525956,I881674);
nand I_30729 (I525768,I525930,I525981);
DFFARX1 I_30730 (I881674,I3563,I525797,I526021,);
nor I_30731 (I526029,I526021,I525964);
DFFARX1 I_30732 (I526029,I3563,I525797,I525762,);
nor I_30733 (I525777,I526021,I525922);
nand I_30734 (I526074,I881689,I881683);
and I_30735 (I526091,I526074,I881677);
DFFARX1 I_30736 (I526091,I3563,I525797,I526117,);
nor I_30737 (I525765,I526117,I526021);
not I_30738 (I526139,I526117);
nor I_30739 (I526156,I526139,I525930);
nor I_30740 (I526173,I525862,I526156);
DFFARX1 I_30741 (I526173,I3563,I525797,I525780,);
nor I_30742 (I526204,I526139,I526021);
nor I_30743 (I526221,I881695,I881683);
nor I_30744 (I525771,I526221,I526204);
not I_30745 (I526252,I526221);
nand I_30746 (I525774,I525981,I526252);
DFFARX1 I_30747 (I526221,I3563,I525797,I525786,);
DFFARX1 I_30748 (I526221,I3563,I525797,I525783,);
not I_30749 (I526338,I3570);
DFFARX1 I_30750 (I862711,I3563,I526338,I526364,);
DFFARX1 I_30751 (I526364,I3563,I526338,I526381,);
not I_30752 (I526330,I526381);
DFFARX1 I_30753 (I862708,I3563,I526338,I526412,);
not I_30754 (I526420,I862708);
nor I_30755 (I526437,I526364,I526420);
not I_30756 (I526454,I862705);
not I_30757 (I526471,I862720);
nand I_30758 (I526488,I526471,I862705);
nor I_30759 (I526505,I526420,I526488);
nor I_30760 (I526522,I526412,I526505);
DFFARX1 I_30761 (I526471,I3563,I526338,I526327,);
nor I_30762 (I526553,I862720,I862714);
nand I_30763 (I526570,I526553,I862702);
nor I_30764 (I526587,I526570,I526454);
nand I_30765 (I526312,I526587,I862708);
DFFARX1 I_30766 (I526570,I3563,I526338,I526324,);
nand I_30767 (I526632,I526454,I862720);
nor I_30768 (I526649,I526454,I862720);
nand I_30769 (I526318,I526437,I526649);
not I_30770 (I526680,I862723);
nor I_30771 (I526697,I526680,I526632);
DFFARX1 I_30772 (I526697,I3563,I526338,I526306,);
nor I_30773 (I526728,I526680,I862702);
and I_30774 (I526745,I526728,I862717);
or I_30775 (I526762,I526745,I862705);
DFFARX1 I_30776 (I526762,I3563,I526338,I526788,);
nor I_30777 (I526796,I526788,I526412);
nor I_30778 (I526315,I526364,I526796);
not I_30779 (I526827,I526788);
nor I_30780 (I526844,I526827,I526522);
DFFARX1 I_30781 (I526844,I3563,I526338,I526321,);
nand I_30782 (I526875,I526827,I526454);
nor I_30783 (I526309,I526680,I526875);
not I_30784 (I526933,I3570);
DFFARX1 I_30785 (I837415,I3563,I526933,I526959,);
DFFARX1 I_30786 (I526959,I3563,I526933,I526976,);
not I_30787 (I526925,I526976);
DFFARX1 I_30788 (I837412,I3563,I526933,I527007,);
not I_30789 (I527015,I837412);
nor I_30790 (I527032,I526959,I527015);
not I_30791 (I527049,I837409);
not I_30792 (I527066,I837424);
nand I_30793 (I527083,I527066,I837409);
nor I_30794 (I527100,I527015,I527083);
nor I_30795 (I527117,I527007,I527100);
DFFARX1 I_30796 (I527066,I3563,I526933,I526922,);
nor I_30797 (I527148,I837424,I837418);
nand I_30798 (I527165,I527148,I837406);
nor I_30799 (I527182,I527165,I527049);
nand I_30800 (I526907,I527182,I837412);
DFFARX1 I_30801 (I527165,I3563,I526933,I526919,);
nand I_30802 (I527227,I527049,I837424);
nor I_30803 (I527244,I527049,I837424);
nand I_30804 (I526913,I527032,I527244);
not I_30805 (I527275,I837427);
nor I_30806 (I527292,I527275,I527227);
DFFARX1 I_30807 (I527292,I3563,I526933,I526901,);
nor I_30808 (I527323,I527275,I837406);
and I_30809 (I527340,I527323,I837421);
or I_30810 (I527357,I527340,I837409);
DFFARX1 I_30811 (I527357,I3563,I526933,I527383,);
nor I_30812 (I527391,I527383,I527007);
nor I_30813 (I526910,I526959,I527391);
not I_30814 (I527422,I527383);
nor I_30815 (I527439,I527422,I527117);
DFFARX1 I_30816 (I527439,I3563,I526933,I526916,);
nand I_30817 (I527470,I527422,I527049);
nor I_30818 (I526904,I527275,I527470);
not I_30819 (I527528,I3570);
DFFARX1 I_30820 (I679230,I3563,I527528,I527554,);
DFFARX1 I_30821 (I527554,I3563,I527528,I527571,);
not I_30822 (I527520,I527571);
DFFARX1 I_30823 (I679224,I3563,I527528,I527602,);
not I_30824 (I527610,I679221);
nor I_30825 (I527627,I527554,I527610);
not I_30826 (I527644,I679233);
not I_30827 (I527661,I679236);
nand I_30828 (I527678,I527661,I679233);
nor I_30829 (I527695,I527610,I527678);
nor I_30830 (I527712,I527602,I527695);
DFFARX1 I_30831 (I527661,I3563,I527528,I527517,);
nor I_30832 (I527743,I679236,I679245);
nand I_30833 (I527760,I527743,I679239);
nor I_30834 (I527777,I527760,I527644);
nand I_30835 (I527502,I527777,I679221);
DFFARX1 I_30836 (I527760,I3563,I527528,I527514,);
nand I_30837 (I527822,I527644,I679236);
nor I_30838 (I527839,I527644,I679236);
nand I_30839 (I527508,I527627,I527839);
not I_30840 (I527870,I679227);
nor I_30841 (I527887,I527870,I527822);
DFFARX1 I_30842 (I527887,I3563,I527528,I527496,);
nor I_30843 (I527918,I527870,I679242);
and I_30844 (I527935,I527918,I679221);
or I_30845 (I527952,I527935,I679224);
DFFARX1 I_30846 (I527952,I3563,I527528,I527978,);
nor I_30847 (I527986,I527978,I527602);
nor I_30848 (I527505,I527554,I527986);
not I_30849 (I528017,I527978);
nor I_30850 (I528034,I528017,I527712);
DFFARX1 I_30851 (I528034,I3563,I527528,I527511,);
nand I_30852 (I528065,I528017,I527644);
nor I_30853 (I527499,I527870,I528065);
not I_30854 (I528123,I3570);
DFFARX1 I_30855 (I197628,I3563,I528123,I528149,);
DFFARX1 I_30856 (I528149,I3563,I528123,I528166,);
not I_30857 (I528115,I528166);
DFFARX1 I_30858 (I197652,I3563,I528123,I528197,);
not I_30859 (I528205,I197646);
nor I_30860 (I528222,I528149,I528205);
not I_30861 (I528239,I197640);
not I_30862 (I528256,I197637);
nand I_30863 (I528273,I528256,I197640);
nor I_30864 (I528290,I528205,I528273);
nor I_30865 (I528307,I528197,I528290);
DFFARX1 I_30866 (I528256,I3563,I528123,I528112,);
nor I_30867 (I528338,I197637,I197631);
nand I_30868 (I528355,I528338,I197649);
nor I_30869 (I528372,I528355,I528239);
nand I_30870 (I528097,I528372,I197646);
DFFARX1 I_30871 (I528355,I3563,I528123,I528109,);
nand I_30872 (I528417,I528239,I197637);
nor I_30873 (I528434,I528239,I197637);
nand I_30874 (I528103,I528222,I528434);
not I_30875 (I528465,I197643);
nor I_30876 (I528482,I528465,I528417);
DFFARX1 I_30877 (I528482,I3563,I528123,I528091,);
nor I_30878 (I528513,I528465,I197628);
and I_30879 (I528530,I528513,I197634);
or I_30880 (I528547,I528530,I197631);
DFFARX1 I_30881 (I528547,I3563,I528123,I528573,);
nor I_30882 (I528581,I528573,I528197);
nor I_30883 (I528100,I528149,I528581);
not I_30884 (I528612,I528573);
nor I_30885 (I528629,I528612,I528307);
DFFARX1 I_30886 (I528629,I3563,I528123,I528106,);
nand I_30887 (I528660,I528612,I528239);
nor I_30888 (I528094,I528465,I528660);
not I_30889 (I528718,I3570);
DFFARX1 I_30890 (I835834,I3563,I528718,I528744,);
DFFARX1 I_30891 (I528744,I3563,I528718,I528761,);
not I_30892 (I528710,I528761);
DFFARX1 I_30893 (I835831,I3563,I528718,I528792,);
not I_30894 (I528800,I835831);
nor I_30895 (I528817,I528744,I528800);
not I_30896 (I528834,I835828);
not I_30897 (I528851,I835843);
nand I_30898 (I528868,I528851,I835828);
nor I_30899 (I528885,I528800,I528868);
nor I_30900 (I528902,I528792,I528885);
DFFARX1 I_30901 (I528851,I3563,I528718,I528707,);
nor I_30902 (I528933,I835843,I835837);
nand I_30903 (I528950,I528933,I835825);
nor I_30904 (I528967,I528950,I528834);
nand I_30905 (I528692,I528967,I835831);
DFFARX1 I_30906 (I528950,I3563,I528718,I528704,);
nand I_30907 (I529012,I528834,I835843);
nor I_30908 (I529029,I528834,I835843);
nand I_30909 (I528698,I528817,I529029);
not I_30910 (I529060,I835846);
nor I_30911 (I529077,I529060,I529012);
DFFARX1 I_30912 (I529077,I3563,I528718,I528686,);
nor I_30913 (I529108,I529060,I835825);
and I_30914 (I529125,I529108,I835840);
or I_30915 (I529142,I529125,I835828);
DFFARX1 I_30916 (I529142,I3563,I528718,I529168,);
nor I_30917 (I529176,I529168,I528792);
nor I_30918 (I528695,I528744,I529176);
not I_30919 (I529207,I529168);
nor I_30920 (I529224,I529207,I528902);
DFFARX1 I_30921 (I529224,I3563,I528718,I528701,);
nand I_30922 (I529255,I529207,I528834);
nor I_30923 (I528689,I529060,I529255);
not I_30924 (I529313,I3570);
DFFARX1 I_30925 (I410806,I3563,I529313,I529339,);
DFFARX1 I_30926 (I529339,I3563,I529313,I529356,);
not I_30927 (I529305,I529356);
DFFARX1 I_30928 (I410794,I3563,I529313,I529387,);
not I_30929 (I529395,I410797);
nor I_30930 (I529412,I529339,I529395);
not I_30931 (I529429,I410800);
not I_30932 (I529446,I410812);
nand I_30933 (I529463,I529446,I410800);
nor I_30934 (I529480,I529395,I529463);
nor I_30935 (I529497,I529387,I529480);
DFFARX1 I_30936 (I529446,I3563,I529313,I529302,);
nor I_30937 (I529528,I410812,I410803);
nand I_30938 (I529545,I529528,I410791);
nor I_30939 (I529562,I529545,I529429);
nand I_30940 (I529287,I529562,I410797);
DFFARX1 I_30941 (I529545,I3563,I529313,I529299,);
nand I_30942 (I529607,I529429,I410812);
nor I_30943 (I529624,I529429,I410812);
nand I_30944 (I529293,I529412,I529624);
not I_30945 (I529655,I410809);
nor I_30946 (I529672,I529655,I529607);
DFFARX1 I_30947 (I529672,I3563,I529313,I529281,);
nor I_30948 (I529703,I529655,I410815);
and I_30949 (I529720,I529703,I410818);
or I_30950 (I529737,I529720,I410791);
DFFARX1 I_30951 (I529737,I3563,I529313,I529763,);
nor I_30952 (I529771,I529763,I529387);
nor I_30953 (I529290,I529339,I529771);
not I_30954 (I529802,I529763);
nor I_30955 (I529819,I529802,I529497);
DFFARX1 I_30956 (I529819,I3563,I529313,I529296,);
nand I_30957 (I529850,I529802,I529429);
nor I_30958 (I529284,I529655,I529850);
not I_30959 (I529908,I3570);
DFFARX1 I_30960 (I1387458,I3563,I529908,I529934,);
DFFARX1 I_30961 (I529934,I3563,I529908,I529951,);
not I_30962 (I529900,I529951);
DFFARX1 I_30963 (I1387464,I3563,I529908,I529982,);
not I_30964 (I529990,I1387479);
nor I_30965 (I530007,I529934,I529990);
not I_30966 (I530024,I1387470);
not I_30967 (I530041,I1387467);
nand I_30968 (I530058,I530041,I1387470);
nor I_30969 (I530075,I529990,I530058);
nor I_30970 (I530092,I529982,I530075);
DFFARX1 I_30971 (I530041,I3563,I529908,I529897,);
nor I_30972 (I530123,I1387467,I1387458);
nand I_30973 (I530140,I530123,I1387482);
nor I_30974 (I530157,I530140,I530024);
nand I_30975 (I529882,I530157,I1387479);
DFFARX1 I_30976 (I530140,I3563,I529908,I529894,);
nand I_30977 (I530202,I530024,I1387467);
nor I_30978 (I530219,I530024,I1387467);
nand I_30979 (I529888,I530007,I530219);
not I_30980 (I530250,I1387476);
nor I_30981 (I530267,I530250,I530202);
DFFARX1 I_30982 (I530267,I3563,I529908,I529876,);
nor I_30983 (I530298,I530250,I1387461);
and I_30984 (I530315,I530298,I1387473);
or I_30985 (I530332,I530315,I1387485);
DFFARX1 I_30986 (I530332,I3563,I529908,I530358,);
nor I_30987 (I530366,I530358,I529982);
nor I_30988 (I529885,I529934,I530366);
not I_30989 (I530397,I530358);
nor I_30990 (I530414,I530397,I530092);
DFFARX1 I_30991 (I530414,I3563,I529908,I529891,);
nand I_30992 (I530445,I530397,I530024);
nor I_30993 (I529879,I530250,I530445);
not I_30994 (I530503,I3570);
DFFARX1 I_30995 (I599460,I3563,I530503,I530529,);
DFFARX1 I_30996 (I530529,I3563,I530503,I530546,);
not I_30997 (I530495,I530546);
DFFARX1 I_30998 (I599472,I3563,I530503,I530577,);
not I_30999 (I530585,I599457);
nor I_31000 (I530602,I530529,I530585);
not I_31001 (I530619,I599475);
not I_31002 (I530636,I599466);
nand I_31003 (I530653,I530636,I599475);
nor I_31004 (I530670,I530585,I530653);
nor I_31005 (I530687,I530577,I530670);
DFFARX1 I_31006 (I530636,I3563,I530503,I530492,);
nor I_31007 (I530718,I599466,I599478);
nand I_31008 (I530735,I530718,I599481);
nor I_31009 (I530752,I530735,I530619);
nand I_31010 (I530477,I530752,I599457);
DFFARX1 I_31011 (I530735,I3563,I530503,I530489,);
nand I_31012 (I530797,I530619,I599466);
nor I_31013 (I530814,I530619,I599466);
nand I_31014 (I530483,I530602,I530814);
not I_31015 (I530845,I599457);
nor I_31016 (I530862,I530845,I530797);
DFFARX1 I_31017 (I530862,I3563,I530503,I530471,);
nor I_31018 (I530893,I530845,I599469);
and I_31019 (I530910,I530893,I599463);
or I_31020 (I530927,I530910,I599460);
DFFARX1 I_31021 (I530927,I3563,I530503,I530953,);
nor I_31022 (I530961,I530953,I530577);
nor I_31023 (I530480,I530529,I530961);
not I_31024 (I530992,I530953);
nor I_31025 (I531009,I530992,I530687);
DFFARX1 I_31026 (I531009,I3563,I530503,I530486,);
nand I_31027 (I531040,I530992,I530619);
nor I_31028 (I530474,I530845,I531040);
not I_31029 (I531098,I3570);
DFFARX1 I_31030 (I313311,I3563,I531098,I531124,);
DFFARX1 I_31031 (I531124,I3563,I531098,I531141,);
not I_31032 (I531090,I531141);
DFFARX1 I_31033 (I313299,I3563,I531098,I531172,);
not I_31034 (I531180,I313302);
nor I_31035 (I531197,I531124,I531180);
not I_31036 (I531214,I313305);
not I_31037 (I531231,I313317);
nand I_31038 (I531248,I531231,I313305);
nor I_31039 (I531265,I531180,I531248);
nor I_31040 (I531282,I531172,I531265);
DFFARX1 I_31041 (I531231,I3563,I531098,I531087,);
nor I_31042 (I531313,I313317,I313308);
nand I_31043 (I531330,I531313,I313296);
nor I_31044 (I531347,I531330,I531214);
nand I_31045 (I531072,I531347,I313302);
DFFARX1 I_31046 (I531330,I3563,I531098,I531084,);
nand I_31047 (I531392,I531214,I313317);
nor I_31048 (I531409,I531214,I313317);
nand I_31049 (I531078,I531197,I531409);
not I_31050 (I531440,I313314);
nor I_31051 (I531457,I531440,I531392);
DFFARX1 I_31052 (I531457,I3563,I531098,I531066,);
nor I_31053 (I531488,I531440,I313320);
and I_31054 (I531505,I531488,I313323);
or I_31055 (I531522,I531505,I313296);
DFFARX1 I_31056 (I531522,I3563,I531098,I531548,);
nor I_31057 (I531556,I531548,I531172);
nor I_31058 (I531075,I531124,I531556);
not I_31059 (I531587,I531548);
nor I_31060 (I531604,I531587,I531282);
DFFARX1 I_31061 (I531604,I3563,I531098,I531081,);
nand I_31062 (I531635,I531587,I531214);
nor I_31063 (I531069,I531440,I531635);
not I_31064 (I531693,I3570);
DFFARX1 I_31065 (I397104,I3563,I531693,I531719,);
DFFARX1 I_31066 (I531719,I3563,I531693,I531736,);
not I_31067 (I531685,I531736);
DFFARX1 I_31068 (I397092,I3563,I531693,I531767,);
not I_31069 (I531775,I397095);
nor I_31070 (I531792,I531719,I531775);
not I_31071 (I531809,I397098);
not I_31072 (I531826,I397110);
nand I_31073 (I531843,I531826,I397098);
nor I_31074 (I531860,I531775,I531843);
nor I_31075 (I531877,I531767,I531860);
DFFARX1 I_31076 (I531826,I3563,I531693,I531682,);
nor I_31077 (I531908,I397110,I397101);
nand I_31078 (I531925,I531908,I397089);
nor I_31079 (I531942,I531925,I531809);
nand I_31080 (I531667,I531942,I397095);
DFFARX1 I_31081 (I531925,I3563,I531693,I531679,);
nand I_31082 (I531987,I531809,I397110);
nor I_31083 (I532004,I531809,I397110);
nand I_31084 (I531673,I531792,I532004);
not I_31085 (I532035,I397107);
nor I_31086 (I532052,I532035,I531987);
DFFARX1 I_31087 (I532052,I3563,I531693,I531661,);
nor I_31088 (I532083,I532035,I397113);
and I_31089 (I532100,I532083,I397116);
or I_31090 (I532117,I532100,I397089);
DFFARX1 I_31091 (I532117,I3563,I531693,I532143,);
nor I_31092 (I532151,I532143,I531767);
nor I_31093 (I531670,I531719,I532151);
not I_31094 (I532182,I532143);
nor I_31095 (I532199,I532182,I531877);
DFFARX1 I_31096 (I532199,I3563,I531693,I531676,);
nand I_31097 (I532230,I532182,I531809);
nor I_31098 (I531664,I532035,I532230);
not I_31099 (I532288,I3570);
DFFARX1 I_31100 (I1136675,I3563,I532288,I532314,);
DFFARX1 I_31101 (I532314,I3563,I532288,I532331,);
not I_31102 (I532280,I532331);
DFFARX1 I_31103 (I1136657,I3563,I532288,I532362,);
not I_31104 (I532370,I1136663);
nor I_31105 (I532387,I532314,I532370);
not I_31106 (I532404,I1136678);
not I_31107 (I532421,I1136669);
nand I_31108 (I532438,I532421,I1136678);
nor I_31109 (I532455,I532370,I532438);
nor I_31110 (I532472,I532362,I532455);
DFFARX1 I_31111 (I532421,I3563,I532288,I532277,);
nor I_31112 (I532503,I1136669,I1136681);
nand I_31113 (I532520,I532503,I1136660);
nor I_31114 (I532537,I532520,I532404);
nand I_31115 (I532262,I532537,I1136663);
DFFARX1 I_31116 (I532520,I3563,I532288,I532274,);
nand I_31117 (I532582,I532404,I1136669);
nor I_31118 (I532599,I532404,I1136669);
nand I_31119 (I532268,I532387,I532599);
not I_31120 (I532630,I1136666);
nor I_31121 (I532647,I532630,I532582);
DFFARX1 I_31122 (I532647,I3563,I532288,I532256,);
nor I_31123 (I532678,I532630,I1136672);
and I_31124 (I532695,I532678,I1136657);
or I_31125 (I532712,I532695,I1136660);
DFFARX1 I_31126 (I532712,I3563,I532288,I532738,);
nor I_31127 (I532746,I532738,I532362);
nor I_31128 (I532265,I532314,I532746);
not I_31129 (I532777,I532738);
nor I_31130 (I532794,I532777,I532472);
DFFARX1 I_31131 (I532794,I3563,I532288,I532271,);
nand I_31132 (I532825,I532777,I532404);
nor I_31133 (I532259,I532630,I532825);
not I_31134 (I532883,I3570);
DFFARX1 I_31135 (I81425,I3563,I532883,I532909,);
DFFARX1 I_31136 (I532909,I3563,I532883,I532926,);
not I_31137 (I532875,I532926);
DFFARX1 I_31138 (I81437,I3563,I532883,I532957,);
not I_31139 (I532965,I81428);
nor I_31140 (I532982,I532909,I532965);
not I_31141 (I532999,I81419);
not I_31142 (I533016,I81416);
nand I_31143 (I533033,I533016,I81419);
nor I_31144 (I533050,I532965,I533033);
nor I_31145 (I533067,I532957,I533050);
DFFARX1 I_31146 (I533016,I3563,I532883,I532872,);
nor I_31147 (I533098,I81416,I81416);
nand I_31148 (I533115,I533098,I81434);
nor I_31149 (I533132,I533115,I532999);
nand I_31150 (I532857,I533132,I81428);
DFFARX1 I_31151 (I533115,I3563,I532883,I532869,);
nand I_31152 (I533177,I532999,I81416);
nor I_31153 (I533194,I532999,I81416);
nand I_31154 (I532863,I532982,I533194);
not I_31155 (I533225,I81440);
nor I_31156 (I533242,I533225,I533177);
DFFARX1 I_31157 (I533242,I3563,I532883,I532851,);
nor I_31158 (I533273,I533225,I81419);
and I_31159 (I533290,I533273,I81422);
or I_31160 (I533307,I533290,I81431);
DFFARX1 I_31161 (I533307,I3563,I532883,I533333,);
nor I_31162 (I533341,I533333,I532957);
nor I_31163 (I532860,I532909,I533341);
not I_31164 (I533372,I533333);
nor I_31165 (I533389,I533372,I533067);
DFFARX1 I_31166 (I533389,I3563,I532883,I532866,);
nand I_31167 (I533420,I533372,I532999);
nor I_31168 (I532854,I533225,I533420);
not I_31169 (I533478,I3570);
DFFARX1 I_31170 (I900655,I3563,I533478,I533504,);
DFFARX1 I_31171 (I533504,I3563,I533478,I533521,);
not I_31172 (I533470,I533521);
DFFARX1 I_31173 (I900652,I3563,I533478,I533552,);
not I_31174 (I533560,I900652);
nor I_31175 (I533577,I533504,I533560);
not I_31176 (I533594,I900649);
not I_31177 (I533611,I900664);
nand I_31178 (I533628,I533611,I900649);
nor I_31179 (I533645,I533560,I533628);
nor I_31180 (I533662,I533552,I533645);
DFFARX1 I_31181 (I533611,I3563,I533478,I533467,);
nor I_31182 (I533693,I900664,I900658);
nand I_31183 (I533710,I533693,I900646);
nor I_31184 (I533727,I533710,I533594);
nand I_31185 (I533452,I533727,I900652);
DFFARX1 I_31186 (I533710,I3563,I533478,I533464,);
nand I_31187 (I533772,I533594,I900664);
nor I_31188 (I533789,I533594,I900664);
nand I_31189 (I533458,I533577,I533789);
not I_31190 (I533820,I900667);
nor I_31191 (I533837,I533820,I533772);
DFFARX1 I_31192 (I533837,I3563,I533478,I533446,);
nor I_31193 (I533868,I533820,I900646);
and I_31194 (I533885,I533868,I900661);
or I_31195 (I533902,I533885,I900649);
DFFARX1 I_31196 (I533902,I3563,I533478,I533928,);
nor I_31197 (I533936,I533928,I533552);
nor I_31198 (I533455,I533504,I533936);
not I_31199 (I533967,I533928);
nor I_31200 (I533984,I533967,I533662);
DFFARX1 I_31201 (I533984,I3563,I533478,I533461,);
nand I_31202 (I534015,I533967,I533594);
nor I_31203 (I533449,I533820,I534015);
not I_31204 (I534073,I3570);
DFFARX1 I_31205 (I1103151,I3563,I534073,I534099,);
DFFARX1 I_31206 (I534099,I3563,I534073,I534116,);
not I_31207 (I534065,I534116);
DFFARX1 I_31208 (I1103133,I3563,I534073,I534147,);
not I_31209 (I534155,I1103139);
nor I_31210 (I534172,I534099,I534155);
not I_31211 (I534189,I1103154);
not I_31212 (I534206,I1103145);
nand I_31213 (I534223,I534206,I1103154);
nor I_31214 (I534240,I534155,I534223);
nor I_31215 (I534257,I534147,I534240);
DFFARX1 I_31216 (I534206,I3563,I534073,I534062,);
nor I_31217 (I534288,I1103145,I1103157);
nand I_31218 (I534305,I534288,I1103136);
nor I_31219 (I534322,I534305,I534189);
nand I_31220 (I534047,I534322,I1103139);
DFFARX1 I_31221 (I534305,I3563,I534073,I534059,);
nand I_31222 (I534367,I534189,I1103145);
nor I_31223 (I534384,I534189,I1103145);
nand I_31224 (I534053,I534172,I534384);
not I_31225 (I534415,I1103142);
nor I_31226 (I534432,I534415,I534367);
DFFARX1 I_31227 (I534432,I3563,I534073,I534041,);
nor I_31228 (I534463,I534415,I1103148);
and I_31229 (I534480,I534463,I1103133);
or I_31230 (I534497,I534480,I1103136);
DFFARX1 I_31231 (I534497,I3563,I534073,I534523,);
nor I_31232 (I534531,I534523,I534147);
nor I_31233 (I534050,I534099,I534531);
not I_31234 (I534562,I534523);
nor I_31235 (I534579,I534562,I534257);
DFFARX1 I_31236 (I534579,I3563,I534073,I534056,);
nand I_31237 (I534610,I534562,I534189);
nor I_31238 (I534044,I534415,I534610);
not I_31239 (I534668,I3570);
DFFARX1 I_31240 (I514882,I3563,I534668,I534694,);
DFFARX1 I_31241 (I534694,I3563,I534668,I534711,);
not I_31242 (I534660,I534711);
DFFARX1 I_31243 (I514906,I3563,I534668,I534742,);
not I_31244 (I534750,I514885);
nor I_31245 (I534767,I534694,I534750);
not I_31246 (I534784,I514891);
not I_31247 (I534801,I514897);
nand I_31248 (I534818,I534801,I514891);
nor I_31249 (I534835,I534750,I534818);
nor I_31250 (I534852,I534742,I534835);
DFFARX1 I_31251 (I534801,I3563,I534668,I534657,);
nor I_31252 (I534883,I514897,I514909);
nand I_31253 (I534900,I534883,I514903);
nor I_31254 (I534917,I534900,I534784);
nand I_31255 (I534642,I534917,I514885);
DFFARX1 I_31256 (I534900,I3563,I534668,I534654,);
nand I_31257 (I534962,I534784,I514897);
nor I_31258 (I534979,I534784,I514897);
nand I_31259 (I534648,I534767,I534979);
not I_31260 (I535010,I514888);
nor I_31261 (I535027,I535010,I534962);
DFFARX1 I_31262 (I535027,I3563,I534668,I534636,);
nor I_31263 (I535058,I535010,I514882);
and I_31264 (I535075,I535058,I514900);
or I_31265 (I535092,I535075,I514894);
DFFARX1 I_31266 (I535092,I3563,I534668,I535118,);
nor I_31267 (I535126,I535118,I534742);
nor I_31268 (I534645,I534694,I535126);
not I_31269 (I535157,I535118);
nor I_31270 (I535174,I535157,I534852);
DFFARX1 I_31271 (I535174,I3563,I534668,I534651,);
nand I_31272 (I535205,I535157,I534784);
nor I_31273 (I534639,I535010,I535205);
not I_31274 (I535263,I3570);
DFFARX1 I_31275 (I370754,I3563,I535263,I535289,);
DFFARX1 I_31276 (I535289,I3563,I535263,I535306,);
not I_31277 (I535255,I535306);
DFFARX1 I_31278 (I370742,I3563,I535263,I535337,);
not I_31279 (I535345,I370745);
nor I_31280 (I535362,I535289,I535345);
not I_31281 (I535379,I370748);
not I_31282 (I535396,I370760);
nand I_31283 (I535413,I535396,I370748);
nor I_31284 (I535430,I535345,I535413);
nor I_31285 (I535447,I535337,I535430);
DFFARX1 I_31286 (I535396,I3563,I535263,I535252,);
nor I_31287 (I535478,I370760,I370751);
nand I_31288 (I535495,I535478,I370739);
nor I_31289 (I535512,I535495,I535379);
nand I_31290 (I535237,I535512,I370745);
DFFARX1 I_31291 (I535495,I3563,I535263,I535249,);
nand I_31292 (I535557,I535379,I370760);
nor I_31293 (I535574,I535379,I370760);
nand I_31294 (I535243,I535362,I535574);
not I_31295 (I535605,I370757);
nor I_31296 (I535622,I535605,I535557);
DFFARX1 I_31297 (I535622,I3563,I535263,I535231,);
nor I_31298 (I535653,I535605,I370763);
and I_31299 (I535670,I535653,I370766);
or I_31300 (I535687,I535670,I370739);
DFFARX1 I_31301 (I535687,I3563,I535263,I535713,);
nor I_31302 (I535721,I535713,I535337);
nor I_31303 (I535240,I535289,I535721);
not I_31304 (I535752,I535713);
nor I_31305 (I535769,I535752,I535447);
DFFARX1 I_31306 (I535769,I3563,I535263,I535246,);
nand I_31307 (I535800,I535752,I535379);
nor I_31308 (I535234,I535605,I535800);
not I_31309 (I535858,I3570);
DFFARX1 I_31310 (I220833,I3563,I535858,I535884,);
DFFARX1 I_31311 (I535884,I3563,I535858,I535901,);
not I_31312 (I535850,I535901);
DFFARX1 I_31313 (I220857,I3563,I535858,I535932,);
not I_31314 (I535940,I220851);
nor I_31315 (I535957,I535884,I535940);
not I_31316 (I535974,I220845);
not I_31317 (I535991,I220842);
nand I_31318 (I536008,I535991,I220845);
nor I_31319 (I536025,I535940,I536008);
nor I_31320 (I536042,I535932,I536025);
DFFARX1 I_31321 (I535991,I3563,I535858,I535847,);
nor I_31322 (I536073,I220842,I220836);
nand I_31323 (I536090,I536073,I220854);
nor I_31324 (I536107,I536090,I535974);
nand I_31325 (I535832,I536107,I220851);
DFFARX1 I_31326 (I536090,I3563,I535858,I535844,);
nand I_31327 (I536152,I535974,I220842);
nor I_31328 (I536169,I535974,I220842);
nand I_31329 (I535838,I535957,I536169);
not I_31330 (I536200,I220848);
nor I_31331 (I536217,I536200,I536152);
DFFARX1 I_31332 (I536217,I3563,I535858,I535826,);
nor I_31333 (I536248,I536200,I220833);
and I_31334 (I536265,I536248,I220839);
or I_31335 (I536282,I536265,I220836);
DFFARX1 I_31336 (I536282,I3563,I535858,I536308,);
nor I_31337 (I536316,I536308,I535932);
nor I_31338 (I535835,I535884,I536316);
not I_31339 (I536347,I536308);
nor I_31340 (I536364,I536347,I536042);
DFFARX1 I_31341 (I536364,I3563,I535858,I535841,);
nand I_31342 (I536395,I536347,I535974);
nor I_31343 (I535829,I536200,I536395);
not I_31344 (I536453,I3570);
DFFARX1 I_31345 (I597148,I3563,I536453,I536479,);
DFFARX1 I_31346 (I536479,I3563,I536453,I536496,);
not I_31347 (I536445,I536496);
DFFARX1 I_31348 (I597160,I3563,I536453,I536527,);
not I_31349 (I536535,I597145);
nor I_31350 (I536552,I536479,I536535);
not I_31351 (I536569,I597163);
not I_31352 (I536586,I597154);
nand I_31353 (I536603,I536586,I597163);
nor I_31354 (I536620,I536535,I536603);
nor I_31355 (I536637,I536527,I536620);
DFFARX1 I_31356 (I536586,I3563,I536453,I536442,);
nor I_31357 (I536668,I597154,I597166);
nand I_31358 (I536685,I536668,I597169);
nor I_31359 (I536702,I536685,I536569);
nand I_31360 (I536427,I536702,I597145);
DFFARX1 I_31361 (I536685,I3563,I536453,I536439,);
nand I_31362 (I536747,I536569,I597154);
nor I_31363 (I536764,I536569,I597154);
nand I_31364 (I536433,I536552,I536764);
not I_31365 (I536795,I597145);
nor I_31366 (I536812,I536795,I536747);
DFFARX1 I_31367 (I536812,I3563,I536453,I536421,);
nor I_31368 (I536843,I536795,I597157);
and I_31369 (I536860,I536843,I597151);
or I_31370 (I536877,I536860,I597148);
DFFARX1 I_31371 (I536877,I3563,I536453,I536903,);
nor I_31372 (I536911,I536903,I536527);
nor I_31373 (I536430,I536479,I536911);
not I_31374 (I536942,I536903);
nor I_31375 (I536959,I536942,I536637);
DFFARX1 I_31376 (I536959,I3563,I536453,I536436,);
nand I_31377 (I536990,I536942,I536569);
nor I_31378 (I536424,I536795,I536990);
not I_31379 (I537048,I3570);
DFFARX1 I_31380 (I513794,I3563,I537048,I537074,);
DFFARX1 I_31381 (I537074,I3563,I537048,I537091,);
not I_31382 (I537040,I537091);
DFFARX1 I_31383 (I513818,I3563,I537048,I537122,);
not I_31384 (I537130,I513797);
nor I_31385 (I537147,I537074,I537130);
not I_31386 (I537164,I513803);
not I_31387 (I537181,I513809);
nand I_31388 (I537198,I537181,I513803);
nor I_31389 (I537215,I537130,I537198);
nor I_31390 (I537232,I537122,I537215);
DFFARX1 I_31391 (I537181,I3563,I537048,I537037,);
nor I_31392 (I537263,I513809,I513821);
nand I_31393 (I537280,I537263,I513815);
nor I_31394 (I537297,I537280,I537164);
nand I_31395 (I537022,I537297,I513797);
DFFARX1 I_31396 (I537280,I3563,I537048,I537034,);
nand I_31397 (I537342,I537164,I513809);
nor I_31398 (I537359,I537164,I513809);
nand I_31399 (I537028,I537147,I537359);
not I_31400 (I537390,I513800);
nor I_31401 (I537407,I537390,I537342);
DFFARX1 I_31402 (I537407,I3563,I537048,I537016,);
nor I_31403 (I537438,I537390,I513794);
and I_31404 (I537455,I537438,I513812);
or I_31405 (I537472,I537455,I513806);
DFFARX1 I_31406 (I537472,I3563,I537048,I537498,);
nor I_31407 (I537506,I537498,I537122);
nor I_31408 (I537025,I537074,I537506);
not I_31409 (I537537,I537498);
nor I_31410 (I537554,I537537,I537232);
DFFARX1 I_31411 (I537554,I3563,I537048,I537031,);
nand I_31412 (I537585,I537537,I537164);
nor I_31413 (I537019,I537390,I537585);
not I_31414 (I537643,I3570);
DFFARX1 I_31415 (I201793,I3563,I537643,I537669,);
DFFARX1 I_31416 (I537669,I3563,I537643,I537686,);
not I_31417 (I537635,I537686);
DFFARX1 I_31418 (I201817,I3563,I537643,I537717,);
not I_31419 (I537725,I201811);
nor I_31420 (I537742,I537669,I537725);
not I_31421 (I537759,I201805);
not I_31422 (I537776,I201802);
nand I_31423 (I537793,I537776,I201805);
nor I_31424 (I537810,I537725,I537793);
nor I_31425 (I537827,I537717,I537810);
DFFARX1 I_31426 (I537776,I3563,I537643,I537632,);
nor I_31427 (I537858,I201802,I201796);
nand I_31428 (I537875,I537858,I201814);
nor I_31429 (I537892,I537875,I537759);
nand I_31430 (I537617,I537892,I201811);
DFFARX1 I_31431 (I537875,I3563,I537643,I537629,);
nand I_31432 (I537937,I537759,I201802);
nor I_31433 (I537954,I537759,I201802);
nand I_31434 (I537623,I537742,I537954);
not I_31435 (I537985,I201808);
nor I_31436 (I538002,I537985,I537937);
DFFARX1 I_31437 (I538002,I3563,I537643,I537611,);
nor I_31438 (I538033,I537985,I201793);
and I_31439 (I538050,I538033,I201799);
or I_31440 (I538067,I538050,I201796);
DFFARX1 I_31441 (I538067,I3563,I537643,I538093,);
nor I_31442 (I538101,I538093,I537717);
nor I_31443 (I537620,I537669,I538101);
not I_31444 (I538132,I538093);
nor I_31445 (I538149,I538132,I537827);
DFFARX1 I_31446 (I538149,I3563,I537643,I537626,);
nand I_31447 (I538180,I538132,I537759);
nor I_31448 (I537614,I537985,I538180);
not I_31449 (I538238,I3570);
DFFARX1 I_31450 (I866400,I3563,I538238,I538264,);
DFFARX1 I_31451 (I538264,I3563,I538238,I538281,);
not I_31452 (I538230,I538281);
DFFARX1 I_31453 (I866397,I3563,I538238,I538312,);
not I_31454 (I538320,I866397);
nor I_31455 (I538337,I538264,I538320);
not I_31456 (I538354,I866394);
not I_31457 (I538371,I866409);
nand I_31458 (I538388,I538371,I866394);
nor I_31459 (I538405,I538320,I538388);
nor I_31460 (I538422,I538312,I538405);
DFFARX1 I_31461 (I538371,I3563,I538238,I538227,);
nor I_31462 (I538453,I866409,I866403);
nand I_31463 (I538470,I538453,I866391);
nor I_31464 (I538487,I538470,I538354);
nand I_31465 (I538212,I538487,I866397);
DFFARX1 I_31466 (I538470,I3563,I538238,I538224,);
nand I_31467 (I538532,I538354,I866409);
nor I_31468 (I538549,I538354,I866409);
nand I_31469 (I538218,I538337,I538549);
not I_31470 (I538580,I866412);
nor I_31471 (I538597,I538580,I538532);
DFFARX1 I_31472 (I538597,I3563,I538238,I538206,);
nor I_31473 (I538628,I538580,I866391);
and I_31474 (I538645,I538628,I866406);
or I_31475 (I538662,I538645,I866394);
DFFARX1 I_31476 (I538662,I3563,I538238,I538688,);
nor I_31477 (I538696,I538688,I538312);
nor I_31478 (I538215,I538264,I538696);
not I_31479 (I538727,I538688);
nor I_31480 (I538744,I538727,I538422);
DFFARX1 I_31481 (I538744,I3563,I538238,I538221,);
nand I_31482 (I538775,I538727,I538354);
nor I_31483 (I538209,I538580,I538775);
not I_31484 (I538833,I3570);
DFFARX1 I_31485 (I410279,I3563,I538833,I538859,);
DFFARX1 I_31486 (I538859,I3563,I538833,I538876,);
not I_31487 (I538825,I538876);
DFFARX1 I_31488 (I410267,I3563,I538833,I538907,);
not I_31489 (I538915,I410270);
nor I_31490 (I538932,I538859,I538915);
not I_31491 (I538949,I410273);
not I_31492 (I538966,I410285);
nand I_31493 (I538983,I538966,I410273);
nor I_31494 (I539000,I538915,I538983);
nor I_31495 (I539017,I538907,I539000);
DFFARX1 I_31496 (I538966,I3563,I538833,I538822,);
nor I_31497 (I539048,I410285,I410276);
nand I_31498 (I539065,I539048,I410264);
nor I_31499 (I539082,I539065,I538949);
nand I_31500 (I538807,I539082,I410270);
DFFARX1 I_31501 (I539065,I3563,I538833,I538819,);
nand I_31502 (I539127,I538949,I410285);
nor I_31503 (I539144,I538949,I410285);
nand I_31504 (I538813,I538932,I539144);
not I_31505 (I539175,I410282);
nor I_31506 (I539192,I539175,I539127);
DFFARX1 I_31507 (I539192,I3563,I538833,I538801,);
nor I_31508 (I539223,I539175,I410288);
and I_31509 (I539240,I539223,I410291);
or I_31510 (I539257,I539240,I410264);
DFFARX1 I_31511 (I539257,I3563,I538833,I539283,);
nor I_31512 (I539291,I539283,I538907);
nor I_31513 (I538810,I538859,I539291);
not I_31514 (I539322,I539283);
nor I_31515 (I539339,I539322,I539017);
DFFARX1 I_31516 (I539339,I3563,I538833,I538816,);
nand I_31517 (I539370,I539322,I538949);
nor I_31518 (I538804,I539175,I539370);
not I_31519 (I539428,I3570);
DFFARX1 I_31520 (I1126271,I3563,I539428,I539454,);
DFFARX1 I_31521 (I539454,I3563,I539428,I539471,);
not I_31522 (I539420,I539471);
DFFARX1 I_31523 (I1126253,I3563,I539428,I539502,);
not I_31524 (I539510,I1126259);
nor I_31525 (I539527,I539454,I539510);
not I_31526 (I539544,I1126274);
not I_31527 (I539561,I1126265);
nand I_31528 (I539578,I539561,I1126274);
nor I_31529 (I539595,I539510,I539578);
nor I_31530 (I539612,I539502,I539595);
DFFARX1 I_31531 (I539561,I3563,I539428,I539417,);
nor I_31532 (I539643,I1126265,I1126277);
nand I_31533 (I539660,I539643,I1126256);
nor I_31534 (I539677,I539660,I539544);
nand I_31535 (I539402,I539677,I1126259);
DFFARX1 I_31536 (I539660,I3563,I539428,I539414,);
nand I_31537 (I539722,I539544,I1126265);
nor I_31538 (I539739,I539544,I1126265);
nand I_31539 (I539408,I539527,I539739);
not I_31540 (I539770,I1126262);
nor I_31541 (I539787,I539770,I539722);
DFFARX1 I_31542 (I539787,I3563,I539428,I539396,);
nor I_31543 (I539818,I539770,I1126268);
and I_31544 (I539835,I539818,I1126253);
or I_31545 (I539852,I539835,I1126256);
DFFARX1 I_31546 (I539852,I3563,I539428,I539878,);
nor I_31547 (I539886,I539878,I539502);
nor I_31548 (I539405,I539454,I539886);
not I_31549 (I539917,I539878);
nor I_31550 (I539934,I539917,I539612);
DFFARX1 I_31551 (I539934,I3563,I539428,I539411,);
nand I_31552 (I539965,I539917,I539544);
nor I_31553 (I539399,I539770,I539965);
not I_31554 (I540023,I3570);
DFFARX1 I_31555 (I217263,I3563,I540023,I540049,);
DFFARX1 I_31556 (I540049,I3563,I540023,I540066,);
not I_31557 (I540015,I540066);
DFFARX1 I_31558 (I217287,I3563,I540023,I540097,);
not I_31559 (I540105,I217281);
nor I_31560 (I540122,I540049,I540105);
not I_31561 (I540139,I217275);
not I_31562 (I540156,I217272);
nand I_31563 (I540173,I540156,I217275);
nor I_31564 (I540190,I540105,I540173);
nor I_31565 (I540207,I540097,I540190);
DFFARX1 I_31566 (I540156,I3563,I540023,I540012,);
nor I_31567 (I540238,I217272,I217266);
nand I_31568 (I540255,I540238,I217284);
nor I_31569 (I540272,I540255,I540139);
nand I_31570 (I539997,I540272,I217281);
DFFARX1 I_31571 (I540255,I3563,I540023,I540009,);
nand I_31572 (I540317,I540139,I217272);
nor I_31573 (I540334,I540139,I217272);
nand I_31574 (I540003,I540122,I540334);
not I_31575 (I540365,I217278);
nor I_31576 (I540382,I540365,I540317);
DFFARX1 I_31577 (I540382,I3563,I540023,I539991,);
nor I_31578 (I540413,I540365,I217263);
and I_31579 (I540430,I540413,I217269);
or I_31580 (I540447,I540430,I217266);
DFFARX1 I_31581 (I540447,I3563,I540023,I540473,);
nor I_31582 (I540481,I540473,I540097);
nor I_31583 (I540000,I540049,I540481);
not I_31584 (I540512,I540473);
nor I_31585 (I540529,I540512,I540207);
DFFARX1 I_31586 (I540529,I3563,I540023,I540006,);
nand I_31587 (I540560,I540512,I540139);
nor I_31588 (I539994,I540365,I540560);
not I_31589 (I540618,I3570);
DFFARX1 I_31590 (I779802,I3563,I540618,I540644,);
DFFARX1 I_31591 (I540644,I3563,I540618,I540661,);
not I_31592 (I540610,I540661);
DFFARX1 I_31593 (I779796,I3563,I540618,I540692,);
not I_31594 (I540700,I779793);
nor I_31595 (I540717,I540644,I540700);
not I_31596 (I540734,I779805);
not I_31597 (I540751,I779808);
nand I_31598 (I540768,I540751,I779805);
nor I_31599 (I540785,I540700,I540768);
nor I_31600 (I540802,I540692,I540785);
DFFARX1 I_31601 (I540751,I3563,I540618,I540607,);
nor I_31602 (I540833,I779808,I779817);
nand I_31603 (I540850,I540833,I779811);
nor I_31604 (I540867,I540850,I540734);
nand I_31605 (I540592,I540867,I779793);
DFFARX1 I_31606 (I540850,I3563,I540618,I540604,);
nand I_31607 (I540912,I540734,I779808);
nor I_31608 (I540929,I540734,I779808);
nand I_31609 (I540598,I540717,I540929);
not I_31610 (I540960,I779799);
nor I_31611 (I540977,I540960,I540912);
DFFARX1 I_31612 (I540977,I3563,I540618,I540586,);
nor I_31613 (I541008,I540960,I779814);
and I_31614 (I541025,I541008,I779793);
or I_31615 (I541042,I541025,I779796);
DFFARX1 I_31616 (I541042,I3563,I540618,I541068,);
nor I_31617 (I541076,I541068,I540692);
nor I_31618 (I540595,I540644,I541076);
not I_31619 (I541107,I541068);
nor I_31620 (I541124,I541107,I540802);
DFFARX1 I_31621 (I541124,I3563,I540618,I540601,);
nand I_31622 (I541155,I541107,I540734);
nor I_31623 (I540589,I540960,I541155);
not I_31624 (I541213,I3570);
DFFARX1 I_31625 (I1319552,I3563,I541213,I541239,);
DFFARX1 I_31626 (I541239,I3563,I541213,I541256,);
not I_31627 (I541205,I541256);
DFFARX1 I_31628 (I1319558,I3563,I541213,I541287,);
not I_31629 (I541295,I1319546);
nor I_31630 (I541312,I541239,I541295);
not I_31631 (I541329,I1319549);
not I_31632 (I541346,I1319555);
nand I_31633 (I541363,I541346,I1319549);
nor I_31634 (I541380,I541295,I541363);
nor I_31635 (I541397,I541287,I541380);
DFFARX1 I_31636 (I541346,I3563,I541213,I541202,);
nor I_31637 (I541428,I1319555,I1319546);
nand I_31638 (I541445,I541428,I1319564);
nor I_31639 (I541462,I541445,I541329);
nand I_31640 (I541187,I541462,I1319546);
DFFARX1 I_31641 (I541445,I3563,I541213,I541199,);
nand I_31642 (I541507,I541329,I1319555);
nor I_31643 (I541524,I541329,I1319555);
nand I_31644 (I541193,I541312,I541524);
not I_31645 (I541555,I1319543);
nor I_31646 (I541572,I541555,I541507);
DFFARX1 I_31647 (I541572,I3563,I541213,I541181,);
nor I_31648 (I541603,I541555,I1319567);
and I_31649 (I541620,I541603,I1319543);
or I_31650 (I541637,I541620,I1319561);
DFFARX1 I_31651 (I541637,I3563,I541213,I541663,);
nor I_31652 (I541671,I541663,I541287);
nor I_31653 (I541190,I541239,I541671);
not I_31654 (I541702,I541663);
nor I_31655 (I541719,I541702,I541397);
DFFARX1 I_31656 (I541719,I3563,I541213,I541196,);
nand I_31657 (I541750,I541702,I541329);
nor I_31658 (I541184,I541555,I541750);
not I_31659 (I541808,I3570);
DFFARX1 I_31660 (I218453,I3563,I541808,I541834,);
DFFARX1 I_31661 (I541834,I3563,I541808,I541851,);
not I_31662 (I541800,I541851);
DFFARX1 I_31663 (I218477,I3563,I541808,I541882,);
not I_31664 (I541890,I218471);
nor I_31665 (I541907,I541834,I541890);
not I_31666 (I541924,I218465);
not I_31667 (I541941,I218462);
nand I_31668 (I541958,I541941,I218465);
nor I_31669 (I541975,I541890,I541958);
nor I_31670 (I541992,I541882,I541975);
DFFARX1 I_31671 (I541941,I3563,I541808,I541797,);
nor I_31672 (I542023,I218462,I218456);
nand I_31673 (I542040,I542023,I218474);
nor I_31674 (I542057,I542040,I541924);
nand I_31675 (I541782,I542057,I218471);
DFFARX1 I_31676 (I542040,I3563,I541808,I541794,);
nand I_31677 (I542102,I541924,I218462);
nor I_31678 (I542119,I541924,I218462);
nand I_31679 (I541788,I541907,I542119);
not I_31680 (I542150,I218468);
nor I_31681 (I542167,I542150,I542102);
DFFARX1 I_31682 (I542167,I3563,I541808,I541776,);
nor I_31683 (I542198,I542150,I218453);
and I_31684 (I542215,I542198,I218459);
or I_31685 (I542232,I542215,I218456);
DFFARX1 I_31686 (I542232,I3563,I541808,I542258,);
nor I_31687 (I542266,I542258,I541882);
nor I_31688 (I541785,I541834,I542266);
not I_31689 (I542297,I542258);
nor I_31690 (I542314,I542297,I541992);
DFFARX1 I_31691 (I542314,I3563,I541808,I541791,);
nand I_31692 (I542345,I542297,I541924);
nor I_31693 (I541779,I542150,I542345);
not I_31694 (I542403,I3570);
DFFARX1 I_31695 (I691946,I3563,I542403,I542429,);
DFFARX1 I_31696 (I542429,I3563,I542403,I542446,);
not I_31697 (I542395,I542446);
DFFARX1 I_31698 (I691940,I3563,I542403,I542477,);
not I_31699 (I542485,I691937);
nor I_31700 (I542502,I542429,I542485);
not I_31701 (I542519,I691949);
not I_31702 (I542536,I691952);
nand I_31703 (I542553,I542536,I691949);
nor I_31704 (I542570,I542485,I542553);
nor I_31705 (I542587,I542477,I542570);
DFFARX1 I_31706 (I542536,I3563,I542403,I542392,);
nor I_31707 (I542618,I691952,I691961);
nand I_31708 (I542635,I542618,I691955);
nor I_31709 (I542652,I542635,I542519);
nand I_31710 (I542377,I542652,I691937);
DFFARX1 I_31711 (I542635,I3563,I542403,I542389,);
nand I_31712 (I542697,I542519,I691952);
nor I_31713 (I542714,I542519,I691952);
nand I_31714 (I542383,I542502,I542714);
not I_31715 (I542745,I691943);
nor I_31716 (I542762,I542745,I542697);
DFFARX1 I_31717 (I542762,I3563,I542403,I542371,);
nor I_31718 (I542793,I542745,I691958);
and I_31719 (I542810,I542793,I691937);
or I_31720 (I542827,I542810,I691940);
DFFARX1 I_31721 (I542827,I3563,I542403,I542853,);
nor I_31722 (I542861,I542853,I542477);
nor I_31723 (I542380,I542429,I542861);
not I_31724 (I542892,I542853);
nor I_31725 (I542909,I542892,I542587);
DFFARX1 I_31726 (I542909,I3563,I542403,I542386,);
nand I_31727 (I542940,I542892,I542519);
nor I_31728 (I542374,I542745,I542940);
not I_31729 (I542998,I3570);
DFFARX1 I_31730 (I167878,I3563,I542998,I543024,);
DFFARX1 I_31731 (I543024,I3563,I542998,I543041,);
not I_31732 (I542990,I543041);
DFFARX1 I_31733 (I167902,I3563,I542998,I543072,);
not I_31734 (I543080,I167896);
nor I_31735 (I543097,I543024,I543080);
not I_31736 (I543114,I167890);
not I_31737 (I543131,I167887);
nand I_31738 (I543148,I543131,I167890);
nor I_31739 (I543165,I543080,I543148);
nor I_31740 (I543182,I543072,I543165);
DFFARX1 I_31741 (I543131,I3563,I542998,I542987,);
nor I_31742 (I543213,I167887,I167881);
nand I_31743 (I543230,I543213,I167899);
nor I_31744 (I543247,I543230,I543114);
nand I_31745 (I542972,I543247,I167896);
DFFARX1 I_31746 (I543230,I3563,I542998,I542984,);
nand I_31747 (I543292,I543114,I167887);
nor I_31748 (I543309,I543114,I167887);
nand I_31749 (I542978,I543097,I543309);
not I_31750 (I543340,I167893);
nor I_31751 (I543357,I543340,I543292);
DFFARX1 I_31752 (I543357,I3563,I542998,I542966,);
nor I_31753 (I543388,I543340,I167878);
and I_31754 (I543405,I543388,I167884);
or I_31755 (I543422,I543405,I167881);
DFFARX1 I_31756 (I543422,I3563,I542998,I543448,);
nor I_31757 (I543456,I543448,I543072);
nor I_31758 (I542975,I543024,I543456);
not I_31759 (I543487,I543448);
nor I_31760 (I543504,I543487,I543182);
DFFARX1 I_31761 (I543504,I3563,I542998,I542981,);
nand I_31762 (I543535,I543487,I543114);
nor I_31763 (I542969,I543340,I543535);
not I_31764 (I543593,I3570);
DFFARX1 I_31765 (I655526,I3563,I543593,I543619,);
DFFARX1 I_31766 (I543619,I3563,I543593,I543636,);
not I_31767 (I543585,I543636);
DFFARX1 I_31768 (I655538,I3563,I543593,I543667,);
not I_31769 (I543675,I655523);
nor I_31770 (I543692,I543619,I543675);
not I_31771 (I543709,I655541);
not I_31772 (I543726,I655532);
nand I_31773 (I543743,I543726,I655541);
nor I_31774 (I543760,I543675,I543743);
nor I_31775 (I543777,I543667,I543760);
DFFARX1 I_31776 (I543726,I3563,I543593,I543582,);
nor I_31777 (I543808,I655532,I655544);
nand I_31778 (I543825,I543808,I655547);
nor I_31779 (I543842,I543825,I543709);
nand I_31780 (I543567,I543842,I655523);
DFFARX1 I_31781 (I543825,I3563,I543593,I543579,);
nand I_31782 (I543887,I543709,I655532);
nor I_31783 (I543904,I543709,I655532);
nand I_31784 (I543573,I543692,I543904);
not I_31785 (I543935,I655523);
nor I_31786 (I543952,I543935,I543887);
DFFARX1 I_31787 (I543952,I3563,I543593,I543561,);
nor I_31788 (I543983,I543935,I655535);
and I_31789 (I544000,I543983,I655529);
or I_31790 (I544017,I544000,I655526);
DFFARX1 I_31791 (I544017,I3563,I543593,I544043,);
nor I_31792 (I544051,I544043,I543667);
nor I_31793 (I543570,I543619,I544051);
not I_31794 (I544082,I544043);
nor I_31795 (I544099,I544082,I543777);
DFFARX1 I_31796 (I544099,I3563,I543593,I543576,);
nand I_31797 (I544130,I544082,I543709);
nor I_31798 (I543564,I543935,I544130);
not I_31799 (I544188,I3570);
DFFARX1 I_31800 (I1355923,I3563,I544188,I544214,);
DFFARX1 I_31801 (I544214,I3563,I544188,I544231,);
not I_31802 (I544180,I544231);
DFFARX1 I_31803 (I1355929,I3563,I544188,I544262,);
not I_31804 (I544270,I1355944);
nor I_31805 (I544287,I544214,I544270);
not I_31806 (I544304,I1355935);
not I_31807 (I544321,I1355932);
nand I_31808 (I544338,I544321,I1355935);
nor I_31809 (I544355,I544270,I544338);
nor I_31810 (I544372,I544262,I544355);
DFFARX1 I_31811 (I544321,I3563,I544188,I544177,);
nor I_31812 (I544403,I1355932,I1355923);
nand I_31813 (I544420,I544403,I1355947);
nor I_31814 (I544437,I544420,I544304);
nand I_31815 (I544162,I544437,I1355944);
DFFARX1 I_31816 (I544420,I3563,I544188,I544174,);
nand I_31817 (I544482,I544304,I1355932);
nor I_31818 (I544499,I544304,I1355932);
nand I_31819 (I544168,I544287,I544499);
not I_31820 (I544530,I1355941);
nor I_31821 (I544547,I544530,I544482);
DFFARX1 I_31822 (I544547,I3563,I544188,I544156,);
nor I_31823 (I544578,I544530,I1355926);
and I_31824 (I544595,I544578,I1355938);
or I_31825 (I544612,I544595,I1355950);
DFFARX1 I_31826 (I544612,I3563,I544188,I544638,);
nor I_31827 (I544646,I544638,I544262);
nor I_31828 (I544165,I544214,I544646);
not I_31829 (I544677,I544638);
nor I_31830 (I544694,I544677,I544372);
DFFARX1 I_31831 (I544694,I3563,I544188,I544171,);
nand I_31832 (I544725,I544677,I544304);
nor I_31833 (I544159,I544530,I544725);
not I_31834 (I544783,I3570);
DFFARX1 I_31835 (I1119913,I3563,I544783,I544809,);
DFFARX1 I_31836 (I544809,I3563,I544783,I544826,);
not I_31837 (I544775,I544826);
DFFARX1 I_31838 (I1119895,I3563,I544783,I544857,);
not I_31839 (I544865,I1119901);
nor I_31840 (I544882,I544809,I544865);
not I_31841 (I544899,I1119916);
not I_31842 (I544916,I1119907);
nand I_31843 (I544933,I544916,I1119916);
nor I_31844 (I544950,I544865,I544933);
nor I_31845 (I544967,I544857,I544950);
DFFARX1 I_31846 (I544916,I3563,I544783,I544772,);
nor I_31847 (I544998,I1119907,I1119919);
nand I_31848 (I545015,I544998,I1119898);
nor I_31849 (I545032,I545015,I544899);
nand I_31850 (I544757,I545032,I1119901);
DFFARX1 I_31851 (I545015,I3563,I544783,I544769,);
nand I_31852 (I545077,I544899,I1119907);
nor I_31853 (I545094,I544899,I1119907);
nand I_31854 (I544763,I544882,I545094);
not I_31855 (I545125,I1119904);
nor I_31856 (I545142,I545125,I545077);
DFFARX1 I_31857 (I545142,I3563,I544783,I544751,);
nor I_31858 (I545173,I545125,I1119910);
and I_31859 (I545190,I545173,I1119895);
or I_31860 (I545207,I545190,I1119898);
DFFARX1 I_31861 (I545207,I3563,I544783,I545233,);
nor I_31862 (I545241,I545233,I544857);
nor I_31863 (I544760,I544809,I545241);
not I_31864 (I545272,I545233);
nor I_31865 (I545289,I545272,I544967);
DFFARX1 I_31866 (I545289,I3563,I544783,I544766,);
nand I_31867 (I545320,I545272,I544899);
nor I_31868 (I544754,I545125,I545320);
not I_31869 (I545378,I3570);
DFFARX1 I_31870 (I645122,I3563,I545378,I545404,);
DFFARX1 I_31871 (I545404,I3563,I545378,I545421,);
not I_31872 (I545370,I545421);
DFFARX1 I_31873 (I645134,I3563,I545378,I545452,);
not I_31874 (I545460,I645119);
nor I_31875 (I545477,I545404,I545460);
not I_31876 (I545494,I645137);
not I_31877 (I545511,I645128);
nand I_31878 (I545528,I545511,I645137);
nor I_31879 (I545545,I545460,I545528);
nor I_31880 (I545562,I545452,I545545);
DFFARX1 I_31881 (I545511,I3563,I545378,I545367,);
nor I_31882 (I545593,I645128,I645140);
nand I_31883 (I545610,I545593,I645143);
nor I_31884 (I545627,I545610,I545494);
nand I_31885 (I545352,I545627,I645119);
DFFARX1 I_31886 (I545610,I3563,I545378,I545364,);
nand I_31887 (I545672,I545494,I645128);
nor I_31888 (I545689,I545494,I645128);
nand I_31889 (I545358,I545477,I545689);
not I_31890 (I545720,I645119);
nor I_31891 (I545737,I545720,I545672);
DFFARX1 I_31892 (I545737,I3563,I545378,I545346,);
nor I_31893 (I545768,I545720,I645131);
and I_31894 (I545785,I545768,I645125);
or I_31895 (I545802,I545785,I645122);
DFFARX1 I_31896 (I545802,I3563,I545378,I545828,);
nor I_31897 (I545836,I545828,I545452);
nor I_31898 (I545355,I545404,I545836);
not I_31899 (I545867,I545828);
nor I_31900 (I545884,I545867,I545562);
DFFARX1 I_31901 (I545884,I3563,I545378,I545361,);
nand I_31902 (I545915,I545867,I545494);
nor I_31903 (I545349,I545720,I545915);
not I_31904 (I545973,I3570);
DFFARX1 I_31905 (I2916,I3563,I545973,I545999,);
DFFARX1 I_31906 (I545999,I3563,I545973,I546016,);
not I_31907 (I545965,I546016);
DFFARX1 I_31908 (I3044,I3563,I545973,I546047,);
not I_31909 (I546055,I1684);
nor I_31910 (I546072,I545999,I546055);
not I_31911 (I546089,I3324);
not I_31912 (I546106,I3204);
nand I_31913 (I546123,I546106,I3324);
nor I_31914 (I546140,I546055,I546123);
nor I_31915 (I546157,I546047,I546140);
DFFARX1 I_31916 (I546106,I3563,I545973,I545962,);
nor I_31917 (I546188,I3204,I2180);
nand I_31918 (I546205,I546188,I3292);
nor I_31919 (I546222,I546205,I546089);
nand I_31920 (I545947,I546222,I1684);
DFFARX1 I_31921 (I546205,I3563,I545973,I545959,);
nand I_31922 (I546267,I546089,I3204);
nor I_31923 (I546284,I546089,I3204);
nand I_31924 (I545953,I546072,I546284);
not I_31925 (I546315,I2596);
nor I_31926 (I546332,I546315,I546267);
DFFARX1 I_31927 (I546332,I3563,I545973,I545941,);
nor I_31928 (I546363,I546315,I1820);
and I_31929 (I546380,I546363,I3364);
or I_31930 (I546397,I546380,I2636);
DFFARX1 I_31931 (I546397,I3563,I545973,I546423,);
nor I_31932 (I546431,I546423,I546047);
nor I_31933 (I545950,I545999,I546431);
not I_31934 (I546462,I546423);
nor I_31935 (I546479,I546462,I546157);
DFFARX1 I_31936 (I546479,I3563,I545973,I545956,);
nand I_31937 (I546510,I546462,I546089);
nor I_31938 (I545944,I546315,I546510);
not I_31939 (I546568,I3570);
DFFARX1 I_31940 (I1000808,I3563,I546568,I546594,);
DFFARX1 I_31941 (I546594,I3563,I546568,I546611,);
not I_31942 (I546560,I546611);
DFFARX1 I_31943 (I1000796,I3563,I546568,I546642,);
not I_31944 (I546650,I1000793);
nor I_31945 (I546667,I546594,I546650);
not I_31946 (I546684,I1000805);
not I_31947 (I546701,I1000802);
nand I_31948 (I546718,I546701,I1000805);
nor I_31949 (I546735,I546650,I546718);
nor I_31950 (I546752,I546642,I546735);
DFFARX1 I_31951 (I546701,I3563,I546568,I546557,);
nor I_31952 (I546783,I1000802,I1000811);
nand I_31953 (I546800,I546783,I1000814);
nor I_31954 (I546817,I546800,I546684);
nand I_31955 (I546542,I546817,I1000793);
DFFARX1 I_31956 (I546800,I3563,I546568,I546554,);
nand I_31957 (I546862,I546684,I1000802);
nor I_31958 (I546879,I546684,I1000802);
nand I_31959 (I546548,I546667,I546879);
not I_31960 (I546910,I1000817);
nor I_31961 (I546927,I546910,I546862);
DFFARX1 I_31962 (I546927,I3563,I546568,I546536,);
nor I_31963 (I546958,I546910,I1000820);
and I_31964 (I546975,I546958,I1000799);
or I_31965 (I546992,I546975,I1000793);
DFFARX1 I_31966 (I546992,I3563,I546568,I547018,);
nor I_31967 (I547026,I547018,I546642);
nor I_31968 (I546545,I546594,I547026);
not I_31969 (I547057,I547018);
nor I_31970 (I547074,I547057,I546752);
DFFARX1 I_31971 (I547074,I3563,I546568,I546551,);
nand I_31972 (I547105,I547057,I546684);
nor I_31973 (I546539,I546910,I547105);
not I_31974 (I547163,I3570);
DFFARX1 I_31975 (I2164,I3563,I547163,I547189,);
DFFARX1 I_31976 (I547189,I3563,I547163,I547206,);
not I_31977 (I547155,I547206);
DFFARX1 I_31978 (I2460,I3563,I547163,I547237,);
not I_31979 (I547245,I2340);
nor I_31980 (I547262,I547189,I547245);
not I_31981 (I547279,I3068);
not I_31982 (I547296,I2948);
nand I_31983 (I547313,I547296,I3068);
nor I_31984 (I547330,I547245,I547313);
nor I_31985 (I547347,I547237,I547330);
DFFARX1 I_31986 (I547296,I3563,I547163,I547152,);
nor I_31987 (I547378,I2948,I1724);
nand I_31988 (I547395,I547378,I3028);
nor I_31989 (I547412,I547395,I547279);
nand I_31990 (I547137,I547412,I2340);
DFFARX1 I_31991 (I547395,I3563,I547163,I547149,);
nand I_31992 (I547457,I547279,I2948);
nor I_31993 (I547474,I547279,I2948);
nand I_31994 (I547143,I547262,I547474);
not I_31995 (I547505,I2612);
nor I_31996 (I547522,I547505,I547457);
DFFARX1 I_31997 (I547522,I3563,I547163,I547131,);
nor I_31998 (I547553,I547505,I3036);
and I_31999 (I547570,I547553,I2436);
or I_32000 (I547587,I547570,I1364);
DFFARX1 I_32001 (I547587,I3563,I547163,I547613,);
nor I_32002 (I547621,I547613,I547237);
nor I_32003 (I547140,I547189,I547621);
not I_32004 (I547652,I547613);
nor I_32005 (I547669,I547652,I547347);
DFFARX1 I_32006 (I547669,I3563,I547163,I547146,);
nand I_32007 (I547700,I547652,I547279);
nor I_32008 (I547134,I547505,I547700);
not I_32009 (I547758,I3570);
DFFARX1 I_32010 (I67196,I3563,I547758,I547784,);
DFFARX1 I_32011 (I547784,I3563,I547758,I547801,);
not I_32012 (I547750,I547801);
DFFARX1 I_32013 (I67208,I3563,I547758,I547832,);
not I_32014 (I547840,I67199);
nor I_32015 (I547857,I547784,I547840);
not I_32016 (I547874,I67190);
not I_32017 (I547891,I67187);
nand I_32018 (I547908,I547891,I67190);
nor I_32019 (I547925,I547840,I547908);
nor I_32020 (I547942,I547832,I547925);
DFFARX1 I_32021 (I547891,I3563,I547758,I547747,);
nor I_32022 (I547973,I67187,I67187);
nand I_32023 (I547990,I547973,I67205);
nor I_32024 (I548007,I547990,I547874);
nand I_32025 (I547732,I548007,I67199);
DFFARX1 I_32026 (I547990,I3563,I547758,I547744,);
nand I_32027 (I548052,I547874,I67187);
nor I_32028 (I548069,I547874,I67187);
nand I_32029 (I547738,I547857,I548069);
not I_32030 (I548100,I67211);
nor I_32031 (I548117,I548100,I548052);
DFFARX1 I_32032 (I548117,I3563,I547758,I547726,);
nor I_32033 (I548148,I548100,I67190);
and I_32034 (I548165,I548148,I67193);
or I_32035 (I548182,I548165,I67202);
DFFARX1 I_32036 (I548182,I3563,I547758,I548208,);
nor I_32037 (I548216,I548208,I547832);
nor I_32038 (I547735,I547784,I548216);
not I_32039 (I548247,I548208);
nor I_32040 (I548264,I548247,I547942);
DFFARX1 I_32041 (I548264,I3563,I547758,I547741,);
nand I_32042 (I548295,I548247,I547874);
nor I_32043 (I547729,I548100,I548295);
not I_32044 (I548353,I3570);
DFFARX1 I_32045 (I110937,I3563,I548353,I548379,);
DFFARX1 I_32046 (I548379,I3563,I548353,I548396,);
not I_32047 (I548345,I548396);
DFFARX1 I_32048 (I110949,I3563,I548353,I548427,);
not I_32049 (I548435,I110940);
nor I_32050 (I548452,I548379,I548435);
not I_32051 (I548469,I110931);
not I_32052 (I548486,I110928);
nand I_32053 (I548503,I548486,I110931);
nor I_32054 (I548520,I548435,I548503);
nor I_32055 (I548537,I548427,I548520);
DFFARX1 I_32056 (I548486,I3563,I548353,I548342,);
nor I_32057 (I548568,I110928,I110928);
nand I_32058 (I548585,I548568,I110946);
nor I_32059 (I548602,I548585,I548469);
nand I_32060 (I548327,I548602,I110940);
DFFARX1 I_32061 (I548585,I3563,I548353,I548339,);
nand I_32062 (I548647,I548469,I110928);
nor I_32063 (I548664,I548469,I110928);
nand I_32064 (I548333,I548452,I548664);
not I_32065 (I548695,I110952);
nor I_32066 (I548712,I548695,I548647);
DFFARX1 I_32067 (I548712,I3563,I548353,I548321,);
nor I_32068 (I548743,I548695,I110931);
and I_32069 (I548760,I548743,I110934);
or I_32070 (I548777,I548760,I110943);
DFFARX1 I_32071 (I548777,I3563,I548353,I548803,);
nor I_32072 (I548811,I548803,I548427);
nor I_32073 (I548330,I548379,I548811);
not I_32074 (I548842,I548803);
nor I_32075 (I548859,I548842,I548537);
DFFARX1 I_32076 (I548859,I3563,I548353,I548336,);
nand I_32077 (I548890,I548842,I548469);
nor I_32078 (I548324,I548695,I548890);
not I_32079 (I548948,I3570);
DFFARX1 I_32080 (I940084,I3563,I548948,I548974,);
DFFARX1 I_32081 (I548974,I3563,I548948,I548991,);
not I_32082 (I548940,I548991);
DFFARX1 I_32083 (I940072,I3563,I548948,I549022,);
not I_32084 (I549030,I940069);
nor I_32085 (I549047,I548974,I549030);
not I_32086 (I549064,I940081);
not I_32087 (I549081,I940078);
nand I_32088 (I549098,I549081,I940081);
nor I_32089 (I549115,I549030,I549098);
nor I_32090 (I549132,I549022,I549115);
DFFARX1 I_32091 (I549081,I3563,I548948,I548937,);
nor I_32092 (I549163,I940078,I940087);
nand I_32093 (I549180,I549163,I940090);
nor I_32094 (I549197,I549180,I549064);
nand I_32095 (I548922,I549197,I940069);
DFFARX1 I_32096 (I549180,I3563,I548948,I548934,);
nand I_32097 (I549242,I549064,I940078);
nor I_32098 (I549259,I549064,I940078);
nand I_32099 (I548928,I549047,I549259);
not I_32100 (I549290,I940093);
nor I_32101 (I549307,I549290,I549242);
DFFARX1 I_32102 (I549307,I3563,I548948,I548916,);
nor I_32103 (I549338,I549290,I940096);
and I_32104 (I549355,I549338,I940075);
or I_32105 (I549372,I549355,I940069);
DFFARX1 I_32106 (I549372,I3563,I548948,I549398,);
nor I_32107 (I549406,I549398,I549022);
nor I_32108 (I548925,I548974,I549406);
not I_32109 (I549437,I549398);
nor I_32110 (I549454,I549437,I549132);
DFFARX1 I_32111 (I549454,I3563,I548948,I548931,);
nand I_32112 (I549485,I549437,I549064);
nor I_32113 (I548919,I549290,I549485);
not I_32114 (I549543,I3570);
DFFARX1 I_32115 (I944606,I3563,I549543,I549569,);
DFFARX1 I_32116 (I549569,I3563,I549543,I549586,);
not I_32117 (I549535,I549586);
DFFARX1 I_32118 (I944594,I3563,I549543,I549617,);
not I_32119 (I549625,I944591);
nor I_32120 (I549642,I549569,I549625);
not I_32121 (I549659,I944603);
not I_32122 (I549676,I944600);
nand I_32123 (I549693,I549676,I944603);
nor I_32124 (I549710,I549625,I549693);
nor I_32125 (I549727,I549617,I549710);
DFFARX1 I_32126 (I549676,I3563,I549543,I549532,);
nor I_32127 (I549758,I944600,I944609);
nand I_32128 (I549775,I549758,I944612);
nor I_32129 (I549792,I549775,I549659);
nand I_32130 (I549517,I549792,I944591);
DFFARX1 I_32131 (I549775,I3563,I549543,I549529,);
nand I_32132 (I549837,I549659,I944600);
nor I_32133 (I549854,I549659,I944600);
nand I_32134 (I549523,I549642,I549854);
not I_32135 (I549885,I944615);
nor I_32136 (I549902,I549885,I549837);
DFFARX1 I_32137 (I549902,I3563,I549543,I549511,);
nor I_32138 (I549933,I549885,I944618);
and I_32139 (I549950,I549933,I944597);
or I_32140 (I549967,I549950,I944591);
DFFARX1 I_32141 (I549967,I3563,I549543,I549993,);
nor I_32142 (I550001,I549993,I549617);
nor I_32143 (I549520,I549569,I550001);
not I_32144 (I550032,I549993);
nor I_32145 (I550049,I550032,I549727);
DFFARX1 I_32146 (I550049,I3563,I549543,I549526,);
nand I_32147 (I550080,I550032,I549659);
nor I_32148 (I549514,I549885,I550080);
not I_32149 (I550138,I3570);
DFFARX1 I_32150 (I894858,I3563,I550138,I550164,);
DFFARX1 I_32151 (I550164,I3563,I550138,I550181,);
not I_32152 (I550130,I550181);
DFFARX1 I_32153 (I894855,I3563,I550138,I550212,);
not I_32154 (I550220,I894855);
nor I_32155 (I550237,I550164,I550220);
not I_32156 (I550254,I894852);
not I_32157 (I550271,I894867);
nand I_32158 (I550288,I550271,I894852);
nor I_32159 (I550305,I550220,I550288);
nor I_32160 (I550322,I550212,I550305);
DFFARX1 I_32161 (I550271,I3563,I550138,I550127,);
nor I_32162 (I550353,I894867,I894861);
nand I_32163 (I550370,I550353,I894849);
nor I_32164 (I550387,I550370,I550254);
nand I_32165 (I550112,I550387,I894855);
DFFARX1 I_32166 (I550370,I3563,I550138,I550124,);
nand I_32167 (I550432,I550254,I894867);
nor I_32168 (I550449,I550254,I894867);
nand I_32169 (I550118,I550237,I550449);
not I_32170 (I550480,I894870);
nor I_32171 (I550497,I550480,I550432);
DFFARX1 I_32172 (I550497,I3563,I550138,I550106,);
nor I_32173 (I550528,I550480,I894849);
and I_32174 (I550545,I550528,I894864);
or I_32175 (I550562,I550545,I894852);
DFFARX1 I_32176 (I550562,I3563,I550138,I550588,);
nor I_32177 (I550596,I550588,I550212);
nor I_32178 (I550115,I550164,I550596);
not I_32179 (I550627,I550588);
nor I_32180 (I550644,I550627,I550322);
DFFARX1 I_32181 (I550644,I3563,I550138,I550121,);
nand I_32182 (I550675,I550627,I550254);
nor I_32183 (I550109,I550480,I550675);
not I_32184 (I550733,I3570);
DFFARX1 I_32185 (I690790,I3563,I550733,I550759,);
DFFARX1 I_32186 (I550759,I3563,I550733,I550776,);
not I_32187 (I550725,I550776);
DFFARX1 I_32188 (I690784,I3563,I550733,I550807,);
not I_32189 (I550815,I690781);
nor I_32190 (I550832,I550759,I550815);
not I_32191 (I550849,I690793);
not I_32192 (I550866,I690796);
nand I_32193 (I550883,I550866,I690793);
nor I_32194 (I550900,I550815,I550883);
nor I_32195 (I550917,I550807,I550900);
DFFARX1 I_32196 (I550866,I3563,I550733,I550722,);
nor I_32197 (I550948,I690796,I690805);
nand I_32198 (I550965,I550948,I690799);
nor I_32199 (I550982,I550965,I550849);
nand I_32200 (I550707,I550982,I690781);
DFFARX1 I_32201 (I550965,I3563,I550733,I550719,);
nand I_32202 (I551027,I550849,I690796);
nor I_32203 (I551044,I550849,I690796);
nand I_32204 (I550713,I550832,I551044);
not I_32205 (I551075,I690787);
nor I_32206 (I551092,I551075,I551027);
DFFARX1 I_32207 (I551092,I3563,I550733,I550701,);
nor I_32208 (I551123,I551075,I690802);
and I_32209 (I551140,I551123,I690781);
or I_32210 (I551157,I551140,I690784);
DFFARX1 I_32211 (I551157,I3563,I550733,I551183,);
nor I_32212 (I551191,I551183,I550807);
nor I_32213 (I550710,I550759,I551191);
not I_32214 (I551222,I551183);
nor I_32215 (I551239,I551222,I550917);
DFFARX1 I_32216 (I551239,I3563,I550733,I550716,);
nand I_32217 (I551270,I551222,I550849);
nor I_32218 (I550704,I551075,I551270);
not I_32219 (I551328,I3570);
DFFARX1 I_32220 (I659000,I3563,I551328,I551354,);
DFFARX1 I_32221 (I551354,I3563,I551328,I551371,);
not I_32222 (I551320,I551371);
DFFARX1 I_32223 (I658994,I3563,I551328,I551402,);
not I_32224 (I551410,I658991);
nor I_32225 (I551427,I551354,I551410);
not I_32226 (I551444,I659003);
not I_32227 (I551461,I659006);
nand I_32228 (I551478,I551461,I659003);
nor I_32229 (I551495,I551410,I551478);
nor I_32230 (I551512,I551402,I551495);
DFFARX1 I_32231 (I551461,I3563,I551328,I551317,);
nor I_32232 (I551543,I659006,I659015);
nand I_32233 (I551560,I551543,I659009);
nor I_32234 (I551577,I551560,I551444);
nand I_32235 (I551302,I551577,I658991);
DFFARX1 I_32236 (I551560,I3563,I551328,I551314,);
nand I_32237 (I551622,I551444,I659006);
nor I_32238 (I551639,I551444,I659006);
nand I_32239 (I551308,I551427,I551639);
not I_32240 (I551670,I658997);
nor I_32241 (I551687,I551670,I551622);
DFFARX1 I_32242 (I551687,I3563,I551328,I551296,);
nor I_32243 (I551718,I551670,I659012);
and I_32244 (I551735,I551718,I658991);
or I_32245 (I551752,I551735,I658994);
DFFARX1 I_32246 (I551752,I3563,I551328,I551778,);
nor I_32247 (I551786,I551778,I551402);
nor I_32248 (I551305,I551354,I551786);
not I_32249 (I551817,I551778);
nor I_32250 (I551834,I551817,I551512);
DFFARX1 I_32251 (I551834,I3563,I551328,I551311,);
nand I_32252 (I551865,I551817,I551444);
nor I_32253 (I551299,I551670,I551865);
not I_32254 (I551923,I3570);
DFFARX1 I_32255 (I740498,I3563,I551923,I551949,);
DFFARX1 I_32256 (I551949,I3563,I551923,I551966,);
not I_32257 (I551915,I551966);
DFFARX1 I_32258 (I740492,I3563,I551923,I551997,);
not I_32259 (I552005,I740489);
nor I_32260 (I552022,I551949,I552005);
not I_32261 (I552039,I740501);
not I_32262 (I552056,I740504);
nand I_32263 (I552073,I552056,I740501);
nor I_32264 (I552090,I552005,I552073);
nor I_32265 (I552107,I551997,I552090);
DFFARX1 I_32266 (I552056,I3563,I551923,I551912,);
nor I_32267 (I552138,I740504,I740513);
nand I_32268 (I552155,I552138,I740507);
nor I_32269 (I552172,I552155,I552039);
nand I_32270 (I551897,I552172,I740489);
DFFARX1 I_32271 (I552155,I3563,I551923,I551909,);
nand I_32272 (I552217,I552039,I740504);
nor I_32273 (I552234,I552039,I740504);
nand I_32274 (I551903,I552022,I552234);
not I_32275 (I552265,I740495);
nor I_32276 (I552282,I552265,I552217);
DFFARX1 I_32277 (I552282,I3563,I551923,I551891,);
nor I_32278 (I552313,I552265,I740510);
and I_32279 (I552330,I552313,I740489);
or I_32280 (I552347,I552330,I740492);
DFFARX1 I_32281 (I552347,I3563,I551923,I552373,);
nor I_32282 (I552381,I552373,I551997);
nor I_32283 (I551900,I551949,I552381);
not I_32284 (I552412,I552373);
nor I_32285 (I552429,I552412,I552107);
DFFARX1 I_32286 (I552429,I3563,I551923,I551906,);
nand I_32287 (I552460,I552412,I552039);
nor I_32288 (I551894,I552265,I552460);
not I_32289 (I552518,I3570);
DFFARX1 I_32290 (I697148,I3563,I552518,I552544,);
DFFARX1 I_32291 (I552544,I3563,I552518,I552561,);
not I_32292 (I552510,I552561);
DFFARX1 I_32293 (I697142,I3563,I552518,I552592,);
not I_32294 (I552600,I697139);
nor I_32295 (I552617,I552544,I552600);
not I_32296 (I552634,I697151);
not I_32297 (I552651,I697154);
nand I_32298 (I552668,I552651,I697151);
nor I_32299 (I552685,I552600,I552668);
nor I_32300 (I552702,I552592,I552685);
DFFARX1 I_32301 (I552651,I3563,I552518,I552507,);
nor I_32302 (I552733,I697154,I697163);
nand I_32303 (I552750,I552733,I697157);
nor I_32304 (I552767,I552750,I552634);
nand I_32305 (I552492,I552767,I697139);
DFFARX1 I_32306 (I552750,I3563,I552518,I552504,);
nand I_32307 (I552812,I552634,I697154);
nor I_32308 (I552829,I552634,I697154);
nand I_32309 (I552498,I552617,I552829);
not I_32310 (I552860,I697145);
nor I_32311 (I552877,I552860,I552812);
DFFARX1 I_32312 (I552877,I3563,I552518,I552486,);
nor I_32313 (I552908,I552860,I697160);
and I_32314 (I552925,I552908,I697139);
or I_32315 (I552942,I552925,I697142);
DFFARX1 I_32316 (I552942,I3563,I552518,I552968,);
nor I_32317 (I552976,I552968,I552592);
nor I_32318 (I552495,I552544,I552976);
not I_32319 (I553007,I552968);
nor I_32320 (I553024,I553007,I552702);
DFFARX1 I_32321 (I553024,I3563,I552518,I552501,);
nand I_32322 (I553055,I553007,I552634);
nor I_32323 (I552489,I552860,I553055);
not I_32324 (I553113,I3570);
DFFARX1 I_32325 (I857441,I3563,I553113,I553139,);
DFFARX1 I_32326 (I553139,I3563,I553113,I553156,);
not I_32327 (I553105,I553156);
DFFARX1 I_32328 (I857438,I3563,I553113,I553187,);
not I_32329 (I553195,I857438);
nor I_32330 (I553212,I553139,I553195);
not I_32331 (I553229,I857435);
not I_32332 (I553246,I857450);
nand I_32333 (I553263,I553246,I857435);
nor I_32334 (I553280,I553195,I553263);
nor I_32335 (I553297,I553187,I553280);
DFFARX1 I_32336 (I553246,I3563,I553113,I553102,);
nor I_32337 (I553328,I857450,I857444);
nand I_32338 (I553345,I553328,I857432);
nor I_32339 (I553362,I553345,I553229);
nand I_32340 (I553087,I553362,I857438);
DFFARX1 I_32341 (I553345,I3563,I553113,I553099,);
nand I_32342 (I553407,I553229,I857450);
nor I_32343 (I553424,I553229,I857450);
nand I_32344 (I553093,I553212,I553424);
not I_32345 (I553455,I857453);
nor I_32346 (I553472,I553455,I553407);
DFFARX1 I_32347 (I553472,I3563,I553113,I553081,);
nor I_32348 (I553503,I553455,I857432);
and I_32349 (I553520,I553503,I857447);
or I_32350 (I553537,I553520,I857435);
DFFARX1 I_32351 (I553537,I3563,I553113,I553563,);
nor I_32352 (I553571,I553563,I553187);
nor I_32353 (I553090,I553139,I553571);
not I_32354 (I553602,I553563);
nor I_32355 (I553619,I553602,I553297);
DFFARX1 I_32356 (I553619,I3563,I553113,I553096,);
nand I_32357 (I553650,I553602,I553229);
nor I_32358 (I553084,I553455,I553650);
not I_32359 (I553708,I3570);
DFFARX1 I_32360 (I114099,I3563,I553708,I553734,);
DFFARX1 I_32361 (I553734,I3563,I553708,I553751,);
not I_32362 (I553700,I553751);
DFFARX1 I_32363 (I114111,I3563,I553708,I553782,);
not I_32364 (I553790,I114102);
nor I_32365 (I553807,I553734,I553790);
not I_32366 (I553824,I114093);
not I_32367 (I553841,I114090);
nand I_32368 (I553858,I553841,I114093);
nor I_32369 (I553875,I553790,I553858);
nor I_32370 (I553892,I553782,I553875);
DFFARX1 I_32371 (I553841,I3563,I553708,I553697,);
nor I_32372 (I553923,I114090,I114090);
nand I_32373 (I553940,I553923,I114108);
nor I_32374 (I553957,I553940,I553824);
nand I_32375 (I553682,I553957,I114102);
DFFARX1 I_32376 (I553940,I3563,I553708,I553694,);
nand I_32377 (I554002,I553824,I114090);
nor I_32378 (I554019,I553824,I114090);
nand I_32379 (I553688,I553807,I554019);
not I_32380 (I554050,I114114);
nor I_32381 (I554067,I554050,I554002);
DFFARX1 I_32382 (I554067,I3563,I553708,I553676,);
nor I_32383 (I554098,I554050,I114093);
and I_32384 (I554115,I554098,I114096);
or I_32385 (I554132,I554115,I114105);
DFFARX1 I_32386 (I554132,I3563,I553708,I554158,);
nor I_32387 (I554166,I554158,I553782);
nor I_32388 (I553685,I553734,I554166);
not I_32389 (I554197,I554158);
nor I_32390 (I554214,I554197,I553892);
DFFARX1 I_32391 (I554214,I3563,I553708,I553691,);
nand I_32392 (I554245,I554197,I553824);
nor I_32393 (I553679,I554050,I554245);
not I_32394 (I554303,I3570);
DFFARX1 I_32395 (I1044090,I3563,I554303,I554329,);
DFFARX1 I_32396 (I554329,I3563,I554303,I554346,);
not I_32397 (I554295,I554346);
DFFARX1 I_32398 (I1044078,I3563,I554303,I554377,);
not I_32399 (I554385,I1044075);
nor I_32400 (I554402,I554329,I554385);
not I_32401 (I554419,I1044087);
not I_32402 (I554436,I1044084);
nand I_32403 (I554453,I554436,I1044087);
nor I_32404 (I554470,I554385,I554453);
nor I_32405 (I554487,I554377,I554470);
DFFARX1 I_32406 (I554436,I3563,I554303,I554292,);
nor I_32407 (I554518,I1044084,I1044093);
nand I_32408 (I554535,I554518,I1044096);
nor I_32409 (I554552,I554535,I554419);
nand I_32410 (I554277,I554552,I1044075);
DFFARX1 I_32411 (I554535,I3563,I554303,I554289,);
nand I_32412 (I554597,I554419,I1044084);
nor I_32413 (I554614,I554419,I1044084);
nand I_32414 (I554283,I554402,I554614);
not I_32415 (I554645,I1044099);
nor I_32416 (I554662,I554645,I554597);
DFFARX1 I_32417 (I554662,I3563,I554303,I554271,);
nor I_32418 (I554693,I554645,I1044102);
and I_32419 (I554710,I554693,I1044081);
or I_32420 (I554727,I554710,I1044075);
DFFARX1 I_32421 (I554727,I3563,I554303,I554753,);
nor I_32422 (I554761,I554753,I554377);
nor I_32423 (I554280,I554329,I554761);
not I_32424 (I554792,I554753);
nor I_32425 (I554809,I554792,I554487);
DFFARX1 I_32426 (I554809,I3563,I554303,I554286,);
nand I_32427 (I554840,I554792,I554419);
nor I_32428 (I554274,I554645,I554840);
not I_32429 (I554898,I3570);
DFFARX1 I_32430 (I1149969,I3563,I554898,I554924,);
DFFARX1 I_32431 (I554924,I3563,I554898,I554941,);
not I_32432 (I554890,I554941);
DFFARX1 I_32433 (I1149951,I3563,I554898,I554972,);
not I_32434 (I554980,I1149957);
nor I_32435 (I554997,I554924,I554980);
not I_32436 (I555014,I1149972);
not I_32437 (I555031,I1149963);
nand I_32438 (I555048,I555031,I1149972);
nor I_32439 (I555065,I554980,I555048);
nor I_32440 (I555082,I554972,I555065);
DFFARX1 I_32441 (I555031,I3563,I554898,I554887,);
nor I_32442 (I555113,I1149963,I1149975);
nand I_32443 (I555130,I555113,I1149954);
nor I_32444 (I555147,I555130,I555014);
nand I_32445 (I554872,I555147,I1149957);
DFFARX1 I_32446 (I555130,I3563,I554898,I554884,);
nand I_32447 (I555192,I555014,I1149963);
nor I_32448 (I555209,I555014,I1149963);
nand I_32449 (I554878,I554997,I555209);
not I_32450 (I555240,I1149960);
nor I_32451 (I555257,I555240,I555192);
DFFARX1 I_32452 (I555257,I3563,I554898,I554866,);
nor I_32453 (I555288,I555240,I1149966);
and I_32454 (I555305,I555288,I1149951);
or I_32455 (I555322,I555305,I1149954);
DFFARX1 I_32456 (I555322,I3563,I554898,I555348,);
nor I_32457 (I555356,I555348,I554972);
nor I_32458 (I554875,I554924,I555356);
not I_32459 (I555387,I555348);
nor I_32460 (I555404,I555387,I555082);
DFFARX1 I_32461 (I555404,I3563,I554898,I554881,);
nand I_32462 (I555435,I555387,I555014);
nor I_32463 (I554869,I555240,I555435);
not I_32464 (I555493,I3570);
DFFARX1 I_32465 (I464290,I3563,I555493,I555519,);
DFFARX1 I_32466 (I555519,I3563,I555493,I555536,);
not I_32467 (I555485,I555536);
DFFARX1 I_32468 (I464314,I3563,I555493,I555567,);
not I_32469 (I555575,I464293);
nor I_32470 (I555592,I555519,I555575);
not I_32471 (I555609,I464299);
not I_32472 (I555626,I464305);
nand I_32473 (I555643,I555626,I464299);
nor I_32474 (I555660,I555575,I555643);
nor I_32475 (I555677,I555567,I555660);
DFFARX1 I_32476 (I555626,I3563,I555493,I555482,);
nor I_32477 (I555708,I464305,I464317);
nand I_32478 (I555725,I555708,I464311);
nor I_32479 (I555742,I555725,I555609);
nand I_32480 (I555467,I555742,I464293);
DFFARX1 I_32481 (I555725,I3563,I555493,I555479,);
nand I_32482 (I555787,I555609,I464305);
nor I_32483 (I555804,I555609,I464305);
nand I_32484 (I555473,I555592,I555804);
not I_32485 (I555835,I464296);
nor I_32486 (I555852,I555835,I555787);
DFFARX1 I_32487 (I555852,I3563,I555493,I555461,);
nor I_32488 (I555883,I555835,I464290);
and I_32489 (I555900,I555883,I464308);
or I_32490 (I555917,I555900,I464302);
DFFARX1 I_32491 (I555917,I3563,I555493,I555943,);
nor I_32492 (I555951,I555943,I555567);
nor I_32493 (I555470,I555519,I555951);
not I_32494 (I555982,I555943);
nor I_32495 (I555999,I555982,I555677);
DFFARX1 I_32496 (I555999,I3563,I555493,I555476,);
nand I_32497 (I556030,I555982,I555609);
nor I_32498 (I555464,I555835,I556030);
not I_32499 (I556088,I3570);
DFFARX1 I_32500 (I1213549,I3563,I556088,I556114,);
DFFARX1 I_32501 (I556114,I3563,I556088,I556131,);
not I_32502 (I556080,I556131);
DFFARX1 I_32503 (I1213531,I3563,I556088,I556162,);
not I_32504 (I556170,I1213537);
nor I_32505 (I556187,I556114,I556170);
not I_32506 (I556204,I1213552);
not I_32507 (I556221,I1213543);
nand I_32508 (I556238,I556221,I1213552);
nor I_32509 (I556255,I556170,I556238);
nor I_32510 (I556272,I556162,I556255);
DFFARX1 I_32511 (I556221,I3563,I556088,I556077,);
nor I_32512 (I556303,I1213543,I1213555);
nand I_32513 (I556320,I556303,I1213534);
nor I_32514 (I556337,I556320,I556204);
nand I_32515 (I556062,I556337,I1213537);
DFFARX1 I_32516 (I556320,I3563,I556088,I556074,);
nand I_32517 (I556382,I556204,I1213543);
nor I_32518 (I556399,I556204,I1213543);
nand I_32519 (I556068,I556187,I556399);
not I_32520 (I556430,I1213540);
nor I_32521 (I556447,I556430,I556382);
DFFARX1 I_32522 (I556447,I3563,I556088,I556056,);
nor I_32523 (I556478,I556430,I1213546);
and I_32524 (I556495,I556478,I1213531);
or I_32525 (I556512,I556495,I1213534);
DFFARX1 I_32526 (I556512,I3563,I556088,I556538,);
nor I_32527 (I556546,I556538,I556162);
nor I_32528 (I556065,I556114,I556546);
not I_32529 (I556577,I556538);
nor I_32530 (I556594,I556577,I556272);
DFFARX1 I_32531 (I556594,I3563,I556088,I556071,);
nand I_32532 (I556625,I556577,I556204);
nor I_32533 (I556059,I556430,I556625);
not I_32534 (I556683,I3570);
DFFARX1 I_32535 (I712754,I3563,I556683,I556709,);
DFFARX1 I_32536 (I556709,I3563,I556683,I556726,);
not I_32537 (I556675,I556726);
DFFARX1 I_32538 (I712748,I3563,I556683,I556757,);
not I_32539 (I556765,I712745);
nor I_32540 (I556782,I556709,I556765);
not I_32541 (I556799,I712757);
not I_32542 (I556816,I712760);
nand I_32543 (I556833,I556816,I712757);
nor I_32544 (I556850,I556765,I556833);
nor I_32545 (I556867,I556757,I556850);
DFFARX1 I_32546 (I556816,I3563,I556683,I556672,);
nor I_32547 (I556898,I712760,I712769);
nand I_32548 (I556915,I556898,I712763);
nor I_32549 (I556932,I556915,I556799);
nand I_32550 (I556657,I556932,I712745);
DFFARX1 I_32551 (I556915,I3563,I556683,I556669,);
nand I_32552 (I556977,I556799,I712760);
nor I_32553 (I556994,I556799,I712760);
nand I_32554 (I556663,I556782,I556994);
not I_32555 (I557025,I712751);
nor I_32556 (I557042,I557025,I556977);
DFFARX1 I_32557 (I557042,I3563,I556683,I556651,);
nor I_32558 (I557073,I557025,I712766);
and I_32559 (I557090,I557073,I712745);
or I_32560 (I557107,I557090,I712748);
DFFARX1 I_32561 (I557107,I3563,I556683,I557133,);
nor I_32562 (I557141,I557133,I556757);
nor I_32563 (I556660,I556709,I557141);
not I_32564 (I557172,I557133);
nor I_32565 (I557189,I557172,I556867);
DFFARX1 I_32566 (I557189,I3563,I556683,I556666,);
nand I_32567 (I557220,I557172,I556799);
nor I_32568 (I556654,I557025,I557220);
not I_32569 (I557278,I3570);
DFFARX1 I_32570 (I715644,I3563,I557278,I557304,);
DFFARX1 I_32571 (I557304,I3563,I557278,I557321,);
not I_32572 (I557270,I557321);
DFFARX1 I_32573 (I715638,I3563,I557278,I557352,);
not I_32574 (I557360,I715635);
nor I_32575 (I557377,I557304,I557360);
not I_32576 (I557394,I715647);
not I_32577 (I557411,I715650);
nand I_32578 (I557428,I557411,I715647);
nor I_32579 (I557445,I557360,I557428);
nor I_32580 (I557462,I557352,I557445);
DFFARX1 I_32581 (I557411,I3563,I557278,I557267,);
nor I_32582 (I557493,I715650,I715659);
nand I_32583 (I557510,I557493,I715653);
nor I_32584 (I557527,I557510,I557394);
nand I_32585 (I557252,I557527,I715635);
DFFARX1 I_32586 (I557510,I3563,I557278,I557264,);
nand I_32587 (I557572,I557394,I715650);
nor I_32588 (I557589,I557394,I715650);
nand I_32589 (I557258,I557377,I557589);
not I_32590 (I557620,I715641);
nor I_32591 (I557637,I557620,I557572);
DFFARX1 I_32592 (I557637,I3563,I557278,I557246,);
nor I_32593 (I557668,I557620,I715656);
and I_32594 (I557685,I557668,I715635);
or I_32595 (I557702,I557685,I715638);
DFFARX1 I_32596 (I557702,I3563,I557278,I557728,);
nor I_32597 (I557736,I557728,I557352);
nor I_32598 (I557255,I557304,I557736);
not I_32599 (I557767,I557728);
nor I_32600 (I557784,I557767,I557462);
DFFARX1 I_32601 (I557784,I3563,I557278,I557261,);
nand I_32602 (I557815,I557767,I557394);
nor I_32603 (I557249,I557620,I557815);
not I_32604 (I557873,I3570);
DFFARX1 I_32605 (I498562,I3563,I557873,I557899,);
DFFARX1 I_32606 (I557899,I3563,I557873,I557916,);
not I_32607 (I557865,I557916);
DFFARX1 I_32608 (I498586,I3563,I557873,I557947,);
not I_32609 (I557955,I498565);
nor I_32610 (I557972,I557899,I557955);
not I_32611 (I557989,I498571);
not I_32612 (I558006,I498577);
nand I_32613 (I558023,I558006,I498571);
nor I_32614 (I558040,I557955,I558023);
nor I_32615 (I558057,I557947,I558040);
DFFARX1 I_32616 (I558006,I3563,I557873,I557862,);
nor I_32617 (I558088,I498577,I498589);
nand I_32618 (I558105,I558088,I498583);
nor I_32619 (I558122,I558105,I557989);
nand I_32620 (I557847,I558122,I498565);
DFFARX1 I_32621 (I558105,I3563,I557873,I557859,);
nand I_32622 (I558167,I557989,I498577);
nor I_32623 (I558184,I557989,I498577);
nand I_32624 (I557853,I557972,I558184);
not I_32625 (I558215,I498568);
nor I_32626 (I558232,I558215,I558167);
DFFARX1 I_32627 (I558232,I3563,I557873,I557841,);
nor I_32628 (I558263,I558215,I498562);
and I_32629 (I558280,I558263,I498580);
or I_32630 (I558297,I558280,I498574);
DFFARX1 I_32631 (I558297,I3563,I557873,I558323,);
nor I_32632 (I558331,I558323,I557947);
nor I_32633 (I557850,I557899,I558331);
not I_32634 (I558362,I558323);
nor I_32635 (I558379,I558362,I558057);
DFFARX1 I_32636 (I558379,I3563,I557873,I557856,);
nand I_32637 (I558410,I558362,I557989);
nor I_32638 (I557844,I558215,I558410);
not I_32639 (I558468,I3570);
DFFARX1 I_32640 (I149935,I3563,I558468,I558494,);
DFFARX1 I_32641 (I558494,I3563,I558468,I558511,);
not I_32642 (I558460,I558511);
DFFARX1 I_32643 (I149947,I3563,I558468,I558542,);
not I_32644 (I558550,I149938);
nor I_32645 (I558567,I558494,I558550);
not I_32646 (I558584,I149929);
not I_32647 (I558601,I149926);
nand I_32648 (I558618,I558601,I149929);
nor I_32649 (I558635,I558550,I558618);
nor I_32650 (I558652,I558542,I558635);
DFFARX1 I_32651 (I558601,I3563,I558468,I558457,);
nor I_32652 (I558683,I149926,I149926);
nand I_32653 (I558700,I558683,I149944);
nor I_32654 (I558717,I558700,I558584);
nand I_32655 (I558442,I558717,I149938);
DFFARX1 I_32656 (I558700,I3563,I558468,I558454,);
nand I_32657 (I558762,I558584,I149926);
nor I_32658 (I558779,I558584,I149926);
nand I_32659 (I558448,I558567,I558779);
not I_32660 (I558810,I149950);
nor I_32661 (I558827,I558810,I558762);
DFFARX1 I_32662 (I558827,I3563,I558468,I558436,);
nor I_32663 (I558858,I558810,I149929);
and I_32664 (I558875,I558858,I149932);
or I_32665 (I558892,I558875,I149941);
DFFARX1 I_32666 (I558892,I3563,I558468,I558918,);
nor I_32667 (I558926,I558918,I558542);
nor I_32668 (I558445,I558494,I558926);
not I_32669 (I558957,I558918);
nor I_32670 (I558974,I558957,I558652);
DFFARX1 I_32671 (I558974,I3563,I558468,I558451,);
nand I_32672 (I559005,I558957,I558584);
nor I_32673 (I558439,I558810,I559005);
not I_32674 (I559063,I3570);
DFFARX1 I_32675 (I1084807,I3563,I559063,I559089,);
DFFARX1 I_32676 (I559089,I3563,I559063,I559106,);
not I_32677 (I559055,I559106);
DFFARX1 I_32678 (I1084810,I3563,I559063,I559137,);
not I_32679 (I559145,I1084813);
nor I_32680 (I559162,I559089,I559145);
not I_32681 (I559179,I1084825);
not I_32682 (I559196,I1084816);
nand I_32683 (I559213,I559196,I1084825);
nor I_32684 (I559230,I559145,I559213);
nor I_32685 (I559247,I559137,I559230);
DFFARX1 I_32686 (I559196,I3563,I559063,I559052,);
nor I_32687 (I559278,I1084816,I1084822);
nand I_32688 (I559295,I559278,I1084810);
nor I_32689 (I559312,I559295,I559179);
nand I_32690 (I559037,I559312,I1084813);
DFFARX1 I_32691 (I559295,I3563,I559063,I559049,);
nand I_32692 (I559357,I559179,I1084816);
nor I_32693 (I559374,I559179,I1084816);
nand I_32694 (I559043,I559162,I559374);
not I_32695 (I559405,I1084813);
nor I_32696 (I559422,I559405,I559357);
DFFARX1 I_32697 (I559422,I3563,I559063,I559031,);
nor I_32698 (I559453,I559405,I1084819);
and I_32699 (I559470,I559453,I1084807);
or I_32700 (I559487,I559470,I1084828);
DFFARX1 I_32701 (I559487,I3563,I559063,I559513,);
nor I_32702 (I559521,I559513,I559137);
nor I_32703 (I559040,I559089,I559521);
not I_32704 (I559552,I559513);
nor I_32705 (I559569,I559552,I559247);
DFFARX1 I_32706 (I559569,I3563,I559063,I559046,);
nand I_32707 (I559600,I559552,I559179);
nor I_32708 (I559034,I559405,I559600);
not I_32709 (I559658,I3570);
DFFARX1 I_32710 (I215478,I3563,I559658,I559684,);
DFFARX1 I_32711 (I559684,I3563,I559658,I559701,);
not I_32712 (I559650,I559701);
DFFARX1 I_32713 (I215502,I3563,I559658,I559732,);
not I_32714 (I559740,I215496);
nor I_32715 (I559757,I559684,I559740);
not I_32716 (I559774,I215490);
not I_32717 (I559791,I215487);
nand I_32718 (I559808,I559791,I215490);
nor I_32719 (I559825,I559740,I559808);
nor I_32720 (I559842,I559732,I559825);
DFFARX1 I_32721 (I559791,I3563,I559658,I559647,);
nor I_32722 (I559873,I215487,I215481);
nand I_32723 (I559890,I559873,I215499);
nor I_32724 (I559907,I559890,I559774);
nand I_32725 (I559632,I559907,I215496);
DFFARX1 I_32726 (I559890,I3563,I559658,I559644,);
nand I_32727 (I559952,I559774,I215487);
nor I_32728 (I559969,I559774,I215487);
nand I_32729 (I559638,I559757,I559969);
not I_32730 (I560000,I215493);
nor I_32731 (I560017,I560000,I559952);
DFFARX1 I_32732 (I560017,I3563,I559658,I559626,);
nor I_32733 (I560048,I560000,I215478);
and I_32734 (I560065,I560048,I215484);
or I_32735 (I560082,I560065,I215481);
DFFARX1 I_32736 (I560082,I3563,I559658,I560108,);
nor I_32737 (I560116,I560108,I559732);
nor I_32738 (I559635,I559684,I560116);
not I_32739 (I560147,I560108);
nor I_32740 (I560164,I560147,I559842);
DFFARX1 I_32741 (I560164,I3563,I559658,I559641,);
nand I_32742 (I560195,I560147,I559774);
nor I_32743 (I559629,I560000,I560195);
not I_32744 (I560253,I3570);
DFFARX1 I_32745 (I224998,I3563,I560253,I560279,);
DFFARX1 I_32746 (I560279,I3563,I560253,I560296,);
not I_32747 (I560245,I560296);
DFFARX1 I_32748 (I225022,I3563,I560253,I560327,);
not I_32749 (I560335,I225016);
nor I_32750 (I560352,I560279,I560335);
not I_32751 (I560369,I225010);
not I_32752 (I560386,I225007);
nand I_32753 (I560403,I560386,I225010);
nor I_32754 (I560420,I560335,I560403);
nor I_32755 (I560437,I560327,I560420);
DFFARX1 I_32756 (I560386,I3563,I560253,I560242,);
nor I_32757 (I560468,I225007,I225001);
nand I_32758 (I560485,I560468,I225019);
nor I_32759 (I560502,I560485,I560369);
nand I_32760 (I560227,I560502,I225016);
DFFARX1 I_32761 (I560485,I3563,I560253,I560239,);
nand I_32762 (I560547,I560369,I225007);
nor I_32763 (I560564,I560369,I225007);
nand I_32764 (I560233,I560352,I560564);
not I_32765 (I560595,I225013);
nor I_32766 (I560612,I560595,I560547);
DFFARX1 I_32767 (I560612,I3563,I560253,I560221,);
nor I_32768 (I560643,I560595,I224998);
and I_32769 (I560660,I560643,I225004);
or I_32770 (I560677,I560660,I225001);
DFFARX1 I_32771 (I560677,I3563,I560253,I560703,);
nor I_32772 (I560711,I560703,I560327);
nor I_32773 (I560230,I560279,I560711);
not I_32774 (I560742,I560703);
nor I_32775 (I560759,I560742,I560437);
DFFARX1 I_32776 (I560759,I3563,I560253,I560236,);
nand I_32777 (I560790,I560742,I560369);
nor I_32778 (I560224,I560595,I560790);
not I_32779 (I560848,I3570);
DFFARX1 I_32780 (I880102,I3563,I560848,I560874,);
DFFARX1 I_32781 (I560874,I3563,I560848,I560891,);
not I_32782 (I560840,I560891);
DFFARX1 I_32783 (I880099,I3563,I560848,I560922,);
not I_32784 (I560930,I880099);
nor I_32785 (I560947,I560874,I560930);
not I_32786 (I560964,I880096);
not I_32787 (I560981,I880111);
nand I_32788 (I560998,I560981,I880096);
nor I_32789 (I561015,I560930,I560998);
nor I_32790 (I561032,I560922,I561015);
DFFARX1 I_32791 (I560981,I3563,I560848,I560837,);
nor I_32792 (I561063,I880111,I880105);
nand I_32793 (I561080,I561063,I880093);
nor I_32794 (I561097,I561080,I560964);
nand I_32795 (I560822,I561097,I880099);
DFFARX1 I_32796 (I561080,I3563,I560848,I560834,);
nand I_32797 (I561142,I560964,I880111);
nor I_32798 (I561159,I560964,I880111);
nand I_32799 (I560828,I560947,I561159);
not I_32800 (I561190,I880114);
nor I_32801 (I561207,I561190,I561142);
DFFARX1 I_32802 (I561207,I3563,I560848,I560816,);
nor I_32803 (I561238,I561190,I880093);
and I_32804 (I561255,I561238,I880108);
or I_32805 (I561272,I561255,I880096);
DFFARX1 I_32806 (I561272,I3563,I560848,I561298,);
nor I_32807 (I561306,I561298,I560922);
nor I_32808 (I560825,I560874,I561306);
not I_32809 (I561337,I561298);
nor I_32810 (I561354,I561337,I561032);
DFFARX1 I_32811 (I561354,I3563,I560848,I560831,);
nand I_32812 (I561385,I561337,I560964);
nor I_32813 (I560819,I561190,I561385);
not I_32814 (I561443,I3570);
DFFARX1 I_32815 (I319635,I3563,I561443,I561469,);
DFFARX1 I_32816 (I561469,I3563,I561443,I561486,);
not I_32817 (I561435,I561486);
DFFARX1 I_32818 (I319623,I3563,I561443,I561517,);
not I_32819 (I561525,I319626);
nor I_32820 (I561542,I561469,I561525);
not I_32821 (I561559,I319629);
not I_32822 (I561576,I319641);
nand I_32823 (I561593,I561576,I319629);
nor I_32824 (I561610,I561525,I561593);
nor I_32825 (I561627,I561517,I561610);
DFFARX1 I_32826 (I561576,I3563,I561443,I561432,);
nor I_32827 (I561658,I319641,I319632);
nand I_32828 (I561675,I561658,I319620);
nor I_32829 (I561692,I561675,I561559);
nand I_32830 (I561417,I561692,I319626);
DFFARX1 I_32831 (I561675,I3563,I561443,I561429,);
nand I_32832 (I561737,I561559,I319641);
nor I_32833 (I561754,I561559,I319641);
nand I_32834 (I561423,I561542,I561754);
not I_32835 (I561785,I319638);
nor I_32836 (I561802,I561785,I561737);
DFFARX1 I_32837 (I561802,I3563,I561443,I561411,);
nor I_32838 (I561833,I561785,I319644);
and I_32839 (I561850,I561833,I319647);
or I_32840 (I561867,I561850,I319620);
DFFARX1 I_32841 (I561867,I3563,I561443,I561893,);
nor I_32842 (I561901,I561893,I561517);
nor I_32843 (I561420,I561469,I561901);
not I_32844 (I561932,I561893);
nor I_32845 (I561949,I561932,I561627);
DFFARX1 I_32846 (I561949,I3563,I561443,I561426,);
nand I_32847 (I561980,I561932,I561559);
nor I_32848 (I561414,I561785,I561980);
not I_32849 (I562038,I3570);
DFFARX1 I_32850 (I1232623,I3563,I562038,I562064,);
DFFARX1 I_32851 (I562064,I3563,I562038,I562081,);
not I_32852 (I562030,I562081);
DFFARX1 I_32853 (I1232605,I3563,I562038,I562112,);
not I_32854 (I562120,I1232611);
nor I_32855 (I562137,I562064,I562120);
not I_32856 (I562154,I1232626);
not I_32857 (I562171,I1232617);
nand I_32858 (I562188,I562171,I1232626);
nor I_32859 (I562205,I562120,I562188);
nor I_32860 (I562222,I562112,I562205);
DFFARX1 I_32861 (I562171,I3563,I562038,I562027,);
nor I_32862 (I562253,I1232617,I1232629);
nand I_32863 (I562270,I562253,I1232608);
nor I_32864 (I562287,I562270,I562154);
nand I_32865 (I562012,I562287,I1232611);
DFFARX1 I_32866 (I562270,I3563,I562038,I562024,);
nand I_32867 (I562332,I562154,I1232617);
nor I_32868 (I562349,I562154,I1232617);
nand I_32869 (I562018,I562137,I562349);
not I_32870 (I562380,I1232614);
nor I_32871 (I562397,I562380,I562332);
DFFARX1 I_32872 (I562397,I3563,I562038,I562006,);
nor I_32873 (I562428,I562380,I1232620);
and I_32874 (I562445,I562428,I1232605);
or I_32875 (I562462,I562445,I1232608);
DFFARX1 I_32876 (I562462,I3563,I562038,I562488,);
nor I_32877 (I562496,I562488,I562112);
nor I_32878 (I562015,I562064,I562496);
not I_32879 (I562527,I562488);
nor I_32880 (I562544,I562527,I562222);
DFFARX1 I_32881 (I562544,I3563,I562038,I562021,);
nand I_32882 (I562575,I562527,I562154);
nor I_32883 (I562009,I562380,I562575);
not I_32884 (I562633,I3570);
DFFARX1 I_32885 (I609864,I3563,I562633,I562659,);
DFFARX1 I_32886 (I562659,I3563,I562633,I562676,);
not I_32887 (I562625,I562676);
DFFARX1 I_32888 (I609876,I3563,I562633,I562707,);
not I_32889 (I562715,I609861);
nor I_32890 (I562732,I562659,I562715);
not I_32891 (I562749,I609879);
not I_32892 (I562766,I609870);
nand I_32893 (I562783,I562766,I609879);
nor I_32894 (I562800,I562715,I562783);
nor I_32895 (I562817,I562707,I562800);
DFFARX1 I_32896 (I562766,I3563,I562633,I562622,);
nor I_32897 (I562848,I609870,I609882);
nand I_32898 (I562865,I562848,I609885);
nor I_32899 (I562882,I562865,I562749);
nand I_32900 (I562607,I562882,I609861);
DFFARX1 I_32901 (I562865,I3563,I562633,I562619,);
nand I_32902 (I562927,I562749,I609870);
nor I_32903 (I562944,I562749,I609870);
nand I_32904 (I562613,I562732,I562944);
not I_32905 (I562975,I609861);
nor I_32906 (I562992,I562975,I562927);
DFFARX1 I_32907 (I562992,I3563,I562633,I562601,);
nor I_32908 (I563023,I562975,I609873);
and I_32909 (I563040,I563023,I609867);
or I_32910 (I563057,I563040,I609864);
DFFARX1 I_32911 (I563057,I3563,I562633,I563083,);
nor I_32912 (I563091,I563083,I562707);
nor I_32913 (I562610,I562659,I563091);
not I_32914 (I563122,I563083);
nor I_32915 (I563139,I563122,I562817);
DFFARX1 I_32916 (I563139,I3563,I562633,I562616,);
nand I_32917 (I563170,I563122,I562749);
nor I_32918 (I562604,I562975,I563170);
not I_32919 (I563228,I3570);
DFFARX1 I_32920 (I469186,I3563,I563228,I563254,);
DFFARX1 I_32921 (I563254,I3563,I563228,I563271,);
not I_32922 (I563220,I563271);
DFFARX1 I_32923 (I469210,I3563,I563228,I563302,);
not I_32924 (I563310,I469189);
nor I_32925 (I563327,I563254,I563310);
not I_32926 (I563344,I469195);
not I_32927 (I563361,I469201);
nand I_32928 (I563378,I563361,I469195);
nor I_32929 (I563395,I563310,I563378);
nor I_32930 (I563412,I563302,I563395);
DFFARX1 I_32931 (I563361,I3563,I563228,I563217,);
nor I_32932 (I563443,I469201,I469213);
nand I_32933 (I563460,I563443,I469207);
nor I_32934 (I563477,I563460,I563344);
nand I_32935 (I563202,I563477,I469189);
DFFARX1 I_32936 (I563460,I3563,I563228,I563214,);
nand I_32937 (I563522,I563344,I469201);
nor I_32938 (I563539,I563344,I469201);
nand I_32939 (I563208,I563327,I563539);
not I_32940 (I563570,I469192);
nor I_32941 (I563587,I563570,I563522);
DFFARX1 I_32942 (I563587,I3563,I563228,I563196,);
nor I_32943 (I563618,I563570,I469186);
and I_32944 (I563635,I563618,I469204);
or I_32945 (I563652,I563635,I469198);
DFFARX1 I_32946 (I563652,I3563,I563228,I563678,);
nor I_32947 (I563686,I563678,I563302);
nor I_32948 (I563205,I563254,I563686);
not I_32949 (I563717,I563678);
nor I_32950 (I563734,I563717,I563412);
DFFARX1 I_32951 (I563734,I3563,I563228,I563211,);
nand I_32952 (I563765,I563717,I563344);
nor I_32953 (I563199,I563570,I563765);
not I_32954 (I563823,I3570);
DFFARX1 I_32955 (I705818,I3563,I563823,I563849,);
DFFARX1 I_32956 (I563849,I3563,I563823,I563866,);
not I_32957 (I563815,I563866);
DFFARX1 I_32958 (I705812,I3563,I563823,I563897,);
not I_32959 (I563905,I705809);
nor I_32960 (I563922,I563849,I563905);
not I_32961 (I563939,I705821);
not I_32962 (I563956,I705824);
nand I_32963 (I563973,I563956,I705821);
nor I_32964 (I563990,I563905,I563973);
nor I_32965 (I564007,I563897,I563990);
DFFARX1 I_32966 (I563956,I3563,I563823,I563812,);
nor I_32967 (I564038,I705824,I705833);
nand I_32968 (I564055,I564038,I705827);
nor I_32969 (I564072,I564055,I563939);
nand I_32970 (I563797,I564072,I705809);
DFFARX1 I_32971 (I564055,I3563,I563823,I563809,);
nand I_32972 (I564117,I563939,I705824);
nor I_32973 (I564134,I563939,I705824);
nand I_32974 (I563803,I563922,I564134);
not I_32975 (I564165,I705815);
nor I_32976 (I564182,I564165,I564117);
DFFARX1 I_32977 (I564182,I3563,I563823,I563791,);
nor I_32978 (I564213,I564165,I705830);
and I_32979 (I564230,I564213,I705809);
or I_32980 (I564247,I564230,I705812);
DFFARX1 I_32981 (I564247,I3563,I563823,I564273,);
nor I_32982 (I564281,I564273,I563897);
nor I_32983 (I563800,I563849,I564281);
not I_32984 (I564312,I564273);
nor I_32985 (I564329,I564312,I564007);
DFFARX1 I_32986 (I564329,I3563,I563823,I563806,);
nand I_32987 (I564360,I564312,I563939);
nor I_32988 (I563794,I564165,I564360);
not I_32989 (I564418,I3570);
DFFARX1 I_32990 (I1310304,I3563,I564418,I564444,);
DFFARX1 I_32991 (I564444,I3563,I564418,I564461,);
not I_32992 (I564410,I564461);
DFFARX1 I_32993 (I1310310,I3563,I564418,I564492,);
not I_32994 (I564500,I1310298);
nor I_32995 (I564517,I564444,I564500);
not I_32996 (I564534,I1310301);
not I_32997 (I564551,I1310307);
nand I_32998 (I564568,I564551,I1310301);
nor I_32999 (I564585,I564500,I564568);
nor I_33000 (I564602,I564492,I564585);
DFFARX1 I_33001 (I564551,I3563,I564418,I564407,);
nor I_33002 (I564633,I1310307,I1310298);
nand I_33003 (I564650,I564633,I1310316);
nor I_33004 (I564667,I564650,I564534);
nand I_33005 (I564392,I564667,I1310298);
DFFARX1 I_33006 (I564650,I3563,I564418,I564404,);
nand I_33007 (I564712,I564534,I1310307);
nor I_33008 (I564729,I564534,I1310307);
nand I_33009 (I564398,I564517,I564729);
not I_33010 (I564760,I1310295);
nor I_33011 (I564777,I564760,I564712);
DFFARX1 I_33012 (I564777,I3563,I564418,I564386,);
nor I_33013 (I564808,I564760,I1310319);
and I_33014 (I564825,I564808,I1310295);
or I_33015 (I564842,I564825,I1310313);
DFFARX1 I_33016 (I564842,I3563,I564418,I564868,);
nor I_33017 (I564876,I564868,I564492);
nor I_33018 (I564395,I564444,I564876);
not I_33019 (I564907,I564868);
nor I_33020 (I564924,I564907,I564602);
DFFARX1 I_33021 (I564924,I3563,I564418,I564401,);
nand I_33022 (I564955,I564907,I564534);
nor I_33023 (I564389,I564760,I564955);
not I_33024 (I565013,I3570);
DFFARX1 I_33025 (I309622,I3563,I565013,I565039,);
DFFARX1 I_33026 (I565039,I3563,I565013,I565056,);
not I_33027 (I565005,I565056);
DFFARX1 I_33028 (I309610,I3563,I565013,I565087,);
not I_33029 (I565095,I309613);
nor I_33030 (I565112,I565039,I565095);
not I_33031 (I565129,I309616);
not I_33032 (I565146,I309628);
nand I_33033 (I565163,I565146,I309616);
nor I_33034 (I565180,I565095,I565163);
nor I_33035 (I565197,I565087,I565180);
DFFARX1 I_33036 (I565146,I3563,I565013,I565002,);
nor I_33037 (I565228,I309628,I309619);
nand I_33038 (I565245,I565228,I309607);
nor I_33039 (I565262,I565245,I565129);
nand I_33040 (I564987,I565262,I309613);
DFFARX1 I_33041 (I565245,I3563,I565013,I564999,);
nand I_33042 (I565307,I565129,I309628);
nor I_33043 (I565324,I565129,I309628);
nand I_33044 (I564993,I565112,I565324);
not I_33045 (I565355,I309625);
nor I_33046 (I565372,I565355,I565307);
DFFARX1 I_33047 (I565372,I3563,I565013,I564981,);
nor I_33048 (I565403,I565355,I309631);
and I_33049 (I565420,I565403,I309634);
or I_33050 (I565437,I565420,I309607);
DFFARX1 I_33051 (I565437,I3563,I565013,I565463,);
nor I_33052 (I565471,I565463,I565087);
nor I_33053 (I564990,I565039,I565471);
not I_33054 (I565502,I565463);
nor I_33055 (I565519,I565502,I565197);
DFFARX1 I_33056 (I565519,I3563,I565013,I564996,);
nand I_33057 (I565550,I565502,I565129);
nor I_33058 (I564984,I565355,I565550);
not I_33059 (I565608,I3570);
DFFARX1 I_33060 (I964632,I3563,I565608,I565634,);
DFFARX1 I_33061 (I565634,I3563,I565608,I565651,);
not I_33062 (I565600,I565651);
DFFARX1 I_33063 (I964620,I3563,I565608,I565682,);
not I_33064 (I565690,I964617);
nor I_33065 (I565707,I565634,I565690);
not I_33066 (I565724,I964629);
not I_33067 (I565741,I964626);
nand I_33068 (I565758,I565741,I964629);
nor I_33069 (I565775,I565690,I565758);
nor I_33070 (I565792,I565682,I565775);
DFFARX1 I_33071 (I565741,I3563,I565608,I565597,);
nor I_33072 (I565823,I964626,I964635);
nand I_33073 (I565840,I565823,I964638);
nor I_33074 (I565857,I565840,I565724);
nand I_33075 (I565582,I565857,I964617);
DFFARX1 I_33076 (I565840,I3563,I565608,I565594,);
nand I_33077 (I565902,I565724,I964626);
nor I_33078 (I565919,I565724,I964626);
nand I_33079 (I565588,I565707,I565919);
not I_33080 (I565950,I964641);
nor I_33081 (I565967,I565950,I565902);
DFFARX1 I_33082 (I565967,I3563,I565608,I565576,);
nor I_33083 (I565998,I565950,I964644);
and I_33084 (I566015,I565998,I964623);
or I_33085 (I566032,I566015,I964617);
DFFARX1 I_33086 (I566032,I3563,I565608,I566058,);
nor I_33087 (I566066,I566058,I565682);
nor I_33088 (I565585,I565634,I566066);
not I_33089 (I566097,I566058);
nor I_33090 (I566114,I566097,I565792);
DFFARX1 I_33091 (I566114,I3563,I565608,I565591,);
nand I_33092 (I566145,I566097,I565724);
nor I_33093 (I565579,I565950,I566145);
not I_33094 (I566203,I3570);
DFFARX1 I_33095 (I290650,I3563,I566203,I566229,);
DFFARX1 I_33096 (I566229,I3563,I566203,I566246,);
not I_33097 (I566195,I566246);
DFFARX1 I_33098 (I290638,I3563,I566203,I566277,);
not I_33099 (I566285,I290641);
nor I_33100 (I566302,I566229,I566285);
not I_33101 (I566319,I290644);
not I_33102 (I566336,I290656);
nand I_33103 (I566353,I566336,I290644);
nor I_33104 (I566370,I566285,I566353);
nor I_33105 (I566387,I566277,I566370);
DFFARX1 I_33106 (I566336,I3563,I566203,I566192,);
nor I_33107 (I566418,I290656,I290647);
nand I_33108 (I566435,I566418,I290635);
nor I_33109 (I566452,I566435,I566319);
nand I_33110 (I566177,I566452,I290641);
DFFARX1 I_33111 (I566435,I3563,I566203,I566189,);
nand I_33112 (I566497,I566319,I290656);
nor I_33113 (I566514,I566319,I290656);
nand I_33114 (I566183,I566302,I566514);
not I_33115 (I566545,I290653);
nor I_33116 (I566562,I566545,I566497);
DFFARX1 I_33117 (I566562,I3563,I566203,I566171,);
nor I_33118 (I566593,I566545,I290659);
and I_33119 (I566610,I566593,I290662);
or I_33120 (I566627,I566610,I290635);
DFFARX1 I_33121 (I566627,I3563,I566203,I566653,);
nor I_33122 (I566661,I566653,I566277);
nor I_33123 (I566180,I566229,I566661);
not I_33124 (I566692,I566653);
nor I_33125 (I566709,I566692,I566387);
DFFARX1 I_33126 (I566709,I3563,I566203,I566186,);
nand I_33127 (I566740,I566692,I566319);
nor I_33128 (I566174,I566545,I566740);
not I_33129 (I566798,I3570);
DFFARX1 I_33130 (I667670,I3563,I566798,I566824,);
DFFARX1 I_33131 (I566824,I3563,I566798,I566841,);
not I_33132 (I566790,I566841);
DFFARX1 I_33133 (I667664,I3563,I566798,I566872,);
not I_33134 (I566880,I667661);
nor I_33135 (I566897,I566824,I566880);
not I_33136 (I566914,I667673);
not I_33137 (I566931,I667676);
nand I_33138 (I566948,I566931,I667673);
nor I_33139 (I566965,I566880,I566948);
nor I_33140 (I566982,I566872,I566965);
DFFARX1 I_33141 (I566931,I3563,I566798,I566787,);
nor I_33142 (I567013,I667676,I667685);
nand I_33143 (I567030,I567013,I667679);
nor I_33144 (I567047,I567030,I566914);
nand I_33145 (I566772,I567047,I667661);
DFFARX1 I_33146 (I567030,I3563,I566798,I566784,);
nand I_33147 (I567092,I566914,I667676);
nor I_33148 (I567109,I566914,I667676);
nand I_33149 (I566778,I566897,I567109);
not I_33150 (I567140,I667667);
nor I_33151 (I567157,I567140,I567092);
DFFARX1 I_33152 (I567157,I3563,I566798,I566766,);
nor I_33153 (I567188,I567140,I667682);
and I_33154 (I567205,I567188,I667661);
or I_33155 (I567222,I567205,I667664);
DFFARX1 I_33156 (I567222,I3563,I566798,I567248,);
nor I_33157 (I567256,I567248,I566872);
nor I_33158 (I566775,I566824,I567256);
not I_33159 (I567287,I567248);
nor I_33160 (I567304,I567287,I566982);
DFFARX1 I_33161 (I567304,I3563,I566798,I566781,);
nand I_33162 (I567335,I567287,I566914);
nor I_33163 (I566769,I567140,I567335);
not I_33164 (I567393,I3570);
DFFARX1 I_33165 (I310149,I3563,I567393,I567419,);
DFFARX1 I_33166 (I567419,I3563,I567393,I567436,);
not I_33167 (I567385,I567436);
DFFARX1 I_33168 (I310137,I3563,I567393,I567467,);
not I_33169 (I567475,I310140);
nor I_33170 (I567492,I567419,I567475);
not I_33171 (I567509,I310143);
not I_33172 (I567526,I310155);
nand I_33173 (I567543,I567526,I310143);
nor I_33174 (I567560,I567475,I567543);
nor I_33175 (I567577,I567467,I567560);
DFFARX1 I_33176 (I567526,I3563,I567393,I567382,);
nor I_33177 (I567608,I310155,I310146);
nand I_33178 (I567625,I567608,I310134);
nor I_33179 (I567642,I567625,I567509);
nand I_33180 (I567367,I567642,I310140);
DFFARX1 I_33181 (I567625,I3563,I567393,I567379,);
nand I_33182 (I567687,I567509,I310155);
nor I_33183 (I567704,I567509,I310155);
nand I_33184 (I567373,I567492,I567704);
not I_33185 (I567735,I310152);
nor I_33186 (I567752,I567735,I567687);
DFFARX1 I_33187 (I567752,I3563,I567393,I567361,);
nor I_33188 (I567783,I567735,I310158);
and I_33189 (I567800,I567783,I310161);
or I_33190 (I567817,I567800,I310134);
DFFARX1 I_33191 (I567817,I3563,I567393,I567843,);
nor I_33192 (I567851,I567843,I567467);
nor I_33193 (I567370,I567419,I567851);
not I_33194 (I567882,I567843);
nor I_33195 (I567899,I567882,I567577);
DFFARX1 I_33196 (I567899,I3563,I567393,I567376,);
nand I_33197 (I567930,I567882,I567509);
nor I_33198 (I567364,I567735,I567930);
not I_33199 (I567988,I3570);
DFFARX1 I_33200 (I960110,I3563,I567988,I568014,);
DFFARX1 I_33201 (I568014,I3563,I567988,I568031,);
not I_33202 (I567980,I568031);
DFFARX1 I_33203 (I960098,I3563,I567988,I568062,);
not I_33204 (I568070,I960095);
nor I_33205 (I568087,I568014,I568070);
not I_33206 (I568104,I960107);
not I_33207 (I568121,I960104);
nand I_33208 (I568138,I568121,I960107);
nor I_33209 (I568155,I568070,I568138);
nor I_33210 (I568172,I568062,I568155);
DFFARX1 I_33211 (I568121,I3563,I567988,I567977,);
nor I_33212 (I568203,I960104,I960113);
nand I_33213 (I568220,I568203,I960116);
nor I_33214 (I568237,I568220,I568104);
nand I_33215 (I567962,I568237,I960095);
DFFARX1 I_33216 (I568220,I3563,I567988,I567974,);
nand I_33217 (I568282,I568104,I960104);
nor I_33218 (I568299,I568104,I960104);
nand I_33219 (I567968,I568087,I568299);
not I_33220 (I568330,I960119);
nor I_33221 (I568347,I568330,I568282);
DFFARX1 I_33222 (I568347,I3563,I567988,I567956,);
nor I_33223 (I568378,I568330,I960122);
and I_33224 (I568395,I568378,I960101);
or I_33225 (I568412,I568395,I960095);
DFFARX1 I_33226 (I568412,I3563,I567988,I568438,);
nor I_33227 (I568446,I568438,I568062);
nor I_33228 (I567965,I568014,I568446);
not I_33229 (I568477,I568438);
nor I_33230 (I568494,I568477,I568172);
DFFARX1 I_33231 (I568494,I3563,I567988,I567971,);
nand I_33232 (I568525,I568477,I568104);
nor I_33233 (I567959,I568330,I568525);
not I_33234 (I568583,I3570);
DFFARX1 I_33235 (I761884,I3563,I568583,I568609,);
DFFARX1 I_33236 (I568609,I3563,I568583,I568626,);
not I_33237 (I568575,I568626);
DFFARX1 I_33238 (I761878,I3563,I568583,I568657,);
not I_33239 (I568665,I761875);
nor I_33240 (I568682,I568609,I568665);
not I_33241 (I568699,I761887);
not I_33242 (I568716,I761890);
nand I_33243 (I568733,I568716,I761887);
nor I_33244 (I568750,I568665,I568733);
nor I_33245 (I568767,I568657,I568750);
DFFARX1 I_33246 (I568716,I3563,I568583,I568572,);
nor I_33247 (I568798,I761890,I761899);
nand I_33248 (I568815,I568798,I761893);
nor I_33249 (I568832,I568815,I568699);
nand I_33250 (I568557,I568832,I761875);
DFFARX1 I_33251 (I568815,I3563,I568583,I568569,);
nand I_33252 (I568877,I568699,I761890);
nor I_33253 (I568894,I568699,I761890);
nand I_33254 (I568563,I568682,I568894);
not I_33255 (I568925,I761881);
nor I_33256 (I568942,I568925,I568877);
DFFARX1 I_33257 (I568942,I3563,I568583,I568551,);
nor I_33258 (I568973,I568925,I761896);
and I_33259 (I568990,I568973,I761875);
or I_33260 (I569007,I568990,I761878);
DFFARX1 I_33261 (I569007,I3563,I568583,I569033,);
nor I_33262 (I569041,I569033,I568657);
nor I_33263 (I568560,I568609,I569041);
not I_33264 (I569072,I569033);
nor I_33265 (I569089,I569072,I568767);
DFFARX1 I_33266 (I569089,I3563,I568583,I568566,);
nand I_33267 (I569120,I569072,I568699);
nor I_33268 (I568554,I568925,I569120);
not I_33269 (I569178,I3570);
DFFARX1 I_33270 (I1244183,I3563,I569178,I569204,);
DFFARX1 I_33271 (I569204,I3563,I569178,I569221,);
not I_33272 (I569170,I569221);
DFFARX1 I_33273 (I1244165,I3563,I569178,I569252,);
not I_33274 (I569260,I1244171);
nor I_33275 (I569277,I569204,I569260);
not I_33276 (I569294,I1244186);
not I_33277 (I569311,I1244177);
nand I_33278 (I569328,I569311,I1244186);
nor I_33279 (I569345,I569260,I569328);
nor I_33280 (I569362,I569252,I569345);
DFFARX1 I_33281 (I569311,I3563,I569178,I569167,);
nor I_33282 (I569393,I1244177,I1244189);
nand I_33283 (I569410,I569393,I1244168);
nor I_33284 (I569427,I569410,I569294);
nand I_33285 (I569152,I569427,I1244171);
DFFARX1 I_33286 (I569410,I3563,I569178,I569164,);
nand I_33287 (I569472,I569294,I1244177);
nor I_33288 (I569489,I569294,I1244177);
nand I_33289 (I569158,I569277,I569489);
not I_33290 (I569520,I1244174);
nor I_33291 (I569537,I569520,I569472);
DFFARX1 I_33292 (I569537,I3563,I569178,I569146,);
nor I_33293 (I569568,I569520,I1244180);
and I_33294 (I569585,I569568,I1244165);
or I_33295 (I569602,I569585,I1244168);
DFFARX1 I_33296 (I569602,I3563,I569178,I569628,);
nor I_33297 (I569636,I569628,I569252);
nor I_33298 (I569155,I569204,I569636);
not I_33299 (I569667,I569628);
nor I_33300 (I569684,I569667,I569362);
DFFARX1 I_33301 (I569684,I3563,I569178,I569161,);
nand I_33302 (I569715,I569667,I569294);
nor I_33303 (I569149,I569520,I569715);
not I_33304 (I569773,I3570);
DFFARX1 I_33305 (I1020188,I3563,I569773,I569799,);
DFFARX1 I_33306 (I569799,I3563,I569773,I569816,);
not I_33307 (I569765,I569816);
DFFARX1 I_33308 (I1020176,I3563,I569773,I569847,);
not I_33309 (I569855,I1020173);
nor I_33310 (I569872,I569799,I569855);
not I_33311 (I569889,I1020185);
not I_33312 (I569906,I1020182);
nand I_33313 (I569923,I569906,I1020185);
nor I_33314 (I569940,I569855,I569923);
nor I_33315 (I569957,I569847,I569940);
DFFARX1 I_33316 (I569906,I3563,I569773,I569762,);
nor I_33317 (I569988,I1020182,I1020191);
nand I_33318 (I570005,I569988,I1020194);
nor I_33319 (I570022,I570005,I569889);
nand I_33320 (I569747,I570022,I1020173);
DFFARX1 I_33321 (I570005,I3563,I569773,I569759,);
nand I_33322 (I570067,I569889,I1020182);
nor I_33323 (I570084,I569889,I1020182);
nand I_33324 (I569753,I569872,I570084);
not I_33325 (I570115,I1020197);
nor I_33326 (I570132,I570115,I570067);
DFFARX1 I_33327 (I570132,I3563,I569773,I569741,);
nor I_33328 (I570163,I570115,I1020200);
and I_33329 (I570180,I570163,I1020179);
or I_33330 (I570197,I570180,I1020173);
DFFARX1 I_33331 (I570197,I3563,I569773,I570223,);
nor I_33332 (I570231,I570223,I569847);
nor I_33333 (I569750,I569799,I570231);
not I_33334 (I570262,I570223);
nor I_33335 (I570279,I570262,I569957);
DFFARX1 I_33336 (I570279,I3563,I569773,I569756,);
nand I_33337 (I570310,I570262,I569889);
nor I_33338 (I569744,I570115,I570310);
not I_33339 (I570368,I3570);
DFFARX1 I_33340 (I339134,I3563,I570368,I570394,);
DFFARX1 I_33341 (I570394,I3563,I570368,I570411,);
not I_33342 (I570360,I570411);
DFFARX1 I_33343 (I339122,I3563,I570368,I570442,);
not I_33344 (I570450,I339125);
nor I_33345 (I570467,I570394,I570450);
not I_33346 (I570484,I339128);
not I_33347 (I570501,I339140);
nand I_33348 (I570518,I570501,I339128);
nor I_33349 (I570535,I570450,I570518);
nor I_33350 (I570552,I570442,I570535);
DFFARX1 I_33351 (I570501,I3563,I570368,I570357,);
nor I_33352 (I570583,I339140,I339131);
nand I_33353 (I570600,I570583,I339119);
nor I_33354 (I570617,I570600,I570484);
nand I_33355 (I570342,I570617,I339125);
DFFARX1 I_33356 (I570600,I3563,I570368,I570354,);
nand I_33357 (I570662,I570484,I339140);
nor I_33358 (I570679,I570484,I339140);
nand I_33359 (I570348,I570467,I570679);
not I_33360 (I570710,I339137);
nor I_33361 (I570727,I570710,I570662);
DFFARX1 I_33362 (I570727,I3563,I570368,I570336,);
nor I_33363 (I570758,I570710,I339143);
and I_33364 (I570775,I570758,I339146);
or I_33365 (I570792,I570775,I339119);
DFFARX1 I_33366 (I570792,I3563,I570368,I570818,);
nor I_33367 (I570826,I570818,I570442);
nor I_33368 (I570345,I570394,I570826);
not I_33369 (I570857,I570818);
nor I_33370 (I570874,I570857,I570552);
DFFARX1 I_33371 (I570874,I3563,I570368,I570351,);
nand I_33372 (I570905,I570857,I570484);
nor I_33373 (I570339,I570710,I570905);
not I_33374 (I570963,I3570);
DFFARX1 I_33375 (I809280,I3563,I570963,I570989,);
DFFARX1 I_33376 (I570989,I3563,I570963,I571006,);
not I_33377 (I570955,I571006);
DFFARX1 I_33378 (I809274,I3563,I570963,I571037,);
not I_33379 (I571045,I809271);
nor I_33380 (I571062,I570989,I571045);
not I_33381 (I571079,I809283);
not I_33382 (I571096,I809286);
nand I_33383 (I571113,I571096,I809283);
nor I_33384 (I571130,I571045,I571113);
nor I_33385 (I571147,I571037,I571130);
DFFARX1 I_33386 (I571096,I3563,I570963,I570952,);
nor I_33387 (I571178,I809286,I809295);
nand I_33388 (I571195,I571178,I809289);
nor I_33389 (I571212,I571195,I571079);
nand I_33390 (I570937,I571212,I809271);
DFFARX1 I_33391 (I571195,I3563,I570963,I570949,);
nand I_33392 (I571257,I571079,I809286);
nor I_33393 (I571274,I571079,I809286);
nand I_33394 (I570943,I571062,I571274);
not I_33395 (I571305,I809277);
nor I_33396 (I571322,I571305,I571257);
DFFARX1 I_33397 (I571322,I3563,I570963,I570931,);
nor I_33398 (I571353,I571305,I809292);
and I_33399 (I571370,I571353,I809271);
or I_33400 (I571387,I571370,I809274);
DFFARX1 I_33401 (I571387,I3563,I570963,I571413,);
nor I_33402 (I571421,I571413,I571037);
nor I_33403 (I570940,I570989,I571421);
not I_33404 (I571452,I571413);
nor I_33405 (I571469,I571452,I571147);
DFFARX1 I_33406 (I571469,I3563,I570963,I570946,);
nand I_33407 (I571500,I571452,I571079);
nor I_33408 (I570934,I571305,I571500);
not I_33409 (I571558,I3570);
DFFARX1 I_33410 (I1042798,I3563,I571558,I571584,);
DFFARX1 I_33411 (I571584,I3563,I571558,I571601,);
not I_33412 (I571550,I571601);
DFFARX1 I_33413 (I1042786,I3563,I571558,I571632,);
not I_33414 (I571640,I1042783);
nor I_33415 (I571657,I571584,I571640);
not I_33416 (I571674,I1042795);
not I_33417 (I571691,I1042792);
nand I_33418 (I571708,I571691,I1042795);
nor I_33419 (I571725,I571640,I571708);
nor I_33420 (I571742,I571632,I571725);
DFFARX1 I_33421 (I571691,I3563,I571558,I571547,);
nor I_33422 (I571773,I1042792,I1042801);
nand I_33423 (I571790,I571773,I1042804);
nor I_33424 (I571807,I571790,I571674);
nand I_33425 (I571532,I571807,I1042783);
DFFARX1 I_33426 (I571790,I3563,I571558,I571544,);
nand I_33427 (I571852,I571674,I1042792);
nor I_33428 (I571869,I571674,I1042792);
nand I_33429 (I571538,I571657,I571869);
not I_33430 (I571900,I1042807);
nor I_33431 (I571917,I571900,I571852);
DFFARX1 I_33432 (I571917,I3563,I571558,I571526,);
nor I_33433 (I571948,I571900,I1042810);
and I_33434 (I571965,I571948,I1042789);
or I_33435 (I571982,I571965,I1042783);
DFFARX1 I_33436 (I571982,I3563,I571558,I572008,);
nor I_33437 (I572016,I572008,I571632);
nor I_33438 (I571535,I571584,I572016);
not I_33439 (I572047,I572008);
nor I_33440 (I572064,I572047,I571742);
DFFARX1 I_33441 (I572064,I3563,I571558,I571541,);
nand I_33442 (I572095,I572047,I571674);
nor I_33443 (I571529,I571900,I572095);
not I_33444 (I572153,I3570);
DFFARX1 I_33445 (I177993,I3563,I572153,I572179,);
DFFARX1 I_33446 (I572179,I3563,I572153,I572196,);
not I_33447 (I572145,I572196);
DFFARX1 I_33448 (I178017,I3563,I572153,I572227,);
not I_33449 (I572235,I178011);
nor I_33450 (I572252,I572179,I572235);
not I_33451 (I572269,I178005);
not I_33452 (I572286,I178002);
nand I_33453 (I572303,I572286,I178005);
nor I_33454 (I572320,I572235,I572303);
nor I_33455 (I572337,I572227,I572320);
DFFARX1 I_33456 (I572286,I3563,I572153,I572142,);
nor I_33457 (I572368,I178002,I177996);
nand I_33458 (I572385,I572368,I178014);
nor I_33459 (I572402,I572385,I572269);
nand I_33460 (I572127,I572402,I178011);
DFFARX1 I_33461 (I572385,I3563,I572153,I572139,);
nand I_33462 (I572447,I572269,I178002);
nor I_33463 (I572464,I572269,I178002);
nand I_33464 (I572133,I572252,I572464);
not I_33465 (I572495,I178008);
nor I_33466 (I572512,I572495,I572447);
DFFARX1 I_33467 (I572512,I3563,I572153,I572121,);
nor I_33468 (I572543,I572495,I177993);
and I_33469 (I572560,I572543,I177999);
or I_33470 (I572577,I572560,I177996);
DFFARX1 I_33471 (I572577,I3563,I572153,I572603,);
nor I_33472 (I572611,I572603,I572227);
nor I_33473 (I572130,I572179,I572611);
not I_33474 (I572642,I572603);
nor I_33475 (I572659,I572642,I572337);
DFFARX1 I_33476 (I572659,I3563,I572153,I572136,);
nand I_33477 (I572690,I572642,I572269);
nor I_33478 (I572124,I572495,I572690);
not I_33479 (I572748,I3570);
DFFARX1 I_33480 (I1261097,I3563,I572748,I572774,);
DFFARX1 I_33481 (I572774,I3563,I572748,I572791,);
not I_33482 (I572740,I572791);
DFFARX1 I_33483 (I1261112,I3563,I572748,I572822,);
not I_33484 (I572830,I1261121);
nor I_33485 (I572847,I572774,I572830);
not I_33486 (I572864,I1261100);
not I_33487 (I572881,I1261106);
nand I_33488 (I572898,I572881,I1261100);
nor I_33489 (I572915,I572830,I572898);
nor I_33490 (I572932,I572822,I572915);
DFFARX1 I_33491 (I572881,I3563,I572748,I572737,);
nor I_33492 (I572963,I1261106,I1261118);
nand I_33493 (I572980,I572963,I1261115);
nor I_33494 (I572997,I572980,I572864);
nand I_33495 (I572722,I572997,I1261121);
DFFARX1 I_33496 (I572980,I3563,I572748,I572734,);
nand I_33497 (I573042,I572864,I1261106);
nor I_33498 (I573059,I572864,I1261106);
nand I_33499 (I572728,I572847,I573059);
not I_33500 (I573090,I1261097);
nor I_33501 (I573107,I573090,I573042);
DFFARX1 I_33502 (I573107,I3563,I572748,I572716,);
nor I_33503 (I573138,I573090,I1261109);
and I_33504 (I573155,I573138,I1261103);
or I_33505 (I573172,I573155,I1261100);
DFFARX1 I_33506 (I573172,I3563,I572748,I573198,);
nor I_33507 (I573206,I573198,I572822);
nor I_33508 (I572725,I572774,I573206);
not I_33509 (I573237,I573198);
nor I_33510 (I573254,I573237,I572932);
DFFARX1 I_33511 (I573254,I3563,I572748,I572731,);
nand I_33512 (I573285,I573237,I572864);
nor I_33513 (I572719,I573090,I573285);
not I_33514 (I573343,I3570);
DFFARX1 I_33515 (I402901,I3563,I573343,I573369,);
DFFARX1 I_33516 (I573369,I3563,I573343,I573386,);
not I_33517 (I573335,I573386);
DFFARX1 I_33518 (I402889,I3563,I573343,I573417,);
not I_33519 (I573425,I402892);
nor I_33520 (I573442,I573369,I573425);
not I_33521 (I573459,I402895);
not I_33522 (I573476,I402907);
nand I_33523 (I573493,I573476,I402895);
nor I_33524 (I573510,I573425,I573493);
nor I_33525 (I573527,I573417,I573510);
DFFARX1 I_33526 (I573476,I3563,I573343,I573332,);
nor I_33527 (I573558,I402907,I402898);
nand I_33528 (I573575,I573558,I402886);
nor I_33529 (I573592,I573575,I573459);
nand I_33530 (I573317,I573592,I402892);
DFFARX1 I_33531 (I573575,I3563,I573343,I573329,);
nand I_33532 (I573637,I573459,I402907);
nor I_33533 (I573654,I573459,I402907);
nand I_33534 (I573323,I573442,I573654);
not I_33535 (I573685,I402904);
nor I_33536 (I573702,I573685,I573637);
DFFARX1 I_33537 (I573702,I3563,I573343,I573311,);
nor I_33538 (I573733,I573685,I402910);
and I_33539 (I573750,I573733,I402913);
or I_33540 (I573767,I573750,I402886);
DFFARX1 I_33541 (I573767,I3563,I573343,I573793,);
nor I_33542 (I573801,I573793,I573417);
nor I_33543 (I573320,I573369,I573801);
not I_33544 (I573832,I573793);
nor I_33545 (I573849,I573832,I573527);
DFFARX1 I_33546 (I573849,I3563,I573343,I573326,);
nand I_33547 (I573880,I573832,I573459);
nor I_33548 (I573314,I573685,I573880);
not I_33549 (I573938,I3570);
DFFARX1 I_33550 (I194058,I3563,I573938,I573964,);
DFFARX1 I_33551 (I573964,I3563,I573938,I573981,);
not I_33552 (I573930,I573981);
DFFARX1 I_33553 (I194082,I3563,I573938,I574012,);
not I_33554 (I574020,I194076);
nor I_33555 (I574037,I573964,I574020);
not I_33556 (I574054,I194070);
not I_33557 (I574071,I194067);
nand I_33558 (I574088,I574071,I194070);
nor I_33559 (I574105,I574020,I574088);
nor I_33560 (I574122,I574012,I574105);
DFFARX1 I_33561 (I574071,I3563,I573938,I573927,);
nor I_33562 (I574153,I194067,I194061);
nand I_33563 (I574170,I574153,I194079);
nor I_33564 (I574187,I574170,I574054);
nand I_33565 (I573912,I574187,I194076);
DFFARX1 I_33566 (I574170,I3563,I573938,I573924,);
nand I_33567 (I574232,I574054,I194067);
nor I_33568 (I574249,I574054,I194067);
nand I_33569 (I573918,I574037,I574249);
not I_33570 (I574280,I194073);
nor I_33571 (I574297,I574280,I574232);
DFFARX1 I_33572 (I574297,I3563,I573938,I573906,);
nor I_33573 (I574328,I574280,I194058);
and I_33574 (I574345,I574328,I194064);
or I_33575 (I574362,I574345,I194061);
DFFARX1 I_33576 (I574362,I3563,I573938,I574388,);
nor I_33577 (I574396,I574388,I574012);
nor I_33578 (I573915,I573964,I574396);
not I_33579 (I574427,I574388);
nor I_33580 (I574444,I574427,I574122);
DFFARX1 I_33581 (I574444,I3563,I573938,I573921,);
nand I_33582 (I574475,I574427,I574054);
nor I_33583 (I573909,I574280,I574475);
not I_33584 (I574533,I3570);
DFFARX1 I_33585 (I931686,I3563,I574533,I574559,);
DFFARX1 I_33586 (I574559,I3563,I574533,I574576,);
not I_33587 (I574525,I574576);
DFFARX1 I_33588 (I931674,I3563,I574533,I574607,);
not I_33589 (I574615,I931671);
nor I_33590 (I574632,I574559,I574615);
not I_33591 (I574649,I931683);
not I_33592 (I574666,I931680);
nand I_33593 (I574683,I574666,I931683);
nor I_33594 (I574700,I574615,I574683);
nor I_33595 (I574717,I574607,I574700);
DFFARX1 I_33596 (I574666,I3563,I574533,I574522,);
nor I_33597 (I574748,I931680,I931689);
nand I_33598 (I574765,I574748,I931692);
nor I_33599 (I574782,I574765,I574649);
nand I_33600 (I574507,I574782,I931671);
DFFARX1 I_33601 (I574765,I3563,I574533,I574519,);
nand I_33602 (I574827,I574649,I931680);
nor I_33603 (I574844,I574649,I931680);
nand I_33604 (I574513,I574632,I574844);
not I_33605 (I574875,I931695);
nor I_33606 (I574892,I574875,I574827);
DFFARX1 I_33607 (I574892,I3563,I574533,I574501,);
nor I_33608 (I574923,I574875,I931698);
and I_33609 (I574940,I574923,I931677);
or I_33610 (I574957,I574940,I931671);
DFFARX1 I_33611 (I574957,I3563,I574533,I574983,);
nor I_33612 (I574991,I574983,I574607);
nor I_33613 (I574510,I574559,I574991);
not I_33614 (I575022,I574983);
nor I_33615 (I575039,I575022,I574717);
DFFARX1 I_33616 (I575039,I3563,I574533,I574516,);
nand I_33617 (I575070,I575022,I574649);
nor I_33618 (I574504,I574875,I575070);
not I_33619 (I575128,I3570);
DFFARX1 I_33620 (I1203723,I3563,I575128,I575154,);
DFFARX1 I_33621 (I575154,I3563,I575128,I575171,);
not I_33622 (I575120,I575171);
DFFARX1 I_33623 (I1203705,I3563,I575128,I575202,);
not I_33624 (I575210,I1203711);
nor I_33625 (I575227,I575154,I575210);
not I_33626 (I575244,I1203726);
not I_33627 (I575261,I1203717);
nand I_33628 (I575278,I575261,I1203726);
nor I_33629 (I575295,I575210,I575278);
nor I_33630 (I575312,I575202,I575295);
DFFARX1 I_33631 (I575261,I3563,I575128,I575117,);
nor I_33632 (I575343,I1203717,I1203729);
nand I_33633 (I575360,I575343,I1203708);
nor I_33634 (I575377,I575360,I575244);
nand I_33635 (I575102,I575377,I1203711);
DFFARX1 I_33636 (I575360,I3563,I575128,I575114,);
nand I_33637 (I575422,I575244,I1203717);
nor I_33638 (I575439,I575244,I1203717);
nand I_33639 (I575108,I575227,I575439);
not I_33640 (I575470,I1203714);
nor I_33641 (I575487,I575470,I575422);
DFFARX1 I_33642 (I575487,I3563,I575128,I575096,);
nor I_33643 (I575518,I575470,I1203720);
and I_33644 (I575535,I575518,I1203705);
or I_33645 (I575552,I575535,I1203708);
DFFARX1 I_33646 (I575552,I3563,I575128,I575578,);
nor I_33647 (I575586,I575578,I575202);
nor I_33648 (I575105,I575154,I575586);
not I_33649 (I575617,I575578);
nor I_33650 (I575634,I575617,I575312);
DFFARX1 I_33651 (I575634,I3563,I575128,I575111,);
nand I_33652 (I575665,I575617,I575244);
nor I_33653 (I575099,I575470,I575665);
not I_33654 (I575723,I3570);
DFFARX1 I_33655 (I508898,I3563,I575723,I575749,);
DFFARX1 I_33656 (I575749,I3563,I575723,I575766,);
not I_33657 (I575715,I575766);
DFFARX1 I_33658 (I508922,I3563,I575723,I575797,);
not I_33659 (I575805,I508901);
nor I_33660 (I575822,I575749,I575805);
not I_33661 (I575839,I508907);
not I_33662 (I575856,I508913);
nand I_33663 (I575873,I575856,I508907);
nor I_33664 (I575890,I575805,I575873);
nor I_33665 (I575907,I575797,I575890);
DFFARX1 I_33666 (I575856,I3563,I575723,I575712,);
nor I_33667 (I575938,I508913,I508925);
nand I_33668 (I575955,I575938,I508919);
nor I_33669 (I575972,I575955,I575839);
nand I_33670 (I575697,I575972,I508901);
DFFARX1 I_33671 (I575955,I3563,I575723,I575709,);
nand I_33672 (I576017,I575839,I508913);
nor I_33673 (I576034,I575839,I508913);
nand I_33674 (I575703,I575822,I576034);
not I_33675 (I576065,I508904);
nor I_33676 (I576082,I576065,I576017);
DFFARX1 I_33677 (I576082,I3563,I575723,I575691,);
nor I_33678 (I576113,I576065,I508898);
and I_33679 (I576130,I576113,I508916);
or I_33680 (I576147,I576130,I508910);
DFFARX1 I_33681 (I576147,I3563,I575723,I576173,);
nor I_33682 (I576181,I576173,I575797);
nor I_33683 (I575700,I575749,I576181);
not I_33684 (I576212,I576173);
nor I_33685 (I576229,I576212,I575907);
DFFARX1 I_33686 (I576229,I3563,I575723,I575706,);
nand I_33687 (I576260,I576212,I575839);
nor I_33688 (I575694,I576065,I576260);
not I_33689 (I576318,I3570);
DFFARX1 I_33690 (I1329231,I3563,I576318,I576344,);
DFFARX1 I_33691 (I576344,I3563,I576318,I576361,);
not I_33692 (I576310,I576361);
DFFARX1 I_33693 (I1329237,I3563,I576318,I576392,);
not I_33694 (I576400,I1329240);
nor I_33695 (I576417,I576344,I576400);
not I_33696 (I576434,I1329243);
not I_33697 (I576451,I1329228);
nand I_33698 (I576468,I576451,I1329243);
nor I_33699 (I576485,I576400,I576468);
nor I_33700 (I576502,I576392,I576485);
DFFARX1 I_33701 (I576451,I3563,I576318,I576307,);
nor I_33702 (I576533,I1329228,I1329234);
nand I_33703 (I576550,I576533,I1329216);
nor I_33704 (I576567,I576550,I576434);
nand I_33705 (I576292,I576567,I1329240);
DFFARX1 I_33706 (I576550,I3563,I576318,I576304,);
nand I_33707 (I576612,I576434,I1329228);
nor I_33708 (I576629,I576434,I1329228);
nand I_33709 (I576298,I576417,I576629);
not I_33710 (I576660,I1329216);
nor I_33711 (I576677,I576660,I576612);
DFFARX1 I_33712 (I576677,I3563,I576318,I576286,);
nor I_33713 (I576708,I576660,I1329225);
and I_33714 (I576725,I576708,I1329222);
or I_33715 (I576742,I576725,I1329219);
DFFARX1 I_33716 (I576742,I3563,I576318,I576768,);
nor I_33717 (I576776,I576768,I576392);
nor I_33718 (I576295,I576344,I576776);
not I_33719 (I576807,I576768);
nor I_33720 (I576824,I576807,I576502);
DFFARX1 I_33721 (I576824,I3563,I576318,I576301,);
nand I_33722 (I576855,I576807,I576434);
nor I_33723 (I576289,I576660,I576855);
not I_33724 (I576913,I3570);
DFFARX1 I_33725 (I834780,I3563,I576913,I576939,);
DFFARX1 I_33726 (I576939,I3563,I576913,I576956,);
not I_33727 (I576905,I576956);
DFFARX1 I_33728 (I834777,I3563,I576913,I576987,);
not I_33729 (I576995,I834777);
nor I_33730 (I577012,I576939,I576995);
not I_33731 (I577029,I834774);
not I_33732 (I577046,I834789);
nand I_33733 (I577063,I577046,I834774);
nor I_33734 (I577080,I576995,I577063);
nor I_33735 (I577097,I576987,I577080);
DFFARX1 I_33736 (I577046,I3563,I576913,I576902,);
nor I_33737 (I577128,I834789,I834783);
nand I_33738 (I577145,I577128,I834771);
nor I_33739 (I577162,I577145,I577029);
nand I_33740 (I576887,I577162,I834777);
DFFARX1 I_33741 (I577145,I3563,I576913,I576899,);
nand I_33742 (I577207,I577029,I834789);
nor I_33743 (I577224,I577029,I834789);
nand I_33744 (I576893,I577012,I577224);
not I_33745 (I577255,I834792);
nor I_33746 (I577272,I577255,I577207);
DFFARX1 I_33747 (I577272,I3563,I576913,I576881,);
nor I_33748 (I577303,I577255,I834771);
and I_33749 (I577320,I577303,I834786);
or I_33750 (I577337,I577320,I834774);
DFFARX1 I_33751 (I577337,I3563,I576913,I577363,);
nor I_33752 (I577371,I577363,I576987);
nor I_33753 (I576890,I576939,I577371);
not I_33754 (I577402,I577363);
nor I_33755 (I577419,I577402,I577097);
DFFARX1 I_33756 (I577419,I3563,I576913,I576896,);
nand I_33757 (I577450,I577402,I577029);
nor I_33758 (I576884,I577255,I577450);
not I_33759 (I577508,I3570);
DFFARX1 I_33760 (I1076392,I3563,I577508,I577534,);
DFFARX1 I_33761 (I577534,I3563,I577508,I577551,);
not I_33762 (I577500,I577551);
DFFARX1 I_33763 (I1076395,I3563,I577508,I577582,);
not I_33764 (I577590,I1076398);
nor I_33765 (I577607,I577534,I577590);
not I_33766 (I577624,I1076410);
not I_33767 (I577641,I1076401);
nand I_33768 (I577658,I577641,I1076410);
nor I_33769 (I577675,I577590,I577658);
nor I_33770 (I577692,I577582,I577675);
DFFARX1 I_33771 (I577641,I3563,I577508,I577497,);
nor I_33772 (I577723,I1076401,I1076407);
nand I_33773 (I577740,I577723,I1076395);
nor I_33774 (I577757,I577740,I577624);
nand I_33775 (I577482,I577757,I1076398);
DFFARX1 I_33776 (I577740,I3563,I577508,I577494,);
nand I_33777 (I577802,I577624,I1076401);
nor I_33778 (I577819,I577624,I1076401);
nand I_33779 (I577488,I577607,I577819);
not I_33780 (I577850,I1076398);
nor I_33781 (I577867,I577850,I577802);
DFFARX1 I_33782 (I577867,I3563,I577508,I577476,);
nor I_33783 (I577898,I577850,I1076404);
and I_33784 (I577915,I577898,I1076392);
or I_33785 (I577932,I577915,I1076413);
DFFARX1 I_33786 (I577932,I3563,I577508,I577958,);
nor I_33787 (I577966,I577958,I577582);
nor I_33788 (I577485,I577534,I577966);
not I_33789 (I577997,I577958);
nor I_33790 (I578014,I577997,I577692);
DFFARX1 I_33791 (I578014,I3563,I577508,I577491,);
nand I_33792 (I578045,I577997,I577624);
nor I_33793 (I577479,I577850,I578045);
not I_33794 (I578103,I3570);
DFFARX1 I_33795 (I230963,I3563,I578103,I578129,);
not I_33796 (I578137,I578129);
DFFARX1 I_33797 (I230948,I3563,I578103,I578163,);
not I_33798 (I578171,I230966);
nand I_33799 (I578188,I578171,I230951);
not I_33800 (I578205,I578188);
nor I_33801 (I578222,I578205,I230948);
nor I_33802 (I578239,I578137,I578222);
DFFARX1 I_33803 (I578239,I3563,I578103,I578089,);
not I_33804 (I578270,I230948);
nand I_33805 (I578287,I578270,I578205);
and I_33806 (I578304,I578270,I230951);
nand I_33807 (I578321,I578304,I230972);
nor I_33808 (I578086,I578321,I578270);
and I_33809 (I578077,I578163,I578321);
not I_33810 (I578366,I578321);
nand I_33811 (I578080,I578163,I578366);
nor I_33812 (I578074,I578129,I578321);
not I_33813 (I578411,I230960);
nor I_33814 (I578428,I578411,I230951);
nand I_33815 (I578445,I578428,I578270);
nor I_33816 (I578083,I578188,I578445);
nor I_33817 (I578476,I578411,I230954);
and I_33818 (I578493,I578476,I230969);
or I_33819 (I578510,I578493,I230957);
DFFARX1 I_33820 (I578510,I3563,I578103,I578536,);
nor I_33821 (I578544,I578536,I578287);
DFFARX1 I_33822 (I578544,I3563,I578103,I578071,);
DFFARX1 I_33823 (I578536,I3563,I578103,I578095,);
not I_33824 (I578589,I578536);
nor I_33825 (I578606,I578589,I578163);
nor I_33826 (I578623,I578428,I578606);
DFFARX1 I_33827 (I578623,I3563,I578103,I578092,);
not I_33828 (I578681,I3570);
DFFARX1 I_33829 (I372853,I3563,I578681,I578707,);
not I_33830 (I578715,I578707);
DFFARX1 I_33831 (I372868,I3563,I578681,I578741,);
not I_33832 (I578749,I372871);
nand I_33833 (I578766,I578749,I372850);
not I_33834 (I578783,I578766);
nor I_33835 (I578800,I578783,I372874);
nor I_33836 (I578817,I578715,I578800);
DFFARX1 I_33837 (I578817,I3563,I578681,I578667,);
not I_33838 (I578848,I372874);
nand I_33839 (I578865,I578848,I578783);
and I_33840 (I578882,I578848,I372856);
nand I_33841 (I578899,I578882,I372847);
nor I_33842 (I578664,I578899,I578848);
and I_33843 (I578655,I578741,I578899);
not I_33844 (I578944,I578899);
nand I_33845 (I578658,I578741,I578944);
nor I_33846 (I578652,I578707,I578899);
not I_33847 (I578989,I372847);
nor I_33848 (I579006,I578989,I372856);
nand I_33849 (I579023,I579006,I578848);
nor I_33850 (I578661,I578766,I579023);
nor I_33851 (I579054,I578989,I372862);
and I_33852 (I579071,I579054,I372865);
or I_33853 (I579088,I579071,I372859);
DFFARX1 I_33854 (I579088,I3563,I578681,I579114,);
nor I_33855 (I579122,I579114,I578865);
DFFARX1 I_33856 (I579122,I3563,I578681,I578649,);
DFFARX1 I_33857 (I579114,I3563,I578681,I578673,);
not I_33858 (I579167,I579114);
nor I_33859 (I579184,I579167,I578741);
nor I_33860 (I579201,I579006,I579184);
DFFARX1 I_33861 (I579201,I3563,I578681,I578670,);
not I_33862 (I579259,I3570);
DFFARX1 I_33863 (I915527,I3563,I579259,I579285,);
not I_33864 (I579293,I579285);
DFFARX1 I_33865 (I915524,I3563,I579259,I579319,);
not I_33866 (I579327,I915521);
nand I_33867 (I579344,I579327,I915548);
not I_33868 (I579361,I579344);
nor I_33869 (I579378,I579361,I915536);
nor I_33870 (I579395,I579293,I579378);
DFFARX1 I_33871 (I579395,I3563,I579259,I579245,);
not I_33872 (I579426,I915536);
nand I_33873 (I579443,I579426,I579361);
and I_33874 (I579460,I579426,I915542);
nand I_33875 (I579477,I579460,I915533);
nor I_33876 (I579242,I579477,I579426);
and I_33877 (I579233,I579319,I579477);
not I_33878 (I579522,I579477);
nand I_33879 (I579236,I579319,I579522);
nor I_33880 (I579230,I579285,I579477);
not I_33881 (I579567,I915530);
nor I_33882 (I579584,I579567,I915542);
nand I_33883 (I579601,I579584,I579426);
nor I_33884 (I579239,I579344,I579601);
nor I_33885 (I579632,I579567,I915545);
and I_33886 (I579649,I579632,I915539);
or I_33887 (I579666,I579649,I915521);
DFFARX1 I_33888 (I579666,I3563,I579259,I579692,);
nor I_33889 (I579700,I579692,I579443);
DFFARX1 I_33890 (I579700,I3563,I579259,I579227,);
DFFARX1 I_33891 (I579692,I3563,I579259,I579251,);
not I_33892 (I579745,I579692);
nor I_33893 (I579762,I579745,I579319);
nor I_33894 (I579779,I579584,I579762);
DFFARX1 I_33895 (I579779,I3563,I579259,I579248,);
not I_33896 (I579837,I3570);
DFFARX1 I_33897 (I1315509,I3563,I579837,I579863,);
not I_33898 (I579871,I579863);
DFFARX1 I_33899 (I1315521,I3563,I579837,I579897,);
not I_33900 (I579905,I1315512);
nand I_33901 (I579922,I579905,I1315500);
not I_33902 (I579939,I579922);
nor I_33903 (I579956,I579939,I1315497);
nor I_33904 (I579973,I579871,I579956);
DFFARX1 I_33905 (I579973,I3563,I579837,I579823,);
not I_33906 (I580004,I1315497);
nand I_33907 (I580021,I580004,I579939);
and I_33908 (I580038,I580004,I1315503);
nand I_33909 (I580055,I580038,I1315500);
nor I_33910 (I579820,I580055,I580004);
and I_33911 (I579811,I579897,I580055);
not I_33912 (I580100,I580055);
nand I_33913 (I579814,I579897,I580100);
nor I_33914 (I579808,I579863,I580055);
not I_33915 (I580145,I1315518);
nor I_33916 (I580162,I580145,I1315503);
nand I_33917 (I580179,I580162,I580004);
nor I_33918 (I579817,I579922,I580179);
nor I_33919 (I580210,I580145,I1315506);
and I_33920 (I580227,I580210,I1315497);
or I_33921 (I580244,I580227,I1315515);
DFFARX1 I_33922 (I580244,I3563,I579837,I580270,);
nor I_33923 (I580278,I580270,I580021);
DFFARX1 I_33924 (I580278,I3563,I579837,I579805,);
DFFARX1 I_33925 (I580270,I3563,I579837,I579829,);
not I_33926 (I580323,I580270);
nor I_33927 (I580340,I580323,I579897);
nor I_33928 (I580357,I580162,I580340);
DFFARX1 I_33929 (I580357,I3563,I579837,I579826,);
not I_33930 (I580415,I3570);
DFFARX1 I_33931 (I1298747,I3563,I580415,I580441,);
not I_33932 (I580449,I580441);
DFFARX1 I_33933 (I1298759,I3563,I580415,I580475,);
not I_33934 (I580483,I1298750);
nand I_33935 (I580500,I580483,I1298738);
not I_33936 (I580517,I580500);
nor I_33937 (I580534,I580517,I1298735);
nor I_33938 (I580551,I580449,I580534);
DFFARX1 I_33939 (I580551,I3563,I580415,I580401,);
not I_33940 (I580582,I1298735);
nand I_33941 (I580599,I580582,I580517);
and I_33942 (I580616,I580582,I1298741);
nand I_33943 (I580633,I580616,I1298738);
nor I_33944 (I580398,I580633,I580582);
and I_33945 (I580389,I580475,I580633);
not I_33946 (I580678,I580633);
nand I_33947 (I580392,I580475,I580678);
nor I_33948 (I580386,I580441,I580633);
not I_33949 (I580723,I1298756);
nor I_33950 (I580740,I580723,I1298741);
nand I_33951 (I580757,I580740,I580582);
nor I_33952 (I580395,I580500,I580757);
nor I_33953 (I580788,I580723,I1298744);
and I_33954 (I580805,I580788,I1298735);
or I_33955 (I580822,I580805,I1298753);
DFFARX1 I_33956 (I580822,I3563,I580415,I580848,);
nor I_33957 (I580856,I580848,I580599);
DFFARX1 I_33958 (I580856,I3563,I580415,I580383,);
DFFARX1 I_33959 (I580848,I3563,I580415,I580407,);
not I_33960 (I580901,I580848);
nor I_33961 (I580918,I580901,I580475);
nor I_33962 (I580935,I580740,I580918);
DFFARX1 I_33963 (I580935,I3563,I580415,I580404,);
not I_33964 (I580993,I3570);
DFFARX1 I_33965 (I726617,I3563,I580993,I581019,);
not I_33966 (I581027,I581019);
DFFARX1 I_33967 (I726629,I3563,I580993,I581053,);
not I_33968 (I581061,I726620);
nand I_33969 (I581078,I581061,I726623);
not I_33970 (I581095,I581078);
nor I_33971 (I581112,I581095,I726626);
nor I_33972 (I581129,I581027,I581112);
DFFARX1 I_33973 (I581129,I3563,I580993,I580979,);
not I_33974 (I581160,I726626);
nand I_33975 (I581177,I581160,I581095);
and I_33976 (I581194,I581160,I726620);
nand I_33977 (I581211,I581194,I726632);
nor I_33978 (I580976,I581211,I581160);
and I_33979 (I580967,I581053,I581211);
not I_33980 (I581256,I581211);
nand I_33981 (I580970,I581053,I581256);
nor I_33982 (I580964,I581019,I581211);
not I_33983 (I581301,I726638);
nor I_33984 (I581318,I581301,I726620);
nand I_33985 (I581335,I581318,I581160);
nor I_33986 (I580973,I581078,I581335);
nor I_33987 (I581366,I581301,I726617);
and I_33988 (I581383,I581366,I726635);
or I_33989 (I581400,I581383,I726641);
DFFARX1 I_33990 (I581400,I3563,I580993,I581426,);
nor I_33991 (I581434,I581426,I581177);
DFFARX1 I_33992 (I581434,I3563,I580993,I580961,);
DFFARX1 I_33993 (I581426,I3563,I580993,I580985,);
not I_33994 (I581479,I581426);
nor I_33995 (I581496,I581479,I581053);
nor I_33996 (I581513,I581318,I581496);
DFFARX1 I_33997 (I581513,I3563,I580993,I580982,);
not I_33998 (I581571,I3570);
DFFARX1 I_33999 (I1235495,I3563,I581571,I581597,);
not I_34000 (I581605,I581597);
DFFARX1 I_34001 (I1235501,I3563,I581571,I581631,);
not I_34002 (I581639,I1235495);
nand I_34003 (I581656,I581639,I1235498);
not I_34004 (I581673,I581656);
nor I_34005 (I581690,I581673,I1235516);
nor I_34006 (I581707,I581605,I581690);
DFFARX1 I_34007 (I581707,I3563,I581571,I581557,);
not I_34008 (I581738,I1235516);
nand I_34009 (I581755,I581738,I581673);
and I_34010 (I581772,I581738,I1235519);
nand I_34011 (I581789,I581772,I1235498);
nor I_34012 (I581554,I581789,I581738);
and I_34013 (I581545,I581631,I581789);
not I_34014 (I581834,I581789);
nand I_34015 (I581548,I581631,I581834);
nor I_34016 (I581542,I581597,I581789);
not I_34017 (I581879,I1235504);
nor I_34018 (I581896,I581879,I1235519);
nand I_34019 (I581913,I581896,I581738);
nor I_34020 (I581551,I581656,I581913);
nor I_34021 (I581944,I581879,I1235510);
and I_34022 (I581961,I581944,I1235507);
or I_34023 (I581978,I581961,I1235513);
DFFARX1 I_34024 (I581978,I3563,I581571,I582004,);
nor I_34025 (I582012,I582004,I581755);
DFFARX1 I_34026 (I582012,I3563,I581571,I581539,);
DFFARX1 I_34027 (I582004,I3563,I581571,I581563,);
not I_34028 (I582057,I582004);
nor I_34029 (I582074,I582057,I581631);
nor I_34030 (I582091,I581896,I582074);
DFFARX1 I_34031 (I582091,I3563,I581571,I581560,);
not I_34032 (I582149,I3570);
DFFARX1 I_34033 (I139410,I3563,I582149,I582175,);
not I_34034 (I582183,I582175);
DFFARX1 I_34035 (I139389,I3563,I582149,I582209,);
not I_34036 (I582217,I139386);
nand I_34037 (I582234,I582217,I139401);
not I_34038 (I582251,I582234);
nor I_34039 (I582268,I582251,I139389);
nor I_34040 (I582285,I582183,I582268);
DFFARX1 I_34041 (I582285,I3563,I582149,I582135,);
not I_34042 (I582316,I139389);
nand I_34043 (I582333,I582316,I582251);
and I_34044 (I582350,I582316,I139392);
nand I_34045 (I582367,I582350,I139407);
nor I_34046 (I582132,I582367,I582316);
and I_34047 (I582123,I582209,I582367);
not I_34048 (I582412,I582367);
nand I_34049 (I582126,I582209,I582412);
nor I_34050 (I582120,I582175,I582367);
not I_34051 (I582457,I139398);
nor I_34052 (I582474,I582457,I139392);
nand I_34053 (I582491,I582474,I582316);
nor I_34054 (I582129,I582234,I582491);
nor I_34055 (I582522,I582457,I139386);
and I_34056 (I582539,I582522,I139395);
or I_34057 (I582556,I582539,I139404);
DFFARX1 I_34058 (I582556,I3563,I582149,I582582,);
nor I_34059 (I582590,I582582,I582333);
DFFARX1 I_34060 (I582590,I3563,I582149,I582117,);
DFFARX1 I_34061 (I582582,I3563,I582149,I582141,);
not I_34062 (I582635,I582582);
nor I_34063 (I582652,I582635,I582209);
nor I_34064 (I582669,I582474,I582652);
DFFARX1 I_34065 (I582669,I3563,I582149,I582138,);
not I_34066 (I582727,I3570);
DFFARX1 I_34067 (I443630,I3563,I582727,I582753,);
not I_34068 (I582761,I582753);
DFFARX1 I_34069 (I443642,I3563,I582727,I582787,);
not I_34070 (I582795,I443618);
nand I_34071 (I582812,I582795,I443645);
not I_34072 (I582829,I582812);
nor I_34073 (I582846,I582829,I443633);
nor I_34074 (I582863,I582761,I582846);
DFFARX1 I_34075 (I582863,I3563,I582727,I582713,);
not I_34076 (I582894,I443633);
nand I_34077 (I582911,I582894,I582829);
and I_34078 (I582928,I582894,I443618);
nand I_34079 (I582945,I582928,I443621);
nor I_34080 (I582710,I582945,I582894);
and I_34081 (I582701,I582787,I582945);
not I_34082 (I582990,I582945);
nand I_34083 (I582704,I582787,I582990);
nor I_34084 (I582698,I582753,I582945);
not I_34085 (I583035,I443627);
nor I_34086 (I583052,I583035,I443618);
nand I_34087 (I583069,I583052,I582894);
nor I_34088 (I582707,I582812,I583069);
nor I_34089 (I583100,I583035,I443636);
and I_34090 (I583117,I583100,I443624);
or I_34091 (I583134,I583117,I443639);
DFFARX1 I_34092 (I583134,I3563,I582727,I583160,);
nor I_34093 (I583168,I583160,I582911);
DFFARX1 I_34094 (I583168,I3563,I582727,I582695,);
DFFARX1 I_34095 (I583160,I3563,I582727,I582719,);
not I_34096 (I583213,I583160);
nor I_34097 (I583230,I583213,I582787);
nor I_34098 (I583247,I583052,I583230);
DFFARX1 I_34099 (I583247,I3563,I582727,I582716,);
not I_34100 (I583305,I3570);
DFFARX1 I_34101 (I1064071,I3563,I583305,I583331,);
not I_34102 (I583339,I583331);
DFFARX1 I_34103 (I1064062,I3563,I583305,I583365,);
not I_34104 (I583373,I1064056);
nand I_34105 (I583390,I583373,I1064068);
not I_34106 (I583407,I583390);
nor I_34107 (I583424,I583407,I1064059);
nor I_34108 (I583441,I583339,I583424);
DFFARX1 I_34109 (I583441,I3563,I583305,I583291,);
not I_34110 (I583472,I1064059);
nand I_34111 (I583489,I583472,I583407);
and I_34112 (I583506,I583472,I1064065);
nand I_34113 (I583523,I583506,I1064050);
nor I_34114 (I583288,I583523,I583472);
and I_34115 (I583279,I583365,I583523);
not I_34116 (I583568,I583523);
nand I_34117 (I583282,I583365,I583568);
nor I_34118 (I583276,I583331,I583523);
not I_34119 (I583613,I1064050);
nor I_34120 (I583630,I583613,I1064065);
nand I_34121 (I583647,I583630,I583472);
nor I_34122 (I583285,I583390,I583647);
nor I_34123 (I583678,I583613,I1064053);
and I_34124 (I583695,I583678,I1064056);
or I_34125 (I583712,I583695,I1064053);
DFFARX1 I_34126 (I583712,I3563,I583305,I583738,);
nor I_34127 (I583746,I583738,I583489);
DFFARX1 I_34128 (I583746,I3563,I583305,I583273,);
DFFARX1 I_34129 (I583738,I3563,I583305,I583297,);
not I_34130 (I583791,I583738);
nor I_34131 (I583808,I583791,I583365);
nor I_34132 (I583825,I583630,I583808);
DFFARX1 I_34133 (I583825,I3563,I583305,I583294,);
not I_34134 (I583883,I3570);
DFFARX1 I_34135 (I222038,I3563,I583883,I583909,);
not I_34136 (I583917,I583909);
DFFARX1 I_34137 (I222023,I3563,I583883,I583943,);
not I_34138 (I583951,I222041);
nand I_34139 (I583968,I583951,I222026);
not I_34140 (I583985,I583968);
nor I_34141 (I584002,I583985,I222023);
nor I_34142 (I584019,I583917,I584002);
DFFARX1 I_34143 (I584019,I3563,I583883,I583869,);
not I_34144 (I584050,I222023);
nand I_34145 (I584067,I584050,I583985);
and I_34146 (I584084,I584050,I222026);
nand I_34147 (I584101,I584084,I222047);
nor I_34148 (I583866,I584101,I584050);
and I_34149 (I583857,I583943,I584101);
not I_34150 (I584146,I584101);
nand I_34151 (I583860,I583943,I584146);
nor I_34152 (I583854,I583909,I584101);
not I_34153 (I584191,I222035);
nor I_34154 (I584208,I584191,I222026);
nand I_34155 (I584225,I584208,I584050);
nor I_34156 (I583863,I583968,I584225);
nor I_34157 (I584256,I584191,I222029);
and I_34158 (I584273,I584256,I222044);
or I_34159 (I584290,I584273,I222032);
DFFARX1 I_34160 (I584290,I3563,I583883,I584316,);
nor I_34161 (I584324,I584316,I584067);
DFFARX1 I_34162 (I584324,I3563,I583883,I583851,);
DFFARX1 I_34163 (I584316,I3563,I583883,I583875,);
not I_34164 (I584369,I584316);
nor I_34165 (I584386,I584369,I583943);
nor I_34166 (I584403,I584208,I584386);
DFFARX1 I_34167 (I584403,I3563,I583883,I583872,);
not I_34168 (I584461,I3570);
DFFARX1 I_34169 (I428942,I3563,I584461,I584487,);
not I_34170 (I584495,I584487);
DFFARX1 I_34171 (I428954,I3563,I584461,I584521,);
not I_34172 (I584529,I428930);
nand I_34173 (I584546,I584529,I428957);
not I_34174 (I584563,I584546);
nor I_34175 (I584580,I584563,I428945);
nor I_34176 (I584597,I584495,I584580);
DFFARX1 I_34177 (I584597,I3563,I584461,I584447,);
not I_34178 (I584628,I428945);
nand I_34179 (I584645,I584628,I584563);
and I_34180 (I584662,I584628,I428930);
nand I_34181 (I584679,I584662,I428933);
nor I_34182 (I584444,I584679,I584628);
and I_34183 (I584435,I584521,I584679);
not I_34184 (I584724,I584679);
nand I_34185 (I584438,I584521,I584724);
nor I_34186 (I584432,I584487,I584679);
not I_34187 (I584769,I428939);
nor I_34188 (I584786,I584769,I428930);
nand I_34189 (I584803,I584786,I584628);
nor I_34190 (I584441,I584546,I584803);
nor I_34191 (I584834,I584769,I428948);
and I_34192 (I584851,I584834,I428936);
or I_34193 (I584868,I584851,I428951);
DFFARX1 I_34194 (I584868,I3563,I584461,I584894,);
nor I_34195 (I584902,I584894,I584645);
DFFARX1 I_34196 (I584902,I3563,I584461,I584429,);
DFFARX1 I_34197 (I584894,I3563,I584461,I584453,);
not I_34198 (I584947,I584894);
nor I_34199 (I584964,I584947,I584521);
nor I_34200 (I584981,I584786,I584964);
DFFARX1 I_34201 (I584981,I3563,I584461,I584450,);
not I_34202 (I585039,I3570);
DFFARX1 I_34203 (I518702,I3563,I585039,I585065,);
not I_34204 (I585073,I585065);
DFFARX1 I_34205 (I518714,I3563,I585039,I585099,);
not I_34206 (I585107,I518690);
nand I_34207 (I585124,I585107,I518717);
not I_34208 (I585141,I585124);
nor I_34209 (I585158,I585141,I518705);
nor I_34210 (I585175,I585073,I585158);
DFFARX1 I_34211 (I585175,I3563,I585039,I585025,);
not I_34212 (I585206,I518705);
nand I_34213 (I585223,I585206,I585141);
and I_34214 (I585240,I585206,I518690);
nand I_34215 (I585257,I585240,I518693);
nor I_34216 (I585022,I585257,I585206);
and I_34217 (I585013,I585099,I585257);
not I_34218 (I585302,I585257);
nand I_34219 (I585016,I585099,I585302);
nor I_34220 (I585010,I585065,I585257);
not I_34221 (I585347,I518699);
nor I_34222 (I585364,I585347,I518690);
nand I_34223 (I585381,I585364,I585206);
nor I_34224 (I585019,I585124,I585381);
nor I_34225 (I585412,I585347,I518708);
and I_34226 (I585429,I585412,I518696);
or I_34227 (I585446,I585429,I518711);
DFFARX1 I_34228 (I585446,I3563,I585039,I585472,);
nor I_34229 (I585480,I585472,I585223);
DFFARX1 I_34230 (I585480,I3563,I585039,I585007,);
DFFARX1 I_34231 (I585472,I3563,I585039,I585031,);
not I_34232 (I585525,I585472);
nor I_34233 (I585542,I585525,I585099);
nor I_34234 (I585559,I585364,I585542);
DFFARX1 I_34235 (I585559,I3563,I585039,I585028,);
not I_34236 (I585617,I3570);
DFFARX1 I_34237 (I743379,I3563,I585617,I585643,);
not I_34238 (I585651,I585643);
DFFARX1 I_34239 (I743391,I3563,I585617,I585677,);
not I_34240 (I585685,I743382);
nand I_34241 (I585702,I585685,I743385);
not I_34242 (I585719,I585702);
nor I_34243 (I585736,I585719,I743388);
nor I_34244 (I585753,I585651,I585736);
DFFARX1 I_34245 (I585753,I3563,I585617,I585603,);
not I_34246 (I585784,I743388);
nand I_34247 (I585801,I585784,I585719);
and I_34248 (I585818,I585784,I743382);
nand I_34249 (I585835,I585818,I743394);
nor I_34250 (I585600,I585835,I585784);
and I_34251 (I585591,I585677,I585835);
not I_34252 (I585880,I585835);
nand I_34253 (I585594,I585677,I585880);
nor I_34254 (I585588,I585643,I585835);
not I_34255 (I585925,I743400);
nor I_34256 (I585942,I585925,I743382);
nand I_34257 (I585959,I585942,I585784);
nor I_34258 (I585597,I585702,I585959);
nor I_34259 (I585990,I585925,I743379);
and I_34260 (I586007,I585990,I743397);
or I_34261 (I586024,I586007,I743403);
DFFARX1 I_34262 (I586024,I3563,I585617,I586050,);
nor I_34263 (I586058,I586050,I585801);
DFFARX1 I_34264 (I586058,I3563,I585617,I585585,);
DFFARX1 I_34265 (I586050,I3563,I585617,I585609,);
not I_34266 (I586103,I586050);
nor I_34267 (I586120,I586103,I585677);
nor I_34268 (I586137,I585942,I586120);
DFFARX1 I_34269 (I586137,I3563,I585617,I585606,);
not I_34270 (I586195,I3570);
DFFARX1 I_34271 (I189908,I3563,I586195,I586221,);
not I_34272 (I586229,I586221);
DFFARX1 I_34273 (I189893,I3563,I586195,I586255,);
not I_34274 (I586263,I189911);
nand I_34275 (I586280,I586263,I189896);
not I_34276 (I586297,I586280);
nor I_34277 (I586314,I586297,I189893);
nor I_34278 (I586331,I586229,I586314);
DFFARX1 I_34279 (I586331,I3563,I586195,I586181,);
not I_34280 (I586362,I189893);
nand I_34281 (I586379,I586362,I586297);
and I_34282 (I586396,I586362,I189896);
nand I_34283 (I586413,I586396,I189917);
nor I_34284 (I586178,I586413,I586362);
and I_34285 (I586169,I586255,I586413);
not I_34286 (I586458,I586413);
nand I_34287 (I586172,I586255,I586458);
nor I_34288 (I586166,I586221,I586413);
not I_34289 (I586503,I189905);
nor I_34290 (I586520,I586503,I189896);
nand I_34291 (I586537,I586520,I586362);
nor I_34292 (I586175,I586280,I586537);
nor I_34293 (I586568,I586503,I189899);
and I_34294 (I586585,I586568,I189914);
or I_34295 (I586602,I586585,I189902);
DFFARX1 I_34296 (I586602,I3563,I586195,I586628,);
nor I_34297 (I586636,I586628,I586379);
DFFARX1 I_34298 (I586636,I3563,I586195,I586163,);
DFFARX1 I_34299 (I586628,I3563,I586195,I586187,);
not I_34300 (I586681,I586628);
nor I_34301 (I586698,I586681,I586255);
nor I_34302 (I586715,I586520,I586698);
DFFARX1 I_34303 (I586715,I3563,I586195,I586184,);
not I_34304 (I586773,I3570);
DFFARX1 I_34305 (I78805,I3563,I586773,I586799,);
not I_34306 (I586807,I586799);
DFFARX1 I_34307 (I78784,I3563,I586773,I586833,);
not I_34308 (I586841,I78781);
nand I_34309 (I586858,I586841,I78796);
not I_34310 (I586875,I586858);
nor I_34311 (I586892,I586875,I78784);
nor I_34312 (I586909,I586807,I586892);
DFFARX1 I_34313 (I586909,I3563,I586773,I586759,);
not I_34314 (I586940,I78784);
nand I_34315 (I586957,I586940,I586875);
and I_34316 (I586974,I586940,I78787);
nand I_34317 (I586991,I586974,I78802);
nor I_34318 (I586756,I586991,I586940);
and I_34319 (I586747,I586833,I586991);
not I_34320 (I587036,I586991);
nand I_34321 (I586750,I586833,I587036);
nor I_34322 (I586744,I586799,I586991);
not I_34323 (I587081,I78793);
nor I_34324 (I587098,I587081,I78787);
nand I_34325 (I587115,I587098,I586940);
nor I_34326 (I586753,I586858,I587115);
nor I_34327 (I587146,I587081,I78781);
and I_34328 (I587163,I587146,I78790);
or I_34329 (I587180,I587163,I78799);
DFFARX1 I_34330 (I587180,I3563,I586773,I587206,);
nor I_34331 (I587214,I587206,I586957);
DFFARX1 I_34332 (I587214,I3563,I586773,I586741,);
DFFARX1 I_34333 (I587206,I3563,I586773,I586765,);
not I_34334 (I587259,I587206);
nor I_34335 (I587276,I587259,I586833);
nor I_34336 (I587293,I587098,I587276);
DFFARX1 I_34337 (I587293,I3563,I586773,I586762,);
not I_34338 (I587351,I3570);
DFFARX1 I_34339 (I27138,I3563,I587351,I587377,);
not I_34340 (I587385,I587377);
DFFARX1 I_34341 (I27141,I3563,I587351,I587411,);
not I_34342 (I587419,I27135);
nand I_34343 (I587436,I587419,I27159);
not I_34344 (I587453,I587436);
nor I_34345 (I587470,I587453,I27138);
nor I_34346 (I587487,I587385,I587470);
DFFARX1 I_34347 (I587487,I3563,I587351,I587337,);
not I_34348 (I587518,I27138);
nand I_34349 (I587535,I587518,I587453);
and I_34350 (I587552,I587518,I27153);
nand I_34351 (I587569,I587552,I27147);
nor I_34352 (I587334,I587569,I587518);
and I_34353 (I587325,I587411,I587569);
not I_34354 (I587614,I587569);
nand I_34355 (I587328,I587411,I587614);
nor I_34356 (I587322,I587377,I587569);
not I_34357 (I587659,I27156);
nor I_34358 (I587676,I587659,I27153);
nand I_34359 (I587693,I587676,I587518);
nor I_34360 (I587331,I587436,I587693);
nor I_34361 (I587724,I587659,I27135);
and I_34362 (I587741,I587724,I27144);
or I_34363 (I587758,I587741,I27150);
DFFARX1 I_34364 (I587758,I3563,I587351,I587784,);
nor I_34365 (I587792,I587784,I587535);
DFFARX1 I_34366 (I587792,I3563,I587351,I587319,);
DFFARX1 I_34367 (I587784,I3563,I587351,I587343,);
not I_34368 (I587837,I587784);
nor I_34369 (I587854,I587837,I587411);
nor I_34370 (I587871,I587676,I587854);
DFFARX1 I_34371 (I587871,I3563,I587351,I587340,);
not I_34372 (I587929,I3570);
DFFARX1 I_34373 (I464846,I3563,I587929,I587955,);
not I_34374 (I587963,I587955);
DFFARX1 I_34375 (I464858,I3563,I587929,I587989,);
not I_34376 (I587997,I464834);
nand I_34377 (I588014,I587997,I464861);
not I_34378 (I588031,I588014);
nor I_34379 (I588048,I588031,I464849);
nor I_34380 (I588065,I587963,I588048);
DFFARX1 I_34381 (I588065,I3563,I587929,I587915,);
not I_34382 (I588096,I464849);
nand I_34383 (I588113,I588096,I588031);
and I_34384 (I588130,I588096,I464834);
nand I_34385 (I588147,I588130,I464837);
nor I_34386 (I587912,I588147,I588096);
and I_34387 (I587903,I587989,I588147);
not I_34388 (I588192,I588147);
nand I_34389 (I587906,I587989,I588192);
nor I_34390 (I587900,I587955,I588147);
not I_34391 (I588237,I464843);
nor I_34392 (I588254,I588237,I464834);
nand I_34393 (I588271,I588254,I588096);
nor I_34394 (I587909,I588014,I588271);
nor I_34395 (I588302,I588237,I464852);
and I_34396 (I588319,I588302,I464840);
or I_34397 (I588336,I588319,I464855);
DFFARX1 I_34398 (I588336,I3563,I587929,I588362,);
nor I_34399 (I588370,I588362,I588113);
DFFARX1 I_34400 (I588370,I3563,I587929,I587897,);
DFFARX1 I_34401 (I588362,I3563,I587929,I587921,);
not I_34402 (I588415,I588362);
nor I_34403 (I588432,I588415,I587989);
nor I_34404 (I588449,I588254,I588432);
DFFARX1 I_34405 (I588449,I3563,I587929,I587918,);
not I_34406 (I588507,I3570);
DFFARX1 I_34407 (I520334,I3563,I588507,I588533,);
not I_34408 (I588541,I588533);
DFFARX1 I_34409 (I520346,I3563,I588507,I588567,);
not I_34410 (I588575,I520322);
nand I_34411 (I588592,I588575,I520349);
not I_34412 (I588609,I588592);
nor I_34413 (I588626,I588609,I520337);
nor I_34414 (I588643,I588541,I588626);
DFFARX1 I_34415 (I588643,I3563,I588507,I588493,);
not I_34416 (I588674,I520337);
nand I_34417 (I588691,I588674,I588609);
and I_34418 (I588708,I588674,I520322);
nand I_34419 (I588725,I588708,I520325);
nor I_34420 (I588490,I588725,I588674);
and I_34421 (I588481,I588567,I588725);
not I_34422 (I588770,I588725);
nand I_34423 (I588484,I588567,I588770);
nor I_34424 (I588478,I588533,I588725);
not I_34425 (I588815,I520331);
nor I_34426 (I588832,I588815,I520322);
nand I_34427 (I588849,I588832,I588674);
nor I_34428 (I588487,I588592,I588849);
nor I_34429 (I588880,I588815,I520340);
and I_34430 (I588897,I588880,I520328);
or I_34431 (I588914,I588897,I520343);
DFFARX1 I_34432 (I588914,I3563,I588507,I588940,);
nor I_34433 (I588948,I588940,I588691);
DFFARX1 I_34434 (I588948,I3563,I588507,I588475,);
DFFARX1 I_34435 (I588940,I3563,I588507,I588499,);
not I_34436 (I588993,I588940);
nor I_34437 (I589010,I588993,I588567);
nor I_34438 (I589027,I588832,I589010);
DFFARX1 I_34439 (I589027,I3563,I588507,I588496,);
not I_34440 (I589085,I3570);
DFFARX1 I_34441 (I664771,I3563,I589085,I589111,);
not I_34442 (I589119,I589111);
DFFARX1 I_34443 (I664783,I3563,I589085,I589145,);
not I_34444 (I589153,I664774);
nand I_34445 (I589170,I589153,I664777);
not I_34446 (I589187,I589170);
nor I_34447 (I589204,I589187,I664780);
nor I_34448 (I589221,I589119,I589204);
DFFARX1 I_34449 (I589221,I3563,I589085,I589071,);
not I_34450 (I589252,I664780);
nand I_34451 (I589269,I589252,I589187);
and I_34452 (I589286,I589252,I664774);
nand I_34453 (I589303,I589286,I664786);
nor I_34454 (I589068,I589303,I589252);
and I_34455 (I589059,I589145,I589303);
not I_34456 (I589348,I589303);
nand I_34457 (I589062,I589145,I589348);
nor I_34458 (I589056,I589111,I589303);
not I_34459 (I589393,I664792);
nor I_34460 (I589410,I589393,I664774);
nand I_34461 (I589427,I589410,I589252);
nor I_34462 (I589065,I589170,I589427);
nor I_34463 (I589458,I589393,I664771);
and I_34464 (I589475,I589458,I664789);
or I_34465 (I589492,I589475,I664795);
DFFARX1 I_34466 (I589492,I3563,I589085,I589518,);
nor I_34467 (I589526,I589518,I589269);
DFFARX1 I_34468 (I589526,I3563,I589085,I589053,);
DFFARX1 I_34469 (I589518,I3563,I589085,I589077,);
not I_34470 (I589571,I589518);
nor I_34471 (I589588,I589571,I589145);
nor I_34472 (I589605,I589410,I589588);
DFFARX1 I_34473 (I589605,I3563,I589085,I589074,);
not I_34474 (I589663,I3570);
DFFARX1 I_34475 (I428398,I3563,I589663,I589689,);
not I_34476 (I589697,I589689);
DFFARX1 I_34477 (I428410,I3563,I589663,I589723,);
not I_34478 (I589731,I428386);
nand I_34479 (I589748,I589731,I428413);
not I_34480 (I589765,I589748);
nor I_34481 (I589782,I589765,I428401);
nor I_34482 (I589799,I589697,I589782);
DFFARX1 I_34483 (I589799,I3563,I589663,I589649,);
not I_34484 (I589830,I428401);
nand I_34485 (I589847,I589830,I589765);
and I_34486 (I589864,I589830,I428386);
nand I_34487 (I589881,I589864,I428389);
nor I_34488 (I589646,I589881,I589830);
and I_34489 (I589637,I589723,I589881);
not I_34490 (I589926,I589881);
nand I_34491 (I589640,I589723,I589926);
nor I_34492 (I589634,I589689,I589881);
not I_34493 (I589971,I428395);
nor I_34494 (I589988,I589971,I428386);
nand I_34495 (I590005,I589988,I589830);
nor I_34496 (I589643,I589748,I590005);
nor I_34497 (I590036,I589971,I428404);
and I_34498 (I590053,I590036,I428392);
or I_34499 (I590070,I590053,I428407);
DFFARX1 I_34500 (I590070,I3563,I589663,I590096,);
nor I_34501 (I590104,I590096,I589847);
DFFARX1 I_34502 (I590104,I3563,I589663,I589631,);
DFFARX1 I_34503 (I590096,I3563,I589663,I589655,);
not I_34504 (I590149,I590096);
nor I_34505 (I590166,I590149,I589723);
nor I_34506 (I590183,I589988,I590166);
DFFARX1 I_34507 (I590183,I3563,I589663,I589652,);
not I_34508 (I590241,I3570);
DFFARX1 I_34509 (I1106023,I3563,I590241,I590267,);
not I_34510 (I590275,I590267);
DFFARX1 I_34511 (I1106029,I3563,I590241,I590301,);
not I_34512 (I590309,I1106023);
nand I_34513 (I590326,I590309,I1106026);
not I_34514 (I590343,I590326);
nor I_34515 (I590360,I590343,I1106044);
nor I_34516 (I590377,I590275,I590360);
DFFARX1 I_34517 (I590377,I3563,I590241,I590227,);
not I_34518 (I590408,I1106044);
nand I_34519 (I590425,I590408,I590343);
and I_34520 (I590442,I590408,I1106047);
nand I_34521 (I590459,I590442,I1106026);
nor I_34522 (I590224,I590459,I590408);
and I_34523 (I590215,I590301,I590459);
not I_34524 (I590504,I590459);
nand I_34525 (I590218,I590301,I590504);
nor I_34526 (I590212,I590267,I590459);
not I_34527 (I590549,I1106032);
nor I_34528 (I590566,I590549,I1106047);
nand I_34529 (I590583,I590566,I590408);
nor I_34530 (I590221,I590326,I590583);
nor I_34531 (I590614,I590549,I1106038);
and I_34532 (I590631,I590614,I1106035);
or I_34533 (I590648,I590631,I1106041);
DFFARX1 I_34534 (I590648,I3563,I590241,I590674,);
nor I_34535 (I590682,I590674,I590425);
DFFARX1 I_34536 (I590682,I3563,I590241,I590209,);
DFFARX1 I_34537 (I590674,I3563,I590241,I590233,);
not I_34538 (I590727,I590674);
nor I_34539 (I590744,I590727,I590301);
nor I_34540 (I590761,I590566,I590744);
DFFARX1 I_34541 (I590761,I3563,I590241,I590230,);
not I_34542 (I590819,I3570);
DFFARX1 I_34543 (I1358303,I3563,I590819,I590845,);
not I_34544 (I590853,I590845);
DFFARX1 I_34545 (I1358303,I3563,I590819,I590879,);
not I_34546 (I590887,I1358327);
nand I_34547 (I590904,I590887,I1358309);
not I_34548 (I590921,I590904);
nor I_34549 (I590938,I590921,I1358324);
nor I_34550 (I590955,I590853,I590938);
DFFARX1 I_34551 (I590955,I3563,I590819,I590805,);
not I_34552 (I590986,I1358324);
nand I_34553 (I591003,I590986,I590921);
and I_34554 (I591020,I590986,I1358306);
nand I_34555 (I591037,I591020,I1358315);
nor I_34556 (I590802,I591037,I590986);
and I_34557 (I590793,I590879,I591037);
not I_34558 (I591082,I591037);
nand I_34559 (I590796,I590879,I591082);
nor I_34560 (I590790,I590845,I591037);
not I_34561 (I591127,I1358312);
nor I_34562 (I591144,I591127,I1358306);
nand I_34563 (I591161,I591144,I590986);
nor I_34564 (I590799,I590904,I591161);
nor I_34565 (I591192,I591127,I1358321);
and I_34566 (I591209,I591192,I1358330);
or I_34567 (I591226,I591209,I1358318);
DFFARX1 I_34568 (I591226,I3563,I590819,I591252,);
nor I_34569 (I591260,I591252,I591003);
DFFARX1 I_34570 (I591260,I3563,I590819,I590787,);
DFFARX1 I_34571 (I591252,I3563,I590819,I590811,);
not I_34572 (I591305,I591252);
nor I_34573 (I591322,I591305,I590879);
nor I_34574 (I591339,I591144,I591322);
DFFARX1 I_34575 (I591339,I3563,I590819,I590808,);
not I_34576 (I591397,I3570);
DFFARX1 I_34577 (I1160355,I3563,I591397,I591423,);
not I_34578 (I591431,I591423);
DFFARX1 I_34579 (I1160361,I3563,I591397,I591457,);
not I_34580 (I591465,I1160355);
nand I_34581 (I591482,I591465,I1160358);
not I_34582 (I591499,I591482);
nor I_34583 (I591516,I591499,I1160376);
nor I_34584 (I591533,I591431,I591516);
DFFARX1 I_34585 (I591533,I3563,I591397,I591383,);
not I_34586 (I591564,I1160376);
nand I_34587 (I591581,I591564,I591499);
and I_34588 (I591598,I591564,I1160379);
nand I_34589 (I591615,I591598,I1160358);
nor I_34590 (I591380,I591615,I591564);
and I_34591 (I591371,I591457,I591615);
not I_34592 (I591660,I591615);
nand I_34593 (I591374,I591457,I591660);
nor I_34594 (I591368,I591423,I591615);
not I_34595 (I591705,I1160364);
nor I_34596 (I591722,I591705,I1160379);
nand I_34597 (I591739,I591722,I591564);
nor I_34598 (I591377,I591482,I591739);
nor I_34599 (I591770,I591705,I1160370);
and I_34600 (I591787,I591770,I1160367);
or I_34601 (I591804,I591787,I1160373);
DFFARX1 I_34602 (I591804,I3563,I591397,I591830,);
nor I_34603 (I591838,I591830,I591581);
DFFARX1 I_34604 (I591838,I3563,I591397,I591365,);
DFFARX1 I_34605 (I591830,I3563,I591397,I591389,);
not I_34606 (I591883,I591830);
nor I_34607 (I591900,I591883,I591457);
nor I_34608 (I591917,I591722,I591900);
DFFARX1 I_34609 (I591917,I3563,I591397,I591386,);
not I_34610 (I591975,I3570);
DFFARX1 I_34611 (I186933,I3563,I591975,I592001,);
not I_34612 (I592009,I592001);
DFFARX1 I_34613 (I186918,I3563,I591975,I592035,);
not I_34614 (I592043,I186936);
nand I_34615 (I592060,I592043,I186921);
not I_34616 (I592077,I592060);
nor I_34617 (I592094,I592077,I186918);
nor I_34618 (I592111,I592009,I592094);
DFFARX1 I_34619 (I592111,I3563,I591975,I591961,);
not I_34620 (I592142,I186918);
nand I_34621 (I592159,I592142,I592077);
and I_34622 (I592176,I592142,I186921);
nand I_34623 (I592193,I592176,I186942);
nor I_34624 (I591958,I592193,I592142);
and I_34625 (I591949,I592035,I592193);
not I_34626 (I592238,I592193);
nand I_34627 (I591952,I592035,I592238);
nor I_34628 (I591946,I592001,I592193);
not I_34629 (I592283,I186930);
nor I_34630 (I592300,I592283,I186921);
nand I_34631 (I592317,I592300,I592142);
nor I_34632 (I591955,I592060,I592317);
nor I_34633 (I592348,I592283,I186924);
and I_34634 (I592365,I592348,I186939);
or I_34635 (I592382,I592365,I186927);
DFFARX1 I_34636 (I592382,I3563,I591975,I592408,);
nor I_34637 (I592416,I592408,I592159);
DFFARX1 I_34638 (I592416,I3563,I591975,I591943,);
DFFARX1 I_34639 (I592408,I3563,I591975,I591967,);
not I_34640 (I592461,I592408);
nor I_34641 (I592478,I592461,I592035);
nor I_34642 (I592495,I592300,I592478);
DFFARX1 I_34643 (I592495,I3563,I591975,I591964,);
not I_34644 (I592553,I3570);
DFFARX1 I_34645 (I1263291,I3563,I592553,I592579,);
not I_34646 (I592587,I592579);
DFFARX1 I_34647 (I1263285,I3563,I592553,I592613,);
not I_34648 (I592621,I1263294);
nand I_34649 (I592638,I592621,I1263273);
not I_34650 (I592655,I592638);
nor I_34651 (I592672,I592655,I1263282);
nor I_34652 (I592689,I592587,I592672);
DFFARX1 I_34653 (I592689,I3563,I592553,I592539,);
not I_34654 (I592720,I1263282);
nand I_34655 (I592737,I592720,I592655);
and I_34656 (I592754,I592720,I1263297);
nand I_34657 (I592771,I592754,I1263276);
nor I_34658 (I592536,I592771,I592720);
and I_34659 (I592527,I592613,I592771);
not I_34660 (I592816,I592771);
nand I_34661 (I592530,I592613,I592816);
nor I_34662 (I592524,I592579,I592771);
not I_34663 (I592861,I1263279);
nor I_34664 (I592878,I592861,I1263297);
nand I_34665 (I592895,I592878,I592720);
nor I_34666 (I592533,I592638,I592895);
nor I_34667 (I592926,I592861,I1263288);
and I_34668 (I592943,I592926,I1263276);
or I_34669 (I592960,I592943,I1263273);
DFFARX1 I_34670 (I592960,I3563,I592553,I592986,);
nor I_34671 (I592994,I592986,I592737);
DFFARX1 I_34672 (I592994,I3563,I592553,I592521,);
DFFARX1 I_34673 (I592986,I3563,I592553,I592545,);
not I_34674 (I593039,I592986);
nor I_34675 (I593056,I593039,I592613);
nor I_34676 (I593073,I592878,I593056);
DFFARX1 I_34677 (I593073,I3563,I592553,I592542,);
not I_34678 (I593131,I3570);
DFFARX1 I_34679 (I303289,I3563,I593131,I593157,);
not I_34680 (I593165,I593157);
DFFARX1 I_34681 (I303304,I3563,I593131,I593191,);
not I_34682 (I593199,I303307);
nand I_34683 (I593216,I593199,I303286);
not I_34684 (I593233,I593216);
nor I_34685 (I593250,I593233,I303310);
nor I_34686 (I593267,I593165,I593250);
DFFARX1 I_34687 (I593267,I3563,I593131,I593117,);
not I_34688 (I593298,I303310);
nand I_34689 (I593315,I593298,I593233);
and I_34690 (I593332,I593298,I303292);
nand I_34691 (I593349,I593332,I303283);
nor I_34692 (I593114,I593349,I593298);
and I_34693 (I593105,I593191,I593349);
not I_34694 (I593394,I593349);
nand I_34695 (I593108,I593191,I593394);
nor I_34696 (I593102,I593157,I593349);
not I_34697 (I593439,I303283);
nor I_34698 (I593456,I593439,I303292);
nand I_34699 (I593473,I593456,I593298);
nor I_34700 (I593111,I593216,I593473);
nor I_34701 (I593504,I593439,I303298);
and I_34702 (I593521,I593504,I303301);
or I_34703 (I593538,I593521,I303295);
DFFARX1 I_34704 (I593538,I3563,I593131,I593564,);
nor I_34705 (I593572,I593564,I593315);
DFFARX1 I_34706 (I593572,I3563,I593131,I593099,);
DFFARX1 I_34707 (I593564,I3563,I593131,I593123,);
not I_34708 (I593617,I593564);
nor I_34709 (I593634,I593617,I593191);
nor I_34710 (I593651,I593456,I593634);
DFFARX1 I_34711 (I593651,I3563,I593131,I593120,);
not I_34712 (I593709,I3570);
DFFARX1 I_34713 (I786151,I3563,I593709,I593735,);
not I_34714 (I593743,I593735);
DFFARX1 I_34715 (I786163,I3563,I593709,I593769,);
not I_34716 (I593777,I786154);
nand I_34717 (I593794,I593777,I786157);
not I_34718 (I593811,I593794);
nor I_34719 (I593828,I593811,I786160);
nor I_34720 (I593845,I593743,I593828);
DFFARX1 I_34721 (I593845,I3563,I593709,I593695,);
not I_34722 (I593876,I786160);
nand I_34723 (I593893,I593876,I593811);
and I_34724 (I593910,I593876,I786154);
nand I_34725 (I593927,I593910,I786166);
nor I_34726 (I593692,I593927,I593876);
and I_34727 (I593683,I593769,I593927);
not I_34728 (I593972,I593927);
nand I_34729 (I593686,I593769,I593972);
nor I_34730 (I593680,I593735,I593927);
not I_34731 (I594017,I786172);
nor I_34732 (I594034,I594017,I786154);
nand I_34733 (I594051,I594034,I593876);
nor I_34734 (I593689,I593794,I594051);
nor I_34735 (I594082,I594017,I786151);
and I_34736 (I594099,I594082,I786169);
or I_34737 (I594116,I594099,I786175);
DFFARX1 I_34738 (I594116,I3563,I593709,I594142,);
nor I_34739 (I594150,I594142,I593893);
DFFARX1 I_34740 (I594150,I3563,I593709,I593677,);
DFFARX1 I_34741 (I594142,I3563,I593709,I593701,);
not I_34742 (I594195,I594142);
nor I_34743 (I594212,I594195,I593769);
nor I_34744 (I594229,I594034,I594212);
DFFARX1 I_34745 (I594229,I3563,I593709,I593698,);
not I_34746 (I594287,I3570);
DFFARX1 I_34747 (I190503,I3563,I594287,I594313,);
not I_34748 (I594321,I594313);
DFFARX1 I_34749 (I190488,I3563,I594287,I594347,);
not I_34750 (I594355,I190506);
nand I_34751 (I594372,I594355,I190491);
not I_34752 (I594389,I594372);
nor I_34753 (I594406,I594389,I190488);
nor I_34754 (I594423,I594321,I594406);
DFFARX1 I_34755 (I594423,I3563,I594287,I594273,);
not I_34756 (I594454,I190488);
nand I_34757 (I594471,I594454,I594389);
and I_34758 (I594488,I594454,I190491);
nand I_34759 (I594505,I594488,I190512);
nor I_34760 (I594270,I594505,I594454);
and I_34761 (I594261,I594347,I594505);
not I_34762 (I594550,I594505);
nand I_34763 (I594264,I594347,I594550);
nor I_34764 (I594258,I594313,I594505);
not I_34765 (I594595,I190500);
nor I_34766 (I594612,I594595,I190491);
nand I_34767 (I594629,I594612,I594454);
nor I_34768 (I594267,I594372,I594629);
nor I_34769 (I594660,I594595,I190494);
and I_34770 (I594677,I594660,I190509);
or I_34771 (I594694,I594677,I190497);
DFFARX1 I_34772 (I594694,I3563,I594287,I594720,);
nor I_34773 (I594728,I594720,I594471);
DFFARX1 I_34774 (I594728,I3563,I594287,I594255,);
DFFARX1 I_34775 (I594720,I3563,I594287,I594279,);
not I_34776 (I594773,I594720);
nor I_34777 (I594790,I594773,I594347);
nor I_34778 (I594807,I594612,I594790);
DFFARX1 I_34779 (I594807,I3563,I594287,I594276,);
not I_34780 (I594865,I3570);
DFFARX1 I_34781 (I375488,I3563,I594865,I594891,);
not I_34782 (I594899,I594891);
DFFARX1 I_34783 (I375503,I3563,I594865,I594925,);
not I_34784 (I594933,I375506);
nand I_34785 (I594950,I594933,I375485);
not I_34786 (I594967,I594950);
nor I_34787 (I594984,I594967,I375509);
nor I_34788 (I595001,I594899,I594984);
DFFARX1 I_34789 (I595001,I3563,I594865,I594851,);
not I_34790 (I595032,I375509);
nand I_34791 (I595049,I595032,I594967);
and I_34792 (I595066,I595032,I375491);
nand I_34793 (I595083,I595066,I375482);
nor I_34794 (I594848,I595083,I595032);
and I_34795 (I594839,I594925,I595083);
not I_34796 (I595128,I595083);
nand I_34797 (I594842,I594925,I595128);
nor I_34798 (I594836,I594891,I595083);
not I_34799 (I595173,I375482);
nor I_34800 (I595190,I595173,I375491);
nand I_34801 (I595207,I595190,I595032);
nor I_34802 (I594845,I594950,I595207);
nor I_34803 (I595238,I595173,I375497);
and I_34804 (I595255,I595238,I375500);
or I_34805 (I595272,I595255,I375494);
DFFARX1 I_34806 (I595272,I3563,I594865,I595298,);
nor I_34807 (I595306,I595298,I595049);
DFFARX1 I_34808 (I595306,I3563,I594865,I594833,);
DFFARX1 I_34809 (I595298,I3563,I594865,I594857,);
not I_34810 (I595351,I595298);
nor I_34811 (I595368,I595351,I594925);
nor I_34812 (I595385,I595190,I595368);
DFFARX1 I_34813 (I595385,I3563,I594865,I594854,);
not I_34814 (I595443,I3570);
DFFARX1 I_34815 (I85129,I3563,I595443,I595469,);
not I_34816 (I595477,I595469);
DFFARX1 I_34817 (I85108,I3563,I595443,I595503,);
not I_34818 (I595511,I85105);
nand I_34819 (I595528,I595511,I85120);
not I_34820 (I595545,I595528);
nor I_34821 (I595562,I595545,I85108);
nor I_34822 (I595579,I595477,I595562);
DFFARX1 I_34823 (I595579,I3563,I595443,I595429,);
not I_34824 (I595610,I85108);
nand I_34825 (I595627,I595610,I595545);
and I_34826 (I595644,I595610,I85111);
nand I_34827 (I595661,I595644,I85126);
nor I_34828 (I595426,I595661,I595610);
and I_34829 (I595417,I595503,I595661);
not I_34830 (I595706,I595661);
nand I_34831 (I595420,I595503,I595706);
nor I_34832 (I595414,I595469,I595661);
not I_34833 (I595751,I85117);
nor I_34834 (I595768,I595751,I85111);
nand I_34835 (I595785,I595768,I595610);
nor I_34836 (I595423,I595528,I595785);
nor I_34837 (I595816,I595751,I85105);
and I_34838 (I595833,I595816,I85114);
or I_34839 (I595850,I595833,I85123);
DFFARX1 I_34840 (I595850,I3563,I595443,I595876,);
nor I_34841 (I595884,I595876,I595627);
DFFARX1 I_34842 (I595884,I3563,I595443,I595411,);
DFFARX1 I_34843 (I595876,I3563,I595443,I595435,);
not I_34844 (I595929,I595876);
nor I_34845 (I595946,I595929,I595503);
nor I_34846 (I595963,I595768,I595946);
DFFARX1 I_34847 (I595963,I3563,I595443,I595432,);
not I_34848 (I596021,I3570);
DFFARX1 I_34849 (I1201971,I3563,I596021,I596047,);
not I_34850 (I596055,I596047);
DFFARX1 I_34851 (I1201977,I3563,I596021,I596081,);
not I_34852 (I596089,I1201971);
nand I_34853 (I596106,I596089,I1201974);
not I_34854 (I596123,I596106);
nor I_34855 (I596140,I596123,I1201992);
nor I_34856 (I596157,I596055,I596140);
DFFARX1 I_34857 (I596157,I3563,I596021,I596007,);
not I_34858 (I596188,I1201992);
nand I_34859 (I596205,I596188,I596123);
and I_34860 (I596222,I596188,I1201995);
nand I_34861 (I596239,I596222,I1201974);
nor I_34862 (I596004,I596239,I596188);
and I_34863 (I595995,I596081,I596239);
not I_34864 (I596284,I596239);
nand I_34865 (I595998,I596081,I596284);
nor I_34866 (I595992,I596047,I596239);
not I_34867 (I596329,I1201980);
nor I_34868 (I596346,I596329,I1201995);
nand I_34869 (I596363,I596346,I596188);
nor I_34870 (I596001,I596106,I596363);
nor I_34871 (I596394,I596329,I1201986);
and I_34872 (I596411,I596394,I1201983);
or I_34873 (I596428,I596411,I1201989);
DFFARX1 I_34874 (I596428,I3563,I596021,I596454,);
nor I_34875 (I596462,I596454,I596205);
DFFARX1 I_34876 (I596462,I3563,I596021,I595989,);
DFFARX1 I_34877 (I596454,I3563,I596021,I596013,);
not I_34878 (I596507,I596454);
nor I_34879 (I596524,I596507,I596081);
nor I_34880 (I596541,I596346,I596524);
DFFARX1 I_34881 (I596541,I3563,I596021,I596010,);
not I_34882 (I596599,I3570);
DFFARX1 I_34883 (I700607,I3563,I596599,I596625,);
not I_34884 (I596633,I596625);
DFFARX1 I_34885 (I700619,I3563,I596599,I596659,);
not I_34886 (I596667,I700610);
nand I_34887 (I596684,I596667,I700613);
not I_34888 (I596701,I596684);
nor I_34889 (I596718,I596701,I700616);
nor I_34890 (I596735,I596633,I596718);
DFFARX1 I_34891 (I596735,I3563,I596599,I596585,);
not I_34892 (I596766,I700616);
nand I_34893 (I596783,I596766,I596701);
and I_34894 (I596800,I596766,I700610);
nand I_34895 (I596817,I596800,I700622);
nor I_34896 (I596582,I596817,I596766);
and I_34897 (I596573,I596659,I596817);
not I_34898 (I596862,I596817);
nand I_34899 (I596576,I596659,I596862);
nor I_34900 (I596570,I596625,I596817);
not I_34901 (I596907,I700628);
nor I_34902 (I596924,I596907,I700610);
nand I_34903 (I596941,I596924,I596766);
nor I_34904 (I596579,I596684,I596941);
nor I_34905 (I596972,I596907,I700607);
and I_34906 (I596989,I596972,I700625);
or I_34907 (I597006,I596989,I700631);
DFFARX1 I_34908 (I597006,I3563,I596599,I597032,);
nor I_34909 (I597040,I597032,I596783);
DFFARX1 I_34910 (I597040,I3563,I596599,I596567,);
DFFARX1 I_34911 (I597032,I3563,I596599,I596591,);
not I_34912 (I597085,I597032);
nor I_34913 (I597102,I597085,I596659);
nor I_34914 (I597119,I596924,I597102);
DFFARX1 I_34915 (I597119,I3563,I596599,I596588,);
not I_34916 (I597177,I3570);
DFFARX1 I_34917 (I186338,I3563,I597177,I597203,);
not I_34918 (I597211,I597203);
DFFARX1 I_34919 (I186323,I3563,I597177,I597237,);
not I_34920 (I597245,I186341);
nand I_34921 (I597262,I597245,I186326);
not I_34922 (I597279,I597262);
nor I_34923 (I597296,I597279,I186323);
nor I_34924 (I597313,I597211,I597296);
DFFARX1 I_34925 (I597313,I3563,I597177,I597163,);
not I_34926 (I597344,I186323);
nand I_34927 (I597361,I597344,I597279);
and I_34928 (I597378,I597344,I186326);
nand I_34929 (I597395,I597378,I186347);
nor I_34930 (I597160,I597395,I597344);
and I_34931 (I597151,I597237,I597395);
not I_34932 (I597440,I597395);
nand I_34933 (I597154,I597237,I597440);
nor I_34934 (I597148,I597203,I597395);
not I_34935 (I597485,I186335);
nor I_34936 (I597502,I597485,I186326);
nand I_34937 (I597519,I597502,I597344);
nor I_34938 (I597157,I597262,I597519);
nor I_34939 (I597550,I597485,I186329);
and I_34940 (I597567,I597550,I186344);
or I_34941 (I597584,I597567,I186332);
DFFARX1 I_34942 (I597584,I3563,I597177,I597610,);
nor I_34943 (I597618,I597610,I597361);
DFFARX1 I_34944 (I597618,I3563,I597177,I597145,);
DFFARX1 I_34945 (I597610,I3563,I597177,I597169,);
not I_34946 (I597663,I597610);
nor I_34947 (I597680,I597663,I597237);
nor I_34948 (I597697,I597502,I597680);
DFFARX1 I_34949 (I597697,I3563,I597177,I597166,);
not I_34950 (I597755,I3570);
DFFARX1 I_34951 (I393406,I3563,I597755,I597781,);
not I_34952 (I597789,I597781);
DFFARX1 I_34953 (I393421,I3563,I597755,I597815,);
not I_34954 (I597823,I393424);
nand I_34955 (I597840,I597823,I393403);
not I_34956 (I597857,I597840);
nor I_34957 (I597874,I597857,I393427);
nor I_34958 (I597891,I597789,I597874);
DFFARX1 I_34959 (I597891,I3563,I597755,I597741,);
not I_34960 (I597922,I393427);
nand I_34961 (I597939,I597922,I597857);
and I_34962 (I597956,I597922,I393409);
nand I_34963 (I597973,I597956,I393400);
nor I_34964 (I597738,I597973,I597922);
and I_34965 (I597729,I597815,I597973);
not I_34966 (I598018,I597973);
nand I_34967 (I597732,I597815,I598018);
nor I_34968 (I597726,I597781,I597973);
not I_34969 (I598063,I393400);
nor I_34970 (I598080,I598063,I393409);
nand I_34971 (I598097,I598080,I597922);
nor I_34972 (I597735,I597840,I598097);
nor I_34973 (I598128,I598063,I393415);
and I_34974 (I598145,I598128,I393418);
or I_34975 (I598162,I598145,I393412);
DFFARX1 I_34976 (I598162,I3563,I597755,I598188,);
nor I_34977 (I598196,I598188,I597939);
DFFARX1 I_34978 (I598196,I3563,I597755,I597723,);
DFFARX1 I_34979 (I598188,I3563,I597755,I597747,);
not I_34980 (I598241,I598188);
nor I_34981 (I598258,I598241,I597815);
nor I_34982 (I598275,I598080,I598258);
DFFARX1 I_34983 (I598275,I3563,I597755,I597744,);
not I_34984 (I598333,I3570);
DFFARX1 I_34985 (I780371,I3563,I598333,I598359,);
not I_34986 (I598367,I598359);
DFFARX1 I_34987 (I780383,I3563,I598333,I598393,);
not I_34988 (I598401,I780374);
nand I_34989 (I598418,I598401,I780377);
not I_34990 (I598435,I598418);
nor I_34991 (I598452,I598435,I780380);
nor I_34992 (I598469,I598367,I598452);
DFFARX1 I_34993 (I598469,I3563,I598333,I598319,);
not I_34994 (I598500,I780380);
nand I_34995 (I598517,I598500,I598435);
and I_34996 (I598534,I598500,I780374);
nand I_34997 (I598551,I598534,I780386);
nor I_34998 (I598316,I598551,I598500);
and I_34999 (I598307,I598393,I598551);
not I_35000 (I598596,I598551);
nand I_35001 (I598310,I598393,I598596);
nor I_35002 (I598304,I598359,I598551);
not I_35003 (I598641,I780392);
nor I_35004 (I598658,I598641,I780374);
nand I_35005 (I598675,I598658,I598500);
nor I_35006 (I598313,I598418,I598675);
nor I_35007 (I598706,I598641,I780371);
and I_35008 (I598723,I598706,I780389);
or I_35009 (I598740,I598723,I780395);
DFFARX1 I_35010 (I598740,I3563,I598333,I598766,);
nor I_35011 (I598774,I598766,I598517);
DFFARX1 I_35012 (I598774,I3563,I598333,I598301,);
DFFARX1 I_35013 (I598766,I3563,I598333,I598325,);
not I_35014 (I598819,I598766);
nor I_35015 (I598836,I598819,I598393);
nor I_35016 (I598853,I598658,I598836);
DFFARX1 I_35017 (I598853,I3563,I598333,I598322,);
not I_35018 (I598911,I3570);
DFFARX1 I_35019 (I349665,I3563,I598911,I598937,);
not I_35020 (I598945,I598937);
DFFARX1 I_35021 (I349680,I3563,I598911,I598971,);
not I_35022 (I598979,I349683);
nand I_35023 (I598996,I598979,I349662);
not I_35024 (I599013,I598996);
nor I_35025 (I599030,I599013,I349686);
nor I_35026 (I599047,I598945,I599030);
DFFARX1 I_35027 (I599047,I3563,I598911,I598897,);
not I_35028 (I599078,I349686);
nand I_35029 (I599095,I599078,I599013);
and I_35030 (I599112,I599078,I349668);
nand I_35031 (I599129,I599112,I349659);
nor I_35032 (I598894,I599129,I599078);
and I_35033 (I598885,I598971,I599129);
not I_35034 (I599174,I599129);
nand I_35035 (I598888,I598971,I599174);
nor I_35036 (I598882,I598937,I599129);
not I_35037 (I599219,I349659);
nor I_35038 (I599236,I599219,I349668);
nand I_35039 (I599253,I599236,I599078);
nor I_35040 (I598891,I598996,I599253);
nor I_35041 (I599284,I599219,I349674);
and I_35042 (I599301,I599284,I349677);
or I_35043 (I599318,I599301,I349671);
DFFARX1 I_35044 (I599318,I3563,I598911,I599344,);
nor I_35045 (I599352,I599344,I599095);
DFFARX1 I_35046 (I599352,I3563,I598911,I598879,);
DFFARX1 I_35047 (I599344,I3563,I598911,I598903,);
not I_35048 (I599397,I599344);
nor I_35049 (I599414,I599397,I598971);
nor I_35050 (I599431,I599236,I599414);
DFFARX1 I_35051 (I599431,I3563,I598911,I598900,);
not I_35052 (I599489,I3570);
DFFARX1 I_35053 (I548919,I3563,I599489,I599515,);
not I_35054 (I599523,I599515);
DFFARX1 I_35055 (I548931,I3563,I599489,I599549,);
not I_35056 (I599557,I548937);
nand I_35057 (I599574,I599557,I548928);
not I_35058 (I599591,I599574);
nor I_35059 (I599608,I599591,I548934);
nor I_35060 (I599625,I599523,I599608);
DFFARX1 I_35061 (I599625,I3563,I599489,I599475,);
not I_35062 (I599656,I548934);
nand I_35063 (I599673,I599656,I599591);
and I_35064 (I599690,I599656,I548925);
nand I_35065 (I599707,I599690,I548916);
nor I_35066 (I599472,I599707,I599656);
and I_35067 (I599463,I599549,I599707);
not I_35068 (I599752,I599707);
nand I_35069 (I599466,I599549,I599752);
nor I_35070 (I599460,I599515,I599707);
not I_35071 (I599797,I548922);
nor I_35072 (I599814,I599797,I548925);
nand I_35073 (I599831,I599814,I599656);
nor I_35074 (I599469,I599574,I599831);
nor I_35075 (I599862,I599797,I548919);
and I_35076 (I599879,I599862,I548916);
or I_35077 (I599896,I599879,I548940);
DFFARX1 I_35078 (I599896,I3563,I599489,I599922,);
nor I_35079 (I599930,I599922,I599673);
DFFARX1 I_35080 (I599930,I3563,I599489,I599457,);
DFFARX1 I_35081 (I599922,I3563,I599489,I599481,);
not I_35082 (I599975,I599922);
nor I_35083 (I599992,I599975,I599549);
nor I_35084 (I600009,I599814,I599992);
DFFARX1 I_35085 (I600009,I3563,I599489,I599478,);
not I_35086 (I600067,I3570);
DFFARX1 I_35087 (I1132033,I3563,I600067,I600093,);
not I_35088 (I600101,I600093);
DFFARX1 I_35089 (I1132039,I3563,I600067,I600127,);
not I_35090 (I600135,I1132033);
nand I_35091 (I600152,I600135,I1132036);
not I_35092 (I600169,I600152);
nor I_35093 (I600186,I600169,I1132054);
nor I_35094 (I600203,I600101,I600186);
DFFARX1 I_35095 (I600203,I3563,I600067,I600053,);
not I_35096 (I600234,I1132054);
nand I_35097 (I600251,I600234,I600169);
and I_35098 (I600268,I600234,I1132057);
nand I_35099 (I600285,I600268,I1132036);
nor I_35100 (I600050,I600285,I600234);
and I_35101 (I600041,I600127,I600285);
not I_35102 (I600330,I600285);
nand I_35103 (I600044,I600127,I600330);
nor I_35104 (I600038,I600093,I600285);
not I_35105 (I600375,I1132042);
nor I_35106 (I600392,I600375,I1132057);
nand I_35107 (I600409,I600392,I600234);
nor I_35108 (I600047,I600152,I600409);
nor I_35109 (I600440,I600375,I1132048);
and I_35110 (I600457,I600440,I1132045);
or I_35111 (I600474,I600457,I1132051);
DFFARX1 I_35112 (I600474,I3563,I600067,I600500,);
nor I_35113 (I600508,I600500,I600251);
DFFARX1 I_35114 (I600508,I3563,I600067,I600035,);
DFFARX1 I_35115 (I600500,I3563,I600067,I600059,);
not I_35116 (I600553,I600500);
nor I_35117 (I600570,I600553,I600127);
nor I_35118 (I600587,I600392,I600570);
DFFARX1 I_35119 (I600587,I3563,I600067,I600056,);
not I_35120 (I600645,I3570);
DFFARX1 I_35121 (I1370798,I3563,I600645,I600671,);
not I_35122 (I600679,I600671);
DFFARX1 I_35123 (I1370798,I3563,I600645,I600705,);
not I_35124 (I600713,I1370822);
nand I_35125 (I600730,I600713,I1370804);
not I_35126 (I600747,I600730);
nor I_35127 (I600764,I600747,I1370819);
nor I_35128 (I600781,I600679,I600764);
DFFARX1 I_35129 (I600781,I3563,I600645,I600631,);
not I_35130 (I600812,I1370819);
nand I_35131 (I600829,I600812,I600747);
and I_35132 (I600846,I600812,I1370801);
nand I_35133 (I600863,I600846,I1370810);
nor I_35134 (I600628,I600863,I600812);
and I_35135 (I600619,I600705,I600863);
not I_35136 (I600908,I600863);
nand I_35137 (I600622,I600705,I600908);
nor I_35138 (I600616,I600671,I600863);
not I_35139 (I600953,I1370807);
nor I_35140 (I600970,I600953,I1370801);
nand I_35141 (I600987,I600970,I600812);
nor I_35142 (I600625,I600730,I600987);
nor I_35143 (I601018,I600953,I1370816);
and I_35144 (I601035,I601018,I1370825);
or I_35145 (I601052,I601035,I1370813);
DFFARX1 I_35146 (I601052,I3563,I600645,I601078,);
nor I_35147 (I601086,I601078,I600829);
DFFARX1 I_35148 (I601086,I3563,I600645,I600613,);
DFFARX1 I_35149 (I601078,I3563,I600645,I600637,);
not I_35150 (I601131,I601078);
nor I_35151 (I601148,I601131,I600705);
nor I_35152 (I601165,I600970,I601148);
DFFARX1 I_35153 (I601165,I3563,I600645,I600634,);
not I_35154 (I601223,I3570);
DFFARX1 I_35155 (I331220,I3563,I601223,I601249,);
not I_35156 (I601257,I601249);
DFFARX1 I_35157 (I331235,I3563,I601223,I601283,);
not I_35158 (I601291,I331238);
nand I_35159 (I601308,I601291,I331217);
not I_35160 (I601325,I601308);
nor I_35161 (I601342,I601325,I331241);
nor I_35162 (I601359,I601257,I601342);
DFFARX1 I_35163 (I601359,I3563,I601223,I601209,);
not I_35164 (I601390,I331241);
nand I_35165 (I601407,I601390,I601325);
and I_35166 (I601424,I601390,I331223);
nand I_35167 (I601441,I601424,I331214);
nor I_35168 (I601206,I601441,I601390);
and I_35169 (I601197,I601283,I601441);
not I_35170 (I601486,I601441);
nand I_35171 (I601200,I601283,I601486);
nor I_35172 (I601194,I601249,I601441);
not I_35173 (I601531,I331214);
nor I_35174 (I601548,I601531,I331223);
nand I_35175 (I601565,I601548,I601390);
nor I_35176 (I601203,I601308,I601565);
nor I_35177 (I601596,I601531,I331229);
and I_35178 (I601613,I601596,I331232);
or I_35179 (I601630,I601613,I331226);
DFFARX1 I_35180 (I601630,I3563,I601223,I601656,);
nor I_35181 (I601664,I601656,I601407);
DFFARX1 I_35182 (I601664,I3563,I601223,I601191,);
DFFARX1 I_35183 (I601656,I3563,I601223,I601215,);
not I_35184 (I601709,I601656);
nor I_35185 (I601726,I601709,I601283);
nor I_35186 (I601743,I601548,I601726);
DFFARX1 I_35187 (I601743,I3563,I601223,I601212,);
not I_35188 (I601801,I3570);
DFFARX1 I_35189 (I314883,I3563,I601801,I601827,);
not I_35190 (I601835,I601827);
DFFARX1 I_35191 (I314898,I3563,I601801,I601861,);
not I_35192 (I601869,I314901);
nand I_35193 (I601886,I601869,I314880);
not I_35194 (I601903,I601886);
nor I_35195 (I601920,I601903,I314904);
nor I_35196 (I601937,I601835,I601920);
DFFARX1 I_35197 (I601937,I3563,I601801,I601787,);
not I_35198 (I601968,I314904);
nand I_35199 (I601985,I601968,I601903);
and I_35200 (I602002,I601968,I314886);
nand I_35201 (I602019,I602002,I314877);
nor I_35202 (I601784,I602019,I601968);
and I_35203 (I601775,I601861,I602019);
not I_35204 (I602064,I602019);
nand I_35205 (I601778,I601861,I602064);
nor I_35206 (I601772,I601827,I602019);
not I_35207 (I602109,I314877);
nor I_35208 (I602126,I602109,I314886);
nand I_35209 (I602143,I602126,I601968);
nor I_35210 (I601781,I601886,I602143);
nor I_35211 (I602174,I602109,I314892);
and I_35212 (I602191,I602174,I314895);
or I_35213 (I602208,I602191,I314889);
DFFARX1 I_35214 (I602208,I3563,I601801,I602234,);
nor I_35215 (I602242,I602234,I601985);
DFFARX1 I_35216 (I602242,I3563,I601801,I601769,);
DFFARX1 I_35217 (I602234,I3563,I601801,I601793,);
not I_35218 (I602287,I602234);
nor I_35219 (I602304,I602287,I601861);
nor I_35220 (I602321,I602126,I602304);
DFFARX1 I_35221 (I602321,I3563,I601801,I601790,);
not I_35222 (I602379,I3570);
DFFARX1 I_35223 (I537614,I3563,I602379,I602405,);
not I_35224 (I602413,I602405);
DFFARX1 I_35225 (I537626,I3563,I602379,I602439,);
not I_35226 (I602447,I537632);
nand I_35227 (I602464,I602447,I537623);
not I_35228 (I602481,I602464);
nor I_35229 (I602498,I602481,I537629);
nor I_35230 (I602515,I602413,I602498);
DFFARX1 I_35231 (I602515,I3563,I602379,I602365,);
not I_35232 (I602546,I537629);
nand I_35233 (I602563,I602546,I602481);
and I_35234 (I602580,I602546,I537620);
nand I_35235 (I602597,I602580,I537611);
nor I_35236 (I602362,I602597,I602546);
and I_35237 (I602353,I602439,I602597);
not I_35238 (I602642,I602597);
nand I_35239 (I602356,I602439,I602642);
nor I_35240 (I602350,I602405,I602597);
not I_35241 (I602687,I537617);
nor I_35242 (I602704,I602687,I537620);
nand I_35243 (I602721,I602704,I602546);
nor I_35244 (I602359,I602464,I602721);
nor I_35245 (I602752,I602687,I537614);
and I_35246 (I602769,I602752,I537611);
or I_35247 (I602786,I602769,I537635);
DFFARX1 I_35248 (I602786,I3563,I602379,I602812,);
nor I_35249 (I602820,I602812,I602563);
DFFARX1 I_35250 (I602820,I3563,I602379,I602347,);
DFFARX1 I_35251 (I602812,I3563,I602379,I602371,);
not I_35252 (I602865,I602812);
nor I_35253 (I602882,I602865,I602439);
nor I_35254 (I602899,I602704,I602882);
DFFARX1 I_35255 (I602899,I3563,I602379,I602368,);
not I_35256 (I602957,I3570);
DFFARX1 I_35257 (I305924,I3563,I602957,I602983,);
not I_35258 (I602991,I602983);
DFFARX1 I_35259 (I305939,I3563,I602957,I603017,);
not I_35260 (I603025,I305942);
nand I_35261 (I603042,I603025,I305921);
not I_35262 (I603059,I603042);
nor I_35263 (I603076,I603059,I305945);
nor I_35264 (I603093,I602991,I603076);
DFFARX1 I_35265 (I603093,I3563,I602957,I602943,);
not I_35266 (I603124,I305945);
nand I_35267 (I603141,I603124,I603059);
and I_35268 (I603158,I603124,I305927);
nand I_35269 (I603175,I603158,I305918);
nor I_35270 (I602940,I603175,I603124);
and I_35271 (I602931,I603017,I603175);
not I_35272 (I603220,I603175);
nand I_35273 (I602934,I603017,I603220);
nor I_35274 (I602928,I602983,I603175);
not I_35275 (I603265,I305918);
nor I_35276 (I603282,I603265,I305927);
nand I_35277 (I603299,I603282,I603124);
nor I_35278 (I602937,I603042,I603299);
nor I_35279 (I603330,I603265,I305933);
and I_35280 (I603347,I603330,I305936);
or I_35281 (I603364,I603347,I305930);
DFFARX1 I_35282 (I603364,I3563,I602957,I603390,);
nor I_35283 (I603398,I603390,I603141);
DFFARX1 I_35284 (I603398,I3563,I602957,I602925,);
DFFARX1 I_35285 (I603390,I3563,I602957,I602949,);
not I_35286 (I603443,I603390);
nor I_35287 (I603460,I603443,I603017);
nor I_35288 (I603477,I603282,I603460);
DFFARX1 I_35289 (I603477,I3563,I602957,I602946,);
not I_35290 (I603535,I3570);
DFFARX1 I_35291 (I1140703,I3563,I603535,I603561,);
not I_35292 (I603569,I603561);
DFFARX1 I_35293 (I1140709,I3563,I603535,I603595,);
not I_35294 (I603603,I1140703);
nand I_35295 (I603620,I603603,I1140706);
not I_35296 (I603637,I603620);
nor I_35297 (I603654,I603637,I1140724);
nor I_35298 (I603671,I603569,I603654);
DFFARX1 I_35299 (I603671,I3563,I603535,I603521,);
not I_35300 (I603702,I1140724);
nand I_35301 (I603719,I603702,I603637);
and I_35302 (I603736,I603702,I1140727);
nand I_35303 (I603753,I603736,I1140706);
nor I_35304 (I603518,I603753,I603702);
and I_35305 (I603509,I603595,I603753);
not I_35306 (I603798,I603753);
nand I_35307 (I603512,I603595,I603798);
nor I_35308 (I603506,I603561,I603753);
not I_35309 (I603843,I1140712);
nor I_35310 (I603860,I603843,I1140727);
nand I_35311 (I603877,I603860,I603702);
nor I_35312 (I603515,I603620,I603877);
nor I_35313 (I603908,I603843,I1140718);
and I_35314 (I603925,I603908,I1140715);
or I_35315 (I603942,I603925,I1140721);
DFFARX1 I_35316 (I603942,I3563,I603535,I603968,);
nor I_35317 (I603976,I603968,I603719);
DFFARX1 I_35318 (I603976,I3563,I603535,I603503,);
DFFARX1 I_35319 (I603968,I3563,I603535,I603527,);
not I_35320 (I604021,I603968);
nor I_35321 (I604038,I604021,I603595);
nor I_35322 (I604055,I603860,I604038);
DFFARX1 I_35323 (I604055,I3563,I603535,I603524,);
not I_35324 (I604113,I3570);
DFFARX1 I_35325 (I3252,I3563,I604113,I604139,);
not I_35326 (I604147,I604139);
DFFARX1 I_35327 (I3060,I3563,I604113,I604173,);
not I_35328 (I604181,I3300);
nand I_35329 (I604198,I604181,I2884);
not I_35330 (I604215,I604198);
nor I_35331 (I604232,I604215,I1412);
nor I_35332 (I604249,I604147,I604232);
DFFARX1 I_35333 (I604249,I3563,I604113,I604099,);
not I_35334 (I604280,I1412);
nand I_35335 (I604297,I604280,I604215);
and I_35336 (I604314,I604280,I1652);
nand I_35337 (I604331,I604314,I1836);
nor I_35338 (I604096,I604331,I604280);
and I_35339 (I604087,I604173,I604331);
not I_35340 (I604376,I604331);
nand I_35341 (I604090,I604173,I604376);
nor I_35342 (I604084,I604139,I604331);
not I_35343 (I604421,I3140);
nor I_35344 (I604438,I604421,I1652);
nand I_35345 (I604455,I604438,I604280);
nor I_35346 (I604093,I604198,I604455);
nor I_35347 (I604486,I604421,I1396);
and I_35348 (I604503,I604486,I2540);
or I_35349 (I604520,I604503,I3268);
DFFARX1 I_35350 (I604520,I3563,I604113,I604546,);
nor I_35351 (I604554,I604546,I604297);
DFFARX1 I_35352 (I604554,I3563,I604113,I604081,);
DFFARX1 I_35353 (I604546,I3563,I604113,I604105,);
not I_35354 (I604599,I604546);
nor I_35355 (I604616,I604599,I604173);
nor I_35356 (I604633,I604438,I604616);
DFFARX1 I_35357 (I604633,I3563,I604113,I604102,);
not I_35358 (I604691,I3570);
DFFARX1 I_35359 (I785573,I3563,I604691,I604717,);
not I_35360 (I604725,I604717);
DFFARX1 I_35361 (I785585,I3563,I604691,I604751,);
not I_35362 (I604759,I785576);
nand I_35363 (I604776,I604759,I785579);
not I_35364 (I604793,I604776);
nor I_35365 (I604810,I604793,I785582);
nor I_35366 (I604827,I604725,I604810);
DFFARX1 I_35367 (I604827,I3563,I604691,I604677,);
not I_35368 (I604858,I785582);
nand I_35369 (I604875,I604858,I604793);
and I_35370 (I604892,I604858,I785576);
nand I_35371 (I604909,I604892,I785588);
nor I_35372 (I604674,I604909,I604858);
and I_35373 (I604665,I604751,I604909);
not I_35374 (I604954,I604909);
nand I_35375 (I604668,I604751,I604954);
nor I_35376 (I604662,I604717,I604909);
not I_35377 (I604999,I785594);
nor I_35378 (I605016,I604999,I785576);
nand I_35379 (I605033,I605016,I604858);
nor I_35380 (I604671,I604776,I605033);
nor I_35381 (I605064,I604999,I785573);
and I_35382 (I605081,I605064,I785591);
or I_35383 (I605098,I605081,I785597);
DFFARX1 I_35384 (I605098,I3563,I604691,I605124,);
nor I_35385 (I605132,I605124,I604875);
DFFARX1 I_35386 (I605132,I3563,I604691,I604659,);
DFFARX1 I_35387 (I605124,I3563,I604691,I604683,);
not I_35388 (I605177,I605124);
nor I_35389 (I605194,I605177,I604751);
nor I_35390 (I605211,I605016,I605194);
DFFARX1 I_35391 (I605211,I3563,I604691,I604680,);
not I_35392 (I605269,I3570);
DFFARX1 I_35393 (I1087633,I3563,I605269,I605295,);
not I_35394 (I605303,I605295);
DFFARX1 I_35395 (I1087624,I3563,I605269,I605329,);
not I_35396 (I605337,I1087618);
nand I_35397 (I605354,I605337,I1087630);
not I_35398 (I605371,I605354);
nor I_35399 (I605388,I605371,I1087621);
nor I_35400 (I605405,I605303,I605388);
DFFARX1 I_35401 (I605405,I3563,I605269,I605255,);
not I_35402 (I605436,I1087621);
nand I_35403 (I605453,I605436,I605371);
and I_35404 (I605470,I605436,I1087627);
nand I_35405 (I605487,I605470,I1087612);
nor I_35406 (I605252,I605487,I605436);
and I_35407 (I605243,I605329,I605487);
not I_35408 (I605532,I605487);
nand I_35409 (I605246,I605329,I605532);
nor I_35410 (I605240,I605295,I605487);
not I_35411 (I605577,I1087612);
nor I_35412 (I605594,I605577,I1087627);
nand I_35413 (I605611,I605594,I605436);
nor I_35414 (I605249,I605354,I605611);
nor I_35415 (I605642,I605577,I1087615);
and I_35416 (I605659,I605642,I1087618);
or I_35417 (I605676,I605659,I1087615);
DFFARX1 I_35418 (I605676,I3563,I605269,I605702,);
nor I_35419 (I605710,I605702,I605453);
DFFARX1 I_35420 (I605710,I3563,I605269,I605237,);
DFFARX1 I_35421 (I605702,I3563,I605269,I605261,);
not I_35422 (I605755,I605702);
nor I_35423 (I605772,I605755,I605329);
nor I_35424 (I605789,I605594,I605772);
DFFARX1 I_35425 (I605789,I3563,I605269,I605258,);
not I_35426 (I605847,I3570);
DFFARX1 I_35427 (I118857,I3563,I605847,I605873,);
not I_35428 (I605881,I605873);
DFFARX1 I_35429 (I118836,I3563,I605847,I605907,);
not I_35430 (I605915,I118833);
nand I_35431 (I605932,I605915,I118848);
not I_35432 (I605949,I605932);
nor I_35433 (I605966,I605949,I118836);
nor I_35434 (I605983,I605881,I605966);
DFFARX1 I_35435 (I605983,I3563,I605847,I605833,);
not I_35436 (I606014,I118836);
nand I_35437 (I606031,I606014,I605949);
and I_35438 (I606048,I606014,I118839);
nand I_35439 (I606065,I606048,I118854);
nor I_35440 (I605830,I606065,I606014);
and I_35441 (I605821,I605907,I606065);
not I_35442 (I606110,I606065);
nand I_35443 (I605824,I605907,I606110);
nor I_35444 (I605818,I605873,I606065);
not I_35445 (I606155,I118845);
nor I_35446 (I606172,I606155,I118839);
nand I_35447 (I606189,I606172,I606014);
nor I_35448 (I605827,I605932,I606189);
nor I_35449 (I606220,I606155,I118833);
and I_35450 (I606237,I606220,I118842);
or I_35451 (I606254,I606237,I118851);
DFFARX1 I_35452 (I606254,I3563,I605847,I606280,);
nor I_35453 (I606288,I606280,I606031);
DFFARX1 I_35454 (I606288,I3563,I605847,I605815,);
DFFARX1 I_35455 (I606280,I3563,I605847,I605839,);
not I_35456 (I606333,I606280);
nor I_35457 (I606350,I606333,I605907);
nor I_35458 (I606367,I606172,I606350);
DFFARX1 I_35459 (I606367,I3563,I605847,I605836,);
not I_35460 (I606425,I3570);
DFFARX1 I_35461 (I833723,I3563,I606425,I606451,);
not I_35462 (I606459,I606451);
DFFARX1 I_35463 (I833723,I3563,I606425,I606485,);
not I_35464 (I606493,I833720);
nand I_35465 (I606510,I606493,I833735);
not I_35466 (I606527,I606510);
nor I_35467 (I606544,I606527,I833729);
nor I_35468 (I606561,I606459,I606544);
DFFARX1 I_35469 (I606561,I3563,I606425,I606411,);
not I_35470 (I606592,I833729);
nand I_35471 (I606609,I606592,I606527);
and I_35472 (I606626,I606592,I833726);
nand I_35473 (I606643,I606626,I833717);
nor I_35474 (I606408,I606643,I606592);
and I_35475 (I606399,I606485,I606643);
not I_35476 (I606688,I606643);
nand I_35477 (I606402,I606485,I606688);
nor I_35478 (I606396,I606451,I606643);
not I_35479 (I606733,I833738);
nor I_35480 (I606750,I606733,I833726);
nand I_35481 (I606767,I606750,I606592);
nor I_35482 (I606405,I606510,I606767);
nor I_35483 (I606798,I606733,I833717);
and I_35484 (I606815,I606798,I833720);
or I_35485 (I606832,I606815,I833732);
DFFARX1 I_35486 (I606832,I3563,I606425,I606858,);
nor I_35487 (I606866,I606858,I606609);
DFFARX1 I_35488 (I606866,I3563,I606425,I606393,);
DFFARX1 I_35489 (I606858,I3563,I606425,I606417,);
not I_35490 (I606911,I606858);
nor I_35491 (I606928,I606911,I606485);
nor I_35492 (I606945,I606750,I606928);
DFFARX1 I_35493 (I606945,I3563,I606425,I606414,);
not I_35494 (I607003,I3570);
DFFARX1 I_35495 (I265473,I3563,I607003,I607029,);
not I_35496 (I607037,I607029);
DFFARX1 I_35497 (I265458,I3563,I607003,I607063,);
not I_35498 (I607071,I265476);
nand I_35499 (I607088,I607071,I265461);
not I_35500 (I607105,I607088);
nor I_35501 (I607122,I607105,I265458);
nor I_35502 (I607139,I607037,I607122);
DFFARX1 I_35503 (I607139,I3563,I607003,I606989,);
not I_35504 (I607170,I265458);
nand I_35505 (I607187,I607170,I607105);
and I_35506 (I607204,I607170,I265461);
nand I_35507 (I607221,I607204,I265482);
nor I_35508 (I606986,I607221,I607170);
and I_35509 (I606977,I607063,I607221);
not I_35510 (I607266,I607221);
nand I_35511 (I606980,I607063,I607266);
nor I_35512 (I606974,I607029,I607221);
not I_35513 (I607311,I265470);
nor I_35514 (I607328,I607311,I265461);
nand I_35515 (I607345,I607328,I607170);
nor I_35516 (I606983,I607088,I607345);
nor I_35517 (I607376,I607311,I265464);
and I_35518 (I607393,I607376,I265479);
or I_35519 (I607410,I607393,I265467);
DFFARX1 I_35520 (I607410,I3563,I607003,I607436,);
nor I_35521 (I607444,I607436,I607187);
DFFARX1 I_35522 (I607444,I3563,I607003,I606971,);
DFFARX1 I_35523 (I607436,I3563,I607003,I606995,);
not I_35524 (I607489,I607436);
nor I_35525 (I607506,I607489,I607063);
nor I_35526 (I607523,I607328,I607506);
DFFARX1 I_35527 (I607523,I3563,I607003,I606992,);
not I_35528 (I607581,I3570);
DFFARX1 I_35529 (I40313,I3563,I607581,I607607,);
not I_35530 (I607615,I607607);
DFFARX1 I_35531 (I40316,I3563,I607581,I607641,);
not I_35532 (I607649,I40310);
nand I_35533 (I607666,I607649,I40334);
not I_35534 (I607683,I607666);
nor I_35535 (I607700,I607683,I40313);
nor I_35536 (I607717,I607615,I607700);
DFFARX1 I_35537 (I607717,I3563,I607581,I607567,);
not I_35538 (I607748,I40313);
nand I_35539 (I607765,I607748,I607683);
and I_35540 (I607782,I607748,I40328);
nand I_35541 (I607799,I607782,I40322);
nor I_35542 (I607564,I607799,I607748);
and I_35543 (I607555,I607641,I607799);
not I_35544 (I607844,I607799);
nand I_35545 (I607558,I607641,I607844);
nor I_35546 (I607552,I607607,I607799);
not I_35547 (I607889,I40331);
nor I_35548 (I607906,I607889,I40328);
nand I_35549 (I607923,I607906,I607748);
nor I_35550 (I607561,I607666,I607923);
nor I_35551 (I607954,I607889,I40310);
and I_35552 (I607971,I607954,I40319);
or I_35553 (I607988,I607971,I40325);
DFFARX1 I_35554 (I607988,I3563,I607581,I608014,);
nor I_35555 (I608022,I608014,I607765);
DFFARX1 I_35556 (I608022,I3563,I607581,I607549,);
DFFARX1 I_35557 (I608014,I3563,I607581,I607573,);
not I_35558 (I608067,I608014);
nor I_35559 (I608084,I608067,I607641);
nor I_35560 (I608101,I607906,I608084);
DFFARX1 I_35561 (I608101,I3563,I607581,I607570,);
not I_35562 (I608159,I3570);
DFFARX1 I_35563 (I119911,I3563,I608159,I608185,);
not I_35564 (I608193,I608185);
DFFARX1 I_35565 (I119890,I3563,I608159,I608219,);
not I_35566 (I608227,I119887);
nand I_35567 (I608244,I608227,I119902);
not I_35568 (I608261,I608244);
nor I_35569 (I608278,I608261,I119890);
nor I_35570 (I608295,I608193,I608278);
DFFARX1 I_35571 (I608295,I3563,I608159,I608145,);
not I_35572 (I608326,I119890);
nand I_35573 (I608343,I608326,I608261);
and I_35574 (I608360,I608326,I119893);
nand I_35575 (I608377,I608360,I119908);
nor I_35576 (I608142,I608377,I608326);
and I_35577 (I608133,I608219,I608377);
not I_35578 (I608422,I608377);
nand I_35579 (I608136,I608219,I608422);
nor I_35580 (I608130,I608185,I608377);
not I_35581 (I608467,I119899);
nor I_35582 (I608484,I608467,I119893);
nand I_35583 (I608501,I608484,I608326);
nor I_35584 (I608139,I608244,I608501);
nor I_35585 (I608532,I608467,I119887);
and I_35586 (I608549,I608532,I119896);
or I_35587 (I608566,I608549,I119905);
DFFARX1 I_35588 (I608566,I3563,I608159,I608592,);
nor I_35589 (I608600,I608592,I608343);
DFFARX1 I_35590 (I608600,I3563,I608159,I608127,);
DFFARX1 I_35591 (I608592,I3563,I608159,I608151,);
not I_35592 (I608645,I608592);
nor I_35593 (I608662,I608645,I608219);
nor I_35594 (I608679,I608484,I608662);
DFFARX1 I_35595 (I608679,I3563,I608159,I608148,);
not I_35596 (I608737,I3570);
DFFARX1 I_35597 (I386028,I3563,I608737,I608763,);
not I_35598 (I608771,I608763);
DFFARX1 I_35599 (I386043,I3563,I608737,I608797,);
not I_35600 (I608805,I386046);
nand I_35601 (I608822,I608805,I386025);
not I_35602 (I608839,I608822);
nor I_35603 (I608856,I608839,I386049);
nor I_35604 (I608873,I608771,I608856);
DFFARX1 I_35605 (I608873,I3563,I608737,I608723,);
not I_35606 (I608904,I386049);
nand I_35607 (I608921,I608904,I608839);
and I_35608 (I608938,I608904,I386031);
nand I_35609 (I608955,I608938,I386022);
nor I_35610 (I608720,I608955,I608904);
and I_35611 (I608711,I608797,I608955);
not I_35612 (I609000,I608955);
nand I_35613 (I608714,I608797,I609000);
nor I_35614 (I608708,I608763,I608955);
not I_35615 (I609045,I386022);
nor I_35616 (I609062,I609045,I386031);
nand I_35617 (I609079,I609062,I608904);
nor I_35618 (I608717,I608822,I609079);
nor I_35619 (I609110,I609045,I386037);
and I_35620 (I609127,I609110,I386040);
or I_35621 (I609144,I609127,I386034);
DFFARX1 I_35622 (I609144,I3563,I608737,I609170,);
nor I_35623 (I609178,I609170,I608921);
DFFARX1 I_35624 (I609178,I3563,I608737,I608705,);
DFFARX1 I_35625 (I609170,I3563,I608737,I608729,);
not I_35626 (I609223,I609170);
nor I_35627 (I609240,I609223,I608797);
nor I_35628 (I609257,I609062,I609240);
DFFARX1 I_35629 (I609257,I3563,I608737,I608726,);
not I_35630 (I609315,I3570);
DFFARX1 I_35631 (I451246,I3563,I609315,I609341,);
not I_35632 (I609349,I609341);
DFFARX1 I_35633 (I451258,I3563,I609315,I609375,);
not I_35634 (I609383,I451234);
nand I_35635 (I609400,I609383,I451261);
not I_35636 (I609417,I609400);
nor I_35637 (I609434,I609417,I451249);
nor I_35638 (I609451,I609349,I609434);
DFFARX1 I_35639 (I609451,I3563,I609315,I609301,);
not I_35640 (I609482,I451249);
nand I_35641 (I609499,I609482,I609417);
and I_35642 (I609516,I609482,I451234);
nand I_35643 (I609533,I609516,I451237);
nor I_35644 (I609298,I609533,I609482);
and I_35645 (I609289,I609375,I609533);
not I_35646 (I609578,I609533);
nand I_35647 (I609292,I609375,I609578);
nor I_35648 (I609286,I609341,I609533);
not I_35649 (I609623,I451243);
nor I_35650 (I609640,I609623,I451234);
nand I_35651 (I609657,I609640,I609482);
nor I_35652 (I609295,I609400,I609657);
nor I_35653 (I609688,I609623,I451252);
and I_35654 (I609705,I609688,I451240);
or I_35655 (I609722,I609705,I451255);
DFFARX1 I_35656 (I609722,I3563,I609315,I609748,);
nor I_35657 (I609756,I609748,I609499);
DFFARX1 I_35658 (I609756,I3563,I609315,I609283,);
DFFARX1 I_35659 (I609748,I3563,I609315,I609307,);
not I_35660 (I609801,I609748);
nor I_35661 (I609818,I609801,I609375);
nor I_35662 (I609835,I609640,I609818);
DFFARX1 I_35663 (I609835,I3563,I609315,I609304,);
not I_35664 (I609893,I3570);
DFFARX1 I_35665 (I494222,I3563,I609893,I609919,);
not I_35666 (I609927,I609919);
DFFARX1 I_35667 (I494234,I3563,I609893,I609953,);
not I_35668 (I609961,I494210);
nand I_35669 (I609978,I609961,I494237);
not I_35670 (I609995,I609978);
nor I_35671 (I610012,I609995,I494225);
nor I_35672 (I610029,I609927,I610012);
DFFARX1 I_35673 (I610029,I3563,I609893,I609879,);
not I_35674 (I610060,I494225);
nand I_35675 (I610077,I610060,I609995);
and I_35676 (I610094,I610060,I494210);
nand I_35677 (I610111,I610094,I494213);
nor I_35678 (I609876,I610111,I610060);
and I_35679 (I609867,I609953,I610111);
not I_35680 (I610156,I610111);
nand I_35681 (I609870,I609953,I610156);
nor I_35682 (I609864,I609919,I610111);
not I_35683 (I610201,I494219);
nor I_35684 (I610218,I610201,I494210);
nand I_35685 (I610235,I610218,I610060);
nor I_35686 (I609873,I609978,I610235);
nor I_35687 (I610266,I610201,I494228);
and I_35688 (I610283,I610266,I494216);
or I_35689 (I610300,I610283,I494231);
DFFARX1 I_35690 (I610300,I3563,I609893,I610326,);
nor I_35691 (I610334,I610326,I610077);
DFFARX1 I_35692 (I610334,I3563,I609893,I609861,);
DFFARX1 I_35693 (I610326,I3563,I609893,I609885,);
not I_35694 (I610379,I610326);
nor I_35695 (I610396,I610379,I609953);
nor I_35696 (I610413,I610218,I610396);
DFFARX1 I_35697 (I610413,I3563,I609893,I609882,);
not I_35698 (I610471,I3570);
DFFARX1 I_35699 (I948473,I3563,I610471,I610497,);
not I_35700 (I610505,I610497);
DFFARX1 I_35701 (I948470,I3563,I610471,I610531,);
not I_35702 (I610539,I948467);
nand I_35703 (I610556,I610539,I948494);
not I_35704 (I610573,I610556);
nor I_35705 (I610590,I610573,I948482);
nor I_35706 (I610607,I610505,I610590);
DFFARX1 I_35707 (I610607,I3563,I610471,I610457,);
not I_35708 (I610638,I948482);
nand I_35709 (I610655,I610638,I610573);
and I_35710 (I610672,I610638,I948488);
nand I_35711 (I610689,I610672,I948479);
nor I_35712 (I610454,I610689,I610638);
and I_35713 (I610445,I610531,I610689);
not I_35714 (I610734,I610689);
nand I_35715 (I610448,I610531,I610734);
nor I_35716 (I610442,I610497,I610689);
not I_35717 (I610779,I948476);
nor I_35718 (I610796,I610779,I948488);
nand I_35719 (I610813,I610796,I610638);
nor I_35720 (I610451,I610556,I610813);
nor I_35721 (I610844,I610779,I948491);
and I_35722 (I610861,I610844,I948485);
or I_35723 (I610878,I610861,I948467);
DFFARX1 I_35724 (I610878,I3563,I610471,I610904,);
nor I_35725 (I610912,I610904,I610655);
DFFARX1 I_35726 (I610912,I3563,I610471,I610439,);
DFFARX1 I_35727 (I610904,I3563,I610471,I610463,);
not I_35728 (I610957,I610904);
nor I_35729 (I610974,I610957,I610531);
nor I_35730 (I610991,I610796,I610974);
DFFARX1 I_35731 (I610991,I3563,I610471,I610460,);
not I_35732 (I611049,I3570);
DFFARX1 I_35733 (I1207751,I3563,I611049,I611075,);
not I_35734 (I611083,I611075);
DFFARX1 I_35735 (I1207757,I3563,I611049,I611109,);
not I_35736 (I611117,I1207751);
nand I_35737 (I611134,I611117,I1207754);
not I_35738 (I611151,I611134);
nor I_35739 (I611168,I611151,I1207772);
nor I_35740 (I611185,I611083,I611168);
DFFARX1 I_35741 (I611185,I3563,I611049,I611035,);
not I_35742 (I611216,I1207772);
nand I_35743 (I611233,I611216,I611151);
and I_35744 (I611250,I611216,I1207775);
nand I_35745 (I611267,I611250,I1207754);
nor I_35746 (I611032,I611267,I611216);
and I_35747 (I611023,I611109,I611267);
not I_35748 (I611312,I611267);
nand I_35749 (I611026,I611109,I611312);
nor I_35750 (I611020,I611075,I611267);
not I_35751 (I611357,I1207760);
nor I_35752 (I611374,I611357,I1207775);
nand I_35753 (I611391,I611374,I611216);
nor I_35754 (I611029,I611134,I611391);
nor I_35755 (I611422,I611357,I1207766);
and I_35756 (I611439,I611422,I1207763);
or I_35757 (I611456,I611439,I1207769);
DFFARX1 I_35758 (I611456,I3563,I611049,I611482,);
nor I_35759 (I611490,I611482,I611233);
DFFARX1 I_35760 (I611490,I3563,I611049,I611017,);
DFFARX1 I_35761 (I611482,I3563,I611049,I611041,);
not I_35762 (I611535,I611482);
nor I_35763 (I611552,I611535,I611109);
nor I_35764 (I611569,I611374,I611552);
DFFARX1 I_35765 (I611569,I3563,I611049,I611038,);
not I_35766 (I611627,I3570);
DFFARX1 I_35767 (I271423,I3563,I611627,I611653,);
not I_35768 (I611661,I611653);
DFFARX1 I_35769 (I271408,I3563,I611627,I611687,);
not I_35770 (I611695,I271426);
nand I_35771 (I611712,I611695,I271411);
not I_35772 (I611729,I611712);
nor I_35773 (I611746,I611729,I271408);
nor I_35774 (I611763,I611661,I611746);
DFFARX1 I_35775 (I611763,I3563,I611627,I611613,);
not I_35776 (I611794,I271408);
nand I_35777 (I611811,I611794,I611729);
and I_35778 (I611828,I611794,I271411);
nand I_35779 (I611845,I611828,I271432);
nor I_35780 (I611610,I611845,I611794);
and I_35781 (I611601,I611687,I611845);
not I_35782 (I611890,I611845);
nand I_35783 (I611604,I611687,I611890);
nor I_35784 (I611598,I611653,I611845);
not I_35785 (I611935,I271420);
nor I_35786 (I611952,I611935,I271411);
nand I_35787 (I611969,I611952,I611794);
nor I_35788 (I611607,I611712,I611969);
nor I_35789 (I612000,I611935,I271414);
and I_35790 (I612017,I612000,I271429);
or I_35791 (I612034,I612017,I271417);
DFFARX1 I_35792 (I612034,I3563,I611627,I612060,);
nor I_35793 (I612068,I612060,I611811);
DFFARX1 I_35794 (I612068,I3563,I611627,I611595,);
DFFARX1 I_35795 (I612060,I3563,I611627,I611619,);
not I_35796 (I612113,I612060);
nor I_35797 (I612130,I612113,I611687);
nor I_35798 (I612147,I611952,I612130);
DFFARX1 I_35799 (I612147,I3563,I611627,I611616,);
not I_35800 (I612205,I3570);
DFFARX1 I_35801 (I452878,I3563,I612205,I612231,);
not I_35802 (I612239,I612231);
DFFARX1 I_35803 (I452890,I3563,I612205,I612265,);
not I_35804 (I612273,I452866);
nand I_35805 (I612290,I612273,I452893);
not I_35806 (I612307,I612290);
nor I_35807 (I612324,I612307,I452881);
nor I_35808 (I612341,I612239,I612324);
DFFARX1 I_35809 (I612341,I3563,I612205,I612191,);
not I_35810 (I612372,I452881);
nand I_35811 (I612389,I612372,I612307);
and I_35812 (I612406,I612372,I452866);
nand I_35813 (I612423,I612406,I452869);
nor I_35814 (I612188,I612423,I612372);
and I_35815 (I612179,I612265,I612423);
not I_35816 (I612468,I612423);
nand I_35817 (I612182,I612265,I612468);
nor I_35818 (I612176,I612231,I612423);
not I_35819 (I612513,I452875);
nor I_35820 (I612530,I612513,I452866);
nand I_35821 (I612547,I612530,I612372);
nor I_35822 (I612185,I612290,I612547);
nor I_35823 (I612578,I612513,I452884);
and I_35824 (I612595,I612578,I452872);
or I_35825 (I612612,I612595,I452887);
DFFARX1 I_35826 (I612612,I3563,I612205,I612638,);
nor I_35827 (I612646,I612638,I612389);
DFFARX1 I_35828 (I612646,I3563,I612205,I612173,);
DFFARX1 I_35829 (I612638,I3563,I612205,I612197,);
not I_35830 (I612691,I612638);
nor I_35831 (I612708,I612691,I612265);
nor I_35832 (I612725,I612530,I612708);
DFFARX1 I_35833 (I612725,I3563,I612205,I612194,);
not I_35834 (I612783,I3570);
DFFARX1 I_35835 (I1354733,I3563,I612783,I612809,);
not I_35836 (I612817,I612809);
DFFARX1 I_35837 (I1354733,I3563,I612783,I612843,);
not I_35838 (I612851,I1354757);
nand I_35839 (I612868,I612851,I1354739);
not I_35840 (I612885,I612868);
nor I_35841 (I612902,I612885,I1354754);
nor I_35842 (I612919,I612817,I612902);
DFFARX1 I_35843 (I612919,I3563,I612783,I612769,);
not I_35844 (I612950,I1354754);
nand I_35845 (I612967,I612950,I612885);
and I_35846 (I612984,I612950,I1354736);
nand I_35847 (I613001,I612984,I1354745);
nor I_35848 (I612766,I613001,I612950);
and I_35849 (I612757,I612843,I613001);
not I_35850 (I613046,I613001);
nand I_35851 (I612760,I612843,I613046);
nor I_35852 (I612754,I612809,I613001);
not I_35853 (I613091,I1354742);
nor I_35854 (I613108,I613091,I1354736);
nand I_35855 (I613125,I613108,I612950);
nor I_35856 (I612763,I612868,I613125);
nor I_35857 (I613156,I613091,I1354751);
and I_35858 (I613173,I613156,I1354760);
or I_35859 (I613190,I613173,I1354748);
DFFARX1 I_35860 (I613190,I3563,I612783,I613216,);
nor I_35861 (I613224,I613216,I612967);
DFFARX1 I_35862 (I613224,I3563,I612783,I612751,);
DFFARX1 I_35863 (I613216,I3563,I612783,I612775,);
not I_35864 (I613269,I613216);
nor I_35865 (I613286,I613269,I612843);
nor I_35866 (I613303,I613108,I613286);
DFFARX1 I_35867 (I613303,I3563,I612783,I612772,);
not I_35868 (I613361,I3570);
DFFARX1 I_35869 (I820548,I3563,I613361,I613387,);
not I_35870 (I613395,I613387);
DFFARX1 I_35871 (I820548,I3563,I613361,I613421,);
not I_35872 (I613429,I820545);
nand I_35873 (I613446,I613429,I820560);
not I_35874 (I613463,I613446);
nor I_35875 (I613480,I613463,I820554);
nor I_35876 (I613497,I613395,I613480);
DFFARX1 I_35877 (I613497,I3563,I613361,I613347,);
not I_35878 (I613528,I820554);
nand I_35879 (I613545,I613528,I613463);
and I_35880 (I613562,I613528,I820551);
nand I_35881 (I613579,I613562,I820542);
nor I_35882 (I613344,I613579,I613528);
and I_35883 (I613335,I613421,I613579);
not I_35884 (I613624,I613579);
nand I_35885 (I613338,I613421,I613624);
nor I_35886 (I613332,I613387,I613579);
not I_35887 (I613669,I820563);
nor I_35888 (I613686,I613669,I820551);
nand I_35889 (I613703,I613686,I613528);
nor I_35890 (I613341,I613446,I613703);
nor I_35891 (I613734,I613669,I820542);
and I_35892 (I613751,I613734,I820545);
or I_35893 (I613768,I613751,I820557);
DFFARX1 I_35894 (I613768,I3563,I613361,I613794,);
nor I_35895 (I613802,I613794,I613545);
DFFARX1 I_35896 (I613802,I3563,I613361,I613329,);
DFFARX1 I_35897 (I613794,I3563,I613361,I613353,);
not I_35898 (I613847,I613794);
nor I_35899 (I613864,I613847,I613421);
nor I_35900 (I613881,I613686,I613864);
DFFARX1 I_35901 (I613881,I3563,I613361,I613350,);
not I_35902 (I613939,I3570);
DFFARX1 I_35903 (I747425,I3563,I613939,I613965,);
not I_35904 (I613973,I613965);
DFFARX1 I_35905 (I747437,I3563,I613939,I613999,);
not I_35906 (I614007,I747428);
nand I_35907 (I614024,I614007,I747431);
not I_35908 (I614041,I614024);
nor I_35909 (I614058,I614041,I747434);
nor I_35910 (I614075,I613973,I614058);
DFFARX1 I_35911 (I614075,I3563,I613939,I613925,);
not I_35912 (I614106,I747434);
nand I_35913 (I614123,I614106,I614041);
and I_35914 (I614140,I614106,I747428);
nand I_35915 (I614157,I614140,I747440);
nor I_35916 (I613922,I614157,I614106);
and I_35917 (I613913,I613999,I614157);
not I_35918 (I614202,I614157);
nand I_35919 (I613916,I613999,I614202);
nor I_35920 (I613910,I613965,I614157);
not I_35921 (I614247,I747446);
nor I_35922 (I614264,I614247,I747428);
nand I_35923 (I614281,I614264,I614106);
nor I_35924 (I613919,I614024,I614281);
nor I_35925 (I614312,I614247,I747425);
and I_35926 (I614329,I614312,I747443);
or I_35927 (I614346,I614329,I747449);
DFFARX1 I_35928 (I614346,I3563,I613939,I614372,);
nor I_35929 (I614380,I614372,I614123);
DFFARX1 I_35930 (I614380,I3563,I613939,I613907,);
DFFARX1 I_35931 (I614372,I3563,I613939,I613931,);
not I_35932 (I614425,I614372);
nor I_35933 (I614442,I614425,I613999);
nor I_35934 (I614459,I614264,I614442);
DFFARX1 I_35935 (I614459,I3563,I613939,I613928,);
not I_35936 (I614517,I3570);
DFFARX1 I_35937 (I1182319,I3563,I614517,I614543,);
not I_35938 (I614551,I614543);
DFFARX1 I_35939 (I1182325,I3563,I614517,I614577,);
not I_35940 (I614585,I1182319);
nand I_35941 (I614602,I614585,I1182322);
not I_35942 (I614619,I614602);
nor I_35943 (I614636,I614619,I1182340);
nor I_35944 (I614653,I614551,I614636);
DFFARX1 I_35945 (I614653,I3563,I614517,I614503,);
not I_35946 (I614684,I1182340);
nand I_35947 (I614701,I614684,I614619);
and I_35948 (I614718,I614684,I1182343);
nand I_35949 (I614735,I614718,I1182322);
nor I_35950 (I614500,I614735,I614684);
and I_35951 (I614491,I614577,I614735);
not I_35952 (I614780,I614735);
nand I_35953 (I614494,I614577,I614780);
nor I_35954 (I614488,I614543,I614735);
not I_35955 (I614825,I1182328);
nor I_35956 (I614842,I614825,I1182343);
nand I_35957 (I614859,I614842,I614684);
nor I_35958 (I614497,I614602,I614859);
nor I_35959 (I614890,I614825,I1182334);
and I_35960 (I614907,I614890,I1182331);
or I_35961 (I614924,I614907,I1182337);
DFFARX1 I_35962 (I614924,I3563,I614517,I614950,);
nor I_35963 (I614958,I614950,I614701);
DFFARX1 I_35964 (I614958,I3563,I614517,I614485,);
DFFARX1 I_35965 (I614950,I3563,I614517,I614509,);
not I_35966 (I615003,I614950);
nor I_35967 (I615020,I615003,I614577);
nor I_35968 (I615037,I614842,I615020);
DFFARX1 I_35969 (I615037,I3563,I614517,I614506,);
not I_35970 (I615095,I3570);
DFFARX1 I_35971 (I1132611,I3563,I615095,I615121,);
not I_35972 (I615129,I615121);
DFFARX1 I_35973 (I1132617,I3563,I615095,I615155,);
not I_35974 (I615163,I1132611);
nand I_35975 (I615180,I615163,I1132614);
not I_35976 (I615197,I615180);
nor I_35977 (I615214,I615197,I1132632);
nor I_35978 (I615231,I615129,I615214);
DFFARX1 I_35979 (I615231,I3563,I615095,I615081,);
not I_35980 (I615262,I1132632);
nand I_35981 (I615279,I615262,I615197);
and I_35982 (I615296,I615262,I1132635);
nand I_35983 (I615313,I615296,I1132614);
nor I_35984 (I615078,I615313,I615262);
and I_35985 (I615069,I615155,I615313);
not I_35986 (I615358,I615313);
nand I_35987 (I615072,I615155,I615358);
nor I_35988 (I615066,I615121,I615313);
not I_35989 (I615403,I1132620);
nor I_35990 (I615420,I615403,I1132635);
nand I_35991 (I615437,I615420,I615262);
nor I_35992 (I615075,I615180,I615437);
nor I_35993 (I615468,I615403,I1132626);
and I_35994 (I615485,I615468,I1132623);
or I_35995 (I615502,I615485,I1132629);
DFFARX1 I_35996 (I615502,I3563,I615095,I615528,);
nor I_35997 (I615536,I615528,I615279);
DFFARX1 I_35998 (I615536,I3563,I615095,I615063,);
DFFARX1 I_35999 (I615528,I3563,I615095,I615087,);
not I_36000 (I615581,I615528);
nor I_36001 (I615598,I615581,I615155);
nor I_36002 (I615615,I615420,I615598);
DFFARX1 I_36003 (I615615,I3563,I615095,I615084,);
not I_36004 (I615673,I3570);
DFFARX1 I_36005 (I1164401,I3563,I615673,I615699,);
not I_36006 (I615707,I615699);
DFFARX1 I_36007 (I1164407,I3563,I615673,I615733,);
not I_36008 (I615741,I1164401);
nand I_36009 (I615758,I615741,I1164404);
not I_36010 (I615775,I615758);
nor I_36011 (I615792,I615775,I1164422);
nor I_36012 (I615809,I615707,I615792);
DFFARX1 I_36013 (I615809,I3563,I615673,I615659,);
not I_36014 (I615840,I1164422);
nand I_36015 (I615857,I615840,I615775);
and I_36016 (I615874,I615840,I1164425);
nand I_36017 (I615891,I615874,I1164404);
nor I_36018 (I615656,I615891,I615840);
and I_36019 (I615647,I615733,I615891);
not I_36020 (I615936,I615891);
nand I_36021 (I615650,I615733,I615936);
nor I_36022 (I615644,I615699,I615891);
not I_36023 (I615981,I1164410);
nor I_36024 (I615998,I615981,I1164425);
nand I_36025 (I616015,I615998,I615840);
nor I_36026 (I615653,I615758,I616015);
nor I_36027 (I616046,I615981,I1164416);
and I_36028 (I616063,I616046,I1164413);
or I_36029 (I616080,I616063,I1164419);
DFFARX1 I_36030 (I616080,I3563,I615673,I616106,);
nor I_36031 (I616114,I616106,I615857);
DFFARX1 I_36032 (I616114,I3563,I615673,I615641,);
DFFARX1 I_36033 (I616106,I3563,I615673,I615665,);
not I_36034 (I616159,I616106);
nor I_36035 (I616176,I616159,I615733);
nor I_36036 (I616193,I615998,I616176);
DFFARX1 I_36037 (I616193,I3563,I615673,I615662,);
not I_36038 (I616251,I3570);
DFFARX1 I_36039 (I413959,I3563,I616251,I616277,);
not I_36040 (I616285,I616277);
DFFARX1 I_36041 (I413974,I3563,I616251,I616311,);
not I_36042 (I616319,I413977);
nand I_36043 (I616336,I616319,I413956);
not I_36044 (I616353,I616336);
nor I_36045 (I616370,I616353,I413980);
nor I_36046 (I616387,I616285,I616370);
DFFARX1 I_36047 (I616387,I3563,I616251,I616237,);
not I_36048 (I616418,I413980);
nand I_36049 (I616435,I616418,I616353);
and I_36050 (I616452,I616418,I413962);
nand I_36051 (I616469,I616452,I413953);
nor I_36052 (I616234,I616469,I616418);
and I_36053 (I616225,I616311,I616469);
not I_36054 (I616514,I616469);
nand I_36055 (I616228,I616311,I616514);
nor I_36056 (I616222,I616277,I616469);
not I_36057 (I616559,I413953);
nor I_36058 (I616576,I616559,I413962);
nand I_36059 (I616593,I616576,I616418);
nor I_36060 (I616231,I616336,I616593);
nor I_36061 (I616624,I616559,I413968);
and I_36062 (I616641,I616624,I413971);
or I_36063 (I616658,I616641,I413965);
DFFARX1 I_36064 (I616658,I3563,I616251,I616684,);
nor I_36065 (I616692,I616684,I616435);
DFFARX1 I_36066 (I616692,I3563,I616251,I616219,);
DFFARX1 I_36067 (I616684,I3563,I616251,I616243,);
not I_36068 (I616737,I616684);
nor I_36069 (I616754,I616737,I616311);
nor I_36070 (I616771,I616576,I616754);
DFFARX1 I_36071 (I616771,I3563,I616251,I616240,);
not I_36072 (I616829,I3570);
DFFARX1 I_36073 (I817386,I3563,I616829,I616855,);
not I_36074 (I616863,I616855);
DFFARX1 I_36075 (I817386,I3563,I616829,I616889,);
not I_36076 (I616897,I817383);
nand I_36077 (I616914,I616897,I817398);
not I_36078 (I616931,I616914);
nor I_36079 (I616948,I616931,I817392);
nor I_36080 (I616965,I616863,I616948);
DFFARX1 I_36081 (I616965,I3563,I616829,I616815,);
not I_36082 (I616996,I817392);
nand I_36083 (I617013,I616996,I616931);
and I_36084 (I617030,I616996,I817389);
nand I_36085 (I617047,I617030,I817380);
nor I_36086 (I616812,I617047,I616996);
and I_36087 (I616803,I616889,I617047);
not I_36088 (I617092,I617047);
nand I_36089 (I616806,I616889,I617092);
nor I_36090 (I616800,I616855,I617047);
not I_36091 (I617137,I817401);
nor I_36092 (I617154,I617137,I817389);
nand I_36093 (I617171,I617154,I616996);
nor I_36094 (I616809,I616914,I617171);
nor I_36095 (I617202,I617137,I817380);
and I_36096 (I617219,I617202,I817383);
or I_36097 (I617236,I617219,I817395);
DFFARX1 I_36098 (I617236,I3563,I616829,I617262,);
nor I_36099 (I617270,I617262,I617013);
DFFARX1 I_36100 (I617270,I3563,I616829,I616797,);
DFFARX1 I_36101 (I617262,I3563,I616829,I616821,);
not I_36102 (I617315,I617262);
nor I_36103 (I617332,I617315,I616889);
nor I_36104 (I617349,I617154,I617332);
DFFARX1 I_36105 (I617349,I3563,I616829,I616818,);
not I_36106 (I617407,I3570);
DFFARX1 I_36107 (I841101,I3563,I617407,I617433,);
not I_36108 (I617441,I617433);
DFFARX1 I_36109 (I841101,I3563,I617407,I617467,);
not I_36110 (I617475,I841098);
nand I_36111 (I617492,I617475,I841113);
not I_36112 (I617509,I617492);
nor I_36113 (I617526,I617509,I841107);
nor I_36114 (I617543,I617441,I617526);
DFFARX1 I_36115 (I617543,I3563,I617407,I617393,);
not I_36116 (I617574,I841107);
nand I_36117 (I617591,I617574,I617509);
and I_36118 (I617608,I617574,I841104);
nand I_36119 (I617625,I617608,I841095);
nor I_36120 (I617390,I617625,I617574);
and I_36121 (I617381,I617467,I617625);
not I_36122 (I617670,I617625);
nand I_36123 (I617384,I617467,I617670);
nor I_36124 (I617378,I617433,I617625);
not I_36125 (I617715,I841116);
nor I_36126 (I617732,I617715,I841104);
nand I_36127 (I617749,I617732,I617574);
nor I_36128 (I617387,I617492,I617749);
nor I_36129 (I617780,I617715,I841095);
and I_36130 (I617797,I617780,I841098);
or I_36131 (I617814,I617797,I841110);
DFFARX1 I_36132 (I617814,I3563,I617407,I617840,);
nor I_36133 (I617848,I617840,I617591);
DFFARX1 I_36134 (I617848,I3563,I617407,I617375,);
DFFARX1 I_36135 (I617840,I3563,I617407,I617399,);
not I_36136 (I617893,I617840);
nor I_36137 (I617910,I617893,I617467);
nor I_36138 (I617927,I617732,I617910);
DFFARX1 I_36139 (I617927,I3563,I617407,I617396,);
not I_36140 (I617985,I3570);
DFFARX1 I_36141 (I1151685,I3563,I617985,I618011,);
not I_36142 (I618019,I618011);
DFFARX1 I_36143 (I1151691,I3563,I617985,I618045,);
not I_36144 (I618053,I1151685);
nand I_36145 (I618070,I618053,I1151688);
not I_36146 (I618087,I618070);
nor I_36147 (I618104,I618087,I1151706);
nor I_36148 (I618121,I618019,I618104);
DFFARX1 I_36149 (I618121,I3563,I617985,I617971,);
not I_36150 (I618152,I1151706);
nand I_36151 (I618169,I618152,I618087);
and I_36152 (I618186,I618152,I1151709);
nand I_36153 (I618203,I618186,I1151688);
nor I_36154 (I617968,I618203,I618152);
and I_36155 (I617959,I618045,I618203);
not I_36156 (I618248,I618203);
nand I_36157 (I617962,I618045,I618248);
nor I_36158 (I617956,I618011,I618203);
not I_36159 (I618293,I1151694);
nor I_36160 (I618310,I618293,I1151709);
nand I_36161 (I618327,I618310,I618152);
nor I_36162 (I617965,I618070,I618327);
nor I_36163 (I618358,I618293,I1151700);
and I_36164 (I618375,I618358,I1151697);
or I_36165 (I618392,I618375,I1151703);
DFFARX1 I_36166 (I618392,I3563,I617985,I618418,);
nor I_36167 (I618426,I618418,I618169);
DFFARX1 I_36168 (I618426,I3563,I617985,I617953,);
DFFARX1 I_36169 (I618418,I3563,I617985,I617977,);
not I_36170 (I618471,I618418);
nor I_36171 (I618488,I618471,I618045);
nor I_36172 (I618505,I618310,I618488);
DFFARX1 I_36173 (I618505,I3563,I617985,I617974,);
not I_36174 (I618563,I3570);
DFFARX1 I_36175 (I175628,I3563,I618563,I618589,);
not I_36176 (I618597,I618589);
DFFARX1 I_36177 (I175613,I3563,I618563,I618623,);
not I_36178 (I618631,I175631);
nand I_36179 (I618648,I618631,I175616);
not I_36180 (I618665,I618648);
nor I_36181 (I618682,I618665,I175613);
nor I_36182 (I618699,I618597,I618682);
DFFARX1 I_36183 (I618699,I3563,I618563,I618549,);
not I_36184 (I618730,I175613);
nand I_36185 (I618747,I618730,I618665);
and I_36186 (I618764,I618730,I175616);
nand I_36187 (I618781,I618764,I175637);
nor I_36188 (I618546,I618781,I618730);
and I_36189 (I618537,I618623,I618781);
not I_36190 (I618826,I618781);
nand I_36191 (I618540,I618623,I618826);
nor I_36192 (I618534,I618589,I618781);
not I_36193 (I618871,I175625);
nor I_36194 (I618888,I618871,I175616);
nand I_36195 (I618905,I618888,I618730);
nor I_36196 (I618543,I618648,I618905);
nor I_36197 (I618936,I618871,I175619);
and I_36198 (I618953,I618936,I175634);
or I_36199 (I618970,I618953,I175622);
DFFARX1 I_36200 (I618970,I3563,I618563,I618996,);
nor I_36201 (I619004,I618996,I618747);
DFFARX1 I_36202 (I619004,I3563,I618563,I618531,);
DFFARX1 I_36203 (I618996,I3563,I618563,I618555,);
not I_36204 (I619049,I618996);
nor I_36205 (I619066,I619049,I618623);
nor I_36206 (I619083,I618888,I619066);
DFFARX1 I_36207 (I619083,I3563,I618563,I618552,);
not I_36208 (I619141,I3570);
DFFARX1 I_36209 (I975605,I3563,I619141,I619167,);
not I_36210 (I619175,I619167);
DFFARX1 I_36211 (I975602,I3563,I619141,I619201,);
not I_36212 (I619209,I975599);
nand I_36213 (I619226,I619209,I975626);
not I_36214 (I619243,I619226);
nor I_36215 (I619260,I619243,I975614);
nor I_36216 (I619277,I619175,I619260);
DFFARX1 I_36217 (I619277,I3563,I619141,I619127,);
not I_36218 (I619308,I975614);
nand I_36219 (I619325,I619308,I619243);
and I_36220 (I619342,I619308,I975620);
nand I_36221 (I619359,I619342,I975611);
nor I_36222 (I619124,I619359,I619308);
and I_36223 (I619115,I619201,I619359);
not I_36224 (I619404,I619359);
nand I_36225 (I619118,I619201,I619404);
nor I_36226 (I619112,I619167,I619359);
not I_36227 (I619449,I975608);
nor I_36228 (I619466,I619449,I975620);
nand I_36229 (I619483,I619466,I619308);
nor I_36230 (I619121,I619226,I619483);
nor I_36231 (I619514,I619449,I975623);
and I_36232 (I619531,I619514,I975617);
or I_36233 (I619548,I619531,I975599);
DFFARX1 I_36234 (I619548,I3563,I619141,I619574,);
nor I_36235 (I619582,I619574,I619325);
DFFARX1 I_36236 (I619582,I3563,I619141,I619109,);
DFFARX1 I_36237 (I619574,I3563,I619141,I619133,);
not I_36238 (I619627,I619574);
nor I_36239 (I619644,I619627,I619201);
nor I_36240 (I619661,I619466,I619644);
DFFARX1 I_36241 (I619661,I3563,I619141,I619130,);
not I_36242 (I619719,I3570);
DFFARX1 I_36243 (I65630,I3563,I619719,I619745,);
not I_36244 (I619753,I619745);
DFFARX1 I_36245 (I65609,I3563,I619719,I619779,);
not I_36246 (I619787,I65606);
nand I_36247 (I619804,I619787,I65621);
not I_36248 (I619821,I619804);
nor I_36249 (I619838,I619821,I65609);
nor I_36250 (I619855,I619753,I619838);
DFFARX1 I_36251 (I619855,I3563,I619719,I619705,);
not I_36252 (I619886,I65609);
nand I_36253 (I619903,I619886,I619821);
and I_36254 (I619920,I619886,I65612);
nand I_36255 (I619937,I619920,I65627);
nor I_36256 (I619702,I619937,I619886);
and I_36257 (I619693,I619779,I619937);
not I_36258 (I619982,I619937);
nand I_36259 (I619696,I619779,I619982);
nor I_36260 (I619690,I619745,I619937);
not I_36261 (I620027,I65618);
nor I_36262 (I620044,I620027,I65612);
nand I_36263 (I620061,I620044,I619886);
nor I_36264 (I619699,I619804,I620061);
nor I_36265 (I620092,I620027,I65606);
and I_36266 (I620109,I620092,I65615);
or I_36267 (I620126,I620109,I65624);
DFFARX1 I_36268 (I620126,I3563,I619719,I620152,);
nor I_36269 (I620160,I620152,I619903);
DFFARX1 I_36270 (I620160,I3563,I619719,I619687,);
DFFARX1 I_36271 (I620152,I3563,I619719,I619711,);
not I_36272 (I620205,I620152);
nor I_36273 (I620222,I620205,I619779);
nor I_36274 (I620239,I620044,I620222);
DFFARX1 I_36275 (I620239,I3563,I619719,I619708,);
not I_36276 (I620297,I3570);
DFFARX1 I_36277 (I1940,I3563,I620297,I620323,);
not I_36278 (I620331,I620323);
DFFARX1 I_36279 (I2716,I3563,I620297,I620357,);
not I_36280 (I620365,I2028);
nand I_36281 (I620382,I620365,I1708);
not I_36282 (I620399,I620382);
nor I_36283 (I620416,I620399,I1476);
nor I_36284 (I620433,I620331,I620416);
DFFARX1 I_36285 (I620433,I3563,I620297,I620283,);
not I_36286 (I620464,I1476);
nand I_36287 (I620481,I620464,I620399);
and I_36288 (I620498,I620464,I2188);
nand I_36289 (I620515,I620498,I3436);
nor I_36290 (I620280,I620515,I620464);
and I_36291 (I620271,I620357,I620515);
not I_36292 (I620560,I620515);
nand I_36293 (I620274,I620357,I620560);
nor I_36294 (I620268,I620323,I620515);
not I_36295 (I620605,I1924);
nor I_36296 (I620622,I620605,I2188);
nand I_36297 (I620639,I620622,I620464);
nor I_36298 (I620277,I620382,I620639);
nor I_36299 (I620670,I620605,I3228);
and I_36300 (I620687,I620670,I2868);
or I_36301 (I620704,I620687,I2692);
DFFARX1 I_36302 (I620704,I3563,I620297,I620730,);
nor I_36303 (I620738,I620730,I620481);
DFFARX1 I_36304 (I620738,I3563,I620297,I620265,);
DFFARX1 I_36305 (I620730,I3563,I620297,I620289,);
not I_36306 (I620783,I620730);
nor I_36307 (I620800,I620783,I620357);
nor I_36308 (I620817,I620622,I620800);
DFFARX1 I_36309 (I620817,I3563,I620297,I620286,);
not I_36310 (I620875,I3570);
DFFARX1 I_36311 (I88291,I3563,I620875,I620901,);
not I_36312 (I620909,I620901);
DFFARX1 I_36313 (I88270,I3563,I620875,I620935,);
not I_36314 (I620943,I88267);
nand I_36315 (I620960,I620943,I88282);
not I_36316 (I620977,I620960);
nor I_36317 (I620994,I620977,I88270);
nor I_36318 (I621011,I620909,I620994);
DFFARX1 I_36319 (I621011,I3563,I620875,I620861,);
not I_36320 (I621042,I88270);
nand I_36321 (I621059,I621042,I620977);
and I_36322 (I621076,I621042,I88273);
nand I_36323 (I621093,I621076,I88288);
nor I_36324 (I620858,I621093,I621042);
and I_36325 (I620849,I620935,I621093);
not I_36326 (I621138,I621093);
nand I_36327 (I620852,I620935,I621138);
nor I_36328 (I620846,I620901,I621093);
not I_36329 (I621183,I88279);
nor I_36330 (I621200,I621183,I88273);
nand I_36331 (I621217,I621200,I621042);
nor I_36332 (I620855,I620960,I621217);
nor I_36333 (I621248,I621183,I88267);
and I_36334 (I621265,I621248,I88276);
or I_36335 (I621282,I621265,I88285);
DFFARX1 I_36336 (I621282,I3563,I620875,I621308,);
nor I_36337 (I621316,I621308,I621059);
DFFARX1 I_36338 (I621316,I3563,I620875,I620843,);
DFFARX1 I_36339 (I621308,I3563,I620875,I620867,);
not I_36340 (I621361,I621308);
nor I_36341 (I621378,I621361,I620935);
nor I_36342 (I621395,I621200,I621378);
DFFARX1 I_36343 (I621395,I3563,I620875,I620864,);
not I_36344 (I621453,I3570);
DFFARX1 I_36345 (I83548,I3563,I621453,I621479,);
not I_36346 (I621487,I621479);
DFFARX1 I_36347 (I83527,I3563,I621453,I621513,);
not I_36348 (I621521,I83524);
nand I_36349 (I621538,I621521,I83539);
not I_36350 (I621555,I621538);
nor I_36351 (I621572,I621555,I83527);
nor I_36352 (I621589,I621487,I621572);
DFFARX1 I_36353 (I621589,I3563,I621453,I621439,);
not I_36354 (I621620,I83527);
nand I_36355 (I621637,I621620,I621555);
and I_36356 (I621654,I621620,I83530);
nand I_36357 (I621671,I621654,I83545);
nor I_36358 (I621436,I621671,I621620);
and I_36359 (I621427,I621513,I621671);
not I_36360 (I621716,I621671);
nand I_36361 (I621430,I621513,I621716);
nor I_36362 (I621424,I621479,I621671);
not I_36363 (I621761,I83536);
nor I_36364 (I621778,I621761,I83530);
nand I_36365 (I621795,I621778,I621620);
nor I_36366 (I621433,I621538,I621795);
nor I_36367 (I621826,I621761,I83524);
and I_36368 (I621843,I621826,I83533);
or I_36369 (I621860,I621843,I83542);
DFFARX1 I_36370 (I621860,I3563,I621453,I621886,);
nor I_36371 (I621894,I621886,I621637);
DFFARX1 I_36372 (I621894,I3563,I621453,I621421,);
DFFARX1 I_36373 (I621886,I3563,I621453,I621445,);
not I_36374 (I621939,I621886);
nor I_36375 (I621956,I621939,I621513);
nor I_36376 (I621973,I621778,I621956);
DFFARX1 I_36377 (I621973,I3563,I621453,I621442,);
not I_36378 (I622031,I3570);
DFFARX1 I_36379 (I1088755,I3563,I622031,I622057,);
not I_36380 (I622065,I622057);
DFFARX1 I_36381 (I1088746,I3563,I622031,I622091,);
not I_36382 (I622099,I1088740);
nand I_36383 (I622116,I622099,I1088752);
not I_36384 (I622133,I622116);
nor I_36385 (I622150,I622133,I1088743);
nor I_36386 (I622167,I622065,I622150);
DFFARX1 I_36387 (I622167,I3563,I622031,I622017,);
not I_36388 (I622198,I1088743);
nand I_36389 (I622215,I622198,I622133);
and I_36390 (I622232,I622198,I1088749);
nand I_36391 (I622249,I622232,I1088734);
nor I_36392 (I622014,I622249,I622198);
and I_36393 (I622005,I622091,I622249);
not I_36394 (I622294,I622249);
nand I_36395 (I622008,I622091,I622294);
nor I_36396 (I622002,I622057,I622249);
not I_36397 (I622339,I1088734);
nor I_36398 (I622356,I622339,I1088749);
nand I_36399 (I622373,I622356,I622198);
nor I_36400 (I622011,I622116,I622373);
nor I_36401 (I622404,I622339,I1088737);
and I_36402 (I622421,I622404,I1088740);
or I_36403 (I622438,I622421,I1088737);
DFFARX1 I_36404 (I622438,I3563,I622031,I622464,);
nor I_36405 (I622472,I622464,I622215);
DFFARX1 I_36406 (I622472,I3563,I622031,I621999,);
DFFARX1 I_36407 (I622464,I3563,I622031,I622023,);
not I_36408 (I622517,I622464);
nor I_36409 (I622534,I622517,I622091);
nor I_36410 (I622551,I622356,I622534);
DFFARX1 I_36411 (I622551,I3563,I622031,I622020,);
not I_36412 (I622609,I3570);
DFFARX1 I_36413 (I1397573,I3563,I622609,I622635,);
not I_36414 (I622643,I622635);
DFFARX1 I_36415 (I1397573,I3563,I622609,I622669,);
not I_36416 (I622677,I1397597);
nand I_36417 (I622694,I622677,I1397579);
not I_36418 (I622711,I622694);
nor I_36419 (I622728,I622711,I1397594);
nor I_36420 (I622745,I622643,I622728);
DFFARX1 I_36421 (I622745,I3563,I622609,I622595,);
not I_36422 (I622776,I1397594);
nand I_36423 (I622793,I622776,I622711);
and I_36424 (I622810,I622776,I1397576);
nand I_36425 (I622827,I622810,I1397585);
nor I_36426 (I622592,I622827,I622776);
and I_36427 (I622583,I622669,I622827);
not I_36428 (I622872,I622827);
nand I_36429 (I622586,I622669,I622872);
nor I_36430 (I622580,I622635,I622827);
not I_36431 (I622917,I1397582);
nor I_36432 (I622934,I622917,I1397576);
nand I_36433 (I622951,I622934,I622776);
nor I_36434 (I622589,I622694,I622951);
nor I_36435 (I622982,I622917,I1397591);
and I_36436 (I622999,I622982,I1397600);
or I_36437 (I623016,I622999,I1397588);
DFFARX1 I_36438 (I623016,I3563,I622609,I623042,);
nor I_36439 (I623050,I623042,I622793);
DFFARX1 I_36440 (I623050,I3563,I622609,I622577,);
DFFARX1 I_36441 (I623042,I3563,I622609,I622601,);
not I_36442 (I623095,I623042);
nor I_36443 (I623112,I623095,I622669);
nor I_36444 (I623129,I622934,I623112);
DFFARX1 I_36445 (I623129,I3563,I622609,I622598,);
not I_36446 (I623187,I3570);
DFFARX1 I_36447 (I506734,I3563,I623187,I623213,);
not I_36448 (I623221,I623213);
DFFARX1 I_36449 (I506746,I3563,I623187,I623247,);
not I_36450 (I623255,I506722);
nand I_36451 (I623272,I623255,I506749);
not I_36452 (I623289,I623272);
nor I_36453 (I623306,I623289,I506737);
nor I_36454 (I623323,I623221,I623306);
DFFARX1 I_36455 (I623323,I3563,I623187,I623173,);
not I_36456 (I623354,I506737);
nand I_36457 (I623371,I623354,I623289);
and I_36458 (I623388,I623354,I506722);
nand I_36459 (I623405,I623388,I506725);
nor I_36460 (I623170,I623405,I623354);
and I_36461 (I623161,I623247,I623405);
not I_36462 (I623450,I623405);
nand I_36463 (I623164,I623247,I623450);
nor I_36464 (I623158,I623213,I623405);
not I_36465 (I623495,I506731);
nor I_36466 (I623512,I623495,I506722);
nand I_36467 (I623529,I623512,I623354);
nor I_36468 (I623167,I623272,I623529);
nor I_36469 (I623560,I623495,I506740);
and I_36470 (I623577,I623560,I506728);
or I_36471 (I623594,I623577,I506743);
DFFARX1 I_36472 (I623594,I3563,I623187,I623620,);
nor I_36473 (I623628,I623620,I623371);
DFFARX1 I_36474 (I623628,I3563,I623187,I623155,);
DFFARX1 I_36475 (I623620,I3563,I623187,I623179,);
not I_36476 (I623673,I623620);
nor I_36477 (I623690,I623673,I623247);
nor I_36478 (I623707,I623512,I623690);
DFFARX1 I_36479 (I623707,I3563,I623187,I623176,);
not I_36480 (I623765,I3570);
DFFARX1 I_36481 (I161354,I3563,I623765,I623791,);
not I_36482 (I623799,I623791);
DFFARX1 I_36483 (I161333,I3563,I623765,I623825,);
not I_36484 (I623833,I161333);
nand I_36485 (I623850,I623833,I161360);
not I_36486 (I623867,I623850);
nor I_36487 (I623884,I623867,I161336);
nor I_36488 (I623901,I623799,I623884);
DFFARX1 I_36489 (I623901,I3563,I623765,I623751,);
not I_36490 (I623932,I161336);
nand I_36491 (I623949,I623932,I623867);
and I_36492 (I623966,I623932,I161357);
nand I_36493 (I623983,I623966,I161339);
nor I_36494 (I623748,I623983,I623932);
and I_36495 (I623739,I623825,I623983);
not I_36496 (I624028,I623983);
nand I_36497 (I623742,I623825,I624028);
nor I_36498 (I623736,I623791,I623983);
not I_36499 (I624073,I161342);
nor I_36500 (I624090,I624073,I161357);
nand I_36501 (I624107,I624090,I623932);
nor I_36502 (I623745,I623850,I624107);
nor I_36503 (I624138,I624073,I161348);
and I_36504 (I624155,I624138,I161345);
or I_36505 (I624172,I624155,I161351);
DFFARX1 I_36506 (I624172,I3563,I623765,I624198,);
nor I_36507 (I624206,I624198,I623949);
DFFARX1 I_36508 (I624206,I3563,I623765,I623733,);
DFFARX1 I_36509 (I624198,I3563,I623765,I623757,);
not I_36510 (I624251,I624198);
nor I_36511 (I624268,I624251,I623825);
nor I_36512 (I624285,I624090,I624268);
DFFARX1 I_36513 (I624285,I3563,I623765,I623754,);
not I_36514 (I624343,I3570);
DFFARX1 I_36515 (I1047241,I3563,I624343,I624369,);
not I_36516 (I624377,I624369);
DFFARX1 I_36517 (I1047232,I3563,I624343,I624403,);
not I_36518 (I624411,I1047226);
nand I_36519 (I624428,I624411,I1047238);
not I_36520 (I624445,I624428);
nor I_36521 (I624462,I624445,I1047229);
nor I_36522 (I624479,I624377,I624462);
DFFARX1 I_36523 (I624479,I3563,I624343,I624329,);
not I_36524 (I624510,I1047229);
nand I_36525 (I624527,I624510,I624445);
and I_36526 (I624544,I624510,I1047235);
nand I_36527 (I624561,I624544,I1047220);
nor I_36528 (I624326,I624561,I624510);
and I_36529 (I624317,I624403,I624561);
not I_36530 (I624606,I624561);
nand I_36531 (I624320,I624403,I624606);
nor I_36532 (I624314,I624369,I624561);
not I_36533 (I624651,I1047220);
nor I_36534 (I624668,I624651,I1047235);
nand I_36535 (I624685,I624668,I624510);
nor I_36536 (I624323,I624428,I624685);
nor I_36537 (I624716,I624651,I1047223);
and I_36538 (I624733,I624716,I1047226);
or I_36539 (I624750,I624733,I1047223);
DFFARX1 I_36540 (I624750,I3563,I624343,I624776,);
nor I_36541 (I624784,I624776,I624527);
DFFARX1 I_36542 (I624784,I3563,I624343,I624311,);
DFFARX1 I_36543 (I624776,I3563,I624343,I624335,);
not I_36544 (I624829,I624776);
nor I_36545 (I624846,I624829,I624403);
nor I_36546 (I624863,I624668,I624846);
DFFARX1 I_36547 (I624863,I3563,I624343,I624332,);
not I_36548 (I624921,I3570);
DFFARX1 I_36549 (I1297591,I3563,I624921,I624947,);
not I_36550 (I624955,I624947);
DFFARX1 I_36551 (I1297603,I3563,I624921,I624981,);
not I_36552 (I624989,I1297594);
nand I_36553 (I625006,I624989,I1297582);
not I_36554 (I625023,I625006);
nor I_36555 (I625040,I625023,I1297579);
nor I_36556 (I625057,I624955,I625040);
DFFARX1 I_36557 (I625057,I3563,I624921,I624907,);
not I_36558 (I625088,I1297579);
nand I_36559 (I625105,I625088,I625023);
and I_36560 (I625122,I625088,I1297585);
nand I_36561 (I625139,I625122,I1297582);
nor I_36562 (I624904,I625139,I625088);
and I_36563 (I624895,I624981,I625139);
not I_36564 (I625184,I625139);
nand I_36565 (I624898,I624981,I625184);
nor I_36566 (I624892,I624947,I625139);
not I_36567 (I625229,I1297600);
nor I_36568 (I625246,I625229,I1297585);
nand I_36569 (I625263,I625246,I625088);
nor I_36570 (I624901,I625006,I625263);
nor I_36571 (I625294,I625229,I1297588);
and I_36572 (I625311,I625294,I1297579);
or I_36573 (I625328,I625311,I1297597);
DFFARX1 I_36574 (I625328,I3563,I624921,I625354,);
nor I_36575 (I625362,I625354,I625105);
DFFARX1 I_36576 (I625362,I3563,I624921,I624889,);
DFFARX1 I_36577 (I625354,I3563,I624921,I624913,);
not I_36578 (I625407,I625354);
nor I_36579 (I625424,I625407,I624981);
nor I_36580 (I625441,I625246,I625424);
DFFARX1 I_36581 (I625441,I3563,I624921,I624910,);
not I_36582 (I625499,I3570);
DFFARX1 I_36583 (I1299903,I3563,I625499,I625525,);
not I_36584 (I625533,I625525);
DFFARX1 I_36585 (I1299915,I3563,I625499,I625559,);
not I_36586 (I625567,I1299906);
nand I_36587 (I625584,I625567,I1299894);
not I_36588 (I625601,I625584);
nor I_36589 (I625618,I625601,I1299891);
nor I_36590 (I625635,I625533,I625618);
DFFARX1 I_36591 (I625635,I3563,I625499,I625485,);
not I_36592 (I625666,I1299891);
nand I_36593 (I625683,I625666,I625601);
and I_36594 (I625700,I625666,I1299897);
nand I_36595 (I625717,I625700,I1299894);
nor I_36596 (I625482,I625717,I625666);
and I_36597 (I625473,I625559,I625717);
not I_36598 (I625762,I625717);
nand I_36599 (I625476,I625559,I625762);
nor I_36600 (I625470,I625525,I625717);
not I_36601 (I625807,I1299912);
nor I_36602 (I625824,I625807,I1299897);
nand I_36603 (I625841,I625824,I625666);
nor I_36604 (I625479,I625584,I625841);
nor I_36605 (I625872,I625807,I1299900);
and I_36606 (I625889,I625872,I1299891);
or I_36607 (I625906,I625889,I1299909);
DFFARX1 I_36608 (I625906,I3563,I625499,I625932,);
nor I_36609 (I625940,I625932,I625683);
DFFARX1 I_36610 (I625940,I3563,I625499,I625467,);
DFFARX1 I_36611 (I625932,I3563,I625499,I625491,);
not I_36612 (I625985,I625932);
nor I_36613 (I626002,I625985,I625559);
nor I_36614 (I626019,I625824,I626002);
DFFARX1 I_36615 (I626019,I3563,I625499,I625488,);
not I_36616 (I626077,I3570);
DFFARX1 I_36617 (I256548,I3563,I626077,I626103,);
not I_36618 (I626111,I626103);
DFFARX1 I_36619 (I256533,I3563,I626077,I626137,);
not I_36620 (I626145,I256551);
nand I_36621 (I626162,I626145,I256536);
not I_36622 (I626179,I626162);
nor I_36623 (I626196,I626179,I256533);
nor I_36624 (I626213,I626111,I626196);
DFFARX1 I_36625 (I626213,I3563,I626077,I626063,);
not I_36626 (I626244,I256533);
nand I_36627 (I626261,I626244,I626179);
and I_36628 (I626278,I626244,I256536);
nand I_36629 (I626295,I626278,I256557);
nor I_36630 (I626060,I626295,I626244);
and I_36631 (I626051,I626137,I626295);
not I_36632 (I626340,I626295);
nand I_36633 (I626054,I626137,I626340);
nor I_36634 (I626048,I626103,I626295);
not I_36635 (I626385,I256545);
nor I_36636 (I626402,I626385,I256536);
nand I_36637 (I626419,I626402,I626244);
nor I_36638 (I626057,I626162,I626419);
nor I_36639 (I626450,I626385,I256539);
and I_36640 (I626467,I626450,I256554);
or I_36641 (I626484,I626467,I256542);
DFFARX1 I_36642 (I626484,I3563,I626077,I626510,);
nor I_36643 (I626518,I626510,I626261);
DFFARX1 I_36644 (I626518,I3563,I626077,I626045,);
DFFARX1 I_36645 (I626510,I3563,I626077,I626069,);
not I_36646 (I626563,I626510);
nor I_36647 (I626580,I626563,I626137);
nor I_36648 (I626597,I626402,I626580);
DFFARX1 I_36649 (I626597,I3563,I626077,I626066,);
not I_36650 (I626655,I3570);
DFFARX1 I_36651 (I1000153,I3563,I626655,I626681,);
not I_36652 (I626689,I626681);
DFFARX1 I_36653 (I1000150,I3563,I626655,I626715,);
not I_36654 (I626723,I1000147);
nand I_36655 (I626740,I626723,I1000174);
not I_36656 (I626757,I626740);
nor I_36657 (I626774,I626757,I1000162);
nor I_36658 (I626791,I626689,I626774);
DFFARX1 I_36659 (I626791,I3563,I626655,I626641,);
not I_36660 (I626822,I1000162);
nand I_36661 (I626839,I626822,I626757);
and I_36662 (I626856,I626822,I1000168);
nand I_36663 (I626873,I626856,I1000159);
nor I_36664 (I626638,I626873,I626822);
and I_36665 (I626629,I626715,I626873);
not I_36666 (I626918,I626873);
nand I_36667 (I626632,I626715,I626918);
nor I_36668 (I626626,I626681,I626873);
not I_36669 (I626963,I1000156);
nor I_36670 (I626980,I626963,I1000168);
nand I_36671 (I626997,I626980,I626822);
nor I_36672 (I626635,I626740,I626997);
nor I_36673 (I627028,I626963,I1000171);
and I_36674 (I627045,I627028,I1000165);
or I_36675 (I627062,I627045,I1000147);
DFFARX1 I_36676 (I627062,I3563,I626655,I627088,);
nor I_36677 (I627096,I627088,I626839);
DFFARX1 I_36678 (I627096,I3563,I626655,I626623,);
DFFARX1 I_36679 (I627088,I3563,I626655,I626647,);
not I_36680 (I627141,I627088);
nor I_36681 (I627158,I627141,I626715);
nor I_36682 (I627175,I626980,I627158);
DFFARX1 I_36683 (I627175,I3563,I626655,I626644,);
not I_36684 (I627233,I3570);
DFFARX1 I_36685 (I349138,I3563,I627233,I627259,);
not I_36686 (I627267,I627259);
DFFARX1 I_36687 (I349153,I3563,I627233,I627293,);
not I_36688 (I627301,I349156);
nand I_36689 (I627318,I627301,I349135);
not I_36690 (I627335,I627318);
nor I_36691 (I627352,I627335,I349159);
nor I_36692 (I627369,I627267,I627352);
DFFARX1 I_36693 (I627369,I3563,I627233,I627219,);
not I_36694 (I627400,I349159);
nand I_36695 (I627417,I627400,I627335);
and I_36696 (I627434,I627400,I349141);
nand I_36697 (I627451,I627434,I349132);
nor I_36698 (I627216,I627451,I627400);
and I_36699 (I627207,I627293,I627451);
not I_36700 (I627496,I627451);
nand I_36701 (I627210,I627293,I627496);
nor I_36702 (I627204,I627259,I627451);
not I_36703 (I627541,I349132);
nor I_36704 (I627558,I627541,I349141);
nand I_36705 (I627575,I627558,I627400);
nor I_36706 (I627213,I627318,I627575);
nor I_36707 (I627606,I627541,I349147);
and I_36708 (I627623,I627606,I349150);
or I_36709 (I627640,I627623,I349144);
DFFARX1 I_36710 (I627640,I3563,I627233,I627666,);
nor I_36711 (I627674,I627666,I627417);
DFFARX1 I_36712 (I627674,I3563,I627233,I627201,);
DFFARX1 I_36713 (I627666,I3563,I627233,I627225,);
not I_36714 (I627719,I627666);
nor I_36715 (I627736,I627719,I627293);
nor I_36716 (I627753,I627558,I627736);
DFFARX1 I_36717 (I627753,I3563,I627233,I627222,);
not I_36718 (I627811,I3570);
DFFARX1 I_36719 (I1274715,I3563,I627811,I627837,);
not I_36720 (I627845,I627837);
DFFARX1 I_36721 (I1274709,I3563,I627811,I627871,);
not I_36722 (I627879,I1274718);
nand I_36723 (I627896,I627879,I1274697);
not I_36724 (I627913,I627896);
nor I_36725 (I627930,I627913,I1274706);
nor I_36726 (I627947,I627845,I627930);
DFFARX1 I_36727 (I627947,I3563,I627811,I627797,);
not I_36728 (I627978,I1274706);
nand I_36729 (I627995,I627978,I627913);
and I_36730 (I628012,I627978,I1274721);
nand I_36731 (I628029,I628012,I1274700);
nor I_36732 (I627794,I628029,I627978);
and I_36733 (I627785,I627871,I628029);
not I_36734 (I628074,I628029);
nand I_36735 (I627788,I627871,I628074);
nor I_36736 (I627782,I627837,I628029);
not I_36737 (I628119,I1274703);
nor I_36738 (I628136,I628119,I1274721);
nand I_36739 (I628153,I628136,I627978);
nor I_36740 (I627791,I627896,I628153);
nor I_36741 (I628184,I628119,I1274712);
and I_36742 (I628201,I628184,I1274700);
or I_36743 (I628218,I628201,I1274697);
DFFARX1 I_36744 (I628218,I3563,I627811,I628244,);
nor I_36745 (I628252,I628244,I627995);
DFFARX1 I_36746 (I628252,I3563,I627811,I627779,);
DFFARX1 I_36747 (I628244,I3563,I627811,I627803,);
not I_36748 (I628297,I628244);
nor I_36749 (I628314,I628297,I627871);
nor I_36750 (I628331,I628136,I628314);
DFFARX1 I_36751 (I628331,I3563,I627811,I627800,);
not I_36752 (I628389,I3570);
DFFARX1 I_36753 (I335436,I3563,I628389,I628415,);
not I_36754 (I628423,I628415);
DFFARX1 I_36755 (I335451,I3563,I628389,I628449,);
not I_36756 (I628457,I335454);
nand I_36757 (I628474,I628457,I335433);
not I_36758 (I628491,I628474);
nor I_36759 (I628508,I628491,I335457);
nor I_36760 (I628525,I628423,I628508);
DFFARX1 I_36761 (I628525,I3563,I628389,I628375,);
not I_36762 (I628556,I335457);
nand I_36763 (I628573,I628556,I628491);
and I_36764 (I628590,I628556,I335439);
nand I_36765 (I628607,I628590,I335430);
nor I_36766 (I628372,I628607,I628556);
and I_36767 (I628363,I628449,I628607);
not I_36768 (I628652,I628607);
nand I_36769 (I628366,I628449,I628652);
nor I_36770 (I628360,I628415,I628607);
not I_36771 (I628697,I335430);
nor I_36772 (I628714,I628697,I335439);
nand I_36773 (I628731,I628714,I628556);
nor I_36774 (I628369,I628474,I628731);
nor I_36775 (I628762,I628697,I335445);
and I_36776 (I628779,I628762,I335448);
or I_36777 (I628796,I628779,I335442);
DFFARX1 I_36778 (I628796,I3563,I628389,I628822,);
nor I_36779 (I628830,I628822,I628573);
DFFARX1 I_36780 (I628830,I3563,I628389,I628357,);
DFFARX1 I_36781 (I628822,I3563,I628389,I628381,);
not I_36782 (I628875,I628822);
nor I_36783 (I628892,I628875,I628449);
nor I_36784 (I628909,I628714,I628892);
DFFARX1 I_36785 (I628909,I3563,I628389,I628378,);
not I_36786 (I628967,I3570);
DFFARX1 I_36787 (I299073,I3563,I628967,I628993,);
not I_36788 (I629001,I628993);
DFFARX1 I_36789 (I299088,I3563,I628967,I629027,);
not I_36790 (I629035,I299091);
nand I_36791 (I629052,I629035,I299070);
not I_36792 (I629069,I629052);
nor I_36793 (I629086,I629069,I299094);
nor I_36794 (I629103,I629001,I629086);
DFFARX1 I_36795 (I629103,I3563,I628967,I628953,);
not I_36796 (I629134,I299094);
nand I_36797 (I629151,I629134,I629069);
and I_36798 (I629168,I629134,I299076);
nand I_36799 (I629185,I629168,I299067);
nor I_36800 (I628950,I629185,I629134);
and I_36801 (I628941,I629027,I629185);
not I_36802 (I629230,I629185);
nand I_36803 (I628944,I629027,I629230);
nor I_36804 (I628938,I628993,I629185);
not I_36805 (I629275,I299067);
nor I_36806 (I629292,I629275,I299076);
nand I_36807 (I629309,I629292,I629134);
nor I_36808 (I628947,I629052,I629309);
nor I_36809 (I629340,I629275,I299082);
and I_36810 (I629357,I629340,I299085);
or I_36811 (I629374,I629357,I299079);
DFFARX1 I_36812 (I629374,I3563,I628967,I629400,);
nor I_36813 (I629408,I629400,I629151);
DFFARX1 I_36814 (I629408,I3563,I628967,I628935,);
DFFARX1 I_36815 (I629400,I3563,I628967,I628959,);
not I_36816 (I629453,I629400);
nor I_36817 (I629470,I629453,I629027);
nor I_36818 (I629487,I629292,I629470);
DFFARX1 I_36819 (I629487,I3563,I628967,I628956,);
not I_36820 (I629545,I3570);
DFFARX1 I_36821 (I1273083,I3563,I629545,I629571,);
not I_36822 (I629579,I629571);
DFFARX1 I_36823 (I1273077,I3563,I629545,I629605,);
not I_36824 (I629613,I1273086);
nand I_36825 (I629630,I629613,I1273065);
not I_36826 (I629647,I629630);
nor I_36827 (I629664,I629647,I1273074);
nor I_36828 (I629681,I629579,I629664);
DFFARX1 I_36829 (I629681,I3563,I629545,I629531,);
not I_36830 (I629712,I1273074);
nand I_36831 (I629729,I629712,I629647);
and I_36832 (I629746,I629712,I1273089);
nand I_36833 (I629763,I629746,I1273068);
nor I_36834 (I629528,I629763,I629712);
and I_36835 (I629519,I629605,I629763);
not I_36836 (I629808,I629763);
nand I_36837 (I629522,I629605,I629808);
nor I_36838 (I629516,I629571,I629763);
not I_36839 (I629853,I1273071);
nor I_36840 (I629870,I629853,I1273089);
nand I_36841 (I629887,I629870,I629712);
nor I_36842 (I629525,I629630,I629887);
nor I_36843 (I629918,I629853,I1273080);
and I_36844 (I629935,I629918,I1273068);
or I_36845 (I629952,I629935,I1273065);
DFFARX1 I_36846 (I629952,I3563,I629545,I629978,);
nor I_36847 (I629986,I629978,I629729);
DFFARX1 I_36848 (I629986,I3563,I629545,I629513,);
DFFARX1 I_36849 (I629978,I3563,I629545,I629537,);
not I_36850 (I630031,I629978);
nor I_36851 (I630048,I630031,I629605);
nor I_36852 (I630065,I629870,I630048);
DFFARX1 I_36853 (I630065,I3563,I629545,I629534,);
not I_36854 (I630123,I3570);
DFFARX1 I_36855 (I1349378,I3563,I630123,I630149,);
not I_36856 (I630157,I630149);
DFFARX1 I_36857 (I1349378,I3563,I630123,I630183,);
not I_36858 (I630191,I1349402);
nand I_36859 (I630208,I630191,I1349384);
not I_36860 (I630225,I630208);
nor I_36861 (I630242,I630225,I1349399);
nor I_36862 (I630259,I630157,I630242);
DFFARX1 I_36863 (I630259,I3563,I630123,I630109,);
not I_36864 (I630290,I1349399);
nand I_36865 (I630307,I630290,I630225);
and I_36866 (I630324,I630290,I1349381);
nand I_36867 (I630341,I630324,I1349390);
nor I_36868 (I630106,I630341,I630290);
and I_36869 (I630097,I630183,I630341);
not I_36870 (I630386,I630341);
nand I_36871 (I630100,I630183,I630386);
nor I_36872 (I630094,I630149,I630341);
not I_36873 (I630431,I1349387);
nor I_36874 (I630448,I630431,I1349381);
nand I_36875 (I630465,I630448,I630290);
nor I_36876 (I630103,I630208,I630465);
nor I_36877 (I630496,I630431,I1349396);
and I_36878 (I630513,I630496,I1349405);
or I_36879 (I630530,I630513,I1349393);
DFFARX1 I_36880 (I630530,I3563,I630123,I630556,);
nor I_36881 (I630564,I630556,I630307);
DFFARX1 I_36882 (I630564,I3563,I630123,I630091,);
DFFARX1 I_36883 (I630556,I3563,I630123,I630115,);
not I_36884 (I630609,I630556);
nor I_36885 (I630626,I630609,I630183);
nor I_36886 (I630643,I630448,I630626);
DFFARX1 I_36887 (I630643,I3563,I630123,I630112,);
not I_36888 (I630701,I3570);
DFFARX1 I_36889 (I1346403,I3563,I630701,I630727,);
not I_36890 (I630735,I630727);
DFFARX1 I_36891 (I1346403,I3563,I630701,I630761,);
not I_36892 (I630769,I1346427);
nand I_36893 (I630786,I630769,I1346409);
not I_36894 (I630803,I630786);
nor I_36895 (I630820,I630803,I1346424);
nor I_36896 (I630837,I630735,I630820);
DFFARX1 I_36897 (I630837,I3563,I630701,I630687,);
not I_36898 (I630868,I1346424);
nand I_36899 (I630885,I630868,I630803);
and I_36900 (I630902,I630868,I1346406);
nand I_36901 (I630919,I630902,I1346415);
nor I_36902 (I630684,I630919,I630868);
and I_36903 (I630675,I630761,I630919);
not I_36904 (I630964,I630919);
nand I_36905 (I630678,I630761,I630964);
nor I_36906 (I630672,I630727,I630919);
not I_36907 (I631009,I1346412);
nor I_36908 (I631026,I631009,I1346406);
nand I_36909 (I631043,I631026,I630868);
nor I_36910 (I630681,I630786,I631043);
nor I_36911 (I631074,I631009,I1346421);
and I_36912 (I631091,I631074,I1346430);
or I_36913 (I631108,I631091,I1346418);
DFFARX1 I_36914 (I631108,I3563,I630701,I631134,);
nor I_36915 (I631142,I631134,I630885);
DFFARX1 I_36916 (I631142,I3563,I630701,I630669,);
DFFARX1 I_36917 (I631134,I3563,I630701,I630693,);
not I_36918 (I631187,I631134);
nor I_36919 (I631204,I631187,I630761);
nor I_36920 (I631221,I631026,I631204);
DFFARX1 I_36921 (I631221,I3563,I630701,I630690,);
not I_36922 (I631279,I3570);
DFFARX1 I_36923 (I118330,I3563,I631279,I631305,);
not I_36924 (I631313,I631305);
DFFARX1 I_36925 (I118309,I3563,I631279,I631339,);
not I_36926 (I631347,I118306);
nand I_36927 (I631364,I631347,I118321);
not I_36928 (I631381,I631364);
nor I_36929 (I631398,I631381,I118309);
nor I_36930 (I631415,I631313,I631398);
DFFARX1 I_36931 (I631415,I3563,I631279,I631265,);
not I_36932 (I631446,I118309);
nand I_36933 (I631463,I631446,I631381);
and I_36934 (I631480,I631446,I118312);
nand I_36935 (I631497,I631480,I118327);
nor I_36936 (I631262,I631497,I631446);
and I_36937 (I631253,I631339,I631497);
not I_36938 (I631542,I631497);
nand I_36939 (I631256,I631339,I631542);
nor I_36940 (I631250,I631305,I631497);
not I_36941 (I631587,I118318);
nor I_36942 (I631604,I631587,I118312);
nand I_36943 (I631621,I631604,I631446);
nor I_36944 (I631259,I631364,I631621);
nor I_36945 (I631652,I631587,I118306);
and I_36946 (I631669,I631652,I118315);
or I_36947 (I631686,I631669,I118324);
DFFARX1 I_36948 (I631686,I3563,I631279,I631712,);
nor I_36949 (I631720,I631712,I631463);
DFFARX1 I_36950 (I631720,I3563,I631279,I631247,);
DFFARX1 I_36951 (I631712,I3563,I631279,I631271,);
not I_36952 (I631765,I631712);
nor I_36953 (I631782,I631765,I631339);
nor I_36954 (I631799,I631604,I631782);
DFFARX1 I_36955 (I631799,I3563,I631279,I631268,);
not I_36956 (I631857,I3570);
DFFARX1 I_36957 (I1389838,I3563,I631857,I631883,);
not I_36958 (I631891,I631883);
DFFARX1 I_36959 (I1389838,I3563,I631857,I631917,);
not I_36960 (I631925,I1389862);
nand I_36961 (I631942,I631925,I1389844);
not I_36962 (I631959,I631942);
nor I_36963 (I631976,I631959,I1389859);
nor I_36964 (I631993,I631891,I631976);
DFFARX1 I_36965 (I631993,I3563,I631857,I631843,);
not I_36966 (I632024,I1389859);
nand I_36967 (I632041,I632024,I631959);
and I_36968 (I632058,I632024,I1389841);
nand I_36969 (I632075,I632058,I1389850);
nor I_36970 (I631840,I632075,I632024);
and I_36971 (I631831,I631917,I632075);
not I_36972 (I632120,I632075);
nand I_36973 (I631834,I631917,I632120);
nor I_36974 (I631828,I631883,I632075);
not I_36975 (I632165,I1389847);
nor I_36976 (I632182,I632165,I1389841);
nand I_36977 (I632199,I632182,I632024);
nor I_36978 (I631837,I631942,I632199);
nor I_36979 (I632230,I632165,I1389856);
and I_36980 (I632247,I632230,I1389865);
or I_36981 (I632264,I632247,I1389853);
DFFARX1 I_36982 (I632264,I3563,I631857,I632290,);
nor I_36983 (I632298,I632290,I632041);
DFFARX1 I_36984 (I632298,I3563,I631857,I631825,);
DFFARX1 I_36985 (I632290,I3563,I631857,I631849,);
not I_36986 (I632343,I632290);
nor I_36987 (I632360,I632343,I631917);
nor I_36988 (I632377,I632182,I632360);
DFFARX1 I_36989 (I632377,I3563,I631857,I631846,);
not I_36990 (I632435,I3570);
DFFARX1 I_36991 (I33989,I3563,I632435,I632461,);
not I_36992 (I632469,I632461);
DFFARX1 I_36993 (I33992,I3563,I632435,I632495,);
not I_36994 (I632503,I33986);
nand I_36995 (I632520,I632503,I34010);
not I_36996 (I632537,I632520);
nor I_36997 (I632554,I632537,I33989);
nor I_36998 (I632571,I632469,I632554);
DFFARX1 I_36999 (I632571,I3563,I632435,I632421,);
not I_37000 (I632602,I33989);
nand I_37001 (I632619,I632602,I632537);
and I_37002 (I632636,I632602,I34004);
nand I_37003 (I632653,I632636,I33998);
nor I_37004 (I632418,I632653,I632602);
and I_37005 (I632409,I632495,I632653);
not I_37006 (I632698,I632653);
nand I_37007 (I632412,I632495,I632698);
nor I_37008 (I632406,I632461,I632653);
not I_37009 (I632743,I34007);
nor I_37010 (I632760,I632743,I34004);
nand I_37011 (I632777,I632760,I632602);
nor I_37012 (I632415,I632520,I632777);
nor I_37013 (I632808,I632743,I33986);
and I_37014 (I632825,I632808,I33995);
or I_37015 (I632842,I632825,I34001);
DFFARX1 I_37016 (I632842,I3563,I632435,I632868,);
nor I_37017 (I632876,I632868,I632619);
DFFARX1 I_37018 (I632876,I3563,I632435,I632403,);
DFFARX1 I_37019 (I632868,I3563,I632435,I632427,);
not I_37020 (I632921,I632868);
nor I_37021 (I632938,I632921,I632495);
nor I_37022 (I632955,I632760,I632938);
DFFARX1 I_37023 (I632955,I3563,I632435,I632424,);
not I_37024 (I633013,I3570);
DFFARX1 I_37025 (I1101977,I3563,I633013,I633039,);
not I_37026 (I633047,I633039);
DFFARX1 I_37027 (I1101983,I3563,I633013,I633073,);
not I_37028 (I633081,I1101977);
nand I_37029 (I633098,I633081,I1101980);
not I_37030 (I633115,I633098);
nor I_37031 (I633132,I633115,I1101998);
nor I_37032 (I633149,I633047,I633132);
DFFARX1 I_37033 (I633149,I3563,I633013,I632999,);
not I_37034 (I633180,I1101998);
nand I_37035 (I633197,I633180,I633115);
and I_37036 (I633214,I633180,I1102001);
nand I_37037 (I633231,I633214,I1101980);
nor I_37038 (I632996,I633231,I633180);
and I_37039 (I632987,I633073,I633231);
not I_37040 (I633276,I633231);
nand I_37041 (I632990,I633073,I633276);
nor I_37042 (I632984,I633039,I633231);
not I_37043 (I633321,I1101986);
nor I_37044 (I633338,I633321,I1102001);
nand I_37045 (I633355,I633338,I633180);
nor I_37046 (I632993,I633098,I633355);
nor I_37047 (I633386,I633321,I1101992);
and I_37048 (I633403,I633386,I1101989);
or I_37049 (I633420,I633403,I1101995);
DFFARX1 I_37050 (I633420,I3563,I633013,I633446,);
nor I_37051 (I633454,I633446,I633197);
DFFARX1 I_37052 (I633454,I3563,I633013,I632981,);
DFFARX1 I_37053 (I633446,I3563,I633013,I633005,);
not I_37054 (I633499,I633446);
nor I_37055 (I633516,I633499,I633073);
nor I_37056 (I633533,I633338,I633516);
DFFARX1 I_37057 (I633533,I3563,I633013,I633002,);
not I_37058 (I633591,I3570);
DFFARX1 I_37059 (I357570,I3563,I633591,I633617,);
not I_37060 (I633625,I633617);
DFFARX1 I_37061 (I357585,I3563,I633591,I633651,);
not I_37062 (I633659,I357588);
nand I_37063 (I633676,I633659,I357567);
not I_37064 (I633693,I633676);
nor I_37065 (I633710,I633693,I357591);
nor I_37066 (I633727,I633625,I633710);
DFFARX1 I_37067 (I633727,I3563,I633591,I633577,);
not I_37068 (I633758,I357591);
nand I_37069 (I633775,I633758,I633693);
and I_37070 (I633792,I633758,I357573);
nand I_37071 (I633809,I633792,I357564);
nor I_37072 (I633574,I633809,I633758);
and I_37073 (I633565,I633651,I633809);
not I_37074 (I633854,I633809);
nand I_37075 (I633568,I633651,I633854);
nor I_37076 (I633562,I633617,I633809);
not I_37077 (I633899,I357564);
nor I_37078 (I633916,I633899,I357573);
nand I_37079 (I633933,I633916,I633758);
nor I_37080 (I633571,I633676,I633933);
nor I_37081 (I633964,I633899,I357579);
and I_37082 (I633981,I633964,I357582);
or I_37083 (I633998,I633981,I357576);
DFFARX1 I_37084 (I633998,I3563,I633591,I634024,);
nor I_37085 (I634032,I634024,I633775);
DFFARX1 I_37086 (I634032,I3563,I633591,I633559,);
DFFARX1 I_37087 (I634024,I3563,I633591,I633583,);
not I_37088 (I634077,I634024);
nor I_37089 (I634094,I634077,I633651);
nor I_37090 (I634111,I633916,I634094);
DFFARX1 I_37091 (I634111,I3563,I633591,I633580,);
not I_37092 (I634169,I3570);
DFFARX1 I_37093 (I918757,I3563,I634169,I634195,);
not I_37094 (I634203,I634195);
DFFARX1 I_37095 (I918754,I3563,I634169,I634229,);
not I_37096 (I634237,I918751);
nand I_37097 (I634254,I634237,I918778);
not I_37098 (I634271,I634254);
nor I_37099 (I634288,I634271,I918766);
nor I_37100 (I634305,I634203,I634288);
DFFARX1 I_37101 (I634305,I3563,I634169,I634155,);
not I_37102 (I634336,I918766);
nand I_37103 (I634353,I634336,I634271);
and I_37104 (I634370,I634336,I918772);
nand I_37105 (I634387,I634370,I918763);
nor I_37106 (I634152,I634387,I634336);
and I_37107 (I634143,I634229,I634387);
not I_37108 (I634432,I634387);
nand I_37109 (I634146,I634229,I634432);
nor I_37110 (I634140,I634195,I634387);
not I_37111 (I634477,I918760);
nor I_37112 (I634494,I634477,I918772);
nand I_37113 (I634511,I634494,I634336);
nor I_37114 (I634149,I634254,I634511);
nor I_37115 (I634542,I634477,I918775);
and I_37116 (I634559,I634542,I918769);
or I_37117 (I634576,I634559,I918751);
DFFARX1 I_37118 (I634576,I3563,I634169,I634602,);
nor I_37119 (I634610,I634602,I634353);
DFFARX1 I_37120 (I634610,I3563,I634169,I634137,);
DFFARX1 I_37121 (I634602,I3563,I634169,I634161,);
not I_37122 (I634655,I634602);
nor I_37123 (I634672,I634655,I634229);
nor I_37124 (I634689,I634494,I634672);
DFFARX1 I_37125 (I634689,I3563,I634169,I634158,);
not I_37126 (I634747,I3570);
DFFARX1 I_37127 (I462126,I3563,I634747,I634773,);
not I_37128 (I634781,I634773);
DFFARX1 I_37129 (I462138,I3563,I634747,I634807,);
not I_37130 (I634815,I462114);
nand I_37131 (I634832,I634815,I462141);
not I_37132 (I634849,I634832);
nor I_37133 (I634866,I634849,I462129);
nor I_37134 (I634883,I634781,I634866);
DFFARX1 I_37135 (I634883,I3563,I634747,I634733,);
not I_37136 (I634914,I462129);
nand I_37137 (I634931,I634914,I634849);
and I_37138 (I634948,I634914,I462114);
nand I_37139 (I634965,I634948,I462117);
nor I_37140 (I634730,I634965,I634914);
and I_37141 (I634721,I634807,I634965);
not I_37142 (I635010,I634965);
nand I_37143 (I634724,I634807,I635010);
nor I_37144 (I634718,I634773,I634965);
not I_37145 (I635055,I462123);
nor I_37146 (I635072,I635055,I462114);
nand I_37147 (I635089,I635072,I634914);
nor I_37148 (I634727,I634832,I635089);
nor I_37149 (I635120,I635055,I462132);
and I_37150 (I635137,I635120,I462120);
or I_37151 (I635154,I635137,I462135);
DFFARX1 I_37152 (I635154,I3563,I634747,I635180,);
nor I_37153 (I635188,I635180,I634931);
DFFARX1 I_37154 (I635188,I3563,I634747,I634715,);
DFFARX1 I_37155 (I635180,I3563,I634747,I634739,);
not I_37156 (I635233,I635180);
nor I_37157 (I635250,I635233,I634807);
nor I_37158 (I635267,I635072,I635250);
DFFARX1 I_37159 (I635267,I3563,I634747,I634736,);
not I_37160 (I635325,I3570);
DFFARX1 I_37161 (I328058,I3563,I635325,I635351,);
not I_37162 (I635359,I635351);
DFFARX1 I_37163 (I328073,I3563,I635325,I635385,);
not I_37164 (I635393,I328076);
nand I_37165 (I635410,I635393,I328055);
not I_37166 (I635427,I635410);
nor I_37167 (I635444,I635427,I328079);
nor I_37168 (I635461,I635359,I635444);
DFFARX1 I_37169 (I635461,I3563,I635325,I635311,);
not I_37170 (I635492,I328079);
nand I_37171 (I635509,I635492,I635427);
and I_37172 (I635526,I635492,I328061);
nand I_37173 (I635543,I635526,I328052);
nor I_37174 (I635308,I635543,I635492);
and I_37175 (I635299,I635385,I635543);
not I_37176 (I635588,I635543);
nand I_37177 (I635302,I635385,I635588);
nor I_37178 (I635296,I635351,I635543);
not I_37179 (I635633,I328052);
nor I_37180 (I635650,I635633,I328061);
nand I_37181 (I635667,I635650,I635492);
nor I_37182 (I635305,I635410,I635667);
nor I_37183 (I635698,I635633,I328067);
and I_37184 (I635715,I635698,I328070);
or I_37185 (I635732,I635715,I328064);
DFFARX1 I_37186 (I635732,I3563,I635325,I635758,);
nor I_37187 (I635766,I635758,I635509);
DFFARX1 I_37188 (I635766,I3563,I635325,I635293,);
DFFARX1 I_37189 (I635758,I3563,I635325,I635317,);
not I_37190 (I635811,I635758);
nor I_37191 (I635828,I635811,I635385);
nor I_37192 (I635845,I635650,I635828);
DFFARX1 I_37193 (I635845,I3563,I635325,I635314,);
not I_37194 (I635903,I3570);
DFFARX1 I_37195 (I732975,I3563,I635903,I635929,);
not I_37196 (I635937,I635929);
DFFARX1 I_37197 (I732987,I3563,I635903,I635963,);
not I_37198 (I635971,I732978);
nand I_37199 (I635988,I635971,I732981);
not I_37200 (I636005,I635988);
nor I_37201 (I636022,I636005,I732984);
nor I_37202 (I636039,I635937,I636022);
DFFARX1 I_37203 (I636039,I3563,I635903,I635889,);
not I_37204 (I636070,I732984);
nand I_37205 (I636087,I636070,I636005);
and I_37206 (I636104,I636070,I732978);
nand I_37207 (I636121,I636104,I732990);
nor I_37208 (I635886,I636121,I636070);
and I_37209 (I635877,I635963,I636121);
not I_37210 (I636166,I636121);
nand I_37211 (I635880,I635963,I636166);
nor I_37212 (I635874,I635929,I636121);
not I_37213 (I636211,I732996);
nor I_37214 (I636228,I636211,I732978);
nand I_37215 (I636245,I636228,I636070);
nor I_37216 (I635883,I635988,I636245);
nor I_37217 (I636276,I636211,I732975);
and I_37218 (I636293,I636276,I732993);
or I_37219 (I636310,I636293,I732999);
DFFARX1 I_37220 (I636310,I3563,I635903,I636336,);
nor I_37221 (I636344,I636336,I636087);
DFFARX1 I_37222 (I636344,I3563,I635903,I635871,);
DFFARX1 I_37223 (I636336,I3563,I635903,I635895,);
not I_37224 (I636389,I636336);
nor I_37225 (I636406,I636389,I635963);
nor I_37226 (I636423,I636228,I636406);
DFFARX1 I_37227 (I636423,I3563,I635903,I635892,);
not I_37228 (I636481,I3570);
DFFARX1 I_37229 (I151004,I3563,I636481,I636507,);
not I_37230 (I636515,I636507);
DFFARX1 I_37231 (I150983,I3563,I636481,I636541,);
not I_37232 (I636549,I150980);
nand I_37233 (I636566,I636549,I150995);
not I_37234 (I636583,I636566);
nor I_37235 (I636600,I636583,I150983);
nor I_37236 (I636617,I636515,I636600);
DFFARX1 I_37237 (I636617,I3563,I636481,I636467,);
not I_37238 (I636648,I150983);
nand I_37239 (I636665,I636648,I636583);
and I_37240 (I636682,I636648,I150986);
nand I_37241 (I636699,I636682,I151001);
nor I_37242 (I636464,I636699,I636648);
and I_37243 (I636455,I636541,I636699);
not I_37244 (I636744,I636699);
nand I_37245 (I636458,I636541,I636744);
nor I_37246 (I636452,I636507,I636699);
not I_37247 (I636789,I150992);
nor I_37248 (I636806,I636789,I150986);
nand I_37249 (I636823,I636806,I636648);
nor I_37250 (I636461,I636566,I636823);
nor I_37251 (I636854,I636789,I150980);
and I_37252 (I636871,I636854,I150989);
or I_37253 (I636888,I636871,I150998);
DFFARX1 I_37254 (I636888,I3563,I636481,I636914,);
nor I_37255 (I636922,I636914,I636665);
DFFARX1 I_37256 (I636922,I3563,I636481,I636449,);
DFFARX1 I_37257 (I636914,I3563,I636481,I636473,);
not I_37258 (I636967,I636914);
nor I_37259 (I636984,I636967,I636541);
nor I_37260 (I637001,I636806,I636984);
DFFARX1 I_37261 (I637001,I3563,I636481,I636470,);
not I_37262 (I637059,I3570);
DFFARX1 I_37263 (I1035037,I3563,I637059,I637085,);
not I_37264 (I637093,I637085);
DFFARX1 I_37265 (I1035034,I3563,I637059,I637119,);
not I_37266 (I637127,I1035031);
nand I_37267 (I637144,I637127,I1035058);
not I_37268 (I637161,I637144);
nor I_37269 (I637178,I637161,I1035046);
nor I_37270 (I637195,I637093,I637178);
DFFARX1 I_37271 (I637195,I3563,I637059,I637045,);
not I_37272 (I637226,I1035046);
nand I_37273 (I637243,I637226,I637161);
and I_37274 (I637260,I637226,I1035052);
nand I_37275 (I637277,I637260,I1035043);
nor I_37276 (I637042,I637277,I637226);
and I_37277 (I637033,I637119,I637277);
not I_37278 (I637322,I637277);
nand I_37279 (I637036,I637119,I637322);
nor I_37280 (I637030,I637085,I637277);
not I_37281 (I637367,I1035040);
nor I_37282 (I637384,I637367,I1035052);
nand I_37283 (I637401,I637384,I637226);
nor I_37284 (I637039,I637144,I637401);
nor I_37285 (I637432,I637367,I1035055);
and I_37286 (I637449,I637432,I1035049);
or I_37287 (I637466,I637449,I1035031);
DFFARX1 I_37288 (I637466,I3563,I637059,I637492,);
nor I_37289 (I637500,I637492,I637243);
DFFARX1 I_37290 (I637500,I3563,I637059,I637027,);
DFFARX1 I_37291 (I637492,I3563,I637059,I637051,);
not I_37292 (I637545,I637492);
nor I_37293 (I637562,I637545,I637119);
nor I_37294 (I637579,I637384,I637562);
DFFARX1 I_37295 (I637579,I3563,I637059,I637048,);
not I_37296 (I637637,I3570);
DFFARX1 I_37297 (I178603,I3563,I637637,I637663,);
not I_37298 (I637671,I637663);
DFFARX1 I_37299 (I178588,I3563,I637637,I637697,);
not I_37300 (I637705,I178606);
nand I_37301 (I637722,I637705,I178591);
not I_37302 (I637739,I637722);
nor I_37303 (I637756,I637739,I178588);
nor I_37304 (I637773,I637671,I637756);
DFFARX1 I_37305 (I637773,I3563,I637637,I637623,);
not I_37306 (I637804,I178588);
nand I_37307 (I637821,I637804,I637739);
and I_37308 (I637838,I637804,I178591);
nand I_37309 (I637855,I637838,I178612);
nor I_37310 (I637620,I637855,I637804);
and I_37311 (I637611,I637697,I637855);
not I_37312 (I637900,I637855);
nand I_37313 (I637614,I637697,I637900);
nor I_37314 (I637608,I637663,I637855);
not I_37315 (I637945,I178600);
nor I_37316 (I637962,I637945,I178591);
nand I_37317 (I637979,I637962,I637804);
nor I_37318 (I637617,I637722,I637979);
nor I_37319 (I638010,I637945,I178594);
and I_37320 (I638027,I638010,I178609);
or I_37321 (I638044,I638027,I178597);
DFFARX1 I_37322 (I638044,I3563,I637637,I638070,);
nor I_37323 (I638078,I638070,I637821);
DFFARX1 I_37324 (I638078,I3563,I637637,I637605,);
DFFARX1 I_37325 (I638070,I3563,I637637,I637629,);
not I_37326 (I638123,I638070);
nor I_37327 (I638140,I638123,I637697);
nor I_37328 (I638157,I637962,I638140);
DFFARX1 I_37329 (I638157,I3563,I637637,I637626,);
not I_37330 (I638215,I3570);
DFFARX1 I_37331 (I979481,I3563,I638215,I638241,);
not I_37332 (I638249,I638241);
DFFARX1 I_37333 (I979478,I3563,I638215,I638275,);
not I_37334 (I638283,I979475);
nand I_37335 (I638300,I638283,I979502);
not I_37336 (I638317,I638300);
nor I_37337 (I638334,I638317,I979490);
nor I_37338 (I638351,I638249,I638334);
DFFARX1 I_37339 (I638351,I3563,I638215,I638201,);
not I_37340 (I638382,I979490);
nand I_37341 (I638399,I638382,I638317);
and I_37342 (I638416,I638382,I979496);
nand I_37343 (I638433,I638416,I979487);
nor I_37344 (I638198,I638433,I638382);
and I_37345 (I638189,I638275,I638433);
not I_37346 (I638478,I638433);
nand I_37347 (I638192,I638275,I638478);
nor I_37348 (I638186,I638241,I638433);
not I_37349 (I638523,I979484);
nor I_37350 (I638540,I638523,I979496);
nand I_37351 (I638557,I638540,I638382);
nor I_37352 (I638195,I638300,I638557);
nor I_37353 (I638588,I638523,I979499);
and I_37354 (I638605,I638588,I979493);
or I_37355 (I638622,I638605,I979475);
DFFARX1 I_37356 (I638622,I3563,I638215,I638648,);
nor I_37357 (I638656,I638648,I638399);
DFFARX1 I_37358 (I638656,I3563,I638215,I638183,);
DFFARX1 I_37359 (I638648,I3563,I638215,I638207,);
not I_37360 (I638701,I638648);
nor I_37361 (I638718,I638701,I638275);
nor I_37362 (I638735,I638540,I638718);
DFFARX1 I_37363 (I638735,I3563,I638215,I638204,);
not I_37364 (I638793,I3570);
DFFARX1 I_37365 (I723149,I3563,I638793,I638819,);
not I_37366 (I638827,I638819);
DFFARX1 I_37367 (I723161,I3563,I638793,I638853,);
not I_37368 (I638861,I723152);
nand I_37369 (I638878,I638861,I723155);
not I_37370 (I638895,I638878);
nor I_37371 (I638912,I638895,I723158);
nor I_37372 (I638929,I638827,I638912);
DFFARX1 I_37373 (I638929,I3563,I638793,I638779,);
not I_37374 (I638960,I723158);
nand I_37375 (I638977,I638960,I638895);
and I_37376 (I638994,I638960,I723152);
nand I_37377 (I639011,I638994,I723164);
nor I_37378 (I638776,I639011,I638960);
and I_37379 (I638767,I638853,I639011);
not I_37380 (I639056,I639011);
nand I_37381 (I638770,I638853,I639056);
nor I_37382 (I638764,I638819,I639011);
not I_37383 (I639101,I723170);
nor I_37384 (I639118,I639101,I723152);
nand I_37385 (I639135,I639118,I638960);
nor I_37386 (I638773,I638878,I639135);
nor I_37387 (I639166,I639101,I723149);
and I_37388 (I639183,I639166,I723167);
or I_37389 (I639200,I639183,I723173);
DFFARX1 I_37390 (I639200,I3563,I638793,I639226,);
nor I_37391 (I639234,I639226,I638977);
DFFARX1 I_37392 (I639234,I3563,I638793,I638761,);
DFFARX1 I_37393 (I639226,I3563,I638793,I638785,);
not I_37394 (I639279,I639226);
nor I_37395 (I639296,I639279,I638853);
nor I_37396 (I639313,I639118,I639296);
DFFARX1 I_37397 (I639313,I3563,I638793,I638782,);
not I_37398 (I639371,I3570);
DFFARX1 I_37399 (I1245339,I3563,I639371,I639397,);
not I_37400 (I639405,I639397);
DFFARX1 I_37401 (I1245333,I3563,I639371,I639431,);
not I_37402 (I639439,I1245342);
nand I_37403 (I639456,I639439,I1245321);
not I_37404 (I639473,I639456);
nor I_37405 (I639490,I639473,I1245330);
nor I_37406 (I639507,I639405,I639490);
DFFARX1 I_37407 (I639507,I3563,I639371,I639357,);
not I_37408 (I639538,I1245330);
nand I_37409 (I639555,I639538,I639473);
and I_37410 (I639572,I639538,I1245345);
nand I_37411 (I639589,I639572,I1245324);
nor I_37412 (I639354,I639589,I639538);
and I_37413 (I639345,I639431,I639589);
not I_37414 (I639634,I639589);
nand I_37415 (I639348,I639431,I639634);
nor I_37416 (I639342,I639397,I639589);
not I_37417 (I639679,I1245327);
nor I_37418 (I639696,I639679,I1245345);
nand I_37419 (I639713,I639696,I639538);
nor I_37420 (I639351,I639456,I639713);
nor I_37421 (I639744,I639679,I1245336);
and I_37422 (I639761,I639744,I1245324);
or I_37423 (I639778,I639761,I1245321);
DFFARX1 I_37424 (I639778,I3563,I639371,I639804,);
nor I_37425 (I639812,I639804,I639555);
DFFARX1 I_37426 (I639812,I3563,I639371,I639339,);
DFFARX1 I_37427 (I639804,I3563,I639371,I639363,);
not I_37428 (I639857,I639804);
nor I_37429 (I639874,I639857,I639431);
nor I_37430 (I639891,I639696,I639874);
DFFARX1 I_37431 (I639891,I3563,I639371,I639360,);
not I_37432 (I639949,I3570);
DFFARX1 I_37433 (I727195,I3563,I639949,I639975,);
not I_37434 (I639983,I639975);
DFFARX1 I_37435 (I727207,I3563,I639949,I640009,);
not I_37436 (I640017,I727198);
nand I_37437 (I640034,I640017,I727201);
not I_37438 (I640051,I640034);
nor I_37439 (I640068,I640051,I727204);
nor I_37440 (I640085,I639983,I640068);
DFFARX1 I_37441 (I640085,I3563,I639949,I639935,);
not I_37442 (I640116,I727204);
nand I_37443 (I640133,I640116,I640051);
and I_37444 (I640150,I640116,I727198);
nand I_37445 (I640167,I640150,I727210);
nor I_37446 (I639932,I640167,I640116);
and I_37447 (I639923,I640009,I640167);
not I_37448 (I640212,I640167);
nand I_37449 (I639926,I640009,I640212);
nor I_37450 (I639920,I639975,I640167);
not I_37451 (I640257,I727216);
nor I_37452 (I640274,I640257,I727198);
nand I_37453 (I640291,I640274,I640116);
nor I_37454 (I639929,I640034,I640291);
nor I_37455 (I640322,I640257,I727195);
and I_37456 (I640339,I640322,I727213);
or I_37457 (I640356,I640339,I727219);
DFFARX1 I_37458 (I640356,I3563,I639949,I640382,);
nor I_37459 (I640390,I640382,I640133);
DFFARX1 I_37460 (I640390,I3563,I639949,I639917,);
DFFARX1 I_37461 (I640382,I3563,I639949,I639941,);
not I_37462 (I640435,I640382);
nor I_37463 (I640452,I640435,I640009);
nor I_37464 (I640469,I640274,I640452);
DFFARX1 I_37465 (I640469,I3563,I639949,I639938,);
not I_37466 (I640527,I3570);
DFFARX1 I_37467 (I180983,I3563,I640527,I640553,);
not I_37468 (I640561,I640553);
DFFARX1 I_37469 (I180968,I3563,I640527,I640587,);
not I_37470 (I640595,I180986);
nand I_37471 (I640612,I640595,I180971);
not I_37472 (I640629,I640612);
nor I_37473 (I640646,I640629,I180968);
nor I_37474 (I640663,I640561,I640646);
DFFARX1 I_37475 (I640663,I3563,I640527,I640513,);
not I_37476 (I640694,I180968);
nand I_37477 (I640711,I640694,I640629);
and I_37478 (I640728,I640694,I180971);
nand I_37479 (I640745,I640728,I180992);
nor I_37480 (I640510,I640745,I640694);
and I_37481 (I640501,I640587,I640745);
not I_37482 (I640790,I640745);
nand I_37483 (I640504,I640587,I640790);
nor I_37484 (I640498,I640553,I640745);
not I_37485 (I640835,I180980);
nor I_37486 (I640852,I640835,I180971);
nand I_37487 (I640869,I640852,I640694);
nor I_37488 (I640507,I640612,I640869);
nor I_37489 (I640900,I640835,I180974);
and I_37490 (I640917,I640900,I180989);
or I_37491 (I640934,I640917,I180977);
DFFARX1 I_37492 (I640934,I3563,I640527,I640960,);
nor I_37493 (I640968,I640960,I640711);
DFFARX1 I_37494 (I640968,I3563,I640527,I640495,);
DFFARX1 I_37495 (I640960,I3563,I640527,I640519,);
not I_37496 (I641013,I640960);
nor I_37497 (I641030,I641013,I640587);
nor I_37498 (I641047,I640852,I641030);
DFFARX1 I_37499 (I641047,I3563,I640527,I640516,);
not I_37500 (I641105,I3570);
DFFARX1 I_37501 (I806381,I3563,I641105,I641131,);
not I_37502 (I641139,I641131);
DFFARX1 I_37503 (I806393,I3563,I641105,I641165,);
not I_37504 (I641173,I806384);
nand I_37505 (I641190,I641173,I806387);
not I_37506 (I641207,I641190);
nor I_37507 (I641224,I641207,I806390);
nor I_37508 (I641241,I641139,I641224);
DFFARX1 I_37509 (I641241,I3563,I641105,I641091,);
not I_37510 (I641272,I806390);
nand I_37511 (I641289,I641272,I641207);
and I_37512 (I641306,I641272,I806384);
nand I_37513 (I641323,I641306,I806396);
nor I_37514 (I641088,I641323,I641272);
and I_37515 (I641079,I641165,I641323);
not I_37516 (I641368,I641323);
nand I_37517 (I641082,I641165,I641368);
nor I_37518 (I641076,I641131,I641323);
not I_37519 (I641413,I806402);
nor I_37520 (I641430,I641413,I806384);
nand I_37521 (I641447,I641430,I641272);
nor I_37522 (I641085,I641190,I641447);
nor I_37523 (I641478,I641413,I806381);
and I_37524 (I641495,I641478,I806399);
or I_37525 (I641512,I641495,I806405);
DFFARX1 I_37526 (I641512,I3563,I641105,I641538,);
nor I_37527 (I641546,I641538,I641289);
DFFARX1 I_37528 (I641546,I3563,I641105,I641073,);
DFFARX1 I_37529 (I641538,I3563,I641105,I641097,);
not I_37530 (I641591,I641538);
nor I_37531 (I641608,I641591,I641165);
nor I_37532 (I641625,I641430,I641608);
DFFARX1 I_37533 (I641625,I3563,I641105,I641094,);
not I_37534 (I641683,I3570);
DFFARX1 I_37535 (I447982,I3563,I641683,I641709,);
not I_37536 (I641717,I641709);
DFFARX1 I_37537 (I447994,I3563,I641683,I641743,);
not I_37538 (I641751,I447970);
nand I_37539 (I641768,I641751,I447997);
not I_37540 (I641785,I641768);
nor I_37541 (I641802,I641785,I447985);
nor I_37542 (I641819,I641717,I641802);
DFFARX1 I_37543 (I641819,I3563,I641683,I641669,);
not I_37544 (I641850,I447985);
nand I_37545 (I641867,I641850,I641785);
and I_37546 (I641884,I641850,I447970);
nand I_37547 (I641901,I641884,I447973);
nor I_37548 (I641666,I641901,I641850);
and I_37549 (I641657,I641743,I641901);
not I_37550 (I641946,I641901);
nand I_37551 (I641660,I641743,I641946);
nor I_37552 (I641654,I641709,I641901);
not I_37553 (I641991,I447979);
nor I_37554 (I642008,I641991,I447970);
nand I_37555 (I642025,I642008,I641850);
nor I_37556 (I641663,I641768,I642025);
nor I_37557 (I642056,I641991,I447988);
and I_37558 (I642073,I642056,I447976);
or I_37559 (I642090,I642073,I447991);
DFFARX1 I_37560 (I642090,I3563,I641683,I642116,);
nor I_37561 (I642124,I642116,I641867);
DFFARX1 I_37562 (I642124,I3563,I641683,I641651,);
DFFARX1 I_37563 (I642116,I3563,I641683,I641675,);
not I_37564 (I642169,I642116);
nor I_37565 (I642186,I642169,I641743);
nor I_37566 (I642203,I642008,I642186);
DFFARX1 I_37567 (I642203,I3563,I641683,I641672,);
not I_37568 (I642261,I3570);
DFFARX1 I_37569 (I1295279,I3563,I642261,I642287,);
not I_37570 (I642295,I642287);
DFFARX1 I_37571 (I1295291,I3563,I642261,I642321,);
not I_37572 (I642329,I1295282);
nand I_37573 (I642346,I642329,I1295270);
not I_37574 (I642363,I642346);
nor I_37575 (I642380,I642363,I1295267);
nor I_37576 (I642397,I642295,I642380);
DFFARX1 I_37577 (I642397,I3563,I642261,I642247,);
not I_37578 (I642428,I1295267);
nand I_37579 (I642445,I642428,I642363);
and I_37580 (I642462,I642428,I1295273);
nand I_37581 (I642479,I642462,I1295270);
nor I_37582 (I642244,I642479,I642428);
and I_37583 (I642235,I642321,I642479);
not I_37584 (I642524,I642479);
nand I_37585 (I642238,I642321,I642524);
nor I_37586 (I642232,I642287,I642479);
not I_37587 (I642569,I1295288);
nor I_37588 (I642586,I642569,I1295273);
nand I_37589 (I642603,I642586,I642428);
nor I_37590 (I642241,I642346,I642603);
nor I_37591 (I642634,I642569,I1295276);
and I_37592 (I642651,I642634,I1295267);
or I_37593 (I642668,I642651,I1295285);
DFFARX1 I_37594 (I642668,I3563,I642261,I642694,);
nor I_37595 (I642702,I642694,I642445);
DFFARX1 I_37596 (I642702,I3563,I642261,I642229,);
DFFARX1 I_37597 (I642694,I3563,I642261,I642253,);
not I_37598 (I642747,I642694);
nor I_37599 (I642764,I642747,I642321);
nor I_37600 (I642781,I642586,I642764);
DFFARX1 I_37601 (I642781,I3563,I642261,I642250,);
not I_37602 (I642839,I3570);
DFFARX1 I_37603 (I662459,I3563,I642839,I642865,);
not I_37604 (I642873,I642865);
DFFARX1 I_37605 (I662471,I3563,I642839,I642899,);
not I_37606 (I642907,I662462);
nand I_37607 (I642924,I642907,I662465);
not I_37608 (I642941,I642924);
nor I_37609 (I642958,I642941,I662468);
nor I_37610 (I642975,I642873,I642958);
DFFARX1 I_37611 (I642975,I3563,I642839,I642825,);
not I_37612 (I643006,I662468);
nand I_37613 (I643023,I643006,I642941);
and I_37614 (I643040,I643006,I662462);
nand I_37615 (I643057,I643040,I662474);
nor I_37616 (I642822,I643057,I643006);
and I_37617 (I642813,I642899,I643057);
not I_37618 (I643102,I643057);
nand I_37619 (I642816,I642899,I643102);
nor I_37620 (I642810,I642865,I643057);
not I_37621 (I643147,I662480);
nor I_37622 (I643164,I643147,I662462);
nand I_37623 (I643181,I643164,I643006);
nor I_37624 (I642819,I642924,I643181);
nor I_37625 (I643212,I643147,I662459);
and I_37626 (I643229,I643212,I662477);
or I_37627 (I643246,I643229,I662483);
DFFARX1 I_37628 (I643246,I3563,I642839,I643272,);
nor I_37629 (I643280,I643272,I643023);
DFFARX1 I_37630 (I643280,I3563,I642839,I642807,);
DFFARX1 I_37631 (I643272,I3563,I642839,I642831,);
not I_37632 (I643325,I643272);
nor I_37633 (I643342,I643325,I642899);
nor I_37634 (I643359,I643164,I643342);
DFFARX1 I_37635 (I643359,I3563,I642839,I642828,);
not I_37636 (I643417,I3570);
DFFARX1 I_37637 (I529284,I3563,I643417,I643443,);
not I_37638 (I643451,I643443);
DFFARX1 I_37639 (I529296,I3563,I643417,I643477,);
not I_37640 (I643485,I529302);
nand I_37641 (I643502,I643485,I529293);
not I_37642 (I643519,I643502);
nor I_37643 (I643536,I643519,I529299);
nor I_37644 (I643553,I643451,I643536);
DFFARX1 I_37645 (I643553,I3563,I643417,I643403,);
not I_37646 (I643584,I529299);
nand I_37647 (I643601,I643584,I643519);
and I_37648 (I643618,I643584,I529290);
nand I_37649 (I643635,I643618,I529281);
nor I_37650 (I643400,I643635,I643584);
and I_37651 (I643391,I643477,I643635);
not I_37652 (I643680,I643635);
nand I_37653 (I643394,I643477,I643680);
nor I_37654 (I643388,I643443,I643635);
not I_37655 (I643725,I529287);
nor I_37656 (I643742,I643725,I529290);
nand I_37657 (I643759,I643742,I643584);
nor I_37658 (I643397,I643502,I643759);
nor I_37659 (I643790,I643725,I529284);
and I_37660 (I643807,I643790,I529281);
or I_37661 (I643824,I643807,I529305);
DFFARX1 I_37662 (I643824,I3563,I643417,I643850,);
nor I_37663 (I643858,I643850,I643601);
DFFARX1 I_37664 (I643858,I3563,I643417,I643385,);
DFFARX1 I_37665 (I643850,I3563,I643417,I643409,);
not I_37666 (I643903,I643850);
nor I_37667 (I643920,I643903,I643477);
nor I_37668 (I643937,I643742,I643920);
DFFARX1 I_37669 (I643937,I3563,I643417,I643406,);
not I_37670 (I643995,I3570);
DFFARX1 I_37671 (I741645,I3563,I643995,I644021,);
not I_37672 (I644029,I644021);
DFFARX1 I_37673 (I741657,I3563,I643995,I644055,);
not I_37674 (I644063,I741648);
nand I_37675 (I644080,I644063,I741651);
not I_37676 (I644097,I644080);
nor I_37677 (I644114,I644097,I741654);
nor I_37678 (I644131,I644029,I644114);
DFFARX1 I_37679 (I644131,I3563,I643995,I643981,);
not I_37680 (I644162,I741654);
nand I_37681 (I644179,I644162,I644097);
and I_37682 (I644196,I644162,I741648);
nand I_37683 (I644213,I644196,I741660);
nor I_37684 (I643978,I644213,I644162);
and I_37685 (I643969,I644055,I644213);
not I_37686 (I644258,I644213);
nand I_37687 (I643972,I644055,I644258);
nor I_37688 (I643966,I644021,I644213);
not I_37689 (I644303,I741666);
nor I_37690 (I644320,I644303,I741648);
nand I_37691 (I644337,I644320,I644162);
nor I_37692 (I643975,I644080,I644337);
nor I_37693 (I644368,I644303,I741645);
and I_37694 (I644385,I644368,I741663);
or I_37695 (I644402,I644385,I741669);
DFFARX1 I_37696 (I644402,I3563,I643995,I644428,);
nor I_37697 (I644436,I644428,I644179);
DFFARX1 I_37698 (I644436,I3563,I643995,I643963,);
DFFARX1 I_37699 (I644428,I3563,I643995,I643987,);
not I_37700 (I644481,I644428);
nor I_37701 (I644498,I644481,I644055);
nor I_37702 (I644515,I644320,I644498);
DFFARX1 I_37703 (I644515,I3563,I643995,I643984,);
not I_37704 (I644573,I3570);
DFFARX1 I_37705 (I1145905,I3563,I644573,I644599,);
not I_37706 (I644607,I644599);
DFFARX1 I_37707 (I1145911,I3563,I644573,I644633,);
not I_37708 (I644641,I1145905);
nand I_37709 (I644658,I644641,I1145908);
not I_37710 (I644675,I644658);
nor I_37711 (I644692,I644675,I1145926);
nor I_37712 (I644709,I644607,I644692);
DFFARX1 I_37713 (I644709,I3563,I644573,I644559,);
not I_37714 (I644740,I1145926);
nand I_37715 (I644757,I644740,I644675);
and I_37716 (I644774,I644740,I1145929);
nand I_37717 (I644791,I644774,I1145908);
nor I_37718 (I644556,I644791,I644740);
and I_37719 (I644547,I644633,I644791);
not I_37720 (I644836,I644791);
nand I_37721 (I644550,I644633,I644836);
nor I_37722 (I644544,I644599,I644791);
not I_37723 (I644881,I1145914);
nor I_37724 (I644898,I644881,I1145929);
nand I_37725 (I644915,I644898,I644740);
nor I_37726 (I644553,I644658,I644915);
nor I_37727 (I644946,I644881,I1145920);
and I_37728 (I644963,I644946,I1145917);
or I_37729 (I644980,I644963,I1145923);
DFFARX1 I_37730 (I644980,I3563,I644573,I645006,);
nor I_37731 (I645014,I645006,I644757);
DFFARX1 I_37732 (I645014,I3563,I644573,I644541,);
DFFARX1 I_37733 (I645006,I3563,I644573,I644565,);
not I_37734 (I645059,I645006);
nor I_37735 (I645076,I645059,I644633);
nor I_37736 (I645093,I644898,I645076);
DFFARX1 I_37737 (I645093,I3563,I644573,I644562,);
not I_37738 (I645151,I3570);
DFFARX1 I_37739 (I46637,I3563,I645151,I645177,);
not I_37740 (I645185,I645177);
DFFARX1 I_37741 (I46640,I3563,I645151,I645211,);
not I_37742 (I645219,I46634);
nand I_37743 (I645236,I645219,I46658);
not I_37744 (I645253,I645236);
nor I_37745 (I645270,I645253,I46637);
nor I_37746 (I645287,I645185,I645270);
DFFARX1 I_37747 (I645287,I3563,I645151,I645137,);
not I_37748 (I645318,I46637);
nand I_37749 (I645335,I645318,I645253);
and I_37750 (I645352,I645318,I46652);
nand I_37751 (I645369,I645352,I46646);
nor I_37752 (I645134,I645369,I645318);
and I_37753 (I645125,I645211,I645369);
not I_37754 (I645414,I645369);
nand I_37755 (I645128,I645211,I645414);
nor I_37756 (I645122,I645177,I645369);
not I_37757 (I645459,I46655);
nor I_37758 (I645476,I645459,I46652);
nand I_37759 (I645493,I645476,I645318);
nor I_37760 (I645131,I645236,I645493);
nor I_37761 (I645524,I645459,I46634);
and I_37762 (I645541,I645524,I46643);
or I_37763 (I645558,I645541,I46649);
DFFARX1 I_37764 (I645558,I3563,I645151,I645584,);
nor I_37765 (I645592,I645584,I645335);
DFFARX1 I_37766 (I645592,I3563,I645151,I645119,);
DFFARX1 I_37767 (I645584,I3563,I645151,I645143,);
not I_37768 (I645637,I645584);
nor I_37769 (I645654,I645637,I645211);
nor I_37770 (I645671,I645476,I645654);
DFFARX1 I_37771 (I645671,I3563,I645151,I645140,);
not I_37772 (I645729,I3570);
DFFARX1 I_37773 (I400257,I3563,I645729,I645755,);
not I_37774 (I645763,I645755);
DFFARX1 I_37775 (I400272,I3563,I645729,I645789,);
not I_37776 (I645797,I400275);
nand I_37777 (I645814,I645797,I400254);
not I_37778 (I645831,I645814);
nor I_37779 (I645848,I645831,I400278);
nor I_37780 (I645865,I645763,I645848);
DFFARX1 I_37781 (I645865,I3563,I645729,I645715,);
not I_37782 (I645896,I400278);
nand I_37783 (I645913,I645896,I645831);
and I_37784 (I645930,I645896,I400260);
nand I_37785 (I645947,I645930,I400251);
nor I_37786 (I645712,I645947,I645896);
and I_37787 (I645703,I645789,I645947);
not I_37788 (I645992,I645947);
nand I_37789 (I645706,I645789,I645992);
nor I_37790 (I645700,I645755,I645947);
not I_37791 (I646037,I400251);
nor I_37792 (I646054,I646037,I400260);
nand I_37793 (I646071,I646054,I645896);
nor I_37794 (I645709,I645814,I646071);
nor I_37795 (I646102,I646037,I400266);
and I_37796 (I646119,I646102,I400269);
or I_37797 (I646136,I646119,I400263);
DFFARX1 I_37798 (I646136,I3563,I645729,I646162,);
nor I_37799 (I646170,I646162,I645913);
DFFARX1 I_37800 (I646170,I3563,I645729,I645697,);
DFFARX1 I_37801 (I646162,I3563,I645729,I645721,);
not I_37802 (I646215,I646162);
nor I_37803 (I646232,I646215,I645789);
nor I_37804 (I646249,I646054,I646232);
DFFARX1 I_37805 (I646249,I3563,I645729,I645718,);
not I_37806 (I646307,I3570);
DFFARX1 I_37807 (I163734,I3563,I646307,I646333,);
not I_37808 (I646341,I646333);
DFFARX1 I_37809 (I163713,I3563,I646307,I646367,);
not I_37810 (I646375,I163713);
nand I_37811 (I646392,I646375,I163740);
not I_37812 (I646409,I646392);
nor I_37813 (I646426,I646409,I163716);
nor I_37814 (I646443,I646341,I646426);
DFFARX1 I_37815 (I646443,I3563,I646307,I646293,);
not I_37816 (I646474,I163716);
nand I_37817 (I646491,I646474,I646409);
and I_37818 (I646508,I646474,I163737);
nand I_37819 (I646525,I646508,I163719);
nor I_37820 (I646290,I646525,I646474);
and I_37821 (I646281,I646367,I646525);
not I_37822 (I646570,I646525);
nand I_37823 (I646284,I646367,I646570);
nor I_37824 (I646278,I646333,I646525);
not I_37825 (I646615,I163722);
nor I_37826 (I646632,I646615,I163737);
nand I_37827 (I646649,I646632,I646474);
nor I_37828 (I646287,I646392,I646649);
nor I_37829 (I646680,I646615,I163728);
and I_37830 (I646697,I646680,I163725);
or I_37831 (I646714,I646697,I163731);
DFFARX1 I_37832 (I646714,I3563,I646307,I646740,);
nor I_37833 (I646748,I646740,I646491);
DFFARX1 I_37834 (I646748,I3563,I646307,I646275,);
DFFARX1 I_37835 (I646740,I3563,I646307,I646299,);
not I_37836 (I646793,I646740);
nor I_37837 (I646810,I646793,I646367);
nor I_37838 (I646827,I646632,I646810);
DFFARX1 I_37839 (I646827,I3563,I646307,I646296,);
not I_37840 (I646885,I3570);
DFFARX1 I_37841 (I1400548,I3563,I646885,I646911,);
not I_37842 (I646919,I646911);
DFFARX1 I_37843 (I1400548,I3563,I646885,I646945,);
not I_37844 (I646953,I1400572);
nand I_37845 (I646970,I646953,I1400554);
not I_37846 (I646987,I646970);
nor I_37847 (I647004,I646987,I1400569);
nor I_37848 (I647021,I646919,I647004);
DFFARX1 I_37849 (I647021,I3563,I646885,I646871,);
not I_37850 (I647052,I1400569);
nand I_37851 (I647069,I647052,I646987);
and I_37852 (I647086,I647052,I1400551);
nand I_37853 (I647103,I647086,I1400560);
nor I_37854 (I646868,I647103,I647052);
and I_37855 (I646859,I646945,I647103);
not I_37856 (I647148,I647103);
nand I_37857 (I646862,I646945,I647148);
nor I_37858 (I646856,I646911,I647103);
not I_37859 (I647193,I1400557);
nor I_37860 (I647210,I647193,I1400551);
nand I_37861 (I647227,I647210,I647052);
nor I_37862 (I646865,I646970,I647227);
nor I_37863 (I647258,I647193,I1400566);
and I_37864 (I647275,I647258,I1400575);
or I_37865 (I647292,I647275,I1400563);
DFFARX1 I_37866 (I647292,I3563,I646885,I647318,);
nor I_37867 (I647326,I647318,I647069);
DFFARX1 I_37868 (I647326,I3563,I646885,I646853,);
DFFARX1 I_37869 (I647318,I3563,I646885,I646877,);
not I_37870 (I647371,I647318);
nor I_37871 (I647388,I647371,I646945);
nor I_37872 (I647405,I647210,I647388);
DFFARX1 I_37873 (I647405,I3563,I646885,I646874,);
not I_37874 (I647463,I3570);
DFFARX1 I_37875 (I977543,I3563,I647463,I647489,);
not I_37876 (I647497,I647489);
DFFARX1 I_37877 (I977540,I3563,I647463,I647523,);
not I_37878 (I647531,I977537);
nand I_37879 (I647548,I647531,I977564);
not I_37880 (I647565,I647548);
nor I_37881 (I647582,I647565,I977552);
nor I_37882 (I647599,I647497,I647582);
DFFARX1 I_37883 (I647599,I3563,I647463,I647449,);
not I_37884 (I647630,I977552);
nand I_37885 (I647647,I647630,I647565);
and I_37886 (I647664,I647630,I977558);
nand I_37887 (I647681,I647664,I977549);
nor I_37888 (I647446,I647681,I647630);
and I_37889 (I647437,I647523,I647681);
not I_37890 (I647726,I647681);
nand I_37891 (I647440,I647523,I647726);
nor I_37892 (I647434,I647489,I647681);
not I_37893 (I647771,I977546);
nor I_37894 (I647788,I647771,I977558);
nand I_37895 (I647805,I647788,I647630);
nor I_37896 (I647443,I647548,I647805);
nor I_37897 (I647836,I647771,I977561);
and I_37898 (I647853,I647836,I977555);
or I_37899 (I647870,I647853,I977537);
DFFARX1 I_37900 (I647870,I3563,I647463,I647896,);
nor I_37901 (I647904,I647896,I647647);
DFFARX1 I_37902 (I647904,I3563,I647463,I647431,);
DFFARX1 I_37903 (I647896,I3563,I647463,I647455,);
not I_37904 (I647949,I647896);
nor I_37905 (I647966,I647949,I647523);
nor I_37906 (I647983,I647788,I647966);
DFFARX1 I_37907 (I647983,I3563,I647463,I647452,);
not I_37908 (I648041,I3570);
DFFARX1 I_37909 (I511630,I3563,I648041,I648067,);
not I_37910 (I648075,I648067);
DFFARX1 I_37911 (I511642,I3563,I648041,I648101,);
not I_37912 (I648109,I511618);
nand I_37913 (I648126,I648109,I511645);
not I_37914 (I648143,I648126);
nor I_37915 (I648160,I648143,I511633);
nor I_37916 (I648177,I648075,I648160);
DFFARX1 I_37917 (I648177,I3563,I648041,I648027,);
not I_37918 (I648208,I511633);
nand I_37919 (I648225,I648208,I648143);
and I_37920 (I648242,I648208,I511618);
nand I_37921 (I648259,I648242,I511621);
nor I_37922 (I648024,I648259,I648208);
and I_37923 (I648015,I648101,I648259);
not I_37924 (I648304,I648259);
nand I_37925 (I648018,I648101,I648304);
nor I_37926 (I648012,I648067,I648259);
not I_37927 (I648349,I511627);
nor I_37928 (I648366,I648349,I511618);
nand I_37929 (I648383,I648366,I648208);
nor I_37930 (I648021,I648126,I648383);
nor I_37931 (I648414,I648349,I511636);
and I_37932 (I648431,I648414,I511624);
or I_37933 (I648448,I648431,I511639);
DFFARX1 I_37934 (I648448,I3563,I648041,I648474,);
nor I_37935 (I648482,I648474,I648225);
DFFARX1 I_37936 (I648482,I3563,I648041,I648009,);
DFFARX1 I_37937 (I648474,I3563,I648041,I648033,);
not I_37938 (I648527,I648474);
nor I_37939 (I648544,I648527,I648101);
nor I_37940 (I648561,I648366,I648544);
DFFARX1 I_37941 (I648561,I3563,I648041,I648030,);
not I_37942 (I648619,I3570);
DFFARX1 I_37943 (I80386,I3563,I648619,I648645,);
not I_37944 (I648653,I648645);
DFFARX1 I_37945 (I80365,I3563,I648619,I648679,);
not I_37946 (I648687,I80362);
nand I_37947 (I648704,I648687,I80377);
not I_37948 (I648721,I648704);
nor I_37949 (I648738,I648721,I80365);
nor I_37950 (I648755,I648653,I648738);
DFFARX1 I_37951 (I648755,I3563,I648619,I648605,);
not I_37952 (I648786,I80365);
nand I_37953 (I648803,I648786,I648721);
and I_37954 (I648820,I648786,I80368);
nand I_37955 (I648837,I648820,I80383);
nor I_37956 (I648602,I648837,I648786);
and I_37957 (I648593,I648679,I648837);
not I_37958 (I648882,I648837);
nand I_37959 (I648596,I648679,I648882);
nor I_37960 (I648590,I648645,I648837);
not I_37961 (I648927,I80374);
nor I_37962 (I648944,I648927,I80368);
nand I_37963 (I648961,I648944,I648786);
nor I_37964 (I648599,I648704,I648961);
nor I_37965 (I648992,I648927,I80362);
and I_37966 (I649009,I648992,I80371);
or I_37967 (I649026,I649009,I80380);
DFFARX1 I_37968 (I649026,I3563,I648619,I649052,);
nor I_37969 (I649060,I649052,I648803);
DFFARX1 I_37970 (I649060,I3563,I648619,I648587,);
DFFARX1 I_37971 (I649052,I3563,I648619,I648611,);
not I_37972 (I649105,I649052);
nor I_37973 (I649122,I649105,I648679);
nor I_37974 (I649139,I648944,I649122);
DFFARX1 I_37975 (I649139,I3563,I648619,I648608,);
not I_37976 (I649197,I3570);
DFFARX1 I_37977 (I458318,I3563,I649197,I649223,);
not I_37978 (I649231,I649223);
DFFARX1 I_37979 (I458330,I3563,I649197,I649257,);
not I_37980 (I649265,I458306);
nand I_37981 (I649282,I649265,I458333);
not I_37982 (I649299,I649282);
nor I_37983 (I649316,I649299,I458321);
nor I_37984 (I649333,I649231,I649316);
DFFARX1 I_37985 (I649333,I3563,I649197,I649183,);
not I_37986 (I649364,I458321);
nand I_37987 (I649381,I649364,I649299);
and I_37988 (I649398,I649364,I458306);
nand I_37989 (I649415,I649398,I458309);
nor I_37990 (I649180,I649415,I649364);
and I_37991 (I649171,I649257,I649415);
not I_37992 (I649460,I649415);
nand I_37993 (I649174,I649257,I649460);
nor I_37994 (I649168,I649223,I649415);
not I_37995 (I649505,I458315);
nor I_37996 (I649522,I649505,I458306);
nand I_37997 (I649539,I649522,I649364);
nor I_37998 (I649177,I649282,I649539);
nor I_37999 (I649570,I649505,I458324);
and I_38000 (I649587,I649570,I458312);
or I_38001 (I649604,I649587,I458327);
DFFARX1 I_38002 (I649604,I3563,I649197,I649630,);
nor I_38003 (I649638,I649630,I649381);
DFFARX1 I_38004 (I649638,I3563,I649197,I649165,);
DFFARX1 I_38005 (I649630,I3563,I649197,I649189,);
not I_38006 (I649683,I649630);
nor I_38007 (I649700,I649683,I649257);
nor I_38008 (I649717,I649522,I649700);
DFFARX1 I_38009 (I649717,I3563,I649197,I649186,);
not I_38010 (I649775,I3570);
DFFARX1 I_38011 (I886423,I3563,I649775,I649801,);
not I_38012 (I649809,I649801);
DFFARX1 I_38013 (I886423,I3563,I649775,I649835,);
not I_38014 (I649843,I886420);
nand I_38015 (I649860,I649843,I886435);
not I_38016 (I649877,I649860);
nor I_38017 (I649894,I649877,I886429);
nor I_38018 (I649911,I649809,I649894);
DFFARX1 I_38019 (I649911,I3563,I649775,I649761,);
not I_38020 (I649942,I886429);
nand I_38021 (I649959,I649942,I649877);
and I_38022 (I649976,I649942,I886426);
nand I_38023 (I649993,I649976,I886417);
nor I_38024 (I649758,I649993,I649942);
and I_38025 (I649749,I649835,I649993);
not I_38026 (I650038,I649993);
nand I_38027 (I649752,I649835,I650038);
nor I_38028 (I649746,I649801,I649993);
not I_38029 (I650083,I886438);
nor I_38030 (I650100,I650083,I886426);
nand I_38031 (I650117,I650100,I649942);
nor I_38032 (I649755,I649860,I650117);
nor I_38033 (I650148,I650083,I886417);
and I_38034 (I650165,I650148,I886420);
or I_38035 (I650182,I650165,I886432);
DFFARX1 I_38036 (I650182,I3563,I649775,I650208,);
nor I_38037 (I650216,I650208,I649959);
DFFARX1 I_38038 (I650216,I3563,I649775,I649743,);
DFFARX1 I_38039 (I650208,I3563,I649775,I649767,);
not I_38040 (I650261,I650208);
nor I_38041 (I650278,I650261,I649835);
nor I_38042 (I650295,I650100,I650278);
DFFARX1 I_38043 (I650295,I3563,I649775,I649764,);
not I_38044 (I650353,I3570);
DFFARX1 I_38045 (I99358,I3563,I650353,I650379,);
not I_38046 (I650387,I650379);
DFFARX1 I_38047 (I99337,I3563,I650353,I650413,);
not I_38048 (I650421,I99334);
nand I_38049 (I650438,I650421,I99349);
not I_38050 (I650455,I650438);
nor I_38051 (I650472,I650455,I99337);
nor I_38052 (I650489,I650387,I650472);
DFFARX1 I_38053 (I650489,I3563,I650353,I650339,);
not I_38054 (I650520,I99337);
nand I_38055 (I650537,I650520,I650455);
and I_38056 (I650554,I650520,I99340);
nand I_38057 (I650571,I650554,I99355);
nor I_38058 (I650336,I650571,I650520);
and I_38059 (I650327,I650413,I650571);
not I_38060 (I650616,I650571);
nand I_38061 (I650330,I650413,I650616);
nor I_38062 (I650324,I650379,I650571);
not I_38063 (I650661,I99346);
nor I_38064 (I650678,I650661,I99340);
nand I_38065 (I650695,I650678,I650520);
nor I_38066 (I650333,I650438,I650695);
nor I_38067 (I650726,I650661,I99334);
and I_38068 (I650743,I650726,I99343);
or I_38069 (I650760,I650743,I99352);
DFFARX1 I_38070 (I650760,I3563,I650353,I650786,);
nor I_38071 (I650794,I650786,I650537);
DFFARX1 I_38072 (I650794,I3563,I650353,I650321,);
DFFARX1 I_38073 (I650786,I3563,I650353,I650345,);
not I_38074 (I650839,I650786);
nor I_38075 (I650856,I650839,I650413);
nor I_38076 (I650873,I650678,I650856);
DFFARX1 I_38077 (I650873,I3563,I650353,I650342,);
not I_38078 (I650931,I3570);
DFFARX1 I_38079 (I31881,I3563,I650931,I650957,);
not I_38080 (I650965,I650957);
DFFARX1 I_38081 (I31884,I3563,I650931,I650991,);
not I_38082 (I650999,I31878);
nand I_38083 (I651016,I650999,I31902);
not I_38084 (I651033,I651016);
nor I_38085 (I651050,I651033,I31881);
nor I_38086 (I651067,I650965,I651050);
DFFARX1 I_38087 (I651067,I3563,I650931,I650917,);
not I_38088 (I651098,I31881);
nand I_38089 (I651115,I651098,I651033);
and I_38090 (I651132,I651098,I31896);
nand I_38091 (I651149,I651132,I31890);
nor I_38092 (I650914,I651149,I651098);
and I_38093 (I650905,I650991,I651149);
not I_38094 (I651194,I651149);
nand I_38095 (I650908,I650991,I651194);
nor I_38096 (I650902,I650957,I651149);
not I_38097 (I651239,I31899);
nor I_38098 (I651256,I651239,I31896);
nand I_38099 (I651273,I651256,I651098);
nor I_38100 (I650911,I651016,I651273);
nor I_38101 (I651304,I651239,I31878);
and I_38102 (I651321,I651304,I31887);
or I_38103 (I651338,I651321,I31893);
DFFARX1 I_38104 (I651338,I3563,I650931,I651364,);
nor I_38105 (I651372,I651364,I651115);
DFFARX1 I_38106 (I651372,I3563,I650931,I650899,);
DFFARX1 I_38107 (I651364,I3563,I650931,I650923,);
not I_38108 (I651417,I651364);
nor I_38109 (I651434,I651417,I650991);
nor I_38110 (I651451,I651256,I651434);
DFFARX1 I_38111 (I651451,I3563,I650931,I650920,);
not I_38112 (I651509,I3570);
DFFARX1 I_38113 (I445262,I3563,I651509,I651535,);
not I_38114 (I651543,I651535);
DFFARX1 I_38115 (I445274,I3563,I651509,I651569,);
not I_38116 (I651577,I445250);
nand I_38117 (I651594,I651577,I445277);
not I_38118 (I651611,I651594);
nor I_38119 (I651628,I651611,I445265);
nor I_38120 (I651645,I651543,I651628);
DFFARX1 I_38121 (I651645,I3563,I651509,I651495,);
not I_38122 (I651676,I445265);
nand I_38123 (I651693,I651676,I651611);
and I_38124 (I651710,I651676,I445250);
nand I_38125 (I651727,I651710,I445253);
nor I_38126 (I651492,I651727,I651676);
and I_38127 (I651483,I651569,I651727);
not I_38128 (I651772,I651727);
nand I_38129 (I651486,I651569,I651772);
nor I_38130 (I651480,I651535,I651727);
not I_38131 (I651817,I445259);
nor I_38132 (I651834,I651817,I445250);
nand I_38133 (I651851,I651834,I651676);
nor I_38134 (I651489,I651594,I651851);
nor I_38135 (I651882,I651817,I445268);
and I_38136 (I651899,I651882,I445256);
or I_38137 (I651916,I651899,I445271);
DFFARX1 I_38138 (I651916,I3563,I651509,I651942,);
nor I_38139 (I651950,I651942,I651693);
DFFARX1 I_38140 (I651950,I3563,I651509,I651477,);
DFFARX1 I_38141 (I651942,I3563,I651509,I651501,);
not I_38142 (I651995,I651942);
nor I_38143 (I652012,I651995,I651569);
nor I_38144 (I652029,I651834,I652012);
DFFARX1 I_38145 (I652029,I3563,I651509,I651498,);
not I_38146 (I652087,I3570);
DFFARX1 I_38147 (I269638,I3563,I652087,I652113,);
not I_38148 (I652121,I652113);
DFFARX1 I_38149 (I269623,I3563,I652087,I652147,);
not I_38150 (I652155,I269641);
nand I_38151 (I652172,I652155,I269626);
not I_38152 (I652189,I652172);
nor I_38153 (I652206,I652189,I269623);
nor I_38154 (I652223,I652121,I652206);
DFFARX1 I_38155 (I652223,I3563,I652087,I652073,);
not I_38156 (I652254,I269623);
nand I_38157 (I652271,I652254,I652189);
and I_38158 (I652288,I652254,I269626);
nand I_38159 (I652305,I652288,I269647);
nor I_38160 (I652070,I652305,I652254);
and I_38161 (I652061,I652147,I652305);
not I_38162 (I652350,I652305);
nand I_38163 (I652064,I652147,I652350);
nor I_38164 (I652058,I652113,I652305);
not I_38165 (I652395,I269635);
nor I_38166 (I652412,I652395,I269626);
nand I_38167 (I652429,I652412,I652254);
nor I_38168 (I652067,I652172,I652429);
nor I_38169 (I652460,I652395,I269629);
and I_38170 (I652477,I652460,I269644);
or I_38171 (I652494,I652477,I269632);
DFFARX1 I_38172 (I652494,I3563,I652087,I652520,);
nor I_38173 (I652528,I652520,I652271);
DFFARX1 I_38174 (I652528,I3563,I652087,I652055,);
DFFARX1 I_38175 (I652520,I3563,I652087,I652079,);
not I_38176 (I652573,I652520);
nor I_38177 (I652590,I652573,I652147);
nor I_38178 (I652607,I652412,I652590);
DFFARX1 I_38179 (I652607,I3563,I652087,I652076,);
not I_38180 (I652665,I3570);
DFFARX1 I_38181 (I408689,I3563,I652665,I652691,);
not I_38182 (I652699,I652691);
DFFARX1 I_38183 (I408704,I3563,I652665,I652725,);
not I_38184 (I652733,I408707);
nand I_38185 (I652750,I652733,I408686);
not I_38186 (I652767,I652750);
nor I_38187 (I652784,I652767,I408710);
nor I_38188 (I652801,I652699,I652784);
DFFARX1 I_38189 (I652801,I3563,I652665,I652651,);
not I_38190 (I652832,I408710);
nand I_38191 (I652849,I652832,I652767);
and I_38192 (I652866,I652832,I408692);
nand I_38193 (I652883,I652866,I408683);
nor I_38194 (I652648,I652883,I652832);
and I_38195 (I652639,I652725,I652883);
not I_38196 (I652928,I652883);
nand I_38197 (I652642,I652725,I652928);
nor I_38198 (I652636,I652691,I652883);
not I_38199 (I652973,I408683);
nor I_38200 (I652990,I652973,I408692);
nand I_38201 (I653007,I652990,I652832);
nor I_38202 (I652645,I652750,I653007);
nor I_38203 (I653038,I652973,I408698);
and I_38204 (I653055,I653038,I408701);
or I_38205 (I653072,I653055,I408695);
DFFARX1 I_38206 (I653072,I3563,I652665,I653098,);
nor I_38207 (I653106,I653098,I652849);
DFFARX1 I_38208 (I653106,I3563,I652665,I652633,);
DFFARX1 I_38209 (I653098,I3563,I652665,I652657,);
not I_38210 (I653151,I653098);
nor I_38211 (I653168,I653151,I652725);
nor I_38212 (I653185,I652990,I653168);
DFFARX1 I_38213 (I653185,I3563,I652665,I652654,);
not I_38214 (I653243,I3570);
DFFARX1 I_38215 (I722571,I3563,I653243,I653269,);
not I_38216 (I653277,I653269);
DFFARX1 I_38217 (I722583,I3563,I653243,I653303,);
not I_38218 (I653311,I722574);
nand I_38219 (I653328,I653311,I722577);
not I_38220 (I653345,I653328);
nor I_38221 (I653362,I653345,I722580);
nor I_38222 (I653379,I653277,I653362);
DFFARX1 I_38223 (I653379,I3563,I653243,I653229,);
not I_38224 (I653410,I722580);
nand I_38225 (I653427,I653410,I653345);
and I_38226 (I653444,I653410,I722574);
nand I_38227 (I653461,I653444,I722586);
nor I_38228 (I653226,I653461,I653410);
and I_38229 (I653217,I653303,I653461);
not I_38230 (I653506,I653461);
nand I_38231 (I653220,I653303,I653506);
nor I_38232 (I653214,I653269,I653461);
not I_38233 (I653551,I722592);
nor I_38234 (I653568,I653551,I722574);
nand I_38235 (I653585,I653568,I653410);
nor I_38236 (I653223,I653328,I653585);
nor I_38237 (I653616,I653551,I722571);
and I_38238 (I653633,I653616,I722589);
or I_38239 (I653650,I653633,I722595);
DFFARX1 I_38240 (I653650,I3563,I653243,I653676,);
nor I_38241 (I653684,I653676,I653427);
DFFARX1 I_38242 (I653684,I3563,I653243,I653211,);
DFFARX1 I_38243 (I653676,I3563,I653243,I653235,);
not I_38244 (I653729,I653676);
nor I_38245 (I653746,I653729,I653303);
nor I_38246 (I653763,I653568,I653746);
DFFARX1 I_38247 (I653763,I3563,I653243,I653232,);
not I_38248 (I653821,I3570);
DFFARX1 I_38249 (I56123,I3563,I653821,I653847,);
not I_38250 (I653855,I653847);
DFFARX1 I_38251 (I56126,I3563,I653821,I653881,);
not I_38252 (I653889,I56120);
nand I_38253 (I653906,I653889,I56144);
not I_38254 (I653923,I653906);
nor I_38255 (I653940,I653923,I56123);
nor I_38256 (I653957,I653855,I653940);
DFFARX1 I_38257 (I653957,I3563,I653821,I653807,);
not I_38258 (I653988,I56123);
nand I_38259 (I654005,I653988,I653923);
and I_38260 (I654022,I653988,I56138);
nand I_38261 (I654039,I654022,I56132);
nor I_38262 (I653804,I654039,I653988);
and I_38263 (I653795,I653881,I654039);
not I_38264 (I654084,I654039);
nand I_38265 (I653798,I653881,I654084);
nor I_38266 (I653792,I653847,I654039);
not I_38267 (I654129,I56141);
nor I_38268 (I654146,I654129,I56138);
nand I_38269 (I654163,I654146,I653988);
nor I_38270 (I653801,I653906,I654163);
nor I_38271 (I654194,I654129,I56120);
and I_38272 (I654211,I654194,I56129);
or I_38273 (I654228,I654211,I56135);
DFFARX1 I_38274 (I654228,I3563,I653821,I654254,);
nor I_38275 (I654262,I654254,I654005);
DFFARX1 I_38276 (I654262,I3563,I653821,I653789,);
DFFARX1 I_38277 (I654254,I3563,I653821,I653813,);
not I_38278 (I654307,I654254);
nor I_38279 (I654324,I654307,I653881);
nor I_38280 (I654341,I654146,I654324);
DFFARX1 I_38281 (I654341,I3563,I653821,I653810,);
not I_38282 (I654399,I3570);
DFFARX1 I_38283 (I18706,I3563,I654399,I654425,);
not I_38284 (I654433,I654425);
DFFARX1 I_38285 (I18709,I3563,I654399,I654459,);
not I_38286 (I654467,I18703);
nand I_38287 (I654484,I654467,I18727);
not I_38288 (I654501,I654484);
nor I_38289 (I654518,I654501,I18706);
nor I_38290 (I654535,I654433,I654518);
DFFARX1 I_38291 (I654535,I3563,I654399,I654385,);
not I_38292 (I654566,I18706);
nand I_38293 (I654583,I654566,I654501);
and I_38294 (I654600,I654566,I18721);
nand I_38295 (I654617,I654600,I18715);
nor I_38296 (I654382,I654617,I654566);
and I_38297 (I654373,I654459,I654617);
not I_38298 (I654662,I654617);
nand I_38299 (I654376,I654459,I654662);
nor I_38300 (I654370,I654425,I654617);
not I_38301 (I654707,I18724);
nor I_38302 (I654724,I654707,I18721);
nand I_38303 (I654741,I654724,I654566);
nor I_38304 (I654379,I654484,I654741);
nor I_38305 (I654772,I654707,I18703);
and I_38306 (I654789,I654772,I18712);
or I_38307 (I654806,I654789,I18718);
DFFARX1 I_38308 (I654806,I3563,I654399,I654832,);
nor I_38309 (I654840,I654832,I654583);
DFFARX1 I_38310 (I654840,I3563,I654399,I654367,);
DFFARX1 I_38311 (I654832,I3563,I654399,I654391,);
not I_38312 (I654885,I654832);
nor I_38313 (I654902,I654885,I654459);
nor I_38314 (I654919,I654724,I654902);
DFFARX1 I_38315 (I654919,I3563,I654399,I654388,);
not I_38316 (I654977,I3570);
DFFARX1 I_38317 (I856911,I3563,I654977,I655003,);
not I_38318 (I655011,I655003);
DFFARX1 I_38319 (I856911,I3563,I654977,I655037,);
not I_38320 (I655045,I856908);
nand I_38321 (I655062,I655045,I856923);
not I_38322 (I655079,I655062);
nor I_38323 (I655096,I655079,I856917);
nor I_38324 (I655113,I655011,I655096);
DFFARX1 I_38325 (I655113,I3563,I654977,I654963,);
not I_38326 (I655144,I856917);
nand I_38327 (I655161,I655144,I655079);
and I_38328 (I655178,I655144,I856914);
nand I_38329 (I655195,I655178,I856905);
nor I_38330 (I654960,I655195,I655144);
and I_38331 (I654951,I655037,I655195);
not I_38332 (I655240,I655195);
nand I_38333 (I654954,I655037,I655240);
nor I_38334 (I654948,I655003,I655195);
not I_38335 (I655285,I856926);
nor I_38336 (I655302,I655285,I856914);
nand I_38337 (I655319,I655302,I655144);
nor I_38338 (I654957,I655062,I655319);
nor I_38339 (I655350,I655285,I856905);
and I_38340 (I655367,I655350,I856908);
or I_38341 (I655384,I655367,I856920);
DFFARX1 I_38342 (I655384,I3563,I654977,I655410,);
nor I_38343 (I655418,I655410,I655161);
DFFARX1 I_38344 (I655418,I3563,I654977,I654945,);
DFFARX1 I_38345 (I655410,I3563,I654977,I654969,);
not I_38346 (I655463,I655410);
nor I_38347 (I655480,I655463,I655037);
nor I_38348 (I655497,I655302,I655480);
DFFARX1 I_38349 (I655497,I3563,I654977,I654966,);
not I_38350 (I655555,I3570);
DFFARX1 I_38351 (I286893,I3563,I655555,I655581,);
not I_38352 (I655589,I655581);
DFFARX1 I_38353 (I286878,I3563,I655555,I655615,);
not I_38354 (I655623,I286896);
nand I_38355 (I655640,I655623,I286881);
not I_38356 (I655657,I655640);
nor I_38357 (I655674,I655657,I286878);
nor I_38358 (I655691,I655589,I655674);
DFFARX1 I_38359 (I655691,I3563,I655555,I655541,);
not I_38360 (I655722,I286878);
nand I_38361 (I655739,I655722,I655657);
and I_38362 (I655756,I655722,I286881);
nand I_38363 (I655773,I655756,I286902);
nor I_38364 (I655538,I655773,I655722);
and I_38365 (I655529,I655615,I655773);
not I_38366 (I655818,I655773);
nand I_38367 (I655532,I655615,I655818);
nor I_38368 (I655526,I655581,I655773);
not I_38369 (I655863,I286890);
nor I_38370 (I655880,I655863,I286881);
nand I_38371 (I655897,I655880,I655722);
nor I_38372 (I655535,I655640,I655897);
nor I_38373 (I655928,I655863,I286884);
and I_38374 (I655945,I655928,I286899);
or I_38375 (I655962,I655945,I286887);
DFFARX1 I_38376 (I655962,I3563,I655555,I655988,);
nor I_38377 (I655996,I655988,I655739);
DFFARX1 I_38378 (I655996,I3563,I655555,I655523,);
DFFARX1 I_38379 (I655988,I3563,I655555,I655547,);
not I_38380 (I656041,I655988);
nor I_38381 (I656058,I656041,I655615);
nor I_38382 (I656075,I655880,I656058);
DFFARX1 I_38383 (I656075,I3563,I655555,I655544,);
not I_38384 (I656133,I3570);
DFFARX1 I_38385 (I558439,I3563,I656133,I656159,);
not I_38386 (I656167,I656159);
DFFARX1 I_38387 (I558451,I3563,I656133,I656193,);
not I_38388 (I656201,I558457);
nand I_38389 (I656218,I656201,I558448);
not I_38390 (I656235,I656218);
nor I_38391 (I656252,I656235,I558454);
nor I_38392 (I656269,I656167,I656252);
DFFARX1 I_38393 (I656269,I3563,I656133,I656119,);
not I_38394 (I656300,I558454);
nand I_38395 (I656317,I656300,I656235);
and I_38396 (I656334,I656300,I558445);
nand I_38397 (I656351,I656334,I558436);
nor I_38398 (I656116,I656351,I656300);
and I_38399 (I656107,I656193,I656351);
not I_38400 (I656396,I656351);
nand I_38401 (I656110,I656193,I656396);
nor I_38402 (I656104,I656159,I656351);
not I_38403 (I656441,I558442);
nor I_38404 (I656458,I656441,I558445);
nand I_38405 (I656475,I656458,I656300);
nor I_38406 (I656113,I656218,I656475);
nor I_38407 (I656506,I656441,I558439);
and I_38408 (I656523,I656506,I558436);
or I_38409 (I656540,I656523,I558460);
DFFARX1 I_38410 (I656540,I3563,I656133,I656566,);
nor I_38411 (I656574,I656566,I656317);
DFFARX1 I_38412 (I656574,I3563,I656133,I656101,);
DFFARX1 I_38413 (I656566,I3563,I656133,I656125,);
not I_38414 (I656619,I656566);
nor I_38415 (I656636,I656619,I656193);
nor I_38416 (I656653,I656458,I656636);
DFFARX1 I_38417 (I656653,I3563,I656133,I656122,);
not I_38418 (I656711,I3570);
DFFARX1 I_38419 (I296965,I3563,I656711,I656737,);
not I_38420 (I656745,I656737);
DFFARX1 I_38421 (I296980,I3563,I656711,I656771,);
not I_38422 (I656779,I296983);
nand I_38423 (I656796,I656779,I296962);
not I_38424 (I656813,I656796);
nor I_38425 (I656830,I656813,I296986);
nor I_38426 (I656847,I656745,I656830);
DFFARX1 I_38427 (I656847,I3563,I656711,I656697,);
not I_38428 (I656878,I296986);
nand I_38429 (I656895,I656878,I656813);
and I_38430 (I656912,I656878,I296968);
nand I_38431 (I656929,I656912,I296959);
nor I_38432 (I656694,I656929,I656878);
and I_38433 (I656685,I656771,I656929);
not I_38434 (I656974,I656929);
nand I_38435 (I656688,I656771,I656974);
nor I_38436 (I656682,I656737,I656929);
not I_38437 (I657019,I296959);
nor I_38438 (I657036,I657019,I296968);
nand I_38439 (I657053,I657036,I656878);
nor I_38440 (I656691,I656796,I657053);
nor I_38441 (I657084,I657019,I296974);
and I_38442 (I657101,I657084,I296977);
or I_38443 (I657118,I657101,I296971);
DFFARX1 I_38444 (I657118,I3563,I656711,I657144,);
nor I_38445 (I657152,I657144,I656895);
DFFARX1 I_38446 (I657152,I3563,I656711,I656679,);
DFFARX1 I_38447 (I657144,I3563,I656711,I656703,);
not I_38448 (I657197,I657144);
nor I_38449 (I657214,I657197,I656771);
nor I_38450 (I657231,I657036,I657214);
DFFARX1 I_38451 (I657231,I3563,I656711,I656700,);
not I_38452 (I657289,I3570);
DFFARX1 I_38453 (I745691,I3563,I657289,I657315,);
not I_38454 (I657323,I657315);
DFFARX1 I_38455 (I745703,I3563,I657289,I657349,);
not I_38456 (I657357,I745694);
nand I_38457 (I657374,I657357,I745697);
not I_38458 (I657391,I657374);
nor I_38459 (I657408,I657391,I745700);
nor I_38460 (I657425,I657323,I657408);
DFFARX1 I_38461 (I657425,I3563,I657289,I657275,);
not I_38462 (I657456,I745700);
nand I_38463 (I657473,I657456,I657391);
and I_38464 (I657490,I657456,I745694);
nand I_38465 (I657507,I657490,I745706);
nor I_38466 (I657272,I657507,I657456);
and I_38467 (I657263,I657349,I657507);
not I_38468 (I657552,I657507);
nand I_38469 (I657266,I657349,I657552);
nor I_38470 (I657260,I657315,I657507);
not I_38471 (I657597,I745712);
nor I_38472 (I657614,I657597,I745694);
nand I_38473 (I657631,I657614,I657456);
nor I_38474 (I657269,I657374,I657631);
nor I_38475 (I657662,I657597,I745691);
and I_38476 (I657679,I657662,I745709);
or I_38477 (I657696,I657679,I745715);
DFFARX1 I_38478 (I657696,I3563,I657289,I657722,);
nor I_38479 (I657730,I657722,I657473);
DFFARX1 I_38480 (I657730,I3563,I657289,I657257,);
DFFARX1 I_38481 (I657722,I3563,I657289,I657281,);
not I_38482 (I657775,I657722);
nor I_38483 (I657792,I657775,I657349);
nor I_38484 (I657809,I657614,I657792);
DFFARX1 I_38485 (I657809,I3563,I657289,I657278,);
not I_38486 (I657867,I3570);
DFFARX1 I_38487 (I192288,I3563,I657867,I657893,);
not I_38488 (I657901,I657893);
DFFARX1 I_38489 (I192273,I3563,I657867,I657927,);
not I_38490 (I657935,I192291);
nand I_38491 (I657952,I657935,I192276);
not I_38492 (I657969,I657952);
nor I_38493 (I657986,I657969,I192273);
nor I_38494 (I658003,I657901,I657986);
DFFARX1 I_38495 (I658003,I3563,I657867,I657853,);
not I_38496 (I658034,I192273);
nand I_38497 (I658051,I658034,I657969);
and I_38498 (I658068,I658034,I192276);
nand I_38499 (I658085,I658068,I192297);
nor I_38500 (I657850,I658085,I658034);
and I_38501 (I657841,I657927,I658085);
not I_38502 (I658130,I658085);
nand I_38503 (I657844,I657927,I658130);
nor I_38504 (I657838,I657893,I658085);
not I_38505 (I658175,I192285);
nor I_38506 (I658192,I658175,I192276);
nand I_38507 (I658209,I658192,I658034);
nor I_38508 (I657847,I657952,I658209);
nor I_38509 (I658240,I658175,I192279);
and I_38510 (I658257,I658240,I192294);
or I_38511 (I658274,I658257,I192282);
DFFARX1 I_38512 (I658274,I3563,I657867,I658300,);
nor I_38513 (I658308,I658300,I658051);
DFFARX1 I_38514 (I658308,I3563,I657867,I657835,);
DFFARX1 I_38515 (I658300,I3563,I657867,I657859,);
not I_38516 (I658353,I658300);
nor I_38517 (I658370,I658353,I657927);
nor I_38518 (I658387,I658192,I658370);
DFFARX1 I_38519 (I658387,I3563,I657867,I657856,);
not I_38520 (I658445,I3570);
DFFARX1 I_38521 (I1247497,I3563,I658445,I658471,);
not I_38522 (I658479,I658471);
nand I_38523 (I658496,I1247500,I1247509);
and I_38524 (I658513,I658496,I1247512);
DFFARX1 I_38525 (I658513,I3563,I658445,I658539,);
not I_38526 (I658547,I1247521);
DFFARX1 I_38527 (I1247503,I3563,I658445,I658573,);
not I_38528 (I658581,I658573);
nor I_38529 (I658598,I658581,I658479);
and I_38530 (I658615,I658598,I1247521);
nor I_38531 (I658632,I658581,I658547);
nor I_38532 (I658428,I658539,I658632);
DFFARX1 I_38533 (I1247500,I3563,I658445,I658672,);
nor I_38534 (I658680,I658672,I658539);
not I_38535 (I658697,I658680);
not I_38536 (I658714,I658672);
nor I_38537 (I658731,I658714,I658615);
DFFARX1 I_38538 (I658731,I3563,I658445,I658431,);
nand I_38539 (I658762,I1247518,I1247497);
and I_38540 (I658779,I658762,I1247515);
DFFARX1 I_38541 (I658779,I3563,I658445,I658805,);
nor I_38542 (I658813,I658805,I658672);
DFFARX1 I_38543 (I658813,I3563,I658445,I658413,);
nand I_38544 (I658844,I658805,I658714);
nand I_38545 (I658422,I658697,I658844);
not I_38546 (I658875,I658805);
nor I_38547 (I658892,I658875,I658615);
DFFARX1 I_38548 (I658892,I3563,I658445,I658434,);
nor I_38549 (I658923,I1247506,I1247497);
or I_38550 (I658425,I658672,I658923);
nor I_38551 (I658416,I658805,I658923);
or I_38552 (I658419,I658539,I658923);
DFFARX1 I_38553 (I658923,I3563,I658445,I658437,);
not I_38554 (I659023,I3570);
DFFARX1 I_38555 (I391316,I3563,I659023,I659049,);
not I_38556 (I659057,I659049);
nand I_38557 (I659074,I391319,I391295);
and I_38558 (I659091,I659074,I391292);
DFFARX1 I_38559 (I659091,I3563,I659023,I659117,);
not I_38560 (I659125,I391298);
DFFARX1 I_38561 (I391292,I3563,I659023,I659151,);
not I_38562 (I659159,I659151);
nor I_38563 (I659176,I659159,I659057);
and I_38564 (I659193,I659176,I391298);
nor I_38565 (I659210,I659159,I659125);
nor I_38566 (I659006,I659117,I659210);
DFFARX1 I_38567 (I391301,I3563,I659023,I659250,);
nor I_38568 (I659258,I659250,I659117);
not I_38569 (I659275,I659258);
not I_38570 (I659292,I659250);
nor I_38571 (I659309,I659292,I659193);
DFFARX1 I_38572 (I659309,I3563,I659023,I659009,);
nand I_38573 (I659340,I391304,I391313);
and I_38574 (I659357,I659340,I391310);
DFFARX1 I_38575 (I659357,I3563,I659023,I659383,);
nor I_38576 (I659391,I659383,I659250);
DFFARX1 I_38577 (I659391,I3563,I659023,I658991,);
nand I_38578 (I659422,I659383,I659292);
nand I_38579 (I659000,I659275,I659422);
not I_38580 (I659453,I659383);
nor I_38581 (I659470,I659453,I659193);
DFFARX1 I_38582 (I659470,I3563,I659023,I659012,);
nor I_38583 (I659501,I391307,I391313);
or I_38584 (I659003,I659250,I659501);
nor I_38585 (I658994,I659383,I659501);
or I_38586 (I658997,I659117,I659501);
DFFARX1 I_38587 (I659501,I3563,I659023,I659015,);
not I_38588 (I659601,I3570);
DFFARX1 I_38589 (I831097,I3563,I659601,I659627,);
not I_38590 (I659635,I659627);
nand I_38591 (I659652,I831085,I831103);
and I_38592 (I659669,I659652,I831100);
DFFARX1 I_38593 (I659669,I3563,I659601,I659695,);
not I_38594 (I659703,I831091);
DFFARX1 I_38595 (I831088,I3563,I659601,I659729,);
not I_38596 (I659737,I659729);
nor I_38597 (I659754,I659737,I659635);
and I_38598 (I659771,I659754,I831091);
nor I_38599 (I659788,I659737,I659703);
nor I_38600 (I659584,I659695,I659788);
DFFARX1 I_38601 (I831082,I3563,I659601,I659828,);
nor I_38602 (I659836,I659828,I659695);
not I_38603 (I659853,I659836);
not I_38604 (I659870,I659828);
nor I_38605 (I659887,I659870,I659771);
DFFARX1 I_38606 (I659887,I3563,I659601,I659587,);
nand I_38607 (I659918,I831082,I831085);
and I_38608 (I659935,I659918,I831088);
DFFARX1 I_38609 (I659935,I3563,I659601,I659961,);
nor I_38610 (I659969,I659961,I659828);
DFFARX1 I_38611 (I659969,I3563,I659601,I659569,);
nand I_38612 (I660000,I659961,I659870);
nand I_38613 (I659578,I659853,I660000);
not I_38614 (I660031,I659961);
nor I_38615 (I660048,I660031,I659771);
DFFARX1 I_38616 (I660048,I3563,I659601,I659590,);
nor I_38617 (I660079,I831094,I831085);
or I_38618 (I659581,I659828,I660079);
nor I_38619 (I659572,I659961,I660079);
or I_38620 (I659575,I659695,I660079);
DFFARX1 I_38621 (I660079,I3563,I659601,I659593,);
not I_38622 (I660179,I3570);
DFFARX1 I_38623 (I642229,I3563,I660179,I660205,);
not I_38624 (I660213,I660205);
nand I_38625 (I660230,I642238,I642247);
and I_38626 (I660247,I660230,I642253);
DFFARX1 I_38627 (I660247,I3563,I660179,I660273,);
not I_38628 (I660281,I642250);
DFFARX1 I_38629 (I642235,I3563,I660179,I660307,);
not I_38630 (I660315,I660307);
nor I_38631 (I660332,I660315,I660213);
and I_38632 (I660349,I660332,I642250);
nor I_38633 (I660366,I660315,I660281);
nor I_38634 (I660162,I660273,I660366);
DFFARX1 I_38635 (I642244,I3563,I660179,I660406,);
nor I_38636 (I660414,I660406,I660273);
not I_38637 (I660431,I660414);
not I_38638 (I660448,I660406);
nor I_38639 (I660465,I660448,I660349);
DFFARX1 I_38640 (I660465,I3563,I660179,I660165,);
nand I_38641 (I660496,I642241,I642232);
and I_38642 (I660513,I660496,I642229);
DFFARX1 I_38643 (I660513,I3563,I660179,I660539,);
nor I_38644 (I660547,I660539,I660406);
DFFARX1 I_38645 (I660547,I3563,I660179,I660147,);
nand I_38646 (I660578,I660539,I660448);
nand I_38647 (I660156,I660431,I660578);
not I_38648 (I660609,I660539);
nor I_38649 (I660626,I660609,I660349);
DFFARX1 I_38650 (I660626,I3563,I660179,I660168,);
nor I_38651 (I660657,I642232,I642232);
or I_38652 (I660159,I660406,I660657);
nor I_38653 (I660150,I660539,I660657);
or I_38654 (I660153,I660273,I660657);
DFFARX1 I_38655 (I660657,I3563,I660179,I660171,);
not I_38656 (I660757,I3570);
DFFARX1 I_38657 (I1098527,I3563,I660757,I660783,);
not I_38658 (I660791,I660783);
nand I_38659 (I660808,I1098509,I1098521);
and I_38660 (I660825,I660808,I1098524);
DFFARX1 I_38661 (I660825,I3563,I660757,I660851,);
not I_38662 (I660859,I1098518);
DFFARX1 I_38663 (I1098515,I3563,I660757,I660885,);
not I_38664 (I660893,I660885);
nor I_38665 (I660910,I660893,I660791);
and I_38666 (I660927,I660910,I1098518);
nor I_38667 (I660944,I660893,I660859);
nor I_38668 (I660740,I660851,I660944);
DFFARX1 I_38669 (I1098533,I3563,I660757,I660984,);
nor I_38670 (I660992,I660984,I660851);
not I_38671 (I661009,I660992);
not I_38672 (I661026,I660984);
nor I_38673 (I661043,I661026,I660927);
DFFARX1 I_38674 (I661043,I3563,I660757,I660743,);
nand I_38675 (I661074,I1098512,I1098512);
and I_38676 (I661091,I661074,I1098509);
DFFARX1 I_38677 (I661091,I3563,I660757,I661117,);
nor I_38678 (I661125,I661117,I660984);
DFFARX1 I_38679 (I661125,I3563,I660757,I660725,);
nand I_38680 (I661156,I661117,I661026);
nand I_38681 (I660734,I661009,I661156);
not I_38682 (I661187,I661117);
nor I_38683 (I661204,I661187,I660927);
DFFARX1 I_38684 (I661204,I3563,I660757,I660746,);
nor I_38685 (I661235,I1098530,I1098512);
or I_38686 (I660737,I660984,I661235);
nor I_38687 (I660728,I661117,I661235);
or I_38688 (I660731,I660851,I661235);
DFFARX1 I_38689 (I661235,I3563,I660757,I660749,);
not I_38690 (I661335,I3570);
DFFARX1 I_38691 (I1119335,I3563,I661335,I661361,);
not I_38692 (I661369,I661361);
nand I_38693 (I661386,I1119317,I1119329);
and I_38694 (I661403,I661386,I1119332);
DFFARX1 I_38695 (I661403,I3563,I661335,I661429,);
not I_38696 (I661437,I1119326);
DFFARX1 I_38697 (I1119323,I3563,I661335,I661463,);
not I_38698 (I661471,I661463);
nor I_38699 (I661488,I661471,I661369);
and I_38700 (I661505,I661488,I1119326);
nor I_38701 (I661522,I661471,I661437);
nor I_38702 (I661318,I661429,I661522);
DFFARX1 I_38703 (I1119341,I3563,I661335,I661562,);
nor I_38704 (I661570,I661562,I661429);
not I_38705 (I661587,I661570);
not I_38706 (I661604,I661562);
nor I_38707 (I661621,I661604,I661505);
DFFARX1 I_38708 (I661621,I3563,I661335,I661321,);
nand I_38709 (I661652,I1119320,I1119320);
and I_38710 (I661669,I661652,I1119317);
DFFARX1 I_38711 (I661669,I3563,I661335,I661695,);
nor I_38712 (I661703,I661695,I661562);
DFFARX1 I_38713 (I661703,I3563,I661335,I661303,);
nand I_38714 (I661734,I661695,I661604);
nand I_38715 (I661312,I661587,I661734);
not I_38716 (I661765,I661695);
nor I_38717 (I661782,I661765,I661505);
DFFARX1 I_38718 (I661782,I3563,I661335,I661324,);
nor I_38719 (I661813,I1119338,I1119320);
or I_38720 (I661315,I661562,I661813);
nor I_38721 (I661306,I661695,I661813);
or I_38722 (I661309,I661429,I661813);
DFFARX1 I_38723 (I661813,I3563,I661335,I661327,);
not I_38724 (I661913,I3570);
DFFARX1 I_38725 (I1090435,I3563,I661913,I661939,);
not I_38726 (I661947,I661939);
nand I_38727 (I661964,I1090417,I1090429);
and I_38728 (I661981,I661964,I1090432);
DFFARX1 I_38729 (I661981,I3563,I661913,I662007,);
not I_38730 (I662015,I1090426);
DFFARX1 I_38731 (I1090423,I3563,I661913,I662041,);
not I_38732 (I662049,I662041);
nor I_38733 (I662066,I662049,I661947);
and I_38734 (I662083,I662066,I1090426);
nor I_38735 (I662100,I662049,I662015);
nor I_38736 (I661896,I662007,I662100);
DFFARX1 I_38737 (I1090441,I3563,I661913,I662140,);
nor I_38738 (I662148,I662140,I662007);
not I_38739 (I662165,I662148);
not I_38740 (I662182,I662140);
nor I_38741 (I662199,I662182,I662083);
DFFARX1 I_38742 (I662199,I3563,I661913,I661899,);
nand I_38743 (I662230,I1090420,I1090420);
and I_38744 (I662247,I662230,I1090417);
DFFARX1 I_38745 (I662247,I3563,I661913,I662273,);
nor I_38746 (I662281,I662273,I662140);
DFFARX1 I_38747 (I662281,I3563,I661913,I661881,);
nand I_38748 (I662312,I662273,I662182);
nand I_38749 (I661890,I662165,I662312);
not I_38750 (I662343,I662273);
nor I_38751 (I662360,I662343,I662083);
DFFARX1 I_38752 (I662360,I3563,I661913,I661902,);
nor I_38753 (I662391,I1090438,I1090420);
or I_38754 (I661893,I662140,I662391);
nor I_38755 (I661884,I662273,I662391);
or I_38756 (I661887,I662007,I662391);
DFFARX1 I_38757 (I662391,I3563,I661913,I661905,);
not I_38758 (I662491,I3570);
DFFARX1 I_38759 (I1081447,I3563,I662491,I662517,);
not I_38760 (I662525,I662517);
nand I_38761 (I662542,I1081444,I1081462);
and I_38762 (I662559,I662542,I1081459);
DFFARX1 I_38763 (I662559,I3563,I662491,I662585,);
not I_38764 (I662593,I1081441);
DFFARX1 I_38765 (I1081444,I3563,I662491,I662619,);
not I_38766 (I662627,I662619);
nor I_38767 (I662644,I662627,I662525);
and I_38768 (I662661,I662644,I1081441);
nor I_38769 (I662678,I662627,I662593);
nor I_38770 (I662474,I662585,I662678);
DFFARX1 I_38771 (I1081453,I3563,I662491,I662718,);
nor I_38772 (I662726,I662718,I662585);
not I_38773 (I662743,I662726);
not I_38774 (I662760,I662718);
nor I_38775 (I662777,I662760,I662661);
DFFARX1 I_38776 (I662777,I3563,I662491,I662477,);
nand I_38777 (I662808,I1081456,I1081441);
and I_38778 (I662825,I662808,I1081447);
DFFARX1 I_38779 (I662825,I3563,I662491,I662851,);
nor I_38780 (I662859,I662851,I662718);
DFFARX1 I_38781 (I662859,I3563,I662491,I662459,);
nand I_38782 (I662890,I662851,I662760);
nand I_38783 (I662468,I662743,I662890);
not I_38784 (I662921,I662851);
nor I_38785 (I662938,I662921,I662661);
DFFARX1 I_38786 (I662938,I3563,I662491,I662480,);
nor I_38787 (I662969,I1081450,I1081441);
or I_38788 (I662471,I662718,I662969);
nor I_38789 (I662462,I662851,I662969);
or I_38790 (I662465,I662585,I662969);
DFFARX1 I_38791 (I662969,I3563,I662491,I662483,);
not I_38792 (I663069,I3570);
DFFARX1 I_38793 (I1074715,I3563,I663069,I663095,);
not I_38794 (I663103,I663095);
nand I_38795 (I663120,I1074712,I1074730);
and I_38796 (I663137,I663120,I1074727);
DFFARX1 I_38797 (I663137,I3563,I663069,I663163,);
not I_38798 (I663171,I1074709);
DFFARX1 I_38799 (I1074712,I3563,I663069,I663197,);
not I_38800 (I663205,I663197);
nor I_38801 (I663222,I663205,I663103);
and I_38802 (I663239,I663222,I1074709);
nor I_38803 (I663256,I663205,I663171);
nor I_38804 (I663052,I663163,I663256);
DFFARX1 I_38805 (I1074721,I3563,I663069,I663296,);
nor I_38806 (I663304,I663296,I663163);
not I_38807 (I663321,I663304);
not I_38808 (I663338,I663296);
nor I_38809 (I663355,I663338,I663239);
DFFARX1 I_38810 (I663355,I3563,I663069,I663055,);
nand I_38811 (I663386,I1074724,I1074709);
and I_38812 (I663403,I663386,I1074715);
DFFARX1 I_38813 (I663403,I3563,I663069,I663429,);
nor I_38814 (I663437,I663429,I663296);
DFFARX1 I_38815 (I663437,I3563,I663069,I663037,);
nand I_38816 (I663468,I663429,I663338);
nand I_38817 (I663046,I663321,I663468);
not I_38818 (I663499,I663429);
nor I_38819 (I663516,I663499,I663239);
DFFARX1 I_38820 (I663516,I3563,I663069,I663058,);
nor I_38821 (I663547,I1074718,I1074709);
or I_38822 (I663049,I663296,I663547);
nor I_38823 (I663040,I663429,I663547);
or I_38824 (I663043,I663163,I663547);
DFFARX1 I_38825 (I663547,I3563,I663069,I663061,);
not I_38826 (I663647,I3570);
DFFARX1 I_38827 (I859555,I3563,I663647,I663673,);
not I_38828 (I663681,I663673);
nand I_38829 (I663698,I859543,I859561);
and I_38830 (I663715,I663698,I859558);
DFFARX1 I_38831 (I663715,I3563,I663647,I663741,);
not I_38832 (I663749,I859549);
DFFARX1 I_38833 (I859546,I3563,I663647,I663775,);
not I_38834 (I663783,I663775);
nor I_38835 (I663800,I663783,I663681);
and I_38836 (I663817,I663800,I859549);
nor I_38837 (I663834,I663783,I663749);
nor I_38838 (I663630,I663741,I663834);
DFFARX1 I_38839 (I859540,I3563,I663647,I663874,);
nor I_38840 (I663882,I663874,I663741);
not I_38841 (I663899,I663882);
not I_38842 (I663916,I663874);
nor I_38843 (I663933,I663916,I663817);
DFFARX1 I_38844 (I663933,I3563,I663647,I663633,);
nand I_38845 (I663964,I859540,I859543);
and I_38846 (I663981,I663964,I859546);
DFFARX1 I_38847 (I663981,I3563,I663647,I664007,);
nor I_38848 (I664015,I664007,I663874);
DFFARX1 I_38849 (I664015,I3563,I663647,I663615,);
nand I_38850 (I664046,I664007,I663916);
nand I_38851 (I663624,I663899,I664046);
not I_38852 (I664077,I664007);
nor I_38853 (I664094,I664077,I663817);
DFFARX1 I_38854 (I664094,I3563,I663647,I663636,);
nor I_38855 (I664125,I859552,I859543);
or I_38856 (I663627,I663874,I664125);
nor I_38857 (I663618,I664007,I664125);
or I_38858 (I663621,I663741,I664125);
DFFARX1 I_38859 (I664125,I3563,I663647,I663639,);
not I_38860 (I664225,I3570);
DFFARX1 I_38861 (I1042161,I3563,I664225,I664251,);
not I_38862 (I664259,I664251);
nand I_38863 (I664276,I1042137,I1042152);
and I_38864 (I664293,I664276,I1042164);
DFFARX1 I_38865 (I664293,I3563,I664225,I664319,);
not I_38866 (I664327,I1042149);
DFFARX1 I_38867 (I1042140,I3563,I664225,I664353,);
not I_38868 (I664361,I664353);
nor I_38869 (I664378,I664361,I664259);
and I_38870 (I664395,I664378,I1042149);
nor I_38871 (I664412,I664361,I664327);
nor I_38872 (I664208,I664319,I664412);
DFFARX1 I_38873 (I1042137,I3563,I664225,I664452,);
nor I_38874 (I664460,I664452,I664319);
not I_38875 (I664477,I664460);
not I_38876 (I664494,I664452);
nor I_38877 (I664511,I664494,I664395);
DFFARX1 I_38878 (I664511,I3563,I664225,I664211,);
nand I_38879 (I664542,I1042155,I1042146);
and I_38880 (I664559,I664542,I1042158);
DFFARX1 I_38881 (I664559,I3563,I664225,I664585,);
nor I_38882 (I664593,I664585,I664452);
DFFARX1 I_38883 (I664593,I3563,I664225,I664193,);
nand I_38884 (I664624,I664585,I664494);
nand I_38885 (I664202,I664477,I664624);
not I_38886 (I664655,I664585);
nor I_38887 (I664672,I664655,I664395);
DFFARX1 I_38888 (I664672,I3563,I664225,I664214,);
nor I_38889 (I664703,I1042143,I1042146);
or I_38890 (I664205,I664452,I664703);
nor I_38891 (I664196,I664585,I664703);
or I_38892 (I664199,I664319,I664703);
DFFARX1 I_38893 (I664703,I3563,I664225,I664217,);
not I_38894 (I664803,I3570);
DFFARX1 I_38895 (I908039,I3563,I664803,I664829,);
not I_38896 (I664837,I664829);
nand I_38897 (I664854,I908027,I908045);
and I_38898 (I664871,I664854,I908042);
DFFARX1 I_38899 (I664871,I3563,I664803,I664897,);
not I_38900 (I664905,I908033);
DFFARX1 I_38901 (I908030,I3563,I664803,I664931,);
not I_38902 (I664939,I664931);
nor I_38903 (I664956,I664939,I664837);
and I_38904 (I664973,I664956,I908033);
nor I_38905 (I664990,I664939,I664905);
nor I_38906 (I664786,I664897,I664990);
DFFARX1 I_38907 (I908024,I3563,I664803,I665030,);
nor I_38908 (I665038,I665030,I664897);
not I_38909 (I665055,I665038);
not I_38910 (I665072,I665030);
nor I_38911 (I665089,I665072,I664973);
DFFARX1 I_38912 (I665089,I3563,I664803,I664789,);
nand I_38913 (I665120,I908024,I908027);
and I_38914 (I665137,I665120,I908030);
DFFARX1 I_38915 (I665137,I3563,I664803,I665163,);
nor I_38916 (I665171,I665163,I665030);
DFFARX1 I_38917 (I665171,I3563,I664803,I664771,);
nand I_38918 (I665202,I665163,I665072);
nand I_38919 (I664780,I665055,I665202);
not I_38920 (I665233,I665163);
nor I_38921 (I665250,I665233,I664973);
DFFARX1 I_38922 (I665250,I3563,I664803,I664792,);
nor I_38923 (I665281,I908036,I908027);
or I_38924 (I664783,I665030,I665281);
nor I_38925 (I664774,I665163,I665281);
or I_38926 (I664777,I664897,I665281);
DFFARX1 I_38927 (I665281,I3563,I664803,I664795,);
not I_38928 (I665381,I3570);
DFFARX1 I_38929 (I515435,I3563,I665381,I665407,);
not I_38930 (I665415,I665407);
nand I_38931 (I665432,I515426,I515444);
and I_38932 (I665449,I665432,I515447);
DFFARX1 I_38933 (I665449,I3563,I665381,I665475,);
not I_38934 (I665483,I515441);
DFFARX1 I_38935 (I515429,I3563,I665381,I665509,);
not I_38936 (I665517,I665509);
nor I_38937 (I665534,I665517,I665415);
and I_38938 (I665551,I665534,I515441);
nor I_38939 (I665568,I665517,I665483);
nor I_38940 (I665364,I665475,I665568);
DFFARX1 I_38941 (I515438,I3563,I665381,I665608,);
nor I_38942 (I665616,I665608,I665475);
not I_38943 (I665633,I665616);
not I_38944 (I665650,I665608);
nor I_38945 (I665667,I665650,I665551);
DFFARX1 I_38946 (I665667,I3563,I665381,I665367,);
nand I_38947 (I665698,I515453,I515450);
and I_38948 (I665715,I665698,I515432);
DFFARX1 I_38949 (I665715,I3563,I665381,I665741,);
nor I_38950 (I665749,I665741,I665608);
DFFARX1 I_38951 (I665749,I3563,I665381,I665349,);
nand I_38952 (I665780,I665741,I665650);
nand I_38953 (I665358,I665633,I665780);
not I_38954 (I665811,I665741);
nor I_38955 (I665828,I665811,I665551);
DFFARX1 I_38956 (I665828,I3563,I665381,I665370,);
nor I_38957 (I665859,I515426,I515450);
or I_38958 (I665361,I665608,I665859);
nor I_38959 (I665352,I665741,I665859);
or I_38960 (I665355,I665475,I665859);
DFFARX1 I_38961 (I665859,I3563,I665381,I665373,);
not I_38962 (I665959,I3570);
DFFARX1 I_38963 (I1157483,I3563,I665959,I665985,);
not I_38964 (I665993,I665985);
nand I_38965 (I666010,I1157465,I1157477);
and I_38966 (I666027,I666010,I1157480);
DFFARX1 I_38967 (I666027,I3563,I665959,I666053,);
not I_38968 (I666061,I1157474);
DFFARX1 I_38969 (I1157471,I3563,I665959,I666087,);
not I_38970 (I666095,I666087);
nor I_38971 (I666112,I666095,I665993);
and I_38972 (I666129,I666112,I1157474);
nor I_38973 (I666146,I666095,I666061);
nor I_38974 (I665942,I666053,I666146);
DFFARX1 I_38975 (I1157489,I3563,I665959,I666186,);
nor I_38976 (I666194,I666186,I666053);
not I_38977 (I666211,I666194);
not I_38978 (I666228,I666186);
nor I_38979 (I666245,I666228,I666129);
DFFARX1 I_38980 (I666245,I3563,I665959,I665945,);
nand I_38981 (I666276,I1157468,I1157468);
and I_38982 (I666293,I666276,I1157465);
DFFARX1 I_38983 (I666293,I3563,I665959,I666319,);
nor I_38984 (I666327,I666319,I666186);
DFFARX1 I_38985 (I666327,I3563,I665959,I665927,);
nand I_38986 (I666358,I666319,I666228);
nand I_38987 (I665936,I666211,I666358);
not I_38988 (I666389,I666319);
nor I_38989 (I666406,I666389,I666129);
DFFARX1 I_38990 (I666406,I3563,I665959,I665948,);
nor I_38991 (I666437,I1157486,I1157468);
or I_38992 (I665939,I666186,I666437);
nor I_38993 (I665930,I666319,I666437);
or I_38994 (I665933,I666053,I666437);
DFFARX1 I_38995 (I666437,I3563,I665959,I665951,);
not I_38996 (I666537,I3570);
DFFARX1 I_38997 (I10719,I3563,I666537,I666563,);
not I_38998 (I666571,I666563);
nand I_38999 (I666588,I10722,I10734);
and I_39000 (I666605,I666588,I10713);
DFFARX1 I_39001 (I666605,I3563,I666537,I666631,);
not I_39002 (I666639,I10713);
DFFARX1 I_39003 (I10716,I3563,I666537,I666665,);
not I_39004 (I666673,I666665);
nor I_39005 (I666690,I666673,I666571);
and I_39006 (I666707,I666690,I10713);
nor I_39007 (I666724,I666673,I666639);
nor I_39008 (I666520,I666631,I666724);
DFFARX1 I_39009 (I10728,I3563,I666537,I666764,);
nor I_39010 (I666772,I666764,I666631);
not I_39011 (I666789,I666772);
not I_39012 (I666806,I666764);
nor I_39013 (I666823,I666806,I666707);
DFFARX1 I_39014 (I666823,I3563,I666537,I666523,);
nand I_39015 (I666854,I10731,I10716);
and I_39016 (I666871,I666854,I10725);
DFFARX1 I_39017 (I666871,I3563,I666537,I666897,);
nor I_39018 (I666905,I666897,I666764);
DFFARX1 I_39019 (I666905,I3563,I666537,I666505,);
nand I_39020 (I666936,I666897,I666806);
nand I_39021 (I666514,I666789,I666936);
not I_39022 (I666967,I666897);
nor I_39023 (I666984,I666967,I666707);
DFFARX1 I_39024 (I666984,I3563,I666537,I666526,);
nor I_39025 (I667015,I10719,I10716);
or I_39026 (I666517,I666764,I667015);
nor I_39027 (I666508,I666897,I667015);
or I_39028 (I666511,I666631,I667015);
DFFARX1 I_39029 (I667015,I3563,I666537,I666529,);
not I_39030 (I667115,I3570);
DFFARX1 I_39031 (I1166731,I3563,I667115,I667141,);
not I_39032 (I667149,I667141);
nand I_39033 (I667166,I1166713,I1166725);
and I_39034 (I667183,I667166,I1166728);
DFFARX1 I_39035 (I667183,I3563,I667115,I667209,);
not I_39036 (I667217,I1166722);
DFFARX1 I_39037 (I1166719,I3563,I667115,I667243,);
not I_39038 (I667251,I667243);
nor I_39039 (I667268,I667251,I667149);
and I_39040 (I667285,I667268,I1166722);
nor I_39041 (I667302,I667251,I667217);
nor I_39042 (I667098,I667209,I667302);
DFFARX1 I_39043 (I1166737,I3563,I667115,I667342,);
nor I_39044 (I667350,I667342,I667209);
not I_39045 (I667367,I667350);
not I_39046 (I667384,I667342);
nor I_39047 (I667401,I667384,I667285);
DFFARX1 I_39048 (I667401,I3563,I667115,I667101,);
nand I_39049 (I667432,I1166716,I1166716);
and I_39050 (I667449,I667432,I1166713);
DFFARX1 I_39051 (I667449,I3563,I667115,I667475,);
nor I_39052 (I667483,I667475,I667342);
DFFARX1 I_39053 (I667483,I3563,I667115,I667083,);
nand I_39054 (I667514,I667475,I667384);
nand I_39055 (I667092,I667367,I667514);
not I_39056 (I667545,I667475);
nor I_39057 (I667562,I667545,I667285);
DFFARX1 I_39058 (I667562,I3563,I667115,I667104,);
nor I_39059 (I667593,I1166734,I1166716);
or I_39060 (I667095,I667342,I667593);
nor I_39061 (I667086,I667475,I667593);
or I_39062 (I667089,I667209,I667593);
DFFARX1 I_39063 (I667593,I3563,I667115,I667107,);
not I_39064 (I667693,I3570);
DFFARX1 I_39065 (I373925,I3563,I667693,I667719,);
not I_39066 (I667727,I667719);
nand I_39067 (I667744,I373928,I373904);
and I_39068 (I667761,I667744,I373901);
DFFARX1 I_39069 (I667761,I3563,I667693,I667787,);
not I_39070 (I667795,I373907);
DFFARX1 I_39071 (I373901,I3563,I667693,I667821,);
not I_39072 (I667829,I667821);
nor I_39073 (I667846,I667829,I667727);
and I_39074 (I667863,I667846,I373907);
nor I_39075 (I667880,I667829,I667795);
nor I_39076 (I667676,I667787,I667880);
DFFARX1 I_39077 (I373910,I3563,I667693,I667920,);
nor I_39078 (I667928,I667920,I667787);
not I_39079 (I667945,I667928);
not I_39080 (I667962,I667920);
nor I_39081 (I667979,I667962,I667863);
DFFARX1 I_39082 (I667979,I3563,I667693,I667679,);
nand I_39083 (I668010,I373913,I373922);
and I_39084 (I668027,I668010,I373919);
DFFARX1 I_39085 (I668027,I3563,I667693,I668053,);
nor I_39086 (I668061,I668053,I667920);
DFFARX1 I_39087 (I668061,I3563,I667693,I667661,);
nand I_39088 (I668092,I668053,I667962);
nand I_39089 (I667670,I667945,I668092);
not I_39090 (I668123,I668053);
nor I_39091 (I668140,I668123,I667863);
DFFARX1 I_39092 (I668140,I3563,I667693,I667682,);
nor I_39093 (I668171,I373916,I373922);
or I_39094 (I667673,I667920,I668171);
nor I_39095 (I667664,I668053,I668171);
or I_39096 (I667667,I667787,I668171);
DFFARX1 I_39097 (I668171,I3563,I667693,I667685,);
not I_39098 (I668271,I3570);
DFFARX1 I_39099 (I1223953,I3563,I668271,I668297,);
not I_39100 (I668305,I668297);
nand I_39101 (I668322,I1223935,I1223947);
and I_39102 (I668339,I668322,I1223950);
DFFARX1 I_39103 (I668339,I3563,I668271,I668365,);
not I_39104 (I668373,I1223944);
DFFARX1 I_39105 (I1223941,I3563,I668271,I668399,);
not I_39106 (I668407,I668399);
nor I_39107 (I668424,I668407,I668305);
and I_39108 (I668441,I668424,I1223944);
nor I_39109 (I668458,I668407,I668373);
nor I_39110 (I668254,I668365,I668458);
DFFARX1 I_39111 (I1223959,I3563,I668271,I668498,);
nor I_39112 (I668506,I668498,I668365);
not I_39113 (I668523,I668506);
not I_39114 (I668540,I668498);
nor I_39115 (I668557,I668540,I668441);
DFFARX1 I_39116 (I668557,I3563,I668271,I668257,);
nand I_39117 (I668588,I1223938,I1223938);
and I_39118 (I668605,I668588,I1223935);
DFFARX1 I_39119 (I668605,I3563,I668271,I668631,);
nor I_39120 (I668639,I668631,I668498);
DFFARX1 I_39121 (I668639,I3563,I668271,I668239,);
nand I_39122 (I668670,I668631,I668540);
nand I_39123 (I668248,I668523,I668670);
not I_39124 (I668701,I668631);
nor I_39125 (I668718,I668701,I668441);
DFFARX1 I_39126 (I668718,I3563,I668271,I668260,);
nor I_39127 (I668749,I1223956,I1223938);
or I_39128 (I668251,I668498,I668749);
nor I_39129 (I668242,I668631,I668749);
or I_39130 (I668245,I668365,I668749);
DFFARX1 I_39131 (I668749,I3563,I668271,I668263,);
not I_39132 (I668849,I3570);
DFFARX1 I_39133 (I1178291,I3563,I668849,I668875,);
not I_39134 (I668883,I668875);
nand I_39135 (I668900,I1178273,I1178285);
and I_39136 (I668917,I668900,I1178288);
DFFARX1 I_39137 (I668917,I3563,I668849,I668943,);
not I_39138 (I668951,I1178282);
DFFARX1 I_39139 (I1178279,I3563,I668849,I668977,);
not I_39140 (I668985,I668977);
nor I_39141 (I669002,I668985,I668883);
and I_39142 (I669019,I669002,I1178282);
nor I_39143 (I669036,I668985,I668951);
nor I_39144 (I668832,I668943,I669036);
DFFARX1 I_39145 (I1178297,I3563,I668849,I669076,);
nor I_39146 (I669084,I669076,I668943);
not I_39147 (I669101,I669084);
not I_39148 (I669118,I669076);
nor I_39149 (I669135,I669118,I669019);
DFFARX1 I_39150 (I669135,I3563,I668849,I668835,);
nand I_39151 (I669166,I1178276,I1178276);
and I_39152 (I669183,I669166,I1178273);
DFFARX1 I_39153 (I669183,I3563,I668849,I669209,);
nor I_39154 (I669217,I669209,I669076);
DFFARX1 I_39155 (I669217,I3563,I668849,I668817,);
nand I_39156 (I669248,I669209,I669118);
nand I_39157 (I668826,I669101,I669248);
not I_39158 (I669279,I669209);
nor I_39159 (I669296,I669279,I669019);
DFFARX1 I_39160 (I669296,I3563,I668849,I668838,);
nor I_39161 (I669327,I1178294,I1178276);
or I_39162 (I668829,I669076,I669327);
nor I_39163 (I668820,I669209,I669327);
or I_39164 (I668823,I668943,I669327);
DFFARX1 I_39165 (I669327,I3563,I668849,I668841,);
not I_39166 (I669427,I3570);
DFFARX1 I_39167 (I1029887,I3563,I669427,I669453,);
not I_39168 (I669461,I669453);
nand I_39169 (I669478,I1029863,I1029878);
and I_39170 (I669495,I669478,I1029890);
DFFARX1 I_39171 (I669495,I3563,I669427,I669521,);
not I_39172 (I669529,I1029875);
DFFARX1 I_39173 (I1029866,I3563,I669427,I669555,);
not I_39174 (I669563,I669555);
nor I_39175 (I669580,I669563,I669461);
and I_39176 (I669597,I669580,I1029875);
nor I_39177 (I669614,I669563,I669529);
nor I_39178 (I669410,I669521,I669614);
DFFARX1 I_39179 (I1029863,I3563,I669427,I669654,);
nor I_39180 (I669662,I669654,I669521);
not I_39181 (I669679,I669662);
not I_39182 (I669696,I669654);
nor I_39183 (I669713,I669696,I669597);
DFFARX1 I_39184 (I669713,I3563,I669427,I669413,);
nand I_39185 (I669744,I1029881,I1029872);
and I_39186 (I669761,I669744,I1029884);
DFFARX1 I_39187 (I669761,I3563,I669427,I669787,);
nor I_39188 (I669795,I669787,I669654);
DFFARX1 I_39189 (I669795,I3563,I669427,I669395,);
nand I_39190 (I669826,I669787,I669696);
nand I_39191 (I669404,I669679,I669826);
not I_39192 (I669857,I669787);
nor I_39193 (I669874,I669857,I669597);
DFFARX1 I_39194 (I669874,I3563,I669427,I669416,);
nor I_39195 (I669905,I1029869,I1029872);
or I_39196 (I669407,I669654,I669905);
nor I_39197 (I669398,I669787,I669905);
or I_39198 (I669401,I669521,I669905);
DFFARX1 I_39199 (I669905,I3563,I669427,I669419,);
not I_39200 (I670005,I3570);
DFFARX1 I_39201 (I656101,I3563,I670005,I670031,);
not I_39202 (I670039,I670031);
nand I_39203 (I670056,I656110,I656119);
and I_39204 (I670073,I670056,I656125);
DFFARX1 I_39205 (I670073,I3563,I670005,I670099,);
not I_39206 (I670107,I656122);
DFFARX1 I_39207 (I656107,I3563,I670005,I670133,);
not I_39208 (I670141,I670133);
nor I_39209 (I670158,I670141,I670039);
and I_39210 (I670175,I670158,I656122);
nor I_39211 (I670192,I670141,I670107);
nor I_39212 (I669988,I670099,I670192);
DFFARX1 I_39213 (I656116,I3563,I670005,I670232,);
nor I_39214 (I670240,I670232,I670099);
not I_39215 (I670257,I670240);
not I_39216 (I670274,I670232);
nor I_39217 (I670291,I670274,I670175);
DFFARX1 I_39218 (I670291,I3563,I670005,I669991,);
nand I_39219 (I670322,I656113,I656104);
and I_39220 (I670339,I670322,I656101);
DFFARX1 I_39221 (I670339,I3563,I670005,I670365,);
nor I_39222 (I670373,I670365,I670232);
DFFARX1 I_39223 (I670373,I3563,I670005,I669973,);
nand I_39224 (I670404,I670365,I670274);
nand I_39225 (I669982,I670257,I670404);
not I_39226 (I670435,I670365);
nor I_39227 (I670452,I670435,I670175);
DFFARX1 I_39228 (I670452,I3563,I670005,I669994,);
nor I_39229 (I670483,I656104,I656104);
or I_39230 (I669985,I670232,I670483);
nor I_39231 (I669976,I670365,I670483);
or I_39232 (I669979,I670099,I670483);
DFFARX1 I_39233 (I670483,I3563,I670005,I669997,);
not I_39234 (I670583,I3570);
DFFARX1 I_39235 (I1252937,I3563,I670583,I670609,);
not I_39236 (I670617,I670609);
nand I_39237 (I670634,I1252940,I1252949);
and I_39238 (I670651,I670634,I1252952);
DFFARX1 I_39239 (I670651,I3563,I670583,I670677,);
not I_39240 (I670685,I1252961);
DFFARX1 I_39241 (I1252943,I3563,I670583,I670711,);
not I_39242 (I670719,I670711);
nor I_39243 (I670736,I670719,I670617);
and I_39244 (I670753,I670736,I1252961);
nor I_39245 (I670770,I670719,I670685);
nor I_39246 (I670566,I670677,I670770);
DFFARX1 I_39247 (I1252940,I3563,I670583,I670810,);
nor I_39248 (I670818,I670810,I670677);
not I_39249 (I670835,I670818);
not I_39250 (I670852,I670810);
nor I_39251 (I670869,I670852,I670753);
DFFARX1 I_39252 (I670869,I3563,I670583,I670569,);
nand I_39253 (I670900,I1252958,I1252937);
and I_39254 (I670917,I670900,I1252955);
DFFARX1 I_39255 (I670917,I3563,I670583,I670943,);
nor I_39256 (I670951,I670943,I670810);
DFFARX1 I_39257 (I670951,I3563,I670583,I670551,);
nand I_39258 (I670982,I670943,I670852);
nand I_39259 (I670560,I670835,I670982);
not I_39260 (I671013,I670943);
nor I_39261 (I671030,I671013,I670753);
DFFARX1 I_39262 (I671030,I3563,I670583,I670572,);
nor I_39263 (I671061,I1252946,I1252937);
or I_39264 (I670563,I670810,I671061);
nor I_39265 (I670554,I670943,I671061);
or I_39266 (I670557,I670677,I671061);
DFFARX1 I_39267 (I671061,I3563,I670583,I670575,);
not I_39268 (I671161,I3570);
DFFARX1 I_39269 (I1169043,I3563,I671161,I671187,);
not I_39270 (I671195,I671187);
nand I_39271 (I671212,I1169025,I1169037);
and I_39272 (I671229,I671212,I1169040);
DFFARX1 I_39273 (I671229,I3563,I671161,I671255,);
not I_39274 (I671263,I1169034);
DFFARX1 I_39275 (I1169031,I3563,I671161,I671289,);
not I_39276 (I671297,I671289);
nor I_39277 (I671314,I671297,I671195);
and I_39278 (I671331,I671314,I1169034);
nor I_39279 (I671348,I671297,I671263);
nor I_39280 (I671144,I671255,I671348);
DFFARX1 I_39281 (I1169049,I3563,I671161,I671388,);
nor I_39282 (I671396,I671388,I671255);
not I_39283 (I671413,I671396);
not I_39284 (I671430,I671388);
nor I_39285 (I671447,I671430,I671331);
DFFARX1 I_39286 (I671447,I3563,I671161,I671147,);
nand I_39287 (I671478,I1169028,I1169028);
and I_39288 (I671495,I671478,I1169025);
DFFARX1 I_39289 (I671495,I3563,I671161,I671521,);
nor I_39290 (I671529,I671521,I671388);
DFFARX1 I_39291 (I671529,I3563,I671161,I671129,);
nand I_39292 (I671560,I671521,I671430);
nand I_39293 (I671138,I671413,I671560);
not I_39294 (I671591,I671521);
nor I_39295 (I671608,I671591,I671331);
DFFARX1 I_39296 (I671608,I3563,I671161,I671150,);
nor I_39297 (I671639,I1169046,I1169028);
or I_39298 (I671141,I671388,I671639);
nor I_39299 (I671132,I671521,I671639);
or I_39300 (I671135,I671255,I671639);
DFFARX1 I_39301 (I671639,I3563,I671161,I671153,);
not I_39302 (I671739,I3570);
DFFARX1 I_39303 (I1364875,I3563,I671739,I671765,);
not I_39304 (I671773,I671765);
nand I_39305 (I671790,I1364860,I1364848);
and I_39306 (I671807,I671790,I1364863);
DFFARX1 I_39307 (I671807,I3563,I671739,I671833,);
not I_39308 (I671841,I1364848);
DFFARX1 I_39309 (I1364866,I3563,I671739,I671867,);
not I_39310 (I671875,I671867);
nor I_39311 (I671892,I671875,I671773);
and I_39312 (I671909,I671892,I1364848);
nor I_39313 (I671926,I671875,I671841);
nor I_39314 (I671722,I671833,I671926);
DFFARX1 I_39315 (I1364854,I3563,I671739,I671966,);
nor I_39316 (I671974,I671966,I671833);
not I_39317 (I671991,I671974);
not I_39318 (I672008,I671966);
nor I_39319 (I672025,I672008,I671909);
DFFARX1 I_39320 (I672025,I3563,I671739,I671725,);
nand I_39321 (I672056,I1364851,I1364857);
and I_39322 (I672073,I672056,I1364872);
DFFARX1 I_39323 (I672073,I3563,I671739,I672099,);
nor I_39324 (I672107,I672099,I671966);
DFFARX1 I_39325 (I672107,I3563,I671739,I671707,);
nand I_39326 (I672138,I672099,I672008);
nand I_39327 (I671716,I671991,I672138);
not I_39328 (I672169,I672099);
nor I_39329 (I672186,I672169,I671909);
DFFARX1 I_39330 (I672186,I3563,I671739,I671728,);
nor I_39331 (I672217,I1364869,I1364857);
or I_39332 (I671719,I671966,I672217);
nor I_39333 (I671710,I672099,I672217);
or I_39334 (I671713,I671833,I672217);
DFFARX1 I_39335 (I672217,I3563,I671739,I671731,);
not I_39336 (I672317,I3570);
DFFARX1 I_39337 (I401329,I3563,I672317,I672343,);
not I_39338 (I672351,I672343);
nand I_39339 (I672368,I401332,I401308);
and I_39340 (I672385,I672368,I401305);
DFFARX1 I_39341 (I672385,I3563,I672317,I672411,);
not I_39342 (I672419,I401311);
DFFARX1 I_39343 (I401305,I3563,I672317,I672445,);
not I_39344 (I672453,I672445);
nor I_39345 (I672470,I672453,I672351);
and I_39346 (I672487,I672470,I401311);
nor I_39347 (I672504,I672453,I672419);
nor I_39348 (I672300,I672411,I672504);
DFFARX1 I_39349 (I401314,I3563,I672317,I672544,);
nor I_39350 (I672552,I672544,I672411);
not I_39351 (I672569,I672552);
not I_39352 (I672586,I672544);
nor I_39353 (I672603,I672586,I672487);
DFFARX1 I_39354 (I672603,I3563,I672317,I672303,);
nand I_39355 (I672634,I401317,I401326);
and I_39356 (I672651,I672634,I401323);
DFFARX1 I_39357 (I672651,I3563,I672317,I672677,);
nor I_39358 (I672685,I672677,I672544);
DFFARX1 I_39359 (I672685,I3563,I672317,I672285,);
nand I_39360 (I672716,I672677,I672586);
nand I_39361 (I672294,I672569,I672716);
not I_39362 (I672747,I672677);
nor I_39363 (I672764,I672747,I672487);
DFFARX1 I_39364 (I672764,I3563,I672317,I672306,);
nor I_39365 (I672795,I401320,I401326);
or I_39366 (I672297,I672544,I672795);
nor I_39367 (I672288,I672677,I672795);
or I_39368 (I672291,I672411,I672795);
DFFARX1 I_39369 (I672795,I3563,I672317,I672309,);
not I_39370 (I672895,I3570);
DFFARX1 I_39371 (I930403,I3563,I672895,I672921,);
not I_39372 (I672929,I672921);
nand I_39373 (I672946,I930379,I930394);
and I_39374 (I672963,I672946,I930406);
DFFARX1 I_39375 (I672963,I3563,I672895,I672989,);
not I_39376 (I672997,I930391);
DFFARX1 I_39377 (I930382,I3563,I672895,I673023,);
not I_39378 (I673031,I673023);
nor I_39379 (I673048,I673031,I672929);
and I_39380 (I673065,I673048,I930391);
nor I_39381 (I673082,I673031,I672997);
nor I_39382 (I672878,I672989,I673082);
DFFARX1 I_39383 (I930379,I3563,I672895,I673122,);
nor I_39384 (I673130,I673122,I672989);
not I_39385 (I673147,I673130);
not I_39386 (I673164,I673122);
nor I_39387 (I673181,I673164,I673065);
DFFARX1 I_39388 (I673181,I3563,I672895,I672881,);
nand I_39389 (I673212,I930397,I930388);
and I_39390 (I673229,I673212,I930400);
DFFARX1 I_39391 (I673229,I3563,I672895,I673255,);
nor I_39392 (I673263,I673255,I673122);
DFFARX1 I_39393 (I673263,I3563,I672895,I672863,);
nand I_39394 (I673294,I673255,I673164);
nand I_39395 (I672872,I673147,I673294);
not I_39396 (I673325,I673255);
nor I_39397 (I673342,I673325,I673065);
DFFARX1 I_39398 (I673342,I3563,I672895,I672884,);
nor I_39399 (I673373,I930385,I930388);
or I_39400 (I672875,I673122,I673373);
nor I_39401 (I672866,I673255,I673373);
or I_39402 (I672869,I672989,I673373);
DFFARX1 I_39403 (I673373,I3563,I672895,I672887,);
not I_39404 (I673473,I3570);
DFFARX1 I_39405 (I1141877,I3563,I673473,I673499,);
not I_39406 (I673507,I673499);
nand I_39407 (I673524,I1141859,I1141871);
and I_39408 (I673541,I673524,I1141874);
DFFARX1 I_39409 (I673541,I3563,I673473,I673567,);
not I_39410 (I673575,I1141868);
DFFARX1 I_39411 (I1141865,I3563,I673473,I673601,);
not I_39412 (I673609,I673601);
nor I_39413 (I673626,I673609,I673507);
and I_39414 (I673643,I673626,I1141868);
nor I_39415 (I673660,I673609,I673575);
nor I_39416 (I673456,I673567,I673660);
DFFARX1 I_39417 (I1141883,I3563,I673473,I673700,);
nor I_39418 (I673708,I673700,I673567);
not I_39419 (I673725,I673708);
not I_39420 (I673742,I673700);
nor I_39421 (I673759,I673742,I673643);
DFFARX1 I_39422 (I673759,I3563,I673473,I673459,);
nand I_39423 (I673790,I1141862,I1141862);
and I_39424 (I673807,I673790,I1141859);
DFFARX1 I_39425 (I673807,I3563,I673473,I673833,);
nor I_39426 (I673841,I673833,I673700);
DFFARX1 I_39427 (I673841,I3563,I673473,I673441,);
nand I_39428 (I673872,I673833,I673742);
nand I_39429 (I673450,I673725,I673872);
not I_39430 (I673903,I673833);
nor I_39431 (I673920,I673903,I673643);
DFFARX1 I_39432 (I673920,I3563,I673473,I673462,);
nor I_39433 (I673951,I1141880,I1141862);
or I_39434 (I673453,I673700,I673951);
nor I_39435 (I673444,I673833,I673951);
or I_39436 (I673447,I673567,I673951);
DFFARX1 I_39437 (I673951,I3563,I673473,I673465,);
not I_39438 (I674051,I3570);
DFFARX1 I_39439 (I401856,I3563,I674051,I674077,);
not I_39440 (I674085,I674077);
nand I_39441 (I674102,I401859,I401835);
and I_39442 (I674119,I674102,I401832);
DFFARX1 I_39443 (I674119,I3563,I674051,I674145,);
not I_39444 (I674153,I401838);
DFFARX1 I_39445 (I401832,I3563,I674051,I674179,);
not I_39446 (I674187,I674179);
nor I_39447 (I674204,I674187,I674085);
and I_39448 (I674221,I674204,I401838);
nor I_39449 (I674238,I674187,I674153);
nor I_39450 (I674034,I674145,I674238);
DFFARX1 I_39451 (I401841,I3563,I674051,I674278,);
nor I_39452 (I674286,I674278,I674145);
not I_39453 (I674303,I674286);
not I_39454 (I674320,I674278);
nor I_39455 (I674337,I674320,I674221);
DFFARX1 I_39456 (I674337,I3563,I674051,I674037,);
nand I_39457 (I674368,I401844,I401853);
and I_39458 (I674385,I674368,I401850);
DFFARX1 I_39459 (I674385,I3563,I674051,I674411,);
nor I_39460 (I674419,I674411,I674278);
DFFARX1 I_39461 (I674419,I3563,I674051,I674019,);
nand I_39462 (I674450,I674411,I674320);
nand I_39463 (I674028,I674303,I674450);
not I_39464 (I674481,I674411);
nor I_39465 (I674498,I674481,I674221);
DFFARX1 I_39466 (I674498,I3563,I674051,I674040,);
nor I_39467 (I674529,I401847,I401853);
or I_39468 (I674031,I674278,I674529);
nor I_39469 (I674022,I674411,I674529);
or I_39470 (I674025,I674145,I674529);
DFFARX1 I_39471 (I674529,I3563,I674051,I674043,);
not I_39472 (I674629,I3570);
DFFARX1 I_39473 (I863771,I3563,I674629,I674655,);
not I_39474 (I674663,I674655);
nand I_39475 (I674680,I863759,I863777);
and I_39476 (I674697,I674680,I863774);
DFFARX1 I_39477 (I674697,I3563,I674629,I674723,);
not I_39478 (I674731,I863765);
DFFARX1 I_39479 (I863762,I3563,I674629,I674757,);
not I_39480 (I674765,I674757);
nor I_39481 (I674782,I674765,I674663);
and I_39482 (I674799,I674782,I863765);
nor I_39483 (I674816,I674765,I674731);
nor I_39484 (I674612,I674723,I674816);
DFFARX1 I_39485 (I863756,I3563,I674629,I674856,);
nor I_39486 (I674864,I674856,I674723);
not I_39487 (I674881,I674864);
not I_39488 (I674898,I674856);
nor I_39489 (I674915,I674898,I674799);
DFFARX1 I_39490 (I674915,I3563,I674629,I674615,);
nand I_39491 (I674946,I863756,I863759);
and I_39492 (I674963,I674946,I863762);
DFFARX1 I_39493 (I674963,I3563,I674629,I674989,);
nor I_39494 (I674997,I674989,I674856);
DFFARX1 I_39495 (I674997,I3563,I674629,I674597,);
nand I_39496 (I675028,I674989,I674898);
nand I_39497 (I674606,I674881,I675028);
not I_39498 (I675059,I674989);
nor I_39499 (I675076,I675059,I674799);
DFFARX1 I_39500 (I675076,I3563,I674629,I674618,);
nor I_39501 (I675107,I863768,I863759);
or I_39502 (I674609,I674856,I675107);
nor I_39503 (I674600,I674989,I675107);
or I_39504 (I674603,I674723,I675107);
DFFARX1 I_39505 (I675107,I3563,I674629,I674621,);
not I_39506 (I675207,I3570);
DFFARX1 I_39507 (I157307,I3563,I675207,I675233,);
not I_39508 (I675241,I675233);
nand I_39509 (I675258,I157316,I157325);
and I_39510 (I675275,I675258,I157304);
DFFARX1 I_39511 (I675275,I3563,I675207,I675301,);
not I_39512 (I675309,I157307);
DFFARX1 I_39513 (I157322,I3563,I675207,I675335,);
not I_39514 (I675343,I675335);
nor I_39515 (I675360,I675343,I675241);
and I_39516 (I675377,I675360,I157307);
nor I_39517 (I675394,I675343,I675309);
nor I_39518 (I675190,I675301,I675394);
DFFARX1 I_39519 (I157313,I3563,I675207,I675434,);
nor I_39520 (I675442,I675434,I675301);
not I_39521 (I675459,I675442);
not I_39522 (I675476,I675434);
nor I_39523 (I675493,I675476,I675377);
DFFARX1 I_39524 (I675493,I3563,I675207,I675193,);
nand I_39525 (I675524,I157328,I157304);
and I_39526 (I675541,I675524,I157310);
DFFARX1 I_39527 (I675541,I3563,I675207,I675567,);
nor I_39528 (I675575,I675567,I675434);
DFFARX1 I_39529 (I675575,I3563,I675207,I675175,);
nand I_39530 (I675606,I675567,I675476);
nand I_39531 (I675184,I675459,I675606);
not I_39532 (I675637,I675567);
nor I_39533 (I675654,I675637,I675377);
DFFARX1 I_39534 (I675654,I3563,I675207,I675196,);
nor I_39535 (I675685,I157319,I157304);
or I_39536 (I675187,I675434,I675685);
nor I_39537 (I675178,I675567,I675685);
or I_39538 (I675181,I675301,I675685);
DFFARX1 I_39539 (I675685,I3563,I675207,I675199,);
not I_39540 (I675785,I3570);
DFFARX1 I_39541 (I1291221,I3563,I675785,I675811,);
not I_39542 (I675819,I675811);
nand I_39543 (I675836,I1291245,I1291227);
and I_39544 (I675853,I675836,I1291233);
DFFARX1 I_39545 (I675853,I3563,I675785,I675879,);
not I_39546 (I675887,I1291239);
DFFARX1 I_39547 (I1291224,I3563,I675785,I675913,);
not I_39548 (I675921,I675913);
nor I_39549 (I675938,I675921,I675819);
and I_39550 (I675955,I675938,I1291239);
nor I_39551 (I675972,I675921,I675887);
nor I_39552 (I675768,I675879,I675972);
DFFARX1 I_39553 (I1291236,I3563,I675785,I676012,);
nor I_39554 (I676020,I676012,I675879);
not I_39555 (I676037,I676020);
not I_39556 (I676054,I676012);
nor I_39557 (I676071,I676054,I675955);
DFFARX1 I_39558 (I676071,I3563,I675785,I675771,);
nand I_39559 (I676102,I1291242,I1291230);
and I_39560 (I676119,I676102,I1291224);
DFFARX1 I_39561 (I676119,I3563,I675785,I676145,);
nor I_39562 (I676153,I676145,I676012);
DFFARX1 I_39563 (I676153,I3563,I675785,I675753,);
nand I_39564 (I676184,I676145,I676054);
nand I_39565 (I675762,I676037,I676184);
not I_39566 (I676215,I676145);
nor I_39567 (I676232,I676215,I675955);
DFFARX1 I_39568 (I676232,I3563,I675785,I675774,);
nor I_39569 (I676263,I1291221,I1291230);
or I_39570 (I675765,I676012,I676263);
nor I_39571 (I675756,I676145,I676263);
or I_39572 (I675759,I675879,I676263);
DFFARX1 I_39573 (I676263,I3563,I675785,I675777,);
not I_39574 (I676363,I3570);
DFFARX1 I_39575 (I821611,I3563,I676363,I676389,);
not I_39576 (I676397,I676389);
nand I_39577 (I676414,I821599,I821617);
and I_39578 (I676431,I676414,I821614);
DFFARX1 I_39579 (I676431,I3563,I676363,I676457,);
not I_39580 (I676465,I821605);
DFFARX1 I_39581 (I821602,I3563,I676363,I676491,);
not I_39582 (I676499,I676491);
nor I_39583 (I676516,I676499,I676397);
and I_39584 (I676533,I676516,I821605);
nor I_39585 (I676550,I676499,I676465);
nor I_39586 (I676346,I676457,I676550);
DFFARX1 I_39587 (I821596,I3563,I676363,I676590,);
nor I_39588 (I676598,I676590,I676457);
not I_39589 (I676615,I676598);
not I_39590 (I676632,I676590);
nor I_39591 (I676649,I676632,I676533);
DFFARX1 I_39592 (I676649,I3563,I676363,I676349,);
nand I_39593 (I676680,I821596,I821599);
and I_39594 (I676697,I676680,I821602);
DFFARX1 I_39595 (I676697,I3563,I676363,I676723,);
nor I_39596 (I676731,I676723,I676590);
DFFARX1 I_39597 (I676731,I3563,I676363,I676331,);
nand I_39598 (I676762,I676723,I676632);
nand I_39599 (I676340,I676615,I676762);
not I_39600 (I676793,I676723);
nor I_39601 (I676810,I676793,I676533);
DFFARX1 I_39602 (I676810,I3563,I676363,I676352,);
nor I_39603 (I676841,I821608,I821599);
or I_39604 (I676343,I676590,I676841);
nor I_39605 (I676334,I676723,I676841);
or I_39606 (I676337,I676457,I676841);
DFFARX1 I_39607 (I676841,I3563,I676363,I676355,);
not I_39608 (I676941,I3570);
DFFARX1 I_39609 (I825827,I3563,I676941,I676967,);
not I_39610 (I676975,I676967);
nand I_39611 (I676992,I825815,I825833);
and I_39612 (I677009,I676992,I825830);
DFFARX1 I_39613 (I677009,I3563,I676941,I677035,);
not I_39614 (I677043,I825821);
DFFARX1 I_39615 (I825818,I3563,I676941,I677069,);
not I_39616 (I677077,I677069);
nor I_39617 (I677094,I677077,I676975);
and I_39618 (I677111,I677094,I825821);
nor I_39619 (I677128,I677077,I677043);
nor I_39620 (I676924,I677035,I677128);
DFFARX1 I_39621 (I825812,I3563,I676941,I677168,);
nor I_39622 (I677176,I677168,I677035);
not I_39623 (I677193,I677176);
not I_39624 (I677210,I677168);
nor I_39625 (I677227,I677210,I677111);
DFFARX1 I_39626 (I677227,I3563,I676941,I676927,);
nand I_39627 (I677258,I825812,I825815);
and I_39628 (I677275,I677258,I825818);
DFFARX1 I_39629 (I677275,I3563,I676941,I677301,);
nor I_39630 (I677309,I677301,I677168);
DFFARX1 I_39631 (I677309,I3563,I676941,I676909,);
nand I_39632 (I677340,I677301,I677210);
nand I_39633 (I676918,I677193,I677340);
not I_39634 (I677371,I677301);
nor I_39635 (I677388,I677371,I677111);
DFFARX1 I_39636 (I677388,I3563,I676941,I676930,);
nor I_39637 (I677419,I825824,I825815);
or I_39638 (I676921,I677168,I677419);
nor I_39639 (I676912,I677301,I677419);
or I_39640 (I676915,I677035,I677419);
DFFARX1 I_39641 (I677419,I3563,I676941,I676933,);
not I_39642 (I677519,I3570);
DFFARX1 I_39643 (I239873,I3563,I677519,I677545,);
not I_39644 (I677553,I677545);
nand I_39645 (I677570,I239876,I239897);
and I_39646 (I677587,I677570,I239885);
DFFARX1 I_39647 (I677587,I3563,I677519,I677613,);
not I_39648 (I677621,I239882);
DFFARX1 I_39649 (I239873,I3563,I677519,I677647,);
not I_39650 (I677655,I677647);
nor I_39651 (I677672,I677655,I677553);
and I_39652 (I677689,I677672,I239882);
nor I_39653 (I677706,I677655,I677621);
nor I_39654 (I677502,I677613,I677706);
DFFARX1 I_39655 (I239891,I3563,I677519,I677746,);
nor I_39656 (I677754,I677746,I677613);
not I_39657 (I677771,I677754);
not I_39658 (I677788,I677746);
nor I_39659 (I677805,I677788,I677689);
DFFARX1 I_39660 (I677805,I3563,I677519,I677505,);
nand I_39661 (I677836,I239876,I239879);
and I_39662 (I677853,I677836,I239888);
DFFARX1 I_39663 (I677853,I3563,I677519,I677879,);
nor I_39664 (I677887,I677879,I677746);
DFFARX1 I_39665 (I677887,I3563,I677519,I677487,);
nand I_39666 (I677918,I677879,I677788);
nand I_39667 (I677496,I677771,I677918);
not I_39668 (I677949,I677879);
nor I_39669 (I677966,I677949,I677689);
DFFARX1 I_39670 (I677966,I3563,I677519,I677508,);
nor I_39671 (I677997,I239894,I239879);
or I_39672 (I677499,I677746,I677997);
nor I_39673 (I677490,I677879,I677997);
or I_39674 (I677493,I677613,I677997);
DFFARX1 I_39675 (I677997,I3563,I677519,I677511,);
not I_39676 (I678097,I3570);
DFFARX1 I_39677 (I377614,I3563,I678097,I678123,);
not I_39678 (I678131,I678123);
nand I_39679 (I678148,I377617,I377593);
and I_39680 (I678165,I678148,I377590);
DFFARX1 I_39681 (I678165,I3563,I678097,I678191,);
not I_39682 (I678199,I377596);
DFFARX1 I_39683 (I377590,I3563,I678097,I678225,);
not I_39684 (I678233,I678225);
nor I_39685 (I678250,I678233,I678131);
and I_39686 (I678267,I678250,I377596);
nor I_39687 (I678284,I678233,I678199);
nor I_39688 (I678080,I678191,I678284);
DFFARX1 I_39689 (I377599,I3563,I678097,I678324,);
nor I_39690 (I678332,I678324,I678191);
not I_39691 (I678349,I678332);
not I_39692 (I678366,I678324);
nor I_39693 (I678383,I678366,I678267);
DFFARX1 I_39694 (I678383,I3563,I678097,I678083,);
nand I_39695 (I678414,I377602,I377611);
and I_39696 (I678431,I678414,I377608);
DFFARX1 I_39697 (I678431,I3563,I678097,I678457,);
nor I_39698 (I678465,I678457,I678324);
DFFARX1 I_39699 (I678465,I3563,I678097,I678065,);
nand I_39700 (I678496,I678457,I678366);
nand I_39701 (I678074,I678349,I678496);
not I_39702 (I678527,I678457);
nor I_39703 (I678544,I678527,I678267);
DFFARX1 I_39704 (I678544,I3563,I678097,I678086,);
nor I_39705 (I678575,I377605,I377611);
or I_39706 (I678077,I678324,I678575);
nor I_39707 (I678068,I678457,I678575);
or I_39708 (I678071,I678191,I678575);
DFFARX1 I_39709 (I678575,I3563,I678097,I678089,);
not I_39710 (I678675,I3570);
DFFARX1 I_39711 (I21877,I3563,I678675,I678701,);
not I_39712 (I678709,I678701);
nand I_39713 (I678726,I21874,I21865);
and I_39714 (I678743,I678726,I21865);
DFFARX1 I_39715 (I678743,I3563,I678675,I678769,);
not I_39716 (I678777,I21868);
DFFARX1 I_39717 (I21883,I3563,I678675,I678803,);
not I_39718 (I678811,I678803);
nor I_39719 (I678828,I678811,I678709);
and I_39720 (I678845,I678828,I21868);
nor I_39721 (I678862,I678811,I678777);
nor I_39722 (I678658,I678769,I678862);
DFFARX1 I_39723 (I21868,I3563,I678675,I678902,);
nor I_39724 (I678910,I678902,I678769);
not I_39725 (I678927,I678910);
not I_39726 (I678944,I678902);
nor I_39727 (I678961,I678944,I678845);
DFFARX1 I_39728 (I678961,I3563,I678675,I678661,);
nand I_39729 (I678992,I21886,I21871);
and I_39730 (I679009,I678992,I21889);
DFFARX1 I_39731 (I679009,I3563,I678675,I679035,);
nor I_39732 (I679043,I679035,I678902);
DFFARX1 I_39733 (I679043,I3563,I678675,I678643,);
nand I_39734 (I679074,I679035,I678944);
nand I_39735 (I678652,I678927,I679074);
not I_39736 (I679105,I679035);
nor I_39737 (I679122,I679105,I678845);
DFFARX1 I_39738 (I679122,I3563,I678675,I678664,);
nor I_39739 (I679153,I21880,I21871);
or I_39740 (I678655,I678902,I679153);
nor I_39741 (I678646,I679035,I679153);
or I_39742 (I678649,I678769,I679153);
DFFARX1 I_39743 (I679153,I3563,I678675,I678667,);
not I_39744 (I679253,I3570);
DFFARX1 I_39745 (I525227,I3563,I679253,I679279,);
not I_39746 (I679287,I679279);
nand I_39747 (I679304,I525218,I525236);
and I_39748 (I679321,I679304,I525239);
DFFARX1 I_39749 (I679321,I3563,I679253,I679347,);
not I_39750 (I679355,I525233);
DFFARX1 I_39751 (I525221,I3563,I679253,I679381,);
not I_39752 (I679389,I679381);
nor I_39753 (I679406,I679389,I679287);
and I_39754 (I679423,I679406,I525233);
nor I_39755 (I679440,I679389,I679355);
nor I_39756 (I679236,I679347,I679440);
DFFARX1 I_39757 (I525230,I3563,I679253,I679480,);
nor I_39758 (I679488,I679480,I679347);
not I_39759 (I679505,I679488);
not I_39760 (I679522,I679480);
nor I_39761 (I679539,I679522,I679423);
DFFARX1 I_39762 (I679539,I3563,I679253,I679239,);
nand I_39763 (I679570,I525245,I525242);
and I_39764 (I679587,I679570,I525224);
DFFARX1 I_39765 (I679587,I3563,I679253,I679613,);
nor I_39766 (I679621,I679613,I679480);
DFFARX1 I_39767 (I679621,I3563,I679253,I679221,);
nand I_39768 (I679652,I679613,I679522);
nand I_39769 (I679230,I679505,I679652);
not I_39770 (I679683,I679613);
nor I_39771 (I679700,I679683,I679423);
DFFARX1 I_39772 (I679700,I3563,I679253,I679242,);
nor I_39773 (I679731,I525218,I525242);
or I_39774 (I679233,I679480,I679731);
nor I_39775 (I679224,I679613,I679731);
or I_39776 (I679227,I679347,I679731);
DFFARX1 I_39777 (I679731,I3563,I679253,I679245,);
not I_39778 (I679831,I3570);
DFFARX1 I_39779 (I1251849,I3563,I679831,I679857,);
not I_39780 (I679865,I679857);
nand I_39781 (I679882,I1251852,I1251861);
and I_39782 (I679899,I679882,I1251864);
DFFARX1 I_39783 (I679899,I3563,I679831,I679925,);
not I_39784 (I679933,I1251873);
DFFARX1 I_39785 (I1251855,I3563,I679831,I679959,);
not I_39786 (I679967,I679959);
nor I_39787 (I679984,I679967,I679865);
and I_39788 (I680001,I679984,I1251873);
nor I_39789 (I680018,I679967,I679933);
nor I_39790 (I679814,I679925,I680018);
DFFARX1 I_39791 (I1251852,I3563,I679831,I680058,);
nor I_39792 (I680066,I680058,I679925);
not I_39793 (I680083,I680066);
not I_39794 (I680100,I680058);
nor I_39795 (I680117,I680100,I680001);
DFFARX1 I_39796 (I680117,I3563,I679831,I679817,);
nand I_39797 (I680148,I1251870,I1251849);
and I_39798 (I680165,I680148,I1251867);
DFFARX1 I_39799 (I680165,I3563,I679831,I680191,);
nor I_39800 (I680199,I680191,I680058);
DFFARX1 I_39801 (I680199,I3563,I679831,I679799,);
nand I_39802 (I680230,I680191,I680100);
nand I_39803 (I679808,I680083,I680230);
not I_39804 (I680261,I680191);
nor I_39805 (I680278,I680261,I680001);
DFFARX1 I_39806 (I680278,I3563,I679831,I679820,);
nor I_39807 (I680309,I1251858,I1251849);
or I_39808 (I679811,I680058,I680309);
nor I_39809 (I679802,I680191,I680309);
or I_39810 (I679805,I679925,I680309);
DFFARX1 I_39811 (I680309,I3563,I679831,I679823,);
not I_39812 (I680409,I3570);
DFFARX1 I_39813 (I499115,I3563,I680409,I680435,);
not I_39814 (I680443,I680435);
nand I_39815 (I680460,I499106,I499124);
and I_39816 (I680477,I680460,I499127);
DFFARX1 I_39817 (I680477,I3563,I680409,I680503,);
not I_39818 (I680511,I499121);
DFFARX1 I_39819 (I499109,I3563,I680409,I680537,);
not I_39820 (I680545,I680537);
nor I_39821 (I680562,I680545,I680443);
and I_39822 (I680579,I680562,I499121);
nor I_39823 (I680596,I680545,I680511);
nor I_39824 (I680392,I680503,I680596);
DFFARX1 I_39825 (I499118,I3563,I680409,I680636,);
nor I_39826 (I680644,I680636,I680503);
not I_39827 (I680661,I680644);
not I_39828 (I680678,I680636);
nor I_39829 (I680695,I680678,I680579);
DFFARX1 I_39830 (I680695,I3563,I680409,I680395,);
nand I_39831 (I680726,I499133,I499130);
and I_39832 (I680743,I680726,I499112);
DFFARX1 I_39833 (I680743,I3563,I680409,I680769,);
nor I_39834 (I680777,I680769,I680636);
DFFARX1 I_39835 (I680777,I3563,I680409,I680377,);
nand I_39836 (I680808,I680769,I680678);
nand I_39837 (I680386,I680661,I680808);
not I_39838 (I680839,I680769);
nor I_39839 (I680856,I680839,I680579);
DFFARX1 I_39840 (I680856,I3563,I680409,I680398,);
nor I_39841 (I680887,I499106,I499130);
or I_39842 (I680389,I680636,I680887);
nor I_39843 (I680380,I680769,I680887);
or I_39844 (I680383,I680503,I680887);
DFFARX1 I_39845 (I680887,I3563,I680409,I680401,);
not I_39846 (I680987,I3570);
DFFARX1 I_39847 (I958827,I3563,I680987,I681013,);
not I_39848 (I681021,I681013);
nand I_39849 (I681038,I958803,I958818);
and I_39850 (I681055,I681038,I958830);
DFFARX1 I_39851 (I681055,I3563,I680987,I681081,);
not I_39852 (I681089,I958815);
DFFARX1 I_39853 (I958806,I3563,I680987,I681115,);
not I_39854 (I681123,I681115);
nor I_39855 (I681140,I681123,I681021);
and I_39856 (I681157,I681140,I958815);
nor I_39857 (I681174,I681123,I681089);
nor I_39858 (I680970,I681081,I681174);
DFFARX1 I_39859 (I958803,I3563,I680987,I681214,);
nor I_39860 (I681222,I681214,I681081);
not I_39861 (I681239,I681222);
not I_39862 (I681256,I681214);
nor I_39863 (I681273,I681256,I681157);
DFFARX1 I_39864 (I681273,I3563,I680987,I680973,);
nand I_39865 (I681304,I958821,I958812);
and I_39866 (I681321,I681304,I958824);
DFFARX1 I_39867 (I681321,I3563,I680987,I681347,);
nor I_39868 (I681355,I681347,I681214);
DFFARX1 I_39869 (I681355,I3563,I680987,I680955,);
nand I_39870 (I681386,I681347,I681256);
nand I_39871 (I680964,I681239,I681386);
not I_39872 (I681417,I681347);
nor I_39873 (I681434,I681417,I681157);
DFFARX1 I_39874 (I681434,I3563,I680987,I680976,);
nor I_39875 (I681465,I958809,I958812);
or I_39876 (I680967,I681214,I681465);
nor I_39877 (I680958,I681347,I681465);
or I_39878 (I680961,I681081,I681465);
DFFARX1 I_39879 (I681465,I3563,I680987,I680979,);
not I_39880 (I681565,I3570);
DFFARX1 I_39881 (I1344645,I3563,I681565,I681591,);
not I_39882 (I681599,I681591);
nand I_39883 (I681616,I1344630,I1344618);
and I_39884 (I681633,I681616,I1344633);
DFFARX1 I_39885 (I681633,I3563,I681565,I681659,);
not I_39886 (I681667,I1344618);
DFFARX1 I_39887 (I1344636,I3563,I681565,I681693,);
not I_39888 (I681701,I681693);
nor I_39889 (I681718,I681701,I681599);
and I_39890 (I681735,I681718,I1344618);
nor I_39891 (I681752,I681701,I681667);
nor I_39892 (I681548,I681659,I681752);
DFFARX1 I_39893 (I1344624,I3563,I681565,I681792,);
nor I_39894 (I681800,I681792,I681659);
not I_39895 (I681817,I681800);
not I_39896 (I681834,I681792);
nor I_39897 (I681851,I681834,I681735);
DFFARX1 I_39898 (I681851,I3563,I681565,I681551,);
nand I_39899 (I681882,I1344621,I1344627);
and I_39900 (I681899,I681882,I1344642);
DFFARX1 I_39901 (I681899,I3563,I681565,I681925,);
nor I_39902 (I681933,I681925,I681792);
DFFARX1 I_39903 (I681933,I3563,I681565,I681533,);
nand I_39904 (I681964,I681925,I681834);
nand I_39905 (I681542,I681817,I681964);
not I_39906 (I681995,I681925);
nor I_39907 (I682012,I681995,I681735);
DFFARX1 I_39908 (I682012,I3563,I681565,I681554,);
nor I_39909 (I682043,I1344639,I1344627);
or I_39910 (I681545,I681792,I682043);
nor I_39911 (I681536,I681925,I682043);
or I_39912 (I681539,I681659,I682043);
DFFARX1 I_39913 (I682043,I3563,I681565,I681557,);
not I_39914 (I682143,I3570);
DFFARX1 I_39915 (I2756,I3563,I682143,I682169,);
not I_39916 (I682177,I682169);
nand I_39917 (I682194,I2156,I1572);
and I_39918 (I682211,I682194,I2012);
DFFARX1 I_39919 (I682211,I3563,I682143,I682237,);
not I_39920 (I682245,I1668);
DFFARX1 I_39921 (I2252,I3563,I682143,I682271,);
not I_39922 (I682279,I682271);
nor I_39923 (I682296,I682279,I682177);
and I_39924 (I682313,I682296,I1668);
nor I_39925 (I682330,I682279,I682245);
nor I_39926 (I682126,I682237,I682330);
DFFARX1 I_39927 (I1508,I3563,I682143,I682370,);
nor I_39928 (I682378,I682370,I682237);
not I_39929 (I682395,I682378);
not I_39930 (I682412,I682370);
nor I_39931 (I682429,I682412,I682313);
DFFARX1 I_39932 (I682429,I3563,I682143,I682129,);
nand I_39933 (I682460,I1932,I3188);
and I_39934 (I682477,I682460,I3404);
DFFARX1 I_39935 (I682477,I3563,I682143,I682503,);
nor I_39936 (I682511,I682503,I682370);
DFFARX1 I_39937 (I682511,I3563,I682143,I682111,);
nand I_39938 (I682542,I682503,I682412);
nand I_39939 (I682120,I682395,I682542);
not I_39940 (I682573,I682503);
nor I_39941 (I682590,I682573,I682313);
DFFARX1 I_39942 (I682590,I3563,I682143,I682132,);
nor I_39943 (I682621,I2116,I3188);
or I_39944 (I682123,I682370,I682621);
nor I_39945 (I682114,I682503,I682621);
or I_39946 (I682117,I682237,I682621);
DFFARX1 I_39947 (I682621,I3563,I682143,I682135,);
not I_39948 (I682721,I3570);
DFFARX1 I_39949 (I153091,I3563,I682721,I682747,);
not I_39950 (I682755,I682747);
nand I_39951 (I682772,I153100,I153109);
and I_39952 (I682789,I682772,I153088);
DFFARX1 I_39953 (I682789,I3563,I682721,I682815,);
not I_39954 (I682823,I153091);
DFFARX1 I_39955 (I153106,I3563,I682721,I682849,);
not I_39956 (I682857,I682849);
nor I_39957 (I682874,I682857,I682755);
and I_39958 (I682891,I682874,I153091);
nor I_39959 (I682908,I682857,I682823);
nor I_39960 (I682704,I682815,I682908);
DFFARX1 I_39961 (I153097,I3563,I682721,I682948,);
nor I_39962 (I682956,I682948,I682815);
not I_39963 (I682973,I682956);
not I_39964 (I682990,I682948);
nor I_39965 (I683007,I682990,I682891);
DFFARX1 I_39966 (I683007,I3563,I682721,I682707,);
nand I_39967 (I683038,I153112,I153088);
and I_39968 (I683055,I683038,I153094);
DFFARX1 I_39969 (I683055,I3563,I682721,I683081,);
nor I_39970 (I683089,I683081,I682948);
DFFARX1 I_39971 (I683089,I3563,I682721,I682689,);
nand I_39972 (I683120,I683081,I682990);
nand I_39973 (I682698,I682973,I683120);
not I_39974 (I683151,I683081);
nor I_39975 (I683168,I683151,I682891);
DFFARX1 I_39976 (I683168,I3563,I682721,I682710,);
nor I_39977 (I683199,I153103,I153088);
or I_39978 (I682701,I682948,I683199);
nor I_39979 (I682692,I683081,I683199);
or I_39980 (I682695,I682815,I683199);
DFFARX1 I_39981 (I683199,I3563,I682721,I682713,);
not I_39982 (I683299,I3570);
DFFARX1 I_39983 (I436555,I3563,I683299,I683325,);
not I_39984 (I683333,I683325);
nand I_39985 (I683350,I436546,I436564);
and I_39986 (I683367,I683350,I436567);
DFFARX1 I_39987 (I683367,I3563,I683299,I683393,);
not I_39988 (I683401,I436561);
DFFARX1 I_39989 (I436549,I3563,I683299,I683427,);
not I_39990 (I683435,I683427);
nor I_39991 (I683452,I683435,I683333);
and I_39992 (I683469,I683452,I436561);
nor I_39993 (I683486,I683435,I683401);
nor I_39994 (I683282,I683393,I683486);
DFFARX1 I_39995 (I436558,I3563,I683299,I683526,);
nor I_39996 (I683534,I683526,I683393);
not I_39997 (I683551,I683534);
not I_39998 (I683568,I683526);
nor I_39999 (I683585,I683568,I683469);
DFFARX1 I_40000 (I683585,I3563,I683299,I683285,);
nand I_40001 (I683616,I436573,I436570);
and I_40002 (I683633,I683616,I436552);
DFFARX1 I_40003 (I683633,I3563,I683299,I683659,);
nor I_40004 (I683667,I683659,I683526);
DFFARX1 I_40005 (I683667,I3563,I683299,I683267,);
nand I_40006 (I683698,I683659,I683568);
nand I_40007 (I683276,I683551,I683698);
not I_40008 (I683729,I683659);
nor I_40009 (I683746,I683729,I683469);
DFFARX1 I_40010 (I683746,I3563,I683299,I683288,);
nor I_40011 (I683777,I436546,I436570);
or I_40012 (I683279,I683526,I683777);
nor I_40013 (I683270,I683659,I683777);
or I_40014 (I683273,I683393,I683777);
DFFARX1 I_40015 (I683777,I3563,I683299,I683291,);
not I_40016 (I683877,I3570);
DFFARX1 I_40017 (I1275241,I3563,I683877,I683903,);
not I_40018 (I683911,I683903);
nand I_40019 (I683928,I1275244,I1275253);
and I_40020 (I683945,I683928,I1275256);
DFFARX1 I_40021 (I683945,I3563,I683877,I683971,);
not I_40022 (I683979,I1275265);
DFFARX1 I_40023 (I1275247,I3563,I683877,I684005,);
not I_40024 (I684013,I684005);
nor I_40025 (I684030,I684013,I683911);
and I_40026 (I684047,I684030,I1275265);
nor I_40027 (I684064,I684013,I683979);
nor I_40028 (I683860,I683971,I684064);
DFFARX1 I_40029 (I1275244,I3563,I683877,I684104,);
nor I_40030 (I684112,I684104,I683971);
not I_40031 (I684129,I684112);
not I_40032 (I684146,I684104);
nor I_40033 (I684163,I684146,I684047);
DFFARX1 I_40034 (I684163,I3563,I683877,I683863,);
nand I_40035 (I684194,I1275262,I1275241);
and I_40036 (I684211,I684194,I1275259);
DFFARX1 I_40037 (I684211,I3563,I683877,I684237,);
nor I_40038 (I684245,I684237,I684104);
DFFARX1 I_40039 (I684245,I3563,I683877,I683845,);
nand I_40040 (I684276,I684237,I684146);
nand I_40041 (I683854,I684129,I684276);
not I_40042 (I684307,I684237);
nor I_40043 (I684324,I684307,I684047);
DFFARX1 I_40044 (I684324,I3563,I683877,I683866,);
nor I_40045 (I684355,I1275250,I1275241);
or I_40046 (I683857,I684104,I684355);
nor I_40047 (I683848,I684237,I684355);
or I_40048 (I683851,I683971,I684355);
DFFARX1 I_40049 (I684355,I3563,I683877,I683869,);
not I_40050 (I684455,I3570);
DFFARX1 I_40051 (I1128005,I3563,I684455,I684481,);
not I_40052 (I684489,I684481);
nand I_40053 (I684506,I1127987,I1127999);
and I_40054 (I684523,I684506,I1128002);
DFFARX1 I_40055 (I684523,I3563,I684455,I684549,);
not I_40056 (I684557,I1127996);
DFFARX1 I_40057 (I1127993,I3563,I684455,I684583,);
not I_40058 (I684591,I684583);
nor I_40059 (I684608,I684591,I684489);
and I_40060 (I684625,I684608,I1127996);
nor I_40061 (I684642,I684591,I684557);
nor I_40062 (I684438,I684549,I684642);
DFFARX1 I_40063 (I1128011,I3563,I684455,I684682,);
nor I_40064 (I684690,I684682,I684549);
not I_40065 (I684707,I684690);
not I_40066 (I684724,I684682);
nor I_40067 (I684741,I684724,I684625);
DFFARX1 I_40068 (I684741,I3563,I684455,I684441,);
nand I_40069 (I684772,I1127990,I1127990);
and I_40070 (I684789,I684772,I1127987);
DFFARX1 I_40071 (I684789,I3563,I684455,I684815,);
nor I_40072 (I684823,I684815,I684682);
DFFARX1 I_40073 (I684823,I3563,I684455,I684423,);
nand I_40074 (I684854,I684815,I684724);
nand I_40075 (I684432,I684707,I684854);
not I_40076 (I684885,I684815);
nor I_40077 (I684902,I684885,I684625);
DFFARX1 I_40078 (I684902,I3563,I684455,I684444,);
nor I_40079 (I684933,I1128008,I1127990);
or I_40080 (I684435,I684682,I684933);
nor I_40081 (I684426,I684815,I684933);
or I_40082 (I684429,I684549,I684933);
DFFARX1 I_40083 (I684933,I3563,I684455,I684447,);
not I_40084 (I685033,I3570);
DFFARX1 I_40085 (I493675,I3563,I685033,I685059,);
not I_40086 (I685067,I685059);
nand I_40087 (I685084,I493666,I493684);
and I_40088 (I685101,I685084,I493687);
DFFARX1 I_40089 (I685101,I3563,I685033,I685127,);
not I_40090 (I685135,I493681);
DFFARX1 I_40091 (I493669,I3563,I685033,I685161,);
not I_40092 (I685169,I685161);
nor I_40093 (I685186,I685169,I685067);
and I_40094 (I685203,I685186,I493681);
nor I_40095 (I685220,I685169,I685135);
nor I_40096 (I685016,I685127,I685220);
DFFARX1 I_40097 (I493678,I3563,I685033,I685260,);
nor I_40098 (I685268,I685260,I685127);
not I_40099 (I685285,I685268);
not I_40100 (I685302,I685260);
nor I_40101 (I685319,I685302,I685203);
DFFARX1 I_40102 (I685319,I3563,I685033,I685019,);
nand I_40103 (I685350,I493693,I493690);
and I_40104 (I685367,I685350,I493672);
DFFARX1 I_40105 (I685367,I3563,I685033,I685393,);
nor I_40106 (I685401,I685393,I685260);
DFFARX1 I_40107 (I685401,I3563,I685033,I685001,);
nand I_40108 (I685432,I685393,I685302);
nand I_40109 (I685010,I685285,I685432);
not I_40110 (I685463,I685393);
nor I_40111 (I685480,I685463,I685203);
DFFARX1 I_40112 (I685480,I3563,I685033,I685022,);
nor I_40113 (I685511,I493666,I493690);
or I_40114 (I685013,I685260,I685511);
nor I_40115 (I685004,I685393,I685511);
or I_40116 (I685007,I685127,I685511);
DFFARX1 I_40117 (I685511,I3563,I685033,I685025,);
not I_40118 (I685611,I3570);
DFFARX1 I_40119 (I1334530,I3563,I685611,I685637,);
not I_40120 (I685645,I685637);
nand I_40121 (I685662,I1334515,I1334503);
and I_40122 (I685679,I685662,I1334518);
DFFARX1 I_40123 (I685679,I3563,I685611,I685705,);
not I_40124 (I685713,I1334503);
DFFARX1 I_40125 (I1334521,I3563,I685611,I685739,);
not I_40126 (I685747,I685739);
nor I_40127 (I685764,I685747,I685645);
and I_40128 (I685781,I685764,I1334503);
nor I_40129 (I685798,I685747,I685713);
nor I_40130 (I685594,I685705,I685798);
DFFARX1 I_40131 (I1334509,I3563,I685611,I685838,);
nor I_40132 (I685846,I685838,I685705);
not I_40133 (I685863,I685846);
not I_40134 (I685880,I685838);
nor I_40135 (I685897,I685880,I685781);
DFFARX1 I_40136 (I685897,I3563,I685611,I685597,);
nand I_40137 (I685928,I1334506,I1334512);
and I_40138 (I685945,I685928,I1334527);
DFFARX1 I_40139 (I685945,I3563,I685611,I685971,);
nor I_40140 (I685979,I685971,I685838);
DFFARX1 I_40141 (I685979,I3563,I685611,I685579,);
nand I_40142 (I686010,I685971,I685880);
nand I_40143 (I685588,I685863,I686010);
not I_40144 (I686041,I685971);
nor I_40145 (I686058,I686041,I685781);
DFFARX1 I_40146 (I686058,I3563,I685611,I685600,);
nor I_40147 (I686089,I1334524,I1334512);
or I_40148 (I685591,I685838,I686089);
nor I_40149 (I685582,I685971,I686089);
or I_40150 (I685585,I685705,I686089);
DFFARX1 I_40151 (I686089,I3563,I685611,I685603,);
not I_40152 (I686189,I3570);
DFFARX1 I_40153 (I847961,I3563,I686189,I686215,);
not I_40154 (I686223,I686215);
nand I_40155 (I686240,I847949,I847967);
and I_40156 (I686257,I686240,I847964);
DFFARX1 I_40157 (I686257,I3563,I686189,I686283,);
not I_40158 (I686291,I847955);
DFFARX1 I_40159 (I847952,I3563,I686189,I686317,);
not I_40160 (I686325,I686317);
nor I_40161 (I686342,I686325,I686223);
and I_40162 (I686359,I686342,I847955);
nor I_40163 (I686376,I686325,I686291);
nor I_40164 (I686172,I686283,I686376);
DFFARX1 I_40165 (I847946,I3563,I686189,I686416,);
nor I_40166 (I686424,I686416,I686283);
not I_40167 (I686441,I686424);
not I_40168 (I686458,I686416);
nor I_40169 (I686475,I686458,I686359);
DFFARX1 I_40170 (I686475,I3563,I686189,I686175,);
nand I_40171 (I686506,I847946,I847949);
and I_40172 (I686523,I686506,I847952);
DFFARX1 I_40173 (I686523,I3563,I686189,I686549,);
nor I_40174 (I686557,I686549,I686416);
DFFARX1 I_40175 (I686557,I3563,I686189,I686157,);
nand I_40176 (I686588,I686549,I686458);
nand I_40177 (I686166,I686441,I686588);
not I_40178 (I686619,I686549);
nor I_40179 (I686636,I686619,I686359);
DFFARX1 I_40180 (I686636,I3563,I686189,I686178,);
nor I_40181 (I686667,I847958,I847949);
or I_40182 (I686169,I686416,I686667);
nor I_40183 (I686160,I686549,I686667);
or I_40184 (I686163,I686283,I686667);
DFFARX1 I_40185 (I686667,I3563,I686189,I686181,);
not I_40186 (I686767,I3570);
DFFARX1 I_40187 (I872730,I3563,I686767,I686793,);
not I_40188 (I686801,I686793);
nand I_40189 (I686818,I872718,I872736);
and I_40190 (I686835,I686818,I872733);
DFFARX1 I_40191 (I686835,I3563,I686767,I686861,);
not I_40192 (I686869,I872724);
DFFARX1 I_40193 (I872721,I3563,I686767,I686895,);
not I_40194 (I686903,I686895);
nor I_40195 (I686920,I686903,I686801);
and I_40196 (I686937,I686920,I872724);
nor I_40197 (I686954,I686903,I686869);
nor I_40198 (I686750,I686861,I686954);
DFFARX1 I_40199 (I872715,I3563,I686767,I686994,);
nor I_40200 (I687002,I686994,I686861);
not I_40201 (I687019,I687002);
not I_40202 (I687036,I686994);
nor I_40203 (I687053,I687036,I686937);
DFFARX1 I_40204 (I687053,I3563,I686767,I686753,);
nand I_40205 (I687084,I872715,I872718);
and I_40206 (I687101,I687084,I872721);
DFFARX1 I_40207 (I687101,I3563,I686767,I687127,);
nor I_40208 (I687135,I687127,I686994);
DFFARX1 I_40209 (I687135,I3563,I686767,I686735,);
nand I_40210 (I687166,I687127,I687036);
nand I_40211 (I686744,I687019,I687166);
not I_40212 (I687197,I687127);
nor I_40213 (I687214,I687197,I686937);
DFFARX1 I_40214 (I687214,I3563,I686767,I686756,);
nor I_40215 (I687245,I872727,I872718);
or I_40216 (I686747,I686994,I687245);
nor I_40217 (I686738,I687127,I687245);
or I_40218 (I686741,I686861,I687245);
DFFARX1 I_40219 (I687245,I3563,I686767,I686759,);
not I_40220 (I687345,I3570);
DFFARX1 I_40221 (I1268169,I3563,I687345,I687371,);
not I_40222 (I687379,I687371);
nand I_40223 (I687396,I1268172,I1268181);
and I_40224 (I687413,I687396,I1268184);
DFFARX1 I_40225 (I687413,I3563,I687345,I687439,);
not I_40226 (I687447,I1268193);
DFFARX1 I_40227 (I1268175,I3563,I687345,I687473,);
not I_40228 (I687481,I687473);
nor I_40229 (I687498,I687481,I687379);
and I_40230 (I687515,I687498,I1268193);
nor I_40231 (I687532,I687481,I687447);
nor I_40232 (I687328,I687439,I687532);
DFFARX1 I_40233 (I1268172,I3563,I687345,I687572,);
nor I_40234 (I687580,I687572,I687439);
not I_40235 (I687597,I687580);
not I_40236 (I687614,I687572);
nor I_40237 (I687631,I687614,I687515);
DFFARX1 I_40238 (I687631,I3563,I687345,I687331,);
nand I_40239 (I687662,I1268190,I1268169);
and I_40240 (I687679,I687662,I1268187);
DFFARX1 I_40241 (I687679,I3563,I687345,I687705,);
nor I_40242 (I687713,I687705,I687572);
DFFARX1 I_40243 (I687713,I3563,I687345,I687313,);
nand I_40244 (I687744,I687705,I687614);
nand I_40245 (I687322,I687597,I687744);
not I_40246 (I687775,I687705);
nor I_40247 (I687792,I687775,I687515);
DFFARX1 I_40248 (I687792,I3563,I687345,I687334,);
nor I_40249 (I687823,I1268178,I1268169);
or I_40250 (I687325,I687572,I687823);
nor I_40251 (I687316,I687705,I687823);
or I_40252 (I687319,I687439,I687823);
DFFARX1 I_40253 (I687823,I3563,I687345,I687337,);
not I_40254 (I687923,I3570);
DFFARX1 I_40255 (I1011799,I3563,I687923,I687949,);
not I_40256 (I687957,I687949);
nand I_40257 (I687974,I1011775,I1011790);
and I_40258 (I687991,I687974,I1011802);
DFFARX1 I_40259 (I687991,I3563,I687923,I688017,);
not I_40260 (I688025,I1011787);
DFFARX1 I_40261 (I1011778,I3563,I687923,I688051,);
not I_40262 (I688059,I688051);
nor I_40263 (I688076,I688059,I687957);
and I_40264 (I688093,I688076,I1011787);
nor I_40265 (I688110,I688059,I688025);
nor I_40266 (I687906,I688017,I688110);
DFFARX1 I_40267 (I1011775,I3563,I687923,I688150,);
nor I_40268 (I688158,I688150,I688017);
not I_40269 (I688175,I688158);
not I_40270 (I688192,I688150);
nor I_40271 (I688209,I688192,I688093);
DFFARX1 I_40272 (I688209,I3563,I687923,I687909,);
nand I_40273 (I688240,I1011793,I1011784);
and I_40274 (I688257,I688240,I1011796);
DFFARX1 I_40275 (I688257,I3563,I687923,I688283,);
nor I_40276 (I688291,I688283,I688150);
DFFARX1 I_40277 (I688291,I3563,I687923,I687891,);
nand I_40278 (I688322,I688283,I688192);
nand I_40279 (I687900,I688175,I688322);
not I_40280 (I688353,I688283);
nor I_40281 (I688370,I688353,I688093);
DFFARX1 I_40282 (I688370,I3563,I687923,I687912,);
nor I_40283 (I688401,I1011781,I1011784);
or I_40284 (I687903,I688150,I688401);
nor I_40285 (I687894,I688283,I688401);
or I_40286 (I687897,I688017,I688401);
DFFARX1 I_40287 (I688401,I3563,I687923,I687915,);
not I_40288 (I688501,I3570);
DFFARX1 I_40289 (I300145,I3563,I688501,I688527,);
not I_40290 (I688535,I688527);
nand I_40291 (I688552,I300148,I300124);
and I_40292 (I688569,I688552,I300121);
DFFARX1 I_40293 (I688569,I3563,I688501,I688595,);
not I_40294 (I688603,I300127);
DFFARX1 I_40295 (I300121,I3563,I688501,I688629,);
not I_40296 (I688637,I688629);
nor I_40297 (I688654,I688637,I688535);
and I_40298 (I688671,I688654,I300127);
nor I_40299 (I688688,I688637,I688603);
nor I_40300 (I688484,I688595,I688688);
DFFARX1 I_40301 (I300130,I3563,I688501,I688728,);
nor I_40302 (I688736,I688728,I688595);
not I_40303 (I688753,I688736);
not I_40304 (I688770,I688728);
nor I_40305 (I688787,I688770,I688671);
DFFARX1 I_40306 (I688787,I3563,I688501,I688487,);
nand I_40307 (I688818,I300133,I300142);
and I_40308 (I688835,I688818,I300139);
DFFARX1 I_40309 (I688835,I3563,I688501,I688861,);
nor I_40310 (I688869,I688861,I688728);
DFFARX1 I_40311 (I688869,I3563,I688501,I688469,);
nand I_40312 (I688900,I688861,I688770);
nand I_40313 (I688478,I688753,I688900);
not I_40314 (I688931,I688861);
nor I_40315 (I688948,I688931,I688671);
DFFARX1 I_40316 (I688948,I3563,I688501,I688490,);
nor I_40317 (I688979,I300136,I300142);
or I_40318 (I688481,I688728,I688979);
nor I_40319 (I688472,I688861,I688979);
or I_40320 (I688475,I688595,I688979);
DFFARX1 I_40321 (I688979,I3563,I688501,I688493,);
not I_40322 (I689079,I3570);
DFFARX1 I_40323 (I982083,I3563,I689079,I689105,);
not I_40324 (I689113,I689105);
nand I_40325 (I689130,I982059,I982074);
and I_40326 (I689147,I689130,I982086);
DFFARX1 I_40327 (I689147,I3563,I689079,I689173,);
not I_40328 (I689181,I982071);
DFFARX1 I_40329 (I982062,I3563,I689079,I689207,);
not I_40330 (I689215,I689207);
nor I_40331 (I689232,I689215,I689113);
and I_40332 (I689249,I689232,I982071);
nor I_40333 (I689266,I689215,I689181);
nor I_40334 (I689062,I689173,I689266);
DFFARX1 I_40335 (I982059,I3563,I689079,I689306,);
nor I_40336 (I689314,I689306,I689173);
not I_40337 (I689331,I689314);
not I_40338 (I689348,I689306);
nor I_40339 (I689365,I689348,I689249);
DFFARX1 I_40340 (I689365,I3563,I689079,I689065,);
nand I_40341 (I689396,I982077,I982068);
and I_40342 (I689413,I689396,I982080);
DFFARX1 I_40343 (I689413,I3563,I689079,I689439,);
nor I_40344 (I689447,I689439,I689306);
DFFARX1 I_40345 (I689447,I3563,I689079,I689047,);
nand I_40346 (I689478,I689439,I689348);
nand I_40347 (I689056,I689331,I689478);
not I_40348 (I689509,I689439);
nor I_40349 (I689526,I689509,I689249);
DFFARX1 I_40350 (I689526,I3563,I689079,I689068,);
nor I_40351 (I689557,I982065,I982068);
or I_40352 (I689059,I689306,I689557);
nor I_40353 (I689050,I689439,I689557);
or I_40354 (I689053,I689173,I689557);
DFFARX1 I_40355 (I689557,I3563,I689079,I689071,);
not I_40356 (I689657,I3570);
DFFARX1 I_40357 (I1043453,I3563,I689657,I689683,);
not I_40358 (I689691,I689683);
nand I_40359 (I689708,I1043429,I1043444);
and I_40360 (I689725,I689708,I1043456);
DFFARX1 I_40361 (I689725,I3563,I689657,I689751,);
not I_40362 (I689759,I1043441);
DFFARX1 I_40363 (I1043432,I3563,I689657,I689785,);
not I_40364 (I689793,I689785);
nor I_40365 (I689810,I689793,I689691);
and I_40366 (I689827,I689810,I1043441);
nor I_40367 (I689844,I689793,I689759);
nor I_40368 (I689640,I689751,I689844);
DFFARX1 I_40369 (I1043429,I3563,I689657,I689884,);
nor I_40370 (I689892,I689884,I689751);
not I_40371 (I689909,I689892);
not I_40372 (I689926,I689884);
nor I_40373 (I689943,I689926,I689827);
DFFARX1 I_40374 (I689943,I3563,I689657,I689643,);
nand I_40375 (I689974,I1043447,I1043438);
and I_40376 (I689991,I689974,I1043450);
DFFARX1 I_40377 (I689991,I3563,I689657,I690017,);
nor I_40378 (I690025,I690017,I689884);
DFFARX1 I_40379 (I690025,I3563,I689657,I689625,);
nand I_40380 (I690056,I690017,I689926);
nand I_40381 (I689634,I689909,I690056);
not I_40382 (I690087,I690017);
nor I_40383 (I690104,I690087,I689827);
DFFARX1 I_40384 (I690104,I3563,I689657,I689646,);
nor I_40385 (I690135,I1043435,I1043438);
or I_40386 (I689637,I689884,I690135);
nor I_40387 (I689628,I690017,I690135);
or I_40388 (I689631,I689751,I690135);
DFFARX1 I_40389 (I690135,I3563,I689657,I689649,);
not I_40390 (I690235,I3570);
DFFARX1 I_40391 (I925235,I3563,I690235,I690261,);
not I_40392 (I690269,I690261);
nand I_40393 (I690286,I925211,I925226);
and I_40394 (I690303,I690286,I925238);
DFFARX1 I_40395 (I690303,I3563,I690235,I690329,);
not I_40396 (I690337,I925223);
DFFARX1 I_40397 (I925214,I3563,I690235,I690363,);
not I_40398 (I690371,I690363);
nor I_40399 (I690388,I690371,I690269);
and I_40400 (I690405,I690388,I925223);
nor I_40401 (I690422,I690371,I690337);
nor I_40402 (I690218,I690329,I690422);
DFFARX1 I_40403 (I925211,I3563,I690235,I690462,);
nor I_40404 (I690470,I690462,I690329);
not I_40405 (I690487,I690470);
not I_40406 (I690504,I690462);
nor I_40407 (I690521,I690504,I690405);
DFFARX1 I_40408 (I690521,I3563,I690235,I690221,);
nand I_40409 (I690552,I925229,I925220);
and I_40410 (I690569,I690552,I925232);
DFFARX1 I_40411 (I690569,I3563,I690235,I690595,);
nor I_40412 (I690603,I690595,I690462);
DFFARX1 I_40413 (I690603,I3563,I690235,I690203,);
nand I_40414 (I690634,I690595,I690504);
nand I_40415 (I690212,I690487,I690634);
not I_40416 (I690665,I690595);
nor I_40417 (I690682,I690665,I690405);
DFFARX1 I_40418 (I690682,I3563,I690235,I690224,);
nor I_40419 (I690713,I925217,I925220);
or I_40420 (I690215,I690462,I690713);
nor I_40421 (I690206,I690595,I690713);
or I_40422 (I690209,I690329,I690713);
DFFARX1 I_40423 (I690713,I3563,I690235,I690227,);
not I_40424 (I690813,I3570);
DFFARX1 I_40425 (I471915,I3563,I690813,I690839,);
not I_40426 (I690847,I690839);
nand I_40427 (I690864,I471906,I471924);
and I_40428 (I690881,I690864,I471927);
DFFARX1 I_40429 (I690881,I3563,I690813,I690907,);
not I_40430 (I690915,I471921);
DFFARX1 I_40431 (I471909,I3563,I690813,I690941,);
not I_40432 (I690949,I690941);
nor I_40433 (I690966,I690949,I690847);
and I_40434 (I690983,I690966,I471921);
nor I_40435 (I691000,I690949,I690915);
nor I_40436 (I690796,I690907,I691000);
DFFARX1 I_40437 (I471918,I3563,I690813,I691040,);
nor I_40438 (I691048,I691040,I690907);
not I_40439 (I691065,I691048);
not I_40440 (I691082,I691040);
nor I_40441 (I691099,I691082,I690983);
DFFARX1 I_40442 (I691099,I3563,I690813,I690799,);
nand I_40443 (I691130,I471933,I471930);
and I_40444 (I691147,I691130,I471912);
DFFARX1 I_40445 (I691147,I3563,I690813,I691173,);
nor I_40446 (I691181,I691173,I691040);
DFFARX1 I_40447 (I691181,I3563,I690813,I690781,);
nand I_40448 (I691212,I691173,I691082);
nand I_40449 (I690790,I691065,I691212);
not I_40450 (I691243,I691173);
nor I_40451 (I691260,I691243,I690983);
DFFARX1 I_40452 (I691260,I3563,I690813,I690802,);
nor I_40453 (I691291,I471906,I471930);
or I_40454 (I690793,I691040,I691291);
nor I_40455 (I690784,I691173,I691291);
or I_40456 (I690787,I690907,I691291);
DFFARX1 I_40457 (I691291,I3563,I690813,I690805,);
not I_40458 (I691391,I3570);
DFFARX1 I_40459 (I346521,I3563,I691391,I691417,);
not I_40460 (I691425,I691417);
nand I_40461 (I691442,I346524,I346500);
and I_40462 (I691459,I691442,I346497);
DFFARX1 I_40463 (I691459,I3563,I691391,I691485,);
not I_40464 (I691493,I346503);
DFFARX1 I_40465 (I346497,I3563,I691391,I691519,);
not I_40466 (I691527,I691519);
nor I_40467 (I691544,I691527,I691425);
and I_40468 (I691561,I691544,I346503);
nor I_40469 (I691578,I691527,I691493);
nor I_40470 (I691374,I691485,I691578);
DFFARX1 I_40471 (I346506,I3563,I691391,I691618,);
nor I_40472 (I691626,I691618,I691485);
not I_40473 (I691643,I691626);
not I_40474 (I691660,I691618);
nor I_40475 (I691677,I691660,I691561);
DFFARX1 I_40476 (I691677,I3563,I691391,I691377,);
nand I_40477 (I691708,I346509,I346518);
and I_40478 (I691725,I691708,I346515);
DFFARX1 I_40479 (I691725,I3563,I691391,I691751,);
nor I_40480 (I691759,I691751,I691618);
DFFARX1 I_40481 (I691759,I3563,I691391,I691359,);
nand I_40482 (I691790,I691751,I691660);
nand I_40483 (I691368,I691643,I691790);
not I_40484 (I691821,I691751);
nor I_40485 (I691838,I691821,I691561);
DFFARX1 I_40486 (I691838,I3563,I691391,I691380,);
nor I_40487 (I691869,I346512,I346518);
or I_40488 (I691371,I691618,I691869);
nor I_40489 (I691362,I691751,I691869);
or I_40490 (I691365,I691485,I691869);
DFFARX1 I_40491 (I691869,I3563,I691391,I691383,);
not I_40492 (I691969,I3570);
DFFARX1 I_40493 (I234518,I3563,I691969,I691995,);
not I_40494 (I692003,I691995);
nand I_40495 (I692020,I234521,I234542);
and I_40496 (I692037,I692020,I234530);
DFFARX1 I_40497 (I692037,I3563,I691969,I692063,);
not I_40498 (I692071,I234527);
DFFARX1 I_40499 (I234518,I3563,I691969,I692097,);
not I_40500 (I692105,I692097);
nor I_40501 (I692122,I692105,I692003);
and I_40502 (I692139,I692122,I234527);
nor I_40503 (I692156,I692105,I692071);
nor I_40504 (I691952,I692063,I692156);
DFFARX1 I_40505 (I234536,I3563,I691969,I692196,);
nor I_40506 (I692204,I692196,I692063);
not I_40507 (I692221,I692204);
not I_40508 (I692238,I692196);
nor I_40509 (I692255,I692238,I692139);
DFFARX1 I_40510 (I692255,I3563,I691969,I691955,);
nand I_40511 (I692286,I234521,I234524);
and I_40512 (I692303,I692286,I234533);
DFFARX1 I_40513 (I692303,I3563,I691969,I692329,);
nor I_40514 (I692337,I692329,I692196);
DFFARX1 I_40515 (I692337,I3563,I691969,I691937,);
nand I_40516 (I692368,I692329,I692238);
nand I_40517 (I691946,I692221,I692368);
not I_40518 (I692399,I692329);
nor I_40519 (I692416,I692399,I692139);
DFFARX1 I_40520 (I692416,I3563,I691969,I691958,);
nor I_40521 (I692447,I234539,I234524);
or I_40522 (I691949,I692196,I692447);
nor I_40523 (I691940,I692329,I692447);
or I_40524 (I691943,I692063,I692447);
DFFARX1 I_40525 (I692447,I3563,I691969,I691961,);
not I_40526 (I692547,I3570);
DFFARX1 I_40527 (I1270889,I3563,I692547,I692573,);
not I_40528 (I692581,I692573);
nand I_40529 (I692598,I1270892,I1270901);
and I_40530 (I692615,I692598,I1270904);
DFFARX1 I_40531 (I692615,I3563,I692547,I692641,);
not I_40532 (I692649,I1270913);
DFFARX1 I_40533 (I1270895,I3563,I692547,I692675,);
not I_40534 (I692683,I692675);
nor I_40535 (I692700,I692683,I692581);
and I_40536 (I692717,I692700,I1270913);
nor I_40537 (I692734,I692683,I692649);
nor I_40538 (I692530,I692641,I692734);
DFFARX1 I_40539 (I1270892,I3563,I692547,I692774,);
nor I_40540 (I692782,I692774,I692641);
not I_40541 (I692799,I692782);
not I_40542 (I692816,I692774);
nor I_40543 (I692833,I692816,I692717);
DFFARX1 I_40544 (I692833,I3563,I692547,I692533,);
nand I_40545 (I692864,I1270910,I1270889);
and I_40546 (I692881,I692864,I1270907);
DFFARX1 I_40547 (I692881,I3563,I692547,I692907,);
nor I_40548 (I692915,I692907,I692774);
DFFARX1 I_40549 (I692915,I3563,I692547,I692515,);
nand I_40550 (I692946,I692907,I692816);
nand I_40551 (I692524,I692799,I692946);
not I_40552 (I692977,I692907);
nor I_40553 (I692994,I692977,I692717);
DFFARX1 I_40554 (I692994,I3563,I692547,I692536,);
nor I_40555 (I693025,I1270898,I1270889);
or I_40556 (I692527,I692774,I693025);
nor I_40557 (I692518,I692907,I693025);
or I_40558 (I692521,I692641,I693025);
DFFARX1 I_40559 (I693025,I3563,I692547,I692539,);
not I_40560 (I693125,I3570);
DFFARX1 I_40561 (I918129,I3563,I693125,I693151,);
not I_40562 (I693159,I693151);
nand I_40563 (I693176,I918105,I918120);
and I_40564 (I693193,I693176,I918132);
DFFARX1 I_40565 (I693193,I3563,I693125,I693219,);
not I_40566 (I693227,I918117);
DFFARX1 I_40567 (I918108,I3563,I693125,I693253,);
not I_40568 (I693261,I693253);
nor I_40569 (I693278,I693261,I693159);
and I_40570 (I693295,I693278,I918117);
nor I_40571 (I693312,I693261,I693227);
nor I_40572 (I693108,I693219,I693312);
DFFARX1 I_40573 (I918105,I3563,I693125,I693352,);
nor I_40574 (I693360,I693352,I693219);
not I_40575 (I693377,I693360);
not I_40576 (I693394,I693352);
nor I_40577 (I693411,I693394,I693295);
DFFARX1 I_40578 (I693411,I3563,I693125,I693111,);
nand I_40579 (I693442,I918123,I918114);
and I_40580 (I693459,I693442,I918126);
DFFARX1 I_40581 (I693459,I3563,I693125,I693485,);
nor I_40582 (I693493,I693485,I693352);
DFFARX1 I_40583 (I693493,I3563,I693125,I693093,);
nand I_40584 (I693524,I693485,I693394);
nand I_40585 (I693102,I693377,I693524);
not I_40586 (I693555,I693485);
nor I_40587 (I693572,I693555,I693295);
DFFARX1 I_40588 (I693572,I3563,I693125,I693114,);
nor I_40589 (I693603,I918111,I918114);
or I_40590 (I693105,I693352,I693603);
nor I_40591 (I693096,I693485,I693603);
or I_40592 (I693099,I693219,I693603);
DFFARX1 I_40593 (I693603,I3563,I693125,I693117,);
not I_40594 (I693703,I3570);
DFFARX1 I_40595 (I812125,I3563,I693703,I693729,);
not I_40596 (I693737,I693729);
nand I_40597 (I693754,I812113,I812131);
and I_40598 (I693771,I693754,I812128);
DFFARX1 I_40599 (I693771,I3563,I693703,I693797,);
not I_40600 (I693805,I812119);
DFFARX1 I_40601 (I812116,I3563,I693703,I693831,);
not I_40602 (I693839,I693831);
nor I_40603 (I693856,I693839,I693737);
and I_40604 (I693873,I693856,I812119);
nor I_40605 (I693890,I693839,I693805);
nor I_40606 (I693686,I693797,I693890);
DFFARX1 I_40607 (I812110,I3563,I693703,I693930,);
nor I_40608 (I693938,I693930,I693797);
not I_40609 (I693955,I693938);
not I_40610 (I693972,I693930);
nor I_40611 (I693989,I693972,I693873);
DFFARX1 I_40612 (I693989,I3563,I693703,I693689,);
nand I_40613 (I694020,I812110,I812113);
and I_40614 (I694037,I694020,I812116);
DFFARX1 I_40615 (I694037,I3563,I693703,I694063,);
nor I_40616 (I694071,I694063,I693930);
DFFARX1 I_40617 (I694071,I3563,I693703,I693671,);
nand I_40618 (I694102,I694063,I693972);
nand I_40619 (I693680,I693955,I694102);
not I_40620 (I694133,I694063);
nor I_40621 (I694150,I694133,I693873);
DFFARX1 I_40622 (I694150,I3563,I693703,I693692,);
nor I_40623 (I694181,I812122,I812113);
or I_40624 (I693683,I693930,I694181);
nor I_40625 (I693674,I694063,I694181);
or I_40626 (I693677,I693797,I694181);
DFFARX1 I_40627 (I694181,I3563,I693703,I693695,);
not I_40628 (I694281,I3570);
DFFARX1 I_40629 (I502379,I3563,I694281,I694307,);
not I_40630 (I694315,I694307);
nand I_40631 (I694332,I502370,I502388);
and I_40632 (I694349,I694332,I502391);
DFFARX1 I_40633 (I694349,I3563,I694281,I694375,);
not I_40634 (I694383,I502385);
DFFARX1 I_40635 (I502373,I3563,I694281,I694409,);
not I_40636 (I694417,I694409);
nor I_40637 (I694434,I694417,I694315);
and I_40638 (I694451,I694434,I502385);
nor I_40639 (I694468,I694417,I694383);
nor I_40640 (I694264,I694375,I694468);
DFFARX1 I_40641 (I502382,I3563,I694281,I694508,);
nor I_40642 (I694516,I694508,I694375);
not I_40643 (I694533,I694516);
not I_40644 (I694550,I694508);
nor I_40645 (I694567,I694550,I694451);
DFFARX1 I_40646 (I694567,I3563,I694281,I694267,);
nand I_40647 (I694598,I502397,I502394);
and I_40648 (I694615,I694598,I502376);
DFFARX1 I_40649 (I694615,I3563,I694281,I694641,);
nor I_40650 (I694649,I694641,I694508);
DFFARX1 I_40651 (I694649,I3563,I694281,I694249,);
nand I_40652 (I694680,I694641,I694550);
nand I_40653 (I694258,I694533,I694680);
not I_40654 (I694711,I694641);
nor I_40655 (I694728,I694711,I694451);
DFFARX1 I_40656 (I694728,I3563,I694281,I694270,);
nor I_40657 (I694759,I502370,I502394);
or I_40658 (I694261,I694508,I694759);
nor I_40659 (I694252,I694641,I694759);
or I_40660 (I694255,I694375,I694759);
DFFARX1 I_40661 (I694759,I3563,I694281,I694273,);
not I_40662 (I694859,I3570);
DFFARX1 I_40663 (I913309,I3563,I694859,I694885,);
not I_40664 (I694893,I694885);
nand I_40665 (I694910,I913297,I913315);
and I_40666 (I694927,I694910,I913312);
DFFARX1 I_40667 (I694927,I3563,I694859,I694953,);
not I_40668 (I694961,I913303);
DFFARX1 I_40669 (I913300,I3563,I694859,I694987,);
not I_40670 (I694995,I694987);
nor I_40671 (I695012,I694995,I694893);
and I_40672 (I695029,I695012,I913303);
nor I_40673 (I695046,I694995,I694961);
nor I_40674 (I694842,I694953,I695046);
DFFARX1 I_40675 (I913294,I3563,I694859,I695086,);
nor I_40676 (I695094,I695086,I694953);
not I_40677 (I695111,I695094);
not I_40678 (I695128,I695086);
nor I_40679 (I695145,I695128,I695029);
DFFARX1 I_40680 (I695145,I3563,I694859,I694845,);
nand I_40681 (I695176,I913294,I913297);
and I_40682 (I695193,I695176,I913300);
DFFARX1 I_40683 (I695193,I3563,I694859,I695219,);
nor I_40684 (I695227,I695219,I695086);
DFFARX1 I_40685 (I695227,I3563,I694859,I694827,);
nand I_40686 (I695258,I695219,I695128);
nand I_40687 (I694836,I695111,I695258);
not I_40688 (I695289,I695219);
nor I_40689 (I695306,I695289,I695029);
DFFARX1 I_40690 (I695306,I3563,I694859,I694848,);
nor I_40691 (I695337,I913306,I913297);
or I_40692 (I694839,I695086,I695337);
nor I_40693 (I694830,I695219,I695337);
or I_40694 (I694833,I694953,I695337);
DFFARX1 I_40695 (I695337,I3563,I694859,I694851,);
not I_40696 (I695437,I3570);
DFFARX1 I_40697 (I1065178,I3563,I695437,I695463,);
not I_40698 (I695471,I695463);
nand I_40699 (I695488,I1065175,I1065193);
and I_40700 (I695505,I695488,I1065190);
DFFARX1 I_40701 (I695505,I3563,I695437,I695531,);
not I_40702 (I695539,I1065172);
DFFARX1 I_40703 (I1065175,I3563,I695437,I695565,);
not I_40704 (I695573,I695565);
nor I_40705 (I695590,I695573,I695471);
and I_40706 (I695607,I695590,I1065172);
nor I_40707 (I695624,I695573,I695539);
nor I_40708 (I695420,I695531,I695624);
DFFARX1 I_40709 (I1065184,I3563,I695437,I695664,);
nor I_40710 (I695672,I695664,I695531);
not I_40711 (I695689,I695672);
not I_40712 (I695706,I695664);
nor I_40713 (I695723,I695706,I695607);
DFFARX1 I_40714 (I695723,I3563,I695437,I695423,);
nand I_40715 (I695754,I1065187,I1065172);
and I_40716 (I695771,I695754,I1065178);
DFFARX1 I_40717 (I695771,I3563,I695437,I695797,);
nor I_40718 (I695805,I695797,I695664);
DFFARX1 I_40719 (I695805,I3563,I695437,I695405,);
nand I_40720 (I695836,I695797,I695706);
nand I_40721 (I695414,I695689,I695836);
not I_40722 (I695867,I695797);
nor I_40723 (I695884,I695867,I695607);
DFFARX1 I_40724 (I695884,I3563,I695437,I695426,);
nor I_40725 (I695915,I1065181,I1065172);
or I_40726 (I695417,I695664,I695915);
nor I_40727 (I695408,I695797,I695915);
or I_40728 (I695411,I695531,I695915);
DFFARX1 I_40729 (I695915,I3563,I695437,I695429,);
not I_40730 (I696015,I3570);
DFFARX1 I_40731 (I610439,I3563,I696015,I696041,);
not I_40732 (I696049,I696041);
nand I_40733 (I696066,I610448,I610457);
and I_40734 (I696083,I696066,I610463);
DFFARX1 I_40735 (I696083,I3563,I696015,I696109,);
not I_40736 (I696117,I610460);
DFFARX1 I_40737 (I610445,I3563,I696015,I696143,);
not I_40738 (I696151,I696143);
nor I_40739 (I696168,I696151,I696049);
and I_40740 (I696185,I696168,I610460);
nor I_40741 (I696202,I696151,I696117);
nor I_40742 (I695998,I696109,I696202);
DFFARX1 I_40743 (I610454,I3563,I696015,I696242,);
nor I_40744 (I696250,I696242,I696109);
not I_40745 (I696267,I696250);
not I_40746 (I696284,I696242);
nor I_40747 (I696301,I696284,I696185);
DFFARX1 I_40748 (I696301,I3563,I696015,I696001,);
nand I_40749 (I696332,I610451,I610442);
and I_40750 (I696349,I696332,I610439);
DFFARX1 I_40751 (I696349,I3563,I696015,I696375,);
nor I_40752 (I696383,I696375,I696242);
DFFARX1 I_40753 (I696383,I3563,I696015,I695983,);
nand I_40754 (I696414,I696375,I696284);
nand I_40755 (I695992,I696267,I696414);
not I_40756 (I696445,I696375);
nor I_40757 (I696462,I696445,I696185);
DFFARX1 I_40758 (I696462,I3563,I696015,I696004,);
nor I_40759 (I696493,I610442,I610442);
or I_40760 (I695995,I696242,I696493);
nor I_40761 (I695986,I696375,I696493);
or I_40762 (I695989,I696109,I696493);
DFFARX1 I_40763 (I696493,I3563,I696015,I696007,);
not I_40764 (I696593,I3570);
DFFARX1 I_40765 (I1049470,I3563,I696593,I696619,);
not I_40766 (I696627,I696619);
nand I_40767 (I696644,I1049467,I1049485);
and I_40768 (I696661,I696644,I1049482);
DFFARX1 I_40769 (I696661,I3563,I696593,I696687,);
not I_40770 (I696695,I1049464);
DFFARX1 I_40771 (I1049467,I3563,I696593,I696721,);
not I_40772 (I696729,I696721);
nor I_40773 (I696746,I696729,I696627);
and I_40774 (I696763,I696746,I1049464);
nor I_40775 (I696780,I696729,I696695);
nor I_40776 (I696576,I696687,I696780);
DFFARX1 I_40777 (I1049476,I3563,I696593,I696820,);
nor I_40778 (I696828,I696820,I696687);
not I_40779 (I696845,I696828);
not I_40780 (I696862,I696820);
nor I_40781 (I696879,I696862,I696763);
DFFARX1 I_40782 (I696879,I3563,I696593,I696579,);
nand I_40783 (I696910,I1049479,I1049464);
and I_40784 (I696927,I696910,I1049470);
DFFARX1 I_40785 (I696927,I3563,I696593,I696953,);
nor I_40786 (I696961,I696953,I696820);
DFFARX1 I_40787 (I696961,I3563,I696593,I696561,);
nand I_40788 (I696992,I696953,I696862);
nand I_40789 (I696570,I696845,I696992);
not I_40790 (I697023,I696953);
nor I_40791 (I697040,I697023,I696763);
DFFARX1 I_40792 (I697040,I3563,I696593,I696582,);
nor I_40793 (I697071,I1049473,I1049464);
or I_40794 (I696573,I696820,I697071);
nor I_40795 (I696564,I696953,I697071);
or I_40796 (I696567,I696687,I697071);
DFFARX1 I_40797 (I697071,I3563,I696593,I696585,);
not I_40798 (I697171,I3570);
DFFARX1 I_40799 (I52443,I3563,I697171,I697197,);
not I_40800 (I697205,I697197);
nand I_40801 (I697222,I52440,I52431);
and I_40802 (I697239,I697222,I52431);
DFFARX1 I_40803 (I697239,I3563,I697171,I697265,);
not I_40804 (I697273,I52434);
DFFARX1 I_40805 (I52449,I3563,I697171,I697299,);
not I_40806 (I697307,I697299);
nor I_40807 (I697324,I697307,I697205);
and I_40808 (I697341,I697324,I52434);
nor I_40809 (I697358,I697307,I697273);
nor I_40810 (I697154,I697265,I697358);
DFFARX1 I_40811 (I52434,I3563,I697171,I697398,);
nor I_40812 (I697406,I697398,I697265);
not I_40813 (I697423,I697406);
not I_40814 (I697440,I697398);
nor I_40815 (I697457,I697440,I697341);
DFFARX1 I_40816 (I697457,I3563,I697171,I697157,);
nand I_40817 (I697488,I52452,I52437);
and I_40818 (I697505,I697488,I52455);
DFFARX1 I_40819 (I697505,I3563,I697171,I697531,);
nor I_40820 (I697539,I697531,I697398);
DFFARX1 I_40821 (I697539,I3563,I697171,I697139,);
nand I_40822 (I697570,I697531,I697440);
nand I_40823 (I697148,I697423,I697570);
not I_40824 (I697601,I697531);
nor I_40825 (I697618,I697601,I697341);
DFFARX1 I_40826 (I697618,I3563,I697171,I697160,);
nor I_40827 (I697649,I52446,I52437);
or I_40828 (I697151,I697398,I697649);
nor I_40829 (I697142,I697531,I697649);
or I_40830 (I697145,I697265,I697649);
DFFARX1 I_40831 (I697649,I3563,I697171,I697163,);
not I_40832 (I697749,I3570);
DFFARX1 I_40833 (I122525,I3563,I697749,I697775,);
not I_40834 (I697783,I697775);
nand I_40835 (I697800,I122534,I122543);
and I_40836 (I697817,I697800,I122522);
DFFARX1 I_40837 (I697817,I3563,I697749,I697843,);
not I_40838 (I697851,I122525);
DFFARX1 I_40839 (I122540,I3563,I697749,I697877,);
not I_40840 (I697885,I697877);
nor I_40841 (I697902,I697885,I697783);
and I_40842 (I697919,I697902,I122525);
nor I_40843 (I697936,I697885,I697851);
nor I_40844 (I697732,I697843,I697936);
DFFARX1 I_40845 (I122531,I3563,I697749,I697976,);
nor I_40846 (I697984,I697976,I697843);
not I_40847 (I698001,I697984);
not I_40848 (I698018,I697976);
nor I_40849 (I698035,I698018,I697919);
DFFARX1 I_40850 (I698035,I3563,I697749,I697735,);
nand I_40851 (I698066,I122546,I122522);
and I_40852 (I698083,I698066,I122528);
DFFARX1 I_40853 (I698083,I3563,I697749,I698109,);
nor I_40854 (I698117,I698109,I697976);
DFFARX1 I_40855 (I698117,I3563,I697749,I697717,);
nand I_40856 (I698148,I698109,I698018);
nand I_40857 (I697726,I698001,I698148);
not I_40858 (I698179,I698109);
nor I_40859 (I698196,I698179,I697919);
DFFARX1 I_40860 (I698196,I3563,I697749,I697738,);
nor I_40861 (I698227,I122537,I122522);
or I_40862 (I697729,I697976,I698227);
nor I_40863 (I697720,I698109,I698227);
or I_40864 (I697723,I697843,I698227);
DFFARX1 I_40865 (I698227,I3563,I697749,I697741,);
not I_40866 (I698327,I3570);
DFFARX1 I_40867 (I1144189,I3563,I698327,I698353,);
not I_40868 (I698361,I698353);
nand I_40869 (I698378,I1144171,I1144183);
and I_40870 (I698395,I698378,I1144186);
DFFARX1 I_40871 (I698395,I3563,I698327,I698421,);
not I_40872 (I698429,I1144180);
DFFARX1 I_40873 (I1144177,I3563,I698327,I698455,);
not I_40874 (I698463,I698455);
nor I_40875 (I698480,I698463,I698361);
and I_40876 (I698497,I698480,I1144180);
nor I_40877 (I698514,I698463,I698429);
nor I_40878 (I698310,I698421,I698514);
DFFARX1 I_40879 (I1144195,I3563,I698327,I698554,);
nor I_40880 (I698562,I698554,I698421);
not I_40881 (I698579,I698562);
not I_40882 (I698596,I698554);
nor I_40883 (I698613,I698596,I698497);
DFFARX1 I_40884 (I698613,I3563,I698327,I698313,);
nand I_40885 (I698644,I1144174,I1144174);
and I_40886 (I698661,I698644,I1144171);
DFFARX1 I_40887 (I698661,I3563,I698327,I698687,);
nor I_40888 (I698695,I698687,I698554);
DFFARX1 I_40889 (I698695,I3563,I698327,I698295,);
nand I_40890 (I698726,I698687,I698596);
nand I_40891 (I698304,I698579,I698726);
not I_40892 (I698757,I698687);
nor I_40893 (I698774,I698757,I698497);
DFFARX1 I_40894 (I698774,I3563,I698327,I698316,);
nor I_40895 (I698805,I1144192,I1144174);
or I_40896 (I698307,I698554,I698805);
nor I_40897 (I698298,I698687,I698805);
or I_40898 (I698301,I698421,I698805);
DFFARX1 I_40899 (I698805,I3563,I698327,I698319,);
not I_40900 (I698905,I3570);
DFFARX1 I_40901 (I1173089,I3563,I698905,I698931,);
not I_40902 (I698939,I698931);
nand I_40903 (I698956,I1173071,I1173083);
and I_40904 (I698973,I698956,I1173086);
DFFARX1 I_40905 (I698973,I3563,I698905,I698999,);
not I_40906 (I699007,I1173080);
DFFARX1 I_40907 (I1173077,I3563,I698905,I699033,);
not I_40908 (I699041,I699033);
nor I_40909 (I699058,I699041,I698939);
and I_40910 (I699075,I699058,I1173080);
nor I_40911 (I699092,I699041,I699007);
nor I_40912 (I698888,I698999,I699092);
DFFARX1 I_40913 (I1173095,I3563,I698905,I699132,);
nor I_40914 (I699140,I699132,I698999);
not I_40915 (I699157,I699140);
not I_40916 (I699174,I699132);
nor I_40917 (I699191,I699174,I699075);
DFFARX1 I_40918 (I699191,I3563,I698905,I698891,);
nand I_40919 (I699222,I1173074,I1173074);
and I_40920 (I699239,I699222,I1173071);
DFFARX1 I_40921 (I699239,I3563,I698905,I699265,);
nor I_40922 (I699273,I699265,I699132);
DFFARX1 I_40923 (I699273,I3563,I698905,I698873,);
nand I_40924 (I699304,I699265,I699174);
nand I_40925 (I698882,I699157,I699304);
not I_40926 (I699335,I699265);
nor I_40927 (I699352,I699335,I699075);
DFFARX1 I_40928 (I699352,I3563,I698905,I698894,);
nor I_40929 (I699383,I1173092,I1173074);
or I_40930 (I698885,I699132,I699383);
nor I_40931 (I698876,I699265,I699383);
or I_40932 (I698879,I698999,I699383);
DFFARX1 I_40933 (I699383,I3563,I698905,I698897,);
not I_40934 (I699483,I3570);
DFFARX1 I_40935 (I594255,I3563,I699483,I699509,);
not I_40936 (I699517,I699509);
nand I_40937 (I699534,I594264,I594273);
and I_40938 (I699551,I699534,I594279);
DFFARX1 I_40939 (I699551,I3563,I699483,I699577,);
not I_40940 (I699585,I594276);
DFFARX1 I_40941 (I594261,I3563,I699483,I699611,);
not I_40942 (I699619,I699611);
nor I_40943 (I699636,I699619,I699517);
and I_40944 (I699653,I699636,I594276);
nor I_40945 (I699670,I699619,I699585);
nor I_40946 (I699466,I699577,I699670);
DFFARX1 I_40947 (I594270,I3563,I699483,I699710,);
nor I_40948 (I699718,I699710,I699577);
not I_40949 (I699735,I699718);
not I_40950 (I699752,I699710);
nor I_40951 (I699769,I699752,I699653);
DFFARX1 I_40952 (I699769,I3563,I699483,I699469,);
nand I_40953 (I699800,I594267,I594258);
and I_40954 (I699817,I699800,I594255);
DFFARX1 I_40955 (I699817,I3563,I699483,I699843,);
nor I_40956 (I699851,I699843,I699710);
DFFARX1 I_40957 (I699851,I3563,I699483,I699451,);
nand I_40958 (I699882,I699843,I699752);
nand I_40959 (I699460,I699735,I699882);
not I_40960 (I699913,I699843);
nor I_40961 (I699930,I699913,I699653);
DFFARX1 I_40962 (I699930,I3563,I699483,I699472,);
nor I_40963 (I699961,I594258,I594258);
or I_40964 (I699463,I699710,I699961);
nor I_40965 (I699454,I699843,I699961);
or I_40966 (I699457,I699577,I699961);
DFFARX1 I_40967 (I699961,I3563,I699483,I699475,);
not I_40968 (I700061,I3570);
DFFARX1 I_40969 (I288024,I3563,I700061,I700087,);
not I_40970 (I700095,I700087);
nand I_40971 (I700112,I288027,I288003);
and I_40972 (I700129,I700112,I288000);
DFFARX1 I_40973 (I700129,I3563,I700061,I700155,);
not I_40974 (I700163,I288006);
DFFARX1 I_40975 (I288000,I3563,I700061,I700189,);
not I_40976 (I700197,I700189);
nor I_40977 (I700214,I700197,I700095);
and I_40978 (I700231,I700214,I288006);
nor I_40979 (I700248,I700197,I700163);
nor I_40980 (I700044,I700155,I700248);
DFFARX1 I_40981 (I288009,I3563,I700061,I700288,);
nor I_40982 (I700296,I700288,I700155);
not I_40983 (I700313,I700296);
not I_40984 (I700330,I700288);
nor I_40985 (I700347,I700330,I700231);
DFFARX1 I_40986 (I700347,I3563,I700061,I700047,);
nand I_40987 (I700378,I288012,I288021);
and I_40988 (I700395,I700378,I288018);
DFFARX1 I_40989 (I700395,I3563,I700061,I700421,);
nor I_40990 (I700429,I700421,I700288);
DFFARX1 I_40991 (I700429,I3563,I700061,I700029,);
nand I_40992 (I700460,I700421,I700330);
nand I_40993 (I700038,I700313,I700460);
not I_40994 (I700491,I700421);
nor I_40995 (I700508,I700491,I700231);
DFFARX1 I_40996 (I700508,I3563,I700061,I700050,);
nor I_40997 (I700539,I288015,I288021);
or I_40998 (I700041,I700288,I700539);
nor I_40999 (I700032,I700421,I700539);
or I_41000 (I700035,I700155,I700539);
DFFARX1 I_41001 (I700539,I3563,I700061,I700053,);
not I_41002 (I700639,I3570);
DFFARX1 I_41003 (I563791,I3563,I700639,I700665,);
not I_41004 (I700673,I700665);
nand I_41005 (I700690,I563806,I563791);
and I_41006 (I700707,I700690,I563794);
DFFARX1 I_41007 (I700707,I3563,I700639,I700733,);
not I_41008 (I700741,I563794);
DFFARX1 I_41009 (I563803,I3563,I700639,I700767,);
not I_41010 (I700775,I700767);
nor I_41011 (I700792,I700775,I700673);
and I_41012 (I700809,I700792,I563794);
nor I_41013 (I700826,I700775,I700741);
nor I_41014 (I700622,I700733,I700826);
DFFARX1 I_41015 (I563797,I3563,I700639,I700866,);
nor I_41016 (I700874,I700866,I700733);
not I_41017 (I700891,I700874);
not I_41018 (I700908,I700866);
nor I_41019 (I700925,I700908,I700809);
DFFARX1 I_41020 (I700925,I3563,I700639,I700625,);
nand I_41021 (I700956,I563800,I563809);
and I_41022 (I700973,I700956,I563815);
DFFARX1 I_41023 (I700973,I3563,I700639,I700999,);
nor I_41024 (I701007,I700999,I700866);
DFFARX1 I_41025 (I701007,I3563,I700639,I700607,);
nand I_41026 (I701038,I700999,I700908);
nand I_41027 (I700616,I700891,I701038);
not I_41028 (I701069,I700999);
nor I_41029 (I701086,I701069,I700809);
DFFARX1 I_41030 (I701086,I3563,I700639,I700628,);
nor I_41031 (I701117,I563812,I563809);
or I_41032 (I700619,I700866,I701117);
nor I_41033 (I700610,I700999,I701117);
or I_41034 (I700613,I700733,I701117);
DFFARX1 I_41035 (I701117,I3563,I700639,I700631,);
not I_41036 (I701217,I3570);
DFFARX1 I_41037 (I542966,I3563,I701217,I701243,);
not I_41038 (I701251,I701243);
nand I_41039 (I701268,I542981,I542966);
and I_41040 (I701285,I701268,I542969);
DFFARX1 I_41041 (I701285,I3563,I701217,I701311,);
not I_41042 (I701319,I542969);
DFFARX1 I_41043 (I542978,I3563,I701217,I701345,);
not I_41044 (I701353,I701345);
nor I_41045 (I701370,I701353,I701251);
and I_41046 (I701387,I701370,I542969);
nor I_41047 (I701404,I701353,I701319);
nor I_41048 (I701200,I701311,I701404);
DFFARX1 I_41049 (I542972,I3563,I701217,I701444,);
nor I_41050 (I701452,I701444,I701311);
not I_41051 (I701469,I701452);
not I_41052 (I701486,I701444);
nor I_41053 (I701503,I701486,I701387);
DFFARX1 I_41054 (I701503,I3563,I701217,I701203,);
nand I_41055 (I701534,I542975,I542984);
and I_41056 (I701551,I701534,I542990);
DFFARX1 I_41057 (I701551,I3563,I701217,I701577,);
nor I_41058 (I701585,I701577,I701444);
DFFARX1 I_41059 (I701585,I3563,I701217,I701185,);
nand I_41060 (I701616,I701577,I701486);
nand I_41061 (I701194,I701469,I701616);
not I_41062 (I701647,I701577);
nor I_41063 (I701664,I701647,I701387);
DFFARX1 I_41064 (I701664,I3563,I701217,I701206,);
nor I_41065 (I701695,I542987,I542984);
or I_41066 (I701197,I701444,I701695);
nor I_41067 (I701188,I701577,I701695);
or I_41068 (I701191,I701311,I701695);
DFFARX1 I_41069 (I701695,I3563,I701217,I701209,);
not I_41070 (I701795,I3570);
DFFARX1 I_41071 (I300672,I3563,I701795,I701821,);
not I_41072 (I701829,I701821);
nand I_41073 (I701846,I300675,I300651);
and I_41074 (I701863,I701846,I300648);
DFFARX1 I_41075 (I701863,I3563,I701795,I701889,);
not I_41076 (I701897,I300654);
DFFARX1 I_41077 (I300648,I3563,I701795,I701923,);
not I_41078 (I701931,I701923);
nor I_41079 (I701948,I701931,I701829);
and I_41080 (I701965,I701948,I300654);
nor I_41081 (I701982,I701931,I701897);
nor I_41082 (I701778,I701889,I701982);
DFFARX1 I_41083 (I300657,I3563,I701795,I702022,);
nor I_41084 (I702030,I702022,I701889);
not I_41085 (I702047,I702030);
not I_41086 (I702064,I702022);
nor I_41087 (I702081,I702064,I701965);
DFFARX1 I_41088 (I702081,I3563,I701795,I701781,);
nand I_41089 (I702112,I300660,I300669);
and I_41090 (I702129,I702112,I300666);
DFFARX1 I_41091 (I702129,I3563,I701795,I702155,);
nor I_41092 (I702163,I702155,I702022);
DFFARX1 I_41093 (I702163,I3563,I701795,I701763,);
nand I_41094 (I702194,I702155,I702064);
nand I_41095 (I701772,I702047,I702194);
not I_41096 (I702225,I702155);
nor I_41097 (I702242,I702225,I701965);
DFFARX1 I_41098 (I702242,I3563,I701795,I701784,);
nor I_41099 (I702273,I300663,I300669);
or I_41100 (I701775,I702022,I702273);
nor I_41101 (I701766,I702155,I702273);
or I_41102 (I701769,I701889,I702273);
DFFARX1 I_41103 (I702273,I3563,I701795,I701787,);
not I_41104 (I702373,I3570);
DFFARX1 I_41105 (I1012445,I3563,I702373,I702399,);
not I_41106 (I702407,I702399);
nand I_41107 (I702424,I1012421,I1012436);
and I_41108 (I702441,I702424,I1012448);
DFFARX1 I_41109 (I702441,I3563,I702373,I702467,);
not I_41110 (I702475,I1012433);
DFFARX1 I_41111 (I1012424,I3563,I702373,I702501,);
not I_41112 (I702509,I702501);
nor I_41113 (I702526,I702509,I702407);
and I_41114 (I702543,I702526,I1012433);
nor I_41115 (I702560,I702509,I702475);
nor I_41116 (I702356,I702467,I702560);
DFFARX1 I_41117 (I1012421,I3563,I702373,I702600,);
nor I_41118 (I702608,I702600,I702467);
not I_41119 (I702625,I702608);
not I_41120 (I702642,I702600);
nor I_41121 (I702659,I702642,I702543);
DFFARX1 I_41122 (I702659,I3563,I702373,I702359,);
nand I_41123 (I702690,I1012439,I1012430);
and I_41124 (I702707,I702690,I1012442);
DFFARX1 I_41125 (I702707,I3563,I702373,I702733,);
nor I_41126 (I702741,I702733,I702600);
DFFARX1 I_41127 (I702741,I3563,I702373,I702341,);
nand I_41128 (I702772,I702733,I702642);
nand I_41129 (I702350,I702625,I702772);
not I_41130 (I702803,I702733);
nor I_41131 (I702820,I702803,I702543);
DFFARX1 I_41132 (I702820,I3563,I702373,I702362,);
nor I_41133 (I702851,I1012427,I1012430);
or I_41134 (I702353,I702600,I702851);
nor I_41135 (I702344,I702733,I702851);
or I_41136 (I702347,I702467,I702851);
DFFARX1 I_41137 (I702851,I3563,I702373,I702365,);
not I_41138 (I702951,I3570);
DFFARX1 I_41139 (I811598,I3563,I702951,I702977,);
not I_41140 (I702985,I702977);
nand I_41141 (I703002,I811586,I811604);
and I_41142 (I703019,I703002,I811601);
DFFARX1 I_41143 (I703019,I3563,I702951,I703045,);
not I_41144 (I703053,I811592);
DFFARX1 I_41145 (I811589,I3563,I702951,I703079,);
not I_41146 (I703087,I703079);
nor I_41147 (I703104,I703087,I702985);
and I_41148 (I703121,I703104,I811592);
nor I_41149 (I703138,I703087,I703053);
nor I_41150 (I702934,I703045,I703138);
DFFARX1 I_41151 (I811583,I3563,I702951,I703178,);
nor I_41152 (I703186,I703178,I703045);
not I_41153 (I703203,I703186);
not I_41154 (I703220,I703178);
nor I_41155 (I703237,I703220,I703121);
DFFARX1 I_41156 (I703237,I3563,I702951,I702937,);
nand I_41157 (I703268,I811583,I811586);
and I_41158 (I703285,I703268,I811589);
DFFARX1 I_41159 (I703285,I3563,I702951,I703311,);
nor I_41160 (I703319,I703311,I703178);
DFFARX1 I_41161 (I703319,I3563,I702951,I702919,);
nand I_41162 (I703350,I703311,I703220);
nand I_41163 (I702928,I703203,I703350);
not I_41164 (I703381,I703311);
nor I_41165 (I703398,I703381,I703121);
DFFARX1 I_41166 (I703398,I3563,I702951,I702940,);
nor I_41167 (I703429,I811595,I811586);
or I_41168 (I702931,I703178,I703429);
nor I_41169 (I702922,I703311,I703429);
or I_41170 (I702925,I703045,I703429);
DFFARX1 I_41171 (I703429,I3563,I702951,I702943,);
not I_41172 (I703529,I3570);
DFFARX1 I_41173 (I991773,I3563,I703529,I703555,);
not I_41174 (I703563,I703555);
nand I_41175 (I703580,I991749,I991764);
and I_41176 (I703597,I703580,I991776);
DFFARX1 I_41177 (I703597,I3563,I703529,I703623,);
not I_41178 (I703631,I991761);
DFFARX1 I_41179 (I991752,I3563,I703529,I703657,);
not I_41180 (I703665,I703657);
nor I_41181 (I703682,I703665,I703563);
and I_41182 (I703699,I703682,I991761);
nor I_41183 (I703716,I703665,I703631);
nor I_41184 (I703512,I703623,I703716);
DFFARX1 I_41185 (I991749,I3563,I703529,I703756,);
nor I_41186 (I703764,I703756,I703623);
not I_41187 (I703781,I703764);
not I_41188 (I703798,I703756);
nor I_41189 (I703815,I703798,I703699);
DFFARX1 I_41190 (I703815,I3563,I703529,I703515,);
nand I_41191 (I703846,I991767,I991758);
and I_41192 (I703863,I703846,I991770);
DFFARX1 I_41193 (I703863,I3563,I703529,I703889,);
nor I_41194 (I703897,I703889,I703756);
DFFARX1 I_41195 (I703897,I3563,I703529,I703497,);
nand I_41196 (I703928,I703889,I703798);
nand I_41197 (I703506,I703781,I703928);
not I_41198 (I703959,I703889);
nor I_41199 (I703976,I703959,I703699);
DFFARX1 I_41200 (I703976,I3563,I703529,I703518,);
nor I_41201 (I704007,I991755,I991758);
or I_41202 (I703509,I703756,I704007);
nor I_41203 (I703500,I703889,I704007);
or I_41204 (I703503,I703623,I704007);
DFFARX1 I_41205 (I704007,I3563,I703529,I703521,);
not I_41206 (I704107,I3570);
DFFARX1 I_41207 (I1141299,I3563,I704107,I704133,);
not I_41208 (I704141,I704133);
nand I_41209 (I704158,I1141281,I1141293);
and I_41210 (I704175,I704158,I1141296);
DFFARX1 I_41211 (I704175,I3563,I704107,I704201,);
not I_41212 (I704209,I1141290);
DFFARX1 I_41213 (I1141287,I3563,I704107,I704235,);
not I_41214 (I704243,I704235);
nor I_41215 (I704260,I704243,I704141);
and I_41216 (I704277,I704260,I1141290);
nor I_41217 (I704294,I704243,I704209);
nor I_41218 (I704090,I704201,I704294);
DFFARX1 I_41219 (I1141305,I3563,I704107,I704334,);
nor I_41220 (I704342,I704334,I704201);
not I_41221 (I704359,I704342);
not I_41222 (I704376,I704334);
nor I_41223 (I704393,I704376,I704277);
DFFARX1 I_41224 (I704393,I3563,I704107,I704093,);
nand I_41225 (I704424,I1141284,I1141284);
and I_41226 (I704441,I704424,I1141281);
DFFARX1 I_41227 (I704441,I3563,I704107,I704467,);
nor I_41228 (I704475,I704467,I704334);
DFFARX1 I_41229 (I704475,I3563,I704107,I704075,);
nand I_41230 (I704506,I704467,I704376);
nand I_41231 (I704084,I704359,I704506);
not I_41232 (I704537,I704467);
nor I_41233 (I704554,I704537,I704277);
DFFARX1 I_41234 (I704554,I3563,I704107,I704096,);
nor I_41235 (I704585,I1141302,I1141284);
or I_41236 (I704087,I704334,I704585);
nor I_41237 (I704078,I704467,I704585);
or I_41238 (I704081,I704201,I704585);
DFFARX1 I_41239 (I704585,I3563,I704107,I704099,);
not I_41240 (I704685,I3570);
DFFARX1 I_41241 (I1290643,I3563,I704685,I704711,);
not I_41242 (I704719,I704711);
nand I_41243 (I704736,I1290667,I1290649);
and I_41244 (I704753,I704736,I1290655);
DFFARX1 I_41245 (I704753,I3563,I704685,I704779,);
not I_41246 (I704787,I1290661);
DFFARX1 I_41247 (I1290646,I3563,I704685,I704813,);
not I_41248 (I704821,I704813);
nor I_41249 (I704838,I704821,I704719);
and I_41250 (I704855,I704838,I1290661);
nor I_41251 (I704872,I704821,I704787);
nor I_41252 (I704668,I704779,I704872);
DFFARX1 I_41253 (I1290658,I3563,I704685,I704912,);
nor I_41254 (I704920,I704912,I704779);
not I_41255 (I704937,I704920);
not I_41256 (I704954,I704912);
nor I_41257 (I704971,I704954,I704855);
DFFARX1 I_41258 (I704971,I3563,I704685,I704671,);
nand I_41259 (I705002,I1290664,I1290652);
and I_41260 (I705019,I705002,I1290646);
DFFARX1 I_41261 (I705019,I3563,I704685,I705045,);
nor I_41262 (I705053,I705045,I704912);
DFFARX1 I_41263 (I705053,I3563,I704685,I704653,);
nand I_41264 (I705084,I705045,I704954);
nand I_41265 (I704662,I704937,I705084);
not I_41266 (I705115,I705045);
nor I_41267 (I705132,I705115,I704855);
DFFARX1 I_41268 (I705132,I3563,I704685,I704674,);
nor I_41269 (I705163,I1290643,I1290652);
or I_41270 (I704665,I704912,I705163);
nor I_41271 (I704656,I705045,I705163);
or I_41272 (I704659,I704779,I705163);
DFFARX1 I_41273 (I705163,I3563,I704685,I704677,);
not I_41274 (I705263,I3570);
DFFARX1 I_41275 (I827408,I3563,I705263,I705289,);
not I_41276 (I705297,I705289);
nand I_41277 (I705314,I827396,I827414);
and I_41278 (I705331,I705314,I827411);
DFFARX1 I_41279 (I705331,I3563,I705263,I705357,);
not I_41280 (I705365,I827402);
DFFARX1 I_41281 (I827399,I3563,I705263,I705391,);
not I_41282 (I705399,I705391);
nor I_41283 (I705416,I705399,I705297);
and I_41284 (I705433,I705416,I827402);
nor I_41285 (I705450,I705399,I705365);
nor I_41286 (I705246,I705357,I705450);
DFFARX1 I_41287 (I827393,I3563,I705263,I705490,);
nor I_41288 (I705498,I705490,I705357);
not I_41289 (I705515,I705498);
not I_41290 (I705532,I705490);
nor I_41291 (I705549,I705532,I705433);
DFFARX1 I_41292 (I705549,I3563,I705263,I705249,);
nand I_41293 (I705580,I827393,I827396);
and I_41294 (I705597,I705580,I827399);
DFFARX1 I_41295 (I705597,I3563,I705263,I705623,);
nor I_41296 (I705631,I705623,I705490);
DFFARX1 I_41297 (I705631,I3563,I705263,I705231,);
nand I_41298 (I705662,I705623,I705532);
nand I_41299 (I705240,I705515,I705662);
not I_41300 (I705693,I705623);
nor I_41301 (I705710,I705693,I705433);
DFFARX1 I_41302 (I705710,I3563,I705263,I705252,);
nor I_41303 (I705741,I827405,I827396);
or I_41304 (I705243,I705490,I705741);
nor I_41305 (I705234,I705623,I705741);
or I_41306 (I705237,I705357,I705741);
DFFARX1 I_41307 (I705741,I3563,I705263,I705255,);
not I_41308 (I705841,I3570);
DFFARX1 I_41309 (I242253,I3563,I705841,I705867,);
not I_41310 (I705875,I705867);
nand I_41311 (I705892,I242256,I242277);
and I_41312 (I705909,I705892,I242265);
DFFARX1 I_41313 (I705909,I3563,I705841,I705935,);
not I_41314 (I705943,I242262);
DFFARX1 I_41315 (I242253,I3563,I705841,I705969,);
not I_41316 (I705977,I705969);
nor I_41317 (I705994,I705977,I705875);
and I_41318 (I706011,I705994,I242262);
nor I_41319 (I706028,I705977,I705943);
nor I_41320 (I705824,I705935,I706028);
DFFARX1 I_41321 (I242271,I3563,I705841,I706068,);
nor I_41322 (I706076,I706068,I705935);
not I_41323 (I706093,I706076);
not I_41324 (I706110,I706068);
nor I_41325 (I706127,I706110,I706011);
DFFARX1 I_41326 (I706127,I3563,I705841,I705827,);
nand I_41327 (I706158,I242256,I242259);
and I_41328 (I706175,I706158,I242268);
DFFARX1 I_41329 (I706175,I3563,I705841,I706201,);
nor I_41330 (I706209,I706201,I706068);
DFFARX1 I_41331 (I706209,I3563,I705841,I705809,);
nand I_41332 (I706240,I706201,I706110);
nand I_41333 (I705818,I706093,I706240);
not I_41334 (I706271,I706201);
nor I_41335 (I706288,I706271,I706011);
DFFARX1 I_41336 (I706288,I3563,I705841,I705830,);
nor I_41337 (I706319,I242274,I242259);
or I_41338 (I705821,I706068,I706319);
nor I_41339 (I705812,I706201,I706319);
or I_41340 (I705815,I705935,I706319);
DFFARX1 I_41341 (I706319,I3563,I705841,I705833,);
not I_41342 (I706419,I3570);
DFFARX1 I_41343 (I1207191,I3563,I706419,I706445,);
not I_41344 (I706453,I706445);
nand I_41345 (I706470,I1207173,I1207185);
and I_41346 (I706487,I706470,I1207188);
DFFARX1 I_41347 (I706487,I3563,I706419,I706513,);
not I_41348 (I706521,I1207182);
DFFARX1 I_41349 (I1207179,I3563,I706419,I706547,);
not I_41350 (I706555,I706547);
nor I_41351 (I706572,I706555,I706453);
and I_41352 (I706589,I706572,I1207182);
nor I_41353 (I706606,I706555,I706521);
nor I_41354 (I706402,I706513,I706606);
DFFARX1 I_41355 (I1207197,I3563,I706419,I706646,);
nor I_41356 (I706654,I706646,I706513);
not I_41357 (I706671,I706654);
not I_41358 (I706688,I706646);
nor I_41359 (I706705,I706688,I706589);
DFFARX1 I_41360 (I706705,I3563,I706419,I706405,);
nand I_41361 (I706736,I1207176,I1207176);
and I_41362 (I706753,I706736,I1207173);
DFFARX1 I_41363 (I706753,I3563,I706419,I706779,);
nor I_41364 (I706787,I706779,I706646);
DFFARX1 I_41365 (I706787,I3563,I706419,I706387,);
nand I_41366 (I706818,I706779,I706688);
nand I_41367 (I706396,I706671,I706818);
not I_41368 (I706849,I706779);
nor I_41369 (I706866,I706849,I706589);
DFFARX1 I_41370 (I706866,I3563,I706419,I706408,);
nor I_41371 (I706897,I1207194,I1207176);
or I_41372 (I706399,I706646,I706897);
nor I_41373 (I706390,I706779,I706897);
or I_41374 (I706393,I706513,I706897);
DFFARX1 I_41375 (I706897,I3563,I706419,I706411,);
not I_41376 (I706997,I3570);
DFFARX1 I_41377 (I332292,I3563,I706997,I707023,);
not I_41378 (I707031,I707023);
nand I_41379 (I707048,I332295,I332271);
and I_41380 (I707065,I707048,I332268);
DFFARX1 I_41381 (I707065,I3563,I706997,I707091,);
not I_41382 (I707099,I332274);
DFFARX1 I_41383 (I332268,I3563,I706997,I707125,);
not I_41384 (I707133,I707125);
nor I_41385 (I707150,I707133,I707031);
and I_41386 (I707167,I707150,I332274);
nor I_41387 (I707184,I707133,I707099);
nor I_41388 (I706980,I707091,I707184);
DFFARX1 I_41389 (I332277,I3563,I706997,I707224,);
nor I_41390 (I707232,I707224,I707091);
not I_41391 (I707249,I707232);
not I_41392 (I707266,I707224);
nor I_41393 (I707283,I707266,I707167);
DFFARX1 I_41394 (I707283,I3563,I706997,I706983,);
nand I_41395 (I707314,I332280,I332289);
and I_41396 (I707331,I707314,I332286);
DFFARX1 I_41397 (I707331,I3563,I706997,I707357,);
nor I_41398 (I707365,I707357,I707224);
DFFARX1 I_41399 (I707365,I3563,I706997,I706965,);
nand I_41400 (I707396,I707357,I707266);
nand I_41401 (I706974,I707249,I707396);
not I_41402 (I707427,I707357);
nor I_41403 (I707444,I707427,I707167);
DFFARX1 I_41404 (I707444,I3563,I706997,I706986,);
nor I_41405 (I707475,I332283,I332289);
or I_41406 (I706977,I707224,I707475);
nor I_41407 (I706968,I707357,I707475);
or I_41408 (I706971,I707091,I707475);
DFFARX1 I_41409 (I707475,I3563,I706997,I706989,);
not I_41410 (I707575,I3570);
DFFARX1 I_41411 (I1378560,I3563,I707575,I707601,);
not I_41412 (I707609,I707601);
nand I_41413 (I707626,I1378545,I1378533);
and I_41414 (I707643,I707626,I1378548);
DFFARX1 I_41415 (I707643,I3563,I707575,I707669,);
not I_41416 (I707677,I1378533);
DFFARX1 I_41417 (I1378551,I3563,I707575,I707703,);
not I_41418 (I707711,I707703);
nor I_41419 (I707728,I707711,I707609);
and I_41420 (I707745,I707728,I1378533);
nor I_41421 (I707762,I707711,I707677);
nor I_41422 (I707558,I707669,I707762);
DFFARX1 I_41423 (I1378539,I3563,I707575,I707802,);
nor I_41424 (I707810,I707802,I707669);
not I_41425 (I707827,I707810);
not I_41426 (I707844,I707802);
nor I_41427 (I707861,I707844,I707745);
DFFARX1 I_41428 (I707861,I3563,I707575,I707561,);
nand I_41429 (I707892,I1378536,I1378542);
and I_41430 (I707909,I707892,I1378557);
DFFARX1 I_41431 (I707909,I3563,I707575,I707935,);
nor I_41432 (I707943,I707935,I707802);
DFFARX1 I_41433 (I707943,I3563,I707575,I707543,);
nand I_41434 (I707974,I707935,I707844);
nand I_41435 (I707552,I707827,I707974);
not I_41436 (I708005,I707935);
nor I_41437 (I708022,I708005,I707745);
DFFARX1 I_41438 (I708022,I3563,I707575,I707564,);
nor I_41439 (I708053,I1378554,I1378542);
or I_41440 (I707555,I707802,I708053);
nor I_41441 (I707546,I707935,I708053);
or I_41442 (I707549,I707669,I708053);
DFFARX1 I_41443 (I708053,I3563,I707575,I707567,);
not I_41444 (I708153,I3570);
DFFARX1 I_41445 (I973685,I3563,I708153,I708179,);
not I_41446 (I708187,I708179);
nand I_41447 (I708204,I973661,I973676);
and I_41448 (I708221,I708204,I973688);
DFFARX1 I_41449 (I708221,I3563,I708153,I708247,);
not I_41450 (I708255,I973673);
DFFARX1 I_41451 (I973664,I3563,I708153,I708281,);
not I_41452 (I708289,I708281);
nor I_41453 (I708306,I708289,I708187);
and I_41454 (I708323,I708306,I973673);
nor I_41455 (I708340,I708289,I708255);
nor I_41456 (I708136,I708247,I708340);
DFFARX1 I_41457 (I973661,I3563,I708153,I708380,);
nor I_41458 (I708388,I708380,I708247);
not I_41459 (I708405,I708388);
not I_41460 (I708422,I708380);
nor I_41461 (I708439,I708422,I708323);
DFFARX1 I_41462 (I708439,I3563,I708153,I708139,);
nand I_41463 (I708470,I973679,I973670);
and I_41464 (I708487,I708470,I973682);
DFFARX1 I_41465 (I708487,I3563,I708153,I708513,);
nor I_41466 (I708521,I708513,I708380);
DFFARX1 I_41467 (I708521,I3563,I708153,I708121,);
nand I_41468 (I708552,I708513,I708422);
nand I_41469 (I708130,I708405,I708552);
not I_41470 (I708583,I708513);
nor I_41471 (I708600,I708583,I708323);
DFFARX1 I_41472 (I708600,I3563,I708153,I708142,);
nor I_41473 (I708631,I973667,I973670);
or I_41474 (I708133,I708380,I708631);
nor I_41475 (I708124,I708513,I708631);
or I_41476 (I708127,I708247,I708631);
DFFARX1 I_41477 (I708631,I3563,I708153,I708145,);
not I_41478 (I708731,I3570);
DFFARX1 I_41479 (I274383,I3563,I708731,I708757,);
not I_41480 (I708765,I708757);
nand I_41481 (I708782,I274386,I274407);
and I_41482 (I708799,I708782,I274395);
DFFARX1 I_41483 (I708799,I3563,I708731,I708825,);
not I_41484 (I708833,I274392);
DFFARX1 I_41485 (I274383,I3563,I708731,I708859,);
not I_41486 (I708867,I708859);
nor I_41487 (I708884,I708867,I708765);
and I_41488 (I708901,I708884,I274392);
nor I_41489 (I708918,I708867,I708833);
nor I_41490 (I708714,I708825,I708918);
DFFARX1 I_41491 (I274401,I3563,I708731,I708958,);
nor I_41492 (I708966,I708958,I708825);
not I_41493 (I708983,I708966);
not I_41494 (I709000,I708958);
nor I_41495 (I709017,I709000,I708901);
DFFARX1 I_41496 (I709017,I3563,I708731,I708717,);
nand I_41497 (I709048,I274386,I274389);
and I_41498 (I709065,I709048,I274398);
DFFARX1 I_41499 (I709065,I3563,I708731,I709091,);
nor I_41500 (I709099,I709091,I708958);
DFFARX1 I_41501 (I709099,I3563,I708731,I708699,);
nand I_41502 (I709130,I709091,I709000);
nand I_41503 (I708708,I708983,I709130);
not I_41504 (I709161,I709091);
nor I_41505 (I709178,I709161,I708901);
DFFARX1 I_41506 (I709178,I3563,I708731,I708720,);
nor I_41507 (I709209,I274404,I274389);
or I_41508 (I708711,I708958,I709209);
nor I_41509 (I708702,I709091,I709209);
or I_41510 (I708705,I708825,I709209);
DFFARX1 I_41511 (I709209,I3563,I708731,I708723,);
not I_41512 (I709309,I3570);
DFFARX1 I_41513 (I816868,I3563,I709309,I709335,);
not I_41514 (I709343,I709335);
nand I_41515 (I709360,I816856,I816874);
and I_41516 (I709377,I709360,I816871);
DFFARX1 I_41517 (I709377,I3563,I709309,I709403,);
not I_41518 (I709411,I816862);
DFFARX1 I_41519 (I816859,I3563,I709309,I709437,);
not I_41520 (I709445,I709437);
nor I_41521 (I709462,I709445,I709343);
and I_41522 (I709479,I709462,I816862);
nor I_41523 (I709496,I709445,I709411);
nor I_41524 (I709292,I709403,I709496);
DFFARX1 I_41525 (I816853,I3563,I709309,I709536,);
nor I_41526 (I709544,I709536,I709403);
not I_41527 (I709561,I709544);
not I_41528 (I709578,I709536);
nor I_41529 (I709595,I709578,I709479);
DFFARX1 I_41530 (I709595,I3563,I709309,I709295,);
nand I_41531 (I709626,I816853,I816856);
and I_41532 (I709643,I709626,I816859);
DFFARX1 I_41533 (I709643,I3563,I709309,I709669,);
nor I_41534 (I709677,I709669,I709536);
DFFARX1 I_41535 (I709677,I3563,I709309,I709277,);
nand I_41536 (I709708,I709669,I709578);
nand I_41537 (I709286,I709561,I709708);
not I_41538 (I709739,I709669);
nor I_41539 (I709756,I709739,I709479);
DFFARX1 I_41540 (I709756,I3563,I709309,I709298,);
nor I_41541 (I709787,I816865,I816856);
or I_41542 (I709289,I709536,I709787);
nor I_41543 (I709280,I709669,I709787);
or I_41544 (I709283,I709403,I709787);
DFFARX1 I_41545 (I709787,I3563,I709309,I709301,);
not I_41546 (I709887,I3570);
DFFARX1 I_41547 (I1374395,I3563,I709887,I709913,);
not I_41548 (I709921,I709913);
nand I_41549 (I709938,I1374380,I1374368);
and I_41550 (I709955,I709938,I1374383);
DFFARX1 I_41551 (I709955,I3563,I709887,I709981,);
not I_41552 (I709989,I1374368);
DFFARX1 I_41553 (I1374386,I3563,I709887,I710015,);
not I_41554 (I710023,I710015);
nor I_41555 (I710040,I710023,I709921);
and I_41556 (I710057,I710040,I1374368);
nor I_41557 (I710074,I710023,I709989);
nor I_41558 (I709870,I709981,I710074);
DFFARX1 I_41559 (I1374374,I3563,I709887,I710114,);
nor I_41560 (I710122,I710114,I709981);
not I_41561 (I710139,I710122);
not I_41562 (I710156,I710114);
nor I_41563 (I710173,I710156,I710057);
DFFARX1 I_41564 (I710173,I3563,I709887,I709873,);
nand I_41565 (I710204,I1374371,I1374377);
and I_41566 (I710221,I710204,I1374392);
DFFARX1 I_41567 (I710221,I3563,I709887,I710247,);
nor I_41568 (I710255,I710247,I710114);
DFFARX1 I_41569 (I710255,I3563,I709887,I709855,);
nand I_41570 (I710286,I710247,I710156);
nand I_41571 (I709864,I710139,I710286);
not I_41572 (I710317,I710247);
nor I_41573 (I710334,I710317,I710057);
DFFARX1 I_41574 (I710334,I3563,I709887,I709876,);
nor I_41575 (I710365,I1374389,I1374377);
or I_41576 (I709867,I710114,I710365);
nor I_41577 (I709858,I710247,I710365);
or I_41578 (I709861,I709981,I710365);
DFFARX1 I_41579 (I710365,I3563,I709887,I709879,);
not I_41580 (I710465,I3570);
DFFARX1 I_41581 (I1026011,I3563,I710465,I710491,);
not I_41582 (I710499,I710491);
nand I_41583 (I710516,I1025987,I1026002);
and I_41584 (I710533,I710516,I1026014);
DFFARX1 I_41585 (I710533,I3563,I710465,I710559,);
not I_41586 (I710567,I1025999);
DFFARX1 I_41587 (I1025990,I3563,I710465,I710593,);
not I_41588 (I710601,I710593);
nor I_41589 (I710618,I710601,I710499);
and I_41590 (I710635,I710618,I1025999);
nor I_41591 (I710652,I710601,I710567);
nor I_41592 (I710448,I710559,I710652);
DFFARX1 I_41593 (I1025987,I3563,I710465,I710692,);
nor I_41594 (I710700,I710692,I710559);
not I_41595 (I710717,I710700);
not I_41596 (I710734,I710692);
nor I_41597 (I710751,I710734,I710635);
DFFARX1 I_41598 (I710751,I3563,I710465,I710451,);
nand I_41599 (I710782,I1026005,I1025996);
and I_41600 (I710799,I710782,I1026008);
DFFARX1 I_41601 (I710799,I3563,I710465,I710825,);
nor I_41602 (I710833,I710825,I710692);
DFFARX1 I_41603 (I710833,I3563,I710465,I710433,);
nand I_41604 (I710864,I710825,I710734);
nand I_41605 (I710442,I710717,I710864);
not I_41606 (I710895,I710825);
nor I_41607 (I710912,I710895,I710635);
DFFARX1 I_41608 (I710912,I3563,I710465,I710454,);
nor I_41609 (I710943,I1025993,I1025996);
or I_41610 (I710445,I710692,I710943);
nor I_41611 (I710436,I710825,I710943);
or I_41612 (I710439,I710559,I710943);
DFFARX1 I_41613 (I710943,I3563,I710465,I710457,);
not I_41614 (I711043,I3570);
DFFARX1 I_41615 (I142024,I3563,I711043,I711069,);
not I_41616 (I711077,I711069);
nand I_41617 (I711094,I142033,I142042);
and I_41618 (I711111,I711094,I142021);
DFFARX1 I_41619 (I711111,I3563,I711043,I711137,);
not I_41620 (I711145,I142024);
DFFARX1 I_41621 (I142039,I3563,I711043,I711171,);
not I_41622 (I711179,I711171);
nor I_41623 (I711196,I711179,I711077);
and I_41624 (I711213,I711196,I142024);
nor I_41625 (I711230,I711179,I711145);
nor I_41626 (I711026,I711137,I711230);
DFFARX1 I_41627 (I142030,I3563,I711043,I711270,);
nor I_41628 (I711278,I711270,I711137);
not I_41629 (I711295,I711278);
not I_41630 (I711312,I711270);
nor I_41631 (I711329,I711312,I711213);
DFFARX1 I_41632 (I711329,I3563,I711043,I711029,);
nand I_41633 (I711360,I142045,I142021);
and I_41634 (I711377,I711360,I142027);
DFFARX1 I_41635 (I711377,I3563,I711043,I711403,);
nor I_41636 (I711411,I711403,I711270);
DFFARX1 I_41637 (I711411,I3563,I711043,I711011,);
nand I_41638 (I711442,I711403,I711312);
nand I_41639 (I711020,I711295,I711442);
not I_41640 (I711473,I711403);
nor I_41641 (I711490,I711473,I711213);
DFFARX1 I_41642 (I711490,I3563,I711043,I711032,);
nor I_41643 (I711521,I142036,I142021);
or I_41644 (I711023,I711270,I711521);
nor I_41645 (I711014,I711403,I711521);
or I_41646 (I711017,I711137,I711521);
DFFARX1 I_41647 (I711521,I3563,I711043,I711035,);
not I_41648 (I711621,I3570);
DFFARX1 I_41649 (I958181,I3563,I711621,I711647,);
not I_41650 (I711655,I711647);
nand I_41651 (I711672,I958157,I958172);
and I_41652 (I711689,I711672,I958184);
DFFARX1 I_41653 (I711689,I3563,I711621,I711715,);
not I_41654 (I711723,I958169);
DFFARX1 I_41655 (I958160,I3563,I711621,I711749,);
not I_41656 (I711757,I711749);
nor I_41657 (I711774,I711757,I711655);
and I_41658 (I711791,I711774,I958169);
nor I_41659 (I711808,I711757,I711723);
nor I_41660 (I711604,I711715,I711808);
DFFARX1 I_41661 (I958157,I3563,I711621,I711848,);
nor I_41662 (I711856,I711848,I711715);
not I_41663 (I711873,I711856);
not I_41664 (I711890,I711848);
nor I_41665 (I711907,I711890,I711791);
DFFARX1 I_41666 (I711907,I3563,I711621,I711607,);
nand I_41667 (I711938,I958175,I958166);
and I_41668 (I711955,I711938,I958178);
DFFARX1 I_41669 (I711955,I3563,I711621,I711981,);
nor I_41670 (I711989,I711981,I711848);
DFFARX1 I_41671 (I711989,I3563,I711621,I711589,);
nand I_41672 (I712020,I711981,I711890);
nand I_41673 (I711598,I711873,I712020);
not I_41674 (I712051,I711981);
nor I_41675 (I712068,I712051,I711791);
DFFARX1 I_41676 (I712068,I3563,I711621,I711610,);
nor I_41677 (I712099,I958163,I958166);
or I_41678 (I711601,I711848,I712099);
nor I_41679 (I711592,I711981,I712099);
or I_41680 (I711595,I711715,I712099);
DFFARX1 I_41681 (I712099,I3563,I711621,I711613,);
not I_41682 (I712199,I3570);
DFFARX1 I_41683 (I433291,I3563,I712199,I712225,);
not I_41684 (I712233,I712225);
nand I_41685 (I712250,I433282,I433300);
and I_41686 (I712267,I712250,I433303);
DFFARX1 I_41687 (I712267,I3563,I712199,I712293,);
not I_41688 (I712301,I433297);
DFFARX1 I_41689 (I433285,I3563,I712199,I712327,);
not I_41690 (I712335,I712327);
nor I_41691 (I712352,I712335,I712233);
and I_41692 (I712369,I712352,I433297);
nor I_41693 (I712386,I712335,I712301);
nor I_41694 (I712182,I712293,I712386);
DFFARX1 I_41695 (I433294,I3563,I712199,I712426,);
nor I_41696 (I712434,I712426,I712293);
not I_41697 (I712451,I712434);
not I_41698 (I712468,I712426);
nor I_41699 (I712485,I712468,I712369);
DFFARX1 I_41700 (I712485,I3563,I712199,I712185,);
nand I_41701 (I712516,I433309,I433306);
and I_41702 (I712533,I712516,I433288);
DFFARX1 I_41703 (I712533,I3563,I712199,I712559,);
nor I_41704 (I712567,I712559,I712426);
DFFARX1 I_41705 (I712567,I3563,I712199,I712167,);
nand I_41706 (I712598,I712559,I712468);
nand I_41707 (I712176,I712451,I712598);
not I_41708 (I712629,I712559);
nor I_41709 (I712646,I712629,I712369);
DFFARX1 I_41710 (I712646,I3563,I712199,I712188,);
nor I_41711 (I712677,I433282,I433306);
or I_41712 (I712179,I712426,I712677);
nor I_41713 (I712170,I712559,I712677);
or I_41714 (I712173,I712293,I712677);
DFFARX1 I_41715 (I712677,I3563,I712199,I712191,);
not I_41716 (I712777,I3570);
DFFARX1 I_41717 (I1058446,I3563,I712777,I712803,);
not I_41718 (I712811,I712803);
nand I_41719 (I712828,I1058443,I1058461);
and I_41720 (I712845,I712828,I1058458);
DFFARX1 I_41721 (I712845,I3563,I712777,I712871,);
not I_41722 (I712879,I1058440);
DFFARX1 I_41723 (I1058443,I3563,I712777,I712905,);
not I_41724 (I712913,I712905);
nor I_41725 (I712930,I712913,I712811);
and I_41726 (I712947,I712930,I1058440);
nor I_41727 (I712964,I712913,I712879);
nor I_41728 (I712760,I712871,I712964);
DFFARX1 I_41729 (I1058452,I3563,I712777,I713004,);
nor I_41730 (I713012,I713004,I712871);
not I_41731 (I713029,I713012);
not I_41732 (I713046,I713004);
nor I_41733 (I713063,I713046,I712947);
DFFARX1 I_41734 (I713063,I3563,I712777,I712763,);
nand I_41735 (I713094,I1058455,I1058440);
and I_41736 (I713111,I713094,I1058446);
DFFARX1 I_41737 (I713111,I3563,I712777,I713137,);
nor I_41738 (I713145,I713137,I713004);
DFFARX1 I_41739 (I713145,I3563,I712777,I712745,);
nand I_41740 (I713176,I713137,I713046);
nand I_41741 (I712754,I713029,I713176);
not I_41742 (I713207,I713137);
nor I_41743 (I713224,I713207,I712947);
DFFARX1 I_41744 (I713224,I3563,I712777,I712766,);
nor I_41745 (I713255,I1058449,I1058440);
or I_41746 (I712757,I713004,I713255);
nor I_41747 (I712748,I713137,I713255);
or I_41748 (I712751,I712871,I713255);
DFFARX1 I_41749 (I713255,I3563,I712777,I712769,);
not I_41750 (I713355,I3570);
DFFARX1 I_41751 (I1074154,I3563,I713355,I713381,);
not I_41752 (I713389,I713381);
nand I_41753 (I713406,I1074151,I1074169);
and I_41754 (I713423,I713406,I1074166);
DFFARX1 I_41755 (I713423,I3563,I713355,I713449,);
not I_41756 (I713457,I1074148);
DFFARX1 I_41757 (I1074151,I3563,I713355,I713483,);
not I_41758 (I713491,I713483);
nor I_41759 (I713508,I713491,I713389);
and I_41760 (I713525,I713508,I1074148);
nor I_41761 (I713542,I713491,I713457);
nor I_41762 (I713338,I713449,I713542);
DFFARX1 I_41763 (I1074160,I3563,I713355,I713582,);
nor I_41764 (I713590,I713582,I713449);
not I_41765 (I713607,I713590);
not I_41766 (I713624,I713582);
nor I_41767 (I713641,I713624,I713525);
DFFARX1 I_41768 (I713641,I3563,I713355,I713341,);
nand I_41769 (I713672,I1074163,I1074148);
and I_41770 (I713689,I713672,I1074154);
DFFARX1 I_41771 (I713689,I3563,I713355,I713715,);
nor I_41772 (I713723,I713715,I713582);
DFFARX1 I_41773 (I713723,I3563,I713355,I713323,);
nand I_41774 (I713754,I713715,I713624);
nand I_41775 (I713332,I713607,I713754);
not I_41776 (I713785,I713715);
nor I_41777 (I713802,I713785,I713525);
DFFARX1 I_41778 (I713802,I3563,I713355,I713344,);
nor I_41779 (I713833,I1074157,I1074148);
or I_41780 (I713335,I713582,I713833);
nor I_41781 (I713326,I713715,I713833);
or I_41782 (I713329,I713449,I713833);
DFFARX1 I_41783 (I713833,I3563,I713355,I713347,);
not I_41784 (I713933,I3570);
DFFARX1 I_41785 (I1182915,I3563,I713933,I713959,);
not I_41786 (I713967,I713959);
nand I_41787 (I713984,I1182897,I1182909);
and I_41788 (I714001,I713984,I1182912);
DFFARX1 I_41789 (I714001,I3563,I713933,I714027,);
not I_41790 (I714035,I1182906);
DFFARX1 I_41791 (I1182903,I3563,I713933,I714061,);
not I_41792 (I714069,I714061);
nor I_41793 (I714086,I714069,I713967);
and I_41794 (I714103,I714086,I1182906);
nor I_41795 (I714120,I714069,I714035);
nor I_41796 (I713916,I714027,I714120);
DFFARX1 I_41797 (I1182921,I3563,I713933,I714160,);
nor I_41798 (I714168,I714160,I714027);
not I_41799 (I714185,I714168);
not I_41800 (I714202,I714160);
nor I_41801 (I714219,I714202,I714103);
DFFARX1 I_41802 (I714219,I3563,I713933,I713919,);
nand I_41803 (I714250,I1182900,I1182900);
and I_41804 (I714267,I714250,I1182897);
DFFARX1 I_41805 (I714267,I3563,I713933,I714293,);
nor I_41806 (I714301,I714293,I714160);
DFFARX1 I_41807 (I714301,I3563,I713933,I713901,);
nand I_41808 (I714332,I714293,I714202);
nand I_41809 (I713910,I714185,I714332);
not I_41810 (I714363,I714293);
nor I_41811 (I714380,I714363,I714103);
DFFARX1 I_41812 (I714380,I3563,I713933,I713922,);
nor I_41813 (I714411,I1182918,I1182900);
or I_41814 (I713913,I714160,I714411);
nor I_41815 (I713904,I714293,I714411);
or I_41816 (I713907,I714027,I714411);
DFFARX1 I_41817 (I714411,I3563,I713933,I713925,);
not I_41818 (I714511,I3570);
DFFARX1 I_41819 (I62974,I3563,I714511,I714537,);
not I_41820 (I714545,I714537);
nand I_41821 (I714562,I62983,I62992);
and I_41822 (I714579,I714562,I62971);
DFFARX1 I_41823 (I714579,I3563,I714511,I714605,);
not I_41824 (I714613,I62974);
DFFARX1 I_41825 (I62989,I3563,I714511,I714639,);
not I_41826 (I714647,I714639);
nor I_41827 (I714664,I714647,I714545);
and I_41828 (I714681,I714664,I62974);
nor I_41829 (I714698,I714647,I714613);
nor I_41830 (I714494,I714605,I714698);
DFFARX1 I_41831 (I62980,I3563,I714511,I714738,);
nor I_41832 (I714746,I714738,I714605);
not I_41833 (I714763,I714746);
not I_41834 (I714780,I714738);
nor I_41835 (I714797,I714780,I714681);
DFFARX1 I_41836 (I714797,I3563,I714511,I714497,);
nand I_41837 (I714828,I62995,I62971);
and I_41838 (I714845,I714828,I62977);
DFFARX1 I_41839 (I714845,I3563,I714511,I714871,);
nor I_41840 (I714879,I714871,I714738);
DFFARX1 I_41841 (I714879,I3563,I714511,I714479,);
nand I_41842 (I714910,I714871,I714780);
nand I_41843 (I714488,I714763,I714910);
not I_41844 (I714941,I714871);
nor I_41845 (I714958,I714941,I714681);
DFFARX1 I_41846 (I714958,I3563,I714511,I714500,);
nor I_41847 (I714989,I62986,I62971);
or I_41848 (I714491,I714738,I714989);
nor I_41849 (I714482,I714871,I714989);
or I_41850 (I714485,I714605,I714989);
DFFARX1 I_41851 (I714989,I3563,I714511,I714503,);
not I_41852 (I715089,I3570);
DFFARX1 I_41853 (I602925,I3563,I715089,I715115,);
not I_41854 (I715123,I715115);
nand I_41855 (I715140,I602934,I602943);
and I_41856 (I715157,I715140,I602949);
DFFARX1 I_41857 (I715157,I3563,I715089,I715183,);
not I_41858 (I715191,I602946);
DFFARX1 I_41859 (I602931,I3563,I715089,I715217,);
not I_41860 (I715225,I715217);
nor I_41861 (I715242,I715225,I715123);
and I_41862 (I715259,I715242,I602946);
nor I_41863 (I715276,I715225,I715191);
nor I_41864 (I715072,I715183,I715276);
DFFARX1 I_41865 (I602940,I3563,I715089,I715316,);
nor I_41866 (I715324,I715316,I715183);
not I_41867 (I715341,I715324);
not I_41868 (I715358,I715316);
nor I_41869 (I715375,I715358,I715259);
DFFARX1 I_41870 (I715375,I3563,I715089,I715075,);
nand I_41871 (I715406,I602937,I602928);
and I_41872 (I715423,I715406,I602925);
DFFARX1 I_41873 (I715423,I3563,I715089,I715449,);
nor I_41874 (I715457,I715449,I715316);
DFFARX1 I_41875 (I715457,I3563,I715089,I715057,);
nand I_41876 (I715488,I715449,I715358);
nand I_41877 (I715066,I715341,I715488);
not I_41878 (I715519,I715449);
nor I_41879 (I715536,I715519,I715259);
DFFARX1 I_41880 (I715536,I3563,I715089,I715078,);
nor I_41881 (I715567,I602928,I602928);
or I_41882 (I715069,I715316,I715567);
nor I_41883 (I715060,I715449,I715567);
or I_41884 (I715063,I715183,I715567);
DFFARX1 I_41885 (I715567,I3563,I715089,I715081,);
not I_41886 (I715667,I3570);
DFFARX1 I_41887 (I570336,I3563,I715667,I715693,);
not I_41888 (I715701,I715693);
nand I_41889 (I715718,I570351,I570336);
and I_41890 (I715735,I715718,I570339);
DFFARX1 I_41891 (I715735,I3563,I715667,I715761,);
not I_41892 (I715769,I570339);
DFFARX1 I_41893 (I570348,I3563,I715667,I715795,);
not I_41894 (I715803,I715795);
nor I_41895 (I715820,I715803,I715701);
and I_41896 (I715837,I715820,I570339);
nor I_41897 (I715854,I715803,I715769);
nor I_41898 (I715650,I715761,I715854);
DFFARX1 I_41899 (I570342,I3563,I715667,I715894,);
nor I_41900 (I715902,I715894,I715761);
not I_41901 (I715919,I715902);
not I_41902 (I715936,I715894);
nor I_41903 (I715953,I715936,I715837);
DFFARX1 I_41904 (I715953,I3563,I715667,I715653,);
nand I_41905 (I715984,I570345,I570354);
and I_41906 (I716001,I715984,I570360);
DFFARX1 I_41907 (I716001,I3563,I715667,I716027,);
nor I_41908 (I716035,I716027,I715894);
DFFARX1 I_41909 (I716035,I3563,I715667,I715635,);
nand I_41910 (I716066,I716027,I715936);
nand I_41911 (I715644,I715919,I716066);
not I_41912 (I716097,I716027);
nor I_41913 (I716114,I716097,I715837);
DFFARX1 I_41914 (I716114,I3563,I715667,I715656,);
nor I_41915 (I716145,I570357,I570354);
or I_41916 (I715647,I715894,I716145);
nor I_41917 (I715638,I716027,I716145);
or I_41918 (I715641,I715761,I716145);
DFFARX1 I_41919 (I716145,I3563,I715667,I715659,);
not I_41920 (I716245,I3570);
DFFARX1 I_41921 (I460491,I3563,I716245,I716271,);
not I_41922 (I716279,I716271);
nand I_41923 (I716296,I460482,I460500);
and I_41924 (I716313,I716296,I460503);
DFFARX1 I_41925 (I716313,I3563,I716245,I716339,);
not I_41926 (I716347,I460497);
DFFARX1 I_41927 (I460485,I3563,I716245,I716373,);
not I_41928 (I716381,I716373);
nor I_41929 (I716398,I716381,I716279);
and I_41930 (I716415,I716398,I460497);
nor I_41931 (I716432,I716381,I716347);
nor I_41932 (I716228,I716339,I716432);
DFFARX1 I_41933 (I460494,I3563,I716245,I716472,);
nor I_41934 (I716480,I716472,I716339);
not I_41935 (I716497,I716480);
not I_41936 (I716514,I716472);
nor I_41937 (I716531,I716514,I716415);
DFFARX1 I_41938 (I716531,I3563,I716245,I716231,);
nand I_41939 (I716562,I460509,I460506);
and I_41940 (I716579,I716562,I460488);
DFFARX1 I_41941 (I716579,I3563,I716245,I716605,);
nor I_41942 (I716613,I716605,I716472);
DFFARX1 I_41943 (I716613,I3563,I716245,I716213,);
nand I_41944 (I716644,I716605,I716514);
nand I_41945 (I716222,I716497,I716644);
not I_41946 (I716675,I716605);
nor I_41947 (I716692,I716675,I716415);
DFFARX1 I_41948 (I716692,I3563,I716245,I716234,);
nor I_41949 (I716723,I460482,I460506);
or I_41950 (I716225,I716472,I716723);
nor I_41951 (I716216,I716605,I716723);
or I_41952 (I716219,I716339,I716723);
DFFARX1 I_41953 (I716723,I3563,I716245,I716237,);
not I_41954 (I716823,I3570);
DFFARX1 I_41955 (I840056,I3563,I716823,I716849,);
not I_41956 (I716857,I716849);
nand I_41957 (I716874,I840044,I840062);
and I_41958 (I716891,I716874,I840059);
DFFARX1 I_41959 (I716891,I3563,I716823,I716917,);
not I_41960 (I716925,I840050);
DFFARX1 I_41961 (I840047,I3563,I716823,I716951,);
not I_41962 (I716959,I716951);
nor I_41963 (I716976,I716959,I716857);
and I_41964 (I716993,I716976,I840050);
nor I_41965 (I717010,I716959,I716925);
nor I_41966 (I716806,I716917,I717010);
DFFARX1 I_41967 (I840041,I3563,I716823,I717050,);
nor I_41968 (I717058,I717050,I716917);
not I_41969 (I717075,I717058);
not I_41970 (I717092,I717050);
nor I_41971 (I717109,I717092,I716993);
DFFARX1 I_41972 (I717109,I3563,I716823,I716809,);
nand I_41973 (I717140,I840041,I840044);
and I_41974 (I717157,I717140,I840047);
DFFARX1 I_41975 (I717157,I3563,I716823,I717183,);
nor I_41976 (I717191,I717183,I717050);
DFFARX1 I_41977 (I717191,I3563,I716823,I716791,);
nand I_41978 (I717222,I717183,I717092);
nand I_41979 (I716800,I717075,I717222);
not I_41980 (I717253,I717183);
nor I_41981 (I717270,I717253,I716993);
DFFARX1 I_41982 (I717270,I3563,I716823,I716812,);
nor I_41983 (I717301,I840053,I840044);
or I_41984 (I716803,I717050,I717301);
nor I_41985 (I716794,I717183,I717301);
or I_41986 (I716797,I716917,I717301);
DFFARX1 I_41987 (I717301,I3563,I716823,I716815,);
not I_41988 (I717401,I3570);
DFFARX1 I_41989 (I1001463,I3563,I717401,I717427,);
not I_41990 (I717435,I717427);
nand I_41991 (I717452,I1001439,I1001454);
and I_41992 (I717469,I717452,I1001466);
DFFARX1 I_41993 (I717469,I3563,I717401,I717495,);
not I_41994 (I717503,I1001451);
DFFARX1 I_41995 (I1001442,I3563,I717401,I717529,);
not I_41996 (I717537,I717529);
nor I_41997 (I717554,I717537,I717435);
and I_41998 (I717571,I717554,I1001451);
nor I_41999 (I717588,I717537,I717503);
nor I_42000 (I717384,I717495,I717588);
DFFARX1 I_42001 (I1001439,I3563,I717401,I717628,);
nor I_42002 (I717636,I717628,I717495);
not I_42003 (I717653,I717636);
not I_42004 (I717670,I717628);
nor I_42005 (I717687,I717670,I717571);
DFFARX1 I_42006 (I717687,I3563,I717401,I717387,);
nand I_42007 (I717718,I1001457,I1001448);
and I_42008 (I717735,I717718,I1001460);
DFFARX1 I_42009 (I717735,I3563,I717401,I717761,);
nor I_42010 (I717769,I717761,I717628);
DFFARX1 I_42011 (I717769,I3563,I717401,I717369,);
nand I_42012 (I717800,I717761,I717670);
nand I_42013 (I717378,I717653,I717800);
not I_42014 (I717831,I717761);
nor I_42015 (I717848,I717831,I717571);
DFFARX1 I_42016 (I717848,I3563,I717401,I717390,);
nor I_42017 (I717879,I1001445,I1001448);
or I_42018 (I717381,I717628,I717879);
nor I_42019 (I717372,I717761,I717879);
or I_42020 (I717375,I717495,I717879);
DFFARX1 I_42021 (I717879,I3563,I717401,I717393,);
not I_42022 (I717979,I3570);
DFFARX1 I_42023 (I374452,I3563,I717979,I718005,);
not I_42024 (I718013,I718005);
nand I_42025 (I718030,I374455,I374431);
and I_42026 (I718047,I718030,I374428);
DFFARX1 I_42027 (I718047,I3563,I717979,I718073,);
not I_42028 (I718081,I374434);
DFFARX1 I_42029 (I374428,I3563,I717979,I718107,);
not I_42030 (I718115,I718107);
nor I_42031 (I718132,I718115,I718013);
and I_42032 (I718149,I718132,I374434);
nor I_42033 (I718166,I718115,I718081);
nor I_42034 (I717962,I718073,I718166);
DFFARX1 I_42035 (I374437,I3563,I717979,I718206,);
nor I_42036 (I718214,I718206,I718073);
not I_42037 (I718231,I718214);
not I_42038 (I718248,I718206);
nor I_42039 (I718265,I718248,I718149);
DFFARX1 I_42040 (I718265,I3563,I717979,I717965,);
nand I_42041 (I718296,I374440,I374449);
and I_42042 (I718313,I718296,I374446);
DFFARX1 I_42043 (I718313,I3563,I717979,I718339,);
nor I_42044 (I718347,I718339,I718206);
DFFARX1 I_42045 (I718347,I3563,I717979,I717947,);
nand I_42046 (I718378,I718339,I718248);
nand I_42047 (I717956,I718231,I718378);
not I_42048 (I718409,I718339);
nor I_42049 (I718426,I718409,I718149);
DFFARX1 I_42050 (I718426,I3563,I717979,I717968,);
nor I_42051 (I718457,I374443,I374449);
or I_42052 (I717959,I718206,I718457);
nor I_42053 (I717950,I718339,I718457);
or I_42054 (I717953,I718073,I718457);
DFFARX1 I_42055 (I718457,I3563,I717979,I717971,);
not I_42056 (I718557,I3570);
DFFARX1 I_42057 (I544751,I3563,I718557,I718583,);
not I_42058 (I718591,I718583);
nand I_42059 (I718608,I544766,I544751);
and I_42060 (I718625,I718608,I544754);
DFFARX1 I_42061 (I718625,I3563,I718557,I718651,);
not I_42062 (I718659,I544754);
DFFARX1 I_42063 (I544763,I3563,I718557,I718685,);
not I_42064 (I718693,I718685);
nor I_42065 (I718710,I718693,I718591);
and I_42066 (I718727,I718710,I544754);
nor I_42067 (I718744,I718693,I718659);
nor I_42068 (I718540,I718651,I718744);
DFFARX1 I_42069 (I544757,I3563,I718557,I718784,);
nor I_42070 (I718792,I718784,I718651);
not I_42071 (I718809,I718792);
not I_42072 (I718826,I718784);
nor I_42073 (I718843,I718826,I718727);
DFFARX1 I_42074 (I718843,I3563,I718557,I718543,);
nand I_42075 (I718874,I544760,I544769);
and I_42076 (I718891,I718874,I544775);
DFFARX1 I_42077 (I718891,I3563,I718557,I718917,);
nor I_42078 (I718925,I718917,I718784);
DFFARX1 I_42079 (I718925,I3563,I718557,I718525,);
nand I_42080 (I718956,I718917,I718826);
nand I_42081 (I718534,I718809,I718956);
not I_42082 (I718987,I718917);
nor I_42083 (I719004,I718987,I718727);
DFFARX1 I_42084 (I719004,I3563,I718557,I718546,);
nor I_42085 (I719035,I544772,I544769);
or I_42086 (I718537,I718784,I719035);
nor I_42087 (I718528,I718917,I719035);
or I_42088 (I718531,I718651,I719035);
DFFARX1 I_42089 (I719035,I3563,I718557,I718549,);
not I_42090 (I719135,I3570);
DFFARX1 I_42091 (I579805,I3563,I719135,I719161,);
not I_42092 (I719169,I719161);
nand I_42093 (I719186,I579814,I579823);
and I_42094 (I719203,I719186,I579829);
DFFARX1 I_42095 (I719203,I3563,I719135,I719229,);
not I_42096 (I719237,I579826);
DFFARX1 I_42097 (I579811,I3563,I719135,I719263,);
not I_42098 (I719271,I719263);
nor I_42099 (I719288,I719271,I719169);
and I_42100 (I719305,I719288,I579826);
nor I_42101 (I719322,I719271,I719237);
nor I_42102 (I719118,I719229,I719322);
DFFARX1 I_42103 (I579820,I3563,I719135,I719362,);
nor I_42104 (I719370,I719362,I719229);
not I_42105 (I719387,I719370);
not I_42106 (I719404,I719362);
nor I_42107 (I719421,I719404,I719305);
DFFARX1 I_42108 (I719421,I3563,I719135,I719121,);
nand I_42109 (I719452,I579817,I579808);
and I_42110 (I719469,I719452,I579805);
DFFARX1 I_42111 (I719469,I3563,I719135,I719495,);
nor I_42112 (I719503,I719495,I719362);
DFFARX1 I_42113 (I719503,I3563,I719135,I719103,);
nand I_42114 (I719534,I719495,I719404);
nand I_42115 (I719112,I719387,I719534);
not I_42116 (I719565,I719495);
nor I_42117 (I719582,I719565,I719305);
DFFARX1 I_42118 (I719582,I3563,I719135,I719124,);
nor I_42119 (I719613,I579808,I579808);
or I_42120 (I719115,I719362,I719613);
nor I_42121 (I719106,I719495,I719613);
or I_42122 (I719109,I719229,I719613);
DFFARX1 I_42123 (I719613,I3563,I719135,I719127,);
not I_42124 (I719713,I3570);
DFFARX1 I_42125 (I180373,I3563,I719713,I719739,);
not I_42126 (I719747,I719739);
nand I_42127 (I719764,I180376,I180397);
and I_42128 (I719781,I719764,I180385);
DFFARX1 I_42129 (I719781,I3563,I719713,I719807,);
not I_42130 (I719815,I180382);
DFFARX1 I_42131 (I180373,I3563,I719713,I719841,);
not I_42132 (I719849,I719841);
nor I_42133 (I719866,I719849,I719747);
and I_42134 (I719883,I719866,I180382);
nor I_42135 (I719900,I719849,I719815);
nor I_42136 (I719696,I719807,I719900);
DFFARX1 I_42137 (I180391,I3563,I719713,I719940,);
nor I_42138 (I719948,I719940,I719807);
not I_42139 (I719965,I719948);
not I_42140 (I719982,I719940);
nor I_42141 (I719999,I719982,I719883);
DFFARX1 I_42142 (I719999,I3563,I719713,I719699,);
nand I_42143 (I720030,I180376,I180379);
and I_42144 (I720047,I720030,I180388);
DFFARX1 I_42145 (I720047,I3563,I719713,I720073,);
nor I_42146 (I720081,I720073,I719940);
DFFARX1 I_42147 (I720081,I3563,I719713,I719681,);
nand I_42148 (I720112,I720073,I719982);
nand I_42149 (I719690,I719965,I720112);
not I_42150 (I720143,I720073);
nor I_42151 (I720160,I720143,I719883);
DFFARX1 I_42152 (I720160,I3563,I719713,I719702,);
nor I_42153 (I720191,I180394,I180379);
or I_42154 (I719693,I719940,I720191);
nor I_42155 (I719684,I720073,I720191);
or I_42156 (I719687,I719807,I720191);
DFFARX1 I_42157 (I720191,I3563,I719713,I719705,);
not I_42158 (I720291,I3570);
DFFARX1 I_42159 (I179183,I3563,I720291,I720317,);
not I_42160 (I720325,I720317);
nand I_42161 (I720342,I179186,I179207);
and I_42162 (I720359,I720342,I179195);
DFFARX1 I_42163 (I720359,I3563,I720291,I720385,);
not I_42164 (I720393,I179192);
DFFARX1 I_42165 (I179183,I3563,I720291,I720419,);
not I_42166 (I720427,I720419);
nor I_42167 (I720444,I720427,I720325);
and I_42168 (I720461,I720444,I179192);
nor I_42169 (I720478,I720427,I720393);
nor I_42170 (I720274,I720385,I720478);
DFFARX1 I_42171 (I179201,I3563,I720291,I720518,);
nor I_42172 (I720526,I720518,I720385);
not I_42173 (I720543,I720526);
not I_42174 (I720560,I720518);
nor I_42175 (I720577,I720560,I720461);
DFFARX1 I_42176 (I720577,I3563,I720291,I720277,);
nand I_42177 (I720608,I179186,I179189);
and I_42178 (I720625,I720608,I179198);
DFFARX1 I_42179 (I720625,I3563,I720291,I720651,);
nor I_42180 (I720659,I720651,I720518);
DFFARX1 I_42181 (I720659,I3563,I720291,I720259,);
nand I_42182 (I720690,I720651,I720560);
nand I_42183 (I720268,I720543,I720690);
not I_42184 (I720721,I720651);
nor I_42185 (I720738,I720721,I720461);
DFFARX1 I_42186 (I720738,I3563,I720291,I720280,);
nor I_42187 (I720769,I179204,I179189);
or I_42188 (I720271,I720518,I720769);
nor I_42189 (I720262,I720651,I720769);
or I_42190 (I720265,I720385,I720769);
DFFARX1 I_42191 (I720769,I3563,I720291,I720283,);
not I_42192 (I720869,I3570);
DFFARX1 I_42193 (I1261641,I3563,I720869,I720895,);
not I_42194 (I720903,I720895);
nand I_42195 (I720920,I1261644,I1261653);
and I_42196 (I720937,I720920,I1261656);
DFFARX1 I_42197 (I720937,I3563,I720869,I720963,);
not I_42198 (I720971,I1261665);
DFFARX1 I_42199 (I1261647,I3563,I720869,I720997,);
not I_42200 (I721005,I720997);
nor I_42201 (I721022,I721005,I720903);
and I_42202 (I721039,I721022,I1261665);
nor I_42203 (I721056,I721005,I720971);
nor I_42204 (I720852,I720963,I721056);
DFFARX1 I_42205 (I1261644,I3563,I720869,I721096,);
nor I_42206 (I721104,I721096,I720963);
not I_42207 (I721121,I721104);
not I_42208 (I721138,I721096);
nor I_42209 (I721155,I721138,I721039);
DFFARX1 I_42210 (I721155,I3563,I720869,I720855,);
nand I_42211 (I721186,I1261662,I1261641);
and I_42212 (I721203,I721186,I1261659);
DFFARX1 I_42213 (I721203,I3563,I720869,I721229,);
nor I_42214 (I721237,I721229,I721096);
DFFARX1 I_42215 (I721237,I3563,I720869,I720837,);
nand I_42216 (I721268,I721229,I721138);
nand I_42217 (I720846,I721121,I721268);
not I_42218 (I721299,I721229);
nor I_42219 (I721316,I721299,I721039);
DFFARX1 I_42220 (I721316,I3563,I720869,I720858,);
nor I_42221 (I721347,I1261650,I1261641);
or I_42222 (I720849,I721096,I721347);
nor I_42223 (I720840,I721229,I721347);
or I_42224 (I720843,I720963,I721347);
DFFARX1 I_42225 (I721347,I3563,I720869,I720861,);
not I_42226 (I721447,I3570);
DFFARX1 I_42227 (I906458,I3563,I721447,I721473,);
not I_42228 (I721481,I721473);
nand I_42229 (I721498,I906446,I906464);
and I_42230 (I721515,I721498,I906461);
DFFARX1 I_42231 (I721515,I3563,I721447,I721541,);
not I_42232 (I721549,I906452);
DFFARX1 I_42233 (I906449,I3563,I721447,I721575,);
not I_42234 (I721583,I721575);
nor I_42235 (I721600,I721583,I721481);
and I_42236 (I721617,I721600,I906452);
nor I_42237 (I721634,I721583,I721549);
nor I_42238 (I721430,I721541,I721634);
DFFARX1 I_42239 (I906443,I3563,I721447,I721674,);
nor I_42240 (I721682,I721674,I721541);
not I_42241 (I721699,I721682);
not I_42242 (I721716,I721674);
nor I_42243 (I721733,I721716,I721617);
DFFARX1 I_42244 (I721733,I3563,I721447,I721433,);
nand I_42245 (I721764,I906443,I906446);
and I_42246 (I721781,I721764,I906449);
DFFARX1 I_42247 (I721781,I3563,I721447,I721807,);
nor I_42248 (I721815,I721807,I721674);
DFFARX1 I_42249 (I721815,I3563,I721447,I721415,);
nand I_42250 (I721846,I721807,I721716);
nand I_42251 (I721424,I721699,I721846);
not I_42252 (I721877,I721807);
nor I_42253 (I721894,I721877,I721617);
DFFARX1 I_42254 (I721894,I3563,I721447,I721436,);
nor I_42255 (I721925,I906455,I906446);
or I_42256 (I721427,I721674,I721925);
nor I_42257 (I721418,I721807,I721925);
or I_42258 (I721421,I721541,I721925);
DFFARX1 I_42259 (I721925,I3563,I721447,I721439,);
not I_42260 (I722025,I3570);
DFFARX1 I_42261 (I71406,I3563,I722025,I722051,);
not I_42262 (I722059,I722051);
nand I_42263 (I722076,I71415,I71424);
and I_42264 (I722093,I722076,I71403);
DFFARX1 I_42265 (I722093,I3563,I722025,I722119,);
not I_42266 (I722127,I71406);
DFFARX1 I_42267 (I71421,I3563,I722025,I722153,);
not I_42268 (I722161,I722153);
nor I_42269 (I722178,I722161,I722059);
and I_42270 (I722195,I722178,I71406);
nor I_42271 (I722212,I722161,I722127);
nor I_42272 (I722008,I722119,I722212);
DFFARX1 I_42273 (I71412,I3563,I722025,I722252,);
nor I_42274 (I722260,I722252,I722119);
not I_42275 (I722277,I722260);
not I_42276 (I722294,I722252);
nor I_42277 (I722311,I722294,I722195);
DFFARX1 I_42278 (I722311,I3563,I722025,I722011,);
nand I_42279 (I722342,I71427,I71403);
and I_42280 (I722359,I722342,I71409);
DFFARX1 I_42281 (I722359,I3563,I722025,I722385,);
nor I_42282 (I722393,I722385,I722252);
DFFARX1 I_42283 (I722393,I3563,I722025,I721993,);
nand I_42284 (I722424,I722385,I722294);
nand I_42285 (I722002,I722277,I722424);
not I_42286 (I722455,I722385);
nor I_42287 (I722472,I722455,I722195);
DFFARX1 I_42288 (I722472,I3563,I722025,I722014,);
nor I_42289 (I722503,I71418,I71403);
or I_42290 (I722005,I722252,I722503);
nor I_42291 (I721996,I722385,I722503);
or I_42292 (I721999,I722119,I722503);
DFFARX1 I_42293 (I722503,I3563,I722025,I722017,);
not I_42294 (I722603,I3570);
DFFARX1 I_42295 (I303834,I3563,I722603,I722629,);
not I_42296 (I722637,I722629);
nand I_42297 (I722654,I303837,I303813);
and I_42298 (I722671,I722654,I303810);
DFFARX1 I_42299 (I722671,I3563,I722603,I722697,);
not I_42300 (I722705,I303816);
DFFARX1 I_42301 (I303810,I3563,I722603,I722731,);
not I_42302 (I722739,I722731);
nor I_42303 (I722756,I722739,I722637);
and I_42304 (I722773,I722756,I303816);
nor I_42305 (I722790,I722739,I722705);
nor I_42306 (I722586,I722697,I722790);
DFFARX1 I_42307 (I303819,I3563,I722603,I722830,);
nor I_42308 (I722838,I722830,I722697);
not I_42309 (I722855,I722838);
not I_42310 (I722872,I722830);
nor I_42311 (I722889,I722872,I722773);
DFFARX1 I_42312 (I722889,I3563,I722603,I722589,);
nand I_42313 (I722920,I303822,I303831);
and I_42314 (I722937,I722920,I303828);
DFFARX1 I_42315 (I722937,I3563,I722603,I722963,);
nor I_42316 (I722971,I722963,I722830);
DFFARX1 I_42317 (I722971,I3563,I722603,I722571,);
nand I_42318 (I723002,I722963,I722872);
nand I_42319 (I722580,I722855,I723002);
not I_42320 (I723033,I722963);
nor I_42321 (I723050,I723033,I722773);
DFFARX1 I_42322 (I723050,I3563,I722603,I722592,);
nor I_42323 (I723081,I303825,I303831);
or I_42324 (I722583,I722830,I723081);
nor I_42325 (I722574,I722963,I723081);
or I_42326 (I722577,I722697,I723081);
DFFARX1 I_42327 (I723081,I3563,I722603,I722595,);
not I_42328 (I723181,I3570);
DFFARX1 I_42329 (I622577,I3563,I723181,I723207,);
not I_42330 (I723215,I723207);
nand I_42331 (I723232,I622586,I622595);
and I_42332 (I723249,I723232,I622601);
DFFARX1 I_42333 (I723249,I3563,I723181,I723275,);
not I_42334 (I723283,I622598);
DFFARX1 I_42335 (I622583,I3563,I723181,I723309,);
not I_42336 (I723317,I723309);
nor I_42337 (I723334,I723317,I723215);
and I_42338 (I723351,I723334,I622598);
nor I_42339 (I723368,I723317,I723283);
nor I_42340 (I723164,I723275,I723368);
DFFARX1 I_42341 (I622592,I3563,I723181,I723408,);
nor I_42342 (I723416,I723408,I723275);
not I_42343 (I723433,I723416);
not I_42344 (I723450,I723408);
nor I_42345 (I723467,I723450,I723351);
DFFARX1 I_42346 (I723467,I3563,I723181,I723167,);
nand I_42347 (I723498,I622589,I622580);
and I_42348 (I723515,I723498,I622577);
DFFARX1 I_42349 (I723515,I3563,I723181,I723541,);
nor I_42350 (I723549,I723541,I723408);
DFFARX1 I_42351 (I723549,I3563,I723181,I723149,);
nand I_42352 (I723580,I723541,I723450);
nand I_42353 (I723158,I723433,I723580);
not I_42354 (I723611,I723541);
nor I_42355 (I723628,I723611,I723351);
DFFARX1 I_42356 (I723628,I3563,I723181,I723170,);
nor I_42357 (I723659,I622580,I622580);
or I_42358 (I723161,I723408,I723659);
nor I_42359 (I723152,I723541,I723659);
or I_42360 (I723155,I723275,I723659);
DFFARX1 I_42361 (I723659,I3563,I723181,I723173,);
not I_42362 (I723759,I3570);
DFFARX1 I_42363 (I90378,I3563,I723759,I723785,);
not I_42364 (I723793,I723785);
nand I_42365 (I723810,I90387,I90396);
and I_42366 (I723827,I723810,I90375);
DFFARX1 I_42367 (I723827,I3563,I723759,I723853,);
not I_42368 (I723861,I90378);
DFFARX1 I_42369 (I90393,I3563,I723759,I723887,);
not I_42370 (I723895,I723887);
nor I_42371 (I723912,I723895,I723793);
and I_42372 (I723929,I723912,I90378);
nor I_42373 (I723946,I723895,I723861);
nor I_42374 (I723742,I723853,I723946);
DFFARX1 I_42375 (I90384,I3563,I723759,I723986,);
nor I_42376 (I723994,I723986,I723853);
not I_42377 (I724011,I723994);
not I_42378 (I724028,I723986);
nor I_42379 (I724045,I724028,I723929);
DFFARX1 I_42380 (I724045,I3563,I723759,I723745,);
nand I_42381 (I724076,I90399,I90375);
and I_42382 (I724093,I724076,I90381);
DFFARX1 I_42383 (I724093,I3563,I723759,I724119,);
nor I_42384 (I724127,I724119,I723986);
DFFARX1 I_42385 (I724127,I3563,I723759,I723727,);
nand I_42386 (I724158,I724119,I724028);
nand I_42387 (I723736,I724011,I724158);
not I_42388 (I724189,I724119);
nor I_42389 (I724206,I724189,I723929);
DFFARX1 I_42390 (I724206,I3563,I723759,I723748,);
nor I_42391 (I724237,I90390,I90375);
or I_42392 (I723739,I723986,I724237);
nor I_42393 (I723730,I724119,I724237);
or I_42394 (I723733,I723853,I724237);
DFFARX1 I_42395 (I724237,I3563,I723759,I723751,);
not I_42396 (I724337,I3570);
DFFARX1 I_42397 (I1249129,I3563,I724337,I724363,);
not I_42398 (I724371,I724363);
nand I_42399 (I724388,I1249132,I1249141);
and I_42400 (I724405,I724388,I1249144);
DFFARX1 I_42401 (I724405,I3563,I724337,I724431,);
not I_42402 (I724439,I1249153);
DFFARX1 I_42403 (I1249135,I3563,I724337,I724465,);
not I_42404 (I724473,I724465);
nor I_42405 (I724490,I724473,I724371);
and I_42406 (I724507,I724490,I1249153);
nor I_42407 (I724524,I724473,I724439);
nor I_42408 (I724320,I724431,I724524);
DFFARX1 I_42409 (I1249132,I3563,I724337,I724564,);
nor I_42410 (I724572,I724564,I724431);
not I_42411 (I724589,I724572);
not I_42412 (I724606,I724564);
nor I_42413 (I724623,I724606,I724507);
DFFARX1 I_42414 (I724623,I3563,I724337,I724323,);
nand I_42415 (I724654,I1249150,I1249129);
and I_42416 (I724671,I724654,I1249147);
DFFARX1 I_42417 (I724671,I3563,I724337,I724697,);
nor I_42418 (I724705,I724697,I724564);
DFFARX1 I_42419 (I724705,I3563,I724337,I724305,);
nand I_42420 (I724736,I724697,I724606);
nand I_42421 (I724314,I724589,I724736);
not I_42422 (I724767,I724697);
nor I_42423 (I724784,I724767,I724507);
DFFARX1 I_42424 (I724784,I3563,I724337,I724326,);
nor I_42425 (I724815,I1249138,I1249129);
or I_42426 (I724317,I724564,I724815);
nor I_42427 (I724308,I724697,I724815);
or I_42428 (I724311,I724431,I724815);
DFFARX1 I_42429 (I724815,I3563,I724337,I724329,);
not I_42430 (I724915,I3570);
DFFARX1 I_42431 (I863244,I3563,I724915,I724941,);
not I_42432 (I724949,I724941);
nand I_42433 (I724966,I863232,I863250);
and I_42434 (I724983,I724966,I863247);
DFFARX1 I_42435 (I724983,I3563,I724915,I725009,);
not I_42436 (I725017,I863238);
DFFARX1 I_42437 (I863235,I3563,I724915,I725043,);
not I_42438 (I725051,I725043);
nor I_42439 (I725068,I725051,I724949);
and I_42440 (I725085,I725068,I863238);
nor I_42441 (I725102,I725051,I725017);
nor I_42442 (I724898,I725009,I725102);
DFFARX1 I_42443 (I863229,I3563,I724915,I725142,);
nor I_42444 (I725150,I725142,I725009);
not I_42445 (I725167,I725150);
not I_42446 (I725184,I725142);
nor I_42447 (I725201,I725184,I725085);
DFFARX1 I_42448 (I725201,I3563,I724915,I724901,);
nand I_42449 (I725232,I863229,I863232);
and I_42450 (I725249,I725232,I863235);
DFFARX1 I_42451 (I725249,I3563,I724915,I725275,);
nor I_42452 (I725283,I725275,I725142);
DFFARX1 I_42453 (I725283,I3563,I724915,I724883,);
nand I_42454 (I725314,I725275,I725184);
nand I_42455 (I724892,I725167,I725314);
not I_42456 (I725345,I725275);
nor I_42457 (I725362,I725345,I725085);
DFFARX1 I_42458 (I725362,I3563,I724915,I724904,);
nor I_42459 (I725393,I863241,I863232);
or I_42460 (I724895,I725142,I725393);
nor I_42461 (I724886,I725275,I725393);
or I_42462 (I724889,I725009,I725393);
DFFARX1 I_42463 (I725393,I3563,I724915,I724907,);
not I_42464 (I725493,I3570);
DFFARX1 I_42465 (I884324,I3563,I725493,I725519,);
not I_42466 (I725527,I725519);
nand I_42467 (I725544,I884312,I884330);
and I_42468 (I725561,I725544,I884327);
DFFARX1 I_42469 (I725561,I3563,I725493,I725587,);
not I_42470 (I725595,I884318);
DFFARX1 I_42471 (I884315,I3563,I725493,I725621,);
not I_42472 (I725629,I725621);
nor I_42473 (I725646,I725629,I725527);
and I_42474 (I725663,I725646,I884318);
nor I_42475 (I725680,I725629,I725595);
nor I_42476 (I725476,I725587,I725680);
DFFARX1 I_42477 (I884309,I3563,I725493,I725720,);
nor I_42478 (I725728,I725720,I725587);
not I_42479 (I725745,I725728);
not I_42480 (I725762,I725720);
nor I_42481 (I725779,I725762,I725663);
DFFARX1 I_42482 (I725779,I3563,I725493,I725479,);
nand I_42483 (I725810,I884309,I884312);
and I_42484 (I725827,I725810,I884315);
DFFARX1 I_42485 (I725827,I3563,I725493,I725853,);
nor I_42486 (I725861,I725853,I725720);
DFFARX1 I_42487 (I725861,I3563,I725493,I725461,);
nand I_42488 (I725892,I725853,I725762);
nand I_42489 (I725470,I725745,I725892);
not I_42490 (I725923,I725853);
nor I_42491 (I725940,I725923,I725663);
DFFARX1 I_42492 (I725940,I3563,I725493,I725482,);
nor I_42493 (I725971,I884321,I884312);
or I_42494 (I725473,I725720,I725971);
nor I_42495 (I725464,I725853,I725971);
or I_42496 (I725467,I725587,I725971);
DFFARX1 I_42497 (I725971,I3563,I725493,I725485,);
not I_42498 (I726071,I3570);
DFFARX1 I_42499 (I469739,I3563,I726071,I726097,);
not I_42500 (I726105,I726097);
nand I_42501 (I726122,I469730,I469748);
and I_42502 (I726139,I726122,I469751);
DFFARX1 I_42503 (I726139,I3563,I726071,I726165,);
not I_42504 (I726173,I469745);
DFFARX1 I_42505 (I469733,I3563,I726071,I726199,);
not I_42506 (I726207,I726199);
nor I_42507 (I726224,I726207,I726105);
and I_42508 (I726241,I726224,I469745);
nor I_42509 (I726258,I726207,I726173);
nor I_42510 (I726054,I726165,I726258);
DFFARX1 I_42511 (I469742,I3563,I726071,I726298,);
nor I_42512 (I726306,I726298,I726165);
not I_42513 (I726323,I726306);
not I_42514 (I726340,I726298);
nor I_42515 (I726357,I726340,I726241);
DFFARX1 I_42516 (I726357,I3563,I726071,I726057,);
nand I_42517 (I726388,I469757,I469754);
and I_42518 (I726405,I726388,I469736);
DFFARX1 I_42519 (I726405,I3563,I726071,I726431,);
nor I_42520 (I726439,I726431,I726298);
DFFARX1 I_42521 (I726439,I3563,I726071,I726039,);
nand I_42522 (I726470,I726431,I726340);
nand I_42523 (I726048,I726323,I726470);
not I_42524 (I726501,I726431);
nor I_42525 (I726518,I726501,I726241);
DFFARX1 I_42526 (I726518,I3563,I726071,I726060,);
nor I_42527 (I726549,I469730,I469754);
or I_42528 (I726051,I726298,I726549);
nor I_42529 (I726042,I726431,I726549);
or I_42530 (I726045,I726165,I726549);
DFFARX1 I_42531 (I726549,I3563,I726071,I726063,);
not I_42532 (I726649,I3570);
DFFARX1 I_42533 (I474091,I3563,I726649,I726675,);
not I_42534 (I726683,I726675);
nand I_42535 (I726700,I474082,I474100);
and I_42536 (I726717,I726700,I474103);
DFFARX1 I_42537 (I726717,I3563,I726649,I726743,);
not I_42538 (I726751,I474097);
DFFARX1 I_42539 (I474085,I3563,I726649,I726777,);
not I_42540 (I726785,I726777);
nor I_42541 (I726802,I726785,I726683);
and I_42542 (I726819,I726802,I474097);
nor I_42543 (I726836,I726785,I726751);
nor I_42544 (I726632,I726743,I726836);
DFFARX1 I_42545 (I474094,I3563,I726649,I726876,);
nor I_42546 (I726884,I726876,I726743);
not I_42547 (I726901,I726884);
not I_42548 (I726918,I726876);
nor I_42549 (I726935,I726918,I726819);
DFFARX1 I_42550 (I726935,I3563,I726649,I726635,);
nand I_42551 (I726966,I474109,I474106);
and I_42552 (I726983,I726966,I474088);
DFFARX1 I_42553 (I726983,I3563,I726649,I727009,);
nor I_42554 (I727017,I727009,I726876);
DFFARX1 I_42555 (I727017,I3563,I726649,I726617,);
nand I_42556 (I727048,I727009,I726918);
nand I_42557 (I726626,I726901,I727048);
not I_42558 (I727079,I727009);
nor I_42559 (I727096,I727079,I726819);
DFFARX1 I_42560 (I727096,I3563,I726649,I726638,);
nor I_42561 (I727127,I474082,I474106);
or I_42562 (I726629,I726876,I727127);
nor I_42563 (I726620,I727009,I727127);
or I_42564 (I726623,I726743,I727127);
DFFARX1 I_42565 (I727127,I3563,I726649,I726641,);
not I_42566 (I727227,I3570);
DFFARX1 I_42567 (I607549,I3563,I727227,I727253,);
not I_42568 (I727261,I727253);
nand I_42569 (I727278,I607558,I607567);
and I_42570 (I727295,I727278,I607573);
DFFARX1 I_42571 (I727295,I3563,I727227,I727321,);
not I_42572 (I727329,I607570);
DFFARX1 I_42573 (I607555,I3563,I727227,I727355,);
not I_42574 (I727363,I727355);
nor I_42575 (I727380,I727363,I727261);
and I_42576 (I727397,I727380,I607570);
nor I_42577 (I727414,I727363,I727329);
nor I_42578 (I727210,I727321,I727414);
DFFARX1 I_42579 (I607564,I3563,I727227,I727454,);
nor I_42580 (I727462,I727454,I727321);
not I_42581 (I727479,I727462);
not I_42582 (I727496,I727454);
nor I_42583 (I727513,I727496,I727397);
DFFARX1 I_42584 (I727513,I3563,I727227,I727213,);
nand I_42585 (I727544,I607561,I607552);
and I_42586 (I727561,I727544,I607549);
DFFARX1 I_42587 (I727561,I3563,I727227,I727587,);
nor I_42588 (I727595,I727587,I727454);
DFFARX1 I_42589 (I727595,I3563,I727227,I727195,);
nand I_42590 (I727626,I727587,I727496);
nand I_42591 (I727204,I727479,I727626);
not I_42592 (I727657,I727587);
nor I_42593 (I727674,I727657,I727397);
DFFARX1 I_42594 (I727674,I3563,I727227,I727216,);
nor I_42595 (I727705,I607552,I607552);
or I_42596 (I727207,I727454,I727705);
nor I_42597 (I727198,I727587,I727705);
or I_42598 (I727201,I727321,I727705);
DFFARX1 I_42599 (I727705,I3563,I727227,I727219,);
not I_42600 (I727805,I3570);
DFFARX1 I_42601 (I835313,I3563,I727805,I727831,);
not I_42602 (I727839,I727831);
nand I_42603 (I727856,I835301,I835319);
and I_42604 (I727873,I727856,I835316);
DFFARX1 I_42605 (I727873,I3563,I727805,I727899,);
not I_42606 (I727907,I835307);
DFFARX1 I_42607 (I835304,I3563,I727805,I727933,);
not I_42608 (I727941,I727933);
nor I_42609 (I727958,I727941,I727839);
and I_42610 (I727975,I727958,I835307);
nor I_42611 (I727992,I727941,I727907);
nor I_42612 (I727788,I727899,I727992);
DFFARX1 I_42613 (I835298,I3563,I727805,I728032,);
nor I_42614 (I728040,I728032,I727899);
not I_42615 (I728057,I728040);
not I_42616 (I728074,I728032);
nor I_42617 (I728091,I728074,I727975);
DFFARX1 I_42618 (I728091,I3563,I727805,I727791,);
nand I_42619 (I728122,I835298,I835301);
and I_42620 (I728139,I728122,I835304);
DFFARX1 I_42621 (I728139,I3563,I727805,I728165,);
nor I_42622 (I728173,I728165,I728032);
DFFARX1 I_42623 (I728173,I3563,I727805,I727773,);
nand I_42624 (I728204,I728165,I728074);
nand I_42625 (I727782,I728057,I728204);
not I_42626 (I728235,I728165);
nor I_42627 (I728252,I728235,I727975);
DFFARX1 I_42628 (I728252,I3563,I727805,I727794,);
nor I_42629 (I728283,I835310,I835301);
or I_42630 (I727785,I728032,I728283);
nor I_42631 (I727776,I728165,I728283);
or I_42632 (I727779,I727899,I728283);
DFFARX1 I_42633 (I728283,I3563,I727805,I727797,);
not I_42634 (I728383,I3570);
DFFARX1 I_42635 (I453963,I3563,I728383,I728409,);
not I_42636 (I728417,I728409);
nand I_42637 (I728434,I453954,I453972);
and I_42638 (I728451,I728434,I453975);
DFFARX1 I_42639 (I728451,I3563,I728383,I728477,);
not I_42640 (I728485,I453969);
DFFARX1 I_42641 (I453957,I3563,I728383,I728511,);
not I_42642 (I728519,I728511);
nor I_42643 (I728536,I728519,I728417);
and I_42644 (I728553,I728536,I453969);
nor I_42645 (I728570,I728519,I728485);
nor I_42646 (I728366,I728477,I728570);
DFFARX1 I_42647 (I453966,I3563,I728383,I728610,);
nor I_42648 (I728618,I728610,I728477);
not I_42649 (I728635,I728618);
not I_42650 (I728652,I728610);
nor I_42651 (I728669,I728652,I728553);
DFFARX1 I_42652 (I728669,I3563,I728383,I728369,);
nand I_42653 (I728700,I453981,I453978);
and I_42654 (I728717,I728700,I453960);
DFFARX1 I_42655 (I728717,I3563,I728383,I728743,);
nor I_42656 (I728751,I728743,I728610);
DFFARX1 I_42657 (I728751,I3563,I728383,I728351,);
nand I_42658 (I728782,I728743,I728652);
nand I_42659 (I728360,I728635,I728782);
not I_42660 (I728813,I728743);
nor I_42661 (I728830,I728813,I728553);
DFFARX1 I_42662 (I728830,I3563,I728383,I728372,);
nor I_42663 (I728861,I453954,I453978);
or I_42664 (I728363,I728610,I728861);
nor I_42665 (I728354,I728743,I728861);
or I_42666 (I728357,I728477,I728861);
DFFARX1 I_42667 (I728861,I3563,I728383,I728375,);
not I_42668 (I728961,I3570);
DFFARX1 I_42669 (I1389270,I3563,I728961,I728987,);
not I_42670 (I728995,I728987);
nand I_42671 (I729012,I1389255,I1389243);
and I_42672 (I729029,I729012,I1389258);
DFFARX1 I_42673 (I729029,I3563,I728961,I729055,);
not I_42674 (I729063,I1389243);
DFFARX1 I_42675 (I1389261,I3563,I728961,I729089,);
not I_42676 (I729097,I729089);
nor I_42677 (I729114,I729097,I728995);
and I_42678 (I729131,I729114,I1389243);
nor I_42679 (I729148,I729097,I729063);
nor I_42680 (I728944,I729055,I729148);
DFFARX1 I_42681 (I1389249,I3563,I728961,I729188,);
nor I_42682 (I729196,I729188,I729055);
not I_42683 (I729213,I729196);
not I_42684 (I729230,I729188);
nor I_42685 (I729247,I729230,I729131);
DFFARX1 I_42686 (I729247,I3563,I728961,I728947,);
nand I_42687 (I729278,I1389246,I1389252);
and I_42688 (I729295,I729278,I1389267);
DFFARX1 I_42689 (I729295,I3563,I728961,I729321,);
nor I_42690 (I729329,I729321,I729188);
DFFARX1 I_42691 (I729329,I3563,I728961,I728929,);
nand I_42692 (I729360,I729321,I729230);
nand I_42693 (I728938,I729213,I729360);
not I_42694 (I729391,I729321);
nor I_42695 (I729408,I729391,I729131);
DFFARX1 I_42696 (I729408,I3563,I728961,I728950,);
nor I_42697 (I729439,I1389264,I1389252);
or I_42698 (I728941,I729188,I729439);
nor I_42699 (I728932,I729321,I729439);
or I_42700 (I728935,I729055,I729439);
DFFARX1 I_42701 (I729439,I3563,I728961,I728953,);
not I_42702 (I729539,I3570);
DFFARX1 I_42703 (I1138409,I3563,I729539,I729565,);
not I_42704 (I729573,I729565);
nand I_42705 (I729590,I1138391,I1138403);
and I_42706 (I729607,I729590,I1138406);
DFFARX1 I_42707 (I729607,I3563,I729539,I729633,);
not I_42708 (I729641,I1138400);
DFFARX1 I_42709 (I1138397,I3563,I729539,I729667,);
not I_42710 (I729675,I729667);
nor I_42711 (I729692,I729675,I729573);
and I_42712 (I729709,I729692,I1138400);
nor I_42713 (I729726,I729675,I729641);
nor I_42714 (I729522,I729633,I729726);
DFFARX1 I_42715 (I1138415,I3563,I729539,I729766,);
nor I_42716 (I729774,I729766,I729633);
not I_42717 (I729791,I729774);
not I_42718 (I729808,I729766);
nor I_42719 (I729825,I729808,I729709);
DFFARX1 I_42720 (I729825,I3563,I729539,I729525,);
nand I_42721 (I729856,I1138394,I1138394);
and I_42722 (I729873,I729856,I1138391);
DFFARX1 I_42723 (I729873,I3563,I729539,I729899,);
nor I_42724 (I729907,I729899,I729766);
DFFARX1 I_42725 (I729907,I3563,I729539,I729507,);
nand I_42726 (I729938,I729899,I729808);
nand I_42727 (I729516,I729791,I729938);
not I_42728 (I729969,I729899);
nor I_42729 (I729986,I729969,I729709);
DFFARX1 I_42730 (I729986,I3563,I729539,I729528,);
nor I_42731 (I730017,I1138412,I1138394);
or I_42732 (I729519,I729766,I730017);
nor I_42733 (I729510,I729899,I730017);
or I_42734 (I729513,I729633,I730017);
DFFARX1 I_42735 (I730017,I3563,I729539,I729531,);
not I_42736 (I730117,I3570);
DFFARX1 I_42737 (I210123,I3563,I730117,I730143,);
not I_42738 (I730151,I730143);
nand I_42739 (I730168,I210126,I210147);
and I_42740 (I730185,I730168,I210135);
DFFARX1 I_42741 (I730185,I3563,I730117,I730211,);
not I_42742 (I730219,I210132);
DFFARX1 I_42743 (I210123,I3563,I730117,I730245,);
not I_42744 (I730253,I730245);
nor I_42745 (I730270,I730253,I730151);
and I_42746 (I730287,I730270,I210132);
nor I_42747 (I730304,I730253,I730219);
nor I_42748 (I730100,I730211,I730304);
DFFARX1 I_42749 (I210141,I3563,I730117,I730344,);
nor I_42750 (I730352,I730344,I730211);
not I_42751 (I730369,I730352);
not I_42752 (I730386,I730344);
nor I_42753 (I730403,I730386,I730287);
DFFARX1 I_42754 (I730403,I3563,I730117,I730103,);
nand I_42755 (I730434,I210126,I210129);
and I_42756 (I730451,I730434,I210138);
DFFARX1 I_42757 (I730451,I3563,I730117,I730477,);
nor I_42758 (I730485,I730477,I730344);
DFFARX1 I_42759 (I730485,I3563,I730117,I730085,);
nand I_42760 (I730516,I730477,I730386);
nand I_42761 (I730094,I730369,I730516);
not I_42762 (I730547,I730477);
nor I_42763 (I730564,I730547,I730287);
DFFARX1 I_42764 (I730564,I3563,I730117,I730106,);
nor I_42765 (I730595,I210144,I210129);
or I_42766 (I730097,I730344,I730595);
nor I_42767 (I730088,I730477,I730595);
or I_42768 (I730091,I730211,I730595);
DFFARX1 I_42769 (I730595,I3563,I730117,I730109,);
not I_42770 (I730695,I3570);
DFFARX1 I_42771 (I882216,I3563,I730695,I730721,);
not I_42772 (I730729,I730721);
nand I_42773 (I730746,I882204,I882222);
and I_42774 (I730763,I730746,I882219);
DFFARX1 I_42775 (I730763,I3563,I730695,I730789,);
not I_42776 (I730797,I882210);
DFFARX1 I_42777 (I882207,I3563,I730695,I730823,);
not I_42778 (I730831,I730823);
nor I_42779 (I730848,I730831,I730729);
and I_42780 (I730865,I730848,I882210);
nor I_42781 (I730882,I730831,I730797);
nor I_42782 (I730678,I730789,I730882);
DFFARX1 I_42783 (I882201,I3563,I730695,I730922,);
nor I_42784 (I730930,I730922,I730789);
not I_42785 (I730947,I730930);
not I_42786 (I730964,I730922);
nor I_42787 (I730981,I730964,I730865);
DFFARX1 I_42788 (I730981,I3563,I730695,I730681,);
nand I_42789 (I731012,I882201,I882204);
and I_42790 (I731029,I731012,I882207);
DFFARX1 I_42791 (I731029,I3563,I730695,I731055,);
nor I_42792 (I731063,I731055,I730922);
DFFARX1 I_42793 (I731063,I3563,I730695,I730663,);
nand I_42794 (I731094,I731055,I730964);
nand I_42795 (I730672,I730947,I731094);
not I_42796 (I731125,I731055);
nor I_42797 (I731142,I731125,I730865);
DFFARX1 I_42798 (I731142,I3563,I730695,I730684,);
nor I_42799 (I731173,I882213,I882204);
or I_42800 (I730675,I730922,I731173);
nor I_42801 (I730666,I731055,I731173);
or I_42802 (I730669,I730789,I731173);
DFFARX1 I_42803 (I731173,I3563,I730695,I730687,);
not I_42804 (I731273,I3570);
DFFARX1 I_42805 (I1301625,I3563,I731273,I731299,);
not I_42806 (I731307,I731299);
nand I_42807 (I731324,I1301649,I1301631);
and I_42808 (I731341,I731324,I1301637);
DFFARX1 I_42809 (I731341,I3563,I731273,I731367,);
not I_42810 (I731375,I1301643);
DFFARX1 I_42811 (I1301628,I3563,I731273,I731401,);
not I_42812 (I731409,I731401);
nor I_42813 (I731426,I731409,I731307);
and I_42814 (I731443,I731426,I1301643);
nor I_42815 (I731460,I731409,I731375);
nor I_42816 (I731256,I731367,I731460);
DFFARX1 I_42817 (I1301640,I3563,I731273,I731500,);
nor I_42818 (I731508,I731500,I731367);
not I_42819 (I731525,I731508);
not I_42820 (I731542,I731500);
nor I_42821 (I731559,I731542,I731443);
DFFARX1 I_42822 (I731559,I3563,I731273,I731259,);
nand I_42823 (I731590,I1301646,I1301634);
and I_42824 (I731607,I731590,I1301628);
DFFARX1 I_42825 (I731607,I3563,I731273,I731633,);
nor I_42826 (I731641,I731633,I731500);
DFFARX1 I_42827 (I731641,I3563,I731273,I731241,);
nand I_42828 (I731672,I731633,I731542);
nand I_42829 (I731250,I731525,I731672);
not I_42830 (I731703,I731633);
nor I_42831 (I731720,I731703,I731443);
DFFARX1 I_42832 (I731720,I3563,I731273,I731262,);
nor I_42833 (I731751,I1301625,I1301634);
or I_42834 (I731253,I731500,I731751);
nor I_42835 (I731244,I731633,I731751);
or I_42836 (I731247,I731367,I731751);
DFFARX1 I_42837 (I731751,I3563,I731273,I731265,);
not I_42838 (I731851,I3570);
DFFARX1 I_42839 (I1204301,I3563,I731851,I731877,);
not I_42840 (I731885,I731877);
nand I_42841 (I731902,I1204283,I1204295);
and I_42842 (I731919,I731902,I1204298);
DFFARX1 I_42843 (I731919,I3563,I731851,I731945,);
not I_42844 (I731953,I1204292);
DFFARX1 I_42845 (I1204289,I3563,I731851,I731979,);
not I_42846 (I731987,I731979);
nor I_42847 (I732004,I731987,I731885);
and I_42848 (I732021,I732004,I1204292);
nor I_42849 (I732038,I731987,I731953);
nor I_42850 (I731834,I731945,I732038);
DFFARX1 I_42851 (I1204307,I3563,I731851,I732078,);
nor I_42852 (I732086,I732078,I731945);
not I_42853 (I732103,I732086);
not I_42854 (I732120,I732078);
nor I_42855 (I732137,I732120,I732021);
DFFARX1 I_42856 (I732137,I3563,I731851,I731837,);
nand I_42857 (I732168,I1204286,I1204286);
and I_42858 (I732185,I732168,I1204283);
DFFARX1 I_42859 (I732185,I3563,I731851,I732211,);
nor I_42860 (I732219,I732211,I732078);
DFFARX1 I_42861 (I732219,I3563,I731851,I731819,);
nand I_42862 (I732250,I732211,I732120);
nand I_42863 (I731828,I732103,I732250);
not I_42864 (I732281,I732211);
nor I_42865 (I732298,I732281,I732021);
DFFARX1 I_42866 (I732298,I3563,I731851,I731840,);
nor I_42867 (I732329,I1204304,I1204286);
or I_42868 (I731831,I732078,I732329);
nor I_42869 (I731822,I732211,I732329);
or I_42870 (I731825,I731945,I732329);
DFFARX1 I_42871 (I732329,I3563,I731851,I731843,);
not I_42872 (I732429,I3570);
DFFARX1 I_42873 (I531661,I3563,I732429,I732455,);
not I_42874 (I732463,I732455);
nand I_42875 (I732480,I531676,I531661);
and I_42876 (I732497,I732480,I531664);
DFFARX1 I_42877 (I732497,I3563,I732429,I732523,);
not I_42878 (I732531,I531664);
DFFARX1 I_42879 (I531673,I3563,I732429,I732557,);
not I_42880 (I732565,I732557);
nor I_42881 (I732582,I732565,I732463);
and I_42882 (I732599,I732582,I531664);
nor I_42883 (I732616,I732565,I732531);
nor I_42884 (I732412,I732523,I732616);
DFFARX1 I_42885 (I531667,I3563,I732429,I732656,);
nor I_42886 (I732664,I732656,I732523);
not I_42887 (I732681,I732664);
not I_42888 (I732698,I732656);
nor I_42889 (I732715,I732698,I732599);
DFFARX1 I_42890 (I732715,I3563,I732429,I732415,);
nand I_42891 (I732746,I531670,I531679);
and I_42892 (I732763,I732746,I531685);
DFFARX1 I_42893 (I732763,I3563,I732429,I732789,);
nor I_42894 (I732797,I732789,I732656);
DFFARX1 I_42895 (I732797,I3563,I732429,I732397,);
nand I_42896 (I732828,I732789,I732698);
nand I_42897 (I732406,I732681,I732828);
not I_42898 (I732859,I732789);
nor I_42899 (I732876,I732859,I732599);
DFFARX1 I_42900 (I732876,I3563,I732429,I732418,);
nor I_42901 (I732907,I531682,I531679);
or I_42902 (I732409,I732656,I732907);
nor I_42903 (I732400,I732789,I732907);
or I_42904 (I732403,I732523,I732907);
DFFARX1 I_42905 (I732907,I3563,I732429,I732421,);
not I_42906 (I733007,I3570);
DFFARX1 I_42907 (I70879,I3563,I733007,I733033,);
not I_42908 (I733041,I733033);
nand I_42909 (I733058,I70888,I70897);
and I_42910 (I733075,I733058,I70876);
DFFARX1 I_42911 (I733075,I3563,I733007,I733101,);
not I_42912 (I733109,I70879);
DFFARX1 I_42913 (I70894,I3563,I733007,I733135,);
not I_42914 (I733143,I733135);
nor I_42915 (I733160,I733143,I733041);
and I_42916 (I733177,I733160,I70879);
nor I_42917 (I733194,I733143,I733109);
nor I_42918 (I732990,I733101,I733194);
DFFARX1 I_42919 (I70885,I3563,I733007,I733234,);
nor I_42920 (I733242,I733234,I733101);
not I_42921 (I733259,I733242);
not I_42922 (I733276,I733234);
nor I_42923 (I733293,I733276,I733177);
DFFARX1 I_42924 (I733293,I3563,I733007,I732993,);
nand I_42925 (I733324,I70900,I70876);
and I_42926 (I733341,I733324,I70882);
DFFARX1 I_42927 (I733341,I3563,I733007,I733367,);
nor I_42928 (I733375,I733367,I733234);
DFFARX1 I_42929 (I733375,I3563,I733007,I732975,);
nand I_42930 (I733406,I733367,I733276);
nand I_42931 (I732984,I733259,I733406);
not I_42932 (I733437,I733367);
nor I_42933 (I733454,I733437,I733177);
DFFARX1 I_42934 (I733454,I3563,I733007,I732996,);
nor I_42935 (I733485,I70891,I70876);
or I_42936 (I732987,I733234,I733485);
nor I_42937 (I732978,I733367,I733485);
or I_42938 (I732981,I733101,I733485);
DFFARX1 I_42939 (I733485,I3563,I733007,I732999,);
not I_42940 (I733585,I3570);
DFFARX1 I_42941 (I1050592,I3563,I733585,I733611,);
not I_42942 (I733619,I733611);
nand I_42943 (I733636,I1050589,I1050607);
and I_42944 (I733653,I733636,I1050604);
DFFARX1 I_42945 (I733653,I3563,I733585,I733679,);
not I_42946 (I733687,I1050586);
DFFARX1 I_42947 (I1050589,I3563,I733585,I733713,);
not I_42948 (I733721,I733713);
nor I_42949 (I733738,I733721,I733619);
and I_42950 (I733755,I733738,I1050586);
nor I_42951 (I733772,I733721,I733687);
nor I_42952 (I733568,I733679,I733772);
DFFARX1 I_42953 (I1050598,I3563,I733585,I733812,);
nor I_42954 (I733820,I733812,I733679);
not I_42955 (I733837,I733820);
not I_42956 (I733854,I733812);
nor I_42957 (I733871,I733854,I733755);
DFFARX1 I_42958 (I733871,I3563,I733585,I733571,);
nand I_42959 (I733902,I1050601,I1050586);
and I_42960 (I733919,I733902,I1050592);
DFFARX1 I_42961 (I733919,I3563,I733585,I733945,);
nor I_42962 (I733953,I733945,I733812);
DFFARX1 I_42963 (I733953,I3563,I733585,I733553,);
nand I_42964 (I733984,I733945,I733854);
nand I_42965 (I733562,I733837,I733984);
not I_42966 (I734015,I733945);
nor I_42967 (I734032,I734015,I733755);
DFFARX1 I_42968 (I734032,I3563,I733585,I733574,);
nor I_42969 (I734063,I1050595,I1050586);
or I_42970 (I733565,I733812,I734063);
nor I_42971 (I733556,I733945,I734063);
or I_42972 (I733559,I733679,I734063);
DFFARX1 I_42973 (I734063,I3563,I733585,I733577,);
not I_42974 (I734163,I3570);
DFFARX1 I_42975 (I552486,I3563,I734163,I734189,);
not I_42976 (I734197,I734189);
nand I_42977 (I734214,I552501,I552486);
and I_42978 (I734231,I734214,I552489);
DFFARX1 I_42979 (I734231,I3563,I734163,I734257,);
not I_42980 (I734265,I552489);
DFFARX1 I_42981 (I552498,I3563,I734163,I734291,);
not I_42982 (I734299,I734291);
nor I_42983 (I734316,I734299,I734197);
and I_42984 (I734333,I734316,I552489);
nor I_42985 (I734350,I734299,I734265);
nor I_42986 (I734146,I734257,I734350);
DFFARX1 I_42987 (I552492,I3563,I734163,I734390,);
nor I_42988 (I734398,I734390,I734257);
not I_42989 (I734415,I734398);
not I_42990 (I734432,I734390);
nor I_42991 (I734449,I734432,I734333);
DFFARX1 I_42992 (I734449,I3563,I734163,I734149,);
nand I_42993 (I734480,I552495,I552504);
and I_42994 (I734497,I734480,I552510);
DFFARX1 I_42995 (I734497,I3563,I734163,I734523,);
nor I_42996 (I734531,I734523,I734390);
DFFARX1 I_42997 (I734531,I3563,I734163,I734131,);
nand I_42998 (I734562,I734523,I734432);
nand I_42999 (I734140,I734415,I734562);
not I_43000 (I734593,I734523);
nor I_43001 (I734610,I734593,I734333);
DFFARX1 I_43002 (I734610,I3563,I734163,I734152,);
nor I_43003 (I734641,I552507,I552504);
or I_43004 (I734143,I734390,I734641);
nor I_43005 (I734134,I734523,I734641);
or I_43006 (I734137,I734257,I734641);
DFFARX1 I_43007 (I734641,I3563,I734163,I734155,);
not I_43008 (I734741,I3570);
DFFARX1 I_43009 (I486059,I3563,I734741,I734767,);
not I_43010 (I734775,I734767);
nand I_43011 (I734792,I486050,I486068);
and I_43012 (I734809,I734792,I486071);
DFFARX1 I_43013 (I734809,I3563,I734741,I734835,);
not I_43014 (I734843,I486065);
DFFARX1 I_43015 (I486053,I3563,I734741,I734869,);
not I_43016 (I734877,I734869);
nor I_43017 (I734894,I734877,I734775);
and I_43018 (I734911,I734894,I486065);
nor I_43019 (I734928,I734877,I734843);
nor I_43020 (I734724,I734835,I734928);
DFFARX1 I_43021 (I486062,I3563,I734741,I734968,);
nor I_43022 (I734976,I734968,I734835);
not I_43023 (I734993,I734976);
not I_43024 (I735010,I734968);
nor I_43025 (I735027,I735010,I734911);
DFFARX1 I_43026 (I735027,I3563,I734741,I734727,);
nand I_43027 (I735058,I486077,I486074);
and I_43028 (I735075,I735058,I486056);
DFFARX1 I_43029 (I735075,I3563,I734741,I735101,);
nor I_43030 (I735109,I735101,I734968);
DFFARX1 I_43031 (I735109,I3563,I734741,I734709,);
nand I_43032 (I735140,I735101,I735010);
nand I_43033 (I734718,I734993,I735140);
not I_43034 (I735171,I735101);
nor I_43035 (I735188,I735171,I734911);
DFFARX1 I_43036 (I735188,I3563,I734741,I734730,);
nor I_43037 (I735219,I486050,I486074);
or I_43038 (I734721,I734968,I735219);
nor I_43039 (I734712,I735101,I735219);
or I_43040 (I734715,I734835,I735219);
DFFARX1 I_43041 (I735219,I3563,I734741,I734733,);
not I_43042 (I735319,I3570);
DFFARX1 I_43043 (I320171,I3563,I735319,I735345,);
not I_43044 (I735353,I735345);
nand I_43045 (I735370,I320174,I320150);
and I_43046 (I735387,I735370,I320147);
DFFARX1 I_43047 (I735387,I3563,I735319,I735413,);
not I_43048 (I735421,I320153);
DFFARX1 I_43049 (I320147,I3563,I735319,I735447,);
not I_43050 (I735455,I735447);
nor I_43051 (I735472,I735455,I735353);
and I_43052 (I735489,I735472,I320153);
nor I_43053 (I735506,I735455,I735421);
nor I_43054 (I735302,I735413,I735506);
DFFARX1 I_43055 (I320156,I3563,I735319,I735546,);
nor I_43056 (I735554,I735546,I735413);
not I_43057 (I735571,I735554);
not I_43058 (I735588,I735546);
nor I_43059 (I735605,I735588,I735489);
DFFARX1 I_43060 (I735605,I3563,I735319,I735305,);
nand I_43061 (I735636,I320159,I320168);
and I_43062 (I735653,I735636,I320165);
DFFARX1 I_43063 (I735653,I3563,I735319,I735679,);
nor I_43064 (I735687,I735679,I735546);
DFFARX1 I_43065 (I735687,I3563,I735319,I735287,);
nand I_43066 (I735718,I735679,I735588);
nand I_43067 (I735296,I735571,I735718);
not I_43068 (I735749,I735679);
nor I_43069 (I735766,I735749,I735489);
DFFARX1 I_43070 (I735766,I3563,I735319,I735308,);
nor I_43071 (I735797,I320162,I320168);
or I_43072 (I735299,I735546,I735797);
nor I_43073 (I735290,I735679,I735797);
or I_43074 (I735293,I735413,I735797);
DFFARX1 I_43075 (I735797,I3563,I735319,I735311,);
not I_43076 (I735897,I3570);
DFFARX1 I_43077 (I1145345,I3563,I735897,I735923,);
not I_43078 (I735931,I735923);
nand I_43079 (I735948,I1145327,I1145339);
and I_43080 (I735965,I735948,I1145342);
DFFARX1 I_43081 (I735965,I3563,I735897,I735991,);
not I_43082 (I735999,I1145336);
DFFARX1 I_43083 (I1145333,I3563,I735897,I736025,);
not I_43084 (I736033,I736025);
nor I_43085 (I736050,I736033,I735931);
and I_43086 (I736067,I736050,I1145336);
nor I_43087 (I736084,I736033,I735999);
nor I_43088 (I735880,I735991,I736084);
DFFARX1 I_43089 (I1145351,I3563,I735897,I736124,);
nor I_43090 (I736132,I736124,I735991);
not I_43091 (I736149,I736132);
not I_43092 (I736166,I736124);
nor I_43093 (I736183,I736166,I736067);
DFFARX1 I_43094 (I736183,I3563,I735897,I735883,);
nand I_43095 (I736214,I1145330,I1145330);
and I_43096 (I736231,I736214,I1145327);
DFFARX1 I_43097 (I736231,I3563,I735897,I736257,);
nor I_43098 (I736265,I736257,I736124);
DFFARX1 I_43099 (I736265,I3563,I735897,I735865,);
nand I_43100 (I736296,I736257,I736166);
nand I_43101 (I735874,I736149,I736296);
not I_43102 (I736327,I736257);
nor I_43103 (I736344,I736327,I736067);
DFFARX1 I_43104 (I736344,I3563,I735897,I735886,);
nor I_43105 (I736375,I1145348,I1145330);
or I_43106 (I735877,I736124,I736375);
nor I_43107 (I735868,I736257,I736375);
or I_43108 (I735871,I735991,I736375);
DFFARX1 I_43109 (I736375,I3563,I735897,I735889,);
not I_43110 (I736475,I3570);
DFFARX1 I_43111 (I920067,I3563,I736475,I736501,);
not I_43112 (I736509,I736501);
nand I_43113 (I736526,I920043,I920058);
and I_43114 (I736543,I736526,I920070);
DFFARX1 I_43115 (I736543,I3563,I736475,I736569,);
not I_43116 (I736577,I920055);
DFFARX1 I_43117 (I920046,I3563,I736475,I736603,);
not I_43118 (I736611,I736603);
nor I_43119 (I736628,I736611,I736509);
and I_43120 (I736645,I736628,I920055);
nor I_43121 (I736662,I736611,I736577);
nor I_43122 (I736458,I736569,I736662);
DFFARX1 I_43123 (I920043,I3563,I736475,I736702,);
nor I_43124 (I736710,I736702,I736569);
not I_43125 (I736727,I736710);
not I_43126 (I736744,I736702);
nor I_43127 (I736761,I736744,I736645);
DFFARX1 I_43128 (I736761,I3563,I736475,I736461,);
nand I_43129 (I736792,I920061,I920052);
and I_43130 (I736809,I736792,I920064);
DFFARX1 I_43131 (I736809,I3563,I736475,I736835,);
nor I_43132 (I736843,I736835,I736702);
DFFARX1 I_43133 (I736843,I3563,I736475,I736443,);
nand I_43134 (I736874,I736835,I736744);
nand I_43135 (I736452,I736727,I736874);
not I_43136 (I736905,I736835);
nor I_43137 (I736922,I736905,I736645);
DFFARX1 I_43138 (I736922,I3563,I736475,I736464,);
nor I_43139 (I736953,I920049,I920052);
or I_43140 (I736455,I736702,I736953);
nor I_43141 (I736446,I736835,I736953);
or I_43142 (I736449,I736569,I736953);
DFFARX1 I_43143 (I736953,I3563,I736475,I736467,);
not I_43144 (I737053,I3570);
DFFARX1 I_43145 (I1201411,I3563,I737053,I737079,);
not I_43146 (I737087,I737079);
nand I_43147 (I737104,I1201393,I1201405);
and I_43148 (I737121,I737104,I1201408);
DFFARX1 I_43149 (I737121,I3563,I737053,I737147,);
not I_43150 (I737155,I1201402);
DFFARX1 I_43151 (I1201399,I3563,I737053,I737181,);
not I_43152 (I737189,I737181);
nor I_43153 (I737206,I737189,I737087);
and I_43154 (I737223,I737206,I1201402);
nor I_43155 (I737240,I737189,I737155);
nor I_43156 (I737036,I737147,I737240);
DFFARX1 I_43157 (I1201417,I3563,I737053,I737280,);
nor I_43158 (I737288,I737280,I737147);
not I_43159 (I737305,I737288);
not I_43160 (I737322,I737280);
nor I_43161 (I737339,I737322,I737223);
DFFARX1 I_43162 (I737339,I3563,I737053,I737039,);
nand I_43163 (I737370,I1201396,I1201396);
and I_43164 (I737387,I737370,I1201393);
DFFARX1 I_43165 (I737387,I3563,I737053,I737413,);
nor I_43166 (I737421,I737413,I737280);
DFFARX1 I_43167 (I737421,I3563,I737053,I737021,);
nand I_43168 (I737452,I737413,I737322);
nand I_43169 (I737030,I737305,I737452);
not I_43170 (I737483,I737413);
nor I_43171 (I737500,I737483,I737223);
DFFARX1 I_43172 (I737500,I3563,I737053,I737042,);
nor I_43173 (I737531,I1201414,I1201396);
or I_43174 (I737033,I737280,I737531);
nor I_43175 (I737024,I737413,I737531);
or I_43176 (I737027,I737147,I737531);
DFFARX1 I_43177 (I737531,I3563,I737053,I737045,);
not I_43178 (I737631,I3570);
DFFARX1 I_43179 (I35052,I3563,I737631,I737657,);
not I_43180 (I737665,I737657);
nand I_43181 (I737682,I35049,I35040);
and I_43182 (I737699,I737682,I35040);
DFFARX1 I_43183 (I737699,I3563,I737631,I737725,);
not I_43184 (I737733,I35043);
DFFARX1 I_43185 (I35058,I3563,I737631,I737759,);
not I_43186 (I737767,I737759);
nor I_43187 (I737784,I737767,I737665);
and I_43188 (I737801,I737784,I35043);
nor I_43189 (I737818,I737767,I737733);
nor I_43190 (I737614,I737725,I737818);
DFFARX1 I_43191 (I35043,I3563,I737631,I737858,);
nor I_43192 (I737866,I737858,I737725);
not I_43193 (I737883,I737866);
not I_43194 (I737900,I737858);
nor I_43195 (I737917,I737900,I737801);
DFFARX1 I_43196 (I737917,I3563,I737631,I737617,);
nand I_43197 (I737948,I35061,I35046);
and I_43198 (I737965,I737948,I35064);
DFFARX1 I_43199 (I737965,I3563,I737631,I737991,);
nor I_43200 (I737999,I737991,I737858);
DFFARX1 I_43201 (I737999,I3563,I737631,I737599,);
nand I_43202 (I738030,I737991,I737900);
nand I_43203 (I737608,I737883,I738030);
not I_43204 (I738061,I737991);
nor I_43205 (I738078,I738061,I737801);
DFFARX1 I_43206 (I738078,I3563,I737631,I737620,);
nor I_43207 (I738109,I35055,I35046);
or I_43208 (I737611,I737858,I738109);
nor I_43209 (I737602,I737991,I738109);
or I_43210 (I737605,I737725,I738109);
DFFARX1 I_43211 (I738109,I3563,I737631,I737623,);
not I_43212 (I738209,I3570);
DFFARX1 I_43213 (I648009,I3563,I738209,I738235,);
not I_43214 (I738243,I738235);
nand I_43215 (I738260,I648018,I648027);
and I_43216 (I738277,I738260,I648033);
DFFARX1 I_43217 (I738277,I3563,I738209,I738303,);
not I_43218 (I738311,I648030);
DFFARX1 I_43219 (I648015,I3563,I738209,I738337,);
not I_43220 (I738345,I738337);
nor I_43221 (I738362,I738345,I738243);
and I_43222 (I738379,I738362,I648030);
nor I_43223 (I738396,I738345,I738311);
nor I_43224 (I738192,I738303,I738396);
DFFARX1 I_43225 (I648024,I3563,I738209,I738436,);
nor I_43226 (I738444,I738436,I738303);
not I_43227 (I738461,I738444);
not I_43228 (I738478,I738436);
nor I_43229 (I738495,I738478,I738379);
DFFARX1 I_43230 (I738495,I3563,I738209,I738195,);
nand I_43231 (I738526,I648021,I648012);
and I_43232 (I738543,I738526,I648009);
DFFARX1 I_43233 (I738543,I3563,I738209,I738569,);
nor I_43234 (I738577,I738569,I738436);
DFFARX1 I_43235 (I738577,I3563,I738209,I738177,);
nand I_43236 (I738608,I738569,I738478);
nand I_43237 (I738186,I738461,I738608);
not I_43238 (I738639,I738569);
nor I_43239 (I738656,I738639,I738379);
DFFARX1 I_43240 (I738656,I3563,I738209,I738198,);
nor I_43241 (I738687,I648012,I648012);
or I_43242 (I738189,I738436,I738687);
nor I_43243 (I738180,I738569,I738687);
or I_43244 (I738183,I738303,I738687);
DFFARX1 I_43245 (I738687,I3563,I738209,I738201,);
not I_43246 (I738787,I3570);
DFFARX1 I_43247 (I1370230,I3563,I738787,I738813,);
not I_43248 (I738821,I738813);
nand I_43249 (I738838,I1370215,I1370203);
and I_43250 (I738855,I738838,I1370218);
DFFARX1 I_43251 (I738855,I3563,I738787,I738881,);
not I_43252 (I738889,I1370203);
DFFARX1 I_43253 (I1370221,I3563,I738787,I738915,);
not I_43254 (I738923,I738915);
nor I_43255 (I738940,I738923,I738821);
and I_43256 (I738957,I738940,I1370203);
nor I_43257 (I738974,I738923,I738889);
nor I_43258 (I738770,I738881,I738974);
DFFARX1 I_43259 (I1370209,I3563,I738787,I739014,);
nor I_43260 (I739022,I739014,I738881);
not I_43261 (I739039,I739022);
not I_43262 (I739056,I739014);
nor I_43263 (I739073,I739056,I738957);
DFFARX1 I_43264 (I739073,I3563,I738787,I738773,);
nand I_43265 (I739104,I1370206,I1370212);
and I_43266 (I739121,I739104,I1370227);
DFFARX1 I_43267 (I739121,I3563,I738787,I739147,);
nor I_43268 (I739155,I739147,I739014);
DFFARX1 I_43269 (I739155,I3563,I738787,I738755,);
nand I_43270 (I739186,I739147,I739056);
nand I_43271 (I738764,I739039,I739186);
not I_43272 (I739217,I739147);
nor I_43273 (I739234,I739217,I738957);
DFFARX1 I_43274 (I739234,I3563,I738787,I738776,);
nor I_43275 (I739265,I1370224,I1370212);
or I_43276 (I738767,I739014,I739265);
nor I_43277 (I738758,I739147,I739265);
or I_43278 (I738761,I738881,I739265);
DFFARX1 I_43279 (I739265,I3563,I738787,I738779,);
not I_43280 (I739365,I3570);
DFFARX1 I_43281 (I1188117,I3563,I739365,I739391,);
not I_43282 (I739399,I739391);
nand I_43283 (I739416,I1188099,I1188111);
and I_43284 (I739433,I739416,I1188114);
DFFARX1 I_43285 (I739433,I3563,I739365,I739459,);
not I_43286 (I739467,I1188108);
DFFARX1 I_43287 (I1188105,I3563,I739365,I739493,);
not I_43288 (I739501,I739493);
nor I_43289 (I739518,I739501,I739399);
and I_43290 (I739535,I739518,I1188108);
nor I_43291 (I739552,I739501,I739467);
nor I_43292 (I739348,I739459,I739552);
DFFARX1 I_43293 (I1188123,I3563,I739365,I739592,);
nor I_43294 (I739600,I739592,I739459);
not I_43295 (I739617,I739600);
not I_43296 (I739634,I739592);
nor I_43297 (I739651,I739634,I739535);
DFFARX1 I_43298 (I739651,I3563,I739365,I739351,);
nand I_43299 (I739682,I1188102,I1188102);
and I_43300 (I739699,I739682,I1188099);
DFFARX1 I_43301 (I739699,I3563,I739365,I739725,);
nor I_43302 (I739733,I739725,I739592);
DFFARX1 I_43303 (I739733,I3563,I739365,I739333,);
nand I_43304 (I739764,I739725,I739634);
nand I_43305 (I739342,I739617,I739764);
not I_43306 (I739795,I739725);
nor I_43307 (I739812,I739795,I739535);
DFFARX1 I_43308 (I739812,I3563,I739365,I739354,);
nor I_43309 (I739843,I1188120,I1188102);
or I_43310 (I739345,I739592,I739843);
nor I_43311 (I739336,I739725,I739843);
or I_43312 (I739339,I739459,I739843);
DFFARX1 I_43313 (I739843,I3563,I739365,I739357,);
not I_43314 (I739943,I3570);
DFFARX1 I_43315 (I554271,I3563,I739943,I739969,);
not I_43316 (I739977,I739969);
nand I_43317 (I739994,I554286,I554271);
and I_43318 (I740011,I739994,I554274);
DFFARX1 I_43319 (I740011,I3563,I739943,I740037,);
not I_43320 (I740045,I554274);
DFFARX1 I_43321 (I554283,I3563,I739943,I740071,);
not I_43322 (I740079,I740071);
nor I_43323 (I740096,I740079,I739977);
and I_43324 (I740113,I740096,I554274);
nor I_43325 (I740130,I740079,I740045);
nor I_43326 (I739926,I740037,I740130);
DFFARX1 I_43327 (I554277,I3563,I739943,I740170,);
nor I_43328 (I740178,I740170,I740037);
not I_43329 (I740195,I740178);
not I_43330 (I740212,I740170);
nor I_43331 (I740229,I740212,I740113);
DFFARX1 I_43332 (I740229,I3563,I739943,I739929,);
nand I_43333 (I740260,I554280,I554289);
and I_43334 (I740277,I740260,I554295);
DFFARX1 I_43335 (I740277,I3563,I739943,I740303,);
nor I_43336 (I740311,I740303,I740170);
DFFARX1 I_43337 (I740311,I3563,I739943,I739911,);
nand I_43338 (I740342,I740303,I740212);
nand I_43339 (I739920,I740195,I740342);
not I_43340 (I740373,I740303);
nor I_43341 (I740390,I740373,I740113);
DFFARX1 I_43342 (I740390,I3563,I739943,I739932,);
nor I_43343 (I740421,I554292,I554289);
or I_43344 (I739923,I740170,I740421);
nor I_43345 (I739914,I740303,I740421);
or I_43346 (I739917,I740037,I740421);
DFFARX1 I_43347 (I740421,I3563,I739943,I739935,);
not I_43348 (I740521,I3570);
DFFARX1 I_43349 (I80892,I3563,I740521,I740547,);
not I_43350 (I740555,I740547);
nand I_43351 (I740572,I80901,I80910);
and I_43352 (I740589,I740572,I80889);
DFFARX1 I_43353 (I740589,I3563,I740521,I740615,);
not I_43354 (I740623,I80892);
DFFARX1 I_43355 (I80907,I3563,I740521,I740649,);
not I_43356 (I740657,I740649);
nor I_43357 (I740674,I740657,I740555);
and I_43358 (I740691,I740674,I80892);
nor I_43359 (I740708,I740657,I740623);
nor I_43360 (I740504,I740615,I740708);
DFFARX1 I_43361 (I80898,I3563,I740521,I740748,);
nor I_43362 (I740756,I740748,I740615);
not I_43363 (I740773,I740756);
not I_43364 (I740790,I740748);
nor I_43365 (I740807,I740790,I740691);
DFFARX1 I_43366 (I740807,I3563,I740521,I740507,);
nand I_43367 (I740838,I80913,I80889);
and I_43368 (I740855,I740838,I80895);
DFFARX1 I_43369 (I740855,I3563,I740521,I740881,);
nor I_43370 (I740889,I740881,I740748);
DFFARX1 I_43371 (I740889,I3563,I740521,I740489,);
nand I_43372 (I740920,I740881,I740790);
nand I_43373 (I740498,I740773,I740920);
not I_43374 (I740951,I740881);
nor I_43375 (I740968,I740951,I740691);
DFFARX1 I_43376 (I740968,I3563,I740521,I740510,);
nor I_43377 (I740999,I80904,I80889);
or I_43378 (I740501,I740748,I740999);
nor I_43379 (I740492,I740881,I740999);
or I_43380 (I740495,I740615,I740999);
DFFARX1 I_43381 (I740999,I3563,I740521,I740513,);
not I_43382 (I741099,I3570);
DFFARX1 I_43383 (I284498,I3563,I741099,I741125,);
not I_43384 (I741133,I741125);
nand I_43385 (I741150,I284501,I284522);
and I_43386 (I741167,I741150,I284510);
DFFARX1 I_43387 (I741167,I3563,I741099,I741193,);
not I_43388 (I741201,I284507);
DFFARX1 I_43389 (I284498,I3563,I741099,I741227,);
not I_43390 (I741235,I741227);
nor I_43391 (I741252,I741235,I741133);
and I_43392 (I741269,I741252,I284507);
nor I_43393 (I741286,I741235,I741201);
nor I_43394 (I741082,I741193,I741286);
DFFARX1 I_43395 (I284516,I3563,I741099,I741326,);
nor I_43396 (I741334,I741326,I741193);
not I_43397 (I741351,I741334);
not I_43398 (I741368,I741326);
nor I_43399 (I741385,I741368,I741269);
DFFARX1 I_43400 (I741385,I3563,I741099,I741085,);
nand I_43401 (I741416,I284501,I284504);
and I_43402 (I741433,I741416,I284513);
DFFARX1 I_43403 (I741433,I3563,I741099,I741459,);
nor I_43404 (I741467,I741459,I741326);
DFFARX1 I_43405 (I741467,I3563,I741099,I741067,);
nand I_43406 (I741498,I741459,I741368);
nand I_43407 (I741076,I741351,I741498);
not I_43408 (I741529,I741459);
nor I_43409 (I741546,I741529,I741269);
DFFARX1 I_43410 (I741546,I3563,I741099,I741088,);
nor I_43411 (I741577,I284519,I284504);
or I_43412 (I741079,I741326,I741577);
nor I_43413 (I741070,I741459,I741577);
or I_43414 (I741073,I741193,I741577);
DFFARX1 I_43415 (I741577,I3563,I741099,I741091,);
not I_43416 (I741677,I3570);
DFFARX1 I_43417 (I993065,I3563,I741677,I741703,);
not I_43418 (I741711,I741703);
nand I_43419 (I741728,I993041,I993056);
and I_43420 (I741745,I741728,I993068);
DFFARX1 I_43421 (I741745,I3563,I741677,I741771,);
not I_43422 (I741779,I993053);
DFFARX1 I_43423 (I993044,I3563,I741677,I741805,);
not I_43424 (I741813,I741805);
nor I_43425 (I741830,I741813,I741711);
and I_43426 (I741847,I741830,I993053);
nor I_43427 (I741864,I741813,I741779);
nor I_43428 (I741660,I741771,I741864);
DFFARX1 I_43429 (I993041,I3563,I741677,I741904,);
nor I_43430 (I741912,I741904,I741771);
not I_43431 (I741929,I741912);
not I_43432 (I741946,I741904);
nor I_43433 (I741963,I741946,I741847);
DFFARX1 I_43434 (I741963,I3563,I741677,I741663,);
nand I_43435 (I741994,I993059,I993050);
and I_43436 (I742011,I741994,I993062);
DFFARX1 I_43437 (I742011,I3563,I741677,I742037,);
nor I_43438 (I742045,I742037,I741904);
DFFARX1 I_43439 (I742045,I3563,I741677,I741645,);
nand I_43440 (I742076,I742037,I741946);
nand I_43441 (I741654,I741929,I742076);
not I_43442 (I742107,I742037);
nor I_43443 (I742124,I742107,I741847);
DFFARX1 I_43444 (I742124,I3563,I741677,I741666,);
nor I_43445 (I742155,I993047,I993050);
or I_43446 (I741657,I741904,I742155);
nor I_43447 (I741648,I742037,I742155);
or I_43448 (I741651,I741771,I742155);
DFFARX1 I_43449 (I742155,I3563,I741677,I741669,);
not I_43450 (I742255,I3570);
DFFARX1 I_43451 (I1070227,I3563,I742255,I742281,);
not I_43452 (I742289,I742281);
nand I_43453 (I742306,I1070224,I1070242);
and I_43454 (I742323,I742306,I1070239);
DFFARX1 I_43455 (I742323,I3563,I742255,I742349,);
not I_43456 (I742357,I1070221);
DFFARX1 I_43457 (I1070224,I3563,I742255,I742383,);
not I_43458 (I742391,I742383);
nor I_43459 (I742408,I742391,I742289);
and I_43460 (I742425,I742408,I1070221);
nor I_43461 (I742442,I742391,I742357);
nor I_43462 (I742238,I742349,I742442);
DFFARX1 I_43463 (I1070233,I3563,I742255,I742482,);
nor I_43464 (I742490,I742482,I742349);
not I_43465 (I742507,I742490);
not I_43466 (I742524,I742482);
nor I_43467 (I742541,I742524,I742425);
DFFARX1 I_43468 (I742541,I3563,I742255,I742241,);
nand I_43469 (I742572,I1070236,I1070221);
and I_43470 (I742589,I742572,I1070227);
DFFARX1 I_43471 (I742589,I3563,I742255,I742615,);
nor I_43472 (I742623,I742615,I742482);
DFFARX1 I_43473 (I742623,I3563,I742255,I742223,);
nand I_43474 (I742654,I742615,I742524);
nand I_43475 (I742232,I742507,I742654);
not I_43476 (I742685,I742615);
nor I_43477 (I742702,I742685,I742425);
DFFARX1 I_43478 (I742702,I3563,I742255,I742244,);
nor I_43479 (I742733,I1070230,I1070221);
or I_43480 (I742235,I742482,I742733);
nor I_43481 (I742226,I742615,I742733);
or I_43482 (I742229,I742349,I742733);
DFFARX1 I_43483 (I742733,I3563,I742255,I742247,);
not I_43484 (I742833,I3570);
DFFARX1 I_43485 (I653211,I3563,I742833,I742859,);
not I_43486 (I742867,I742859);
nand I_43487 (I742884,I653220,I653229);
and I_43488 (I742901,I742884,I653235);
DFFARX1 I_43489 (I742901,I3563,I742833,I742927,);
not I_43490 (I742935,I653232);
DFFARX1 I_43491 (I653217,I3563,I742833,I742961,);
not I_43492 (I742969,I742961);
nor I_43493 (I742986,I742969,I742867);
and I_43494 (I743003,I742986,I653232);
nor I_43495 (I743020,I742969,I742935);
nor I_43496 (I742816,I742927,I743020);
DFFARX1 I_43497 (I653226,I3563,I742833,I743060,);
nor I_43498 (I743068,I743060,I742927);
not I_43499 (I743085,I743068);
not I_43500 (I743102,I743060);
nor I_43501 (I743119,I743102,I743003);
DFFARX1 I_43502 (I743119,I3563,I742833,I742819,);
nand I_43503 (I743150,I653223,I653214);
and I_43504 (I743167,I743150,I653211);
DFFARX1 I_43505 (I743167,I3563,I742833,I743193,);
nor I_43506 (I743201,I743193,I743060);
DFFARX1 I_43507 (I743201,I3563,I742833,I742801,);
nand I_43508 (I743232,I743193,I743102);
nand I_43509 (I742810,I743085,I743232);
not I_43510 (I743263,I743193);
nor I_43511 (I743280,I743263,I743003);
DFFARX1 I_43512 (I743280,I3563,I742833,I742822,);
nor I_43513 (I743311,I653214,I653214);
or I_43514 (I742813,I743060,I743311);
nor I_43515 (I742804,I743193,I743311);
or I_43516 (I742807,I742927,I743311);
DFFARX1 I_43517 (I743311,I3563,I742833,I742825,);
not I_43518 (I743411,I3570);
DFFARX1 I_43519 (I389208,I3563,I743411,I743437,);
not I_43520 (I743445,I743437);
nand I_43521 (I743462,I389211,I389187);
and I_43522 (I743479,I743462,I389184);
DFFARX1 I_43523 (I743479,I3563,I743411,I743505,);
not I_43524 (I743513,I389190);
DFFARX1 I_43525 (I389184,I3563,I743411,I743539,);
not I_43526 (I743547,I743539);
nor I_43527 (I743564,I743547,I743445);
and I_43528 (I743581,I743564,I389190);
nor I_43529 (I743598,I743547,I743513);
nor I_43530 (I743394,I743505,I743598);
DFFARX1 I_43531 (I389193,I3563,I743411,I743638,);
nor I_43532 (I743646,I743638,I743505);
not I_43533 (I743663,I743646);
not I_43534 (I743680,I743638);
nor I_43535 (I743697,I743680,I743581);
DFFARX1 I_43536 (I743697,I3563,I743411,I743397,);
nand I_43537 (I743728,I389196,I389205);
and I_43538 (I743745,I743728,I389202);
DFFARX1 I_43539 (I743745,I3563,I743411,I743771,);
nor I_43540 (I743779,I743771,I743638);
DFFARX1 I_43541 (I743779,I3563,I743411,I743379,);
nand I_43542 (I743810,I743771,I743680);
nand I_43543 (I743388,I743663,I743810);
not I_43544 (I743841,I743771);
nor I_43545 (I743858,I743841,I743581);
DFFARX1 I_43546 (I743858,I3563,I743411,I743400,);
nor I_43547 (I743889,I389199,I389205);
or I_43548 (I743391,I743638,I743889);
nor I_43549 (I743382,I743771,I743889);
or I_43550 (I743385,I743505,I743889);
DFFARX1 I_43551 (I743889,I3563,I743411,I743403,);
not I_43552 (I743989,I3570);
DFFARX1 I_43553 (I167283,I3563,I743989,I744015,);
not I_43554 (I744023,I744015);
nand I_43555 (I744040,I167286,I167307);
and I_43556 (I744057,I744040,I167295);
DFFARX1 I_43557 (I744057,I3563,I743989,I744083,);
not I_43558 (I744091,I167292);
DFFARX1 I_43559 (I167283,I3563,I743989,I744117,);
not I_43560 (I744125,I744117);
nor I_43561 (I744142,I744125,I744023);
and I_43562 (I744159,I744142,I167292);
nor I_43563 (I744176,I744125,I744091);
nor I_43564 (I743972,I744083,I744176);
DFFARX1 I_43565 (I167301,I3563,I743989,I744216,);
nor I_43566 (I744224,I744216,I744083);
not I_43567 (I744241,I744224);
not I_43568 (I744258,I744216);
nor I_43569 (I744275,I744258,I744159);
DFFARX1 I_43570 (I744275,I3563,I743989,I743975,);
nand I_43571 (I744306,I167286,I167289);
and I_43572 (I744323,I744306,I167298);
DFFARX1 I_43573 (I744323,I3563,I743989,I744349,);
nor I_43574 (I744357,I744349,I744216);
DFFARX1 I_43575 (I744357,I3563,I743989,I743957,);
nand I_43576 (I744388,I744349,I744258);
nand I_43577 (I743966,I744241,I744388);
not I_43578 (I744419,I744349);
nor I_43579 (I744436,I744419,I744159);
DFFARX1 I_43580 (I744436,I3563,I743989,I743978,);
nor I_43581 (I744467,I167304,I167289);
or I_43582 (I743969,I744216,I744467);
nor I_43583 (I743960,I744349,I744467);
or I_43584 (I743963,I744083,I744467);
DFFARX1 I_43585 (I744467,I3563,I743989,I743981,);
not I_43586 (I744567,I3570);
DFFARX1 I_43587 (I467563,I3563,I744567,I744593,);
not I_43588 (I744601,I744593);
nand I_43589 (I744618,I467554,I467572);
and I_43590 (I744635,I744618,I467575);
DFFARX1 I_43591 (I744635,I3563,I744567,I744661,);
not I_43592 (I744669,I467569);
DFFARX1 I_43593 (I467557,I3563,I744567,I744695,);
not I_43594 (I744703,I744695);
nor I_43595 (I744720,I744703,I744601);
and I_43596 (I744737,I744720,I467569);
nor I_43597 (I744754,I744703,I744669);
nor I_43598 (I744550,I744661,I744754);
DFFARX1 I_43599 (I467566,I3563,I744567,I744794,);
nor I_43600 (I744802,I744794,I744661);
not I_43601 (I744819,I744802);
not I_43602 (I744836,I744794);
nor I_43603 (I744853,I744836,I744737);
DFFARX1 I_43604 (I744853,I3563,I744567,I744553,);
nand I_43605 (I744884,I467581,I467578);
and I_43606 (I744901,I744884,I467560);
DFFARX1 I_43607 (I744901,I3563,I744567,I744927,);
nor I_43608 (I744935,I744927,I744794);
DFFARX1 I_43609 (I744935,I3563,I744567,I744535,);
nand I_43610 (I744966,I744927,I744836);
nand I_43611 (I744544,I744819,I744966);
not I_43612 (I744997,I744927);
nor I_43613 (I745014,I744997,I744737);
DFFARX1 I_43614 (I745014,I3563,I744567,I744556,);
nor I_43615 (I745045,I467554,I467578);
or I_43616 (I744547,I744794,I745045);
nor I_43617 (I744538,I744927,I745045);
or I_43618 (I744541,I744661,I745045);
DFFARX1 I_43619 (I745045,I3563,I744567,I744559,);
not I_43620 (I745145,I3570);
DFFARX1 I_43621 (I501835,I3563,I745145,I745171,);
not I_43622 (I745179,I745171);
nand I_43623 (I745196,I501826,I501844);
and I_43624 (I745213,I745196,I501847);
DFFARX1 I_43625 (I745213,I3563,I745145,I745239,);
not I_43626 (I745247,I501841);
DFFARX1 I_43627 (I501829,I3563,I745145,I745273,);
not I_43628 (I745281,I745273);
nor I_43629 (I745298,I745281,I745179);
and I_43630 (I745315,I745298,I501841);
nor I_43631 (I745332,I745281,I745247);
nor I_43632 (I745128,I745239,I745332);
DFFARX1 I_43633 (I501838,I3563,I745145,I745372,);
nor I_43634 (I745380,I745372,I745239);
not I_43635 (I745397,I745380);
not I_43636 (I745414,I745372);
nor I_43637 (I745431,I745414,I745315);
DFFARX1 I_43638 (I745431,I3563,I745145,I745131,);
nand I_43639 (I745462,I501853,I501850);
and I_43640 (I745479,I745462,I501832);
DFFARX1 I_43641 (I745479,I3563,I745145,I745505,);
nor I_43642 (I745513,I745505,I745372);
DFFARX1 I_43643 (I745513,I3563,I745145,I745113,);
nand I_43644 (I745544,I745505,I745414);
nand I_43645 (I745122,I745397,I745544);
not I_43646 (I745575,I745505);
nor I_43647 (I745592,I745575,I745315);
DFFARX1 I_43648 (I745592,I3563,I745145,I745134,);
nor I_43649 (I745623,I501826,I501850);
or I_43650 (I745125,I745372,I745623);
nor I_43651 (I745116,I745505,I745623);
or I_43652 (I745119,I745239,I745623);
DFFARX1 I_43653 (I745623,I3563,I745145,I745137,);
not I_43654 (I745723,I3570);
DFFARX1 I_43655 (I156780,I3563,I745723,I745749,);
not I_43656 (I745757,I745749);
nand I_43657 (I745774,I156789,I156798);
and I_43658 (I745791,I745774,I156777);
DFFARX1 I_43659 (I745791,I3563,I745723,I745817,);
not I_43660 (I745825,I156780);
DFFARX1 I_43661 (I156795,I3563,I745723,I745851,);
not I_43662 (I745859,I745851);
nor I_43663 (I745876,I745859,I745757);
and I_43664 (I745893,I745876,I156780);
nor I_43665 (I745910,I745859,I745825);
nor I_43666 (I745706,I745817,I745910);
DFFARX1 I_43667 (I156786,I3563,I745723,I745950,);
nor I_43668 (I745958,I745950,I745817);
not I_43669 (I745975,I745958);
not I_43670 (I745992,I745950);
nor I_43671 (I746009,I745992,I745893);
DFFARX1 I_43672 (I746009,I3563,I745723,I745709,);
nand I_43673 (I746040,I156801,I156777);
and I_43674 (I746057,I746040,I156783);
DFFARX1 I_43675 (I746057,I3563,I745723,I746083,);
nor I_43676 (I746091,I746083,I745950);
DFFARX1 I_43677 (I746091,I3563,I745723,I745691,);
nand I_43678 (I746122,I746083,I745992);
nand I_43679 (I745700,I745975,I746122);
not I_43680 (I746153,I746083);
nor I_43681 (I746170,I746153,I745893);
DFFARX1 I_43682 (I746170,I3563,I745723,I745712,);
nor I_43683 (I746201,I156792,I156777);
or I_43684 (I745703,I745950,I746201);
nor I_43685 (I745694,I746083,I746201);
or I_43686 (I745697,I745817,I746201);
DFFARX1 I_43687 (I746201,I3563,I745723,I745715,);
not I_43688 (I746301,I3570);
DFFARX1 I_43689 (I1314341,I3563,I746301,I746327,);
not I_43690 (I746335,I746327);
nand I_43691 (I746352,I1314365,I1314347);
and I_43692 (I746369,I746352,I1314353);
DFFARX1 I_43693 (I746369,I3563,I746301,I746395,);
not I_43694 (I746403,I1314359);
DFFARX1 I_43695 (I1314344,I3563,I746301,I746429,);
not I_43696 (I746437,I746429);
nor I_43697 (I746454,I746437,I746335);
and I_43698 (I746471,I746454,I1314359);
nor I_43699 (I746488,I746437,I746403);
nor I_43700 (I746284,I746395,I746488);
DFFARX1 I_43701 (I1314356,I3563,I746301,I746528,);
nor I_43702 (I746536,I746528,I746395);
not I_43703 (I746553,I746536);
not I_43704 (I746570,I746528);
nor I_43705 (I746587,I746570,I746471);
DFFARX1 I_43706 (I746587,I3563,I746301,I746287,);
nand I_43707 (I746618,I1314362,I1314350);
and I_43708 (I746635,I746618,I1314344);
DFFARX1 I_43709 (I746635,I3563,I746301,I746661,);
nor I_43710 (I746669,I746661,I746528);
DFFARX1 I_43711 (I746669,I3563,I746301,I746269,);
nand I_43712 (I746700,I746661,I746570);
nand I_43713 (I746278,I746553,I746700);
not I_43714 (I746731,I746661);
nor I_43715 (I746748,I746731,I746471);
DFFARX1 I_43716 (I746748,I3563,I746301,I746290,);
nor I_43717 (I746779,I1314341,I1314350);
or I_43718 (I746281,I746528,I746779);
nor I_43719 (I746272,I746661,I746779);
or I_43720 (I746275,I746395,I746779);
DFFARX1 I_43721 (I746779,I3563,I746301,I746293,);
not I_43722 (I746879,I3570);
DFFARX1 I_43723 (I1376180,I3563,I746879,I746905,);
not I_43724 (I746913,I746905);
nand I_43725 (I746930,I1376165,I1376153);
and I_43726 (I746947,I746930,I1376168);
DFFARX1 I_43727 (I746947,I3563,I746879,I746973,);
not I_43728 (I746981,I1376153);
DFFARX1 I_43729 (I1376171,I3563,I746879,I747007,);
not I_43730 (I747015,I747007);
nor I_43731 (I747032,I747015,I746913);
and I_43732 (I747049,I747032,I1376153);
nor I_43733 (I747066,I747015,I746981);
nor I_43734 (I746862,I746973,I747066);
DFFARX1 I_43735 (I1376159,I3563,I746879,I747106,);
nor I_43736 (I747114,I747106,I746973);
not I_43737 (I747131,I747114);
not I_43738 (I747148,I747106);
nor I_43739 (I747165,I747148,I747049);
DFFARX1 I_43740 (I747165,I3563,I746879,I746865,);
nand I_43741 (I747196,I1376156,I1376162);
and I_43742 (I747213,I747196,I1376177);
DFFARX1 I_43743 (I747213,I3563,I746879,I747239,);
nor I_43744 (I747247,I747239,I747106);
DFFARX1 I_43745 (I747247,I3563,I746879,I746847,);
nand I_43746 (I747278,I747239,I747148);
nand I_43747 (I746856,I747131,I747278);
not I_43748 (I747309,I747239);
nor I_43749 (I747326,I747309,I747049);
DFFARX1 I_43750 (I747326,I3563,I746879,I746868,);
nor I_43751 (I747357,I1376174,I1376162);
or I_43752 (I746859,I747106,I747357);
nor I_43753 (I746850,I747239,I747357);
or I_43754 (I746853,I746973,I747357);
DFFARX1 I_43755 (I747357,I3563,I746879,I746871,);
not I_43756 (I747457,I3570);
DFFARX1 I_43757 (I564386,I3563,I747457,I747483,);
not I_43758 (I747491,I747483);
nand I_43759 (I747508,I564401,I564386);
and I_43760 (I747525,I747508,I564389);
DFFARX1 I_43761 (I747525,I3563,I747457,I747551,);
not I_43762 (I747559,I564389);
DFFARX1 I_43763 (I564398,I3563,I747457,I747585,);
not I_43764 (I747593,I747585);
nor I_43765 (I747610,I747593,I747491);
and I_43766 (I747627,I747610,I564389);
nor I_43767 (I747644,I747593,I747559);
nor I_43768 (I747440,I747551,I747644);
DFFARX1 I_43769 (I564392,I3563,I747457,I747684,);
nor I_43770 (I747692,I747684,I747551);
not I_43771 (I747709,I747692);
not I_43772 (I747726,I747684);
nor I_43773 (I747743,I747726,I747627);
DFFARX1 I_43774 (I747743,I3563,I747457,I747443,);
nand I_43775 (I747774,I564395,I564404);
and I_43776 (I747791,I747774,I564410);
DFFARX1 I_43777 (I747791,I3563,I747457,I747817,);
nor I_43778 (I747825,I747817,I747684);
DFFARX1 I_43779 (I747825,I3563,I747457,I747425,);
nand I_43780 (I747856,I747817,I747726);
nand I_43781 (I747434,I747709,I747856);
not I_43782 (I747887,I747817);
nor I_43783 (I747904,I747887,I747627);
DFFARX1 I_43784 (I747904,I3563,I747457,I747446,);
nor I_43785 (I747935,I564407,I564404);
or I_43786 (I747437,I747684,I747935);
nor I_43787 (I747428,I747817,I747935);
or I_43788 (I747431,I747551,I747935);
DFFARX1 I_43789 (I747935,I3563,I747457,I747449,);
not I_43790 (I748035,I3570);
DFFARX1 I_43791 (I1338100,I3563,I748035,I748061,);
not I_43792 (I748069,I748061);
nand I_43793 (I748086,I1338085,I1338073);
and I_43794 (I748103,I748086,I1338088);
DFFARX1 I_43795 (I748103,I3563,I748035,I748129,);
not I_43796 (I748137,I1338073);
DFFARX1 I_43797 (I1338091,I3563,I748035,I748163,);
not I_43798 (I748171,I748163);
nor I_43799 (I748188,I748171,I748069);
and I_43800 (I748205,I748188,I1338073);
nor I_43801 (I748222,I748171,I748137);
nor I_43802 (I748018,I748129,I748222);
DFFARX1 I_43803 (I1338079,I3563,I748035,I748262,);
nor I_43804 (I748270,I748262,I748129);
not I_43805 (I748287,I748270);
not I_43806 (I748304,I748262);
nor I_43807 (I748321,I748304,I748205);
DFFARX1 I_43808 (I748321,I3563,I748035,I748021,);
nand I_43809 (I748352,I1338076,I1338082);
and I_43810 (I748369,I748352,I1338097);
DFFARX1 I_43811 (I748369,I3563,I748035,I748395,);
nor I_43812 (I748403,I748395,I748262);
DFFARX1 I_43813 (I748403,I3563,I748035,I748003,);
nand I_43814 (I748434,I748395,I748304);
nand I_43815 (I748012,I748287,I748434);
not I_43816 (I748465,I748395);
nor I_43817 (I748482,I748465,I748205);
DFFARX1 I_43818 (I748482,I3563,I748035,I748024,);
nor I_43819 (I748513,I1338094,I1338082);
or I_43820 (I748015,I748262,I748513);
nor I_43821 (I748006,I748395,I748513);
or I_43822 (I748009,I748129,I748513);
DFFARX1 I_43823 (I748513,I3563,I748035,I748027,);
not I_43824 (I748613,I3570);
DFFARX1 I_43825 (I1236669,I3563,I748613,I748639,);
not I_43826 (I748647,I748639);
nand I_43827 (I748664,I1236651,I1236663);
and I_43828 (I748681,I748664,I1236666);
DFFARX1 I_43829 (I748681,I3563,I748613,I748707,);
not I_43830 (I748715,I1236660);
DFFARX1 I_43831 (I1236657,I3563,I748613,I748741,);
not I_43832 (I748749,I748741);
nor I_43833 (I748766,I748749,I748647);
and I_43834 (I748783,I748766,I1236660);
nor I_43835 (I748800,I748749,I748715);
nor I_43836 (I748596,I748707,I748800);
DFFARX1 I_43837 (I1236675,I3563,I748613,I748840,);
nor I_43838 (I748848,I748840,I748707);
not I_43839 (I748865,I748848);
not I_43840 (I748882,I748840);
nor I_43841 (I748899,I748882,I748783);
DFFARX1 I_43842 (I748899,I3563,I748613,I748599,);
nand I_43843 (I748930,I1236654,I1236654);
and I_43844 (I748947,I748930,I1236651);
DFFARX1 I_43845 (I748947,I3563,I748613,I748973,);
nor I_43846 (I748981,I748973,I748840);
DFFARX1 I_43847 (I748981,I3563,I748613,I748581,);
nand I_43848 (I749012,I748973,I748882);
nand I_43849 (I748590,I748865,I749012);
not I_43850 (I749043,I748973);
nor I_43851 (I749060,I749043,I748783);
DFFARX1 I_43852 (I749060,I3563,I748613,I748602,);
nor I_43853 (I749091,I1236672,I1236654);
or I_43854 (I748593,I748840,I749091);
nor I_43855 (I748584,I748973,I749091);
or I_43856 (I748587,I748707,I749091);
DFFARX1 I_43857 (I749091,I3563,I748613,I748605,);
not I_43858 (I749191,I3570);
DFFARX1 I_43859 (I1279593,I3563,I749191,I749217,);
not I_43860 (I749225,I749217);
nand I_43861 (I749242,I1279596,I1279605);
and I_43862 (I749259,I749242,I1279608);
DFFARX1 I_43863 (I749259,I3563,I749191,I749285,);
not I_43864 (I749293,I1279617);
DFFARX1 I_43865 (I1279599,I3563,I749191,I749319,);
not I_43866 (I749327,I749319);
nor I_43867 (I749344,I749327,I749225);
and I_43868 (I749361,I749344,I1279617);
nor I_43869 (I749378,I749327,I749293);
nor I_43870 (I749174,I749285,I749378);
DFFARX1 I_43871 (I1279596,I3563,I749191,I749418,);
nor I_43872 (I749426,I749418,I749285);
not I_43873 (I749443,I749426);
not I_43874 (I749460,I749418);
nor I_43875 (I749477,I749460,I749361);
DFFARX1 I_43876 (I749477,I3563,I749191,I749177,);
nand I_43877 (I749508,I1279614,I1279593);
and I_43878 (I749525,I749508,I1279611);
DFFARX1 I_43879 (I749525,I3563,I749191,I749551,);
nor I_43880 (I749559,I749551,I749418);
DFFARX1 I_43881 (I749559,I3563,I749191,I749159,);
nand I_43882 (I749590,I749551,I749460);
nand I_43883 (I749168,I749443,I749590);
not I_43884 (I749621,I749551);
nor I_43885 (I749638,I749621,I749361);
DFFARX1 I_43886 (I749638,I3563,I749191,I749180,);
nor I_43887 (I749669,I1279602,I1279593);
or I_43888 (I749171,I749418,I749669);
nor I_43889 (I749162,I749551,I749669);
or I_43890 (I749165,I749285,I749669);
DFFARX1 I_43891 (I749669,I3563,I749191,I749183,);
not I_43892 (I749769,I3570);
DFFARX1 I_43893 (I1292955,I3563,I749769,I749795,);
not I_43894 (I749803,I749795);
nand I_43895 (I749820,I1292979,I1292961);
and I_43896 (I749837,I749820,I1292967);
DFFARX1 I_43897 (I749837,I3563,I749769,I749863,);
not I_43898 (I749871,I1292973);
DFFARX1 I_43899 (I1292958,I3563,I749769,I749897,);
not I_43900 (I749905,I749897);
nor I_43901 (I749922,I749905,I749803);
and I_43902 (I749939,I749922,I1292973);
nor I_43903 (I749956,I749905,I749871);
nor I_43904 (I749752,I749863,I749956);
DFFARX1 I_43905 (I1292970,I3563,I749769,I749996,);
nor I_43906 (I750004,I749996,I749863);
not I_43907 (I750021,I750004);
not I_43908 (I750038,I749996);
nor I_43909 (I750055,I750038,I749939);
DFFARX1 I_43910 (I750055,I3563,I749769,I749755,);
nand I_43911 (I750086,I1292976,I1292964);
and I_43912 (I750103,I750086,I1292958);
DFFARX1 I_43913 (I750103,I3563,I749769,I750129,);
nor I_43914 (I750137,I750129,I749996);
DFFARX1 I_43915 (I750137,I3563,I749769,I749737,);
nand I_43916 (I750168,I750129,I750038);
nand I_43917 (I749746,I750021,I750168);
not I_43918 (I750199,I750129);
nor I_43919 (I750216,I750199,I749939);
DFFARX1 I_43920 (I750216,I3563,I749769,I749758,);
nor I_43921 (I750247,I1292955,I1292964);
or I_43922 (I749749,I749996,I750247);
nor I_43923 (I749740,I750129,I750247);
or I_43924 (I749743,I749863,I750247);
DFFARX1 I_43925 (I750247,I3563,I749769,I749761,);
not I_43926 (I750347,I3570);
DFFARX1 I_43927 (I453419,I3563,I750347,I750373,);
not I_43928 (I750381,I750373);
nand I_43929 (I750398,I453410,I453428);
and I_43930 (I750415,I750398,I453431);
DFFARX1 I_43931 (I750415,I3563,I750347,I750441,);
not I_43932 (I750449,I453425);
DFFARX1 I_43933 (I453413,I3563,I750347,I750475,);
not I_43934 (I750483,I750475);
nor I_43935 (I750500,I750483,I750381);
and I_43936 (I750517,I750500,I453425);
nor I_43937 (I750534,I750483,I750449);
nor I_43938 (I750330,I750441,I750534);
DFFARX1 I_43939 (I453422,I3563,I750347,I750574,);
nor I_43940 (I750582,I750574,I750441);
not I_43941 (I750599,I750582);
not I_43942 (I750616,I750574);
nor I_43943 (I750633,I750616,I750517);
DFFARX1 I_43944 (I750633,I3563,I750347,I750333,);
nand I_43945 (I750664,I453437,I453434);
and I_43946 (I750681,I750664,I453416);
DFFARX1 I_43947 (I750681,I3563,I750347,I750707,);
nor I_43948 (I750715,I750707,I750574);
DFFARX1 I_43949 (I750715,I3563,I750347,I750315,);
nand I_43950 (I750746,I750707,I750616);
nand I_43951 (I750324,I750599,I750746);
not I_43952 (I750777,I750707);
nor I_43953 (I750794,I750777,I750517);
DFFARX1 I_43954 (I750794,I3563,I750347,I750336,);
nor I_43955 (I750825,I453410,I453434);
or I_43956 (I750327,I750574,I750825);
nor I_43957 (I750318,I750707,I750825);
or I_43958 (I750321,I750441,I750825);
DFFARX1 I_43959 (I750825,I3563,I750347,I750339,);
not I_43960 (I750925,I3570);
DFFARX1 I_43961 (I826354,I3563,I750925,I750951,);
not I_43962 (I750959,I750951);
nand I_43963 (I750976,I826342,I826360);
and I_43964 (I750993,I750976,I826357);
DFFARX1 I_43965 (I750993,I3563,I750925,I751019,);
not I_43966 (I751027,I826348);
DFFARX1 I_43967 (I826345,I3563,I750925,I751053,);
not I_43968 (I751061,I751053);
nor I_43969 (I751078,I751061,I750959);
and I_43970 (I751095,I751078,I826348);
nor I_43971 (I751112,I751061,I751027);
nor I_43972 (I750908,I751019,I751112);
DFFARX1 I_43973 (I826339,I3563,I750925,I751152,);
nor I_43974 (I751160,I751152,I751019);
not I_43975 (I751177,I751160);
not I_43976 (I751194,I751152);
nor I_43977 (I751211,I751194,I751095);
DFFARX1 I_43978 (I751211,I3563,I750925,I750911,);
nand I_43979 (I751242,I826339,I826342);
and I_43980 (I751259,I751242,I826345);
DFFARX1 I_43981 (I751259,I3563,I750925,I751285,);
nor I_43982 (I751293,I751285,I751152);
DFFARX1 I_43983 (I751293,I3563,I750925,I750893,);
nand I_43984 (I751324,I751285,I751194);
nand I_43985 (I750902,I751177,I751324);
not I_43986 (I751355,I751285);
nor I_43987 (I751372,I751355,I751095);
DFFARX1 I_43988 (I751372,I3563,I750925,I750914,);
nor I_43989 (I751403,I826351,I826342);
or I_43990 (I750905,I751152,I751403);
nor I_43991 (I750896,I751285,I751403);
or I_43992 (I750899,I751019,I751403);
DFFARX1 I_43993 (I751403,I3563,I750925,I750917,);
not I_43994 (I751503,I3570);
DFFARX1 I_43995 (I523051,I3563,I751503,I751529,);
not I_43996 (I751537,I751529);
nand I_43997 (I751554,I523042,I523060);
and I_43998 (I751571,I751554,I523063);
DFFARX1 I_43999 (I751571,I3563,I751503,I751597,);
not I_44000 (I751605,I523057);
DFFARX1 I_44001 (I523045,I3563,I751503,I751631,);
not I_44002 (I751639,I751631);
nor I_44003 (I751656,I751639,I751537);
and I_44004 (I751673,I751656,I523057);
nor I_44005 (I751690,I751639,I751605);
nor I_44006 (I751486,I751597,I751690);
DFFARX1 I_44007 (I523054,I3563,I751503,I751730,);
nor I_44008 (I751738,I751730,I751597);
not I_44009 (I751755,I751738);
not I_44010 (I751772,I751730);
nor I_44011 (I751789,I751772,I751673);
DFFARX1 I_44012 (I751789,I3563,I751503,I751489,);
nand I_44013 (I751820,I523069,I523066);
and I_44014 (I751837,I751820,I523048);
DFFARX1 I_44015 (I751837,I3563,I751503,I751863,);
nor I_44016 (I751871,I751863,I751730);
DFFARX1 I_44017 (I751871,I3563,I751503,I751471,);
nand I_44018 (I751902,I751863,I751772);
nand I_44019 (I751480,I751755,I751902);
not I_44020 (I751933,I751863);
nor I_44021 (I751950,I751933,I751673);
DFFARX1 I_44022 (I751950,I3563,I751503,I751492,);
nor I_44023 (I751981,I523042,I523066);
or I_44024 (I751483,I751730,I751981);
nor I_44025 (I751474,I751863,I751981);
or I_44026 (I751477,I751597,I751981);
DFFARX1 I_44027 (I751981,I3563,I751503,I751495,);
not I_44028 (I752081,I3570);
DFFARX1 I_44029 (I1241871,I3563,I752081,I752107,);
not I_44030 (I752115,I752107);
nand I_44031 (I752132,I1241853,I1241865);
and I_44032 (I752149,I752132,I1241868);
DFFARX1 I_44033 (I752149,I3563,I752081,I752175,);
not I_44034 (I752183,I1241862);
DFFARX1 I_44035 (I1241859,I3563,I752081,I752209,);
not I_44036 (I752217,I752209);
nor I_44037 (I752234,I752217,I752115);
and I_44038 (I752251,I752234,I1241862);
nor I_44039 (I752268,I752217,I752183);
nor I_44040 (I752064,I752175,I752268);
DFFARX1 I_44041 (I1241877,I3563,I752081,I752308,);
nor I_44042 (I752316,I752308,I752175);
not I_44043 (I752333,I752316);
not I_44044 (I752350,I752308);
nor I_44045 (I752367,I752350,I752251);
DFFARX1 I_44046 (I752367,I3563,I752081,I752067,);
nand I_44047 (I752398,I1241856,I1241856);
and I_44048 (I752415,I752398,I1241853);
DFFARX1 I_44049 (I752415,I3563,I752081,I752441,);
nor I_44050 (I752449,I752441,I752308);
DFFARX1 I_44051 (I752449,I3563,I752081,I752049,);
nand I_44052 (I752480,I752441,I752350);
nand I_44053 (I752058,I752333,I752480);
not I_44054 (I752511,I752441);
nor I_44055 (I752528,I752511,I752251);
DFFARX1 I_44056 (I752528,I3563,I752081,I752070,);
nor I_44057 (I752559,I1241874,I1241856);
or I_44058 (I752061,I752308,I752559);
nor I_44059 (I752052,I752441,I752559);
or I_44060 (I752055,I752175,I752559);
DFFARX1 I_44061 (I752559,I3563,I752081,I752073,);
not I_44062 (I752659,I3570);
DFFARX1 I_44063 (I1259465,I3563,I752659,I752685,);
not I_44064 (I752693,I752685);
nand I_44065 (I752710,I1259468,I1259477);
and I_44066 (I752727,I752710,I1259480);
DFFARX1 I_44067 (I752727,I3563,I752659,I752753,);
not I_44068 (I752761,I1259489);
DFFARX1 I_44069 (I1259471,I3563,I752659,I752787,);
not I_44070 (I752795,I752787);
nor I_44071 (I752812,I752795,I752693);
and I_44072 (I752829,I752812,I1259489);
nor I_44073 (I752846,I752795,I752761);
nor I_44074 (I752642,I752753,I752846);
DFFARX1 I_44075 (I1259468,I3563,I752659,I752886,);
nor I_44076 (I752894,I752886,I752753);
not I_44077 (I752911,I752894);
not I_44078 (I752928,I752886);
nor I_44079 (I752945,I752928,I752829);
DFFARX1 I_44080 (I752945,I3563,I752659,I752645,);
nand I_44081 (I752976,I1259486,I1259465);
and I_44082 (I752993,I752976,I1259483);
DFFARX1 I_44083 (I752993,I3563,I752659,I753019,);
nor I_44084 (I753027,I753019,I752886);
DFFARX1 I_44085 (I753027,I3563,I752659,I752627,);
nand I_44086 (I753058,I753019,I752928);
nand I_44087 (I752636,I752911,I753058);
not I_44088 (I753089,I753019);
nor I_44089 (I753106,I753089,I752829);
DFFARX1 I_44090 (I753106,I3563,I752659,I752648,);
nor I_44091 (I753137,I1259474,I1259465);
or I_44092 (I752639,I752886,I753137);
nor I_44093 (I752630,I753019,I753137);
or I_44094 (I752633,I752753,I753137);
DFFARX1 I_44095 (I753137,I3563,I752659,I752651,);
not I_44096 (I753237,I3570);
DFFARX1 I_44097 (I960765,I3563,I753237,I753263,);
not I_44098 (I753271,I753263);
nand I_44099 (I753288,I960741,I960756);
and I_44100 (I753305,I753288,I960768);
DFFARX1 I_44101 (I753305,I3563,I753237,I753331,);
not I_44102 (I753339,I960753);
DFFARX1 I_44103 (I960744,I3563,I753237,I753365,);
not I_44104 (I753373,I753365);
nor I_44105 (I753390,I753373,I753271);
and I_44106 (I753407,I753390,I960753);
nor I_44107 (I753424,I753373,I753339);
nor I_44108 (I753220,I753331,I753424);
DFFARX1 I_44109 (I960741,I3563,I753237,I753464,);
nor I_44110 (I753472,I753464,I753331);
not I_44111 (I753489,I753472);
not I_44112 (I753506,I753464);
nor I_44113 (I753523,I753506,I753407);
DFFARX1 I_44114 (I753523,I3563,I753237,I753223,);
nand I_44115 (I753554,I960759,I960750);
and I_44116 (I753571,I753554,I960762);
DFFARX1 I_44117 (I753571,I3563,I753237,I753597,);
nor I_44118 (I753605,I753597,I753464);
DFFARX1 I_44119 (I753605,I3563,I753237,I753205,);
nand I_44120 (I753636,I753597,I753506);
nand I_44121 (I753214,I753489,I753636);
not I_44122 (I753667,I753597);
nor I_44123 (I753684,I753667,I753407);
DFFARX1 I_44124 (I753684,I3563,I753237,I753226,);
nor I_44125 (I753715,I960747,I960750);
or I_44126 (I753217,I753464,I753715);
nor I_44127 (I753208,I753597,I753715);
or I_44128 (I753211,I753331,I753715);
DFFARX1 I_44129 (I753715,I3563,I753237,I753229,);
not I_44130 (I753815,I3570);
DFFARX1 I_44131 (I323333,I3563,I753815,I753841,);
not I_44132 (I753849,I753841);
nand I_44133 (I753866,I323336,I323312);
and I_44134 (I753883,I753866,I323309);
DFFARX1 I_44135 (I753883,I3563,I753815,I753909,);
not I_44136 (I753917,I323315);
DFFARX1 I_44137 (I323309,I3563,I753815,I753943,);
not I_44138 (I753951,I753943);
nor I_44139 (I753968,I753951,I753849);
and I_44140 (I753985,I753968,I323315);
nor I_44141 (I754002,I753951,I753917);
nor I_44142 (I753798,I753909,I754002);
DFFARX1 I_44143 (I323318,I3563,I753815,I754042,);
nor I_44144 (I754050,I754042,I753909);
not I_44145 (I754067,I754050);
not I_44146 (I754084,I754042);
nor I_44147 (I754101,I754084,I753985);
DFFARX1 I_44148 (I754101,I3563,I753815,I753801,);
nand I_44149 (I754132,I323321,I323330);
and I_44150 (I754149,I754132,I323327);
DFFARX1 I_44151 (I754149,I3563,I753815,I754175,);
nor I_44152 (I754183,I754175,I754042);
DFFARX1 I_44153 (I754183,I3563,I753815,I753783,);
nand I_44154 (I754214,I754175,I754084);
nand I_44155 (I753792,I754067,I754214);
not I_44156 (I754245,I754175);
nor I_44157 (I754262,I754245,I753985);
DFFARX1 I_44158 (I754262,I3563,I753815,I753804,);
nor I_44159 (I754293,I323324,I323330);
or I_44160 (I753795,I754042,I754293);
nor I_44161 (I753786,I754175,I754293);
or I_44162 (I753789,I753909,I754293);
DFFARX1 I_44163 (I754293,I3563,I753815,I753807,);
not I_44164 (I754393,I3570);
DFFARX1 I_44165 (I359696,I3563,I754393,I754419,);
not I_44166 (I754427,I754419);
nand I_44167 (I754444,I359699,I359675);
and I_44168 (I754461,I754444,I359672);
DFFARX1 I_44169 (I754461,I3563,I754393,I754487,);
not I_44170 (I754495,I359678);
DFFARX1 I_44171 (I359672,I3563,I754393,I754521,);
not I_44172 (I754529,I754521);
nor I_44173 (I754546,I754529,I754427);
and I_44174 (I754563,I754546,I359678);
nor I_44175 (I754580,I754529,I754495);
nor I_44176 (I754376,I754487,I754580);
DFFARX1 I_44177 (I359681,I3563,I754393,I754620,);
nor I_44178 (I754628,I754620,I754487);
not I_44179 (I754645,I754628);
not I_44180 (I754662,I754620);
nor I_44181 (I754679,I754662,I754563);
DFFARX1 I_44182 (I754679,I3563,I754393,I754379,);
nand I_44183 (I754710,I359684,I359693);
and I_44184 (I754727,I754710,I359690);
DFFARX1 I_44185 (I754727,I3563,I754393,I754753,);
nor I_44186 (I754761,I754753,I754620);
DFFARX1 I_44187 (I754761,I3563,I754393,I754361,);
nand I_44188 (I754792,I754753,I754662);
nand I_44189 (I754370,I754645,I754792);
not I_44190 (I754823,I754753);
nor I_44191 (I754840,I754823,I754563);
DFFARX1 I_44192 (I754840,I3563,I754393,I754382,);
nor I_44193 (I754871,I359687,I359693);
or I_44194 (I754373,I754620,I754871);
nor I_44195 (I754364,I754753,I754871);
or I_44196 (I754367,I754487,I754871);
DFFARX1 I_44197 (I754871,I3563,I754393,I754385,);
not I_44198 (I754971,I3570);
DFFARX1 I_44199 (I69825,I3563,I754971,I754997,);
not I_44200 (I755005,I754997);
nand I_44201 (I755022,I69834,I69843);
and I_44202 (I755039,I755022,I69822);
DFFARX1 I_44203 (I755039,I3563,I754971,I755065,);
not I_44204 (I755073,I69825);
DFFARX1 I_44205 (I69840,I3563,I754971,I755099,);
not I_44206 (I755107,I755099);
nor I_44207 (I755124,I755107,I755005);
and I_44208 (I755141,I755124,I69825);
nor I_44209 (I755158,I755107,I755073);
nor I_44210 (I754954,I755065,I755158);
DFFARX1 I_44211 (I69831,I3563,I754971,I755198,);
nor I_44212 (I755206,I755198,I755065);
not I_44213 (I755223,I755206);
not I_44214 (I755240,I755198);
nor I_44215 (I755257,I755240,I755141);
DFFARX1 I_44216 (I755257,I3563,I754971,I754957,);
nand I_44217 (I755288,I69846,I69822);
and I_44218 (I755305,I755288,I69828);
DFFARX1 I_44219 (I755305,I3563,I754971,I755331,);
nor I_44220 (I755339,I755331,I755198);
DFFARX1 I_44221 (I755339,I3563,I754971,I754939,);
nand I_44222 (I755370,I755331,I755240);
nand I_44223 (I754948,I755223,I755370);
not I_44224 (I755401,I755331);
nor I_44225 (I755418,I755401,I755141);
DFFARX1 I_44226 (I755418,I3563,I754971,I754960,);
nor I_44227 (I755449,I69837,I69822);
or I_44228 (I754951,I755198,I755449);
nor I_44229 (I754942,I755331,I755449);
or I_44230 (I754945,I755065,I755449);
DFFARX1 I_44231 (I755449,I3563,I754971,I754963,);
not I_44232 (I755549,I3570);
DFFARX1 I_44233 (I36633,I3563,I755549,I755575,);
not I_44234 (I755583,I755575);
nand I_44235 (I755600,I36630,I36621);
and I_44236 (I755617,I755600,I36621);
DFFARX1 I_44237 (I755617,I3563,I755549,I755643,);
not I_44238 (I755651,I36624);
DFFARX1 I_44239 (I36639,I3563,I755549,I755677,);
not I_44240 (I755685,I755677);
nor I_44241 (I755702,I755685,I755583);
and I_44242 (I755719,I755702,I36624);
nor I_44243 (I755736,I755685,I755651);
nor I_44244 (I755532,I755643,I755736);
DFFARX1 I_44245 (I36624,I3563,I755549,I755776,);
nor I_44246 (I755784,I755776,I755643);
not I_44247 (I755801,I755784);
not I_44248 (I755818,I755776);
nor I_44249 (I755835,I755818,I755719);
DFFARX1 I_44250 (I755835,I3563,I755549,I755535,);
nand I_44251 (I755866,I36642,I36627);
and I_44252 (I755883,I755866,I36645);
DFFARX1 I_44253 (I755883,I3563,I755549,I755909,);
nor I_44254 (I755917,I755909,I755776);
DFFARX1 I_44255 (I755917,I3563,I755549,I755517,);
nand I_44256 (I755948,I755909,I755818);
nand I_44257 (I755526,I755801,I755948);
not I_44258 (I755979,I755909);
nor I_44259 (I755996,I755979,I755719);
DFFARX1 I_44260 (I755996,I3563,I755549,I755538,);
nor I_44261 (I756027,I36636,I36627);
or I_44262 (I755529,I755776,I756027);
nor I_44263 (I755520,I755909,I756027);
or I_44264 (I755523,I755643,I756027);
DFFARX1 I_44265 (I756027,I3563,I755549,I755541,);
not I_44266 (I756127,I3570);
DFFARX1 I_44267 (I84054,I3563,I756127,I756153,);
not I_44268 (I756161,I756153);
nand I_44269 (I756178,I84063,I84072);
and I_44270 (I756195,I756178,I84051);
DFFARX1 I_44271 (I756195,I3563,I756127,I756221,);
not I_44272 (I756229,I84054);
DFFARX1 I_44273 (I84069,I3563,I756127,I756255,);
not I_44274 (I756263,I756255);
nor I_44275 (I756280,I756263,I756161);
and I_44276 (I756297,I756280,I84054);
nor I_44277 (I756314,I756263,I756229);
nor I_44278 (I756110,I756221,I756314);
DFFARX1 I_44279 (I84060,I3563,I756127,I756354,);
nor I_44280 (I756362,I756354,I756221);
not I_44281 (I756379,I756362);
not I_44282 (I756396,I756354);
nor I_44283 (I756413,I756396,I756297);
DFFARX1 I_44284 (I756413,I3563,I756127,I756113,);
nand I_44285 (I756444,I84075,I84051);
and I_44286 (I756461,I756444,I84057);
DFFARX1 I_44287 (I756461,I3563,I756127,I756487,);
nor I_44288 (I756495,I756487,I756354);
DFFARX1 I_44289 (I756495,I3563,I756127,I756095,);
nand I_44290 (I756526,I756487,I756396);
nand I_44291 (I756104,I756379,I756526);
not I_44292 (I756557,I756487);
nor I_44293 (I756574,I756557,I756297);
DFFARX1 I_44294 (I756574,I3563,I756127,I756116,);
nor I_44295 (I756605,I84066,I84051);
or I_44296 (I756107,I756354,I756605);
nor I_44297 (I756098,I756487,I756605);
or I_44298 (I756101,I756221,I756605);
DFFARX1 I_44299 (I756605,I3563,I756127,I756119,);
not I_44300 (I756705,I3570);
DFFARX1 I_44301 (I1123381,I3563,I756705,I756731,);
not I_44302 (I756739,I756731);
nand I_44303 (I756756,I1123363,I1123375);
and I_44304 (I756773,I756756,I1123378);
DFFARX1 I_44305 (I756773,I3563,I756705,I756799,);
not I_44306 (I756807,I1123372);
DFFARX1 I_44307 (I1123369,I3563,I756705,I756833,);
not I_44308 (I756841,I756833);
nor I_44309 (I756858,I756841,I756739);
and I_44310 (I756875,I756858,I1123372);
nor I_44311 (I756892,I756841,I756807);
nor I_44312 (I756688,I756799,I756892);
DFFARX1 I_44313 (I1123387,I3563,I756705,I756932,);
nor I_44314 (I756940,I756932,I756799);
not I_44315 (I756957,I756940);
not I_44316 (I756974,I756932);
nor I_44317 (I756991,I756974,I756875);
DFFARX1 I_44318 (I756991,I3563,I756705,I756691,);
nand I_44319 (I757022,I1123366,I1123366);
and I_44320 (I757039,I757022,I1123363);
DFFARX1 I_44321 (I757039,I3563,I756705,I757065,);
nor I_44322 (I757073,I757065,I756932);
DFFARX1 I_44323 (I757073,I3563,I756705,I756673,);
nand I_44324 (I757104,I757065,I756974);
nand I_44325 (I756682,I756957,I757104);
not I_44326 (I757135,I757065);
nor I_44327 (I757152,I757135,I756875);
DFFARX1 I_44328 (I757152,I3563,I756705,I756694,);
nor I_44329 (I757183,I1123384,I1123366);
or I_44330 (I756685,I756932,I757183);
nor I_44331 (I756676,I757065,I757183);
or I_44332 (I756679,I756799,I757183);
DFFARX1 I_44333 (I757183,I3563,I756705,I756697,);
not I_44334 (I757283,I3570);
DFFARX1 I_44335 (I515979,I3563,I757283,I757309,);
not I_44336 (I757317,I757309);
nand I_44337 (I757334,I515970,I515988);
and I_44338 (I757351,I757334,I515991);
DFFARX1 I_44339 (I757351,I3563,I757283,I757377,);
not I_44340 (I757385,I515985);
DFFARX1 I_44341 (I515973,I3563,I757283,I757411,);
not I_44342 (I757419,I757411);
nor I_44343 (I757436,I757419,I757317);
and I_44344 (I757453,I757436,I515985);
nor I_44345 (I757470,I757419,I757385);
nor I_44346 (I757266,I757377,I757470);
DFFARX1 I_44347 (I515982,I3563,I757283,I757510,);
nor I_44348 (I757518,I757510,I757377);
not I_44349 (I757535,I757518);
not I_44350 (I757552,I757510);
nor I_44351 (I757569,I757552,I757453);
DFFARX1 I_44352 (I757569,I3563,I757283,I757269,);
nand I_44353 (I757600,I515997,I515994);
and I_44354 (I757617,I757600,I515976);
DFFARX1 I_44355 (I757617,I3563,I757283,I757643,);
nor I_44356 (I757651,I757643,I757510);
DFFARX1 I_44357 (I757651,I3563,I757283,I757251,);
nand I_44358 (I757682,I757643,I757552);
nand I_44359 (I757260,I757535,I757682);
not I_44360 (I757713,I757643);
nor I_44361 (I757730,I757713,I757453);
DFFARX1 I_44362 (I757730,I3563,I757283,I757272,);
nor I_44363 (I757761,I515970,I515994);
or I_44364 (I757263,I757510,I757761);
nor I_44365 (I757254,I757643,I757761);
or I_44366 (I757257,I757377,I757761);
DFFARX1 I_44367 (I757761,I3563,I757283,I757275,);
not I_44368 (I757861,I3570);
DFFARX1 I_44369 (I252963,I3563,I757861,I757887,);
not I_44370 (I757895,I757887);
nand I_44371 (I757912,I252966,I252987);
and I_44372 (I757929,I757912,I252975);
DFFARX1 I_44373 (I757929,I3563,I757861,I757955,);
not I_44374 (I757963,I252972);
DFFARX1 I_44375 (I252963,I3563,I757861,I757989,);
not I_44376 (I757997,I757989);
nor I_44377 (I758014,I757997,I757895);
and I_44378 (I758031,I758014,I252972);
nor I_44379 (I758048,I757997,I757963);
nor I_44380 (I757844,I757955,I758048);
DFFARX1 I_44381 (I252981,I3563,I757861,I758088,);
nor I_44382 (I758096,I758088,I757955);
not I_44383 (I758113,I758096);
not I_44384 (I758130,I758088);
nor I_44385 (I758147,I758130,I758031);
DFFARX1 I_44386 (I758147,I3563,I757861,I757847,);
nand I_44387 (I758178,I252966,I252969);
and I_44388 (I758195,I758178,I252978);
DFFARX1 I_44389 (I758195,I3563,I757861,I758221,);
nor I_44390 (I758229,I758221,I758088);
DFFARX1 I_44391 (I758229,I3563,I757861,I757829,);
nand I_44392 (I758260,I758221,I758130);
nand I_44393 (I757838,I758113,I758260);
not I_44394 (I758291,I758221);
nor I_44395 (I758308,I758291,I758031);
DFFARX1 I_44396 (I758308,I3563,I757861,I757850,);
nor I_44397 (I758339,I252984,I252969);
or I_44398 (I757841,I758088,I758339);
nor I_44399 (I757832,I758221,I758339);
or I_44400 (I757835,I757955,I758339);
DFFARX1 I_44401 (I758339,I3563,I757861,I757853,);
not I_44402 (I758439,I3570);
DFFARX1 I_44403 (I609283,I3563,I758439,I758465,);
not I_44404 (I758473,I758465);
nand I_44405 (I758490,I609292,I609301);
and I_44406 (I758507,I758490,I609307);
DFFARX1 I_44407 (I758507,I3563,I758439,I758533,);
not I_44408 (I758541,I609304);
DFFARX1 I_44409 (I609289,I3563,I758439,I758567,);
not I_44410 (I758575,I758567);
nor I_44411 (I758592,I758575,I758473);
and I_44412 (I758609,I758592,I609304);
nor I_44413 (I758626,I758575,I758541);
nor I_44414 (I758422,I758533,I758626);
DFFARX1 I_44415 (I609298,I3563,I758439,I758666,);
nor I_44416 (I758674,I758666,I758533);
not I_44417 (I758691,I758674);
not I_44418 (I758708,I758666);
nor I_44419 (I758725,I758708,I758609);
DFFARX1 I_44420 (I758725,I3563,I758439,I758425,);
nand I_44421 (I758756,I609295,I609286);
and I_44422 (I758773,I758756,I609283);
DFFARX1 I_44423 (I758773,I3563,I758439,I758799,);
nor I_44424 (I758807,I758799,I758666);
DFFARX1 I_44425 (I758807,I3563,I758439,I758407,);
nand I_44426 (I758838,I758799,I758708);
nand I_44427 (I758416,I758691,I758838);
not I_44428 (I758869,I758799);
nor I_44429 (I758886,I758869,I758609);
DFFARX1 I_44430 (I758886,I3563,I758439,I758428,);
nor I_44431 (I758917,I609286,I609286);
or I_44432 (I758419,I758666,I758917);
nor I_44433 (I758410,I758799,I758917);
or I_44434 (I758413,I758533,I758917);
DFFARX1 I_44435 (I758917,I3563,I758439,I758431,);
not I_44436 (I759017,I3570);
DFFARX1 I_44437 (I1394625,I3563,I759017,I759043,);
not I_44438 (I759051,I759043);
nand I_44439 (I759068,I1394610,I1394598);
and I_44440 (I759085,I759068,I1394613);
DFFARX1 I_44441 (I759085,I3563,I759017,I759111,);
not I_44442 (I759119,I1394598);
DFFARX1 I_44443 (I1394616,I3563,I759017,I759145,);
not I_44444 (I759153,I759145);
nor I_44445 (I759170,I759153,I759051);
and I_44446 (I759187,I759170,I1394598);
nor I_44447 (I759204,I759153,I759119);
nor I_44448 (I759000,I759111,I759204);
DFFARX1 I_44449 (I1394604,I3563,I759017,I759244,);
nor I_44450 (I759252,I759244,I759111);
not I_44451 (I759269,I759252);
not I_44452 (I759286,I759244);
nor I_44453 (I759303,I759286,I759187);
DFFARX1 I_44454 (I759303,I3563,I759017,I759003,);
nand I_44455 (I759334,I1394601,I1394607);
and I_44456 (I759351,I759334,I1394622);
DFFARX1 I_44457 (I759351,I3563,I759017,I759377,);
nor I_44458 (I759385,I759377,I759244);
DFFARX1 I_44459 (I759385,I3563,I759017,I758985,);
nand I_44460 (I759416,I759377,I759286);
nand I_44461 (I758994,I759269,I759416);
not I_44462 (I759447,I759377);
nor I_44463 (I759464,I759447,I759187);
DFFARX1 I_44464 (I759464,I3563,I759017,I759006,);
nor I_44465 (I759495,I1394619,I1394607);
or I_44466 (I758997,I759244,I759495);
nor I_44467 (I758988,I759377,I759495);
or I_44468 (I758991,I759111,I759495);
DFFARX1 I_44469 (I759495,I3563,I759017,I759009,);
not I_44470 (I759595,I3570);
DFFARX1 I_44471 (I1342265,I3563,I759595,I759621,);
not I_44472 (I759629,I759621);
nand I_44473 (I759646,I1342250,I1342238);
and I_44474 (I759663,I759646,I1342253);
DFFARX1 I_44475 (I759663,I3563,I759595,I759689,);
not I_44476 (I759697,I1342238);
DFFARX1 I_44477 (I1342256,I3563,I759595,I759723,);
not I_44478 (I759731,I759723);
nor I_44479 (I759748,I759731,I759629);
and I_44480 (I759765,I759748,I1342238);
nor I_44481 (I759782,I759731,I759697);
nor I_44482 (I759578,I759689,I759782);
DFFARX1 I_44483 (I1342244,I3563,I759595,I759822,);
nor I_44484 (I759830,I759822,I759689);
not I_44485 (I759847,I759830);
not I_44486 (I759864,I759822);
nor I_44487 (I759881,I759864,I759765);
DFFARX1 I_44488 (I759881,I3563,I759595,I759581,);
nand I_44489 (I759912,I1342241,I1342247);
and I_44490 (I759929,I759912,I1342262);
DFFARX1 I_44491 (I759929,I3563,I759595,I759955,);
nor I_44492 (I759963,I759955,I759822);
DFFARX1 I_44493 (I759963,I3563,I759595,I759563,);
nand I_44494 (I759994,I759955,I759864);
nand I_44495 (I759572,I759847,I759994);
not I_44496 (I760025,I759955);
nor I_44497 (I760042,I760025,I759765);
DFFARX1 I_44498 (I760042,I3563,I759595,I759584,);
nor I_44499 (I760073,I1342259,I1342247);
or I_44500 (I759575,I759822,I760073);
nor I_44501 (I759566,I759955,I760073);
or I_44502 (I759569,I759689,I760073);
DFFARX1 I_44503 (I760073,I3563,I759595,I759587,);
not I_44504 (I760173,I3570);
DFFARX1 I_44505 (I309104,I3563,I760173,I760199,);
not I_44506 (I760207,I760199);
nand I_44507 (I760224,I309107,I309083);
and I_44508 (I760241,I760224,I309080);
DFFARX1 I_44509 (I760241,I3563,I760173,I760267,);
not I_44510 (I760275,I309086);
DFFARX1 I_44511 (I309080,I3563,I760173,I760301,);
not I_44512 (I760309,I760301);
nor I_44513 (I760326,I760309,I760207);
and I_44514 (I760343,I760326,I309086);
nor I_44515 (I760360,I760309,I760275);
nor I_44516 (I760156,I760267,I760360);
DFFARX1 I_44517 (I309089,I3563,I760173,I760400,);
nor I_44518 (I760408,I760400,I760267);
not I_44519 (I760425,I760408);
not I_44520 (I760442,I760400);
nor I_44521 (I760459,I760442,I760343);
DFFARX1 I_44522 (I760459,I3563,I760173,I760159,);
nand I_44523 (I760490,I309092,I309101);
and I_44524 (I760507,I760490,I309098);
DFFARX1 I_44525 (I760507,I3563,I760173,I760533,);
nor I_44526 (I760541,I760533,I760400);
DFFARX1 I_44527 (I760541,I3563,I760173,I760141,);
nand I_44528 (I760572,I760533,I760442);
nand I_44529 (I760150,I760425,I760572);
not I_44530 (I760603,I760533);
nor I_44531 (I760620,I760603,I760343);
DFFARX1 I_44532 (I760620,I3563,I760173,I760162,);
nor I_44533 (I760651,I309095,I309101);
or I_44534 (I760153,I760400,I760651);
nor I_44535 (I760144,I760533,I760651);
or I_44536 (I760147,I760267,I760651);
DFFARX1 I_44537 (I760651,I3563,I760173,I760165,);
not I_44538 (I760751,I3570);
DFFARX1 I_44539 (I27674,I3563,I760751,I760777,);
not I_44540 (I760785,I760777);
nand I_44541 (I760802,I27671,I27662);
and I_44542 (I760819,I760802,I27662);
DFFARX1 I_44543 (I760819,I3563,I760751,I760845,);
not I_44544 (I760853,I27665);
DFFARX1 I_44545 (I27680,I3563,I760751,I760879,);
not I_44546 (I760887,I760879);
nor I_44547 (I760904,I760887,I760785);
and I_44548 (I760921,I760904,I27665);
nor I_44549 (I760938,I760887,I760853);
nor I_44550 (I760734,I760845,I760938);
DFFARX1 I_44551 (I27665,I3563,I760751,I760978,);
nor I_44552 (I760986,I760978,I760845);
not I_44553 (I761003,I760986);
not I_44554 (I761020,I760978);
nor I_44555 (I761037,I761020,I760921);
DFFARX1 I_44556 (I761037,I3563,I760751,I760737,);
nand I_44557 (I761068,I27683,I27668);
and I_44558 (I761085,I761068,I27686);
DFFARX1 I_44559 (I761085,I3563,I760751,I761111,);
nor I_44560 (I761119,I761111,I760978);
DFFARX1 I_44561 (I761119,I3563,I760751,I760719,);
nand I_44562 (I761150,I761111,I761020);
nand I_44563 (I760728,I761003,I761150);
not I_44564 (I761181,I761111);
nor I_44565 (I761198,I761181,I760921);
DFFARX1 I_44566 (I761198,I3563,I760751,I760740,);
nor I_44567 (I761229,I27677,I27668);
or I_44568 (I760731,I760978,I761229);
nor I_44569 (I760722,I761111,I761229);
or I_44570 (I760725,I760845,I761229);
DFFARX1 I_44571 (I761229,I3563,I760751,I760743,);
not I_44572 (I761329,I3570);
DFFARX1 I_44573 (I582695,I3563,I761329,I761355,);
not I_44574 (I761363,I761355);
nand I_44575 (I761380,I582704,I582713);
and I_44576 (I761397,I761380,I582719);
DFFARX1 I_44577 (I761397,I3563,I761329,I761423,);
not I_44578 (I761431,I582716);
DFFARX1 I_44579 (I582701,I3563,I761329,I761457,);
not I_44580 (I761465,I761457);
nor I_44581 (I761482,I761465,I761363);
and I_44582 (I761499,I761482,I582716);
nor I_44583 (I761516,I761465,I761431);
nor I_44584 (I761312,I761423,I761516);
DFFARX1 I_44585 (I582710,I3563,I761329,I761556,);
nor I_44586 (I761564,I761556,I761423);
not I_44587 (I761581,I761564);
not I_44588 (I761598,I761556);
nor I_44589 (I761615,I761598,I761499);
DFFARX1 I_44590 (I761615,I3563,I761329,I761315,);
nand I_44591 (I761646,I582707,I582698);
and I_44592 (I761663,I761646,I582695);
DFFARX1 I_44593 (I761663,I3563,I761329,I761689,);
nor I_44594 (I761697,I761689,I761556);
DFFARX1 I_44595 (I761697,I3563,I761329,I761297,);
nand I_44596 (I761728,I761689,I761598);
nand I_44597 (I761306,I761581,I761728);
not I_44598 (I761759,I761689);
nor I_44599 (I761776,I761759,I761499);
DFFARX1 I_44600 (I761776,I3563,I761329,I761318,);
nor I_44601 (I761807,I582698,I582698);
or I_44602 (I761309,I761556,I761807);
nor I_44603 (I761300,I761689,I761807);
or I_44604 (I761303,I761423,I761807);
DFFARX1 I_44605 (I761807,I3563,I761329,I761321,);
not I_44606 (I761907,I3570);
DFFARX1 I_44607 (I1176557,I3563,I761907,I761933,);
not I_44608 (I761941,I761933);
nand I_44609 (I761958,I1176539,I1176551);
and I_44610 (I761975,I761958,I1176554);
DFFARX1 I_44611 (I761975,I3563,I761907,I762001,);
not I_44612 (I762009,I1176548);
DFFARX1 I_44613 (I1176545,I3563,I761907,I762035,);
not I_44614 (I762043,I762035);
nor I_44615 (I762060,I762043,I761941);
and I_44616 (I762077,I762060,I1176548);
nor I_44617 (I762094,I762043,I762009);
nor I_44618 (I761890,I762001,I762094);
DFFARX1 I_44619 (I1176563,I3563,I761907,I762134,);
nor I_44620 (I762142,I762134,I762001);
not I_44621 (I762159,I762142);
not I_44622 (I762176,I762134);
nor I_44623 (I762193,I762176,I762077);
DFFARX1 I_44624 (I762193,I3563,I761907,I761893,);
nand I_44625 (I762224,I1176542,I1176542);
and I_44626 (I762241,I762224,I1176539);
DFFARX1 I_44627 (I762241,I3563,I761907,I762267,);
nor I_44628 (I762275,I762267,I762134);
DFFARX1 I_44629 (I762275,I3563,I761907,I761875,);
nand I_44630 (I762306,I762267,I762176);
nand I_44631 (I761884,I762159,I762306);
not I_44632 (I762337,I762267);
nor I_44633 (I762354,I762337,I762077);
DFFARX1 I_44634 (I762354,I3563,I761907,I761896,);
nor I_44635 (I762385,I1176560,I1176542);
or I_44636 (I761887,I762134,I762385);
nor I_44637 (I761878,I762267,I762385);
or I_44638 (I761881,I762001,I762385);
DFFARX1 I_44639 (I762385,I3563,I761907,I761899,);
not I_44640 (I762485,I3570);
DFFARX1 I_44641 (I641651,I3563,I762485,I762511,);
not I_44642 (I762519,I762511);
nand I_44643 (I762536,I641660,I641669);
and I_44644 (I762553,I762536,I641675);
DFFARX1 I_44645 (I762553,I3563,I762485,I762579,);
not I_44646 (I762587,I641672);
DFFARX1 I_44647 (I641657,I3563,I762485,I762613,);
not I_44648 (I762621,I762613);
nor I_44649 (I762638,I762621,I762519);
and I_44650 (I762655,I762638,I641672);
nor I_44651 (I762672,I762621,I762587);
nor I_44652 (I762468,I762579,I762672);
DFFARX1 I_44653 (I641666,I3563,I762485,I762712,);
nor I_44654 (I762720,I762712,I762579);
not I_44655 (I762737,I762720);
not I_44656 (I762754,I762712);
nor I_44657 (I762771,I762754,I762655);
DFFARX1 I_44658 (I762771,I3563,I762485,I762471,);
nand I_44659 (I762802,I641663,I641654);
and I_44660 (I762819,I762802,I641651);
DFFARX1 I_44661 (I762819,I3563,I762485,I762845,);
nor I_44662 (I762853,I762845,I762712);
DFFARX1 I_44663 (I762853,I3563,I762485,I762453,);
nand I_44664 (I762884,I762845,I762754);
nand I_44665 (I762462,I762737,I762884);
not I_44666 (I762915,I762845);
nor I_44667 (I762932,I762915,I762655);
DFFARX1 I_44668 (I762932,I3563,I762485,I762474,);
nor I_44669 (I762963,I641654,I641654);
or I_44670 (I762465,I762712,I762963);
nor I_44671 (I762456,I762845,I762963);
or I_44672 (I762459,I762579,I762963);
DFFARX1 I_44673 (I762963,I3563,I762485,I762477,);
not I_44674 (I763063,I3570);
DFFARX1 I_44675 (I386573,I3563,I763063,I763089,);
not I_44676 (I763097,I763089);
nand I_44677 (I763114,I386576,I386552);
and I_44678 (I763131,I763114,I386549);
DFFARX1 I_44679 (I763131,I3563,I763063,I763157,);
not I_44680 (I763165,I386555);
DFFARX1 I_44681 (I386549,I3563,I763063,I763191,);
not I_44682 (I763199,I763191);
nor I_44683 (I763216,I763199,I763097);
and I_44684 (I763233,I763216,I386555);
nor I_44685 (I763250,I763199,I763165);
nor I_44686 (I763046,I763157,I763250);
DFFARX1 I_44687 (I386558,I3563,I763063,I763290,);
nor I_44688 (I763298,I763290,I763157);
not I_44689 (I763315,I763298);
not I_44690 (I763332,I763290);
nor I_44691 (I763349,I763332,I763233);
DFFARX1 I_44692 (I763349,I3563,I763063,I763049,);
nand I_44693 (I763380,I386561,I386570);
and I_44694 (I763397,I763380,I386567);
DFFARX1 I_44695 (I763397,I3563,I763063,I763423,);
nor I_44696 (I763431,I763423,I763290);
DFFARX1 I_44697 (I763431,I3563,I763063,I763031,);
nand I_44698 (I763462,I763423,I763332);
nand I_44699 (I763040,I763315,I763462);
not I_44700 (I763493,I763423);
nor I_44701 (I763510,I763493,I763233);
DFFARX1 I_44702 (I763510,I3563,I763063,I763052,);
nor I_44703 (I763541,I386564,I386570);
or I_44704 (I763043,I763290,I763541);
nor I_44705 (I763034,I763423,I763541);
or I_44706 (I763037,I763157,I763541);
DFFARX1 I_44707 (I763541,I3563,I763063,I763055,);
not I_44708 (I763641,I3570);
DFFARX1 I_44709 (I1155749,I3563,I763641,I763667,);
not I_44710 (I763675,I763667);
nand I_44711 (I763692,I1155731,I1155743);
and I_44712 (I763709,I763692,I1155746);
DFFARX1 I_44713 (I763709,I3563,I763641,I763735,);
not I_44714 (I763743,I1155740);
DFFARX1 I_44715 (I1155737,I3563,I763641,I763769,);
not I_44716 (I763777,I763769);
nor I_44717 (I763794,I763777,I763675);
and I_44718 (I763811,I763794,I1155740);
nor I_44719 (I763828,I763777,I763743);
nor I_44720 (I763624,I763735,I763828);
DFFARX1 I_44721 (I1155755,I3563,I763641,I763868,);
nor I_44722 (I763876,I763868,I763735);
not I_44723 (I763893,I763876);
not I_44724 (I763910,I763868);
nor I_44725 (I763927,I763910,I763811);
DFFARX1 I_44726 (I763927,I3563,I763641,I763627,);
nand I_44727 (I763958,I1155734,I1155734);
and I_44728 (I763975,I763958,I1155731);
DFFARX1 I_44729 (I763975,I3563,I763641,I764001,);
nor I_44730 (I764009,I764001,I763868);
DFFARX1 I_44731 (I764009,I3563,I763641,I763609,);
nand I_44732 (I764040,I764001,I763910);
nand I_44733 (I763618,I763893,I764040);
not I_44734 (I764071,I764001);
nor I_44735 (I764088,I764071,I763811);
DFFARX1 I_44736 (I764088,I3563,I763641,I763630,);
nor I_44737 (I764119,I1155752,I1155734);
or I_44738 (I763621,I763868,I764119);
nor I_44739 (I763612,I764001,I764119);
or I_44740 (I763615,I763735,I764119);
DFFARX1 I_44741 (I764119,I3563,I763641,I763633,);
not I_44742 (I764219,I3570);
DFFARX1 I_44743 (I1304515,I3563,I764219,I764245,);
not I_44744 (I764253,I764245);
nand I_44745 (I764270,I1304539,I1304521);
and I_44746 (I764287,I764270,I1304527);
DFFARX1 I_44747 (I764287,I3563,I764219,I764313,);
not I_44748 (I764321,I1304533);
DFFARX1 I_44749 (I1304518,I3563,I764219,I764347,);
not I_44750 (I764355,I764347);
nor I_44751 (I764372,I764355,I764253);
and I_44752 (I764389,I764372,I1304533);
nor I_44753 (I764406,I764355,I764321);
nor I_44754 (I764202,I764313,I764406);
DFFARX1 I_44755 (I1304530,I3563,I764219,I764446,);
nor I_44756 (I764454,I764446,I764313);
not I_44757 (I764471,I764454);
not I_44758 (I764488,I764446);
nor I_44759 (I764505,I764488,I764389);
DFFARX1 I_44760 (I764505,I3563,I764219,I764205,);
nand I_44761 (I764536,I1304536,I1304524);
and I_44762 (I764553,I764536,I1304518);
DFFARX1 I_44763 (I764553,I3563,I764219,I764579,);
nor I_44764 (I764587,I764579,I764446);
DFFARX1 I_44765 (I764587,I3563,I764219,I764187,);
nand I_44766 (I764618,I764579,I764488);
nand I_44767 (I764196,I764471,I764618);
not I_44768 (I764649,I764579);
nor I_44769 (I764666,I764649,I764389);
DFFARX1 I_44770 (I764666,I3563,I764219,I764208,);
nor I_44771 (I764697,I1304515,I1304524);
or I_44772 (I764199,I764446,I764697);
nor I_44773 (I764190,I764579,I764697);
or I_44774 (I764193,I764313,I764697);
DFFARX1 I_44775 (I764697,I3563,I764219,I764211,);
not I_44776 (I764797,I3570);
DFFARX1 I_44777 (I192868,I3563,I764797,I764823,);
not I_44778 (I764831,I764823);
nand I_44779 (I764848,I192871,I192892);
and I_44780 (I764865,I764848,I192880);
DFFARX1 I_44781 (I764865,I3563,I764797,I764891,);
not I_44782 (I764899,I192877);
DFFARX1 I_44783 (I192868,I3563,I764797,I764925,);
not I_44784 (I764933,I764925);
nor I_44785 (I764950,I764933,I764831);
and I_44786 (I764967,I764950,I192877);
nor I_44787 (I764984,I764933,I764899);
nor I_44788 (I764780,I764891,I764984);
DFFARX1 I_44789 (I192886,I3563,I764797,I765024,);
nor I_44790 (I765032,I765024,I764891);
not I_44791 (I765049,I765032);
not I_44792 (I765066,I765024);
nor I_44793 (I765083,I765066,I764967);
DFFARX1 I_44794 (I765083,I3563,I764797,I764783,);
nand I_44795 (I765114,I192871,I192874);
and I_44796 (I765131,I765114,I192883);
DFFARX1 I_44797 (I765131,I3563,I764797,I765157,);
nor I_44798 (I765165,I765157,I765024);
DFFARX1 I_44799 (I765165,I3563,I764797,I764765,);
nand I_44800 (I765196,I765157,I765066);
nand I_44801 (I764774,I765049,I765196);
not I_44802 (I765227,I765157);
nor I_44803 (I765244,I765227,I764967);
DFFARX1 I_44804 (I765244,I3563,I764797,I764786,);
nor I_44805 (I765275,I192889,I192874);
or I_44806 (I764777,I765024,I765275);
nor I_44807 (I764768,I765157,I765275);
or I_44808 (I764771,I764891,I765275);
DFFARX1 I_44809 (I765275,I3563,I764797,I764789,);
not I_44810 (I765375,I3570);
DFFARX1 I_44811 (I221428,I3563,I765375,I765401,);
not I_44812 (I765409,I765401);
nand I_44813 (I765426,I221431,I221452);
and I_44814 (I765443,I765426,I221440);
DFFARX1 I_44815 (I765443,I3563,I765375,I765469,);
not I_44816 (I765477,I221437);
DFFARX1 I_44817 (I221428,I3563,I765375,I765503,);
not I_44818 (I765511,I765503);
nor I_44819 (I765528,I765511,I765409);
and I_44820 (I765545,I765528,I221437);
nor I_44821 (I765562,I765511,I765477);
nor I_44822 (I765358,I765469,I765562);
DFFARX1 I_44823 (I221446,I3563,I765375,I765602,);
nor I_44824 (I765610,I765602,I765469);
not I_44825 (I765627,I765610);
not I_44826 (I765644,I765602);
nor I_44827 (I765661,I765644,I765545);
DFFARX1 I_44828 (I765661,I3563,I765375,I765361,);
nand I_44829 (I765692,I221431,I221434);
and I_44830 (I765709,I765692,I221443);
DFFARX1 I_44831 (I765709,I3563,I765375,I765735,);
nor I_44832 (I765743,I765735,I765602);
DFFARX1 I_44833 (I765743,I3563,I765375,I765343,);
nand I_44834 (I765774,I765735,I765644);
nand I_44835 (I765352,I765627,I765774);
not I_44836 (I765805,I765735);
nor I_44837 (I765822,I765805,I765545);
DFFARX1 I_44838 (I765822,I3563,I765375,I765364,);
nor I_44839 (I765853,I221449,I221434);
or I_44840 (I765355,I765602,I765853);
nor I_44841 (I765346,I765735,I765853);
or I_44842 (I765349,I765469,I765853);
DFFARX1 I_44843 (I765853,I3563,I765375,I765367,);
not I_44844 (I765953,I3570);
DFFARX1 I_44845 (I1106619,I3563,I765953,I765979,);
not I_44846 (I765987,I765979);
nand I_44847 (I766004,I1106601,I1106613);
and I_44848 (I766021,I766004,I1106616);
DFFARX1 I_44849 (I766021,I3563,I765953,I766047,);
not I_44850 (I766055,I1106610);
DFFARX1 I_44851 (I1106607,I3563,I765953,I766081,);
not I_44852 (I766089,I766081);
nor I_44853 (I766106,I766089,I765987);
and I_44854 (I766123,I766106,I1106610);
nor I_44855 (I766140,I766089,I766055);
nor I_44856 (I765936,I766047,I766140);
DFFARX1 I_44857 (I1106625,I3563,I765953,I766180,);
nor I_44858 (I766188,I766180,I766047);
not I_44859 (I766205,I766188);
not I_44860 (I766222,I766180);
nor I_44861 (I766239,I766222,I766123);
DFFARX1 I_44862 (I766239,I3563,I765953,I765939,);
nand I_44863 (I766270,I1106604,I1106604);
and I_44864 (I766287,I766270,I1106601);
DFFARX1 I_44865 (I766287,I3563,I765953,I766313,);
nor I_44866 (I766321,I766313,I766180);
DFFARX1 I_44867 (I766321,I3563,I765953,I765921,);
nand I_44868 (I766352,I766313,I766222);
nand I_44869 (I765930,I766205,I766352);
not I_44870 (I766383,I766313);
nor I_44871 (I766400,I766383,I766123);
DFFARX1 I_44872 (I766400,I3563,I765953,I765942,);
nor I_44873 (I766431,I1106622,I1106604);
or I_44874 (I765933,I766180,I766431);
nor I_44875 (I765924,I766313,I766431);
or I_44876 (I765927,I766047,I766431);
DFFARX1 I_44877 (I766431,I3563,I765953,I765945,);
not I_44878 (I766531,I3570);
DFFARX1 I_44879 (I481707,I3563,I766531,I766557,);
not I_44880 (I766565,I766557);
nand I_44881 (I766582,I481698,I481716);
and I_44882 (I766599,I766582,I481719);
DFFARX1 I_44883 (I766599,I3563,I766531,I766625,);
not I_44884 (I766633,I481713);
DFFARX1 I_44885 (I481701,I3563,I766531,I766659,);
not I_44886 (I766667,I766659);
nor I_44887 (I766684,I766667,I766565);
and I_44888 (I766701,I766684,I481713);
nor I_44889 (I766718,I766667,I766633);
nor I_44890 (I766514,I766625,I766718);
DFFARX1 I_44891 (I481710,I3563,I766531,I766758,);
nor I_44892 (I766766,I766758,I766625);
not I_44893 (I766783,I766766);
not I_44894 (I766800,I766758);
nor I_44895 (I766817,I766800,I766701);
DFFARX1 I_44896 (I766817,I3563,I766531,I766517,);
nand I_44897 (I766848,I481725,I481722);
and I_44898 (I766865,I766848,I481704);
DFFARX1 I_44899 (I766865,I3563,I766531,I766891,);
nor I_44900 (I766899,I766891,I766758);
DFFARX1 I_44901 (I766899,I3563,I766531,I766499,);
nand I_44902 (I766930,I766891,I766800);
nand I_44903 (I766508,I766783,I766930);
not I_44904 (I766961,I766891);
nor I_44905 (I766978,I766961,I766701);
DFFARX1 I_44906 (I766978,I3563,I766531,I766520,);
nor I_44907 (I767009,I481698,I481722);
or I_44908 (I766511,I766758,I767009);
nor I_44909 (I766502,I766891,I767009);
or I_44910 (I766505,I766625,I767009);
DFFARX1 I_44911 (I767009,I3563,I766531,I766523,);
not I_44912 (I767109,I3570);
DFFARX1 I_44913 (I350737,I3563,I767109,I767135,);
not I_44914 (I767143,I767135);
nand I_44915 (I767160,I350740,I350716);
and I_44916 (I767177,I767160,I350713);
DFFARX1 I_44917 (I767177,I3563,I767109,I767203,);
not I_44918 (I767211,I350719);
DFFARX1 I_44919 (I350713,I3563,I767109,I767237,);
not I_44920 (I767245,I767237);
nor I_44921 (I767262,I767245,I767143);
and I_44922 (I767279,I767262,I350719);
nor I_44923 (I767296,I767245,I767211);
nor I_44924 (I767092,I767203,I767296);
DFFARX1 I_44925 (I350722,I3563,I767109,I767336,);
nor I_44926 (I767344,I767336,I767203);
not I_44927 (I767361,I767344);
not I_44928 (I767378,I767336);
nor I_44929 (I767395,I767378,I767279);
DFFARX1 I_44930 (I767395,I3563,I767109,I767095,);
nand I_44931 (I767426,I350725,I350734);
and I_44932 (I767443,I767426,I350731);
DFFARX1 I_44933 (I767443,I3563,I767109,I767469,);
nor I_44934 (I767477,I767469,I767336);
DFFARX1 I_44935 (I767477,I3563,I767109,I767077,);
nand I_44936 (I767508,I767469,I767378);
nand I_44937 (I767086,I767361,I767508);
not I_44938 (I767539,I767469);
nor I_44939 (I767556,I767539,I767279);
DFFARX1 I_44940 (I767556,I3563,I767109,I767098,);
nor I_44941 (I767587,I350728,I350734);
or I_44942 (I767089,I767336,I767587);
nor I_44943 (I767080,I767469,I767587);
or I_44944 (I767083,I767203,I767587);
DFFARX1 I_44945 (I767587,I3563,I767109,I767101,);
not I_44946 (I767687,I3570);
DFFARX1 I_44947 (I1312607,I3563,I767687,I767713,);
not I_44948 (I767721,I767713);
nand I_44949 (I767738,I1312631,I1312613);
and I_44950 (I767755,I767738,I1312619);
DFFARX1 I_44951 (I767755,I3563,I767687,I767781,);
not I_44952 (I767789,I1312625);
DFFARX1 I_44953 (I1312610,I3563,I767687,I767815,);
not I_44954 (I767823,I767815);
nor I_44955 (I767840,I767823,I767721);
and I_44956 (I767857,I767840,I1312625);
nor I_44957 (I767874,I767823,I767789);
nor I_44958 (I767670,I767781,I767874);
DFFARX1 I_44959 (I1312622,I3563,I767687,I767914,);
nor I_44960 (I767922,I767914,I767781);
not I_44961 (I767939,I767922);
not I_44962 (I767956,I767914);
nor I_44963 (I767973,I767956,I767857);
DFFARX1 I_44964 (I767973,I3563,I767687,I767673,);
nand I_44965 (I768004,I1312628,I1312616);
and I_44966 (I768021,I768004,I1312610);
DFFARX1 I_44967 (I768021,I3563,I767687,I768047,);
nor I_44968 (I768055,I768047,I767914);
DFFARX1 I_44969 (I768055,I3563,I767687,I767655,);
nand I_44970 (I768086,I768047,I767956);
nand I_44971 (I767664,I767939,I768086);
not I_44972 (I768117,I768047);
nor I_44973 (I768134,I768117,I767857);
DFFARX1 I_44974 (I768134,I3563,I767687,I767676,);
nor I_44975 (I768165,I1312607,I1312616);
or I_44976 (I767667,I767914,I768165);
nor I_44977 (I767658,I768047,I768165);
or I_44978 (I767661,I767781,I768165);
DFFARX1 I_44979 (I768165,I3563,I767687,I767679,);
not I_44980 (I768265,I3570);
DFFARX1 I_44981 (I596567,I3563,I768265,I768291,);
not I_44982 (I768299,I768291);
nand I_44983 (I768316,I596576,I596585);
and I_44984 (I768333,I768316,I596591);
DFFARX1 I_44985 (I768333,I3563,I768265,I768359,);
not I_44986 (I768367,I596588);
DFFARX1 I_44987 (I596573,I3563,I768265,I768393,);
not I_44988 (I768401,I768393);
nor I_44989 (I768418,I768401,I768299);
and I_44990 (I768435,I768418,I596588);
nor I_44991 (I768452,I768401,I768367);
nor I_44992 (I768248,I768359,I768452);
DFFARX1 I_44993 (I596582,I3563,I768265,I768492,);
nor I_44994 (I768500,I768492,I768359);
not I_44995 (I768517,I768500);
not I_44996 (I768534,I768492);
nor I_44997 (I768551,I768534,I768435);
DFFARX1 I_44998 (I768551,I3563,I768265,I768251,);
nand I_44999 (I768582,I596579,I596570);
and I_45000 (I768599,I768582,I596567);
DFFARX1 I_45001 (I768599,I3563,I768265,I768625,);
nor I_45002 (I768633,I768625,I768492);
DFFARX1 I_45003 (I768633,I3563,I768265,I768233,);
nand I_45004 (I768664,I768625,I768534);
nand I_45005 (I768242,I768517,I768664);
not I_45006 (I768695,I768625);
nor I_45007 (I768712,I768695,I768435);
DFFARX1 I_45008 (I768712,I3563,I768265,I768254,);
nor I_45009 (I768743,I596570,I596570);
or I_45010 (I768245,I768492,I768743);
nor I_45011 (I768236,I768625,I768743);
or I_45012 (I768239,I768359,I768743);
DFFARX1 I_45013 (I768743,I3563,I768265,I768257,);
not I_45014 (I768843,I3570);
DFFARX1 I_45015 (I532851,I3563,I768843,I768869,);
not I_45016 (I768877,I768869);
nand I_45017 (I768894,I532866,I532851);
and I_45018 (I768911,I768894,I532854);
DFFARX1 I_45019 (I768911,I3563,I768843,I768937,);
not I_45020 (I768945,I532854);
DFFARX1 I_45021 (I532863,I3563,I768843,I768971,);
not I_45022 (I768979,I768971);
nor I_45023 (I768996,I768979,I768877);
and I_45024 (I769013,I768996,I532854);
nor I_45025 (I769030,I768979,I768945);
nor I_45026 (I768826,I768937,I769030);
DFFARX1 I_45027 (I532857,I3563,I768843,I769070,);
nor I_45028 (I769078,I769070,I768937);
not I_45029 (I769095,I769078);
not I_45030 (I769112,I769070);
nor I_45031 (I769129,I769112,I769013);
DFFARX1 I_45032 (I769129,I3563,I768843,I768829,);
nand I_45033 (I769160,I532860,I532869);
and I_45034 (I769177,I769160,I532875);
DFFARX1 I_45035 (I769177,I3563,I768843,I769203,);
nor I_45036 (I769211,I769203,I769070);
DFFARX1 I_45037 (I769211,I3563,I768843,I768811,);
nand I_45038 (I769242,I769203,I769112);
nand I_45039 (I768820,I769095,I769242);
not I_45040 (I769273,I769203);
nor I_45041 (I769290,I769273,I769013);
DFFARX1 I_45042 (I769290,I3563,I768843,I768832,);
nor I_45043 (I769321,I532872,I532869);
or I_45044 (I768823,I769070,I769321);
nor I_45045 (I768814,I769203,I769321);
or I_45046 (I768817,I768937,I769321);
DFFARX1 I_45047 (I769321,I3563,I768843,I768835,);
not I_45048 (I769421,I3570);
DFFARX1 I_45049 (I1379155,I3563,I769421,I769447,);
not I_45050 (I769455,I769447);
nand I_45051 (I769472,I1379140,I1379128);
and I_45052 (I769489,I769472,I1379143);
DFFARX1 I_45053 (I769489,I3563,I769421,I769515,);
not I_45054 (I769523,I1379128);
DFFARX1 I_45055 (I1379146,I3563,I769421,I769549,);
not I_45056 (I769557,I769549);
nor I_45057 (I769574,I769557,I769455);
and I_45058 (I769591,I769574,I1379128);
nor I_45059 (I769608,I769557,I769523);
nor I_45060 (I769404,I769515,I769608);
DFFARX1 I_45061 (I1379134,I3563,I769421,I769648,);
nor I_45062 (I769656,I769648,I769515);
not I_45063 (I769673,I769656);
not I_45064 (I769690,I769648);
nor I_45065 (I769707,I769690,I769591);
DFFARX1 I_45066 (I769707,I3563,I769421,I769407,);
nand I_45067 (I769738,I1379131,I1379137);
and I_45068 (I769755,I769738,I1379152);
DFFARX1 I_45069 (I769755,I3563,I769421,I769781,);
nor I_45070 (I769789,I769781,I769648);
DFFARX1 I_45071 (I769789,I3563,I769421,I769389,);
nand I_45072 (I769820,I769781,I769690);
nand I_45073 (I769398,I769673,I769820);
not I_45074 (I769851,I769781);
nor I_45075 (I769868,I769851,I769591);
DFFARX1 I_45076 (I769868,I3563,I769421,I769410,);
nor I_45077 (I769899,I1379149,I1379137);
or I_45078 (I769401,I769648,I769899);
nor I_45079 (I769392,I769781,I769899);
or I_45080 (I769395,I769515,I769899);
DFFARX1 I_45081 (I769899,I3563,I769421,I769413,);
not I_45082 (I769999,I3570);
DFFARX1 I_45083 (I1392840,I3563,I769999,I770025,);
not I_45084 (I770033,I770025);
nand I_45085 (I770050,I1392825,I1392813);
and I_45086 (I770067,I770050,I1392828);
DFFARX1 I_45087 (I770067,I3563,I769999,I770093,);
not I_45088 (I770101,I1392813);
DFFARX1 I_45089 (I1392831,I3563,I769999,I770127,);
not I_45090 (I770135,I770127);
nor I_45091 (I770152,I770135,I770033);
and I_45092 (I770169,I770152,I1392813);
nor I_45093 (I770186,I770135,I770101);
nor I_45094 (I769982,I770093,I770186);
DFFARX1 I_45095 (I1392819,I3563,I769999,I770226,);
nor I_45096 (I770234,I770226,I770093);
not I_45097 (I770251,I770234);
not I_45098 (I770268,I770226);
nor I_45099 (I770285,I770268,I770169);
DFFARX1 I_45100 (I770285,I3563,I769999,I769985,);
nand I_45101 (I770316,I1392816,I1392822);
and I_45102 (I770333,I770316,I1392837);
DFFARX1 I_45103 (I770333,I3563,I769999,I770359,);
nor I_45104 (I770367,I770359,I770226);
DFFARX1 I_45105 (I770367,I3563,I769999,I769967,);
nand I_45106 (I770398,I770359,I770268);
nand I_45107 (I769976,I770251,I770398);
not I_45108 (I770429,I770359);
nor I_45109 (I770446,I770429,I770169);
DFFARX1 I_45110 (I770446,I3563,I769999,I769988,);
nor I_45111 (I770477,I1392834,I1392822);
or I_45112 (I769979,I770226,I770477);
nor I_45113 (I769970,I770359,I770477);
or I_45114 (I769973,I770093,I770477);
DFFARX1 I_45115 (I770477,I3563,I769999,I769991,);
not I_45116 (I770577,I3570);
DFFARX1 I_45117 (I1280137,I3563,I770577,I770603,);
not I_45118 (I770611,I770603);
nand I_45119 (I770628,I1280140,I1280149);
and I_45120 (I770645,I770628,I1280152);
DFFARX1 I_45121 (I770645,I3563,I770577,I770671,);
not I_45122 (I770679,I1280161);
DFFARX1 I_45123 (I1280143,I3563,I770577,I770705,);
not I_45124 (I770713,I770705);
nor I_45125 (I770730,I770713,I770611);
and I_45126 (I770747,I770730,I1280161);
nor I_45127 (I770764,I770713,I770679);
nor I_45128 (I770560,I770671,I770764);
DFFARX1 I_45129 (I1280140,I3563,I770577,I770804,);
nor I_45130 (I770812,I770804,I770671);
not I_45131 (I770829,I770812);
not I_45132 (I770846,I770804);
nor I_45133 (I770863,I770846,I770747);
DFFARX1 I_45134 (I770863,I3563,I770577,I770563,);
nand I_45135 (I770894,I1280158,I1280137);
and I_45136 (I770911,I770894,I1280155);
DFFARX1 I_45137 (I770911,I3563,I770577,I770937,);
nor I_45138 (I770945,I770937,I770804);
DFFARX1 I_45139 (I770945,I3563,I770577,I770545,);
nand I_45140 (I770976,I770937,I770846);
nand I_45141 (I770554,I770829,I770976);
not I_45142 (I771007,I770937);
nor I_45143 (I771024,I771007,I770747);
DFFARX1 I_45144 (I771024,I3563,I770577,I770566,);
nor I_45145 (I771055,I1280146,I1280137);
or I_45146 (I770557,I770804,I771055);
nor I_45147 (I770548,I770937,I771055);
or I_45148 (I770551,I770671,I771055);
DFFARX1 I_45149 (I771055,I3563,I770577,I770569,);
not I_45150 (I771155,I3570);
DFFARX1 I_45151 (I13694,I3563,I771155,I771181,);
not I_45152 (I771189,I771181);
nand I_45153 (I771206,I13697,I13709);
and I_45154 (I771223,I771206,I13688);
DFFARX1 I_45155 (I771223,I3563,I771155,I771249,);
not I_45156 (I771257,I13688);
DFFARX1 I_45157 (I13691,I3563,I771155,I771283,);
not I_45158 (I771291,I771283);
nor I_45159 (I771308,I771291,I771189);
and I_45160 (I771325,I771308,I13688);
nor I_45161 (I771342,I771291,I771257);
nor I_45162 (I771138,I771249,I771342);
DFFARX1 I_45163 (I13703,I3563,I771155,I771382,);
nor I_45164 (I771390,I771382,I771249);
not I_45165 (I771407,I771390);
not I_45166 (I771424,I771382);
nor I_45167 (I771441,I771424,I771325);
DFFARX1 I_45168 (I771441,I3563,I771155,I771141,);
nand I_45169 (I771472,I13706,I13691);
and I_45170 (I771489,I771472,I13700);
DFFARX1 I_45171 (I771489,I3563,I771155,I771515,);
nor I_45172 (I771523,I771515,I771382);
DFFARX1 I_45173 (I771523,I3563,I771155,I771123,);
nand I_45174 (I771554,I771515,I771424);
nand I_45175 (I771132,I771407,I771554);
not I_45176 (I771585,I771515);
nor I_45177 (I771602,I771585,I771325);
DFFARX1 I_45178 (I771602,I3563,I771155,I771144,);
nor I_45179 (I771633,I13694,I13691);
or I_45180 (I771135,I771382,I771633);
nor I_45181 (I771126,I771515,I771633);
or I_45182 (I771129,I771249,I771633);
DFFARX1 I_45183 (I771633,I3563,I771155,I771147,);
not I_45184 (I771733,I3570);
DFFARX1 I_45185 (I1288331,I3563,I771733,I771759,);
not I_45186 (I771767,I771759);
nand I_45187 (I771784,I1288355,I1288337);
and I_45188 (I771801,I771784,I1288343);
DFFARX1 I_45189 (I771801,I3563,I771733,I771827,);
not I_45190 (I771835,I1288349);
DFFARX1 I_45191 (I1288334,I3563,I771733,I771861,);
not I_45192 (I771869,I771861);
nor I_45193 (I771886,I771869,I771767);
and I_45194 (I771903,I771886,I1288349);
nor I_45195 (I771920,I771869,I771835);
nor I_45196 (I771716,I771827,I771920);
DFFARX1 I_45197 (I1288346,I3563,I771733,I771960,);
nor I_45198 (I771968,I771960,I771827);
not I_45199 (I771985,I771968);
not I_45200 (I772002,I771960);
nor I_45201 (I772019,I772002,I771903);
DFFARX1 I_45202 (I772019,I3563,I771733,I771719,);
nand I_45203 (I772050,I1288352,I1288340);
and I_45204 (I772067,I772050,I1288334);
DFFARX1 I_45205 (I772067,I3563,I771733,I772093,);
nor I_45206 (I772101,I772093,I771960);
DFFARX1 I_45207 (I772101,I3563,I771733,I771701,);
nand I_45208 (I772132,I772093,I772002);
nand I_45209 (I771710,I771985,I772132);
not I_45210 (I772163,I772093);
nor I_45211 (I772180,I772163,I771903);
DFFARX1 I_45212 (I772180,I3563,I771733,I771722,);
nor I_45213 (I772211,I1288331,I1288340);
or I_45214 (I771713,I771960,I772211);
nor I_45215 (I771704,I772093,I772211);
or I_45216 (I771707,I771827,I772211);
DFFARX1 I_45217 (I772211,I3563,I771733,I771725,);
not I_45218 (I772311,I3570);
DFFARX1 I_45219 (I110404,I3563,I772311,I772337,);
not I_45220 (I772345,I772337);
nand I_45221 (I772362,I110413,I110422);
and I_45222 (I772379,I772362,I110401);
DFFARX1 I_45223 (I772379,I3563,I772311,I772405,);
not I_45224 (I772413,I110404);
DFFARX1 I_45225 (I110419,I3563,I772311,I772439,);
not I_45226 (I772447,I772439);
nor I_45227 (I772464,I772447,I772345);
and I_45228 (I772481,I772464,I110404);
nor I_45229 (I772498,I772447,I772413);
nor I_45230 (I772294,I772405,I772498);
DFFARX1 I_45231 (I110410,I3563,I772311,I772538,);
nor I_45232 (I772546,I772538,I772405);
not I_45233 (I772563,I772546);
not I_45234 (I772580,I772538);
nor I_45235 (I772597,I772580,I772481);
DFFARX1 I_45236 (I772597,I3563,I772311,I772297,);
nand I_45237 (I772628,I110425,I110401);
and I_45238 (I772645,I772628,I110407);
DFFARX1 I_45239 (I772645,I3563,I772311,I772671,);
nor I_45240 (I772679,I772671,I772538);
DFFARX1 I_45241 (I772679,I3563,I772311,I772279,);
nand I_45242 (I772710,I772671,I772580);
nand I_45243 (I772288,I772563,I772710);
not I_45244 (I772741,I772671);
nor I_45245 (I772758,I772741,I772481);
DFFARX1 I_45246 (I772758,I3563,I772311,I772300,);
nor I_45247 (I772789,I110416,I110401);
or I_45248 (I772291,I772538,I772789);
nor I_45249 (I772282,I772671,I772789);
or I_45250 (I772285,I772405,I772789);
DFFARX1 I_45251 (I772789,I3563,I772311,I772303,);
not I_45252 (I772889,I3570);
DFFARX1 I_45253 (I1080886,I3563,I772889,I772915,);
not I_45254 (I772923,I772915);
nand I_45255 (I772940,I1080883,I1080901);
and I_45256 (I772957,I772940,I1080898);
DFFARX1 I_45257 (I772957,I3563,I772889,I772983,);
not I_45258 (I772991,I1080880);
DFFARX1 I_45259 (I1080883,I3563,I772889,I773017,);
not I_45260 (I773025,I773017);
nor I_45261 (I773042,I773025,I772923);
and I_45262 (I773059,I773042,I1080880);
nor I_45263 (I773076,I773025,I772991);
nor I_45264 (I772872,I772983,I773076);
DFFARX1 I_45265 (I1080892,I3563,I772889,I773116,);
nor I_45266 (I773124,I773116,I772983);
not I_45267 (I773141,I773124);
not I_45268 (I773158,I773116);
nor I_45269 (I773175,I773158,I773059);
DFFARX1 I_45270 (I773175,I3563,I772889,I772875,);
nand I_45271 (I773206,I1080895,I1080880);
and I_45272 (I773223,I773206,I1080886);
DFFARX1 I_45273 (I773223,I3563,I772889,I773249,);
nor I_45274 (I773257,I773249,I773116);
DFFARX1 I_45275 (I773257,I3563,I772889,I772857,);
nand I_45276 (I773288,I773249,I773158);
nand I_45277 (I772866,I773141,I773288);
not I_45278 (I773319,I773249);
nor I_45279 (I773336,I773319,I773059);
DFFARX1 I_45280 (I773336,I3563,I772889,I772878,);
nor I_45281 (I773367,I1080889,I1080880);
or I_45282 (I772869,I773116,I773367);
nor I_45283 (I772860,I773249,I773367);
or I_45284 (I772863,I772983,I773367);
DFFARX1 I_45285 (I773367,I3563,I772889,I772881,);
not I_45286 (I773467,I3570);
DFFARX1 I_45287 (I1309139,I3563,I773467,I773493,);
not I_45288 (I773501,I773493);
nand I_45289 (I773518,I1309163,I1309145);
and I_45290 (I773535,I773518,I1309151);
DFFARX1 I_45291 (I773535,I3563,I773467,I773561,);
not I_45292 (I773569,I1309157);
DFFARX1 I_45293 (I1309142,I3563,I773467,I773595,);
not I_45294 (I773603,I773595);
nor I_45295 (I773620,I773603,I773501);
and I_45296 (I773637,I773620,I1309157);
nor I_45297 (I773654,I773603,I773569);
nor I_45298 (I773450,I773561,I773654);
DFFARX1 I_45299 (I1309154,I3563,I773467,I773694,);
nor I_45300 (I773702,I773694,I773561);
not I_45301 (I773719,I773702);
not I_45302 (I773736,I773694);
nor I_45303 (I773753,I773736,I773637);
DFFARX1 I_45304 (I773753,I3563,I773467,I773453,);
nand I_45305 (I773784,I1309160,I1309148);
and I_45306 (I773801,I773784,I1309142);
DFFARX1 I_45307 (I773801,I3563,I773467,I773827,);
nor I_45308 (I773835,I773827,I773694);
DFFARX1 I_45309 (I773835,I3563,I773467,I773435,);
nand I_45310 (I773866,I773827,I773736);
nand I_45311 (I773444,I773719,I773866);
not I_45312 (I773897,I773827);
nor I_45313 (I773914,I773897,I773637);
DFFARX1 I_45314 (I773914,I3563,I773467,I773456,);
nor I_45315 (I773945,I1309139,I1309148);
or I_45316 (I773447,I773694,I773945);
nor I_45317 (I773438,I773827,I773945);
or I_45318 (I773441,I773561,I773945);
DFFARX1 I_45319 (I773945,I3563,I773467,I773459,);
not I_45320 (I774045,I3570);
DFFARX1 I_45321 (I159560,I3563,I774045,I774071,);
not I_45322 (I774079,I774071);
nand I_45323 (I774096,I159575,I159548);
and I_45324 (I774113,I774096,I159563);
DFFARX1 I_45325 (I774113,I3563,I774045,I774139,);
not I_45326 (I774147,I159566);
DFFARX1 I_45327 (I159551,I3563,I774045,I774173,);
not I_45328 (I774181,I774173);
nor I_45329 (I774198,I774181,I774079);
and I_45330 (I774215,I774198,I159566);
nor I_45331 (I774232,I774181,I774147);
nor I_45332 (I774028,I774139,I774232);
DFFARX1 I_45333 (I159557,I3563,I774045,I774272,);
nor I_45334 (I774280,I774272,I774139);
not I_45335 (I774297,I774280);
not I_45336 (I774314,I774272);
nor I_45337 (I774331,I774314,I774215);
DFFARX1 I_45338 (I774331,I3563,I774045,I774031,);
nand I_45339 (I774362,I159572,I159554);
and I_45340 (I774379,I774362,I159569);
DFFARX1 I_45341 (I774379,I3563,I774045,I774405,);
nor I_45342 (I774413,I774405,I774272);
DFFARX1 I_45343 (I774413,I3563,I774045,I774013,);
nand I_45344 (I774444,I774405,I774314);
nand I_45345 (I774022,I774297,I774444);
not I_45346 (I774475,I774405);
nor I_45347 (I774492,I774475,I774215);
DFFARX1 I_45348 (I774492,I3563,I774045,I774034,);
nor I_45349 (I774523,I159548,I159554);
or I_45350 (I774025,I774272,I774523);
nor I_45351 (I774016,I774405,I774523);
or I_45352 (I774019,I774139,I774523);
DFFARX1 I_45353 (I774523,I3563,I774045,I774037,);
not I_45354 (I774623,I3570);
DFFARX1 I_45355 (I912782,I3563,I774623,I774649,);
not I_45356 (I774657,I774649);
nand I_45357 (I774674,I912770,I912788);
and I_45358 (I774691,I774674,I912785);
DFFARX1 I_45359 (I774691,I3563,I774623,I774717,);
not I_45360 (I774725,I912776);
DFFARX1 I_45361 (I912773,I3563,I774623,I774751,);
not I_45362 (I774759,I774751);
nor I_45363 (I774776,I774759,I774657);
and I_45364 (I774793,I774776,I912776);
nor I_45365 (I774810,I774759,I774725);
nor I_45366 (I774606,I774717,I774810);
DFFARX1 I_45367 (I912767,I3563,I774623,I774850,);
nor I_45368 (I774858,I774850,I774717);
not I_45369 (I774875,I774858);
not I_45370 (I774892,I774850);
nor I_45371 (I774909,I774892,I774793);
DFFARX1 I_45372 (I774909,I3563,I774623,I774609,);
nand I_45373 (I774940,I912767,I912770);
and I_45374 (I774957,I774940,I912773);
DFFARX1 I_45375 (I774957,I3563,I774623,I774983,);
nor I_45376 (I774991,I774983,I774850);
DFFARX1 I_45377 (I774991,I3563,I774623,I774591,);
nand I_45378 (I775022,I774983,I774892);
nand I_45379 (I774600,I774875,I775022);
not I_45380 (I775053,I774983);
nor I_45381 (I775070,I775053,I774793);
DFFARX1 I_45382 (I775070,I3563,I774623,I774612,);
nor I_45383 (I775101,I912779,I912770);
or I_45384 (I774603,I774850,I775101);
nor I_45385 (I774594,I774983,I775101);
or I_45386 (I774597,I774717,I775101);
DFFARX1 I_45387 (I775101,I3563,I774623,I774615,);
not I_45388 (I775201,I3570);
DFFARX1 I_45389 (I283308,I3563,I775201,I775227,);
not I_45390 (I775235,I775227);
nand I_45391 (I775252,I283311,I283332);
and I_45392 (I775269,I775252,I283320);
DFFARX1 I_45393 (I775269,I3563,I775201,I775295,);
not I_45394 (I775303,I283317);
DFFARX1 I_45395 (I283308,I3563,I775201,I775329,);
not I_45396 (I775337,I775329);
nor I_45397 (I775354,I775337,I775235);
and I_45398 (I775371,I775354,I283317);
nor I_45399 (I775388,I775337,I775303);
nor I_45400 (I775184,I775295,I775388);
DFFARX1 I_45401 (I283326,I3563,I775201,I775428,);
nor I_45402 (I775436,I775428,I775295);
not I_45403 (I775453,I775436);
not I_45404 (I775470,I775428);
nor I_45405 (I775487,I775470,I775371);
DFFARX1 I_45406 (I775487,I3563,I775201,I775187,);
nand I_45407 (I775518,I283311,I283314);
and I_45408 (I775535,I775518,I283323);
DFFARX1 I_45409 (I775535,I3563,I775201,I775561,);
nor I_45410 (I775569,I775561,I775428);
DFFARX1 I_45411 (I775569,I3563,I775201,I775169,);
nand I_45412 (I775600,I775561,I775470);
nand I_45413 (I775178,I775453,I775600);
not I_45414 (I775631,I775561);
nor I_45415 (I775648,I775631,I775371);
DFFARX1 I_45416 (I775648,I3563,I775201,I775190,);
nor I_45417 (I775679,I283329,I283314);
or I_45418 (I775181,I775428,I775679);
nor I_45419 (I775172,I775561,I775679);
or I_45420 (I775175,I775295,I775679);
DFFARX1 I_45421 (I775679,I3563,I775201,I775193,);
not I_45422 (I775779,I3570);
DFFARX1 I_45423 (I91432,I3563,I775779,I775805,);
not I_45424 (I775813,I775805);
nand I_45425 (I775830,I91441,I91450);
and I_45426 (I775847,I775830,I91429);
DFFARX1 I_45427 (I775847,I3563,I775779,I775873,);
not I_45428 (I775881,I91432);
DFFARX1 I_45429 (I91447,I3563,I775779,I775907,);
not I_45430 (I775915,I775907);
nor I_45431 (I775932,I775915,I775813);
and I_45432 (I775949,I775932,I91432);
nor I_45433 (I775966,I775915,I775881);
nor I_45434 (I775762,I775873,I775966);
DFFARX1 I_45435 (I91438,I3563,I775779,I776006,);
nor I_45436 (I776014,I776006,I775873);
not I_45437 (I776031,I776014);
not I_45438 (I776048,I776006);
nor I_45439 (I776065,I776048,I775949);
DFFARX1 I_45440 (I776065,I3563,I775779,I775765,);
nand I_45441 (I776096,I91453,I91429);
and I_45442 (I776113,I776096,I91435);
DFFARX1 I_45443 (I776113,I3563,I775779,I776139,);
nor I_45444 (I776147,I776139,I776006);
DFFARX1 I_45445 (I776147,I3563,I775779,I775747,);
nand I_45446 (I776178,I776139,I776048);
nand I_45447 (I775756,I776031,I776178);
not I_45448 (I776209,I776139);
nor I_45449 (I776226,I776209,I775949);
DFFARX1 I_45450 (I776226,I3563,I775779,I775768,);
nor I_45451 (I776257,I91444,I91429);
or I_45452 (I775759,I776006,I776257);
nor I_45453 (I775750,I776139,I776257);
or I_45454 (I775753,I775873,I776257);
DFFARX1 I_45455 (I776257,I3563,I775779,I775771,);
not I_45456 (I776357,I3570);
DFFARX1 I_45457 (I1179447,I3563,I776357,I776383,);
not I_45458 (I776391,I776383);
nand I_45459 (I776408,I1179429,I1179441);
and I_45460 (I776425,I776408,I1179444);
DFFARX1 I_45461 (I776425,I3563,I776357,I776451,);
not I_45462 (I776459,I1179438);
DFFARX1 I_45463 (I1179435,I3563,I776357,I776485,);
not I_45464 (I776493,I776485);
nor I_45465 (I776510,I776493,I776391);
and I_45466 (I776527,I776510,I1179438);
nor I_45467 (I776544,I776493,I776459);
nor I_45468 (I776340,I776451,I776544);
DFFARX1 I_45469 (I1179453,I3563,I776357,I776584,);
nor I_45470 (I776592,I776584,I776451);
not I_45471 (I776609,I776592);
not I_45472 (I776626,I776584);
nor I_45473 (I776643,I776626,I776527);
DFFARX1 I_45474 (I776643,I3563,I776357,I776343,);
nand I_45475 (I776674,I1179432,I1179432);
and I_45476 (I776691,I776674,I1179429);
DFFARX1 I_45477 (I776691,I3563,I776357,I776717,);
nor I_45478 (I776725,I776717,I776584);
DFFARX1 I_45479 (I776725,I3563,I776357,I776325,);
nand I_45480 (I776756,I776717,I776626);
nand I_45481 (I776334,I776609,I776756);
not I_45482 (I776787,I776717);
nor I_45483 (I776804,I776787,I776527);
DFFARX1 I_45484 (I776804,I3563,I776357,I776346,);
nor I_45485 (I776835,I1179450,I1179432);
or I_45486 (I776337,I776584,I776835);
nor I_45487 (I776328,I776717,I776835);
or I_45488 (I776331,I776451,I776835);
DFFARX1 I_45489 (I776835,I3563,I776357,I776349,);
not I_45490 (I776935,I3570);
DFFARX1 I_45491 (I16080,I3563,I776935,I776961,);
not I_45492 (I776969,I776961);
nand I_45493 (I776986,I16077,I16068);
and I_45494 (I777003,I776986,I16068);
DFFARX1 I_45495 (I777003,I3563,I776935,I777029,);
not I_45496 (I777037,I16071);
DFFARX1 I_45497 (I16086,I3563,I776935,I777063,);
not I_45498 (I777071,I777063);
nor I_45499 (I777088,I777071,I776969);
and I_45500 (I777105,I777088,I16071);
nor I_45501 (I777122,I777071,I777037);
nor I_45502 (I776918,I777029,I777122);
DFFARX1 I_45503 (I16071,I3563,I776935,I777162,);
nor I_45504 (I777170,I777162,I777029);
not I_45505 (I777187,I777170);
not I_45506 (I777204,I777162);
nor I_45507 (I777221,I777204,I777105);
DFFARX1 I_45508 (I777221,I3563,I776935,I776921,);
nand I_45509 (I777252,I16089,I16074);
and I_45510 (I777269,I777252,I16092);
DFFARX1 I_45511 (I777269,I3563,I776935,I777295,);
nor I_45512 (I777303,I777295,I777162);
DFFARX1 I_45513 (I777303,I3563,I776935,I776903,);
nand I_45514 (I777334,I777295,I777204);
nand I_45515 (I776912,I777187,I777334);
not I_45516 (I777365,I777295);
nor I_45517 (I777382,I777365,I777105);
DFFARX1 I_45518 (I777382,I3563,I776935,I776924,);
nor I_45519 (I777413,I16083,I16074);
or I_45520 (I776915,I777162,I777413);
nor I_45521 (I776906,I777295,I777413);
or I_45522 (I776909,I777029,I777413);
DFFARX1 I_45523 (I777413,I3563,I776935,I776927,);
not I_45524 (I777513,I3570);
DFFARX1 I_45525 (I1375585,I3563,I777513,I777539,);
not I_45526 (I777547,I777539);
nand I_45527 (I777564,I1375570,I1375558);
and I_45528 (I777581,I777564,I1375573);
DFFARX1 I_45529 (I777581,I3563,I777513,I777607,);
not I_45530 (I777615,I1375558);
DFFARX1 I_45531 (I1375576,I3563,I777513,I777641,);
not I_45532 (I777649,I777641);
nor I_45533 (I777666,I777649,I777547);
and I_45534 (I777683,I777666,I1375558);
nor I_45535 (I777700,I777649,I777615);
nor I_45536 (I777496,I777607,I777700);
DFFARX1 I_45537 (I1375564,I3563,I777513,I777740,);
nor I_45538 (I777748,I777740,I777607);
not I_45539 (I777765,I777748);
not I_45540 (I777782,I777740);
nor I_45541 (I777799,I777782,I777683);
DFFARX1 I_45542 (I777799,I3563,I777513,I777499,);
nand I_45543 (I777830,I1375561,I1375567);
and I_45544 (I777847,I777830,I1375582);
DFFARX1 I_45545 (I777847,I3563,I777513,I777873,);
nor I_45546 (I777881,I777873,I777740);
DFFARX1 I_45547 (I777881,I3563,I777513,I777481,);
nand I_45548 (I777912,I777873,I777782);
nand I_45549 (I777490,I777765,I777912);
not I_45550 (I777943,I777873);
nor I_45551 (I777960,I777943,I777683);
DFFARX1 I_45552 (I777960,I3563,I777513,I777502,);
nor I_45553 (I777991,I1375579,I1375567);
or I_45554 (I777493,I777740,I777991);
nor I_45555 (I777484,I777873,I777991);
or I_45556 (I777487,I777607,I777991);
DFFARX1 I_45557 (I777991,I3563,I777513,I777505,);
not I_45558 (I778091,I3570);
DFFARX1 I_45559 (I374979,I3563,I778091,I778117,);
not I_45560 (I778125,I778117);
nand I_45561 (I778142,I374982,I374958);
and I_45562 (I778159,I778142,I374955);
DFFARX1 I_45563 (I778159,I3563,I778091,I778185,);
not I_45564 (I778193,I374961);
DFFARX1 I_45565 (I374955,I3563,I778091,I778219,);
not I_45566 (I778227,I778219);
nor I_45567 (I778244,I778227,I778125);
and I_45568 (I778261,I778244,I374961);
nor I_45569 (I778278,I778227,I778193);
nor I_45570 (I778074,I778185,I778278);
DFFARX1 I_45571 (I374964,I3563,I778091,I778318,);
nor I_45572 (I778326,I778318,I778185);
not I_45573 (I778343,I778326);
not I_45574 (I778360,I778318);
nor I_45575 (I778377,I778360,I778261);
DFFARX1 I_45576 (I778377,I3563,I778091,I778077,);
nand I_45577 (I778408,I374967,I374976);
and I_45578 (I778425,I778408,I374973);
DFFARX1 I_45579 (I778425,I3563,I778091,I778451,);
nor I_45580 (I778459,I778451,I778318);
DFFARX1 I_45581 (I778459,I3563,I778091,I778059,);
nand I_45582 (I778490,I778451,I778360);
nand I_45583 (I778068,I778343,I778490);
not I_45584 (I778521,I778451);
nor I_45585 (I778538,I778521,I778261);
DFFARX1 I_45586 (I778538,I3563,I778091,I778080,);
nor I_45587 (I778569,I374970,I374976);
or I_45588 (I778071,I778318,I778569);
nor I_45589 (I778062,I778451,I778569);
or I_45590 (I778065,I778185,I778569);
DFFARX1 I_45591 (I778569,I3563,I778091,I778083,);
not I_45592 (I778669,I3570);
DFFARX1 I_45593 (I1326987,I3563,I778669,I778695,);
not I_45594 (I778703,I778695);
nand I_45595 (I778720,I1326975,I1326993);
and I_45596 (I778737,I778720,I1326984);
DFFARX1 I_45597 (I778737,I3563,I778669,I778763,);
not I_45598 (I778771,I1326999);
DFFARX1 I_45599 (I1326996,I3563,I778669,I778797,);
not I_45600 (I778805,I778797);
nor I_45601 (I778822,I778805,I778703);
and I_45602 (I778839,I778822,I1326999);
nor I_45603 (I778856,I778805,I778771);
nor I_45604 (I778652,I778763,I778856);
DFFARX1 I_45605 (I1326978,I3563,I778669,I778896,);
nor I_45606 (I778904,I778896,I778763);
not I_45607 (I778921,I778904);
not I_45608 (I778938,I778896);
nor I_45609 (I778955,I778938,I778839);
DFFARX1 I_45610 (I778955,I3563,I778669,I778655,);
nand I_45611 (I778986,I1326972,I1326972);
and I_45612 (I779003,I778986,I1326981);
DFFARX1 I_45613 (I779003,I3563,I778669,I779029,);
nor I_45614 (I779037,I779029,I778896);
DFFARX1 I_45615 (I779037,I3563,I778669,I778637,);
nand I_45616 (I779068,I779029,I778938);
nand I_45617 (I778646,I778921,I779068);
not I_45618 (I779099,I779029);
nor I_45619 (I779116,I779099,I778839);
DFFARX1 I_45620 (I779116,I3563,I778669,I778658,);
nor I_45621 (I779147,I1326990,I1326972);
or I_45622 (I778649,I778896,I779147);
nor I_45623 (I778640,I779029,I779147);
or I_45624 (I778643,I778763,I779147);
DFFARX1 I_45625 (I779147,I3563,I778669,I778661,);
not I_45626 (I779247,I3570);
DFFARX1 I_45627 (I204173,I3563,I779247,I779273,);
not I_45628 (I779281,I779273);
nand I_45629 (I779298,I204176,I204197);
and I_45630 (I779315,I779298,I204185);
DFFARX1 I_45631 (I779315,I3563,I779247,I779341,);
not I_45632 (I779349,I204182);
DFFARX1 I_45633 (I204173,I3563,I779247,I779375,);
not I_45634 (I779383,I779375);
nor I_45635 (I779400,I779383,I779281);
and I_45636 (I779417,I779400,I204182);
nor I_45637 (I779434,I779383,I779349);
nor I_45638 (I779230,I779341,I779434);
DFFARX1 I_45639 (I204191,I3563,I779247,I779474,);
nor I_45640 (I779482,I779474,I779341);
not I_45641 (I779499,I779482);
not I_45642 (I779516,I779474);
nor I_45643 (I779533,I779516,I779417);
DFFARX1 I_45644 (I779533,I3563,I779247,I779233,);
nand I_45645 (I779564,I204176,I204179);
and I_45646 (I779581,I779564,I204188);
DFFARX1 I_45647 (I779581,I3563,I779247,I779607,);
nor I_45648 (I779615,I779607,I779474);
DFFARX1 I_45649 (I779615,I3563,I779247,I779215,);
nand I_45650 (I779646,I779607,I779516);
nand I_45651 (I779224,I779499,I779646);
not I_45652 (I779677,I779607);
nor I_45653 (I779694,I779677,I779417);
DFFARX1 I_45654 (I779694,I3563,I779247,I779236,);
nor I_45655 (I779725,I204194,I204179);
or I_45656 (I779227,I779474,I779725);
nor I_45657 (I779218,I779607,I779725);
or I_45658 (I779221,I779341,I779725);
DFFARX1 I_45659 (I779725,I3563,I779247,I779239,);
not I_45660 (I779825,I3570);
DFFARX1 I_45661 (I866933,I3563,I779825,I779851,);
not I_45662 (I779859,I779851);
nand I_45663 (I779876,I866921,I866939);
and I_45664 (I779893,I779876,I866936);
DFFARX1 I_45665 (I779893,I3563,I779825,I779919,);
not I_45666 (I779927,I866927);
DFFARX1 I_45667 (I866924,I3563,I779825,I779953,);
not I_45668 (I779961,I779953);
nor I_45669 (I779978,I779961,I779859);
and I_45670 (I779995,I779978,I866927);
nor I_45671 (I780012,I779961,I779927);
nor I_45672 (I779808,I779919,I780012);
DFFARX1 I_45673 (I866918,I3563,I779825,I780052,);
nor I_45674 (I780060,I780052,I779919);
not I_45675 (I780077,I780060);
not I_45676 (I780094,I780052);
nor I_45677 (I780111,I780094,I779995);
DFFARX1 I_45678 (I780111,I3563,I779825,I779811,);
nand I_45679 (I780142,I866918,I866921);
and I_45680 (I780159,I780142,I866924);
DFFARX1 I_45681 (I780159,I3563,I779825,I780185,);
nor I_45682 (I780193,I780185,I780052);
DFFARX1 I_45683 (I780193,I3563,I779825,I779793,);
nand I_45684 (I780224,I780185,I780094);
nand I_45685 (I779802,I780077,I780224);
not I_45686 (I780255,I780185);
nor I_45687 (I780272,I780255,I779995);
DFFARX1 I_45688 (I780272,I3563,I779825,I779814,);
nor I_45689 (I780303,I866930,I866921);
or I_45690 (I779805,I780052,I780303);
nor I_45691 (I779796,I780185,I780303);
or I_45692 (I779799,I779919,I780303);
DFFARX1 I_45693 (I780303,I3563,I779825,I779817,);
not I_45694 (I780403,I3570);
DFFARX1 I_45695 (I1302203,I3563,I780403,I780429,);
not I_45696 (I780437,I780429);
nand I_45697 (I780454,I1302227,I1302209);
and I_45698 (I780471,I780454,I1302215);
DFFARX1 I_45699 (I780471,I3563,I780403,I780497,);
not I_45700 (I780505,I1302221);
DFFARX1 I_45701 (I1302206,I3563,I780403,I780531,);
not I_45702 (I780539,I780531);
nor I_45703 (I780556,I780539,I780437);
and I_45704 (I780573,I780556,I1302221);
nor I_45705 (I780590,I780539,I780505);
nor I_45706 (I780386,I780497,I780590);
DFFARX1 I_45707 (I1302218,I3563,I780403,I780630,);
nor I_45708 (I780638,I780630,I780497);
not I_45709 (I780655,I780638);
not I_45710 (I780672,I780630);
nor I_45711 (I780689,I780672,I780573);
DFFARX1 I_45712 (I780689,I3563,I780403,I780389,);
nand I_45713 (I780720,I1302224,I1302212);
and I_45714 (I780737,I780720,I1302206);
DFFARX1 I_45715 (I780737,I3563,I780403,I780763,);
nor I_45716 (I780771,I780763,I780630);
DFFARX1 I_45717 (I780771,I3563,I780403,I780371,);
nand I_45718 (I780802,I780763,I780672);
nand I_45719 (I780380,I780655,I780802);
not I_45720 (I780833,I780763);
nor I_45721 (I780850,I780833,I780573);
DFFARX1 I_45722 (I780850,I3563,I780403,I780392,);
nor I_45723 (I780881,I1302203,I1302212);
or I_45724 (I780383,I780630,I780881);
nor I_45725 (I780374,I780763,I780881);
or I_45726 (I780377,I780497,I780881);
DFFARX1 I_45727 (I780881,I3563,I780403,I780395,);
not I_45728 (I780981,I3570);
DFFARX1 I_45729 (I1285577,I3563,I780981,I781007,);
not I_45730 (I781015,I781007);
nand I_45731 (I781032,I1285580,I1285589);
and I_45732 (I781049,I781032,I1285592);
DFFARX1 I_45733 (I781049,I3563,I780981,I781075,);
not I_45734 (I781083,I1285601);
DFFARX1 I_45735 (I1285583,I3563,I780981,I781109,);
not I_45736 (I781117,I781109);
nor I_45737 (I781134,I781117,I781015);
and I_45738 (I781151,I781134,I1285601);
nor I_45739 (I781168,I781117,I781083);
nor I_45740 (I780964,I781075,I781168);
DFFARX1 I_45741 (I1285580,I3563,I780981,I781208,);
nor I_45742 (I781216,I781208,I781075);
not I_45743 (I781233,I781216);
not I_45744 (I781250,I781208);
nor I_45745 (I781267,I781250,I781151);
DFFARX1 I_45746 (I781267,I3563,I780981,I780967,);
nand I_45747 (I781298,I1285598,I1285577);
and I_45748 (I781315,I781298,I1285595);
DFFARX1 I_45749 (I781315,I3563,I780981,I781341,);
nor I_45750 (I781349,I781341,I781208);
DFFARX1 I_45751 (I781349,I3563,I780981,I780949,);
nand I_45752 (I781380,I781341,I781250);
nand I_45753 (I780958,I781233,I781380);
not I_45754 (I781411,I781341);
nor I_45755 (I781428,I781411,I781151);
DFFARX1 I_45756 (I781428,I3563,I780981,I780970,);
nor I_45757 (I781459,I1285586,I1285577);
or I_45758 (I780961,I781208,I781459);
nor I_45759 (I780952,I781341,I781459);
or I_45760 (I780955,I781075,I781459);
DFFARX1 I_45761 (I781459,I3563,I780981,I780973,);
not I_45762 (I781559,I3570);
DFFARX1 I_45763 (I846380,I3563,I781559,I781585,);
not I_45764 (I781593,I781585);
nand I_45765 (I781610,I846368,I846386);
and I_45766 (I781627,I781610,I846383);
DFFARX1 I_45767 (I781627,I3563,I781559,I781653,);
not I_45768 (I781661,I846374);
DFFARX1 I_45769 (I846371,I3563,I781559,I781687,);
not I_45770 (I781695,I781687);
nor I_45771 (I781712,I781695,I781593);
and I_45772 (I781729,I781712,I846374);
nor I_45773 (I781746,I781695,I781661);
nor I_45774 (I781542,I781653,I781746);
DFFARX1 I_45775 (I846365,I3563,I781559,I781786,);
nor I_45776 (I781794,I781786,I781653);
not I_45777 (I781811,I781794);
not I_45778 (I781828,I781786);
nor I_45779 (I781845,I781828,I781729);
DFFARX1 I_45780 (I781845,I3563,I781559,I781545,);
nand I_45781 (I781876,I846365,I846368);
and I_45782 (I781893,I781876,I846371);
DFFARX1 I_45783 (I781893,I3563,I781559,I781919,);
nor I_45784 (I781927,I781919,I781786);
DFFARX1 I_45785 (I781927,I3563,I781559,I781527,);
nand I_45786 (I781958,I781919,I781828);
nand I_45787 (I781536,I781811,I781958);
not I_45788 (I781989,I781919);
nor I_45789 (I782006,I781989,I781729);
DFFARX1 I_45790 (I782006,I3563,I781559,I781548,);
nor I_45791 (I782037,I846377,I846368);
or I_45792 (I781539,I781786,I782037);
nor I_45793 (I781530,I781919,I782037);
or I_45794 (I781533,I781653,I782037);
DFFARX1 I_45795 (I782037,I3563,I781559,I781551,);
not I_45796 (I782137,I3570);
DFFARX1 I_45797 (I470827,I3563,I782137,I782163,);
not I_45798 (I782171,I782163);
nand I_45799 (I782188,I470818,I470836);
and I_45800 (I782205,I782188,I470839);
DFFARX1 I_45801 (I782205,I3563,I782137,I782231,);
not I_45802 (I782239,I470833);
DFFARX1 I_45803 (I470821,I3563,I782137,I782265,);
not I_45804 (I782273,I782265);
nor I_45805 (I782290,I782273,I782171);
and I_45806 (I782307,I782290,I470833);
nor I_45807 (I782324,I782273,I782239);
nor I_45808 (I782120,I782231,I782324);
DFFARX1 I_45809 (I470830,I3563,I782137,I782364,);
nor I_45810 (I782372,I782364,I782231);
not I_45811 (I782389,I782372);
not I_45812 (I782406,I782364);
nor I_45813 (I782423,I782406,I782307);
DFFARX1 I_45814 (I782423,I3563,I782137,I782123,);
nand I_45815 (I782454,I470845,I470842);
and I_45816 (I782471,I782454,I470824);
DFFARX1 I_45817 (I782471,I3563,I782137,I782497,);
nor I_45818 (I782505,I782497,I782364);
DFFARX1 I_45819 (I782505,I3563,I782137,I782105,);
nand I_45820 (I782536,I782497,I782406);
nand I_45821 (I782114,I782389,I782536);
not I_45822 (I782567,I782497);
nor I_45823 (I782584,I782567,I782307);
DFFARX1 I_45824 (I782584,I3563,I782137,I782126,);
nor I_45825 (I782615,I470818,I470842);
or I_45826 (I782117,I782364,I782615);
nor I_45827 (I782108,I782497,I782615);
or I_45828 (I782111,I782231,I782615);
DFFARX1 I_45829 (I782615,I3563,I782137,I782129,);
not I_45830 (I782715,I3570);
DFFARX1 I_45831 (I197033,I3563,I782715,I782741,);
not I_45832 (I782749,I782741);
nand I_45833 (I782766,I197036,I197057);
and I_45834 (I782783,I782766,I197045);
DFFARX1 I_45835 (I782783,I3563,I782715,I782809,);
not I_45836 (I782817,I197042);
DFFARX1 I_45837 (I197033,I3563,I782715,I782843,);
not I_45838 (I782851,I782843);
nor I_45839 (I782868,I782851,I782749);
and I_45840 (I782885,I782868,I197042);
nor I_45841 (I782902,I782851,I782817);
nor I_45842 (I782698,I782809,I782902);
DFFARX1 I_45843 (I197051,I3563,I782715,I782942,);
nor I_45844 (I782950,I782942,I782809);
not I_45845 (I782967,I782950);
not I_45846 (I782984,I782942);
nor I_45847 (I783001,I782984,I782885);
DFFARX1 I_45848 (I783001,I3563,I782715,I782701,);
nand I_45849 (I783032,I197036,I197039);
and I_45850 (I783049,I783032,I197048);
DFFARX1 I_45851 (I783049,I3563,I782715,I783075,);
nor I_45852 (I783083,I783075,I782942);
DFFARX1 I_45853 (I783083,I3563,I782715,I782683,);
nand I_45854 (I783114,I783075,I782984);
nand I_45855 (I782692,I782967,I783114);
not I_45856 (I783145,I783075);
nor I_45857 (I783162,I783145,I782885);
DFFARX1 I_45858 (I783162,I3563,I782715,I782704,);
nor I_45859 (I783193,I197054,I197039);
or I_45860 (I782695,I782942,I783193);
nor I_45861 (I782686,I783075,I783193);
or I_45862 (I782689,I782809,I783193);
DFFARX1 I_45863 (I783193,I3563,I782715,I782707,);
not I_45864 (I783293,I3570);
DFFARX1 I_45865 (I405545,I3563,I783293,I783319,);
not I_45866 (I783327,I783319);
nand I_45867 (I783344,I405548,I405524);
and I_45868 (I783361,I783344,I405521);
DFFARX1 I_45869 (I783361,I3563,I783293,I783387,);
not I_45870 (I783395,I405527);
DFFARX1 I_45871 (I405521,I3563,I783293,I783421,);
not I_45872 (I783429,I783421);
nor I_45873 (I783446,I783429,I783327);
and I_45874 (I783463,I783446,I405527);
nor I_45875 (I783480,I783429,I783395);
nor I_45876 (I783276,I783387,I783480);
DFFARX1 I_45877 (I405530,I3563,I783293,I783520,);
nor I_45878 (I783528,I783520,I783387);
not I_45879 (I783545,I783528);
not I_45880 (I783562,I783520);
nor I_45881 (I783579,I783562,I783463);
DFFARX1 I_45882 (I783579,I3563,I783293,I783279,);
nand I_45883 (I783610,I405533,I405542);
and I_45884 (I783627,I783610,I405539);
DFFARX1 I_45885 (I783627,I3563,I783293,I783653,);
nor I_45886 (I783661,I783653,I783520);
DFFARX1 I_45887 (I783661,I3563,I783293,I783261,);
nand I_45888 (I783692,I783653,I783562);
nand I_45889 (I783270,I783545,I783692);
not I_45890 (I783723,I783653);
nor I_45891 (I783740,I783723,I783463);
DFFARX1 I_45892 (I783740,I3563,I783293,I783282,);
nor I_45893 (I783771,I405536,I405542);
or I_45894 (I783273,I783520,I783771);
nor I_45895 (I783264,I783653,I783771);
or I_45896 (I783267,I783387,I783771);
DFFARX1 I_45897 (I783771,I3563,I783293,I783285,);
not I_45898 (I783871,I3570);
DFFARX1 I_45899 (I1282857,I3563,I783871,I783897,);
not I_45900 (I783905,I783897);
nand I_45901 (I783922,I1282860,I1282869);
and I_45902 (I783939,I783922,I1282872);
DFFARX1 I_45903 (I783939,I3563,I783871,I783965,);
not I_45904 (I783973,I1282881);
DFFARX1 I_45905 (I1282863,I3563,I783871,I783999,);
not I_45906 (I784007,I783999);
nor I_45907 (I784024,I784007,I783905);
and I_45908 (I784041,I784024,I1282881);
nor I_45909 (I784058,I784007,I783973);
nor I_45910 (I783854,I783965,I784058);
DFFARX1 I_45911 (I1282860,I3563,I783871,I784098,);
nor I_45912 (I784106,I784098,I783965);
not I_45913 (I784123,I784106);
not I_45914 (I784140,I784098);
nor I_45915 (I784157,I784140,I784041);
DFFARX1 I_45916 (I784157,I3563,I783871,I783857,);
nand I_45917 (I784188,I1282878,I1282857);
and I_45918 (I784205,I784188,I1282875);
DFFARX1 I_45919 (I784205,I3563,I783871,I784231,);
nor I_45920 (I784239,I784231,I784098);
DFFARX1 I_45921 (I784239,I3563,I783871,I783839,);
nand I_45922 (I784270,I784231,I784140);
nand I_45923 (I783848,I784123,I784270);
not I_45924 (I784301,I784231);
nor I_45925 (I784318,I784301,I784041);
DFFARX1 I_45926 (I784318,I3563,I783871,I783860,);
nor I_45927 (I784349,I1282866,I1282857);
or I_45928 (I783851,I784098,I784349);
nor I_45929 (I783842,I784231,I784349);
or I_45930 (I783845,I783965,I784349);
DFFARX1 I_45931 (I784349,I3563,I783871,I783863,);
not I_45932 (I784449,I3570);
DFFARX1 I_45933 (I1064617,I3563,I784449,I784475,);
not I_45934 (I784483,I784475);
nand I_45935 (I784500,I1064614,I1064632);
and I_45936 (I784517,I784500,I1064629);
DFFARX1 I_45937 (I784517,I3563,I784449,I784543,);
not I_45938 (I784551,I1064611);
DFFARX1 I_45939 (I1064614,I3563,I784449,I784577,);
not I_45940 (I784585,I784577);
nor I_45941 (I784602,I784585,I784483);
and I_45942 (I784619,I784602,I1064611);
nor I_45943 (I784636,I784585,I784551);
nor I_45944 (I784432,I784543,I784636);
DFFARX1 I_45945 (I1064623,I3563,I784449,I784676,);
nor I_45946 (I784684,I784676,I784543);
not I_45947 (I784701,I784684);
not I_45948 (I784718,I784676);
nor I_45949 (I784735,I784718,I784619);
DFFARX1 I_45950 (I784735,I3563,I784449,I784435,);
nand I_45951 (I784766,I1064626,I1064611);
and I_45952 (I784783,I784766,I1064617);
DFFARX1 I_45953 (I784783,I3563,I784449,I784809,);
nor I_45954 (I784817,I784809,I784676);
DFFARX1 I_45955 (I784817,I3563,I784449,I784417,);
nand I_45956 (I784848,I784809,I784718);
nand I_45957 (I784426,I784701,I784848);
not I_45958 (I784879,I784809);
nor I_45959 (I784896,I784879,I784619);
DFFARX1 I_45960 (I784896,I3563,I784449,I784438,);
nor I_45961 (I784927,I1064620,I1064611);
or I_45962 (I784429,I784676,I784927);
nor I_45963 (I784420,I784809,I784927);
or I_45964 (I784423,I784543,I784927);
DFFARX1 I_45965 (I784927,I3563,I784449,I784441,);
not I_45966 (I785027,I3570);
DFFARX1 I_45967 (I326495,I3563,I785027,I785053,);
not I_45968 (I785061,I785053);
nand I_45969 (I785078,I326498,I326474);
and I_45970 (I785095,I785078,I326471);
DFFARX1 I_45971 (I785095,I3563,I785027,I785121,);
not I_45972 (I785129,I326477);
DFFARX1 I_45973 (I326471,I3563,I785027,I785155,);
not I_45974 (I785163,I785155);
nor I_45975 (I785180,I785163,I785061);
and I_45976 (I785197,I785180,I326477);
nor I_45977 (I785214,I785163,I785129);
nor I_45978 (I785010,I785121,I785214);
DFFARX1 I_45979 (I326480,I3563,I785027,I785254,);
nor I_45980 (I785262,I785254,I785121);
not I_45981 (I785279,I785262);
not I_45982 (I785296,I785254);
nor I_45983 (I785313,I785296,I785197);
DFFARX1 I_45984 (I785313,I3563,I785027,I785013,);
nand I_45985 (I785344,I326483,I326492);
and I_45986 (I785361,I785344,I326489);
DFFARX1 I_45987 (I785361,I3563,I785027,I785387,);
nor I_45988 (I785395,I785387,I785254);
DFFARX1 I_45989 (I785395,I3563,I785027,I784995,);
nand I_45990 (I785426,I785387,I785296);
nand I_45991 (I785004,I785279,I785426);
not I_45992 (I785457,I785387);
nor I_45993 (I785474,I785457,I785197);
DFFARX1 I_45994 (I785474,I3563,I785027,I785016,);
nor I_45995 (I785505,I326486,I326492);
or I_45996 (I785007,I785254,I785505);
nor I_45997 (I784998,I785387,I785505);
or I_45998 (I785001,I785121,I785505);
DFFARX1 I_45999 (I785505,I3563,I785027,I785019,);
not I_46000 (I785605,I3570);
DFFARX1 I_46001 (I456683,I3563,I785605,I785631,);
not I_46002 (I785639,I785631);
nand I_46003 (I785656,I456674,I456692);
and I_46004 (I785673,I785656,I456695);
DFFARX1 I_46005 (I785673,I3563,I785605,I785699,);
not I_46006 (I785707,I456689);
DFFARX1 I_46007 (I456677,I3563,I785605,I785733,);
not I_46008 (I785741,I785733);
nor I_46009 (I785758,I785741,I785639);
and I_46010 (I785775,I785758,I456689);
nor I_46011 (I785792,I785741,I785707);
nor I_46012 (I785588,I785699,I785792);
DFFARX1 I_46013 (I456686,I3563,I785605,I785832,);
nor I_46014 (I785840,I785832,I785699);
not I_46015 (I785857,I785840);
not I_46016 (I785874,I785832);
nor I_46017 (I785891,I785874,I785775);
DFFARX1 I_46018 (I785891,I3563,I785605,I785591,);
nand I_46019 (I785922,I456701,I456698);
and I_46020 (I785939,I785922,I456680);
DFFARX1 I_46021 (I785939,I3563,I785605,I785965,);
nor I_46022 (I785973,I785965,I785832);
DFFARX1 I_46023 (I785973,I3563,I785605,I785573,);
nand I_46024 (I786004,I785965,I785874);
nand I_46025 (I785582,I785857,I786004);
not I_46026 (I786035,I785965);
nor I_46027 (I786052,I786035,I785775);
DFFARX1 I_46028 (I786052,I3563,I785605,I785594,);
nor I_46029 (I786083,I456674,I456698);
or I_46030 (I785585,I785832,I786083);
nor I_46031 (I785576,I785965,I786083);
or I_46032 (I785579,I785699,I786083);
DFFARX1 I_46033 (I786083,I3563,I785605,I785597,);
not I_46034 (I786183,I3570);
DFFARX1 I_46035 (I1073593,I3563,I786183,I786209,);
not I_46036 (I786217,I786209);
nand I_46037 (I786234,I1073590,I1073608);
and I_46038 (I786251,I786234,I1073605);
DFFARX1 I_46039 (I786251,I3563,I786183,I786277,);
not I_46040 (I786285,I1073587);
DFFARX1 I_46041 (I1073590,I3563,I786183,I786311,);
not I_46042 (I786319,I786311);
nor I_46043 (I786336,I786319,I786217);
and I_46044 (I786353,I786336,I1073587);
nor I_46045 (I786370,I786319,I786285);
nor I_46046 (I786166,I786277,I786370);
DFFARX1 I_46047 (I1073599,I3563,I786183,I786410,);
nor I_46048 (I786418,I786410,I786277);
not I_46049 (I786435,I786418);
not I_46050 (I786452,I786410);
nor I_46051 (I786469,I786452,I786353);
DFFARX1 I_46052 (I786469,I3563,I786183,I786169,);
nand I_46053 (I786500,I1073602,I1073587);
and I_46054 (I786517,I786500,I1073593);
DFFARX1 I_46055 (I786517,I3563,I786183,I786543,);
nor I_46056 (I786551,I786543,I786410);
DFFARX1 I_46057 (I786551,I3563,I786183,I786151,);
nand I_46058 (I786582,I786543,I786452);
nand I_46059 (I786160,I786435,I786582);
not I_46060 (I786613,I786543);
nor I_46061 (I786630,I786613,I786353);
DFFARX1 I_46062 (I786630,I3563,I786183,I786172,);
nor I_46063 (I786661,I1073596,I1073587);
or I_46064 (I786163,I786410,I786661);
nor I_46065 (I786154,I786543,I786661);
or I_46066 (I786157,I786277,I786661);
DFFARX1 I_46067 (I786661,I3563,I786183,I786175,);
not I_46068 (I786761,I3570);
DFFARX1 I_46069 (I291713,I3563,I786761,I786787,);
not I_46070 (I786795,I786787);
nand I_46071 (I786812,I291716,I291692);
and I_46072 (I786829,I786812,I291689);
DFFARX1 I_46073 (I786829,I3563,I786761,I786855,);
not I_46074 (I786863,I291695);
DFFARX1 I_46075 (I291689,I3563,I786761,I786889,);
not I_46076 (I786897,I786889);
nor I_46077 (I786914,I786897,I786795);
and I_46078 (I786931,I786914,I291695);
nor I_46079 (I786948,I786897,I786863);
nor I_46080 (I786744,I786855,I786948);
DFFARX1 I_46081 (I291698,I3563,I786761,I786988,);
nor I_46082 (I786996,I786988,I786855);
not I_46083 (I787013,I786996);
not I_46084 (I787030,I786988);
nor I_46085 (I787047,I787030,I786931);
DFFARX1 I_46086 (I787047,I3563,I786761,I786747,);
nand I_46087 (I787078,I291701,I291710);
and I_46088 (I787095,I787078,I291707);
DFFARX1 I_46089 (I787095,I3563,I786761,I787121,);
nor I_46090 (I787129,I787121,I786988);
DFFARX1 I_46091 (I787129,I3563,I786761,I786729,);
nand I_46092 (I787160,I787121,I787030);
nand I_46093 (I786738,I787013,I787160);
not I_46094 (I787191,I787121);
nor I_46095 (I787208,I787191,I786931);
DFFARX1 I_46096 (I787208,I3563,I786761,I786750,);
nor I_46097 (I787239,I291704,I291710);
or I_46098 (I786741,I786988,I787239);
nor I_46099 (I786732,I787121,I787239);
or I_46100 (I786735,I786855,I787239);
DFFARX1 I_46101 (I787239,I3563,I786761,I786753,);
not I_46102 (I787339,I3570);
DFFARX1 I_46103 (I1230311,I3563,I787339,I787365,);
not I_46104 (I787373,I787365);
nand I_46105 (I787390,I1230293,I1230305);
and I_46106 (I787407,I787390,I1230308);
DFFARX1 I_46107 (I787407,I3563,I787339,I787433,);
not I_46108 (I787441,I1230302);
DFFARX1 I_46109 (I1230299,I3563,I787339,I787467,);
not I_46110 (I787475,I787467);
nor I_46111 (I787492,I787475,I787373);
and I_46112 (I787509,I787492,I1230302);
nor I_46113 (I787526,I787475,I787441);
nor I_46114 (I787322,I787433,I787526);
DFFARX1 I_46115 (I1230317,I3563,I787339,I787566,);
nor I_46116 (I787574,I787566,I787433);
not I_46117 (I787591,I787574);
not I_46118 (I787608,I787566);
nor I_46119 (I787625,I787608,I787509);
DFFARX1 I_46120 (I787625,I3563,I787339,I787325,);
nand I_46121 (I787656,I1230296,I1230296);
and I_46122 (I787673,I787656,I1230293);
DFFARX1 I_46123 (I787673,I3563,I787339,I787699,);
nor I_46124 (I787707,I787699,I787566);
DFFARX1 I_46125 (I787707,I3563,I787339,I787307,);
nand I_46126 (I787738,I787699,I787608);
nand I_46127 (I787316,I787591,I787738);
not I_46128 (I787769,I787699);
nor I_46129 (I787786,I787769,I787509);
DFFARX1 I_46130 (I787786,I3563,I787339,I787328,);
nor I_46131 (I787817,I1230314,I1230296);
or I_46132 (I787319,I787566,I787817);
nor I_46133 (I787310,I787699,I787817);
or I_46134 (I787313,I787433,I787817);
DFFARX1 I_46135 (I787817,I3563,I787339,I787331,);
not I_46136 (I787917,I3570);
DFFARX1 I_46137 (I1351785,I3563,I787917,I787943,);
not I_46138 (I787951,I787943);
nand I_46139 (I787968,I1351770,I1351758);
and I_46140 (I787985,I787968,I1351773);
DFFARX1 I_46141 (I787985,I3563,I787917,I788011,);
not I_46142 (I788019,I1351758);
DFFARX1 I_46143 (I1351776,I3563,I787917,I788045,);
not I_46144 (I788053,I788045);
nor I_46145 (I788070,I788053,I787951);
and I_46146 (I788087,I788070,I1351758);
nor I_46147 (I788104,I788053,I788019);
nor I_46148 (I787900,I788011,I788104);
DFFARX1 I_46149 (I1351764,I3563,I787917,I788144,);
nor I_46150 (I788152,I788144,I788011);
not I_46151 (I788169,I788152);
not I_46152 (I788186,I788144);
nor I_46153 (I788203,I788186,I788087);
DFFARX1 I_46154 (I788203,I3563,I787917,I787903,);
nand I_46155 (I788234,I1351761,I1351767);
and I_46156 (I788251,I788234,I1351782);
DFFARX1 I_46157 (I788251,I3563,I787917,I788277,);
nor I_46158 (I788285,I788277,I788144);
DFFARX1 I_46159 (I788285,I3563,I787917,I787885,);
nand I_46160 (I788316,I788277,I788186);
nand I_46161 (I787894,I788169,I788316);
not I_46162 (I788347,I788277);
nor I_46163 (I788364,I788347,I788087);
DFFARX1 I_46164 (I788364,I3563,I787917,I787906,);
nor I_46165 (I788395,I1351779,I1351767);
or I_46166 (I787897,I788144,I788395);
nor I_46167 (I787888,I788277,I788395);
or I_46168 (I787891,I788011,I788395);
DFFARX1 I_46169 (I788395,I3563,I787917,I787909,);
not I_46170 (I788495,I3570);
DFFARX1 I_46171 (I195843,I3563,I788495,I788521,);
not I_46172 (I788529,I788521);
nand I_46173 (I788546,I195846,I195867);
and I_46174 (I788563,I788546,I195855);
DFFARX1 I_46175 (I788563,I3563,I788495,I788589,);
not I_46176 (I788597,I195852);
DFFARX1 I_46177 (I195843,I3563,I788495,I788623,);
not I_46178 (I788631,I788623);
nor I_46179 (I788648,I788631,I788529);
and I_46180 (I788665,I788648,I195852);
nor I_46181 (I788682,I788631,I788597);
nor I_46182 (I788478,I788589,I788682);
DFFARX1 I_46183 (I195861,I3563,I788495,I788722,);
nor I_46184 (I788730,I788722,I788589);
not I_46185 (I788747,I788730);
not I_46186 (I788764,I788722);
nor I_46187 (I788781,I788764,I788665);
DFFARX1 I_46188 (I788781,I3563,I788495,I788481,);
nand I_46189 (I788812,I195846,I195849);
and I_46190 (I788829,I788812,I195858);
DFFARX1 I_46191 (I788829,I3563,I788495,I788855,);
nor I_46192 (I788863,I788855,I788722);
DFFARX1 I_46193 (I788863,I3563,I788495,I788463,);
nand I_46194 (I788894,I788855,I788764);
nand I_46195 (I788472,I788747,I788894);
not I_46196 (I788925,I788855);
nor I_46197 (I788942,I788925,I788665);
DFFARX1 I_46198 (I788942,I3563,I788495,I788484,);
nor I_46199 (I788973,I195864,I195849);
or I_46200 (I788475,I788722,I788973);
nor I_46201 (I788466,I788855,I788973);
or I_46202 (I788469,I788589,I788973);
DFFARX1 I_46203 (I788973,I3563,I788495,I788487,);
not I_46204 (I789073,I3570);
DFFARX1 I_46205 (I554866,I3563,I789073,I789099,);
not I_46206 (I789107,I789099);
nand I_46207 (I789124,I554881,I554866);
and I_46208 (I789141,I789124,I554869);
DFFARX1 I_46209 (I789141,I3563,I789073,I789167,);
not I_46210 (I789175,I554869);
DFFARX1 I_46211 (I554878,I3563,I789073,I789201,);
not I_46212 (I789209,I789201);
nor I_46213 (I789226,I789209,I789107);
and I_46214 (I789243,I789226,I554869);
nor I_46215 (I789260,I789209,I789175);
nor I_46216 (I789056,I789167,I789260);
DFFARX1 I_46217 (I554872,I3563,I789073,I789300,);
nor I_46218 (I789308,I789300,I789167);
not I_46219 (I789325,I789308);
not I_46220 (I789342,I789300);
nor I_46221 (I789359,I789342,I789243);
DFFARX1 I_46222 (I789359,I3563,I789073,I789059,);
nand I_46223 (I789390,I554875,I554884);
and I_46224 (I789407,I789390,I554890);
DFFARX1 I_46225 (I789407,I3563,I789073,I789433,);
nor I_46226 (I789441,I789433,I789300);
DFFARX1 I_46227 (I789441,I3563,I789073,I789041,);
nand I_46228 (I789472,I789433,I789342);
nand I_46229 (I789050,I789325,I789472);
not I_46230 (I789503,I789433);
nor I_46231 (I789520,I789503,I789243);
DFFARX1 I_46232 (I789520,I3563,I789073,I789062,);
nor I_46233 (I789551,I554887,I554884);
or I_46234 (I789053,I789300,I789551);
nor I_46235 (I789044,I789433,I789551);
or I_46236 (I789047,I789167,I789551);
DFFARX1 I_46237 (I789551,I3563,I789073,I789065,);
not I_46238 (I789651,I3570);
DFFARX1 I_46239 (I636449,I3563,I789651,I789677,);
not I_46240 (I789685,I789677);
nand I_46241 (I789702,I636458,I636467);
and I_46242 (I789719,I789702,I636473);
DFFARX1 I_46243 (I789719,I3563,I789651,I789745,);
not I_46244 (I789753,I636470);
DFFARX1 I_46245 (I636455,I3563,I789651,I789779,);
not I_46246 (I789787,I789779);
nor I_46247 (I789804,I789787,I789685);
and I_46248 (I789821,I789804,I636470);
nor I_46249 (I789838,I789787,I789753);
nor I_46250 (I789634,I789745,I789838);
DFFARX1 I_46251 (I636464,I3563,I789651,I789878,);
nor I_46252 (I789886,I789878,I789745);
not I_46253 (I789903,I789886);
not I_46254 (I789920,I789878);
nor I_46255 (I789937,I789920,I789821);
DFFARX1 I_46256 (I789937,I3563,I789651,I789637,);
nand I_46257 (I789968,I636461,I636452);
and I_46258 (I789985,I789968,I636449);
DFFARX1 I_46259 (I789985,I3563,I789651,I790011,);
nor I_46260 (I790019,I790011,I789878);
DFFARX1 I_46261 (I790019,I3563,I789651,I789619,);
nand I_46262 (I790050,I790011,I789920);
nand I_46263 (I789628,I789903,I790050);
not I_46264 (I790081,I790011);
nor I_46265 (I790098,I790081,I789821);
DFFARX1 I_46266 (I790098,I3563,I789651,I789640,);
nor I_46267 (I790129,I636452,I636452);
or I_46268 (I789631,I789878,I790129);
nor I_46269 (I789622,I790011,I790129);
or I_46270 (I789625,I789745,I790129);
DFFARX1 I_46271 (I790129,I3563,I789651,I789643,);
not I_46272 (I790229,I3570);
DFFARX1 I_46273 (I109877,I3563,I790229,I790255,);
not I_46274 (I790263,I790255);
nand I_46275 (I790280,I109886,I109895);
and I_46276 (I790297,I790280,I109874);
DFFARX1 I_46277 (I790297,I3563,I790229,I790323,);
not I_46278 (I790331,I109877);
DFFARX1 I_46279 (I109892,I3563,I790229,I790357,);
not I_46280 (I790365,I790357);
nor I_46281 (I790382,I790365,I790263);
and I_46282 (I790399,I790382,I109877);
nor I_46283 (I790416,I790365,I790331);
nor I_46284 (I790212,I790323,I790416);
DFFARX1 I_46285 (I109883,I3563,I790229,I790456,);
nor I_46286 (I790464,I790456,I790323);
not I_46287 (I790481,I790464);
not I_46288 (I790498,I790456);
nor I_46289 (I790515,I790498,I790399);
DFFARX1 I_46290 (I790515,I3563,I790229,I790215,);
nand I_46291 (I790546,I109898,I109874);
and I_46292 (I790563,I790546,I109880);
DFFARX1 I_46293 (I790563,I3563,I790229,I790589,);
nor I_46294 (I790597,I790589,I790456);
DFFARX1 I_46295 (I790597,I3563,I790229,I790197,);
nand I_46296 (I790628,I790589,I790498);
nand I_46297 (I790206,I790481,I790628);
not I_46298 (I790659,I790589);
nor I_46299 (I790676,I790659,I790399);
DFFARX1 I_46300 (I790676,I3563,I790229,I790218,);
nor I_46301 (I790707,I109889,I109874);
or I_46302 (I790209,I790456,I790707);
nor I_46303 (I790200,I790589,I790707);
or I_46304 (I790203,I790323,I790707);
DFFARX1 I_46305 (I790707,I3563,I790229,I790221,);
not I_46306 (I790807,I3570);
DFFARX1 I_46307 (I396059,I3563,I790807,I790833,);
not I_46308 (I790841,I790833);
nand I_46309 (I790858,I396062,I396038);
and I_46310 (I790875,I790858,I396035);
DFFARX1 I_46311 (I790875,I3563,I790807,I790901,);
not I_46312 (I790909,I396041);
DFFARX1 I_46313 (I396035,I3563,I790807,I790935,);
not I_46314 (I790943,I790935);
nor I_46315 (I790960,I790943,I790841);
and I_46316 (I790977,I790960,I396041);
nor I_46317 (I790994,I790943,I790909);
nor I_46318 (I790790,I790901,I790994);
DFFARX1 I_46319 (I396044,I3563,I790807,I791034,);
nor I_46320 (I791042,I791034,I790901);
not I_46321 (I791059,I791042);
not I_46322 (I791076,I791034);
nor I_46323 (I791093,I791076,I790977);
DFFARX1 I_46324 (I791093,I3563,I790807,I790793,);
nand I_46325 (I791124,I396047,I396056);
and I_46326 (I791141,I791124,I396053);
DFFARX1 I_46327 (I791141,I3563,I790807,I791167,);
nor I_46328 (I791175,I791167,I791034);
DFFARX1 I_46329 (I791175,I3563,I790807,I790775,);
nand I_46330 (I791206,I791167,I791076);
nand I_46331 (I790784,I791059,I791206);
not I_46332 (I791237,I791167);
nor I_46333 (I791254,I791237,I790977);
DFFARX1 I_46334 (I791254,I3563,I790807,I790796,);
nor I_46335 (I791285,I396050,I396056);
or I_46336 (I790787,I791034,I791285);
nor I_46337 (I790778,I791167,I791285);
or I_46338 (I790781,I790901,I791285);
DFFARX1 I_46339 (I791285,I3563,I790807,I790799,);
not I_46340 (I791385,I3570);
DFFARX1 I_46341 (I343359,I3563,I791385,I791411,);
not I_46342 (I791419,I791411);
nand I_46343 (I791436,I343362,I343338);
and I_46344 (I791453,I791436,I343335);
DFFARX1 I_46345 (I791453,I3563,I791385,I791479,);
not I_46346 (I791487,I343341);
DFFARX1 I_46347 (I343335,I3563,I791385,I791513,);
not I_46348 (I791521,I791513);
nor I_46349 (I791538,I791521,I791419);
and I_46350 (I791555,I791538,I343341);
nor I_46351 (I791572,I791521,I791487);
nor I_46352 (I791368,I791479,I791572);
DFFARX1 I_46353 (I343344,I3563,I791385,I791612,);
nor I_46354 (I791620,I791612,I791479);
not I_46355 (I791637,I791620);
not I_46356 (I791654,I791612);
nor I_46357 (I791671,I791654,I791555);
DFFARX1 I_46358 (I791671,I3563,I791385,I791371,);
nand I_46359 (I791702,I343347,I343356);
and I_46360 (I791719,I791702,I343353);
DFFARX1 I_46361 (I791719,I3563,I791385,I791745,);
nor I_46362 (I791753,I791745,I791612);
DFFARX1 I_46363 (I791753,I3563,I791385,I791353,);
nand I_46364 (I791784,I791745,I791654);
nand I_46365 (I791362,I791637,I791784);
not I_46366 (I791815,I791745);
nor I_46367 (I791832,I791815,I791555);
DFFARX1 I_46368 (I791832,I3563,I791385,I791374,);
nor I_46369 (I791863,I343350,I343356);
or I_46370 (I791365,I791612,I791863);
nor I_46371 (I791356,I791745,I791863);
or I_46372 (I791359,I791479,I791863);
DFFARX1 I_46373 (I791863,I3563,I791385,I791377,);
not I_46374 (I791963,I3570);
DFFARX1 I_46375 (I531066,I3563,I791963,I791989,);
not I_46376 (I791997,I791989);
nand I_46377 (I792014,I531081,I531066);
and I_46378 (I792031,I792014,I531069);
DFFARX1 I_46379 (I792031,I3563,I791963,I792057,);
not I_46380 (I792065,I531069);
DFFARX1 I_46381 (I531078,I3563,I791963,I792091,);
not I_46382 (I792099,I792091);
nor I_46383 (I792116,I792099,I791997);
and I_46384 (I792133,I792116,I531069);
nor I_46385 (I792150,I792099,I792065);
nor I_46386 (I791946,I792057,I792150);
DFFARX1 I_46387 (I531072,I3563,I791963,I792190,);
nor I_46388 (I792198,I792190,I792057);
not I_46389 (I792215,I792198);
not I_46390 (I792232,I792190);
nor I_46391 (I792249,I792232,I792133);
DFFARX1 I_46392 (I792249,I3563,I791963,I791949,);
nand I_46393 (I792280,I531075,I531084);
and I_46394 (I792297,I792280,I531090);
DFFARX1 I_46395 (I792297,I3563,I791963,I792323,);
nor I_46396 (I792331,I792323,I792190);
DFFARX1 I_46397 (I792331,I3563,I791963,I791931,);
nand I_46398 (I792362,I792323,I792232);
nand I_46399 (I791940,I792215,I792362);
not I_46400 (I792393,I792323);
nor I_46401 (I792410,I792393,I792133);
DFFARX1 I_46402 (I792410,I3563,I791963,I791952,);
nor I_46403 (I792441,I531087,I531084);
or I_46404 (I791943,I792190,I792441);
nor I_46405 (I791934,I792323,I792441);
or I_46406 (I791937,I792057,I792441);
DFFARX1 I_46407 (I792441,I3563,I791963,I791955,);
not I_46408 (I792541,I3570);
DFFARX1 I_46409 (I1143611,I3563,I792541,I792567,);
not I_46410 (I792575,I792567);
nand I_46411 (I792592,I1143593,I1143605);
and I_46412 (I792609,I792592,I1143608);
DFFARX1 I_46413 (I792609,I3563,I792541,I792635,);
not I_46414 (I792643,I1143602);
DFFARX1 I_46415 (I1143599,I3563,I792541,I792669,);
not I_46416 (I792677,I792669);
nor I_46417 (I792694,I792677,I792575);
and I_46418 (I792711,I792694,I1143602);
nor I_46419 (I792728,I792677,I792643);
nor I_46420 (I792524,I792635,I792728);
DFFARX1 I_46421 (I1143617,I3563,I792541,I792768,);
nor I_46422 (I792776,I792768,I792635);
not I_46423 (I792793,I792776);
not I_46424 (I792810,I792768);
nor I_46425 (I792827,I792810,I792711);
DFFARX1 I_46426 (I792827,I3563,I792541,I792527,);
nand I_46427 (I792858,I1143596,I1143596);
and I_46428 (I792875,I792858,I1143593);
DFFARX1 I_46429 (I792875,I3563,I792541,I792901,);
nor I_46430 (I792909,I792901,I792768);
DFFARX1 I_46431 (I792909,I3563,I792541,I792509,);
nand I_46432 (I792940,I792901,I792810);
nand I_46433 (I792518,I792793,I792940);
not I_46434 (I792971,I792901);
nor I_46435 (I792988,I792971,I792711);
DFFARX1 I_46436 (I792988,I3563,I792541,I792530,);
nor I_46437 (I793019,I1143614,I1143596);
or I_46438 (I792521,I792768,I793019);
nor I_46439 (I792512,I792901,I793019);
or I_46440 (I792515,I792635,I793019);
DFFARX1 I_46441 (I793019,I3563,I792541,I792533,);
not I_46442 (I793119,I3570);
DFFARX1 I_46443 (I324387,I3563,I793119,I793145,);
not I_46444 (I793153,I793145);
nand I_46445 (I793170,I324390,I324366);
and I_46446 (I793187,I793170,I324363);
DFFARX1 I_46447 (I793187,I3563,I793119,I793213,);
not I_46448 (I793221,I324369);
DFFARX1 I_46449 (I324363,I3563,I793119,I793247,);
not I_46450 (I793255,I793247);
nor I_46451 (I793272,I793255,I793153);
and I_46452 (I793289,I793272,I324369);
nor I_46453 (I793306,I793255,I793221);
nor I_46454 (I793102,I793213,I793306);
DFFARX1 I_46455 (I324372,I3563,I793119,I793346,);
nor I_46456 (I793354,I793346,I793213);
not I_46457 (I793371,I793354);
not I_46458 (I793388,I793346);
nor I_46459 (I793405,I793388,I793289);
DFFARX1 I_46460 (I793405,I3563,I793119,I793105,);
nand I_46461 (I793436,I324375,I324384);
and I_46462 (I793453,I793436,I324381);
DFFARX1 I_46463 (I793453,I3563,I793119,I793479,);
nor I_46464 (I793487,I793479,I793346);
DFFARX1 I_46465 (I793487,I3563,I793119,I793087,);
nand I_46466 (I793518,I793479,I793388);
nand I_46467 (I793096,I793371,I793518);
not I_46468 (I793549,I793479);
nor I_46469 (I793566,I793549,I793289);
DFFARX1 I_46470 (I793566,I3563,I793119,I793108,);
nor I_46471 (I793597,I324378,I324384);
or I_46472 (I793099,I793346,I793597);
nor I_46473 (I793090,I793479,I793597);
or I_46474 (I793093,I793213,I793597);
DFFARX1 I_46475 (I793597,I3563,I793119,I793111,);
not I_46476 (I793697,I3570);
DFFARX1 I_46477 (I1189851,I3563,I793697,I793723,);
not I_46478 (I793731,I793723);
nand I_46479 (I793748,I1189833,I1189845);
and I_46480 (I793765,I793748,I1189848);
DFFARX1 I_46481 (I793765,I3563,I793697,I793791,);
not I_46482 (I793799,I1189842);
DFFARX1 I_46483 (I1189839,I3563,I793697,I793825,);
not I_46484 (I793833,I793825);
nor I_46485 (I793850,I793833,I793731);
and I_46486 (I793867,I793850,I1189842);
nor I_46487 (I793884,I793833,I793799);
nor I_46488 (I793680,I793791,I793884);
DFFARX1 I_46489 (I1189857,I3563,I793697,I793924,);
nor I_46490 (I793932,I793924,I793791);
not I_46491 (I793949,I793932);
not I_46492 (I793966,I793924);
nor I_46493 (I793983,I793966,I793867);
DFFARX1 I_46494 (I793983,I3563,I793697,I793683,);
nand I_46495 (I794014,I1189836,I1189836);
and I_46496 (I794031,I794014,I1189833);
DFFARX1 I_46497 (I794031,I3563,I793697,I794057,);
nor I_46498 (I794065,I794057,I793924);
DFFARX1 I_46499 (I794065,I3563,I793697,I793665,);
nand I_46500 (I794096,I794057,I793966);
nand I_46501 (I793674,I793949,I794096);
not I_46502 (I794127,I794057);
nor I_46503 (I794144,I794127,I793867);
DFFARX1 I_46504 (I794144,I3563,I793697,I793686,);
nor I_46505 (I794175,I1189854,I1189836);
or I_46506 (I793677,I793924,I794175);
nor I_46507 (I793668,I794057,I794175);
or I_46508 (I793671,I793791,I794175);
DFFARX1 I_46509 (I794175,I3563,I793697,I793689,);
not I_46510 (I794275,I3570);
DFFARX1 I_46511 (I1300469,I3563,I794275,I794301,);
not I_46512 (I794309,I794301);
nand I_46513 (I794326,I1300493,I1300475);
and I_46514 (I794343,I794326,I1300481);
DFFARX1 I_46515 (I794343,I3563,I794275,I794369,);
not I_46516 (I794377,I1300487);
DFFARX1 I_46517 (I1300472,I3563,I794275,I794403,);
not I_46518 (I794411,I794403);
nor I_46519 (I794428,I794411,I794309);
and I_46520 (I794445,I794428,I1300487);
nor I_46521 (I794462,I794411,I794377);
nor I_46522 (I794258,I794369,I794462);
DFFARX1 I_46523 (I1300484,I3563,I794275,I794502,);
nor I_46524 (I794510,I794502,I794369);
not I_46525 (I794527,I794510);
not I_46526 (I794544,I794502);
nor I_46527 (I794561,I794544,I794445);
DFFARX1 I_46528 (I794561,I3563,I794275,I794261,);
nand I_46529 (I794592,I1300490,I1300478);
and I_46530 (I794609,I794592,I1300472);
DFFARX1 I_46531 (I794609,I3563,I794275,I794635,);
nor I_46532 (I794643,I794635,I794502);
DFFARX1 I_46533 (I794643,I3563,I794275,I794243,);
nand I_46534 (I794674,I794635,I794544);
nand I_46535 (I794252,I794527,I794674);
not I_46536 (I794705,I794635);
nor I_46537 (I794722,I794705,I794445);
DFFARX1 I_46538 (I794722,I3563,I794275,I794264,);
nor I_46539 (I794753,I1300469,I1300478);
or I_46540 (I794255,I794502,I794753);
nor I_46541 (I794246,I794635,I794753);
or I_46542 (I794249,I794369,I794753);
DFFARX1 I_46543 (I794753,I3563,I794275,I794267,);
not I_46544 (I794853,I3570);
DFFARX1 I_46545 (I533446,I3563,I794853,I794879,);
not I_46546 (I794887,I794879);
nand I_46547 (I794904,I533461,I533446);
and I_46548 (I794921,I794904,I533449);
DFFARX1 I_46549 (I794921,I3563,I794853,I794947,);
not I_46550 (I794955,I533449);
DFFARX1 I_46551 (I533458,I3563,I794853,I794981,);
not I_46552 (I794989,I794981);
nor I_46553 (I795006,I794989,I794887);
and I_46554 (I795023,I795006,I533449);
nor I_46555 (I795040,I794989,I794955);
nor I_46556 (I794836,I794947,I795040);
DFFARX1 I_46557 (I533452,I3563,I794853,I795080,);
nor I_46558 (I795088,I795080,I794947);
not I_46559 (I795105,I795088);
not I_46560 (I795122,I795080);
nor I_46561 (I795139,I795122,I795023);
DFFARX1 I_46562 (I795139,I3563,I794853,I794839,);
nand I_46563 (I795170,I533455,I533464);
and I_46564 (I795187,I795170,I533470);
DFFARX1 I_46565 (I795187,I3563,I794853,I795213,);
nor I_46566 (I795221,I795213,I795080);
DFFARX1 I_46567 (I795221,I3563,I794853,I794821,);
nand I_46568 (I795252,I795213,I795122);
nand I_46569 (I794830,I795105,I795252);
not I_46570 (I795283,I795213);
nor I_46571 (I795300,I795283,I795023);
DFFARX1 I_46572 (I795300,I3563,I794853,I794842,);
nor I_46573 (I795331,I533467,I533464);
or I_46574 (I794833,I795080,I795331);
nor I_46575 (I794824,I795213,I795331);
or I_46576 (I794827,I794947,I795331);
DFFARX1 I_46577 (I795331,I3563,I794853,I794845,);
not I_46578 (I795431,I3570);
DFFARX1 I_46579 (I563196,I3563,I795431,I795457,);
not I_46580 (I795465,I795457);
nand I_46581 (I795482,I563211,I563196);
and I_46582 (I795499,I795482,I563199);
DFFARX1 I_46583 (I795499,I3563,I795431,I795525,);
not I_46584 (I795533,I563199);
DFFARX1 I_46585 (I563208,I3563,I795431,I795559,);
not I_46586 (I795567,I795559);
nor I_46587 (I795584,I795567,I795465);
and I_46588 (I795601,I795584,I563199);
nor I_46589 (I795618,I795567,I795533);
nor I_46590 (I795414,I795525,I795618);
DFFARX1 I_46591 (I563202,I3563,I795431,I795658,);
nor I_46592 (I795666,I795658,I795525);
not I_46593 (I795683,I795666);
not I_46594 (I795700,I795658);
nor I_46595 (I795717,I795700,I795601);
DFFARX1 I_46596 (I795717,I3563,I795431,I795417,);
nand I_46597 (I795748,I563205,I563214);
and I_46598 (I795765,I795748,I563220);
DFFARX1 I_46599 (I795765,I3563,I795431,I795791,);
nor I_46600 (I795799,I795791,I795658);
DFFARX1 I_46601 (I795799,I3563,I795431,I795399,);
nand I_46602 (I795830,I795791,I795700);
nand I_46603 (I795408,I795683,I795830);
not I_46604 (I795861,I795791);
nor I_46605 (I795878,I795861,I795601);
DFFARX1 I_46606 (I795878,I3563,I795431,I795420,);
nor I_46607 (I795909,I563217,I563214);
or I_46608 (I795411,I795658,I795909);
nor I_46609 (I795402,I795791,I795909);
or I_46610 (I795405,I795525,I795909);
DFFARX1 I_46611 (I795909,I3563,I795431,I795423,);
not I_46612 (I796009,I3570);
DFFARX1 I_46613 (I567361,I3563,I796009,I796035,);
not I_46614 (I796043,I796035);
nand I_46615 (I796060,I567376,I567361);
and I_46616 (I796077,I796060,I567364);
DFFARX1 I_46617 (I796077,I3563,I796009,I796103,);
not I_46618 (I796111,I567364);
DFFARX1 I_46619 (I567373,I3563,I796009,I796137,);
not I_46620 (I796145,I796137);
nor I_46621 (I796162,I796145,I796043);
and I_46622 (I796179,I796162,I567364);
nor I_46623 (I796196,I796145,I796111);
nor I_46624 (I795992,I796103,I796196);
DFFARX1 I_46625 (I567367,I3563,I796009,I796236,);
nor I_46626 (I796244,I796236,I796103);
not I_46627 (I796261,I796244);
not I_46628 (I796278,I796236);
nor I_46629 (I796295,I796278,I796179);
DFFARX1 I_46630 (I796295,I3563,I796009,I795995,);
nand I_46631 (I796326,I567370,I567379);
and I_46632 (I796343,I796326,I567385);
DFFARX1 I_46633 (I796343,I3563,I796009,I796369,);
nor I_46634 (I796377,I796369,I796236);
DFFARX1 I_46635 (I796377,I3563,I796009,I795977,);
nand I_46636 (I796408,I796369,I796278);
nand I_46637 (I795986,I796261,I796408);
not I_46638 (I796439,I796369);
nor I_46639 (I796456,I796439,I796179);
DFFARX1 I_46640 (I796456,I3563,I796009,I795998,);
nor I_46641 (I796487,I567382,I567379);
or I_46642 (I795989,I796236,I796487);
nor I_46643 (I795980,I796369,I796487);
or I_46644 (I795983,I796103,I796487);
DFFARX1 I_46645 (I796487,I3563,I796009,I796001,);
not I_46646 (I796587,I3570);
DFFARX1 I_46647 (I1174245,I3563,I796587,I796613,);
not I_46648 (I796621,I796613);
nand I_46649 (I796638,I1174227,I1174239);
and I_46650 (I796655,I796638,I1174242);
DFFARX1 I_46651 (I796655,I3563,I796587,I796681,);
not I_46652 (I796689,I1174236);
DFFARX1 I_46653 (I1174233,I3563,I796587,I796715,);
not I_46654 (I796723,I796715);
nor I_46655 (I796740,I796723,I796621);
and I_46656 (I796757,I796740,I1174236);
nor I_46657 (I796774,I796723,I796689);
nor I_46658 (I796570,I796681,I796774);
DFFARX1 I_46659 (I1174251,I3563,I796587,I796814,);
nor I_46660 (I796822,I796814,I796681);
not I_46661 (I796839,I796822);
not I_46662 (I796856,I796814);
nor I_46663 (I796873,I796856,I796757);
DFFARX1 I_46664 (I796873,I3563,I796587,I796573,);
nand I_46665 (I796904,I1174230,I1174230);
and I_46666 (I796921,I796904,I1174227);
DFFARX1 I_46667 (I796921,I3563,I796587,I796947,);
nor I_46668 (I796955,I796947,I796814);
DFFARX1 I_46669 (I796955,I3563,I796587,I796555,);
nand I_46670 (I796986,I796947,I796856);
nand I_46671 (I796564,I796839,I796986);
not I_46672 (I797017,I796947);
nor I_46673 (I797034,I797017,I796757);
DFFARX1 I_46674 (I797034,I3563,I796587,I796576,);
nor I_46675 (I797065,I1174248,I1174230);
or I_46676 (I796567,I796814,I797065);
nor I_46677 (I796558,I796947,I797065);
or I_46678 (I796561,I796681,I797065);
DFFARX1 I_46679 (I797065,I3563,I796587,I796579,);
not I_46680 (I797165,I3570);
DFFARX1 I_46681 (I322279,I3563,I797165,I797191,);
not I_46682 (I797199,I797191);
nand I_46683 (I797216,I322282,I322258);
and I_46684 (I797233,I797216,I322255);
DFFARX1 I_46685 (I797233,I3563,I797165,I797259,);
not I_46686 (I797267,I322261);
DFFARX1 I_46687 (I322255,I3563,I797165,I797293,);
not I_46688 (I797301,I797293);
nor I_46689 (I797318,I797301,I797199);
and I_46690 (I797335,I797318,I322261);
nor I_46691 (I797352,I797301,I797267);
nor I_46692 (I797148,I797259,I797352);
DFFARX1 I_46693 (I322264,I3563,I797165,I797392,);
nor I_46694 (I797400,I797392,I797259);
not I_46695 (I797417,I797400);
not I_46696 (I797434,I797392);
nor I_46697 (I797451,I797434,I797335);
DFFARX1 I_46698 (I797451,I3563,I797165,I797151,);
nand I_46699 (I797482,I322267,I322276);
and I_46700 (I797499,I797482,I322273);
DFFARX1 I_46701 (I797499,I3563,I797165,I797525,);
nor I_46702 (I797533,I797525,I797392);
DFFARX1 I_46703 (I797533,I3563,I797165,I797133,);
nand I_46704 (I797564,I797525,I797434);
nand I_46705 (I797142,I797417,I797564);
not I_46706 (I797595,I797525);
nor I_46707 (I797612,I797595,I797335);
DFFARX1 I_46708 (I797612,I3563,I797165,I797154,);
nor I_46709 (I797643,I322270,I322276);
or I_46710 (I797145,I797392,I797643);
nor I_46711 (I797136,I797525,I797643);
or I_46712 (I797139,I797259,I797643);
DFFARX1 I_46713 (I797643,I3563,I797165,I797157,);
not I_46714 (I797743,I3570);
DFFARX1 I_46715 (I1382725,I3563,I797743,I797769,);
not I_46716 (I797777,I797769);
nand I_46717 (I797794,I1382710,I1382698);
and I_46718 (I797811,I797794,I1382713);
DFFARX1 I_46719 (I797811,I3563,I797743,I797837,);
not I_46720 (I797845,I1382698);
DFFARX1 I_46721 (I1382716,I3563,I797743,I797871,);
not I_46722 (I797879,I797871);
nor I_46723 (I797896,I797879,I797777);
and I_46724 (I797913,I797896,I1382698);
nor I_46725 (I797930,I797879,I797845);
nor I_46726 (I797726,I797837,I797930);
DFFARX1 I_46727 (I1382704,I3563,I797743,I797970,);
nor I_46728 (I797978,I797970,I797837);
not I_46729 (I797995,I797978);
not I_46730 (I798012,I797970);
nor I_46731 (I798029,I798012,I797913);
DFFARX1 I_46732 (I798029,I3563,I797743,I797729,);
nand I_46733 (I798060,I1382701,I1382707);
and I_46734 (I798077,I798060,I1382722);
DFFARX1 I_46735 (I798077,I3563,I797743,I798103,);
nor I_46736 (I798111,I798103,I797970);
DFFARX1 I_46737 (I798111,I3563,I797743,I797711,);
nand I_46738 (I798142,I798103,I798012);
nand I_46739 (I797720,I797995,I798142);
not I_46740 (I798173,I798103);
nor I_46741 (I798190,I798173,I797913);
DFFARX1 I_46742 (I798190,I3563,I797743,I797732,);
nor I_46743 (I798221,I1382719,I1382707);
or I_46744 (I797723,I797970,I798221);
nor I_46745 (I797714,I798103,I798221);
or I_46746 (I797717,I797837,I798221);
DFFARX1 I_46747 (I798221,I3563,I797743,I797735,);
not I_46748 (I798321,I3570);
DFFARX1 I_46749 (I297510,I3563,I798321,I798347,);
not I_46750 (I798355,I798347);
nand I_46751 (I798372,I297513,I297489);
and I_46752 (I798389,I798372,I297486);
DFFARX1 I_46753 (I798389,I3563,I798321,I798415,);
not I_46754 (I798423,I297492);
DFFARX1 I_46755 (I297486,I3563,I798321,I798449,);
not I_46756 (I798457,I798449);
nor I_46757 (I798474,I798457,I798355);
and I_46758 (I798491,I798474,I297492);
nor I_46759 (I798508,I798457,I798423);
nor I_46760 (I798304,I798415,I798508);
DFFARX1 I_46761 (I297495,I3563,I798321,I798548,);
nor I_46762 (I798556,I798548,I798415);
not I_46763 (I798573,I798556);
not I_46764 (I798590,I798548);
nor I_46765 (I798607,I798590,I798491);
DFFARX1 I_46766 (I798607,I3563,I798321,I798307,);
nand I_46767 (I798638,I297498,I297507);
and I_46768 (I798655,I798638,I297504);
DFFARX1 I_46769 (I798655,I3563,I798321,I798681,);
nor I_46770 (I798689,I798681,I798548);
DFFARX1 I_46771 (I798689,I3563,I798321,I798289,);
nand I_46772 (I798720,I798681,I798590);
nand I_46773 (I798298,I798573,I798720);
not I_46774 (I798751,I798681);
nor I_46775 (I798768,I798751,I798491);
DFFARX1 I_46776 (I798768,I3563,I798321,I798310,);
nor I_46777 (I798799,I297501,I297507);
or I_46778 (I798301,I798548,I798799);
nor I_46779 (I798292,I798681,I798799);
or I_46780 (I798295,I798415,I798799);
DFFARX1 I_46781 (I798799,I3563,I798321,I798313,);
not I_46782 (I798899,I3570);
DFFARX1 I_46783 (I861663,I3563,I798899,I798925,);
not I_46784 (I798933,I798925);
nand I_46785 (I798950,I861651,I861669);
and I_46786 (I798967,I798950,I861666);
DFFARX1 I_46787 (I798967,I3563,I798899,I798993,);
not I_46788 (I799001,I861657);
DFFARX1 I_46789 (I861654,I3563,I798899,I799027,);
not I_46790 (I799035,I799027);
nor I_46791 (I799052,I799035,I798933);
and I_46792 (I799069,I799052,I861657);
nor I_46793 (I799086,I799035,I799001);
nor I_46794 (I798882,I798993,I799086);
DFFARX1 I_46795 (I861648,I3563,I798899,I799126,);
nor I_46796 (I799134,I799126,I798993);
not I_46797 (I799151,I799134);
not I_46798 (I799168,I799126);
nor I_46799 (I799185,I799168,I799069);
DFFARX1 I_46800 (I799185,I3563,I798899,I798885,);
nand I_46801 (I799216,I861648,I861651);
and I_46802 (I799233,I799216,I861654);
DFFARX1 I_46803 (I799233,I3563,I798899,I799259,);
nor I_46804 (I799267,I799259,I799126);
DFFARX1 I_46805 (I799267,I3563,I798899,I798867,);
nand I_46806 (I799298,I799259,I799168);
nand I_46807 (I798876,I799151,I799298);
not I_46808 (I799329,I799259);
nor I_46809 (I799346,I799329,I799069);
DFFARX1 I_46810 (I799346,I3563,I798899,I798888,);
nor I_46811 (I799377,I861660,I861651);
or I_46812 (I798879,I799126,I799377);
nor I_46813 (I798870,I799259,I799377);
or I_46814 (I798873,I798993,I799377);
DFFARX1 I_46815 (I799377,I3563,I798899,I798891,);
not I_46816 (I799477,I3570);
DFFARX1 I_46817 (I360223,I3563,I799477,I799503,);
not I_46818 (I799511,I799503);
nand I_46819 (I799528,I360226,I360202);
and I_46820 (I799545,I799528,I360199);
DFFARX1 I_46821 (I799545,I3563,I799477,I799571,);
not I_46822 (I799579,I360205);
DFFARX1 I_46823 (I360199,I3563,I799477,I799605,);
not I_46824 (I799613,I799605);
nor I_46825 (I799630,I799613,I799511);
and I_46826 (I799647,I799630,I360205);
nor I_46827 (I799664,I799613,I799579);
nor I_46828 (I799460,I799571,I799664);
DFFARX1 I_46829 (I360208,I3563,I799477,I799704,);
nor I_46830 (I799712,I799704,I799571);
not I_46831 (I799729,I799712);
not I_46832 (I799746,I799704);
nor I_46833 (I799763,I799746,I799647);
DFFARX1 I_46834 (I799763,I3563,I799477,I799463,);
nand I_46835 (I799794,I360211,I360220);
and I_46836 (I799811,I799794,I360217);
DFFARX1 I_46837 (I799811,I3563,I799477,I799837,);
nor I_46838 (I799845,I799837,I799704);
DFFARX1 I_46839 (I799845,I3563,I799477,I799445,);
nand I_46840 (I799876,I799837,I799746);
nand I_46841 (I799454,I799729,I799876);
not I_46842 (I799907,I799837);
nor I_46843 (I799924,I799907,I799647);
DFFARX1 I_46844 (I799924,I3563,I799477,I799466,);
nor I_46845 (I799955,I360214,I360220);
or I_46846 (I799457,I799704,I799955);
nor I_46847 (I799448,I799837,I799955);
or I_46848 (I799451,I799571,I799955);
DFFARX1 I_46849 (I799955,I3563,I799477,I799469,);
not I_46850 (I800055,I3570);
DFFARX1 I_46851 (I581539,I3563,I800055,I800081,);
not I_46852 (I800089,I800081);
nand I_46853 (I800106,I581548,I581557);
and I_46854 (I800123,I800106,I581563);
DFFARX1 I_46855 (I800123,I3563,I800055,I800149,);
not I_46856 (I800157,I581560);
DFFARX1 I_46857 (I581545,I3563,I800055,I800183,);
not I_46858 (I800191,I800183);
nor I_46859 (I800208,I800191,I800089);
and I_46860 (I800225,I800208,I581560);
nor I_46861 (I800242,I800191,I800157);
nor I_46862 (I800038,I800149,I800242);
DFFARX1 I_46863 (I581554,I3563,I800055,I800282,);
nor I_46864 (I800290,I800282,I800149);
not I_46865 (I800307,I800290);
not I_46866 (I800324,I800282);
nor I_46867 (I800341,I800324,I800225);
DFFARX1 I_46868 (I800341,I3563,I800055,I800041,);
nand I_46869 (I800372,I581551,I581542);
and I_46870 (I800389,I800372,I581539);
DFFARX1 I_46871 (I800389,I3563,I800055,I800415,);
nor I_46872 (I800423,I800415,I800282);
DFFARX1 I_46873 (I800423,I3563,I800055,I800023,);
nand I_46874 (I800454,I800415,I800324);
nand I_46875 (I800032,I800307,I800454);
not I_46876 (I800485,I800415);
nor I_46877 (I800502,I800485,I800225);
DFFARX1 I_46878 (I800502,I3563,I800055,I800044,);
nor I_46879 (I800533,I581542,I581542);
or I_46880 (I800035,I800282,I800533);
nor I_46881 (I800026,I800415,I800533);
or I_46882 (I800029,I800149,I800533);
DFFARX1 I_46883 (I800533,I3563,I800055,I800047,);
not I_46884 (I800633,I3570);
DFFARX1 I_46885 (I923297,I3563,I800633,I800659,);
not I_46886 (I800667,I800659);
nand I_46887 (I800684,I923273,I923288);
and I_46888 (I800701,I800684,I923300);
DFFARX1 I_46889 (I800701,I3563,I800633,I800727,);
not I_46890 (I800735,I923285);
DFFARX1 I_46891 (I923276,I3563,I800633,I800761,);
not I_46892 (I800769,I800761);
nor I_46893 (I800786,I800769,I800667);
and I_46894 (I800803,I800786,I923285);
nor I_46895 (I800820,I800769,I800735);
nor I_46896 (I800616,I800727,I800820);
DFFARX1 I_46897 (I923273,I3563,I800633,I800860,);
nor I_46898 (I800868,I800860,I800727);
not I_46899 (I800885,I800868);
not I_46900 (I800902,I800860);
nor I_46901 (I800919,I800902,I800803);
DFFARX1 I_46902 (I800919,I3563,I800633,I800619,);
nand I_46903 (I800950,I923291,I923282);
and I_46904 (I800967,I800950,I923294);
DFFARX1 I_46905 (I800967,I3563,I800633,I800993,);
nor I_46906 (I801001,I800993,I800860);
DFFARX1 I_46907 (I801001,I3563,I800633,I800601,);
nand I_46908 (I801032,I800993,I800902);
nand I_46909 (I800610,I800885,I801032);
not I_46910 (I801063,I800993);
nor I_46911 (I801080,I801063,I800803);
DFFARX1 I_46912 (I801080,I3563,I800633,I800622,);
nor I_46913 (I801111,I923279,I923282);
or I_46914 (I800613,I800860,I801111);
nor I_46915 (I800604,I800993,I801111);
or I_46916 (I800607,I800727,I801111);
DFFARX1 I_46917 (I801111,I3563,I800633,I800625,);
not I_46918 (I801211,I3570);
DFFARX1 I_46919 (I524139,I3563,I801211,I801237,);
not I_46920 (I801245,I801237);
nand I_46921 (I801262,I524130,I524148);
and I_46922 (I801279,I801262,I524151);
DFFARX1 I_46923 (I801279,I3563,I801211,I801305,);
not I_46924 (I801313,I524145);
DFFARX1 I_46925 (I524133,I3563,I801211,I801339,);
not I_46926 (I801347,I801339);
nor I_46927 (I801364,I801347,I801245);
and I_46928 (I801381,I801364,I524145);
nor I_46929 (I801398,I801347,I801313);
nor I_46930 (I801194,I801305,I801398);
DFFARX1 I_46931 (I524142,I3563,I801211,I801438,);
nor I_46932 (I801446,I801438,I801305);
not I_46933 (I801463,I801446);
not I_46934 (I801480,I801438);
nor I_46935 (I801497,I801480,I801381);
DFFARX1 I_46936 (I801497,I3563,I801211,I801197,);
nand I_46937 (I801528,I524157,I524154);
and I_46938 (I801545,I801528,I524136);
DFFARX1 I_46939 (I801545,I3563,I801211,I801571,);
nor I_46940 (I801579,I801571,I801438);
DFFARX1 I_46941 (I801579,I3563,I801211,I801179,);
nand I_46942 (I801610,I801571,I801480);
nand I_46943 (I801188,I801463,I801610);
not I_46944 (I801641,I801571);
nor I_46945 (I801658,I801641,I801381);
DFFARX1 I_46946 (I801658,I3563,I801211,I801200,);
nor I_46947 (I801689,I524130,I524154);
or I_46948 (I801191,I801438,I801689);
nor I_46949 (I801182,I801571,I801689);
or I_46950 (I801185,I801305,I801689);
DFFARX1 I_46951 (I801689,I3563,I801211,I801203,);
not I_46952 (I801789,I3570);
DFFARX1 I_46953 (I156253,I3563,I801789,I801815,);
not I_46954 (I801823,I801815);
nand I_46955 (I801840,I156262,I156271);
and I_46956 (I801857,I801840,I156250);
DFFARX1 I_46957 (I801857,I3563,I801789,I801883,);
not I_46958 (I801891,I156253);
DFFARX1 I_46959 (I156268,I3563,I801789,I801917,);
not I_46960 (I801925,I801917);
nor I_46961 (I801942,I801925,I801823);
and I_46962 (I801959,I801942,I156253);
nor I_46963 (I801976,I801925,I801891);
nor I_46964 (I801772,I801883,I801976);
DFFARX1 I_46965 (I156259,I3563,I801789,I802016,);
nor I_46966 (I802024,I802016,I801883);
not I_46967 (I802041,I802024);
not I_46968 (I802058,I802016);
nor I_46969 (I802075,I802058,I801959);
DFFARX1 I_46970 (I802075,I3563,I801789,I801775,);
nand I_46971 (I802106,I156274,I156250);
and I_46972 (I802123,I802106,I156256);
DFFARX1 I_46973 (I802123,I3563,I801789,I802149,);
nor I_46974 (I802157,I802149,I802016);
DFFARX1 I_46975 (I802157,I3563,I801789,I801757,);
nand I_46976 (I802188,I802149,I802058);
nand I_46977 (I801766,I802041,I802188);
not I_46978 (I802219,I802149);
nor I_46979 (I802236,I802219,I801959);
DFFARX1 I_46980 (I802236,I3563,I801789,I801778,);
nor I_46981 (I802267,I156265,I156250);
or I_46982 (I801769,I802016,I802267);
nor I_46983 (I801760,I802149,I802267);
or I_46984 (I801763,I801883,I802267);
DFFARX1 I_46985 (I802267,I3563,I801789,I801781,);
not I_46986 (I802367,I3570);
DFFARX1 I_46987 (I236898,I3563,I802367,I802393,);
not I_46988 (I802401,I802393);
nand I_46989 (I802418,I236901,I236922);
and I_46990 (I802435,I802418,I236910);
DFFARX1 I_46991 (I802435,I3563,I802367,I802461,);
not I_46992 (I802469,I236907);
DFFARX1 I_46993 (I236898,I3563,I802367,I802495,);
not I_46994 (I802503,I802495);
nor I_46995 (I802520,I802503,I802401);
and I_46996 (I802537,I802520,I236907);
nor I_46997 (I802554,I802503,I802469);
nor I_46998 (I802350,I802461,I802554);
DFFARX1 I_46999 (I236916,I3563,I802367,I802594,);
nor I_47000 (I802602,I802594,I802461);
not I_47001 (I802619,I802602);
not I_47002 (I802636,I802594);
nor I_47003 (I802653,I802636,I802537);
DFFARX1 I_47004 (I802653,I3563,I802367,I802353,);
nand I_47005 (I802684,I236901,I236904);
and I_47006 (I802701,I802684,I236913);
DFFARX1 I_47007 (I802701,I3563,I802367,I802727,);
nor I_47008 (I802735,I802727,I802594);
DFFARX1 I_47009 (I802735,I3563,I802367,I802335,);
nand I_47010 (I802766,I802727,I802636);
nand I_47011 (I802344,I802619,I802766);
not I_47012 (I802797,I802727);
nor I_47013 (I802814,I802797,I802537);
DFFARX1 I_47014 (I802814,I3563,I802367,I802356,);
nor I_47015 (I802845,I236919,I236904);
or I_47016 (I802347,I802594,I802845);
nor I_47017 (I802338,I802727,I802845);
or I_47018 (I802341,I802461,I802845);
DFFARX1 I_47019 (I802845,I3563,I802367,I802359,);
not I_47020 (I802945,I3570);
DFFARX1 I_47021 (I950429,I3563,I802945,I802971,);
not I_47022 (I802979,I802971);
nand I_47023 (I802996,I950405,I950420);
and I_47024 (I803013,I802996,I950432);
DFFARX1 I_47025 (I803013,I3563,I802945,I803039,);
not I_47026 (I803047,I950417);
DFFARX1 I_47027 (I950408,I3563,I802945,I803073,);
not I_47028 (I803081,I803073);
nor I_47029 (I803098,I803081,I802979);
and I_47030 (I803115,I803098,I950417);
nor I_47031 (I803132,I803081,I803047);
nor I_47032 (I802928,I803039,I803132);
DFFARX1 I_47033 (I950405,I3563,I802945,I803172,);
nor I_47034 (I803180,I803172,I803039);
not I_47035 (I803197,I803180);
not I_47036 (I803214,I803172);
nor I_47037 (I803231,I803214,I803115);
DFFARX1 I_47038 (I803231,I3563,I802945,I802931,);
nand I_47039 (I803262,I950423,I950414);
and I_47040 (I803279,I803262,I950426);
DFFARX1 I_47041 (I803279,I3563,I802945,I803305,);
nor I_47042 (I803313,I803305,I803172);
DFFARX1 I_47043 (I803313,I3563,I802945,I802913,);
nand I_47044 (I803344,I803305,I803214);
nand I_47045 (I802922,I803197,I803344);
not I_47046 (I803375,I803305);
nor I_47047 (I803392,I803375,I803115);
DFFARX1 I_47048 (I803392,I3563,I802945,I802934,);
nor I_47049 (I803423,I950411,I950414);
or I_47050 (I802925,I803172,I803423);
nor I_47051 (I802916,I803305,I803423);
or I_47052 (I802919,I803039,I803423);
DFFARX1 I_47053 (I803423,I3563,I802945,I802937,);
not I_47054 (I803523,I3570);
DFFARX1 I_47055 (I970455,I3563,I803523,I803549,);
not I_47056 (I803557,I803549);
nand I_47057 (I803574,I970431,I970446);
and I_47058 (I803591,I803574,I970458);
DFFARX1 I_47059 (I803591,I3563,I803523,I803617,);
not I_47060 (I803625,I970443);
DFFARX1 I_47061 (I970434,I3563,I803523,I803651,);
not I_47062 (I803659,I803651);
nor I_47063 (I803676,I803659,I803557);
and I_47064 (I803693,I803676,I970443);
nor I_47065 (I803710,I803659,I803625);
nor I_47066 (I803506,I803617,I803710);
DFFARX1 I_47067 (I970431,I3563,I803523,I803750,);
nor I_47068 (I803758,I803750,I803617);
not I_47069 (I803775,I803758);
not I_47070 (I803792,I803750);
nor I_47071 (I803809,I803792,I803693);
DFFARX1 I_47072 (I803809,I3563,I803523,I803509,);
nand I_47073 (I803840,I970449,I970440);
and I_47074 (I803857,I803840,I970452);
DFFARX1 I_47075 (I803857,I3563,I803523,I803883,);
nor I_47076 (I803891,I803883,I803750);
DFFARX1 I_47077 (I803891,I3563,I803523,I803491,);
nand I_47078 (I803922,I803883,I803792);
nand I_47079 (I803500,I803775,I803922);
not I_47080 (I803953,I803883);
nor I_47081 (I803970,I803953,I803693);
DFFARX1 I_47082 (I803970,I3563,I803523,I803512,);
nor I_47083 (I804001,I970437,I970440);
or I_47084 (I803503,I803750,I804001);
nor I_47085 (I803494,I803883,I804001);
or I_47086 (I803497,I803617,I804001);
DFFARX1 I_47087 (I804001,I3563,I803523,I803515,);
not I_47088 (I804101,I3570);
DFFARX1 I_47089 (I588475,I3563,I804101,I804127,);
not I_47090 (I804135,I804127);
nand I_47091 (I804152,I588484,I588493);
and I_47092 (I804169,I804152,I588499);
DFFARX1 I_47093 (I804169,I3563,I804101,I804195,);
not I_47094 (I804203,I588496);
DFFARX1 I_47095 (I588481,I3563,I804101,I804229,);
not I_47096 (I804237,I804229);
nor I_47097 (I804254,I804237,I804135);
and I_47098 (I804271,I804254,I588496);
nor I_47099 (I804288,I804237,I804203);
nor I_47100 (I804084,I804195,I804288);
DFFARX1 I_47101 (I588490,I3563,I804101,I804328,);
nor I_47102 (I804336,I804328,I804195);
not I_47103 (I804353,I804336);
not I_47104 (I804370,I804328);
nor I_47105 (I804387,I804370,I804271);
DFFARX1 I_47106 (I804387,I3563,I804101,I804087,);
nand I_47107 (I804418,I588487,I588478);
and I_47108 (I804435,I804418,I588475);
DFFARX1 I_47109 (I804435,I3563,I804101,I804461,);
nor I_47110 (I804469,I804461,I804328);
DFFARX1 I_47111 (I804469,I3563,I804101,I804069,);
nand I_47112 (I804500,I804461,I804370);
nand I_47113 (I804078,I804353,I804500);
not I_47114 (I804531,I804461);
nor I_47115 (I804548,I804531,I804271);
DFFARX1 I_47116 (I804548,I3563,I804101,I804090,);
nor I_47117 (I804579,I588478,I588478);
or I_47118 (I804081,I804328,I804579);
nor I_47119 (I804072,I804461,I804579);
or I_47120 (I804075,I804195,I804579);
DFFARX1 I_47121 (I804579,I3563,I804101,I804093,);
not I_47122 (I804679,I3570);
DFFARX1 I_47123 (I416612,I3563,I804679,I804705,);
not I_47124 (I804713,I804705);
nand I_47125 (I804730,I416615,I416591);
and I_47126 (I804747,I804730,I416588);
DFFARX1 I_47127 (I804747,I3563,I804679,I804773,);
not I_47128 (I804781,I416594);
DFFARX1 I_47129 (I416588,I3563,I804679,I804807,);
not I_47130 (I804815,I804807);
nor I_47131 (I804832,I804815,I804713);
and I_47132 (I804849,I804832,I416594);
nor I_47133 (I804866,I804815,I804781);
nor I_47134 (I804662,I804773,I804866);
DFFARX1 I_47135 (I416597,I3563,I804679,I804906,);
nor I_47136 (I804914,I804906,I804773);
not I_47137 (I804931,I804914);
not I_47138 (I804948,I804906);
nor I_47139 (I804965,I804948,I804849);
DFFARX1 I_47140 (I804965,I3563,I804679,I804665,);
nand I_47141 (I804996,I416600,I416609);
and I_47142 (I805013,I804996,I416606);
DFFARX1 I_47143 (I805013,I3563,I804679,I805039,);
nor I_47144 (I805047,I805039,I804906);
DFFARX1 I_47145 (I805047,I3563,I804679,I804647,);
nand I_47146 (I805078,I805039,I804948);
nand I_47147 (I804656,I804931,I805078);
not I_47148 (I805109,I805039);
nor I_47149 (I805126,I805109,I804849);
DFFARX1 I_47150 (I805126,I3563,I804679,I804668,);
nor I_47151 (I805157,I416603,I416609);
or I_47152 (I804659,I804906,I805157);
nor I_47153 (I804650,I805039,I805157);
or I_47154 (I804653,I804773,I805157);
DFFARX1 I_47155 (I805157,I3563,I804679,I804671,);
not I_47156 (I805257,I3570);
DFFARX1 I_47157 (I345467,I3563,I805257,I805283,);
not I_47158 (I805291,I805283);
nand I_47159 (I805308,I345470,I345446);
and I_47160 (I805325,I805308,I345443);
DFFARX1 I_47161 (I805325,I3563,I805257,I805351,);
not I_47162 (I805359,I345449);
DFFARX1 I_47163 (I345443,I3563,I805257,I805385,);
not I_47164 (I805393,I805385);
nor I_47165 (I805410,I805393,I805291);
and I_47166 (I805427,I805410,I345449);
nor I_47167 (I805444,I805393,I805359);
nor I_47168 (I805240,I805351,I805444);
DFFARX1 I_47169 (I345452,I3563,I805257,I805484,);
nor I_47170 (I805492,I805484,I805351);
not I_47171 (I805509,I805492);
not I_47172 (I805526,I805484);
nor I_47173 (I805543,I805526,I805427);
DFFARX1 I_47174 (I805543,I3563,I805257,I805243,);
nand I_47175 (I805574,I345455,I345464);
and I_47176 (I805591,I805574,I345461);
DFFARX1 I_47177 (I805591,I3563,I805257,I805617,);
nor I_47178 (I805625,I805617,I805484);
DFFARX1 I_47179 (I805625,I3563,I805257,I805225,);
nand I_47180 (I805656,I805617,I805526);
nand I_47181 (I805234,I805509,I805656);
not I_47182 (I805687,I805617);
nor I_47183 (I805704,I805687,I805427);
DFFARX1 I_47184 (I805704,I3563,I805257,I805246,);
nor I_47185 (I805735,I345458,I345464);
or I_47186 (I805237,I805484,I805735);
nor I_47187 (I805228,I805617,I805735);
or I_47188 (I805231,I805351,I805735);
DFFARX1 I_47189 (I805735,I3563,I805257,I805249,);
not I_47190 (I805835,I3570);
DFFARX1 I_47191 (I993711,I3563,I805835,I805861,);
not I_47192 (I805869,I805861);
nand I_47193 (I805886,I993687,I993702);
and I_47194 (I805903,I805886,I993714);
DFFARX1 I_47195 (I805903,I3563,I805835,I805929,);
not I_47196 (I805937,I993699);
DFFARX1 I_47197 (I993690,I3563,I805835,I805963,);
not I_47198 (I805971,I805963);
nor I_47199 (I805988,I805971,I805869);
and I_47200 (I806005,I805988,I993699);
nor I_47201 (I806022,I805971,I805937);
nor I_47202 (I805818,I805929,I806022);
DFFARX1 I_47203 (I993687,I3563,I805835,I806062,);
nor I_47204 (I806070,I806062,I805929);
not I_47205 (I806087,I806070);
not I_47206 (I806104,I806062);
nor I_47207 (I806121,I806104,I806005);
DFFARX1 I_47208 (I806121,I3563,I805835,I805821,);
nand I_47209 (I806152,I993705,I993696);
and I_47210 (I806169,I806152,I993708);
DFFARX1 I_47211 (I806169,I3563,I805835,I806195,);
nor I_47212 (I806203,I806195,I806062);
DFFARX1 I_47213 (I806203,I3563,I805835,I805803,);
nand I_47214 (I806234,I806195,I806104);
nand I_47215 (I805812,I806087,I806234);
not I_47216 (I806265,I806195);
nor I_47217 (I806282,I806265,I806005);
DFFARX1 I_47218 (I806282,I3563,I805835,I805824,);
nor I_47219 (I806313,I993693,I993696);
or I_47220 (I805815,I806062,I806313);
nor I_47221 (I805806,I806195,I806313);
or I_47222 (I805809,I805929,I806313);
DFFARX1 I_47223 (I806313,I3563,I805835,I805827,);
not I_47224 (I806413,I3570);
DFFARX1 I_47225 (I935571,I3563,I806413,I806439,);
not I_47226 (I806447,I806439);
nand I_47227 (I806464,I935547,I935562);
and I_47228 (I806481,I806464,I935574);
DFFARX1 I_47229 (I806481,I3563,I806413,I806507,);
not I_47230 (I806515,I935559);
DFFARX1 I_47231 (I935550,I3563,I806413,I806541,);
not I_47232 (I806549,I806541);
nor I_47233 (I806566,I806549,I806447);
and I_47234 (I806583,I806566,I935559);
nor I_47235 (I806600,I806549,I806515);
nor I_47236 (I806396,I806507,I806600);
DFFARX1 I_47237 (I935547,I3563,I806413,I806640,);
nor I_47238 (I806648,I806640,I806507);
not I_47239 (I806665,I806648);
not I_47240 (I806682,I806640);
nor I_47241 (I806699,I806682,I806583);
DFFARX1 I_47242 (I806699,I3563,I806413,I806399,);
nand I_47243 (I806730,I935565,I935556);
and I_47244 (I806747,I806730,I935568);
DFFARX1 I_47245 (I806747,I3563,I806413,I806773,);
nor I_47246 (I806781,I806773,I806640);
DFFARX1 I_47247 (I806781,I3563,I806413,I806381,);
nand I_47248 (I806812,I806773,I806682);
nand I_47249 (I806390,I806665,I806812);
not I_47250 (I806843,I806773);
nor I_47251 (I806860,I806843,I806583);
DFFARX1 I_47252 (I806860,I3563,I806413,I806402,);
nor I_47253 (I806891,I935553,I935556);
or I_47254 (I806393,I806640,I806891);
nor I_47255 (I806384,I806773,I806891);
or I_47256 (I806387,I806507,I806891);
DFFARX1 I_47257 (I806891,I3563,I806413,I806405,);
not I_47258 (I806991,I3570);
DFFARX1 I_47259 (I406072,I3563,I806991,I807017,);
not I_47260 (I807025,I807017);
nand I_47261 (I807042,I406075,I406051);
and I_47262 (I807059,I807042,I406048);
DFFARX1 I_47263 (I807059,I3563,I806991,I807085,);
not I_47264 (I807093,I406054);
DFFARX1 I_47265 (I406048,I3563,I806991,I807119,);
not I_47266 (I807127,I807119);
nor I_47267 (I807144,I807127,I807025);
and I_47268 (I807161,I807144,I406054);
nor I_47269 (I807178,I807127,I807093);
nor I_47270 (I806974,I807085,I807178);
DFFARX1 I_47271 (I406057,I3563,I806991,I807218,);
nor I_47272 (I807226,I807218,I807085);
not I_47273 (I807243,I807226);
not I_47274 (I807260,I807218);
nor I_47275 (I807277,I807260,I807161);
DFFARX1 I_47276 (I807277,I3563,I806991,I806977,);
nand I_47277 (I807308,I406060,I406069);
and I_47278 (I807325,I807308,I406066);
DFFARX1 I_47279 (I807325,I3563,I806991,I807351,);
nor I_47280 (I807359,I807351,I807218);
DFFARX1 I_47281 (I807359,I3563,I806991,I806959,);
nand I_47282 (I807390,I807351,I807260);
nand I_47283 (I806968,I807243,I807390);
not I_47284 (I807421,I807351);
nor I_47285 (I807438,I807421,I807161);
DFFARX1 I_47286 (I807438,I3563,I806991,I806980,);
nor I_47287 (I807469,I406063,I406069);
or I_47288 (I806971,I807218,I807469);
nor I_47289 (I806962,I807351,I807469);
or I_47290 (I806965,I807085,I807469);
DFFARX1 I_47291 (I807469,I3563,I806991,I806983,);
not I_47292 (I807569,I3570);
DFFARX1 I_47293 (I162535,I3563,I807569,I807595,);
not I_47294 (I807603,I807595);
nand I_47295 (I807620,I162550,I162523);
and I_47296 (I807637,I807620,I162538);
DFFARX1 I_47297 (I807637,I3563,I807569,I807663,);
not I_47298 (I807671,I162541);
DFFARX1 I_47299 (I162526,I3563,I807569,I807697,);
not I_47300 (I807705,I807697);
nor I_47301 (I807722,I807705,I807603);
and I_47302 (I807739,I807722,I162541);
nor I_47303 (I807756,I807705,I807671);
nor I_47304 (I807552,I807663,I807756);
DFFARX1 I_47305 (I162532,I3563,I807569,I807796,);
nor I_47306 (I807804,I807796,I807663);
not I_47307 (I807821,I807804);
not I_47308 (I807838,I807796);
nor I_47309 (I807855,I807838,I807739);
DFFARX1 I_47310 (I807855,I3563,I807569,I807555,);
nand I_47311 (I807886,I162547,I162529);
and I_47312 (I807903,I807886,I162544);
DFFARX1 I_47313 (I807903,I3563,I807569,I807929,);
nor I_47314 (I807937,I807929,I807796);
DFFARX1 I_47315 (I807937,I3563,I807569,I807537,);
nand I_47316 (I807968,I807929,I807838);
nand I_47317 (I807546,I807821,I807968);
not I_47318 (I807999,I807929);
nor I_47319 (I808016,I807999,I807739);
DFFARX1 I_47320 (I808016,I3563,I807569,I807558,);
nor I_47321 (I808047,I162523,I162529);
or I_47322 (I807549,I807796,I808047);
nor I_47323 (I807540,I807929,I808047);
or I_47324 (I807543,I807663,I808047);
DFFARX1 I_47325 (I808047,I3563,I807569,I807561,);
not I_47326 (I808147,I3570);
DFFARX1 I_47327 (I26620,I3563,I808147,I808173,);
not I_47328 (I808181,I808173);
nand I_47329 (I808198,I26617,I26608);
and I_47330 (I808215,I808198,I26608);
DFFARX1 I_47331 (I808215,I3563,I808147,I808241,);
not I_47332 (I808249,I26611);
DFFARX1 I_47333 (I26626,I3563,I808147,I808275,);
not I_47334 (I808283,I808275);
nor I_47335 (I808300,I808283,I808181);
and I_47336 (I808317,I808300,I26611);
nor I_47337 (I808334,I808283,I808249);
nor I_47338 (I808130,I808241,I808334);
DFFARX1 I_47339 (I26611,I3563,I808147,I808374,);
nor I_47340 (I808382,I808374,I808241);
not I_47341 (I808399,I808382);
not I_47342 (I808416,I808374);
nor I_47343 (I808433,I808416,I808317);
DFFARX1 I_47344 (I808433,I3563,I808147,I808133,);
nand I_47345 (I808464,I26629,I26614);
and I_47346 (I808481,I808464,I26632);
DFFARX1 I_47347 (I808481,I3563,I808147,I808507,);
nor I_47348 (I808515,I808507,I808374);
DFFARX1 I_47349 (I808515,I3563,I808147,I808115,);
nand I_47350 (I808546,I808507,I808416);
nand I_47351 (I808124,I808399,I808546);
not I_47352 (I808577,I808507);
nor I_47353 (I808594,I808577,I808317);
DFFARX1 I_47354 (I808594,I3563,I808147,I808136,);
nor I_47355 (I808625,I26623,I26614);
or I_47356 (I808127,I808374,I808625);
nor I_47357 (I808118,I808507,I808625);
or I_47358 (I808121,I808241,I808625);
DFFARX1 I_47359 (I808625,I3563,I808147,I808139,);
not I_47360 (I808725,I3570);
DFFARX1 I_47361 (I1401765,I3563,I808725,I808751,);
not I_47362 (I808759,I808751);
nand I_47363 (I808776,I1401750,I1401738);
and I_47364 (I808793,I808776,I1401753);
DFFARX1 I_47365 (I808793,I3563,I808725,I808819,);
not I_47366 (I808827,I1401738);
DFFARX1 I_47367 (I1401756,I3563,I808725,I808853,);
not I_47368 (I808861,I808853);
nor I_47369 (I808878,I808861,I808759);
and I_47370 (I808895,I808878,I1401738);
nor I_47371 (I808912,I808861,I808827);
nor I_47372 (I808708,I808819,I808912);
DFFARX1 I_47373 (I1401744,I3563,I808725,I808952,);
nor I_47374 (I808960,I808952,I808819);
not I_47375 (I808977,I808960);
not I_47376 (I808994,I808952);
nor I_47377 (I809011,I808994,I808895);
DFFARX1 I_47378 (I809011,I3563,I808725,I808711,);
nand I_47379 (I809042,I1401741,I1401747);
and I_47380 (I809059,I809042,I1401762);
DFFARX1 I_47381 (I809059,I3563,I808725,I809085,);
nor I_47382 (I809093,I809085,I808952);
DFFARX1 I_47383 (I809093,I3563,I808725,I808693,);
nand I_47384 (I809124,I809085,I808994);
nand I_47385 (I808702,I808977,I809124);
not I_47386 (I809155,I809085);
nor I_47387 (I809172,I809155,I808895);
DFFARX1 I_47388 (I809172,I3563,I808725,I808714,);
nor I_47389 (I809203,I1401759,I1401747);
or I_47390 (I808705,I808952,I809203);
nor I_47391 (I808696,I809085,I809203);
or I_47392 (I808699,I808819,I809203);
DFFARX1 I_47393 (I809203,I3563,I808725,I808717,);
not I_47394 (I809303,I3570);
DFFARX1 I_47395 (I1287753,I3563,I809303,I809329,);
not I_47396 (I809337,I809329);
nand I_47397 (I809354,I1287777,I1287759);
and I_47398 (I809371,I809354,I1287765);
DFFARX1 I_47399 (I809371,I3563,I809303,I809397,);
not I_47400 (I809405,I1287771);
DFFARX1 I_47401 (I1287756,I3563,I809303,I809431,);
not I_47402 (I809439,I809431);
nor I_47403 (I809456,I809439,I809337);
and I_47404 (I809473,I809456,I1287771);
nor I_47405 (I809490,I809439,I809405);
nor I_47406 (I809286,I809397,I809490);
DFFARX1 I_47407 (I1287768,I3563,I809303,I809530,);
nor I_47408 (I809538,I809530,I809397);
not I_47409 (I809555,I809538);
not I_47410 (I809572,I809530);
nor I_47411 (I809589,I809572,I809473);
DFFARX1 I_47412 (I809589,I3563,I809303,I809289,);
nand I_47413 (I809620,I1287774,I1287762);
and I_47414 (I809637,I809620,I1287756);
DFFARX1 I_47415 (I809637,I3563,I809303,I809663,);
nor I_47416 (I809671,I809663,I809530);
DFFARX1 I_47417 (I809671,I3563,I809303,I809271,);
nand I_47418 (I809702,I809663,I809572);
nand I_47419 (I809280,I809555,I809702);
not I_47420 (I809733,I809663);
nor I_47421 (I809750,I809733,I809473);
DFFARX1 I_47422 (I809750,I3563,I809303,I809292,);
nor I_47423 (I809781,I1287753,I1287762);
or I_47424 (I809283,I809530,I809781);
nor I_47425 (I809274,I809663,I809781);
or I_47426 (I809277,I809397,I809781);
DFFARX1 I_47427 (I809781,I3563,I809303,I809295,);
not I_47428 (I809881,I3570);
DFFARX1 I_47429 (I949137,I3563,I809881,I809907,);
not I_47430 (I809915,I809907);
nand I_47431 (I809932,I949113,I949128);
and I_47432 (I809949,I809932,I949140);
DFFARX1 I_47433 (I809949,I3563,I809881,I809975,);
not I_47434 (I809983,I949125);
DFFARX1 I_47435 (I949116,I3563,I809881,I810009,);
not I_47436 (I810017,I810009);
nor I_47437 (I810034,I810017,I809915);
and I_47438 (I810051,I810034,I949125);
nor I_47439 (I810068,I810017,I809983);
nor I_47440 (I809864,I809975,I810068);
DFFARX1 I_47441 (I949113,I3563,I809881,I810108,);
nor I_47442 (I810116,I810108,I809975);
not I_47443 (I810133,I810116);
not I_47444 (I810150,I810108);
nor I_47445 (I810167,I810150,I810051);
DFFARX1 I_47446 (I810167,I3563,I809881,I809867,);
nand I_47447 (I810198,I949131,I949122);
and I_47448 (I810215,I810198,I949134);
DFFARX1 I_47449 (I810215,I3563,I809881,I810241,);
nor I_47450 (I810249,I810241,I810108);
DFFARX1 I_47451 (I810249,I3563,I809881,I809849,);
nand I_47452 (I810280,I810241,I810150);
nand I_47453 (I809858,I810133,I810280);
not I_47454 (I810311,I810241);
nor I_47455 (I810328,I810311,I810051);
DFFARX1 I_47456 (I810328,I3563,I809881,I809870,);
nor I_47457 (I810359,I949119,I949122);
or I_47458 (I809861,I810108,I810359);
nor I_47459 (I809852,I810241,I810359);
or I_47460 (I809855,I809975,I810359);
DFFARX1 I_47461 (I810359,I3563,I809881,I809873,);
not I_47462 (I810459,I3570);
DFFARX1 I_47463 (I902242,I3563,I810459,I810485,);
not I_47464 (I810493,I810485);
nand I_47465 (I810510,I902230,I902248);
and I_47466 (I810527,I810510,I902245);
DFFARX1 I_47467 (I810527,I3563,I810459,I810553,);
not I_47468 (I810561,I902236);
DFFARX1 I_47469 (I902233,I3563,I810459,I810587,);
not I_47470 (I810595,I810587);
nor I_47471 (I810612,I810595,I810493);
and I_47472 (I810629,I810612,I902236);
nor I_47473 (I810646,I810595,I810561);
nor I_47474 (I810442,I810553,I810646);
DFFARX1 I_47475 (I902227,I3563,I810459,I810686,);
nor I_47476 (I810694,I810686,I810553);
not I_47477 (I810711,I810694);
not I_47478 (I810728,I810686);
nor I_47479 (I810745,I810728,I810629);
DFFARX1 I_47480 (I810745,I3563,I810459,I810445,);
nand I_47481 (I810776,I902227,I902230);
and I_47482 (I810793,I810776,I902233);
DFFARX1 I_47483 (I810793,I3563,I810459,I810819,);
nor I_47484 (I810827,I810819,I810686);
DFFARX1 I_47485 (I810827,I3563,I810459,I810427,);
nand I_47486 (I810858,I810819,I810728);
nand I_47487 (I810436,I810711,I810858);
not I_47488 (I810889,I810819);
nor I_47489 (I810906,I810889,I810629);
DFFARX1 I_47490 (I810906,I3563,I810459,I810448,);
nor I_47491 (I810937,I902239,I902230);
or I_47492 (I810439,I810686,I810937);
nor I_47493 (I810430,I810819,I810937);
or I_47494 (I810433,I810553,I810937);
DFFARX1 I_47495 (I810937,I3563,I810459,I810451,);
not I_47496 (I811037,I3570);
DFFARX1 I_47497 (I421355,I3563,I811037,I811063,);
not I_47498 (I811071,I811063);
nand I_47499 (I811088,I421358,I421334);
and I_47500 (I811105,I811088,I421331);
DFFARX1 I_47501 (I811105,I3563,I811037,I811131,);
not I_47502 (I811139,I421337);
DFFARX1 I_47503 (I421331,I3563,I811037,I811165,);
not I_47504 (I811173,I811165);
nor I_47505 (I811190,I811173,I811071);
and I_47506 (I811207,I811190,I421337);
nor I_47507 (I811224,I811173,I811139);
nor I_47508 (I811020,I811131,I811224);
DFFARX1 I_47509 (I421340,I3563,I811037,I811264,);
nor I_47510 (I811272,I811264,I811131);
not I_47511 (I811289,I811272);
not I_47512 (I811306,I811264);
nor I_47513 (I811323,I811306,I811207);
DFFARX1 I_47514 (I811323,I3563,I811037,I811023,);
nand I_47515 (I811354,I421343,I421352);
and I_47516 (I811371,I811354,I421349);
DFFARX1 I_47517 (I811371,I3563,I811037,I811397,);
nor I_47518 (I811405,I811397,I811264);
DFFARX1 I_47519 (I811405,I3563,I811037,I811005,);
nand I_47520 (I811436,I811397,I811306);
nand I_47521 (I811014,I811289,I811436);
not I_47522 (I811467,I811397);
nor I_47523 (I811484,I811467,I811207);
DFFARX1 I_47524 (I811484,I3563,I811037,I811026,);
nor I_47525 (I811515,I421346,I421352);
or I_47526 (I811017,I811264,I811515);
nor I_47527 (I811008,I811397,I811515);
or I_47528 (I811011,I811131,I811515);
DFFARX1 I_47529 (I811515,I3563,I811037,I811029,);
not I_47530 (I811612,I3570);
DFFARX1 I_47531 (I392355,I3563,I811612,I811638,);
not I_47532 (I811646,I811638);
nand I_47533 (I811663,I392346,I392346);
and I_47534 (I811680,I811663,I392364);
DFFARX1 I_47535 (I811680,I3563,I811612,I811706,);
DFFARX1 I_47536 (I811706,I3563,I811612,I811601,);
DFFARX1 I_47537 (I392367,I3563,I811612,I811737,);
nand I_47538 (I811745,I811737,I392349);
not I_47539 (I811762,I811745);
DFFARX1 I_47540 (I811762,I3563,I811612,I811788,);
not I_47541 (I811796,I811788);
nor I_47542 (I811604,I811646,I811796);
DFFARX1 I_47543 (I392361,I3563,I811612,I811836,);
nor I_47544 (I811595,I811836,I811706);
nor I_47545 (I811586,I811836,I811762);
nand I_47546 (I811872,I392373,I392352);
and I_47547 (I811889,I811872,I392358);
DFFARX1 I_47548 (I811889,I3563,I811612,I811915,);
not I_47549 (I811923,I811915);
nand I_47550 (I811940,I811923,I811836);
nand I_47551 (I811589,I811923,I811745);
nor I_47552 (I811971,I392370,I392352);
and I_47553 (I811988,I811836,I811971);
nor I_47554 (I812005,I811923,I811988);
DFFARX1 I_47555 (I812005,I3563,I811612,I811598,);
nor I_47556 (I812036,I811638,I811971);
DFFARX1 I_47557 (I812036,I3563,I811612,I811583,);
nor I_47558 (I812067,I811915,I811971);
not I_47559 (I812084,I812067);
nand I_47560 (I811592,I812084,I811940);
not I_47561 (I812139,I3570);
DFFARX1 I_47562 (I73535,I3563,I812139,I812165,);
not I_47563 (I812173,I812165);
nand I_47564 (I812190,I73511,I73520);
and I_47565 (I812207,I812190,I73514);
DFFARX1 I_47566 (I812207,I3563,I812139,I812233,);
DFFARX1 I_47567 (I812233,I3563,I812139,I812128,);
DFFARX1 I_47568 (I73532,I3563,I812139,I812264,);
nand I_47569 (I812272,I812264,I73523);
not I_47570 (I812289,I812272);
DFFARX1 I_47571 (I812289,I3563,I812139,I812315,);
not I_47572 (I812323,I812315);
nor I_47573 (I812131,I812173,I812323);
DFFARX1 I_47574 (I73517,I3563,I812139,I812363,);
nor I_47575 (I812122,I812363,I812233);
nor I_47576 (I812113,I812363,I812289);
nand I_47577 (I812399,I73529,I73526);
and I_47578 (I812416,I812399,I73514);
DFFARX1 I_47579 (I812416,I3563,I812139,I812442,);
not I_47580 (I812450,I812442);
nand I_47581 (I812467,I812450,I812363);
nand I_47582 (I812116,I812450,I812272);
nor I_47583 (I812498,I73511,I73526);
and I_47584 (I812515,I812363,I812498);
nor I_47585 (I812532,I812450,I812515);
DFFARX1 I_47586 (I812532,I3563,I812139,I812125,);
nor I_47587 (I812563,I812165,I812498);
DFFARX1 I_47588 (I812563,I3563,I812139,I812110,);
nor I_47589 (I812594,I812442,I812498);
not I_47590 (I812611,I812594);
nand I_47591 (I812119,I812611,I812467);
not I_47592 (I812666,I3570);
DFFARX1 I_47593 (I1083133,I3563,I812666,I812692,);
not I_47594 (I812700,I812692);
nand I_47595 (I812717,I1083142,I1083130);
and I_47596 (I812734,I812717,I1083127);
DFFARX1 I_47597 (I812734,I3563,I812666,I812760,);
DFFARX1 I_47598 (I812760,I3563,I812666,I812655,);
DFFARX1 I_47599 (I1083127,I3563,I812666,I812791,);
nand I_47600 (I812799,I812791,I1083124);
not I_47601 (I812816,I812799);
DFFARX1 I_47602 (I812816,I3563,I812666,I812842,);
not I_47603 (I812850,I812842);
nor I_47604 (I812658,I812700,I812850);
DFFARX1 I_47605 (I1083130,I3563,I812666,I812890,);
nor I_47606 (I812649,I812890,I812760);
nor I_47607 (I812640,I812890,I812816);
nand I_47608 (I812926,I1083145,I1083136);
and I_47609 (I812943,I812926,I1083139);
DFFARX1 I_47610 (I812943,I3563,I812666,I812969,);
not I_47611 (I812977,I812969);
nand I_47612 (I812994,I812977,I812890);
nand I_47613 (I812643,I812977,I812799);
nor I_47614 (I813025,I1083124,I1083136);
and I_47615 (I813042,I812890,I813025);
nor I_47616 (I813059,I812977,I813042);
DFFARX1 I_47617 (I813059,I3563,I812666,I812652,);
nor I_47618 (I813090,I812692,I813025);
DFFARX1 I_47619 (I813090,I3563,I812666,I812637,);
nor I_47620 (I813121,I812969,I813025);
not I_47621 (I813138,I813121);
nand I_47622 (I812646,I813138,I812994);
not I_47623 (I813193,I3570);
DFFARX1 I_47624 (I213699,I3563,I813193,I813219,);
not I_47625 (I813227,I813219);
nand I_47626 (I813244,I213696,I213714);
and I_47627 (I813261,I813244,I213705);
DFFARX1 I_47628 (I813261,I3563,I813193,I813287,);
DFFARX1 I_47629 (I813287,I3563,I813193,I813182,);
DFFARX1 I_47630 (I213711,I3563,I813193,I813318,);
nand I_47631 (I813326,I813318,I213708);
not I_47632 (I813343,I813326);
DFFARX1 I_47633 (I813343,I3563,I813193,I813369,);
not I_47634 (I813377,I813369);
nor I_47635 (I813185,I813227,I813377);
DFFARX1 I_47636 (I213702,I3563,I813193,I813417,);
nor I_47637 (I813176,I813417,I813287);
nor I_47638 (I813167,I813417,I813343);
nand I_47639 (I813453,I213693,I213717);
and I_47640 (I813470,I813453,I213696);
DFFARX1 I_47641 (I813470,I3563,I813193,I813496,);
not I_47642 (I813504,I813496);
nand I_47643 (I813521,I813504,I813417);
nand I_47644 (I813170,I813504,I813326);
nor I_47645 (I813552,I213693,I213717);
and I_47646 (I813569,I813417,I813552);
nor I_47647 (I813586,I813504,I813569);
DFFARX1 I_47648 (I813586,I3563,I813193,I813179,);
nor I_47649 (I813617,I813219,I813552);
DFFARX1 I_47650 (I813617,I3563,I813193,I813164,);
nor I_47651 (I813648,I813496,I813552);
not I_47652 (I813665,I813648);
nand I_47653 (I813173,I813665,I813521);
not I_47654 (I813720,I3570);
DFFARX1 I_47655 (I1134363,I3563,I813720,I813746,);
not I_47656 (I813754,I813746);
nand I_47657 (I813771,I1134345,I1134345);
and I_47658 (I813788,I813771,I1134351);
DFFARX1 I_47659 (I813788,I3563,I813720,I813814,);
DFFARX1 I_47660 (I813814,I3563,I813720,I813709,);
DFFARX1 I_47661 (I1134348,I3563,I813720,I813845,);
nand I_47662 (I813853,I813845,I1134357);
not I_47663 (I813870,I813853);
DFFARX1 I_47664 (I813870,I3563,I813720,I813896,);
not I_47665 (I813904,I813896);
nor I_47666 (I813712,I813754,I813904);
DFFARX1 I_47667 (I1134369,I3563,I813720,I813944,);
nor I_47668 (I813703,I813944,I813814);
nor I_47669 (I813694,I813944,I813870);
nand I_47670 (I813980,I1134360,I1134354);
and I_47671 (I813997,I813980,I1134348);
DFFARX1 I_47672 (I813997,I3563,I813720,I814023,);
not I_47673 (I814031,I814023);
nand I_47674 (I814048,I814031,I813944);
nand I_47675 (I813697,I814031,I813853);
nor I_47676 (I814079,I1134366,I1134354);
and I_47677 (I814096,I813944,I814079);
nor I_47678 (I814113,I814031,I814096);
DFFARX1 I_47679 (I814113,I3563,I813720,I813706,);
nor I_47680 (I814144,I813746,I814079);
DFFARX1 I_47681 (I814144,I3563,I813720,I813691,);
nor I_47682 (I814175,I814023,I814079);
not I_47683 (I814192,I814175);
nand I_47684 (I813700,I814192,I814048);
not I_47685 (I814247,I3570);
DFFARX1 I_47686 (I721993,I3563,I814247,I814273,);
not I_47687 (I814281,I814273);
nand I_47688 (I814298,I721996,I721993);
and I_47689 (I814315,I814298,I722005);
DFFARX1 I_47690 (I814315,I3563,I814247,I814341,);
DFFARX1 I_47691 (I814341,I3563,I814247,I814236,);
DFFARX1 I_47692 (I722002,I3563,I814247,I814372,);
nand I_47693 (I814380,I814372,I722008);
not I_47694 (I814397,I814380);
DFFARX1 I_47695 (I814397,I3563,I814247,I814423,);
not I_47696 (I814431,I814423);
nor I_47697 (I814239,I814281,I814431);
DFFARX1 I_47698 (I722017,I3563,I814247,I814471,);
nor I_47699 (I814230,I814471,I814341);
nor I_47700 (I814221,I814471,I814397);
nand I_47701 (I814507,I722011,I721999);
and I_47702 (I814524,I814507,I721996);
DFFARX1 I_47703 (I814524,I3563,I814247,I814550,);
not I_47704 (I814558,I814550);
nand I_47705 (I814575,I814558,I814471);
nand I_47706 (I814224,I814558,I814380);
nor I_47707 (I814606,I722014,I721999);
and I_47708 (I814623,I814471,I814606);
nor I_47709 (I814640,I814558,I814623);
DFFARX1 I_47710 (I814640,I3563,I814247,I814233,);
nor I_47711 (I814671,I814273,I814606);
DFFARX1 I_47712 (I814671,I3563,I814247,I814218,);
nor I_47713 (I814702,I814550,I814606);
not I_47714 (I814719,I814702);
nand I_47715 (I814227,I814719,I814575);
not I_47716 (I814774,I3570);
DFFARX1 I_47717 (I723727,I3563,I814774,I814800,);
not I_47718 (I814808,I814800);
nand I_47719 (I814825,I723730,I723727);
and I_47720 (I814842,I814825,I723739);
DFFARX1 I_47721 (I814842,I3563,I814774,I814868,);
DFFARX1 I_47722 (I814868,I3563,I814774,I814763,);
DFFARX1 I_47723 (I723736,I3563,I814774,I814899,);
nand I_47724 (I814907,I814899,I723742);
not I_47725 (I814924,I814907);
DFFARX1 I_47726 (I814924,I3563,I814774,I814950,);
not I_47727 (I814958,I814950);
nor I_47728 (I814766,I814808,I814958);
DFFARX1 I_47729 (I723751,I3563,I814774,I814998,);
nor I_47730 (I814757,I814998,I814868);
nor I_47731 (I814748,I814998,I814924);
nand I_47732 (I815034,I723745,I723733);
and I_47733 (I815051,I815034,I723730);
DFFARX1 I_47734 (I815051,I3563,I814774,I815077,);
not I_47735 (I815085,I815077);
nand I_47736 (I815102,I815085,I814998);
nand I_47737 (I814751,I815085,I814907);
nor I_47738 (I815133,I723748,I723733);
and I_47739 (I815150,I814998,I815133);
nor I_47740 (I815167,I815085,I815150);
DFFARX1 I_47741 (I815167,I3563,I814774,I814760,);
nor I_47742 (I815198,I814800,I815133);
DFFARX1 I_47743 (I815198,I3563,I814774,I814745,);
nor I_47744 (I815229,I815077,I815133);
not I_47745 (I815246,I815229);
nand I_47746 (I814754,I815246,I815102);
not I_47747 (I815301,I3570);
DFFARX1 I_47748 (I394463,I3563,I815301,I815327,);
not I_47749 (I815335,I815327);
nand I_47750 (I815352,I394454,I394454);
and I_47751 (I815369,I815352,I394472);
DFFARX1 I_47752 (I815369,I3563,I815301,I815395,);
DFFARX1 I_47753 (I815395,I3563,I815301,I815290,);
DFFARX1 I_47754 (I394475,I3563,I815301,I815426,);
nand I_47755 (I815434,I815426,I394457);
not I_47756 (I815451,I815434);
DFFARX1 I_47757 (I815451,I3563,I815301,I815477,);
not I_47758 (I815485,I815477);
nor I_47759 (I815293,I815335,I815485);
DFFARX1 I_47760 (I394469,I3563,I815301,I815525,);
nor I_47761 (I815284,I815525,I815395);
nor I_47762 (I815275,I815525,I815451);
nand I_47763 (I815561,I394481,I394460);
and I_47764 (I815578,I815561,I394466);
DFFARX1 I_47765 (I815578,I3563,I815301,I815604,);
not I_47766 (I815612,I815604);
nand I_47767 (I815629,I815612,I815525);
nand I_47768 (I815278,I815612,I815434);
nor I_47769 (I815660,I394478,I394460);
and I_47770 (I815677,I815525,I815660);
nor I_47771 (I815694,I815612,I815677);
DFFARX1 I_47772 (I815694,I3563,I815301,I815287,);
nor I_47773 (I815725,I815327,I815660);
DFFARX1 I_47774 (I815725,I3563,I815301,I815272,);
nor I_47775 (I815756,I815604,I815660);
not I_47776 (I815773,I815756);
nand I_47777 (I815281,I815773,I815629);
not I_47778 (I815828,I3570);
DFFARX1 I_47779 (I1045370,I3563,I815828,I815854,);
not I_47780 (I815862,I815854);
nand I_47781 (I815879,I1045385,I1045367);
and I_47782 (I815896,I815879,I1045367);
DFFARX1 I_47783 (I815896,I3563,I815828,I815922,);
DFFARX1 I_47784 (I815922,I3563,I815828,I815817,);
DFFARX1 I_47785 (I1045376,I3563,I815828,I815953,);
nand I_47786 (I815961,I815953,I1045394);
not I_47787 (I815978,I815961);
DFFARX1 I_47788 (I815978,I3563,I815828,I816004,);
not I_47789 (I816012,I816004);
nor I_47790 (I815820,I815862,I816012);
DFFARX1 I_47791 (I1045391,I3563,I815828,I816052,);
nor I_47792 (I815811,I816052,I815922);
nor I_47793 (I815802,I816052,I815978);
nand I_47794 (I816088,I1045388,I1045379);
and I_47795 (I816105,I816088,I1045373);
DFFARX1 I_47796 (I816105,I3563,I815828,I816131,);
not I_47797 (I816139,I816131);
nand I_47798 (I816156,I816139,I816052);
nand I_47799 (I815805,I816139,I815961);
nor I_47800 (I816187,I1045382,I1045379);
and I_47801 (I816204,I816052,I816187);
nor I_47802 (I816221,I816139,I816204);
DFFARX1 I_47803 (I816221,I3563,I815828,I815814,);
nor I_47804 (I816252,I815854,I816187);
DFFARX1 I_47805 (I816252,I3563,I815828,I815799,);
nor I_47806 (I816283,I816131,I816187);
not I_47807 (I816300,I816283);
nand I_47808 (I815808,I816300,I816156);
not I_47809 (I816355,I3570);
DFFARX1 I_47810 (I223814,I3563,I816355,I816381,);
not I_47811 (I816389,I816381);
nand I_47812 (I816406,I223811,I223829);
and I_47813 (I816423,I816406,I223820);
DFFARX1 I_47814 (I816423,I3563,I816355,I816449,);
DFFARX1 I_47815 (I816449,I3563,I816355,I816344,);
DFFARX1 I_47816 (I223826,I3563,I816355,I816480,);
nand I_47817 (I816488,I816480,I223823);
not I_47818 (I816505,I816488);
DFFARX1 I_47819 (I816505,I3563,I816355,I816531,);
not I_47820 (I816539,I816531);
nor I_47821 (I816347,I816389,I816539);
DFFARX1 I_47822 (I223817,I3563,I816355,I816579,);
nor I_47823 (I816338,I816579,I816449);
nor I_47824 (I816329,I816579,I816505);
nand I_47825 (I816615,I223808,I223832);
and I_47826 (I816632,I816615,I223811);
DFFARX1 I_47827 (I816632,I3563,I816355,I816658,);
not I_47828 (I816666,I816658);
nand I_47829 (I816683,I816666,I816579);
nand I_47830 (I816332,I816666,I816488);
nor I_47831 (I816714,I223808,I223832);
and I_47832 (I816731,I816579,I816714);
nor I_47833 (I816748,I816666,I816731);
DFFARX1 I_47834 (I816748,I3563,I816355,I816341,);
nor I_47835 (I816779,I816381,I816714);
DFFARX1 I_47836 (I816779,I3563,I816355,I816326,);
nor I_47837 (I816810,I816658,I816714);
not I_47838 (I816827,I816810);
nand I_47839 (I816335,I816827,I816683);
not I_47840 (I816882,I3570);
DFFARX1 I_47841 (I445800,I3563,I816882,I816908,);
not I_47842 (I816916,I816908);
nand I_47843 (I816933,I445797,I445806);
and I_47844 (I816950,I816933,I445815);
DFFARX1 I_47845 (I816950,I3563,I816882,I816976,);
DFFARX1 I_47846 (I816976,I3563,I816882,I816871,);
DFFARX1 I_47847 (I445818,I3563,I816882,I817007,);
nand I_47848 (I817015,I817007,I445821);
not I_47849 (I817032,I817015);
DFFARX1 I_47850 (I817032,I3563,I816882,I817058,);
not I_47851 (I817066,I817058);
nor I_47852 (I816874,I816916,I817066);
DFFARX1 I_47853 (I445794,I3563,I816882,I817106,);
nor I_47854 (I816865,I817106,I816976);
nor I_47855 (I816856,I817106,I817032);
nand I_47856 (I817142,I445809,I445812);
and I_47857 (I817159,I817142,I445803);
DFFARX1 I_47858 (I817159,I3563,I816882,I817185,);
not I_47859 (I817193,I817185);
nand I_47860 (I817210,I817193,I817106);
nand I_47861 (I816859,I817193,I817015);
nor I_47862 (I817241,I445794,I445812);
and I_47863 (I817258,I817106,I817241);
nor I_47864 (I817275,I817193,I817258);
DFFARX1 I_47865 (I817275,I3563,I816882,I816868,);
nor I_47866 (I817306,I816908,I817241);
DFFARX1 I_47867 (I817306,I3563,I816882,I816853,);
nor I_47868 (I817337,I817185,I817241);
not I_47869 (I817354,I817337);
nand I_47870 (I816862,I817354,I817210);
not I_47871 (I817409,I3570);
DFFARX1 I_47872 (I1209503,I3563,I817409,I817435,);
not I_47873 (I817443,I817435);
nand I_47874 (I817460,I1209485,I1209485);
and I_47875 (I817477,I817460,I1209491);
DFFARX1 I_47876 (I817477,I3563,I817409,I817503,);
DFFARX1 I_47877 (I817503,I3563,I817409,I817398,);
DFFARX1 I_47878 (I1209488,I3563,I817409,I817534,);
nand I_47879 (I817542,I817534,I1209497);
not I_47880 (I817559,I817542);
DFFARX1 I_47881 (I817559,I3563,I817409,I817585,);
not I_47882 (I817593,I817585);
nor I_47883 (I817401,I817443,I817593);
DFFARX1 I_47884 (I1209509,I3563,I817409,I817633,);
nor I_47885 (I817392,I817633,I817503);
nor I_47886 (I817383,I817633,I817559);
nand I_47887 (I817669,I1209500,I1209494);
and I_47888 (I817686,I817669,I1209488);
DFFARX1 I_47889 (I817686,I3563,I817409,I817712,);
not I_47890 (I817720,I817712);
nand I_47891 (I817737,I817720,I817633);
nand I_47892 (I817386,I817720,I817542);
nor I_47893 (I817768,I1209506,I1209494);
and I_47894 (I817785,I817633,I817768);
nor I_47895 (I817802,I817720,I817785);
DFFARX1 I_47896 (I817802,I3563,I817409,I817395,);
nor I_47897 (I817833,I817435,I817768);
DFFARX1 I_47898 (I817833,I3563,I817409,I817380,);
nor I_47899 (I817864,I817712,I817768);
not I_47900 (I817881,I817864);
nand I_47901 (I817389,I817881,I817737);
not I_47902 (I817936,I3570);
DFFARX1 I_47903 (I438184,I3563,I817936,I817962,);
not I_47904 (I817970,I817962);
nand I_47905 (I817987,I438181,I438190);
and I_47906 (I818004,I817987,I438199);
DFFARX1 I_47907 (I818004,I3563,I817936,I818030,);
DFFARX1 I_47908 (I818030,I3563,I817936,I817925,);
DFFARX1 I_47909 (I438202,I3563,I817936,I818061,);
nand I_47910 (I818069,I818061,I438205);
not I_47911 (I818086,I818069);
DFFARX1 I_47912 (I818086,I3563,I817936,I818112,);
not I_47913 (I818120,I818112);
nor I_47914 (I817928,I817970,I818120);
DFFARX1 I_47915 (I438178,I3563,I817936,I818160,);
nor I_47916 (I817919,I818160,I818030);
nor I_47917 (I817910,I818160,I818086);
nand I_47918 (I818196,I438193,I438196);
and I_47919 (I818213,I818196,I438187);
DFFARX1 I_47920 (I818213,I3563,I817936,I818239,);
not I_47921 (I818247,I818239);
nand I_47922 (I818264,I818247,I818160);
nand I_47923 (I817913,I818247,I818069);
nor I_47924 (I818295,I438178,I438196);
and I_47925 (I818312,I818160,I818295);
nor I_47926 (I818329,I818247,I818312);
DFFARX1 I_47927 (I818329,I3563,I817936,I817922,);
nor I_47928 (I818360,I817962,I818295);
DFFARX1 I_47929 (I818360,I3563,I817936,I817907,);
nor I_47930 (I818391,I818239,I818295);
not I_47931 (I818408,I818391);
nand I_47932 (I817916,I818408,I818264);
not I_47933 (I818463,I3570);
DFFARX1 I_47934 (I980124,I3563,I818463,I818489,);
not I_47935 (I818497,I818489);
nand I_47936 (I818514,I980139,I980121);
and I_47937 (I818531,I818514,I980121);
DFFARX1 I_47938 (I818531,I3563,I818463,I818557,);
DFFARX1 I_47939 (I818557,I3563,I818463,I818452,);
DFFARX1 I_47940 (I980130,I3563,I818463,I818588,);
nand I_47941 (I818596,I818588,I980148);
not I_47942 (I818613,I818596);
DFFARX1 I_47943 (I818613,I3563,I818463,I818639,);
not I_47944 (I818647,I818639);
nor I_47945 (I818455,I818497,I818647);
DFFARX1 I_47946 (I980145,I3563,I818463,I818687,);
nor I_47947 (I818446,I818687,I818557);
nor I_47948 (I818437,I818687,I818613);
nand I_47949 (I818723,I980142,I980133);
and I_47950 (I818740,I818723,I980127);
DFFARX1 I_47951 (I818740,I3563,I818463,I818766,);
not I_47952 (I818774,I818766);
nand I_47953 (I818791,I818774,I818687);
nand I_47954 (I818440,I818774,I818596);
nor I_47955 (I818822,I980136,I980133);
and I_47956 (I818839,I818687,I818822);
nor I_47957 (I818856,I818774,I818839);
DFFARX1 I_47958 (I818856,I3563,I818463,I818449,);
nor I_47959 (I818887,I818489,I818822);
DFFARX1 I_47960 (I818887,I3563,I818463,I818434,);
nor I_47961 (I818918,I818766,I818822);
not I_47962 (I818935,I818918);
nand I_47963 (I818443,I818935,I818791);
not I_47964 (I818990,I3570);
DFFARX1 I_47965 (I295387,I3563,I818990,I819016,);
not I_47966 (I819024,I819016);
nand I_47967 (I819041,I295378,I295378);
and I_47968 (I819058,I819041,I295396);
DFFARX1 I_47969 (I819058,I3563,I818990,I819084,);
DFFARX1 I_47970 (I819084,I3563,I818990,I818979,);
DFFARX1 I_47971 (I295399,I3563,I818990,I819115,);
nand I_47972 (I819123,I819115,I295381);
not I_47973 (I819140,I819123);
DFFARX1 I_47974 (I819140,I3563,I818990,I819166,);
not I_47975 (I819174,I819166);
nor I_47976 (I818982,I819024,I819174);
DFFARX1 I_47977 (I295393,I3563,I818990,I819214,);
nor I_47978 (I818973,I819214,I819084);
nor I_47979 (I818964,I819214,I819140);
nand I_47980 (I819250,I295405,I295384);
and I_47981 (I819267,I819250,I295390);
DFFARX1 I_47982 (I819267,I3563,I818990,I819293,);
not I_47983 (I819301,I819293);
nand I_47984 (I819318,I819301,I819214);
nand I_47985 (I818967,I819301,I819123);
nor I_47986 (I819349,I295402,I295384);
and I_47987 (I819366,I819214,I819349);
nor I_47988 (I819383,I819301,I819366);
DFFARX1 I_47989 (I819383,I3563,I818990,I818976,);
nor I_47990 (I819414,I819016,I819349);
DFFARX1 I_47991 (I819414,I3563,I818990,I818961,);
nor I_47992 (I819445,I819293,I819349);
not I_47993 (I819462,I819445);
nand I_47994 (I818970,I819462,I819318);
not I_47995 (I819517,I3570);
DFFARX1 I_47996 (I42427,I3563,I819517,I819543,);
not I_47997 (I819551,I819543);
nand I_47998 (I819568,I42439,I42442);
and I_47999 (I819585,I819568,I42418);
DFFARX1 I_48000 (I819585,I3563,I819517,I819611,);
DFFARX1 I_48001 (I819611,I3563,I819517,I819506,);
DFFARX1 I_48002 (I42436,I3563,I819517,I819642,);
nand I_48003 (I819650,I819642,I42424);
not I_48004 (I819667,I819650);
DFFARX1 I_48005 (I819667,I3563,I819517,I819693,);
not I_48006 (I819701,I819693);
nor I_48007 (I819509,I819551,I819701);
DFFARX1 I_48008 (I42421,I3563,I819517,I819741,);
nor I_48009 (I819500,I819741,I819611);
nor I_48010 (I819491,I819741,I819667);
nand I_48011 (I819777,I42430,I42421);
and I_48012 (I819794,I819777,I42418);
DFFARX1 I_48013 (I819794,I3563,I819517,I819820,);
not I_48014 (I819828,I819820);
nand I_48015 (I819845,I819828,I819741);
nand I_48016 (I819494,I819828,I819650);
nor I_48017 (I819876,I42433,I42421);
and I_48018 (I819893,I819741,I819876);
nor I_48019 (I819910,I819828,I819893);
DFFARX1 I_48020 (I819910,I3563,I819517,I819503,);
nor I_48021 (I819941,I819543,I819876);
DFFARX1 I_48022 (I819941,I3563,I819517,I819488,);
nor I_48023 (I819972,I819820,I819876);
not I_48024 (I819989,I819972);
nand I_48025 (I819497,I819989,I819845);
not I_48026 (I820044,I3570);
DFFARX1 I_48027 (I666505,I3563,I820044,I820070,);
not I_48028 (I820078,I820070);
nand I_48029 (I820095,I666508,I666505);
and I_48030 (I820112,I820095,I666517);
DFFARX1 I_48031 (I820112,I3563,I820044,I820138,);
DFFARX1 I_48032 (I820138,I3563,I820044,I820033,);
DFFARX1 I_48033 (I666514,I3563,I820044,I820169,);
nand I_48034 (I820177,I820169,I666520);
not I_48035 (I820194,I820177);
DFFARX1 I_48036 (I820194,I3563,I820044,I820220,);
not I_48037 (I820228,I820220);
nor I_48038 (I820036,I820078,I820228);
DFFARX1 I_48039 (I666529,I3563,I820044,I820268,);
nor I_48040 (I820027,I820268,I820138);
nor I_48041 (I820018,I820268,I820194);
nand I_48042 (I820304,I666523,I666511);
and I_48043 (I820321,I820304,I666508);
DFFARX1 I_48044 (I820321,I3563,I820044,I820347,);
not I_48045 (I820355,I820347);
nand I_48046 (I820372,I820355,I820268);
nand I_48047 (I820021,I820355,I820177);
nor I_48048 (I820403,I666526,I666511);
and I_48049 (I820420,I820268,I820403);
nor I_48050 (I820437,I820355,I820420);
DFFARX1 I_48051 (I820437,I3563,I820044,I820030,);
nor I_48052 (I820468,I820070,I820403);
DFFARX1 I_48053 (I820468,I3563,I820044,I820015,);
nor I_48054 (I820499,I820347,I820403);
not I_48055 (I820516,I820499);
nand I_48056 (I820024,I820516,I820372);
not I_48057 (I820571,I3570);
DFFARX1 I_48058 (I500200,I3563,I820571,I820597,);
not I_48059 (I820605,I820597);
nand I_48060 (I820622,I500197,I500206);
and I_48061 (I820639,I820622,I500215);
DFFARX1 I_48062 (I820639,I3563,I820571,I820665,);
DFFARX1 I_48063 (I820665,I3563,I820571,I820560,);
DFFARX1 I_48064 (I500218,I3563,I820571,I820696,);
nand I_48065 (I820704,I820696,I500221);
not I_48066 (I820721,I820704);
DFFARX1 I_48067 (I820721,I3563,I820571,I820747,);
not I_48068 (I820755,I820747);
nor I_48069 (I820563,I820605,I820755);
DFFARX1 I_48070 (I500194,I3563,I820571,I820795,);
nor I_48071 (I820554,I820795,I820665);
nor I_48072 (I820545,I820795,I820721);
nand I_48073 (I820831,I500209,I500212);
and I_48074 (I820848,I820831,I500203);
DFFARX1 I_48075 (I820848,I3563,I820571,I820874,);
not I_48076 (I820882,I820874);
nand I_48077 (I820899,I820882,I820795);
nand I_48078 (I820548,I820882,I820704);
nor I_48079 (I820930,I500194,I500212);
and I_48080 (I820947,I820795,I820930);
nor I_48081 (I820964,I820882,I820947);
DFFARX1 I_48082 (I820964,I3563,I820571,I820557,);
nor I_48083 (I820995,I820597,I820930);
DFFARX1 I_48084 (I820995,I3563,I820571,I820542,);
nor I_48085 (I821026,I820874,I820930);
not I_48086 (I821043,I821026);
nand I_48087 (I820551,I821043,I820899);
not I_48088 (I821098,I3570);
DFFARX1 I_48089 (I1264917,I3563,I821098,I821124,);
not I_48090 (I821132,I821124);
nand I_48091 (I821149,I1264923,I1264905);
and I_48092 (I821166,I821149,I1264914);
DFFARX1 I_48093 (I821166,I3563,I821098,I821192,);
DFFARX1 I_48094 (I821192,I3563,I821098,I821087,);
DFFARX1 I_48095 (I1264920,I3563,I821098,I821223,);
nand I_48096 (I821231,I821223,I1264908);
not I_48097 (I821248,I821231);
DFFARX1 I_48098 (I821248,I3563,I821098,I821274,);
not I_48099 (I821282,I821274);
nor I_48100 (I821090,I821132,I821282);
DFFARX1 I_48101 (I1264926,I3563,I821098,I821322,);
nor I_48102 (I821081,I821322,I821192);
nor I_48103 (I821072,I821322,I821248);
nand I_48104 (I821358,I1264905,I1264911);
and I_48105 (I821375,I821358,I1264929);
DFFARX1 I_48106 (I821375,I3563,I821098,I821401,);
not I_48107 (I821409,I821401);
nand I_48108 (I821426,I821409,I821322);
nand I_48109 (I821075,I821409,I821231);
nor I_48110 (I821457,I1264908,I1264911);
and I_48111 (I821474,I821322,I821457);
nor I_48112 (I821491,I821409,I821474);
DFFARX1 I_48113 (I821491,I3563,I821098,I821084,);
nor I_48114 (I821522,I821124,I821457);
DFFARX1 I_48115 (I821522,I3563,I821098,I821069,);
nor I_48116 (I821553,I821401,I821457);
not I_48117 (I821570,I821553);
nand I_48118 (I821078,I821570,I821426);
not I_48119 (I821625,I3570);
DFFARX1 I_48120 (I406584,I3563,I821625,I821651,);
not I_48121 (I821659,I821651);
nand I_48122 (I821676,I406575,I406575);
and I_48123 (I821693,I821676,I406593);
DFFARX1 I_48124 (I821693,I3563,I821625,I821719,);
DFFARX1 I_48125 (I821719,I3563,I821625,I821614,);
DFFARX1 I_48126 (I406596,I3563,I821625,I821750,);
nand I_48127 (I821758,I821750,I406578);
not I_48128 (I821775,I821758);
DFFARX1 I_48129 (I821775,I3563,I821625,I821801,);
not I_48130 (I821809,I821801);
nor I_48131 (I821617,I821659,I821809);
DFFARX1 I_48132 (I406590,I3563,I821625,I821849,);
nor I_48133 (I821608,I821849,I821719);
nor I_48134 (I821599,I821849,I821775);
nand I_48135 (I821885,I406602,I406581);
and I_48136 (I821902,I821885,I406587);
DFFARX1 I_48137 (I821902,I3563,I821625,I821928,);
not I_48138 (I821936,I821928);
nand I_48139 (I821953,I821936,I821849);
nand I_48140 (I821602,I821936,I821758);
nor I_48141 (I821984,I406599,I406581);
and I_48142 (I822001,I821849,I821984);
nor I_48143 (I822018,I821936,I822001);
DFFARX1 I_48144 (I822018,I3563,I821625,I821611,);
nor I_48145 (I822049,I821651,I821984);
DFFARX1 I_48146 (I822049,I3563,I821625,I821596,);
nor I_48147 (I822080,I821928,I821984);
not I_48148 (I822097,I822080);
nand I_48149 (I821605,I822097,I821953);
not I_48150 (I822152,I3570);
DFFARX1 I_48151 (I1138987,I3563,I822152,I822178,);
not I_48152 (I822186,I822178);
nand I_48153 (I822203,I1138969,I1138969);
and I_48154 (I822220,I822203,I1138975);
DFFARX1 I_48155 (I822220,I3563,I822152,I822246,);
DFFARX1 I_48156 (I822246,I3563,I822152,I822141,);
DFFARX1 I_48157 (I1138972,I3563,I822152,I822277,);
nand I_48158 (I822285,I822277,I1138981);
not I_48159 (I822302,I822285);
DFFARX1 I_48160 (I822302,I3563,I822152,I822328,);
not I_48161 (I822336,I822328);
nor I_48162 (I822144,I822186,I822336);
DFFARX1 I_48163 (I1138993,I3563,I822152,I822376,);
nor I_48164 (I822135,I822376,I822246);
nor I_48165 (I822126,I822376,I822302);
nand I_48166 (I822412,I1138984,I1138978);
and I_48167 (I822429,I822412,I1138972);
DFFARX1 I_48168 (I822429,I3563,I822152,I822455,);
not I_48169 (I822463,I822455);
nand I_48170 (I822480,I822463,I822376);
nand I_48171 (I822129,I822463,I822285);
nor I_48172 (I822511,I1138990,I1138978);
and I_48173 (I822528,I822376,I822511);
nor I_48174 (I822545,I822463,I822528);
DFFARX1 I_48175 (I822545,I3563,I822152,I822138,);
nor I_48176 (I822576,I822178,I822511);
DFFARX1 I_48177 (I822576,I3563,I822152,I822123,);
nor I_48178 (I822607,I822455,I822511);
not I_48179 (I822624,I822607);
nand I_48180 (I822132,I822624,I822480);
not I_48181 (I822679,I3570);
DFFARX1 I_48182 (I32414,I3563,I822679,I822705,);
not I_48183 (I822713,I822705);
nand I_48184 (I822730,I32426,I32429);
and I_48185 (I822747,I822730,I32405);
DFFARX1 I_48186 (I822747,I3563,I822679,I822773,);
DFFARX1 I_48187 (I822773,I3563,I822679,I822668,);
DFFARX1 I_48188 (I32423,I3563,I822679,I822804,);
nand I_48189 (I822812,I822804,I32411);
not I_48190 (I822829,I822812);
DFFARX1 I_48191 (I822829,I3563,I822679,I822855,);
not I_48192 (I822863,I822855);
nor I_48193 (I822671,I822713,I822863);
DFFARX1 I_48194 (I32408,I3563,I822679,I822903,);
nor I_48195 (I822662,I822903,I822773);
nor I_48196 (I822653,I822903,I822829);
nand I_48197 (I822939,I32417,I32408);
and I_48198 (I822956,I822939,I32405);
DFFARX1 I_48199 (I822956,I3563,I822679,I822982,);
not I_48200 (I822990,I822982);
nand I_48201 (I823007,I822990,I822903);
nand I_48202 (I822656,I822990,I822812);
nor I_48203 (I823038,I32420,I32408);
and I_48204 (I823055,I822903,I823038);
nor I_48205 (I823072,I822990,I823055);
DFFARX1 I_48206 (I823072,I3563,I822679,I822665,);
nor I_48207 (I823103,I822705,I823038);
DFFARX1 I_48208 (I823103,I3563,I822679,I822650,);
nor I_48209 (I823134,I822982,I823038);
not I_48210 (I823151,I823134);
nand I_48211 (I822659,I823151,I823007);
not I_48212 (I823206,I3570);
DFFARX1 I_48213 (I1094481,I3563,I823206,I823232,);
not I_48214 (I823240,I823232);
nand I_48215 (I823257,I1094463,I1094463);
and I_48216 (I823274,I823257,I1094469);
DFFARX1 I_48217 (I823274,I3563,I823206,I823300,);
DFFARX1 I_48218 (I823300,I3563,I823206,I823195,);
DFFARX1 I_48219 (I1094466,I3563,I823206,I823331,);
nand I_48220 (I823339,I823331,I1094475);
not I_48221 (I823356,I823339);
DFFARX1 I_48222 (I823356,I3563,I823206,I823382,);
not I_48223 (I823390,I823382);
nor I_48224 (I823198,I823240,I823390);
DFFARX1 I_48225 (I1094487,I3563,I823206,I823430,);
nor I_48226 (I823189,I823430,I823300);
nor I_48227 (I823180,I823430,I823356);
nand I_48228 (I823466,I1094478,I1094472);
and I_48229 (I823483,I823466,I1094466);
DFFARX1 I_48230 (I823483,I3563,I823206,I823509,);
not I_48231 (I823517,I823509);
nand I_48232 (I823534,I823517,I823430);
nand I_48233 (I823183,I823517,I823339);
nor I_48234 (I823565,I1094484,I1094472);
and I_48235 (I823582,I823430,I823565);
nor I_48236 (I823599,I823517,I823582);
DFFARX1 I_48237 (I823599,I3563,I823206,I823192,);
nor I_48238 (I823630,I823232,I823565);
DFFARX1 I_48239 (I823630,I3563,I823206,I823177,);
nor I_48240 (I823661,I823509,I823565);
not I_48241 (I823678,I823661);
nand I_48242 (I823186,I823678,I823534);
not I_48243 (I823733,I3570);
DFFARX1 I_48244 (I112533,I3563,I823733,I823759,);
not I_48245 (I823767,I823759);
nand I_48246 (I823784,I112509,I112518);
and I_48247 (I823801,I823784,I112512);
DFFARX1 I_48248 (I823801,I3563,I823733,I823827,);
DFFARX1 I_48249 (I823827,I3563,I823733,I823722,);
DFFARX1 I_48250 (I112530,I3563,I823733,I823858,);
nand I_48251 (I823866,I823858,I112521);
not I_48252 (I823883,I823866);
DFFARX1 I_48253 (I823883,I3563,I823733,I823909,);
not I_48254 (I823917,I823909);
nor I_48255 (I823725,I823767,I823917);
DFFARX1 I_48256 (I112515,I3563,I823733,I823957,);
nor I_48257 (I823716,I823957,I823827);
nor I_48258 (I823707,I823957,I823883);
nand I_48259 (I823993,I112527,I112524);
and I_48260 (I824010,I823993,I112512);
DFFARX1 I_48261 (I824010,I3563,I823733,I824036,);
not I_48262 (I824044,I824036);
nand I_48263 (I824061,I824044,I823957);
nand I_48264 (I823710,I824044,I823866);
nor I_48265 (I824092,I112509,I112524);
and I_48266 (I824109,I823957,I824092);
nor I_48267 (I824126,I824044,I824109);
DFFARX1 I_48268 (I824126,I3563,I823733,I823719,);
nor I_48269 (I824157,I823759,I824092);
DFFARX1 I_48270 (I824157,I3563,I823733,I823704,);
nor I_48271 (I824188,I824036,I824092);
not I_48272 (I824205,I824188);
nand I_48273 (I823713,I824205,I824061);
not I_48274 (I824260,I3570);
DFFARX1 I_48275 (I804647,I3563,I824260,I824286,);
not I_48276 (I824294,I824286);
nand I_48277 (I824311,I804650,I804647);
and I_48278 (I824328,I824311,I804659);
DFFARX1 I_48279 (I824328,I3563,I824260,I824354,);
DFFARX1 I_48280 (I824354,I3563,I824260,I824249,);
DFFARX1 I_48281 (I804656,I3563,I824260,I824385,);
nand I_48282 (I824393,I824385,I804662);
not I_48283 (I824410,I824393);
DFFARX1 I_48284 (I824410,I3563,I824260,I824436,);
not I_48285 (I824444,I824436);
nor I_48286 (I824252,I824294,I824444);
DFFARX1 I_48287 (I804671,I3563,I824260,I824484,);
nor I_48288 (I824243,I824484,I824354);
nor I_48289 (I824234,I824484,I824410);
nand I_48290 (I824520,I804665,I804653);
and I_48291 (I824537,I824520,I804650);
DFFARX1 I_48292 (I824537,I3563,I824260,I824563,);
not I_48293 (I824571,I824563);
nand I_48294 (I824588,I824571,I824484);
nand I_48295 (I824237,I824571,I824393);
nor I_48296 (I824619,I804668,I804653);
and I_48297 (I824636,I824484,I824619);
nor I_48298 (I824653,I824571,I824636);
DFFARX1 I_48299 (I824653,I3563,I824260,I824246,);
nor I_48300 (I824684,I824286,I824619);
DFFARX1 I_48301 (I824684,I3563,I824260,I824231,);
nor I_48302 (I824715,I824563,I824619);
not I_48303 (I824732,I824715);
nand I_48304 (I824240,I824732,I824588);
not I_48305 (I824787,I3570);
DFFARX1 I_48306 (I135721,I3563,I824787,I824813,);
not I_48307 (I824821,I824813);
nand I_48308 (I824838,I135697,I135706);
and I_48309 (I824855,I824838,I135700);
DFFARX1 I_48310 (I824855,I3563,I824787,I824881,);
DFFARX1 I_48311 (I824881,I3563,I824787,I824776,);
DFFARX1 I_48312 (I135718,I3563,I824787,I824912,);
nand I_48313 (I824920,I824912,I135709);
not I_48314 (I824937,I824920);
DFFARX1 I_48315 (I824937,I3563,I824787,I824963,);
not I_48316 (I824971,I824963);
nor I_48317 (I824779,I824821,I824971);
DFFARX1 I_48318 (I135703,I3563,I824787,I825011,);
nor I_48319 (I824770,I825011,I824881);
nor I_48320 (I824761,I825011,I824937);
nand I_48321 (I825047,I135715,I135712);
and I_48322 (I825064,I825047,I135700);
DFFARX1 I_48323 (I825064,I3563,I824787,I825090,);
not I_48324 (I825098,I825090);
nand I_48325 (I825115,I825098,I825011);
nand I_48326 (I824764,I825098,I824920);
nor I_48327 (I825146,I135697,I135712);
and I_48328 (I825163,I825011,I825146);
nor I_48329 (I825180,I825098,I825163);
DFFARX1 I_48330 (I825180,I3563,I824787,I824773,);
nor I_48331 (I825211,I824813,I825146);
DFFARX1 I_48332 (I825211,I3563,I824787,I824758,);
nor I_48333 (I825242,I825090,I825146);
not I_48334 (I825259,I825242);
nand I_48335 (I824767,I825259,I825115);
not I_48336 (I825314,I3570);
DFFARX1 I_48337 (I4778,I3563,I825314,I825340,);
not I_48338 (I825348,I825340);
nand I_48339 (I825365,I4784,I4766);
and I_48340 (I825382,I825365,I4775);
DFFARX1 I_48341 (I825382,I3563,I825314,I825408,);
DFFARX1 I_48342 (I825408,I3563,I825314,I825303,);
DFFARX1 I_48343 (I4766,I3563,I825314,I825439,);
nand I_48344 (I825447,I825439,I4769);
not I_48345 (I825464,I825447);
DFFARX1 I_48346 (I825464,I3563,I825314,I825490,);
not I_48347 (I825498,I825490);
nor I_48348 (I825306,I825348,I825498);
DFFARX1 I_48349 (I4769,I3563,I825314,I825538,);
nor I_48350 (I825297,I825538,I825408);
nor I_48351 (I825288,I825538,I825464);
nand I_48352 (I825574,I4772,I4781);
and I_48353 (I825591,I825574,I4763);
DFFARX1 I_48354 (I825591,I3563,I825314,I825617,);
not I_48355 (I825625,I825617);
nand I_48356 (I825642,I825625,I825538);
nand I_48357 (I825291,I825625,I825447);
nor I_48358 (I825673,I4763,I4781);
and I_48359 (I825690,I825538,I825673);
nor I_48360 (I825707,I825625,I825690);
DFFARX1 I_48361 (I825707,I3563,I825314,I825300,);
nor I_48362 (I825738,I825340,I825673);
DFFARX1 I_48363 (I825738,I3563,I825314,I825285,);
nor I_48364 (I825769,I825617,I825673);
not I_48365 (I825786,I825769);
nand I_48366 (I825294,I825786,I825642);
not I_48367 (I825841,I3570);
DFFARX1 I_48368 (I373383,I3563,I825841,I825867,);
not I_48369 (I825875,I825867);
nand I_48370 (I825892,I373374,I373374);
and I_48371 (I825909,I825892,I373392);
DFFARX1 I_48372 (I825909,I3563,I825841,I825935,);
DFFARX1 I_48373 (I825935,I3563,I825841,I825830,);
DFFARX1 I_48374 (I373395,I3563,I825841,I825966,);
nand I_48375 (I825974,I825966,I373377);
not I_48376 (I825991,I825974);
DFFARX1 I_48377 (I825991,I3563,I825841,I826017,);
not I_48378 (I826025,I826017);
nor I_48379 (I825833,I825875,I826025);
DFFARX1 I_48380 (I373389,I3563,I825841,I826065,);
nor I_48381 (I825824,I826065,I825935);
nor I_48382 (I825815,I826065,I825991);
nand I_48383 (I826101,I373401,I373380);
and I_48384 (I826118,I826101,I373386);
DFFARX1 I_48385 (I826118,I3563,I825841,I826144,);
not I_48386 (I826152,I826144);
nand I_48387 (I826169,I826152,I826065);
nand I_48388 (I825818,I826152,I825974);
nor I_48389 (I826200,I373398,I373380);
and I_48390 (I826217,I826065,I826200);
nor I_48391 (I826234,I826152,I826217);
DFFARX1 I_48392 (I826234,I3563,I825841,I825827,);
nor I_48393 (I826265,I825867,I826200);
DFFARX1 I_48394 (I826265,I3563,I825841,I825812,);
nor I_48395 (I826296,I826144,I826200);
not I_48396 (I826313,I826296);
nand I_48397 (I825821,I826313,I826169);
not I_48398 (I826368,I3570);
DFFARX1 I_48399 (I388139,I3563,I826368,I826394,);
not I_48400 (I826402,I826394);
nand I_48401 (I826419,I388130,I388130);
and I_48402 (I826436,I826419,I388148);
DFFARX1 I_48403 (I826436,I3563,I826368,I826462,);
DFFARX1 I_48404 (I826462,I3563,I826368,I826357,);
DFFARX1 I_48405 (I388151,I3563,I826368,I826493,);
nand I_48406 (I826501,I826493,I388133);
not I_48407 (I826518,I826501);
DFFARX1 I_48408 (I826518,I3563,I826368,I826544,);
not I_48409 (I826552,I826544);
nor I_48410 (I826360,I826402,I826552);
DFFARX1 I_48411 (I388145,I3563,I826368,I826592,);
nor I_48412 (I826351,I826592,I826462);
nor I_48413 (I826342,I826592,I826518);
nand I_48414 (I826628,I388157,I388136);
and I_48415 (I826645,I826628,I388142);
DFFARX1 I_48416 (I826645,I3563,I826368,I826671,);
not I_48417 (I826679,I826671);
nand I_48418 (I826696,I826679,I826592);
nand I_48419 (I826345,I826679,I826501);
nor I_48420 (I826727,I388154,I388136);
and I_48421 (I826744,I826592,I826727);
nor I_48422 (I826761,I826679,I826744);
DFFARX1 I_48423 (I826761,I3563,I826368,I826354,);
nor I_48424 (I826792,I826394,I826727);
DFFARX1 I_48425 (I826792,I3563,I826368,I826339,);
nor I_48426 (I826823,I826671,I826727);
not I_48427 (I826840,I826823);
nand I_48428 (I826348,I826840,I826696);
not I_48429 (I826895,I3570);
DFFARX1 I_48430 (I963328,I3563,I826895,I826921,);
not I_48431 (I826929,I826921);
nand I_48432 (I826946,I963343,I963325);
and I_48433 (I826963,I826946,I963325);
DFFARX1 I_48434 (I826963,I3563,I826895,I826989,);
DFFARX1 I_48435 (I826989,I3563,I826895,I826884,);
DFFARX1 I_48436 (I963334,I3563,I826895,I827020,);
nand I_48437 (I827028,I827020,I963352);
not I_48438 (I827045,I827028);
DFFARX1 I_48439 (I827045,I3563,I826895,I827071,);
not I_48440 (I827079,I827071);
nor I_48441 (I826887,I826929,I827079);
DFFARX1 I_48442 (I963349,I3563,I826895,I827119,);
nor I_48443 (I826878,I827119,I826989);
nor I_48444 (I826869,I827119,I827045);
nand I_48445 (I827155,I963346,I963337);
and I_48446 (I827172,I827155,I963331);
DFFARX1 I_48447 (I827172,I3563,I826895,I827198,);
not I_48448 (I827206,I827198);
nand I_48449 (I827223,I827206,I827119);
nand I_48450 (I826872,I827206,I827028);
nor I_48451 (I827254,I963340,I963337);
and I_48452 (I827271,I827119,I827254);
nor I_48453 (I827288,I827206,I827271);
DFFARX1 I_48454 (I827288,I3563,I826895,I826881,);
nor I_48455 (I827319,I826921,I827254);
DFFARX1 I_48456 (I827319,I3563,I826895,I826866,);
nor I_48457 (I827350,I827198,I827254);
not I_48458 (I827367,I827350);
nand I_48459 (I826875,I827367,I827223);
not I_48460 (I827422,I3570);
DFFARX1 I_48461 (I1405323,I3563,I827422,I827448,);
not I_48462 (I827456,I827448);
nand I_48463 (I827473,I1405320,I1405329);
and I_48464 (I827490,I827473,I1405308);
DFFARX1 I_48465 (I827490,I3563,I827422,I827516,);
DFFARX1 I_48466 (I827516,I3563,I827422,I827411,);
DFFARX1 I_48467 (I1405311,I3563,I827422,I827547,);
nand I_48468 (I827555,I827547,I1405326);
not I_48469 (I827572,I827555);
DFFARX1 I_48470 (I827572,I3563,I827422,I827598,);
not I_48471 (I827606,I827598);
nor I_48472 (I827414,I827456,I827606);
DFFARX1 I_48473 (I1405332,I3563,I827422,I827646,);
nor I_48474 (I827405,I827646,I827516);
nor I_48475 (I827396,I827646,I827572);
nand I_48476 (I827682,I1405314,I1405335);
and I_48477 (I827699,I827682,I1405317);
DFFARX1 I_48478 (I827699,I3563,I827422,I827725,);
not I_48479 (I827733,I827725);
nand I_48480 (I827750,I827733,I827646);
nand I_48481 (I827399,I827733,I827555);
nor I_48482 (I827781,I1405308,I1405335);
and I_48483 (I827798,I827646,I827781);
nor I_48484 (I827815,I827733,I827798);
DFFARX1 I_48485 (I827815,I3563,I827422,I827408,);
nor I_48486 (I827846,I827448,I827781);
DFFARX1 I_48487 (I827846,I3563,I827422,I827393,);
nor I_48488 (I827877,I827725,I827781);
not I_48489 (I827894,I827877);
nand I_48490 (I827402,I827894,I827750);
not I_48491 (I827949,I3570);
DFFARX1 I_48492 (I1211815,I3563,I827949,I827975,);
not I_48493 (I827983,I827975);
nand I_48494 (I828000,I1211797,I1211797);
and I_48495 (I828017,I828000,I1211803);
DFFARX1 I_48496 (I828017,I3563,I827949,I828043,);
DFFARX1 I_48497 (I828043,I3563,I827949,I827938,);
DFFARX1 I_48498 (I1211800,I3563,I827949,I828074,);
nand I_48499 (I828082,I828074,I1211809);
not I_48500 (I828099,I828082);
DFFARX1 I_48501 (I828099,I3563,I827949,I828125,);
not I_48502 (I828133,I828125);
nor I_48503 (I827941,I827983,I828133);
DFFARX1 I_48504 (I1211821,I3563,I827949,I828173,);
nor I_48505 (I827932,I828173,I828043);
nor I_48506 (I827923,I828173,I828099);
nand I_48507 (I828209,I1211812,I1211806);
and I_48508 (I828226,I828209,I1211800);
DFFARX1 I_48509 (I828226,I3563,I827949,I828252,);
not I_48510 (I828260,I828252);
nand I_48511 (I828277,I828260,I828173);
nand I_48512 (I827926,I828260,I828082);
nor I_48513 (I828308,I1211818,I1211806);
and I_48514 (I828325,I828173,I828308);
nor I_48515 (I828342,I828260,I828325);
DFFARX1 I_48516 (I828342,I3563,I827949,I827935,);
nor I_48517 (I828373,I827975,I828308);
DFFARX1 I_48518 (I828373,I3563,I827949,I827920,);
nor I_48519 (I828404,I828252,I828308);
not I_48520 (I828421,I828404);
nand I_48521 (I827929,I828421,I828277);
not I_48522 (I828476,I3570);
DFFARX1 I_48523 (I592536,I3563,I828476,I828502,);
not I_48524 (I828510,I828502);
nand I_48525 (I828527,I592521,I592542);
and I_48526 (I828544,I828527,I592530);
DFFARX1 I_48527 (I828544,I3563,I828476,I828570,);
DFFARX1 I_48528 (I828570,I3563,I828476,I828465,);
DFFARX1 I_48529 (I592524,I3563,I828476,I828601,);
nand I_48530 (I828609,I828601,I592533);
not I_48531 (I828626,I828609);
DFFARX1 I_48532 (I828626,I3563,I828476,I828652,);
not I_48533 (I828660,I828652);
nor I_48534 (I828468,I828510,I828660);
DFFARX1 I_48535 (I592539,I3563,I828476,I828700,);
nor I_48536 (I828459,I828700,I828570);
nor I_48537 (I828450,I828700,I828626);
nand I_48538 (I828736,I592521,I592524);
and I_48539 (I828753,I828736,I592545);
DFFARX1 I_48540 (I828753,I3563,I828476,I828779,);
not I_48541 (I828787,I828779);
nand I_48542 (I828804,I828787,I828700);
nand I_48543 (I828453,I828787,I828609);
nor I_48544 (I828835,I592527,I592524);
and I_48545 (I828852,I828700,I828835);
nor I_48546 (I828869,I828787,I828852);
DFFARX1 I_48547 (I828869,I3563,I828476,I828462,);
nor I_48548 (I828900,I828502,I828835);
DFFARX1 I_48549 (I828900,I3563,I828476,I828447,);
nor I_48550 (I828931,I828779,I828835);
not I_48551 (I828948,I828931);
nand I_48552 (I828456,I828948,I828804);
not I_48553 (I829003,I3570);
DFFARX1 I_48554 (I1305111,I3563,I829003,I829029,);
not I_48555 (I829037,I829029);
nand I_48556 (I829054,I1305093,I1305096);
and I_48557 (I829071,I829054,I1305108);
DFFARX1 I_48558 (I829071,I3563,I829003,I829097,);
DFFARX1 I_48559 (I829097,I3563,I829003,I828992,);
DFFARX1 I_48560 (I1305117,I3563,I829003,I829128,);
nand I_48561 (I829136,I829128,I1305102);
not I_48562 (I829153,I829136);
DFFARX1 I_48563 (I829153,I3563,I829003,I829179,);
not I_48564 (I829187,I829179);
nor I_48565 (I828995,I829037,I829187);
DFFARX1 I_48566 (I1305114,I3563,I829003,I829227,);
nor I_48567 (I828986,I829227,I829097);
nor I_48568 (I828977,I829227,I829153);
nand I_48569 (I829263,I1305105,I1305099);
and I_48570 (I829280,I829263,I1305093);
DFFARX1 I_48571 (I829280,I3563,I829003,I829306,);
not I_48572 (I829314,I829306);
nand I_48573 (I829331,I829314,I829227);
nand I_48574 (I828980,I829314,I829136);
nor I_48575 (I829362,I1305096,I1305099);
and I_48576 (I829379,I829227,I829362);
nor I_48577 (I829396,I829314,I829379);
DFFARX1 I_48578 (I829396,I3563,I829003,I828989,);
nor I_48579 (I829427,I829029,I829362);
DFFARX1 I_48580 (I829427,I3563,I829003,I828974,);
nor I_48581 (I829458,I829306,I829362);
not I_48582 (I829475,I829458);
nand I_48583 (I828983,I829475,I829331);
not I_48584 (I829530,I3570);
DFFARX1 I_48585 (I333331,I3563,I829530,I829556,);
not I_48586 (I829564,I829556);
nand I_48587 (I829581,I333322,I333322);
and I_48588 (I829598,I829581,I333340);
DFFARX1 I_48589 (I829598,I3563,I829530,I829624,);
DFFARX1 I_48590 (I829624,I3563,I829530,I829519,);
DFFARX1 I_48591 (I333343,I3563,I829530,I829655,);
nand I_48592 (I829663,I829655,I333325);
not I_48593 (I829680,I829663);
DFFARX1 I_48594 (I829680,I3563,I829530,I829706,);
not I_48595 (I829714,I829706);
nor I_48596 (I829522,I829564,I829714);
DFFARX1 I_48597 (I333337,I3563,I829530,I829754,);
nor I_48598 (I829513,I829754,I829624);
nor I_48599 (I829504,I829754,I829680);
nand I_48600 (I829790,I333349,I333328);
and I_48601 (I829807,I829790,I333334);
DFFARX1 I_48602 (I829807,I3563,I829530,I829833,);
not I_48603 (I829841,I829833);
nand I_48604 (I829858,I829841,I829754);
nand I_48605 (I829507,I829841,I829663);
nor I_48606 (I829889,I333346,I333328);
and I_48607 (I829906,I829754,I829889);
nor I_48608 (I829923,I829841,I829906);
DFFARX1 I_48609 (I829923,I3563,I829530,I829516,);
nor I_48610 (I829954,I829556,I829889);
DFFARX1 I_48611 (I829954,I3563,I829530,I829501,);
nor I_48612 (I829985,I829833,I829889);
not I_48613 (I830002,I829985);
nand I_48614 (I829510,I830002,I829858);
not I_48615 (I830057,I3570);
DFFARX1 I_48616 (I366005,I3563,I830057,I830083,);
not I_48617 (I830091,I830083);
nand I_48618 (I830108,I365996,I365996);
and I_48619 (I830125,I830108,I366014);
DFFARX1 I_48620 (I830125,I3563,I830057,I830151,);
DFFARX1 I_48621 (I830151,I3563,I830057,I830046,);
DFFARX1 I_48622 (I366017,I3563,I830057,I830182,);
nand I_48623 (I830190,I830182,I365999);
not I_48624 (I830207,I830190);
DFFARX1 I_48625 (I830207,I3563,I830057,I830233,);
not I_48626 (I830241,I830233);
nor I_48627 (I830049,I830091,I830241);
DFFARX1 I_48628 (I366011,I3563,I830057,I830281,);
nor I_48629 (I830040,I830281,I830151);
nor I_48630 (I830031,I830281,I830207);
nand I_48631 (I830317,I366023,I366002);
and I_48632 (I830334,I830317,I366008);
DFFARX1 I_48633 (I830334,I3563,I830057,I830360,);
not I_48634 (I830368,I830360);
nand I_48635 (I830385,I830368,I830281);
nand I_48636 (I830034,I830368,I830190);
nor I_48637 (I830416,I366020,I366002);
and I_48638 (I830433,I830281,I830416);
nor I_48639 (I830450,I830368,I830433);
DFFARX1 I_48640 (I830450,I3563,I830057,I830043,);
nor I_48641 (I830481,I830083,I830416);
DFFARX1 I_48642 (I830481,I3563,I830057,I830028,);
nor I_48643 (I830512,I830360,I830416);
not I_48644 (I830529,I830512);
nand I_48645 (I830037,I830529,I830385);
not I_48646 (I830584,I3570);
DFFARX1 I_48647 (I345979,I3563,I830584,I830610,);
not I_48648 (I830618,I830610);
nand I_48649 (I830635,I345970,I345970);
and I_48650 (I830652,I830635,I345988);
DFFARX1 I_48651 (I830652,I3563,I830584,I830678,);
DFFARX1 I_48652 (I830678,I3563,I830584,I830573,);
DFFARX1 I_48653 (I345991,I3563,I830584,I830709,);
nand I_48654 (I830717,I830709,I345973);
not I_48655 (I830734,I830717);
DFFARX1 I_48656 (I830734,I3563,I830584,I830760,);
not I_48657 (I830768,I830760);
nor I_48658 (I830576,I830618,I830768);
DFFARX1 I_48659 (I345985,I3563,I830584,I830808,);
nor I_48660 (I830567,I830808,I830678);
nor I_48661 (I830558,I830808,I830734);
nand I_48662 (I830844,I345997,I345976);
and I_48663 (I830861,I830844,I345982);
DFFARX1 I_48664 (I830861,I3563,I830584,I830887,);
not I_48665 (I830895,I830887);
nand I_48666 (I830912,I830895,I830808);
nand I_48667 (I830561,I830895,I830717);
nor I_48668 (I830943,I345994,I345976);
and I_48669 (I830960,I830808,I830943);
nor I_48670 (I830977,I830895,I830960);
DFFARX1 I_48671 (I830977,I3563,I830584,I830570,);
nor I_48672 (I831008,I830610,I830943);
DFFARX1 I_48673 (I831008,I3563,I830584,I830555,);
nor I_48674 (I831039,I830887,I830943);
not I_48675 (I831056,I831039);
nand I_48676 (I830564,I831056,I830912);
not I_48677 (I831111,I3570);
DFFARX1 I_48678 (I1104307,I3563,I831111,I831137,);
not I_48679 (I831145,I831137);
nand I_48680 (I831162,I1104289,I1104289);
and I_48681 (I831179,I831162,I1104295);
DFFARX1 I_48682 (I831179,I3563,I831111,I831205,);
DFFARX1 I_48683 (I831205,I3563,I831111,I831100,);
DFFARX1 I_48684 (I1104292,I3563,I831111,I831236,);
nand I_48685 (I831244,I831236,I1104301);
not I_48686 (I831261,I831244);
DFFARX1 I_48687 (I831261,I3563,I831111,I831287,);
not I_48688 (I831295,I831287);
nor I_48689 (I831103,I831145,I831295);
DFFARX1 I_48690 (I1104313,I3563,I831111,I831335,);
nor I_48691 (I831094,I831335,I831205);
nor I_48692 (I831085,I831335,I831261);
nand I_48693 (I831371,I1104304,I1104298);
and I_48694 (I831388,I831371,I1104292);
DFFARX1 I_48695 (I831388,I3563,I831111,I831414,);
not I_48696 (I831422,I831414);
nand I_48697 (I831439,I831422,I831335);
nand I_48698 (I831088,I831422,I831244);
nor I_48699 (I831470,I1104310,I1104298);
and I_48700 (I831487,I831335,I831470);
nor I_48701 (I831504,I831422,I831487);
DFFARX1 I_48702 (I831504,I3563,I831111,I831097,);
nor I_48703 (I831535,I831137,I831470);
DFFARX1 I_48704 (I831535,I3563,I831111,I831082,);
nor I_48705 (I831566,I831414,I831470);
not I_48706 (I831583,I831566);
nand I_48707 (I831091,I831583,I831439);
not I_48708 (I831638,I3570);
DFFARX1 I_48709 (I943948,I3563,I831638,I831664,);
not I_48710 (I831672,I831664);
nand I_48711 (I831689,I943963,I943945);
and I_48712 (I831706,I831689,I943945);
DFFARX1 I_48713 (I831706,I3563,I831638,I831732,);
DFFARX1 I_48714 (I831732,I3563,I831638,I831627,);
DFFARX1 I_48715 (I943954,I3563,I831638,I831763,);
nand I_48716 (I831771,I831763,I943972);
not I_48717 (I831788,I831771);
DFFARX1 I_48718 (I831788,I3563,I831638,I831814,);
not I_48719 (I831822,I831814);
nor I_48720 (I831630,I831672,I831822);
DFFARX1 I_48721 (I943969,I3563,I831638,I831862,);
nor I_48722 (I831621,I831862,I831732);
nor I_48723 (I831612,I831862,I831788);
nand I_48724 (I831898,I943966,I943957);
and I_48725 (I831915,I831898,I943951);
DFFARX1 I_48726 (I831915,I3563,I831638,I831941,);
not I_48727 (I831949,I831941);
nand I_48728 (I831966,I831949,I831862);
nand I_48729 (I831615,I831949,I831771);
nor I_48730 (I831997,I943960,I943957);
and I_48731 (I832014,I831862,I831997);
nor I_48732 (I832031,I831949,I832014);
DFFARX1 I_48733 (I832031,I3563,I831638,I831624,);
nor I_48734 (I832062,I831664,I831997);
DFFARX1 I_48735 (I832062,I3563,I831638,I831609,);
nor I_48736 (I832093,I831941,I831997);
not I_48737 (I832110,I832093);
nand I_48738 (I831618,I832110,I831966);
not I_48739 (I832165,I3570);
DFFARX1 I_48740 (I340182,I3563,I832165,I832191,);
not I_48741 (I832199,I832191);
nand I_48742 (I832216,I340173,I340173);
and I_48743 (I832233,I832216,I340191);
DFFARX1 I_48744 (I832233,I3563,I832165,I832259,);
DFFARX1 I_48745 (I832259,I3563,I832165,I832154,);
DFFARX1 I_48746 (I340194,I3563,I832165,I832290,);
nand I_48747 (I832298,I832290,I340176);
not I_48748 (I832315,I832298);
DFFARX1 I_48749 (I832315,I3563,I832165,I832341,);
not I_48750 (I832349,I832341);
nor I_48751 (I832157,I832199,I832349);
DFFARX1 I_48752 (I340188,I3563,I832165,I832389,);
nor I_48753 (I832148,I832389,I832259);
nor I_48754 (I832139,I832389,I832315);
nand I_48755 (I832425,I340200,I340179);
and I_48756 (I832442,I832425,I340185);
DFFARX1 I_48757 (I832442,I3563,I832165,I832468,);
not I_48758 (I832476,I832468);
nand I_48759 (I832493,I832476,I832389);
nand I_48760 (I832142,I832476,I832298);
nor I_48761 (I832524,I340197,I340179);
and I_48762 (I832541,I832389,I832524);
nor I_48763 (I832558,I832476,I832541);
DFFARX1 I_48764 (I832558,I3563,I832165,I832151,);
nor I_48765 (I832589,I832191,I832524);
DFFARX1 I_48766 (I832589,I3563,I832165,I832136,);
nor I_48767 (I832620,I832468,I832524);
not I_48768 (I832637,I832620);
nand I_48769 (I832145,I832637,I832493);
not I_48770 (I832692,I3570);
DFFARX1 I_48771 (I462664,I3563,I832692,I832718,);
not I_48772 (I832726,I832718);
nand I_48773 (I832743,I462661,I462670);
and I_48774 (I832760,I832743,I462679);
DFFARX1 I_48775 (I832760,I3563,I832692,I832786,);
DFFARX1 I_48776 (I832786,I3563,I832692,I832681,);
DFFARX1 I_48777 (I462682,I3563,I832692,I832817,);
nand I_48778 (I832825,I832817,I462685);
not I_48779 (I832842,I832825);
DFFARX1 I_48780 (I832842,I3563,I832692,I832868,);
not I_48781 (I832876,I832868);
nor I_48782 (I832684,I832726,I832876);
DFFARX1 I_48783 (I462658,I3563,I832692,I832916,);
nor I_48784 (I832675,I832916,I832786);
nor I_48785 (I832666,I832916,I832842);
nand I_48786 (I832952,I462673,I462676);
and I_48787 (I832969,I832952,I462667);
DFFARX1 I_48788 (I832969,I3563,I832692,I832995,);
not I_48789 (I833003,I832995);
nand I_48790 (I833020,I833003,I832916);
nand I_48791 (I832669,I833003,I832825);
nor I_48792 (I833051,I462658,I462676);
and I_48793 (I833068,I832916,I833051);
nor I_48794 (I833085,I833003,I833068);
DFFARX1 I_48795 (I833085,I3563,I832692,I832678,);
nor I_48796 (I833116,I832718,I833051);
DFFARX1 I_48797 (I833116,I3563,I832692,I832663,);
nor I_48798 (I833147,I832995,I833051);
not I_48799 (I833164,I833147);
nand I_48800 (I832672,I833164,I833020);
not I_48801 (I833219,I3570);
DFFARX1 I_48802 (I1167309,I3563,I833219,I833245,);
not I_48803 (I833253,I833245);
nand I_48804 (I833270,I1167291,I1167291);
and I_48805 (I833287,I833270,I1167297);
DFFARX1 I_48806 (I833287,I3563,I833219,I833313,);
DFFARX1 I_48807 (I833313,I3563,I833219,I833208,);
DFFARX1 I_48808 (I1167294,I3563,I833219,I833344,);
nand I_48809 (I833352,I833344,I1167303);
not I_48810 (I833369,I833352);
DFFARX1 I_48811 (I833369,I3563,I833219,I833395,);
not I_48812 (I833403,I833395);
nor I_48813 (I833211,I833253,I833403);
DFFARX1 I_48814 (I1167315,I3563,I833219,I833443,);
nor I_48815 (I833202,I833443,I833313);
nor I_48816 (I833193,I833443,I833369);
nand I_48817 (I833479,I1167306,I1167300);
and I_48818 (I833496,I833479,I1167294);
DFFARX1 I_48819 (I833496,I3563,I833219,I833522,);
not I_48820 (I833530,I833522);
nand I_48821 (I833547,I833530,I833443);
nand I_48822 (I833196,I833530,I833352);
nor I_48823 (I833578,I1167312,I1167300);
and I_48824 (I833595,I833443,I833578);
nor I_48825 (I833612,I833530,I833595);
DFFARX1 I_48826 (I833612,I3563,I833219,I833205,);
nor I_48827 (I833643,I833245,I833578);
DFFARX1 I_48828 (I833643,I3563,I833219,I833190,);
nor I_48829 (I833674,I833522,I833578);
not I_48830 (I833691,I833674);
nand I_48831 (I833199,I833691,I833547);
not I_48832 (I833746,I3570);
DFFARX1 I_48833 (I298022,I3563,I833746,I833772,);
not I_48834 (I833780,I833772);
nand I_48835 (I833797,I298013,I298013);
and I_48836 (I833814,I833797,I298031);
DFFARX1 I_48837 (I833814,I3563,I833746,I833840,);
DFFARX1 I_48838 (I833840,I3563,I833746,I833735,);
DFFARX1 I_48839 (I298034,I3563,I833746,I833871,);
nand I_48840 (I833879,I833871,I298016);
not I_48841 (I833896,I833879);
DFFARX1 I_48842 (I833896,I3563,I833746,I833922,);
not I_48843 (I833930,I833922);
nor I_48844 (I833738,I833780,I833930);
DFFARX1 I_48845 (I298028,I3563,I833746,I833970,);
nor I_48846 (I833729,I833970,I833840);
nor I_48847 (I833720,I833970,I833896);
nand I_48848 (I834006,I298040,I298019);
and I_48849 (I834023,I834006,I298025);
DFFARX1 I_48850 (I834023,I3563,I833746,I834049,);
not I_48851 (I834057,I834049);
nand I_48852 (I834074,I834057,I833970);
nand I_48853 (I833723,I834057,I833879);
nor I_48854 (I834105,I298037,I298019);
and I_48855 (I834122,I833970,I834105);
nor I_48856 (I834139,I834057,I834122);
DFFARX1 I_48857 (I834139,I3563,I833746,I833732,);
nor I_48858 (I834170,I833772,I834105);
DFFARX1 I_48859 (I834170,I3563,I833746,I833717,);
nor I_48860 (I834201,I834049,I834105);
not I_48861 (I834218,I834201);
nand I_48862 (I833726,I834218,I834074);
not I_48863 (I834273,I3570);
DFFARX1 I_48864 (I1269813,I3563,I834273,I834299,);
not I_48865 (I834307,I834299);
nand I_48866 (I834324,I1269819,I1269801);
and I_48867 (I834341,I834324,I1269810);
DFFARX1 I_48868 (I834341,I3563,I834273,I834367,);
DFFARX1 I_48869 (I834367,I3563,I834273,I834262,);
DFFARX1 I_48870 (I1269816,I3563,I834273,I834398,);
nand I_48871 (I834406,I834398,I1269804);
not I_48872 (I834423,I834406);
DFFARX1 I_48873 (I834423,I3563,I834273,I834449,);
not I_48874 (I834457,I834449);
nor I_48875 (I834265,I834307,I834457);
DFFARX1 I_48876 (I1269822,I3563,I834273,I834497,);
nor I_48877 (I834256,I834497,I834367);
nor I_48878 (I834247,I834497,I834423);
nand I_48879 (I834533,I1269801,I1269807);
and I_48880 (I834550,I834533,I1269825);
DFFARX1 I_48881 (I834550,I3563,I834273,I834576,);
not I_48882 (I834584,I834576);
nand I_48883 (I834601,I834584,I834497);
nand I_48884 (I834250,I834584,I834406);
nor I_48885 (I834632,I1269804,I1269807);
and I_48886 (I834649,I834497,I834632);
nor I_48887 (I834666,I834584,I834649);
DFFARX1 I_48888 (I834666,I3563,I834273,I834259,);
nor I_48889 (I834697,I834299,I834632);
DFFARX1 I_48890 (I834697,I3563,I834273,I834244,);
nor I_48891 (I834728,I834576,I834632);
not I_48892 (I834745,I834728);
nand I_48893 (I834253,I834745,I834601);
not I_48894 (I834800,I3570);
DFFARX1 I_48895 (I1009194,I3563,I834800,I834826,);
not I_48896 (I834834,I834826);
nand I_48897 (I834851,I1009209,I1009191);
and I_48898 (I834868,I834851,I1009191);
DFFARX1 I_48899 (I834868,I3563,I834800,I834894,);
DFFARX1 I_48900 (I834894,I3563,I834800,I834789,);
DFFARX1 I_48901 (I1009200,I3563,I834800,I834925,);
nand I_48902 (I834933,I834925,I1009218);
not I_48903 (I834950,I834933);
DFFARX1 I_48904 (I834950,I3563,I834800,I834976,);
not I_48905 (I834984,I834976);
nor I_48906 (I834792,I834834,I834984);
DFFARX1 I_48907 (I1009215,I3563,I834800,I835024,);
nor I_48908 (I834783,I835024,I834894);
nor I_48909 (I834774,I835024,I834950);
nand I_48910 (I835060,I1009212,I1009203);
and I_48911 (I835077,I835060,I1009197);
DFFARX1 I_48912 (I835077,I3563,I834800,I835103,);
not I_48913 (I835111,I835103);
nand I_48914 (I835128,I835111,I835024);
nand I_48915 (I834777,I835111,I834933);
nor I_48916 (I835159,I1009206,I1009203);
and I_48917 (I835176,I835024,I835159);
nor I_48918 (I835193,I835111,I835176);
DFFARX1 I_48919 (I835193,I3563,I834800,I834786,);
nor I_48920 (I835224,I834826,I835159);
DFFARX1 I_48921 (I835224,I3563,I834800,I834771,);
nor I_48922 (I835255,I835103,I835159);
not I_48923 (I835272,I835255);
nand I_48924 (I834780,I835272,I835128);
not I_48925 (I835327,I3570);
DFFARX1 I_48926 (I1019530,I3563,I835327,I835353,);
not I_48927 (I835361,I835353);
nand I_48928 (I835378,I1019545,I1019527);
and I_48929 (I835395,I835378,I1019527);
DFFARX1 I_48930 (I835395,I3563,I835327,I835421,);
DFFARX1 I_48931 (I835421,I3563,I835327,I835316,);
DFFARX1 I_48932 (I1019536,I3563,I835327,I835452,);
nand I_48933 (I835460,I835452,I1019554);
not I_48934 (I835477,I835460);
DFFARX1 I_48935 (I835477,I3563,I835327,I835503,);
not I_48936 (I835511,I835503);
nor I_48937 (I835319,I835361,I835511);
DFFARX1 I_48938 (I1019551,I3563,I835327,I835551,);
nor I_48939 (I835310,I835551,I835421);
nor I_48940 (I835301,I835551,I835477);
nand I_48941 (I835587,I1019548,I1019539);
and I_48942 (I835604,I835587,I1019533);
DFFARX1 I_48943 (I835604,I3563,I835327,I835630,);
not I_48944 (I835638,I835630);
nand I_48945 (I835655,I835638,I835551);
nand I_48946 (I835304,I835638,I835460);
nor I_48947 (I835686,I1019542,I1019539);
and I_48948 (I835703,I835551,I835686);
nor I_48949 (I835720,I835638,I835703);
DFFARX1 I_48950 (I835720,I3563,I835327,I835313,);
nor I_48951 (I835751,I835353,I835686);
DFFARX1 I_48952 (I835751,I3563,I835327,I835298,);
nor I_48953 (I835782,I835630,I835686);
not I_48954 (I835799,I835782);
nand I_48955 (I835307,I835799,I835655);
not I_48956 (I835854,I3570);
DFFARX1 I_48957 (I781527,I3563,I835854,I835880,);
not I_48958 (I835888,I835880);
nand I_48959 (I835905,I781530,I781527);
and I_48960 (I835922,I835905,I781539);
DFFARX1 I_48961 (I835922,I3563,I835854,I835948,);
DFFARX1 I_48962 (I835948,I3563,I835854,I835843,);
DFFARX1 I_48963 (I781536,I3563,I835854,I835979,);
nand I_48964 (I835987,I835979,I781542);
not I_48965 (I836004,I835987);
DFFARX1 I_48966 (I836004,I3563,I835854,I836030,);
not I_48967 (I836038,I836030);
nor I_48968 (I835846,I835888,I836038);
DFFARX1 I_48969 (I781551,I3563,I835854,I836078,);
nor I_48970 (I835837,I836078,I835948);
nor I_48971 (I835828,I836078,I836004);
nand I_48972 (I836114,I781545,I781533);
and I_48973 (I836131,I836114,I781530);
DFFARX1 I_48974 (I836131,I3563,I835854,I836157,);
not I_48975 (I836165,I836157);
nand I_48976 (I836182,I836165,I836078);
nand I_48977 (I835831,I836165,I835987);
nor I_48978 (I836213,I781548,I781533);
and I_48979 (I836230,I836078,I836213);
nor I_48980 (I836247,I836165,I836230);
DFFARX1 I_48981 (I836247,I3563,I835854,I835840,);
nor I_48982 (I836278,I835880,I836213);
DFFARX1 I_48983 (I836278,I3563,I835854,I835825,);
nor I_48984 (I836309,I836157,I836213);
not I_48985 (I836326,I836309);
nand I_48986 (I835834,I836326,I836182);
not I_48987 (I836381,I3570);
DFFARX1 I_48988 (I380761,I3563,I836381,I836407,);
not I_48989 (I836415,I836407);
nand I_48990 (I836432,I380752,I380752);
and I_48991 (I836449,I836432,I380770);
DFFARX1 I_48992 (I836449,I3563,I836381,I836475,);
DFFARX1 I_48993 (I836475,I3563,I836381,I836370,);
DFFARX1 I_48994 (I380773,I3563,I836381,I836506,);
nand I_48995 (I836514,I836506,I380755);
not I_48996 (I836531,I836514);
DFFARX1 I_48997 (I836531,I3563,I836381,I836557,);
not I_48998 (I836565,I836557);
nor I_48999 (I836373,I836415,I836565);
DFFARX1 I_49000 (I380767,I3563,I836381,I836605,);
nor I_49001 (I836364,I836605,I836475);
nor I_49002 (I836355,I836605,I836531);
nand I_49003 (I836641,I380779,I380758);
and I_49004 (I836658,I836641,I380764);
DFFARX1 I_49005 (I836658,I3563,I836381,I836684,);
not I_49006 (I836692,I836684);
nand I_49007 (I836709,I836692,I836605);
nand I_49008 (I836358,I836692,I836514);
nor I_49009 (I836740,I380776,I380758);
and I_49010 (I836757,I836605,I836740);
nor I_49011 (I836774,I836692,I836757);
DFFARX1 I_49012 (I836774,I3563,I836381,I836367,);
nor I_49013 (I836805,I836407,I836740);
DFFARX1 I_49014 (I836805,I3563,I836381,I836352,);
nor I_49015 (I836836,I836684,I836740);
not I_49016 (I836853,I836836);
nand I_49017 (I836361,I836853,I836709);
not I_49018 (I836908,I3570);
DFFARX1 I_49019 (I320683,I3563,I836908,I836934,);
not I_49020 (I836942,I836934);
nand I_49021 (I836959,I320674,I320674);
and I_49022 (I836976,I836959,I320692);
DFFARX1 I_49023 (I836976,I3563,I836908,I837002,);
DFFARX1 I_49024 (I837002,I3563,I836908,I836897,);
DFFARX1 I_49025 (I320695,I3563,I836908,I837033,);
nand I_49026 (I837041,I837033,I320677);
not I_49027 (I837058,I837041);
DFFARX1 I_49028 (I837058,I3563,I836908,I837084,);
not I_49029 (I837092,I837084);
nor I_49030 (I836900,I836942,I837092);
DFFARX1 I_49031 (I320689,I3563,I836908,I837132,);
nor I_49032 (I836891,I837132,I837002);
nor I_49033 (I836882,I837132,I837058);
nand I_49034 (I837168,I320701,I320680);
and I_49035 (I837185,I837168,I320686);
DFFARX1 I_49036 (I837185,I3563,I836908,I837211,);
not I_49037 (I837219,I837211);
nand I_49038 (I837236,I837219,I837132);
nand I_49039 (I836885,I837219,I837041);
nor I_49040 (I837267,I320698,I320680);
and I_49041 (I837284,I837132,I837267);
nor I_49042 (I837301,I837219,I837284);
DFFARX1 I_49043 (I837301,I3563,I836908,I836894,);
nor I_49044 (I837332,I836934,I837267);
DFFARX1 I_49045 (I837332,I3563,I836908,I836879,);
nor I_49046 (I837363,I837211,I837267);
not I_49047 (I837380,I837363);
nand I_49048 (I836888,I837380,I837236);
not I_49049 (I837435,I3570);
DFFARX1 I_49050 (I1171355,I3563,I837435,I837461,);
not I_49051 (I837469,I837461);
nand I_49052 (I837486,I1171337,I1171337);
and I_49053 (I837503,I837486,I1171343);
DFFARX1 I_49054 (I837503,I3563,I837435,I837529,);
DFFARX1 I_49055 (I837529,I3563,I837435,I837424,);
DFFARX1 I_49056 (I1171340,I3563,I837435,I837560,);
nand I_49057 (I837568,I837560,I1171349);
not I_49058 (I837585,I837568);
DFFARX1 I_49059 (I837585,I3563,I837435,I837611,);
not I_49060 (I837619,I837611);
nor I_49061 (I837427,I837469,I837619);
DFFARX1 I_49062 (I1171361,I3563,I837435,I837659,);
nor I_49063 (I837418,I837659,I837529);
nor I_49064 (I837409,I837659,I837585);
nand I_49065 (I837695,I1171352,I1171346);
and I_49066 (I837712,I837695,I1171340);
DFFARX1 I_49067 (I837712,I3563,I837435,I837738,);
not I_49068 (I837746,I837738);
nand I_49069 (I837763,I837746,I837659);
nand I_49070 (I837412,I837746,I837568);
nor I_49071 (I837794,I1171358,I1171346);
and I_49072 (I837811,I837659,I837794);
nor I_49073 (I837828,I837746,I837811);
DFFARX1 I_49074 (I837828,I3563,I837435,I837421,);
nor I_49075 (I837859,I837461,I837794);
DFFARX1 I_49076 (I837859,I3563,I837435,I837406,);
nor I_49077 (I837890,I837738,I837794);
not I_49078 (I837907,I837890);
nand I_49079 (I837415,I837907,I837763);
not I_49080 (I837962,I3570);
DFFARX1 I_49081 (I1396398,I3563,I837962,I837988,);
not I_49082 (I837996,I837988);
nand I_49083 (I838013,I1396395,I1396404);
and I_49084 (I838030,I838013,I1396383);
DFFARX1 I_49085 (I838030,I3563,I837962,I838056,);
DFFARX1 I_49086 (I838056,I3563,I837962,I837951,);
DFFARX1 I_49087 (I1396386,I3563,I837962,I838087,);
nand I_49088 (I838095,I838087,I1396401);
not I_49089 (I838112,I838095);
DFFARX1 I_49090 (I838112,I3563,I837962,I838138,);
not I_49091 (I838146,I838138);
nor I_49092 (I837954,I837996,I838146);
DFFARX1 I_49093 (I1396407,I3563,I837962,I838186,);
nor I_49094 (I837945,I838186,I838056);
nor I_49095 (I837936,I838186,I838112);
nand I_49096 (I838222,I1396389,I1396410);
and I_49097 (I838239,I838222,I1396392);
DFFARX1 I_49098 (I838239,I3563,I837962,I838265,);
not I_49099 (I838273,I838265);
nand I_49100 (I838290,I838273,I838186);
nand I_49101 (I837939,I838273,I838095);
nor I_49102 (I838321,I1396383,I1396410);
and I_49103 (I838338,I838186,I838321);
nor I_49104 (I838355,I838273,I838338);
DFFARX1 I_49105 (I838355,I3563,I837962,I837948,);
nor I_49106 (I838386,I837988,I838321);
DFFARX1 I_49107 (I838386,I3563,I837962,I837933,);
nor I_49108 (I838417,I838265,I838321);
not I_49109 (I838434,I838417);
nand I_49110 (I837942,I838434,I838290);
not I_49111 (I838489,I3570);
DFFARX1 I_49112 (I652070,I3563,I838489,I838515,);
not I_49113 (I838523,I838515);
nand I_49114 (I838540,I652055,I652076);
and I_49115 (I838557,I838540,I652064);
DFFARX1 I_49116 (I838557,I3563,I838489,I838583,);
DFFARX1 I_49117 (I838583,I3563,I838489,I838478,);
DFFARX1 I_49118 (I652058,I3563,I838489,I838614,);
nand I_49119 (I838622,I838614,I652067);
not I_49120 (I838639,I838622);
DFFARX1 I_49121 (I838639,I3563,I838489,I838665,);
not I_49122 (I838673,I838665);
nor I_49123 (I838481,I838523,I838673);
DFFARX1 I_49124 (I652073,I3563,I838489,I838713,);
nor I_49125 (I838472,I838713,I838583);
nor I_49126 (I838463,I838713,I838639);
nand I_49127 (I838749,I652055,I652058);
and I_49128 (I838766,I838749,I652079);
DFFARX1 I_49129 (I838766,I3563,I838489,I838792,);
not I_49130 (I838800,I838792);
nand I_49131 (I838817,I838800,I838713);
nand I_49132 (I838466,I838800,I838622);
nor I_49133 (I838848,I652061,I652058);
and I_49134 (I838865,I838713,I838848);
nor I_49135 (I838882,I838800,I838865);
DFFARX1 I_49136 (I838882,I3563,I838489,I838475,);
nor I_49137 (I838913,I838515,I838848);
DFFARX1 I_49138 (I838913,I3563,I838489,I838460,);
nor I_49139 (I838944,I838792,I838848);
not I_49140 (I838961,I838944);
nand I_49141 (I838469,I838961,I838817);
not I_49142 (I839016,I3570);
DFFARX1 I_49143 (I245829,I3563,I839016,I839042,);
not I_49144 (I839050,I839042);
nand I_49145 (I839067,I245826,I245844);
and I_49146 (I839084,I839067,I245835);
DFFARX1 I_49147 (I839084,I3563,I839016,I839110,);
DFFARX1 I_49148 (I839110,I3563,I839016,I839005,);
DFFARX1 I_49149 (I245841,I3563,I839016,I839141,);
nand I_49150 (I839149,I839141,I245838);
not I_49151 (I839166,I839149);
DFFARX1 I_49152 (I839166,I3563,I839016,I839192,);
not I_49153 (I839200,I839192);
nor I_49154 (I839008,I839050,I839200);
DFFARX1 I_49155 (I245832,I3563,I839016,I839240,);
nor I_49156 (I838999,I839240,I839110);
nor I_49157 (I838990,I839240,I839166);
nand I_49158 (I839276,I245823,I245847);
and I_49159 (I839293,I839276,I245826);
DFFARX1 I_49160 (I839293,I3563,I839016,I839319,);
not I_49161 (I839327,I839319);
nand I_49162 (I839344,I839327,I839240);
nand I_49163 (I838993,I839327,I839149);
nor I_49164 (I839375,I245823,I245847);
and I_49165 (I839392,I839240,I839375);
nor I_49166 (I839409,I839327,I839392);
DFFARX1 I_49167 (I839409,I3563,I839016,I839002,);
nor I_49168 (I839440,I839042,I839375);
DFFARX1 I_49169 (I839440,I3563,I839016,I838987,);
nor I_49170 (I839471,I839319,I839375);
not I_49171 (I839488,I839471);
nand I_49172 (I838996,I839488,I839344);
not I_49173 (I839543,I3570);
DFFARX1 I_49174 (I2772,I3563,I839543,I839569,);
not I_49175 (I839577,I839569);
nand I_49176 (I839594,I1700,I3052);
and I_49177 (I839611,I839594,I1780);
DFFARX1 I_49178 (I839611,I3563,I839543,I839637,);
DFFARX1 I_49179 (I839637,I3563,I839543,I839532,);
DFFARX1 I_49180 (I2260,I3563,I839543,I839668,);
nand I_49181 (I839676,I839668,I3084);
not I_49182 (I839693,I839676);
DFFARX1 I_49183 (I839693,I3563,I839543,I839719,);
not I_49184 (I839727,I839719);
nor I_49185 (I839535,I839577,I839727);
DFFARX1 I_49186 (I2204,I3563,I839543,I839767,);
nor I_49187 (I839526,I839767,I839637);
nor I_49188 (I839517,I839767,I839693);
nand I_49189 (I839803,I2324,I2932);
and I_49190 (I839820,I839803,I2836);
DFFARX1 I_49191 (I839820,I3563,I839543,I839846,);
not I_49192 (I839854,I839846);
nand I_49193 (I839871,I839854,I839767);
nand I_49194 (I839520,I839854,I839676);
nor I_49195 (I839902,I1764,I2932);
and I_49196 (I839919,I839767,I839902);
nor I_49197 (I839936,I839854,I839919);
DFFARX1 I_49198 (I839936,I3563,I839543,I839529,);
nor I_49199 (I839967,I839569,I839902);
DFFARX1 I_49200 (I839967,I3563,I839543,I839514,);
nor I_49201 (I839998,I839846,I839902);
not I_49202 (I840015,I839998);
nand I_49203 (I839523,I840015,I839871);
not I_49204 (I840070,I3570);
DFFARX1 I_49205 (I448520,I3563,I840070,I840096,);
not I_49206 (I840104,I840096);
nand I_49207 (I840121,I448517,I448526);
and I_49208 (I840138,I840121,I448535);
DFFARX1 I_49209 (I840138,I3563,I840070,I840164,);
DFFARX1 I_49210 (I840164,I3563,I840070,I840059,);
DFFARX1 I_49211 (I448538,I3563,I840070,I840195,);
nand I_49212 (I840203,I840195,I448541);
not I_49213 (I840220,I840203);
DFFARX1 I_49214 (I840220,I3563,I840070,I840246,);
not I_49215 (I840254,I840246);
nor I_49216 (I840062,I840104,I840254);
DFFARX1 I_49217 (I448514,I3563,I840070,I840294,);
nor I_49218 (I840053,I840294,I840164);
nor I_49219 (I840044,I840294,I840220);
nand I_49220 (I840330,I448529,I448532);
and I_49221 (I840347,I840330,I448523);
DFFARX1 I_49222 (I840347,I3563,I840070,I840373,);
not I_49223 (I840381,I840373);
nand I_49224 (I840398,I840381,I840294);
nand I_49225 (I840047,I840381,I840203);
nor I_49226 (I840429,I448514,I448532);
and I_49227 (I840446,I840294,I840429);
nor I_49228 (I840463,I840381,I840446);
DFFARX1 I_49229 (I840463,I3563,I840070,I840056,);
nor I_49230 (I840494,I840096,I840429);
DFFARX1 I_49231 (I840494,I3563,I840070,I840041,);
nor I_49232 (I840525,I840373,I840429);
not I_49233 (I840542,I840525);
nand I_49234 (I840050,I840542,I840398);
not I_49235 (I840597,I3570);
DFFARX1 I_49236 (I1048912,I3563,I840597,I840623,);
not I_49237 (I840631,I840623);
nand I_49238 (I840648,I1048921,I1048909);
and I_49239 (I840665,I840648,I1048906);
DFFARX1 I_49240 (I840665,I3563,I840597,I840691,);
DFFARX1 I_49241 (I840691,I3563,I840597,I840586,);
DFFARX1 I_49242 (I1048906,I3563,I840597,I840722,);
nand I_49243 (I840730,I840722,I1048903);
not I_49244 (I840747,I840730);
DFFARX1 I_49245 (I840747,I3563,I840597,I840773,);
not I_49246 (I840781,I840773);
nor I_49247 (I840589,I840631,I840781);
DFFARX1 I_49248 (I1048909,I3563,I840597,I840821,);
nor I_49249 (I840580,I840821,I840691);
nor I_49250 (I840571,I840821,I840747);
nand I_49251 (I840857,I1048924,I1048915);
and I_49252 (I840874,I840857,I1048918);
DFFARX1 I_49253 (I840874,I3563,I840597,I840900,);
not I_49254 (I840908,I840900);
nand I_49255 (I840925,I840908,I840821);
nand I_49256 (I840574,I840908,I840730);
nor I_49257 (I840956,I1048903,I1048915);
and I_49258 (I840973,I840821,I840956);
nor I_49259 (I840990,I840908,I840973);
DFFARX1 I_49260 (I840990,I3563,I840597,I840583,);
nor I_49261 (I841021,I840623,I840956);
DFFARX1 I_49262 (I841021,I3563,I840597,I840568,);
nor I_49263 (I841052,I840900,I840956);
not I_49264 (I841069,I841052);
nand I_49265 (I840577,I841069,I840925);
not I_49266 (I841124,I3570);
DFFARX1 I_49267 (I354411,I3563,I841124,I841150,);
not I_49268 (I841158,I841150);
nand I_49269 (I841175,I354402,I354402);
and I_49270 (I841192,I841175,I354420);
DFFARX1 I_49271 (I841192,I3563,I841124,I841218,);
DFFARX1 I_49272 (I841218,I3563,I841124,I841113,);
DFFARX1 I_49273 (I354423,I3563,I841124,I841249,);
nand I_49274 (I841257,I841249,I354405);
not I_49275 (I841274,I841257);
DFFARX1 I_49276 (I841274,I3563,I841124,I841300,);
not I_49277 (I841308,I841300);
nor I_49278 (I841116,I841158,I841308);
DFFARX1 I_49279 (I354417,I3563,I841124,I841348,);
nor I_49280 (I841107,I841348,I841218);
nor I_49281 (I841098,I841348,I841274);
nand I_49282 (I841384,I354429,I354408);
and I_49283 (I841401,I841384,I354414);
DFFARX1 I_49284 (I841401,I3563,I841124,I841427,);
not I_49285 (I841435,I841427);
nand I_49286 (I841452,I841435,I841348);
nand I_49287 (I841101,I841435,I841257);
nor I_49288 (I841483,I354426,I354408);
and I_49289 (I841500,I841348,I841483);
nor I_49290 (I841517,I841435,I841500);
DFFARX1 I_49291 (I841517,I3563,I841124,I841110,);
nor I_49292 (I841548,I841150,I841483);
DFFARX1 I_49293 (I841548,I3563,I841124,I841095,);
nor I_49294 (I841579,I841427,I841483);
not I_49295 (I841596,I841579);
nand I_49296 (I841104,I841596,I841452);
not I_49297 (I841651,I3570);
DFFARX1 I_49298 (I1318983,I3563,I841651,I841677,);
not I_49299 (I841685,I841677);
nand I_49300 (I841702,I1318965,I1318968);
and I_49301 (I841719,I841702,I1318980);
DFFARX1 I_49302 (I841719,I3563,I841651,I841745,);
DFFARX1 I_49303 (I841745,I3563,I841651,I841640,);
DFFARX1 I_49304 (I1318989,I3563,I841651,I841776,);
nand I_49305 (I841784,I841776,I1318974);
not I_49306 (I841801,I841784);
DFFARX1 I_49307 (I841801,I3563,I841651,I841827,);
not I_49308 (I841835,I841827);
nor I_49309 (I841643,I841685,I841835);
DFFARX1 I_49310 (I1318986,I3563,I841651,I841875,);
nor I_49311 (I841634,I841875,I841745);
nor I_49312 (I841625,I841875,I841801);
nand I_49313 (I841911,I1318977,I1318971);
and I_49314 (I841928,I841911,I1318965);
DFFARX1 I_49315 (I841928,I3563,I841651,I841954,);
not I_49316 (I841962,I841954);
nand I_49317 (I841979,I841962,I841875);
nand I_49318 (I841628,I841962,I841784);
nor I_49319 (I842010,I1318968,I1318971);
and I_49320 (I842027,I841875,I842010);
nor I_49321 (I842044,I841962,I842027);
DFFARX1 I_49322 (I842044,I3563,I841651,I841637,);
nor I_49323 (I842075,I841677,I842010);
DFFARX1 I_49324 (I842075,I3563,I841651,I841622,);
nor I_49325 (I842106,I841954,I842010);
not I_49326 (I842123,I842106);
nand I_49327 (I841631,I842123,I841979);
not I_49328 (I842178,I3570);
DFFARX1 I_49329 (I922630,I3563,I842178,I842204,);
not I_49330 (I842212,I842204);
nand I_49331 (I842229,I922645,I922627);
and I_49332 (I842246,I842229,I922627);
DFFARX1 I_49333 (I842246,I3563,I842178,I842272,);
DFFARX1 I_49334 (I842272,I3563,I842178,I842167,);
DFFARX1 I_49335 (I922636,I3563,I842178,I842303,);
nand I_49336 (I842311,I842303,I922654);
not I_49337 (I842328,I842311);
DFFARX1 I_49338 (I842328,I3563,I842178,I842354,);
not I_49339 (I842362,I842354);
nor I_49340 (I842170,I842212,I842362);
DFFARX1 I_49341 (I922651,I3563,I842178,I842402,);
nor I_49342 (I842161,I842402,I842272);
nor I_49343 (I842152,I842402,I842328);
nand I_49344 (I842438,I922648,I922639);
and I_49345 (I842455,I842438,I922633);
DFFARX1 I_49346 (I842455,I3563,I842178,I842481,);
not I_49347 (I842489,I842481);
nand I_49348 (I842506,I842489,I842402);
nand I_49349 (I842155,I842489,I842311);
nor I_49350 (I842537,I922642,I922639);
and I_49351 (I842554,I842402,I842537);
nor I_49352 (I842571,I842489,I842554);
DFFARX1 I_49353 (I842571,I3563,I842178,I842164,);
nor I_49354 (I842602,I842204,I842537);
DFFARX1 I_49355 (I842602,I3563,I842178,I842149,);
nor I_49356 (I842633,I842481,I842537);
not I_49357 (I842650,I842633);
nand I_49358 (I842158,I842650,I842506);
not I_49359 (I842705,I3570);
DFFARX1 I_49360 (I30833,I3563,I842705,I842731,);
not I_49361 (I842739,I842731);
nand I_49362 (I842756,I30845,I30848);
and I_49363 (I842773,I842756,I30824);
DFFARX1 I_49364 (I842773,I3563,I842705,I842799,);
DFFARX1 I_49365 (I842799,I3563,I842705,I842694,);
DFFARX1 I_49366 (I30842,I3563,I842705,I842830,);
nand I_49367 (I842838,I842830,I30830);
not I_49368 (I842855,I842838);
DFFARX1 I_49369 (I842855,I3563,I842705,I842881,);
not I_49370 (I842889,I842881);
nor I_49371 (I842697,I842739,I842889);
DFFARX1 I_49372 (I30827,I3563,I842705,I842929,);
nor I_49373 (I842688,I842929,I842799);
nor I_49374 (I842679,I842929,I842855);
nand I_49375 (I842965,I30836,I30827);
and I_49376 (I842982,I842965,I30824);
DFFARX1 I_49377 (I842982,I3563,I842705,I843008,);
not I_49378 (I843016,I843008);
nand I_49379 (I843033,I843016,I842929);
nand I_49380 (I842682,I843016,I842838);
nor I_49381 (I843064,I30839,I30827);
and I_49382 (I843081,I842929,I843064);
nor I_49383 (I843098,I843016,I843081);
DFFARX1 I_49384 (I843098,I3563,I842705,I842691,);
nor I_49385 (I843129,I842731,I843064);
DFFARX1 I_49386 (I843129,I3563,I842705,I842676,);
nor I_49387 (I843160,I843008,I843064);
not I_49388 (I843177,I843160);
nand I_49389 (I842685,I843177,I843033);
not I_49390 (I843232,I3570);
DFFARX1 I_49391 (I1076962,I3563,I843232,I843258,);
not I_49392 (I843266,I843258);
nand I_49393 (I843283,I1076971,I1076959);
and I_49394 (I843300,I843283,I1076956);
DFFARX1 I_49395 (I843300,I3563,I843232,I843326,);
DFFARX1 I_49396 (I843326,I3563,I843232,I843221,);
DFFARX1 I_49397 (I1076956,I3563,I843232,I843357,);
nand I_49398 (I843365,I843357,I1076953);
not I_49399 (I843382,I843365);
DFFARX1 I_49400 (I843382,I3563,I843232,I843408,);
not I_49401 (I843416,I843408);
nor I_49402 (I843224,I843266,I843416);
DFFARX1 I_49403 (I1076959,I3563,I843232,I843456,);
nor I_49404 (I843215,I843456,I843326);
nor I_49405 (I843206,I843456,I843382);
nand I_49406 (I843492,I1076974,I1076965);
and I_49407 (I843509,I843492,I1076968);
DFFARX1 I_49408 (I843509,I3563,I843232,I843535,);
not I_49409 (I843543,I843535);
nand I_49410 (I843560,I843543,I843456);
nand I_49411 (I843209,I843543,I843365);
nor I_49412 (I843591,I1076953,I1076965);
and I_49413 (I843608,I843456,I843591);
nor I_49414 (I843625,I843543,I843608);
DFFARX1 I_49415 (I843625,I3563,I843232,I843218,);
nor I_49416 (I843656,I843258,I843591);
DFFARX1 I_49417 (I843656,I3563,I843232,I843203,);
nor I_49418 (I843687,I843535,I843591);
not I_49419 (I843704,I843687);
nand I_49420 (I843212,I843704,I843560);
not I_49421 (I843759,I3570);
DFFARX1 I_49422 (I750315,I3563,I843759,I843785,);
not I_49423 (I843793,I843785);
nand I_49424 (I843810,I750318,I750315);
and I_49425 (I843827,I843810,I750327);
DFFARX1 I_49426 (I843827,I3563,I843759,I843853,);
DFFARX1 I_49427 (I843853,I3563,I843759,I843748,);
DFFARX1 I_49428 (I750324,I3563,I843759,I843884,);
nand I_49429 (I843892,I843884,I750330);
not I_49430 (I843909,I843892);
DFFARX1 I_49431 (I843909,I3563,I843759,I843935,);
not I_49432 (I843943,I843935);
nor I_49433 (I843751,I843793,I843943);
DFFARX1 I_49434 (I750339,I3563,I843759,I843983,);
nor I_49435 (I843742,I843983,I843853);
nor I_49436 (I843733,I843983,I843909);
nand I_49437 (I844019,I750333,I750321);
and I_49438 (I844036,I844019,I750318);
DFFARX1 I_49439 (I844036,I3563,I843759,I844062,);
not I_49440 (I844070,I844062);
nand I_49441 (I844087,I844070,I843983);
nand I_49442 (I843736,I844070,I843892);
nor I_49443 (I844118,I750336,I750321);
and I_49444 (I844135,I843983,I844118);
nor I_49445 (I844152,I844070,I844135);
DFFARX1 I_49446 (I844152,I3563,I843759,I843745,);
nor I_49447 (I844183,I843785,I844118);
DFFARX1 I_49448 (I844183,I3563,I843759,I843730,);
nor I_49449 (I844214,I844062,I844118);
not I_49450 (I844231,I844214);
nand I_49451 (I843739,I844231,I844087);
not I_49452 (I844286,I3570);
DFFARX1 I_49453 (I526907,I3563,I844286,I844312,);
not I_49454 (I844320,I844312);
nand I_49455 (I844337,I526925,I526916);
and I_49456 (I844354,I844337,I526919);
DFFARX1 I_49457 (I844354,I3563,I844286,I844380,);
DFFARX1 I_49458 (I844380,I3563,I844286,I844275,);
DFFARX1 I_49459 (I526913,I3563,I844286,I844411,);
nand I_49460 (I844419,I844411,I526904);
not I_49461 (I844436,I844419);
DFFARX1 I_49462 (I844436,I3563,I844286,I844462,);
not I_49463 (I844470,I844462);
nor I_49464 (I844278,I844320,I844470);
DFFARX1 I_49465 (I526910,I3563,I844286,I844510,);
nor I_49466 (I844269,I844510,I844380);
nor I_49467 (I844260,I844510,I844436);
nand I_49468 (I844546,I526904,I526901);
and I_49469 (I844563,I844546,I526922);
DFFARX1 I_49470 (I844563,I3563,I844286,I844589,);
not I_49471 (I844597,I844589);
nand I_49472 (I844614,I844597,I844510);
nand I_49473 (I844263,I844597,I844419);
nor I_49474 (I844645,I526901,I526901);
and I_49475 (I844662,I844510,I844645);
nor I_49476 (I844679,I844597,I844662);
DFFARX1 I_49477 (I844679,I3563,I844286,I844272,);
nor I_49478 (I844710,I844312,I844645);
DFFARX1 I_49479 (I844710,I3563,I844286,I844257,);
nor I_49480 (I844741,I844589,I844645);
not I_49481 (I844758,I844741);
nand I_49482 (I844266,I844758,I844614);
not I_49483 (I844813,I3570);
DFFARX1 I_49484 (I19766,I3563,I844813,I844839,);
not I_49485 (I844847,I844839);
nand I_49486 (I844864,I19778,I19781);
and I_49487 (I844881,I844864,I19757);
DFFARX1 I_49488 (I844881,I3563,I844813,I844907,);
DFFARX1 I_49489 (I844907,I3563,I844813,I844802,);
DFFARX1 I_49490 (I19775,I3563,I844813,I844938,);
nand I_49491 (I844946,I844938,I19763);
not I_49492 (I844963,I844946);
DFFARX1 I_49493 (I844963,I3563,I844813,I844989,);
not I_49494 (I844997,I844989);
nor I_49495 (I844805,I844847,I844997);
DFFARX1 I_49496 (I19760,I3563,I844813,I845037,);
nor I_49497 (I844796,I845037,I844907);
nor I_49498 (I844787,I845037,I844963);
nand I_49499 (I845073,I19769,I19760);
and I_49500 (I845090,I845073,I19757);
DFFARX1 I_49501 (I845090,I3563,I844813,I845116,);
not I_49502 (I845124,I845116);
nand I_49503 (I845141,I845124,I845037);
nand I_49504 (I844790,I845124,I844946);
nor I_49505 (I845172,I19772,I19760);
and I_49506 (I845189,I845037,I845172);
nor I_49507 (I845206,I845124,I845189);
DFFARX1 I_49508 (I845206,I3563,I844813,I844799,);
nor I_49509 (I845237,I844839,I845172);
DFFARX1 I_49510 (I845237,I3563,I844813,I844784,);
nor I_49511 (I845268,I845116,I845172);
not I_49512 (I845285,I845268);
nand I_49513 (I844793,I845285,I845141);
not I_49514 (I845340,I3570);
DFFARX1 I_49515 (I631262,I3563,I845340,I845366,);
not I_49516 (I845374,I845366);
nand I_49517 (I845391,I631247,I631268);
and I_49518 (I845408,I845391,I631256);
DFFARX1 I_49519 (I845408,I3563,I845340,I845434,);
DFFARX1 I_49520 (I845434,I3563,I845340,I845329,);
DFFARX1 I_49521 (I631250,I3563,I845340,I845465,);
nand I_49522 (I845473,I845465,I631259);
not I_49523 (I845490,I845473);
DFFARX1 I_49524 (I845490,I3563,I845340,I845516,);
not I_49525 (I845524,I845516);
nor I_49526 (I845332,I845374,I845524);
DFFARX1 I_49527 (I631265,I3563,I845340,I845564,);
nor I_49528 (I845323,I845564,I845434);
nor I_49529 (I845314,I845564,I845490);
nand I_49530 (I845600,I631247,I631250);
and I_49531 (I845617,I845600,I631271);
DFFARX1 I_49532 (I845617,I3563,I845340,I845643,);
not I_49533 (I845651,I845643);
nand I_49534 (I845668,I845651,I845564);
nand I_49535 (I845317,I845651,I845473);
nor I_49536 (I845699,I631253,I631250);
and I_49537 (I845716,I845564,I845699);
nor I_49538 (I845733,I845651,I845716);
DFFARX1 I_49539 (I845733,I3563,I845340,I845326,);
nor I_49540 (I845764,I845366,I845699);
DFFARX1 I_49541 (I845764,I3563,I845340,I845311,);
nor I_49542 (I845795,I845643,I845699);
not I_49543 (I845812,I845795);
nand I_49544 (I845320,I845812,I845668);
not I_49545 (I845867,I3570);
DFFARX1 I_49546 (I643978,I3563,I845867,I845893,);
not I_49547 (I845901,I845893);
nand I_49548 (I845918,I643963,I643984);
and I_49549 (I845935,I845918,I643972);
DFFARX1 I_49550 (I845935,I3563,I845867,I845961,);
DFFARX1 I_49551 (I845961,I3563,I845867,I845856,);
DFFARX1 I_49552 (I643966,I3563,I845867,I845992,);
nand I_49553 (I846000,I845992,I643975);
not I_49554 (I846017,I846000);
DFFARX1 I_49555 (I846017,I3563,I845867,I846043,);
not I_49556 (I846051,I846043);
nor I_49557 (I845859,I845901,I846051);
DFFARX1 I_49558 (I643981,I3563,I845867,I846091,);
nor I_49559 (I845850,I846091,I845961);
nor I_49560 (I845841,I846091,I846017);
nand I_49561 (I846127,I643963,I643966);
and I_49562 (I846144,I846127,I643987);
DFFARX1 I_49563 (I846144,I3563,I845867,I846170,);
not I_49564 (I846178,I846170);
nand I_49565 (I846195,I846178,I846091);
nand I_49566 (I845844,I846178,I846000);
nor I_49567 (I846226,I643969,I643966);
and I_49568 (I846243,I846091,I846226);
nor I_49569 (I846260,I846178,I846243);
DFFARX1 I_49570 (I846260,I3563,I845867,I845853,);
nor I_49571 (I846291,I845893,I846226);
DFFARX1 I_49572 (I846291,I3563,I845867,I845838,);
nor I_49573 (I846322,I846170,I846226);
not I_49574 (I846339,I846322);
nand I_49575 (I845847,I846339,I846195);
not I_49576 (I846394,I3570);
DFFARX1 I_49577 (I312251,I3563,I846394,I846420,);
not I_49578 (I846428,I846420);
nand I_49579 (I846445,I312242,I312242);
and I_49580 (I846462,I846445,I312260);
DFFARX1 I_49581 (I846462,I3563,I846394,I846488,);
DFFARX1 I_49582 (I846488,I3563,I846394,I846383,);
DFFARX1 I_49583 (I312263,I3563,I846394,I846519,);
nand I_49584 (I846527,I846519,I312245);
not I_49585 (I846544,I846527);
DFFARX1 I_49586 (I846544,I3563,I846394,I846570,);
not I_49587 (I846578,I846570);
nor I_49588 (I846386,I846428,I846578);
DFFARX1 I_49589 (I312257,I3563,I846394,I846618,);
nor I_49590 (I846377,I846618,I846488);
nor I_49591 (I846368,I846618,I846544);
nand I_49592 (I846654,I312269,I312248);
and I_49593 (I846671,I846654,I312254);
DFFARX1 I_49594 (I846671,I3563,I846394,I846697,);
not I_49595 (I846705,I846697);
nand I_49596 (I846722,I846705,I846618);
nand I_49597 (I846371,I846705,I846527);
nor I_49598 (I846753,I312266,I312248);
and I_49599 (I846770,I846618,I846753);
nor I_49600 (I846787,I846705,I846770);
DFFARX1 I_49601 (I846787,I3563,I846394,I846380,);
nor I_49602 (I846818,I846420,I846753);
DFFARX1 I_49603 (I846818,I3563,I846394,I846365,);
nor I_49604 (I846849,I846697,I846753);
not I_49605 (I846866,I846849);
nand I_49606 (I846374,I846866,I846722);
not I_49607 (I846921,I3570);
DFFARX1 I_49608 (I1217017,I3563,I846921,I846947,);
not I_49609 (I846955,I846947);
nand I_49610 (I846972,I1216999,I1216999);
and I_49611 (I846989,I846972,I1217005);
DFFARX1 I_49612 (I846989,I3563,I846921,I847015,);
DFFARX1 I_49613 (I847015,I3563,I846921,I846910,);
DFFARX1 I_49614 (I1217002,I3563,I846921,I847046,);
nand I_49615 (I847054,I847046,I1217011);
not I_49616 (I847071,I847054);
DFFARX1 I_49617 (I847071,I3563,I846921,I847097,);
not I_49618 (I847105,I847097);
nor I_49619 (I846913,I846955,I847105);
DFFARX1 I_49620 (I1217023,I3563,I846921,I847145,);
nor I_49621 (I846904,I847145,I847015);
nor I_49622 (I846895,I847145,I847071);
nand I_49623 (I847181,I1217014,I1217008);
and I_49624 (I847198,I847181,I1217002);
DFFARX1 I_49625 (I847198,I3563,I846921,I847224,);
not I_49626 (I847232,I847224);
nand I_49627 (I847249,I847232,I847145);
nand I_49628 (I846898,I847232,I847054);
nor I_49629 (I847280,I1217020,I1217008);
and I_49630 (I847297,I847145,I847280);
nor I_49631 (I847314,I847232,I847297);
DFFARX1 I_49632 (I847314,I3563,I846921,I846907,);
nor I_49633 (I847345,I846947,I847280);
DFFARX1 I_49634 (I847345,I3563,I846921,I846892,);
nor I_49635 (I847376,I847224,I847280);
not I_49636 (I847393,I847376);
nand I_49637 (I846901,I847393,I847249);
not I_49638 (I847448,I3570);
DFFARX1 I_49639 (I549517,I3563,I847448,I847474,);
not I_49640 (I847482,I847474);
nand I_49641 (I847499,I549535,I549526);
and I_49642 (I847516,I847499,I549529);
DFFARX1 I_49643 (I847516,I3563,I847448,I847542,);
DFFARX1 I_49644 (I847542,I3563,I847448,I847437,);
DFFARX1 I_49645 (I549523,I3563,I847448,I847573,);
nand I_49646 (I847581,I847573,I549514);
not I_49647 (I847598,I847581);
DFFARX1 I_49648 (I847598,I3563,I847448,I847624,);
not I_49649 (I847632,I847624);
nor I_49650 (I847440,I847482,I847632);
DFFARX1 I_49651 (I549520,I3563,I847448,I847672,);
nor I_49652 (I847431,I847672,I847542);
nor I_49653 (I847422,I847672,I847598);
nand I_49654 (I847708,I549514,I549511);
and I_49655 (I847725,I847708,I549532);
DFFARX1 I_49656 (I847725,I3563,I847448,I847751,);
not I_49657 (I847759,I847751);
nand I_49658 (I847776,I847759,I847672);
nand I_49659 (I847425,I847759,I847581);
nor I_49660 (I847807,I549511,I549511);
and I_49661 (I847824,I847672,I847807);
nor I_49662 (I847841,I847759,I847824);
DFFARX1 I_49663 (I847841,I3563,I847448,I847434,);
nor I_49664 (I847872,I847474,I847807);
DFFARX1 I_49665 (I847872,I3563,I847448,I847419,);
nor I_49666 (I847903,I847751,I847807);
not I_49667 (I847920,I847903);
nand I_49668 (I847428,I847920,I847776);
not I_49669 (I847975,I3570);
DFFARX1 I_49670 (I544162,I3563,I847975,I848001,);
not I_49671 (I848009,I848001);
nand I_49672 (I848026,I544180,I544171);
and I_49673 (I848043,I848026,I544174);
DFFARX1 I_49674 (I848043,I3563,I847975,I848069,);
DFFARX1 I_49675 (I848069,I3563,I847975,I847964,);
DFFARX1 I_49676 (I544168,I3563,I847975,I848100,);
nand I_49677 (I848108,I848100,I544159);
not I_49678 (I848125,I848108);
DFFARX1 I_49679 (I848125,I3563,I847975,I848151,);
not I_49680 (I848159,I848151);
nor I_49681 (I847967,I848009,I848159);
DFFARX1 I_49682 (I544165,I3563,I847975,I848199,);
nor I_49683 (I847958,I848199,I848069);
nor I_49684 (I847949,I848199,I848125);
nand I_49685 (I848235,I544159,I544156);
and I_49686 (I848252,I848235,I544177);
DFFARX1 I_49687 (I848252,I3563,I847975,I848278,);
not I_49688 (I848286,I848278);
nand I_49689 (I848303,I848286,I848199);
nand I_49690 (I847952,I848286,I848108);
nor I_49691 (I848334,I544156,I544156);
and I_49692 (I848351,I848199,I848334);
nor I_49693 (I848368,I848286,I848351);
DFFARX1 I_49694 (I848368,I3563,I847975,I847961,);
nor I_49695 (I848399,I848001,I848334);
DFFARX1 I_49696 (I848399,I3563,I847975,I847946,);
nor I_49697 (I848430,I848278,I848334);
not I_49698 (I848447,I848430);
nand I_49699 (I847955,I848447,I848303);
not I_49700 (I848502,I3570);
DFFARX1 I_49701 (I976248,I3563,I848502,I848528,);
not I_49702 (I848536,I848528);
nand I_49703 (I848553,I976263,I976245);
and I_49704 (I848570,I848553,I976245);
DFFARX1 I_49705 (I848570,I3563,I848502,I848596,);
DFFARX1 I_49706 (I848596,I3563,I848502,I848491,);
DFFARX1 I_49707 (I976254,I3563,I848502,I848627,);
nand I_49708 (I848635,I848627,I976272);
not I_49709 (I848652,I848635);
DFFARX1 I_49710 (I848652,I3563,I848502,I848678,);
not I_49711 (I848686,I848678);
nor I_49712 (I848494,I848536,I848686);
DFFARX1 I_49713 (I976269,I3563,I848502,I848726,);
nor I_49714 (I848485,I848726,I848596);
nor I_49715 (I848476,I848726,I848652);
nand I_49716 (I848762,I976266,I976257);
and I_49717 (I848779,I848762,I976251);
DFFARX1 I_49718 (I848779,I3563,I848502,I848805,);
not I_49719 (I848813,I848805);
nand I_49720 (I848830,I848813,I848726);
nand I_49721 (I848479,I848813,I848635);
nor I_49722 (I848861,I976260,I976257);
and I_49723 (I848878,I848726,I848861);
nor I_49724 (I848895,I848813,I848878);
DFFARX1 I_49725 (I848895,I3563,I848502,I848488,);
nor I_49726 (I848926,I848528,I848861);
DFFARX1 I_49727 (I848926,I3563,I848502,I848473,);
nor I_49728 (I848957,I848805,I848861);
not I_49729 (I848974,I848957);
nand I_49730 (I848482,I848974,I848830);
not I_49731 (I849029,I3570);
DFFARX1 I_49732 (I363370,I3563,I849029,I849055,);
not I_49733 (I849063,I849055);
nand I_49734 (I849080,I363361,I363361);
and I_49735 (I849097,I849080,I363379);
DFFARX1 I_49736 (I849097,I3563,I849029,I849123,);
DFFARX1 I_49737 (I849123,I3563,I849029,I849018,);
DFFARX1 I_49738 (I363382,I3563,I849029,I849154,);
nand I_49739 (I849162,I849154,I363364);
not I_49740 (I849179,I849162);
DFFARX1 I_49741 (I849179,I3563,I849029,I849205,);
not I_49742 (I849213,I849205);
nor I_49743 (I849021,I849063,I849213);
DFFARX1 I_49744 (I363376,I3563,I849029,I849253,);
nor I_49745 (I849012,I849253,I849123);
nor I_49746 (I849003,I849253,I849179);
nand I_49747 (I849289,I363388,I363367);
and I_49748 (I849306,I849289,I363373);
DFFARX1 I_49749 (I849306,I3563,I849029,I849332,);
not I_49750 (I849340,I849332);
nand I_49751 (I849357,I849340,I849253);
nand I_49752 (I849006,I849340,I849162);
nor I_49753 (I849388,I363385,I363367);
and I_49754 (I849405,I849253,I849388);
nor I_49755 (I849422,I849340,I849405);
DFFARX1 I_49756 (I849422,I3563,I849029,I849015,);
nor I_49757 (I849453,I849055,I849388);
DFFARX1 I_49758 (I849453,I3563,I849029,I849000,);
nor I_49759 (I849484,I849332,I849388);
not I_49760 (I849501,I849484);
nand I_49761 (I849009,I849501,I849357);
not I_49762 (I849556,I3570);
DFFARX1 I_49763 (I458856,I3563,I849556,I849582,);
not I_49764 (I849590,I849582);
nand I_49765 (I849607,I458853,I458862);
and I_49766 (I849624,I849607,I458871);
DFFARX1 I_49767 (I849624,I3563,I849556,I849650,);
DFFARX1 I_49768 (I849650,I3563,I849556,I849545,);
DFFARX1 I_49769 (I458874,I3563,I849556,I849681,);
nand I_49770 (I849689,I849681,I458877);
not I_49771 (I849706,I849689);
DFFARX1 I_49772 (I849706,I3563,I849556,I849732,);
not I_49773 (I849740,I849732);
nor I_49774 (I849548,I849590,I849740);
DFFARX1 I_49775 (I458850,I3563,I849556,I849780,);
nor I_49776 (I849539,I849780,I849650);
nor I_49777 (I849530,I849780,I849706);
nand I_49778 (I849816,I458865,I458868);
and I_49779 (I849833,I849816,I458859);
DFFARX1 I_49780 (I849833,I3563,I849556,I849859,);
not I_49781 (I849867,I849859);
nand I_49782 (I849884,I849867,I849780);
nand I_49783 (I849533,I849867,I849689);
nor I_49784 (I849915,I458850,I458868);
and I_49785 (I849932,I849780,I849915);
nor I_49786 (I849949,I849867,I849932);
DFFARX1 I_49787 (I849949,I3563,I849556,I849542,);
nor I_49788 (I849980,I849582,I849915);
DFFARX1 I_49789 (I849980,I3563,I849556,I849527,);
nor I_49790 (I850011,I849859,I849915);
not I_49791 (I850028,I850011);
nand I_49792 (I849536,I850028,I849884);
not I_49793 (I850083,I3570);
DFFARX1 I_49794 (I1303377,I3563,I850083,I850109,);
not I_49795 (I850117,I850109);
nand I_49796 (I850134,I1303359,I1303362);
and I_49797 (I850151,I850134,I1303374);
DFFARX1 I_49798 (I850151,I3563,I850083,I850177,);
DFFARX1 I_49799 (I850177,I3563,I850083,I850072,);
DFFARX1 I_49800 (I1303383,I3563,I850083,I850208,);
nand I_49801 (I850216,I850208,I1303368);
not I_49802 (I850233,I850216);
DFFARX1 I_49803 (I850233,I3563,I850083,I850259,);
not I_49804 (I850267,I850259);
nor I_49805 (I850075,I850117,I850267);
DFFARX1 I_49806 (I1303380,I3563,I850083,I850307,);
nor I_49807 (I850066,I850307,I850177);
nor I_49808 (I850057,I850307,I850233);
nand I_49809 (I850343,I1303371,I1303365);
and I_49810 (I850360,I850343,I1303359);
DFFARX1 I_49811 (I850360,I3563,I850083,I850386,);
not I_49812 (I850394,I850386);
nand I_49813 (I850411,I850394,I850307);
nand I_49814 (I850060,I850394,I850216);
nor I_49815 (I850442,I1303362,I1303365);
and I_49816 (I850459,I850307,I850442);
nor I_49817 (I850476,I850394,I850459);
DFFARX1 I_49818 (I850476,I3563,I850083,I850069,);
nor I_49819 (I850507,I850109,I850442);
DFFARX1 I_49820 (I850507,I3563,I850083,I850054,);
nor I_49821 (I850538,I850386,I850442);
not I_49822 (I850555,I850538);
nand I_49823 (I850063,I850555,I850411);
not I_49824 (I850610,I3570);
DFFARX1 I_49825 (I1314937,I3563,I850610,I850636,);
not I_49826 (I850644,I850636);
nand I_49827 (I850661,I1314919,I1314922);
and I_49828 (I850678,I850661,I1314934);
DFFARX1 I_49829 (I850678,I3563,I850610,I850704,);
DFFARX1 I_49830 (I850704,I3563,I850610,I850599,);
DFFARX1 I_49831 (I1314943,I3563,I850610,I850735,);
nand I_49832 (I850743,I850735,I1314928);
not I_49833 (I850760,I850743);
DFFARX1 I_49834 (I850760,I3563,I850610,I850786,);
not I_49835 (I850794,I850786);
nor I_49836 (I850602,I850644,I850794);
DFFARX1 I_49837 (I1314940,I3563,I850610,I850834,);
nor I_49838 (I850593,I850834,I850704);
nor I_49839 (I850584,I850834,I850760);
nand I_49840 (I850870,I1314931,I1314925);
and I_49841 (I850887,I850870,I1314919);
DFFARX1 I_49842 (I850887,I3563,I850610,I850913,);
not I_49843 (I850921,I850913);
nand I_49844 (I850938,I850921,I850834);
nand I_49845 (I850587,I850921,I850743);
nor I_49846 (I850969,I1314922,I1314925);
and I_49847 (I850986,I850834,I850969);
nor I_49848 (I851003,I850921,I850986);
DFFARX1 I_49849 (I851003,I3563,I850610,I850596,);
nor I_49850 (I851034,I850636,I850969);
DFFARX1 I_49851 (I851034,I3563,I850610,I850581,);
nor I_49852 (I851065,I850913,I850969);
not I_49853 (I851082,I851065);
nand I_49854 (I850590,I851082,I850938);
not I_49855 (I851137,I3570);
DFFARX1 I_49856 (I7753,I3563,I851137,I851163,);
not I_49857 (I851171,I851163);
nand I_49858 (I851188,I7759,I7741);
and I_49859 (I851205,I851188,I7750);
DFFARX1 I_49860 (I851205,I3563,I851137,I851231,);
DFFARX1 I_49861 (I851231,I3563,I851137,I851126,);
DFFARX1 I_49862 (I7741,I3563,I851137,I851262,);
nand I_49863 (I851270,I851262,I7744);
not I_49864 (I851287,I851270);
DFFARX1 I_49865 (I851287,I3563,I851137,I851313,);
not I_49866 (I851321,I851313);
nor I_49867 (I851129,I851171,I851321);
DFFARX1 I_49868 (I7744,I3563,I851137,I851361,);
nor I_49869 (I851120,I851361,I851231);
nor I_49870 (I851111,I851361,I851287);
nand I_49871 (I851397,I7747,I7756);
and I_49872 (I851414,I851397,I7738);
DFFARX1 I_49873 (I851414,I3563,I851137,I851440,);
not I_49874 (I851448,I851440);
nand I_49875 (I851465,I851448,I851361);
nand I_49876 (I851114,I851448,I851270);
nor I_49877 (I851496,I7738,I7756);
and I_49878 (I851513,I851361,I851496);
nor I_49879 (I851530,I851448,I851513);
DFFARX1 I_49880 (I851530,I3563,I851137,I851123,);
nor I_49881 (I851561,I851163,I851496);
DFFARX1 I_49882 (I851561,I3563,I851137,I851108,);
nor I_49883 (I851592,I851440,I851496);
not I_49884 (I851609,I851592);
nand I_49885 (I851117,I851609,I851465);
not I_49886 (I851664,I3570);
DFFARX1 I_49887 (I1222797,I3563,I851664,I851690,);
not I_49888 (I851698,I851690);
nand I_49889 (I851715,I1222779,I1222779);
and I_49890 (I851732,I851715,I1222785);
DFFARX1 I_49891 (I851732,I3563,I851664,I851758,);
DFFARX1 I_49892 (I851758,I3563,I851664,I851653,);
DFFARX1 I_49893 (I1222782,I3563,I851664,I851789,);
nand I_49894 (I851797,I851789,I1222791);
not I_49895 (I851814,I851797);
DFFARX1 I_49896 (I851814,I3563,I851664,I851840,);
not I_49897 (I851848,I851840);
nor I_49898 (I851656,I851698,I851848);
DFFARX1 I_49899 (I1222803,I3563,I851664,I851888,);
nor I_49900 (I851647,I851888,I851758);
nor I_49901 (I851638,I851888,I851814);
nand I_49902 (I851924,I1222794,I1222788);
and I_49903 (I851941,I851924,I1222782);
DFFARX1 I_49904 (I851941,I3563,I851664,I851967,);
not I_49905 (I851975,I851967);
nand I_49906 (I851992,I851975,I851888);
nand I_49907 (I851641,I851975,I851797);
nor I_49908 (I852023,I1222800,I1222788);
and I_49909 (I852040,I851888,I852023);
nor I_49910 (I852057,I851975,I852040);
DFFARX1 I_49911 (I852057,I3563,I851664,I851650,);
nor I_49912 (I852088,I851690,I852023);
DFFARX1 I_49913 (I852088,I3563,I851664,I851635,);
nor I_49914 (I852119,I851967,I852023);
not I_49915 (I852136,I852119);
nand I_49916 (I851644,I852136,I851992);
not I_49917 (I852191,I3570);
DFFARX1 I_49918 (I129397,I3563,I852191,I852217,);
not I_49919 (I852225,I852217);
nand I_49920 (I852242,I129373,I129382);
and I_49921 (I852259,I852242,I129376);
DFFARX1 I_49922 (I852259,I3563,I852191,I852285,);
DFFARX1 I_49923 (I852285,I3563,I852191,I852180,);
DFFARX1 I_49924 (I129394,I3563,I852191,I852316,);
nand I_49925 (I852324,I852316,I129385);
not I_49926 (I852341,I852324);
DFFARX1 I_49927 (I852341,I3563,I852191,I852367,);
not I_49928 (I852375,I852367);
nor I_49929 (I852183,I852225,I852375);
DFFARX1 I_49930 (I129379,I3563,I852191,I852415,);
nor I_49931 (I852174,I852415,I852285);
nor I_49932 (I852165,I852415,I852341);
nand I_49933 (I852451,I129391,I129388);
and I_49934 (I852468,I852451,I129376);
DFFARX1 I_49935 (I852468,I3563,I852191,I852494,);
not I_49936 (I852502,I852494);
nand I_49937 (I852519,I852502,I852415);
nand I_49938 (I852168,I852502,I852324);
nor I_49939 (I852550,I129373,I129388);
and I_49940 (I852567,I852415,I852550);
nor I_49941 (I852584,I852502,I852567);
DFFARX1 I_49942 (I852584,I3563,I852191,I852177,);
nor I_49943 (I852615,I852217,I852550);
DFFARX1 I_49944 (I852615,I3563,I852191,I852162,);
nor I_49945 (I852646,I852494,I852550);
not I_49946 (I852663,I852646);
nand I_49947 (I852171,I852663,I852519);
not I_49948 (I852718,I3570);
DFFARX1 I_49949 (I1148235,I3563,I852718,I852744,);
not I_49950 (I852752,I852744);
nand I_49951 (I852769,I1148217,I1148217);
and I_49952 (I852786,I852769,I1148223);
DFFARX1 I_49953 (I852786,I3563,I852718,I852812,);
DFFARX1 I_49954 (I852812,I3563,I852718,I852707,);
DFFARX1 I_49955 (I1148220,I3563,I852718,I852843,);
nand I_49956 (I852851,I852843,I1148229);
not I_49957 (I852868,I852851);
DFFARX1 I_49958 (I852868,I3563,I852718,I852894,);
not I_49959 (I852902,I852894);
nor I_49960 (I852710,I852752,I852902);
DFFARX1 I_49961 (I1148241,I3563,I852718,I852942,);
nor I_49962 (I852701,I852942,I852812);
nor I_49963 (I852692,I852942,I852868);
nand I_49964 (I852978,I1148232,I1148226);
and I_49965 (I852995,I852978,I1148220);
DFFARX1 I_49966 (I852995,I3563,I852718,I853021,);
not I_49967 (I853029,I853021);
nand I_49968 (I853046,I853029,I852942);
nand I_49969 (I852695,I853029,I852851);
nor I_49970 (I853077,I1148238,I1148226);
and I_49971 (I853094,I852942,I853077);
nor I_49972 (I853111,I853029,I853094);
DFFARX1 I_49973 (I853111,I3563,I852718,I852704,);
nor I_49974 (I853142,I852744,I853077);
DFFARX1 I_49975 (I853142,I3563,I852718,I852689,);
nor I_49976 (I853173,I853021,I853077);
not I_49977 (I853190,I853173);
nand I_49978 (I852698,I853190,I853046);
not I_49979 (I853245,I3570);
DFFARX1 I_49980 (I802913,I3563,I853245,I853271,);
not I_49981 (I853279,I853271);
nand I_49982 (I853296,I802916,I802913);
and I_49983 (I853313,I853296,I802925);
DFFARX1 I_49984 (I853313,I3563,I853245,I853339,);
DFFARX1 I_49985 (I853339,I3563,I853245,I853234,);
DFFARX1 I_49986 (I802922,I3563,I853245,I853370,);
nand I_49987 (I853378,I853370,I802928);
not I_49988 (I853395,I853378);
DFFARX1 I_49989 (I853395,I3563,I853245,I853421,);
not I_49990 (I853429,I853421);
nor I_49991 (I853237,I853279,I853429);
DFFARX1 I_49992 (I802937,I3563,I853245,I853469,);
nor I_49993 (I853228,I853469,I853339);
nor I_49994 (I853219,I853469,I853395);
nand I_49995 (I853505,I802931,I802919);
and I_49996 (I853522,I853505,I802916);
DFFARX1 I_49997 (I853522,I3563,I853245,I853548,);
not I_49998 (I853556,I853548);
nand I_49999 (I853573,I853556,I853469);
nand I_50000 (I853222,I853556,I853378);
nor I_50001 (I853604,I802934,I802919);
and I_50002 (I853621,I853469,I853604);
nor I_50003 (I853638,I853556,I853621);
DFFARX1 I_50004 (I853638,I3563,I853245,I853231,);
nor I_50005 (I853669,I853271,I853604);
DFFARX1 I_50006 (I853669,I3563,I853245,I853216,);
nor I_50007 (I853700,I853548,I853604);
not I_50008 (I853717,I853700);
nand I_50009 (I853225,I853717,I853573);
not I_50010 (I853772,I3570);
DFFARX1 I_50011 (I338074,I3563,I853772,I853798,);
not I_50012 (I853806,I853798);
nand I_50013 (I853823,I338065,I338065);
and I_50014 (I853840,I853823,I338083);
DFFARX1 I_50015 (I853840,I3563,I853772,I853866,);
DFFARX1 I_50016 (I853866,I3563,I853772,I853761,);
DFFARX1 I_50017 (I338086,I3563,I853772,I853897,);
nand I_50018 (I853905,I853897,I338068);
not I_50019 (I853922,I853905);
DFFARX1 I_50020 (I853922,I3563,I853772,I853948,);
not I_50021 (I853956,I853948);
nor I_50022 (I853764,I853806,I853956);
DFFARX1 I_50023 (I338080,I3563,I853772,I853996,);
nor I_50024 (I853755,I853996,I853866);
nor I_50025 (I853746,I853996,I853922);
nand I_50026 (I854032,I338092,I338071);
and I_50027 (I854049,I854032,I338077);
DFFARX1 I_50028 (I854049,I3563,I853772,I854075,);
not I_50029 (I854083,I854075);
nand I_50030 (I854100,I854083,I853996);
nand I_50031 (I853749,I854083,I853905);
nor I_50032 (I854131,I338089,I338071);
and I_50033 (I854148,I853996,I854131);
nor I_50034 (I854165,I854083,I854148);
DFFARX1 I_50035 (I854165,I3563,I853772,I853758,);
nor I_50036 (I854196,I853798,I854131);
DFFARX1 I_50037 (I854196,I3563,I853772,I853743,);
nor I_50038 (I854227,I854075,I854131);
not I_50039 (I854244,I854227);
nand I_50040 (I853752,I854244,I854100);
not I_50041 (I854299,I3570);
DFFARX1 I_50042 (I1399373,I3563,I854299,I854325,);
not I_50043 (I854333,I854325);
nand I_50044 (I854350,I1399370,I1399379);
and I_50045 (I854367,I854350,I1399358);
DFFARX1 I_50046 (I854367,I3563,I854299,I854393,);
DFFARX1 I_50047 (I854393,I3563,I854299,I854288,);
DFFARX1 I_50048 (I1399361,I3563,I854299,I854424,);
nand I_50049 (I854432,I854424,I1399376);
not I_50050 (I854449,I854432);
DFFARX1 I_50051 (I854449,I3563,I854299,I854475,);
not I_50052 (I854483,I854475);
nor I_50053 (I854291,I854333,I854483);
DFFARX1 I_50054 (I1399382,I3563,I854299,I854523,);
nor I_50055 (I854282,I854523,I854393);
nor I_50056 (I854273,I854523,I854449);
nand I_50057 (I854559,I1399364,I1399385);
and I_50058 (I854576,I854559,I1399367);
DFFARX1 I_50059 (I854576,I3563,I854299,I854602,);
not I_50060 (I854610,I854602);
nand I_50061 (I854627,I854610,I854523);
nand I_50062 (I854276,I854610,I854432);
nor I_50063 (I854658,I1399358,I1399385);
and I_50064 (I854675,I854523,I854658);
nor I_50065 (I854692,I854610,I854675);
DFFARX1 I_50066 (I854692,I3563,I854299,I854285,);
nor I_50067 (I854723,I854325,I854658);
DFFARX1 I_50068 (I854723,I3563,I854299,I854270,);
nor I_50069 (I854754,I854602,I854658);
not I_50070 (I854771,I854754);
nand I_50071 (I854279,I854771,I854627);
not I_50072 (I854826,I3570);
DFFARX1 I_50073 (I237499,I3563,I854826,I854852,);
not I_50074 (I854860,I854852);
nand I_50075 (I854877,I237496,I237514);
and I_50076 (I854894,I854877,I237505);
DFFARX1 I_50077 (I854894,I3563,I854826,I854920,);
DFFARX1 I_50078 (I854920,I3563,I854826,I854815,);
DFFARX1 I_50079 (I237511,I3563,I854826,I854951,);
nand I_50080 (I854959,I854951,I237508);
not I_50081 (I854976,I854959);
DFFARX1 I_50082 (I854976,I3563,I854826,I855002,);
not I_50083 (I855010,I855002);
nor I_50084 (I854818,I854860,I855010);
DFFARX1 I_50085 (I237502,I3563,I854826,I855050,);
nor I_50086 (I854809,I855050,I854920);
nor I_50087 (I854800,I855050,I854976);
nand I_50088 (I855086,I237493,I237517);
and I_50089 (I855103,I855086,I237496);
DFFARX1 I_50090 (I855103,I3563,I854826,I855129,);
not I_50091 (I855137,I855129);
nand I_50092 (I855154,I855137,I855050);
nand I_50093 (I854803,I855137,I854959);
nor I_50094 (I855185,I237493,I237517);
and I_50095 (I855202,I855050,I855185);
nor I_50096 (I855219,I855137,I855202);
DFFARX1 I_50097 (I855219,I3563,I854826,I854812,);
nor I_50098 (I855250,I854852,I855185);
DFFARX1 I_50099 (I855250,I3563,I854826,I854797,);
nor I_50100 (I855281,I855129,I855185);
not I_50101 (I855298,I855281);
nand I_50102 (I854806,I855298,I855154);
not I_50103 (I855353,I3570);
DFFARX1 I_50104 (I1024052,I3563,I855353,I855379,);
not I_50105 (I855387,I855379);
nand I_50106 (I855404,I1024067,I1024049);
and I_50107 (I855421,I855404,I1024049);
DFFARX1 I_50108 (I855421,I3563,I855353,I855447,);
DFFARX1 I_50109 (I855447,I3563,I855353,I855342,);
DFFARX1 I_50110 (I1024058,I3563,I855353,I855478,);
nand I_50111 (I855486,I855478,I1024076);
not I_50112 (I855503,I855486);
DFFARX1 I_50113 (I855503,I3563,I855353,I855529,);
not I_50114 (I855537,I855529);
nor I_50115 (I855345,I855387,I855537);
DFFARX1 I_50116 (I1024073,I3563,I855353,I855577,);
nor I_50117 (I855336,I855577,I855447);
nor I_50118 (I855327,I855577,I855503);
nand I_50119 (I855613,I1024070,I1024061);
and I_50120 (I855630,I855613,I1024055);
DFFARX1 I_50121 (I855630,I3563,I855353,I855656,);
not I_50122 (I855664,I855656);
nand I_50123 (I855681,I855664,I855577);
nand I_50124 (I855330,I855664,I855486);
nor I_50125 (I855712,I1024064,I1024061);
and I_50126 (I855729,I855577,I855712);
nor I_50127 (I855746,I855664,I855729);
DFFARX1 I_50128 (I855746,I3563,I855353,I855339,);
nor I_50129 (I855777,I855379,I855712);
DFFARX1 I_50130 (I855777,I3563,I855353,I855324,);
nor I_50131 (I855808,I855656,I855712);
not I_50132 (I855825,I855808);
nand I_50133 (I855333,I855825,I855681);
not I_50134 (I855880,I3570);
DFFARX1 I_50135 (I219054,I3563,I855880,I855906,);
not I_50136 (I855914,I855906);
nand I_50137 (I855931,I219051,I219069);
and I_50138 (I855948,I855931,I219060);
DFFARX1 I_50139 (I855948,I3563,I855880,I855974,);
DFFARX1 I_50140 (I855974,I3563,I855880,I855869,);
DFFARX1 I_50141 (I219066,I3563,I855880,I856005,);
nand I_50142 (I856013,I856005,I219063);
not I_50143 (I856030,I856013);
DFFARX1 I_50144 (I856030,I3563,I855880,I856056,);
not I_50145 (I856064,I856056);
nor I_50146 (I855872,I855914,I856064);
DFFARX1 I_50147 (I219057,I3563,I855880,I856104,);
nor I_50148 (I855863,I856104,I855974);
nor I_50149 (I855854,I856104,I856030);
nand I_50150 (I856140,I219048,I219072);
and I_50151 (I856157,I856140,I219051);
DFFARX1 I_50152 (I856157,I3563,I855880,I856183,);
not I_50153 (I856191,I856183);
nand I_50154 (I856208,I856191,I856104);
nand I_50155 (I855857,I856191,I856013);
nor I_50156 (I856239,I219048,I219072);
and I_50157 (I856256,I856104,I856239);
nor I_50158 (I856273,I856191,I856256);
DFFARX1 I_50159 (I856273,I3563,I855880,I855866,);
nor I_50160 (I856304,I855906,I856239);
DFFARX1 I_50161 (I856304,I3563,I855880,I855851,);
nor I_50162 (I856335,I856183,I856239);
not I_50163 (I856352,I856335);
nand I_50164 (I855860,I856352,I856208);
not I_50165 (I856407,I3570);
DFFARX1 I_50166 (I196444,I3563,I856407,I856433,);
not I_50167 (I856441,I856433);
nand I_50168 (I856458,I196441,I196459);
and I_50169 (I856475,I856458,I196450);
DFFARX1 I_50170 (I856475,I3563,I856407,I856501,);
DFFARX1 I_50171 (I856501,I3563,I856407,I856396,);
DFFARX1 I_50172 (I196456,I3563,I856407,I856532,);
nand I_50173 (I856540,I856532,I196453);
not I_50174 (I856557,I856540);
DFFARX1 I_50175 (I856557,I3563,I856407,I856583,);
not I_50176 (I856591,I856583);
nor I_50177 (I856399,I856441,I856591);
DFFARX1 I_50178 (I196447,I3563,I856407,I856631,);
nor I_50179 (I856390,I856631,I856501);
nor I_50180 (I856381,I856631,I856557);
nand I_50181 (I856667,I196438,I196462);
and I_50182 (I856684,I856667,I196441);
DFFARX1 I_50183 (I856684,I3563,I856407,I856710,);
not I_50184 (I856718,I856710);
nand I_50185 (I856735,I856718,I856631);
nand I_50186 (I856384,I856718,I856540);
nor I_50187 (I856766,I196438,I196462);
and I_50188 (I856783,I856631,I856766);
nor I_50189 (I856800,I856718,I856783);
DFFARX1 I_50190 (I856800,I3563,I856407,I856393,);
nor I_50191 (I856831,I856433,I856766);
DFFARX1 I_50192 (I856831,I3563,I856407,I856378,);
nor I_50193 (I856862,I856710,I856766);
not I_50194 (I856879,I856862);
nand I_50195 (I856387,I856879,I856735);
not I_50196 (I856934,I3570);
DFFARX1 I_50197 (I606986,I3563,I856934,I856960,);
not I_50198 (I856968,I856960);
nand I_50199 (I856985,I606971,I606992);
and I_50200 (I857002,I856985,I606980);
DFFARX1 I_50201 (I857002,I3563,I856934,I857028,);
DFFARX1 I_50202 (I857028,I3563,I856934,I856923,);
DFFARX1 I_50203 (I606974,I3563,I856934,I857059,);
nand I_50204 (I857067,I857059,I606983);
not I_50205 (I857084,I857067);
DFFARX1 I_50206 (I857084,I3563,I856934,I857110,);
not I_50207 (I857118,I857110);
nor I_50208 (I856926,I856968,I857118);
DFFARX1 I_50209 (I606989,I3563,I856934,I857158,);
nor I_50210 (I856917,I857158,I857028);
nor I_50211 (I856908,I857158,I857084);
nand I_50212 (I857194,I606971,I606974);
and I_50213 (I857211,I857194,I606995);
DFFARX1 I_50214 (I857211,I3563,I856934,I857237,);
not I_50215 (I857245,I857237);
nand I_50216 (I857262,I857245,I857158);
nand I_50217 (I856911,I857245,I857067);
nor I_50218 (I857293,I606977,I606974);
and I_50219 (I857310,I857158,I857293);
nor I_50220 (I857327,I857245,I857310);
DFFARX1 I_50221 (I857327,I3563,I856934,I856920,);
nor I_50222 (I857358,I856960,I857293);
DFFARX1 I_50223 (I857358,I3563,I856934,I856905,);
nor I_50224 (I857389,I857237,I857293);
not I_50225 (I857406,I857389);
nand I_50226 (I856914,I857406,I857262);
not I_50227 (I857461,I3570);
DFFARX1 I_50228 (I1085938,I3563,I857461,I857487,);
not I_50229 (I857495,I857487);
nand I_50230 (I857512,I1085947,I1085935);
and I_50231 (I857529,I857512,I1085932);
DFFARX1 I_50232 (I857529,I3563,I857461,I857555,);
DFFARX1 I_50233 (I857555,I3563,I857461,I857450,);
DFFARX1 I_50234 (I1085932,I3563,I857461,I857586,);
nand I_50235 (I857594,I857586,I1085929);
not I_50236 (I857611,I857594);
DFFARX1 I_50237 (I857611,I3563,I857461,I857637,);
not I_50238 (I857645,I857637);
nor I_50239 (I857453,I857495,I857645);
DFFARX1 I_50240 (I1085935,I3563,I857461,I857685,);
nor I_50241 (I857444,I857685,I857555);
nor I_50242 (I857435,I857685,I857611);
nand I_50243 (I857721,I1085950,I1085941);
and I_50244 (I857738,I857721,I1085944);
DFFARX1 I_50245 (I857738,I3563,I857461,I857764,);
not I_50246 (I857772,I857764);
nand I_50247 (I857789,I857772,I857685);
nand I_50248 (I857438,I857772,I857594);
nor I_50249 (I857820,I1085929,I1085941);
and I_50250 (I857837,I857685,I857820);
nor I_50251 (I857854,I857772,I857837);
DFFARX1 I_50252 (I857854,I3563,I857461,I857447,);
nor I_50253 (I857885,I857487,I857820);
DFFARX1 I_50254 (I857885,I3563,I857461,I857432,);
nor I_50255 (I857916,I857764,I857820);
not I_50256 (I857933,I857916);
nand I_50257 (I857441,I857933,I857789);
not I_50258 (I857988,I3570);
DFFARX1 I_50259 (I768811,I3563,I857988,I858014,);
not I_50260 (I858022,I858014);
nand I_50261 (I858039,I768814,I768811);
and I_50262 (I858056,I858039,I768823);
DFFARX1 I_50263 (I858056,I3563,I857988,I858082,);
DFFARX1 I_50264 (I858082,I3563,I857988,I857977,);
DFFARX1 I_50265 (I768820,I3563,I857988,I858113,);
nand I_50266 (I858121,I858113,I768826);
not I_50267 (I858138,I858121);
DFFARX1 I_50268 (I858138,I3563,I857988,I858164,);
not I_50269 (I858172,I858164);
nor I_50270 (I857980,I858022,I858172);
DFFARX1 I_50271 (I768835,I3563,I857988,I858212,);
nor I_50272 (I857971,I858212,I858082);
nor I_50273 (I857962,I858212,I858138);
nand I_50274 (I858248,I768829,I768817);
and I_50275 (I858265,I858248,I768814);
DFFARX1 I_50276 (I858265,I3563,I857988,I858291,);
not I_50277 (I858299,I858291);
nand I_50278 (I858316,I858299,I858212);
nand I_50279 (I857965,I858299,I858121);
nor I_50280 (I858347,I768832,I768817);
and I_50281 (I858364,I858212,I858347);
nor I_50282 (I858381,I858299,I858364);
DFFARX1 I_50283 (I858381,I3563,I857988,I857974,);
nor I_50284 (I858412,I858014,I858347);
DFFARX1 I_50285 (I858412,I3563,I857988,I857959,);
nor I_50286 (I858443,I858291,I858347);
not I_50287 (I858460,I858443);
nand I_50288 (I857968,I858460,I858316);
not I_50289 (I858515,I3570);
DFFARX1 I_50290 (I278554,I3563,I858515,I858541,);
not I_50291 (I858549,I858541);
nand I_50292 (I858566,I278551,I278569);
and I_50293 (I858583,I858566,I278560);
DFFARX1 I_50294 (I858583,I3563,I858515,I858609,);
DFFARX1 I_50295 (I858609,I3563,I858515,I858504,);
DFFARX1 I_50296 (I278566,I3563,I858515,I858640,);
nand I_50297 (I858648,I858640,I278563);
not I_50298 (I858665,I858648);
DFFARX1 I_50299 (I858665,I3563,I858515,I858691,);
not I_50300 (I858699,I858691);
nor I_50301 (I858507,I858549,I858699);
DFFARX1 I_50302 (I278557,I3563,I858515,I858739,);
nor I_50303 (I858498,I858739,I858609);
nor I_50304 (I858489,I858739,I858665);
nand I_50305 (I858775,I278548,I278572);
and I_50306 (I858792,I858775,I278551);
DFFARX1 I_50307 (I858792,I3563,I858515,I858818,);
not I_50308 (I858826,I858818);
nand I_50309 (I858843,I858826,I858739);
nand I_50310 (I858492,I858826,I858648);
nor I_50311 (I858874,I278548,I278572);
and I_50312 (I858891,I858739,I858874);
nor I_50313 (I858908,I858826,I858891);
DFFARX1 I_50314 (I858908,I3563,I858515,I858501,);
nor I_50315 (I858939,I858541,I858874);
DFFARX1 I_50316 (I858939,I3563,I858515,I858486,);
nor I_50317 (I858970,I858818,I858874);
not I_50318 (I858987,I858970);
nand I_50319 (I858495,I858987,I858843);
not I_50320 (I859042,I3570);
DFFARX1 I_50321 (I919400,I3563,I859042,I859068,);
not I_50322 (I859076,I859068);
nand I_50323 (I859093,I919415,I919397);
and I_50324 (I859110,I859093,I919397);
DFFARX1 I_50325 (I859110,I3563,I859042,I859136,);
DFFARX1 I_50326 (I859136,I3563,I859042,I859031,);
DFFARX1 I_50327 (I919406,I3563,I859042,I859167,);
nand I_50328 (I859175,I859167,I919424);
not I_50329 (I859192,I859175);
DFFARX1 I_50330 (I859192,I3563,I859042,I859218,);
not I_50331 (I859226,I859218);
nor I_50332 (I859034,I859076,I859226);
DFFARX1 I_50333 (I919421,I3563,I859042,I859266,);
nor I_50334 (I859025,I859266,I859136);
nor I_50335 (I859016,I859266,I859192);
nand I_50336 (I859302,I919418,I919409);
and I_50337 (I859319,I859302,I919403);
DFFARX1 I_50338 (I859319,I3563,I859042,I859345,);
not I_50339 (I859353,I859345);
nand I_50340 (I859370,I859353,I859266);
nand I_50341 (I859019,I859353,I859175);
nor I_50342 (I859401,I919412,I919409);
and I_50343 (I859418,I859266,I859401);
nor I_50344 (I859435,I859353,I859418);
DFFARX1 I_50345 (I859435,I3563,I859042,I859028,);
nor I_50346 (I859466,I859068,I859401);
DFFARX1 I_50347 (I859466,I3563,I859042,I859013,);
nor I_50348 (I859497,I859345,I859401);
not I_50349 (I859514,I859497);
nand I_50350 (I859022,I859514,I859370);
not I_50351 (I859569,I3570);
DFFARX1 I_50352 (I1104885,I3563,I859569,I859595,);
not I_50353 (I859603,I859595);
nand I_50354 (I859620,I1104867,I1104867);
and I_50355 (I859637,I859620,I1104873);
DFFARX1 I_50356 (I859637,I3563,I859569,I859663,);
DFFARX1 I_50357 (I859663,I3563,I859569,I859558,);
DFFARX1 I_50358 (I1104870,I3563,I859569,I859694,);
nand I_50359 (I859702,I859694,I1104879);
not I_50360 (I859719,I859702);
DFFARX1 I_50361 (I859719,I3563,I859569,I859745,);
not I_50362 (I859753,I859745);
nor I_50363 (I859561,I859603,I859753);
DFFARX1 I_50364 (I1104891,I3563,I859569,I859793,);
nor I_50365 (I859552,I859793,I859663);
nor I_50366 (I859543,I859793,I859719);
nand I_50367 (I859829,I1104882,I1104876);
and I_50368 (I859846,I859829,I1104870);
DFFARX1 I_50369 (I859846,I3563,I859569,I859872,);
not I_50370 (I859880,I859872);
nand I_50371 (I859897,I859880,I859793);
nand I_50372 (I859546,I859880,I859702);
nor I_50373 (I859928,I1104888,I1104876);
and I_50374 (I859945,I859793,I859928);
nor I_50375 (I859962,I859880,I859945);
DFFARX1 I_50376 (I859962,I3563,I859569,I859555,);
nor I_50377 (I859993,I859595,I859928);
DFFARX1 I_50378 (I859993,I3563,I859569,I859540,);
nor I_50379 (I860024,I859872,I859928);
not I_50380 (I860041,I860024);
nand I_50381 (I859549,I860041,I859897);
not I_50382 (I860096,I3570);
DFFARX1 I_50383 (I96723,I3563,I860096,I860122,);
not I_50384 (I860130,I860122);
nand I_50385 (I860147,I96699,I96708);
and I_50386 (I860164,I860147,I96702);
DFFARX1 I_50387 (I860164,I3563,I860096,I860190,);
DFFARX1 I_50388 (I860190,I3563,I860096,I860085,);
DFFARX1 I_50389 (I96720,I3563,I860096,I860221,);
nand I_50390 (I860229,I860221,I96711);
not I_50391 (I860246,I860229);
DFFARX1 I_50392 (I860246,I3563,I860096,I860272,);
not I_50393 (I860280,I860272);
nor I_50394 (I860088,I860130,I860280);
DFFARX1 I_50395 (I96705,I3563,I860096,I860320,);
nor I_50396 (I860079,I860320,I860190);
nor I_50397 (I860070,I860320,I860246);
nand I_50398 (I860356,I96717,I96714);
and I_50399 (I860373,I860356,I96702);
DFFARX1 I_50400 (I860373,I3563,I860096,I860399,);
not I_50401 (I860407,I860399);
nand I_50402 (I860424,I860407,I860320);
nand I_50403 (I860073,I860407,I860229);
nor I_50404 (I860455,I96699,I96714);
and I_50405 (I860472,I860320,I860455);
nor I_50406 (I860489,I860407,I860472);
DFFARX1 I_50407 (I860489,I3563,I860096,I860082,);
nor I_50408 (I860520,I860122,I860455);
DFFARX1 I_50409 (I860520,I3563,I860096,I860067,);
nor I_50410 (I860551,I860399,I860455);
not I_50411 (I860568,I860551);
nand I_50412 (I860076,I860568,I860424);
not I_50413 (I860623,I3570);
DFFARX1 I_50414 (I286289,I3563,I860623,I860649,);
not I_50415 (I860657,I860649);
nand I_50416 (I860674,I286286,I286304);
and I_50417 (I860691,I860674,I286295);
DFFARX1 I_50418 (I860691,I3563,I860623,I860717,);
DFFARX1 I_50419 (I860717,I3563,I860623,I860612,);
DFFARX1 I_50420 (I286301,I3563,I860623,I860748,);
nand I_50421 (I860756,I860748,I286298);
not I_50422 (I860773,I860756);
DFFARX1 I_50423 (I860773,I3563,I860623,I860799,);
not I_50424 (I860807,I860799);
nor I_50425 (I860615,I860657,I860807);
DFFARX1 I_50426 (I286292,I3563,I860623,I860847,);
nor I_50427 (I860606,I860847,I860717);
nor I_50428 (I860597,I860847,I860773);
nand I_50429 (I860883,I286283,I286307);
and I_50430 (I860900,I860883,I286286);
DFFARX1 I_50431 (I860900,I3563,I860623,I860926,);
not I_50432 (I860934,I860926);
nand I_50433 (I860951,I860934,I860847);
nand I_50434 (I860600,I860934,I860756);
nor I_50435 (I860982,I286283,I286307);
and I_50436 (I860999,I860847,I860982);
nor I_50437 (I861016,I860934,I860999);
DFFARX1 I_50438 (I861016,I3563,I860623,I860609,);
nor I_50439 (I861047,I860649,I860982);
DFFARX1 I_50440 (I861047,I3563,I860623,I860594,);
nor I_50441 (I861078,I860926,I860982);
not I_50442 (I861095,I861078);
nand I_50443 (I860603,I861095,I860951);
not I_50444 (I861150,I3570);
DFFARX1 I_50445 (I623170,I3563,I861150,I861176,);
not I_50446 (I861184,I861176);
nand I_50447 (I861201,I623155,I623176);
and I_50448 (I861218,I861201,I623164);
DFFARX1 I_50449 (I861218,I3563,I861150,I861244,);
DFFARX1 I_50450 (I861244,I3563,I861150,I861139,);
DFFARX1 I_50451 (I623158,I3563,I861150,I861275,);
nand I_50452 (I861283,I861275,I623167);
not I_50453 (I861300,I861283);
DFFARX1 I_50454 (I861300,I3563,I861150,I861326,);
not I_50455 (I861334,I861326);
nor I_50456 (I861142,I861184,I861334);
DFFARX1 I_50457 (I623173,I3563,I861150,I861374,);
nor I_50458 (I861133,I861374,I861244);
nor I_50459 (I861124,I861374,I861300);
nand I_50460 (I861410,I623155,I623158);
and I_50461 (I861427,I861410,I623179);
DFFARX1 I_50462 (I861427,I3563,I861150,I861453,);
not I_50463 (I861461,I861453);
nand I_50464 (I861478,I861461,I861374);
nand I_50465 (I861127,I861461,I861283);
nor I_50466 (I861509,I623161,I623158);
and I_50467 (I861526,I861374,I861509);
nor I_50468 (I861543,I861461,I861526);
DFFARX1 I_50469 (I861543,I3563,I861150,I861136,);
nor I_50470 (I861574,I861176,I861509);
DFFARX1 I_50471 (I861574,I3563,I861150,I861121,);
nor I_50472 (I861605,I861453,I861509);
not I_50473 (I861622,I861605);
nand I_50474 (I861130,I861622,I861478);
not I_50475 (I861677,I3570);
DFFARX1 I_50476 (I976894,I3563,I861677,I861703,);
not I_50477 (I861711,I861703);
nand I_50478 (I861728,I976909,I976891);
and I_50479 (I861745,I861728,I976891);
DFFARX1 I_50480 (I861745,I3563,I861677,I861771,);
DFFARX1 I_50481 (I861771,I3563,I861677,I861666,);
DFFARX1 I_50482 (I976900,I3563,I861677,I861802,);
nand I_50483 (I861810,I861802,I976918);
not I_50484 (I861827,I861810);
DFFARX1 I_50485 (I861827,I3563,I861677,I861853,);
not I_50486 (I861861,I861853);
nor I_50487 (I861669,I861711,I861861);
DFFARX1 I_50488 (I976915,I3563,I861677,I861901,);
nor I_50489 (I861660,I861901,I861771);
nor I_50490 (I861651,I861901,I861827);
nand I_50491 (I861937,I976912,I976903);
and I_50492 (I861954,I861937,I976897);
DFFARX1 I_50493 (I861954,I3563,I861677,I861980,);
not I_50494 (I861988,I861980);
nand I_50495 (I862005,I861988,I861901);
nand I_50496 (I861654,I861988,I861810);
nor I_50497 (I862036,I976906,I976903);
and I_50498 (I862053,I861901,I862036);
nor I_50499 (I862070,I861988,I862053);
DFFARX1 I_50500 (I862070,I3563,I861677,I861663,);
nor I_50501 (I862101,I861703,I862036);
DFFARX1 I_50502 (I862101,I3563,I861677,I861648,);
nor I_50503 (I862132,I861980,I862036);
not I_50504 (I862149,I862132);
nand I_50505 (I861657,I862149,I862005);
not I_50506 (I862204,I3570);
DFFARX1 I_50507 (I59833,I3563,I862204,I862230,);
not I_50508 (I862238,I862230);
nand I_50509 (I862255,I59809,I59818);
and I_50510 (I862272,I862255,I59812);
DFFARX1 I_50511 (I862272,I3563,I862204,I862298,);
DFFARX1 I_50512 (I862298,I3563,I862204,I862193,);
DFFARX1 I_50513 (I59830,I3563,I862204,I862329,);
nand I_50514 (I862337,I862329,I59821);
not I_50515 (I862354,I862337);
DFFARX1 I_50516 (I862354,I3563,I862204,I862380,);
not I_50517 (I862388,I862380);
nor I_50518 (I862196,I862238,I862388);
DFFARX1 I_50519 (I59815,I3563,I862204,I862428,);
nor I_50520 (I862187,I862428,I862298);
nor I_50521 (I862178,I862428,I862354);
nand I_50522 (I862464,I59827,I59824);
and I_50523 (I862481,I862464,I59812);
DFFARX1 I_50524 (I862481,I3563,I862204,I862507,);
not I_50525 (I862515,I862507);
nand I_50526 (I862532,I862515,I862428);
nand I_50527 (I862181,I862515,I862337);
nor I_50528 (I862563,I59809,I59824);
and I_50529 (I862580,I862428,I862563);
nor I_50530 (I862597,I862515,I862580);
DFFARX1 I_50531 (I862597,I3563,I862204,I862190,);
nor I_50532 (I862628,I862230,I862563);
DFFARX1 I_50533 (I862628,I3563,I862204,I862175,);
nor I_50534 (I862659,I862507,I862563);
not I_50535 (I862676,I862659);
nand I_50536 (I862184,I862676,I862532);
not I_50537 (I862731,I3570);
DFFARX1 I_50538 (I1165575,I3563,I862731,I862757,);
not I_50539 (I862765,I862757);
nand I_50540 (I862782,I1165557,I1165557);
and I_50541 (I862799,I862782,I1165563);
DFFARX1 I_50542 (I862799,I3563,I862731,I862825,);
DFFARX1 I_50543 (I862825,I3563,I862731,I862720,);
DFFARX1 I_50544 (I1165560,I3563,I862731,I862856,);
nand I_50545 (I862864,I862856,I1165569);
not I_50546 (I862881,I862864);
DFFARX1 I_50547 (I862881,I3563,I862731,I862907,);
not I_50548 (I862915,I862907);
nor I_50549 (I862723,I862765,I862915);
DFFARX1 I_50550 (I1165581,I3563,I862731,I862955,);
nor I_50551 (I862714,I862955,I862825);
nor I_50552 (I862705,I862955,I862881);
nand I_50553 (I862991,I1165572,I1165566);
and I_50554 (I863008,I862991,I1165560);
DFFARX1 I_50555 (I863008,I3563,I862731,I863034,);
not I_50556 (I863042,I863034);
nand I_50557 (I863059,I863042,I862955);
nand I_50558 (I862708,I863042,I862864);
nor I_50559 (I863090,I1165578,I1165566);
and I_50560 (I863107,I862955,I863090);
nor I_50561 (I863124,I863042,I863107);
DFFARX1 I_50562 (I863124,I3563,I862731,I862717,);
nor I_50563 (I863155,I862757,I863090);
DFFARX1 I_50564 (I863155,I3563,I862731,I862702,);
nor I_50565 (I863186,I863034,I863090);
not I_50566 (I863203,I863186);
nand I_50567 (I862711,I863203,I863059);
not I_50568 (I863258,I3570);
DFFARX1 I_50569 (I1197943,I3563,I863258,I863284,);
not I_50570 (I863292,I863284);
nand I_50571 (I863309,I1197925,I1197925);
and I_50572 (I863326,I863309,I1197931);
DFFARX1 I_50573 (I863326,I3563,I863258,I863352,);
DFFARX1 I_50574 (I863352,I3563,I863258,I863247,);
DFFARX1 I_50575 (I1197928,I3563,I863258,I863383,);
nand I_50576 (I863391,I863383,I1197937);
not I_50577 (I863408,I863391);
DFFARX1 I_50578 (I863408,I3563,I863258,I863434,);
not I_50579 (I863442,I863434);
nor I_50580 (I863250,I863292,I863442);
DFFARX1 I_50581 (I1197949,I3563,I863258,I863482,);
nor I_50582 (I863241,I863482,I863352);
nor I_50583 (I863232,I863482,I863408);
nand I_50584 (I863518,I1197940,I1197934);
and I_50585 (I863535,I863518,I1197928);
DFFARX1 I_50586 (I863535,I3563,I863258,I863561,);
not I_50587 (I863569,I863561);
nand I_50588 (I863586,I863569,I863482);
nand I_50589 (I863235,I863569,I863391);
nor I_50590 (I863617,I1197946,I1197934);
and I_50591 (I863634,I863482,I863617);
nor I_50592 (I863651,I863569,I863634);
DFFARX1 I_50593 (I863651,I3563,I863258,I863244,);
nor I_50594 (I863682,I863284,I863617);
DFFARX1 I_50595 (I863682,I3563,I863258,I863229,);
nor I_50596 (I863713,I863561,I863617);
not I_50597 (I863730,I863713);
nand I_50598 (I863238,I863730,I863586);
not I_50599 (I863785,I3570);
DFFARX1 I_50600 (I126762,I3563,I863785,I863811,);
not I_50601 (I863819,I863811);
nand I_50602 (I863836,I126738,I126747);
and I_50603 (I863853,I863836,I126741);
DFFARX1 I_50604 (I863853,I3563,I863785,I863879,);
DFFARX1 I_50605 (I863879,I3563,I863785,I863774,);
DFFARX1 I_50606 (I126759,I3563,I863785,I863910,);
nand I_50607 (I863918,I863910,I126750);
not I_50608 (I863935,I863918);
DFFARX1 I_50609 (I863935,I3563,I863785,I863961,);
not I_50610 (I863969,I863961);
nor I_50611 (I863777,I863819,I863969);
DFFARX1 I_50612 (I126744,I3563,I863785,I864009,);
nor I_50613 (I863768,I864009,I863879);
nor I_50614 (I863759,I864009,I863935);
nand I_50615 (I864045,I126756,I126753);
and I_50616 (I864062,I864045,I126741);
DFFARX1 I_50617 (I864062,I3563,I863785,I864088,);
not I_50618 (I864096,I864088);
nand I_50619 (I864113,I864096,I864009);
nand I_50620 (I863762,I864096,I863918);
nor I_50621 (I864144,I126738,I126753);
and I_50622 (I864161,I864009,I864144);
nor I_50623 (I864178,I864096,I864161);
DFFARX1 I_50624 (I864178,I3563,I863785,I863771,);
nor I_50625 (I864209,I863811,I864144);
DFFARX1 I_50626 (I864209,I3563,I863785,I863756,);
nor I_50627 (I864240,I864088,I864144);
not I_50628 (I864257,I864240);
nand I_50629 (I863765,I864257,I864113);
not I_50630 (I864312,I3570);
DFFARX1 I_50631 (I1067425,I3563,I864312,I864338,);
not I_50632 (I864346,I864338);
nand I_50633 (I864363,I1067434,I1067422);
and I_50634 (I864380,I864363,I1067419);
DFFARX1 I_50635 (I864380,I3563,I864312,I864406,);
DFFARX1 I_50636 (I864406,I3563,I864312,I864301,);
DFFARX1 I_50637 (I1067419,I3563,I864312,I864437,);
nand I_50638 (I864445,I864437,I1067416);
not I_50639 (I864462,I864445);
DFFARX1 I_50640 (I864462,I3563,I864312,I864488,);
not I_50641 (I864496,I864488);
nor I_50642 (I864304,I864346,I864496);
DFFARX1 I_50643 (I1067422,I3563,I864312,I864536,);
nor I_50644 (I864295,I864536,I864406);
nor I_50645 (I864286,I864536,I864462);
nand I_50646 (I864572,I1067437,I1067428);
and I_50647 (I864589,I864572,I1067431);
DFFARX1 I_50648 (I864589,I3563,I864312,I864615,);
not I_50649 (I864623,I864615);
nand I_50650 (I864640,I864623,I864536);
nand I_50651 (I864289,I864623,I864445);
nor I_50652 (I864671,I1067416,I1067428);
and I_50653 (I864688,I864536,I864671);
nor I_50654 (I864705,I864623,I864688);
DFFARX1 I_50655 (I864705,I3563,I864312,I864298,);
nor I_50656 (I864736,I864338,I864671);
DFFARX1 I_50657 (I864736,I3563,I864312,I864283,);
nor I_50658 (I864767,I864615,I864671);
not I_50659 (I864784,I864767);
nand I_50660 (I864292,I864784,I864640);
not I_50661 (I864839,I3570);
DFFARX1 I_50662 (I172049,I3563,I864839,I864865,);
not I_50663 (I864873,I864865);
nand I_50664 (I864890,I172046,I172064);
and I_50665 (I864907,I864890,I172055);
DFFARX1 I_50666 (I864907,I3563,I864839,I864933,);
DFFARX1 I_50667 (I864933,I3563,I864839,I864828,);
DFFARX1 I_50668 (I172061,I3563,I864839,I864964,);
nand I_50669 (I864972,I864964,I172058);
not I_50670 (I864989,I864972);
DFFARX1 I_50671 (I864989,I3563,I864839,I865015,);
not I_50672 (I865023,I865015);
nor I_50673 (I864831,I864873,I865023);
DFFARX1 I_50674 (I172052,I3563,I864839,I865063,);
nor I_50675 (I864822,I865063,I864933);
nor I_50676 (I864813,I865063,I864989);
nand I_50677 (I865099,I172043,I172067);
and I_50678 (I865116,I865099,I172046);
DFFARX1 I_50679 (I865116,I3563,I864839,I865142,);
not I_50680 (I865150,I865142);
nand I_50681 (I865167,I865150,I865063);
nand I_50682 (I864816,I865150,I864972);
nor I_50683 (I865198,I172043,I172067);
and I_50684 (I865215,I865063,I865198);
nor I_50685 (I865232,I865150,I865215);
DFFARX1 I_50686 (I865232,I3563,I864839,I864825,);
nor I_50687 (I865263,I864865,I865198);
DFFARX1 I_50688 (I865263,I3563,I864839,I864810,);
nor I_50689 (I865294,I865142,I865198);
not I_50690 (I865311,I865294);
nand I_50691 (I864819,I865311,I865167);
not I_50692 (I865366,I3570);
DFFARX1 I_50693 (I1095637,I3563,I865366,I865392,);
not I_50694 (I865400,I865392);
nand I_50695 (I865417,I1095619,I1095619);
and I_50696 (I865434,I865417,I1095625);
DFFARX1 I_50697 (I865434,I3563,I865366,I865460,);
DFFARX1 I_50698 (I865460,I3563,I865366,I865355,);
DFFARX1 I_50699 (I1095622,I3563,I865366,I865491,);
nand I_50700 (I865499,I865491,I1095631);
not I_50701 (I865516,I865499);
DFFARX1 I_50702 (I865516,I3563,I865366,I865542,);
not I_50703 (I865550,I865542);
nor I_50704 (I865358,I865400,I865550);
DFFARX1 I_50705 (I1095643,I3563,I865366,I865590,);
nor I_50706 (I865349,I865590,I865460);
nor I_50707 (I865340,I865590,I865516);
nand I_50708 (I865626,I1095634,I1095628);
and I_50709 (I865643,I865626,I1095622);
DFFARX1 I_50710 (I865643,I3563,I865366,I865669,);
not I_50711 (I865677,I865669);
nand I_50712 (I865694,I865677,I865590);
nand I_50713 (I865343,I865677,I865499);
nor I_50714 (I865725,I1095640,I1095628);
and I_50715 (I865742,I865590,I865725);
nor I_50716 (I865759,I865677,I865742);
DFFARX1 I_50717 (I865759,I3563,I865366,I865352,);
nor I_50718 (I865790,I865392,I865725);
DFFARX1 I_50719 (I865790,I3563,I865366,I865337,);
nor I_50720 (I865821,I865669,I865725);
not I_50721 (I865838,I865821);
nand I_50722 (I865346,I865838,I865694);
not I_50723 (I865893,I3570);
DFFARX1 I_50724 (I1004672,I3563,I865893,I865919,);
not I_50725 (I865927,I865919);
nand I_50726 (I865944,I1004687,I1004669);
and I_50727 (I865961,I865944,I1004669);
DFFARX1 I_50728 (I865961,I3563,I865893,I865987,);
DFFARX1 I_50729 (I865987,I3563,I865893,I865882,);
DFFARX1 I_50730 (I1004678,I3563,I865893,I866018,);
nand I_50731 (I866026,I866018,I1004696);
not I_50732 (I866043,I866026);
DFFARX1 I_50733 (I866043,I3563,I865893,I866069,);
not I_50734 (I866077,I866069);
nor I_50735 (I865885,I865927,I866077);
DFFARX1 I_50736 (I1004693,I3563,I865893,I866117,);
nor I_50737 (I865876,I866117,I865987);
nor I_50738 (I865867,I866117,I866043);
nand I_50739 (I866153,I1004690,I1004681);
and I_50740 (I866170,I866153,I1004675);
DFFARX1 I_50741 (I866170,I3563,I865893,I866196,);
not I_50742 (I866204,I866196);
nand I_50743 (I866221,I866204,I866117);
nand I_50744 (I865870,I866204,I866026);
nor I_50745 (I866252,I1004684,I1004681);
and I_50746 (I866269,I866117,I866252);
nor I_50747 (I866286,I866204,I866269);
DFFARX1 I_50748 (I866286,I3563,I865893,I865879,);
nor I_50749 (I866317,I865919,I866252);
DFFARX1 I_50750 (I866317,I3563,I865893,I865864,);
nor I_50751 (I866348,I866196,I866252);
not I_50752 (I866365,I866348);
nand I_50753 (I865873,I866365,I866221);
not I_50754 (I866420,I3570);
DFFARX1 I_50755 (I943302,I3563,I866420,I866446,);
not I_50756 (I866454,I866446);
nand I_50757 (I866471,I943317,I943299);
and I_50758 (I866488,I866471,I943299);
DFFARX1 I_50759 (I866488,I3563,I866420,I866514,);
DFFARX1 I_50760 (I866514,I3563,I866420,I866409,);
DFFARX1 I_50761 (I943308,I3563,I866420,I866545,);
nand I_50762 (I866553,I866545,I943326);
not I_50763 (I866570,I866553);
DFFARX1 I_50764 (I866570,I3563,I866420,I866596,);
not I_50765 (I866604,I866596);
nor I_50766 (I866412,I866454,I866604);
DFFARX1 I_50767 (I943323,I3563,I866420,I866644,);
nor I_50768 (I866403,I866644,I866514);
nor I_50769 (I866394,I866644,I866570);
nand I_50770 (I866680,I943320,I943311);
and I_50771 (I866697,I866680,I943305);
DFFARX1 I_50772 (I866697,I3563,I866420,I866723,);
not I_50773 (I866731,I866723);
nand I_50774 (I866748,I866731,I866644);
nand I_50775 (I866397,I866731,I866553);
nor I_50776 (I866779,I943314,I943311);
and I_50777 (I866796,I866644,I866779);
nor I_50778 (I866813,I866731,I866796);
DFFARX1 I_50779 (I866813,I3563,I866420,I866406,);
nor I_50780 (I866844,I866446,I866779);
DFFARX1 I_50781 (I866844,I3563,I866420,I866391,);
nor I_50782 (I866875,I866723,I866779);
not I_50783 (I866892,I866875);
nand I_50784 (I866400,I866892,I866748);
not I_50785 (I866947,I3570);
DFFARX1 I_50786 (I315940,I3563,I866947,I866973,);
not I_50787 (I866981,I866973);
nand I_50788 (I866998,I315931,I315931);
and I_50789 (I867015,I866998,I315949);
DFFARX1 I_50790 (I867015,I3563,I866947,I867041,);
DFFARX1 I_50791 (I867041,I3563,I866947,I866936,);
DFFARX1 I_50792 (I315952,I3563,I866947,I867072,);
nand I_50793 (I867080,I867072,I315934);
not I_50794 (I867097,I867080);
DFFARX1 I_50795 (I867097,I3563,I866947,I867123,);
not I_50796 (I867131,I867123);
nor I_50797 (I866939,I866981,I867131);
DFFARX1 I_50798 (I315946,I3563,I866947,I867171,);
nor I_50799 (I866930,I867171,I867041);
nor I_50800 (I866921,I867171,I867097);
nand I_50801 (I867207,I315958,I315937);
and I_50802 (I867224,I867207,I315943);
DFFARX1 I_50803 (I867224,I3563,I866947,I867250,);
not I_50804 (I867258,I867250);
nand I_50805 (I867275,I867258,I867171);
nand I_50806 (I866924,I867258,I867080);
nor I_50807 (I867306,I315955,I315937);
and I_50808 (I867323,I867171,I867306);
nor I_50809 (I867340,I867258,I867323);
DFFARX1 I_50810 (I867340,I3563,I866947,I866933,);
nor I_50811 (I867371,I866973,I867306);
DFFARX1 I_50812 (I867371,I3563,I866947,I866918,);
nor I_50813 (I867402,I867250,I867306);
not I_50814 (I867419,I867402);
nand I_50815 (I866927,I867419,I867275);
not I_50816 (I867474,I3570);
DFFARX1 I_50817 (I1339873,I3563,I867474,I867500,);
not I_50818 (I867508,I867500);
nand I_50819 (I867525,I1339870,I1339879);
and I_50820 (I867542,I867525,I1339858);
DFFARX1 I_50821 (I867542,I3563,I867474,I867568,);
DFFARX1 I_50822 (I867568,I3563,I867474,I867463,);
DFFARX1 I_50823 (I1339861,I3563,I867474,I867599,);
nand I_50824 (I867607,I867599,I1339876);
not I_50825 (I867624,I867607);
DFFARX1 I_50826 (I867624,I3563,I867474,I867650,);
not I_50827 (I867658,I867650);
nor I_50828 (I867466,I867508,I867658);
DFFARX1 I_50829 (I1339882,I3563,I867474,I867698,);
nor I_50830 (I867457,I867698,I867568);
nor I_50831 (I867448,I867698,I867624);
nand I_50832 (I867734,I1339864,I1339885);
and I_50833 (I867751,I867734,I1339867);
DFFARX1 I_50834 (I867751,I3563,I867474,I867777,);
not I_50835 (I867785,I867777);
nand I_50836 (I867802,I867785,I867698);
nand I_50837 (I867451,I867785,I867607);
nor I_50838 (I867833,I1339858,I1339885);
and I_50839 (I867850,I867698,I867833);
nor I_50840 (I867867,I867785,I867850);
DFFARX1 I_50841 (I867867,I3563,I867474,I867460,);
nor I_50842 (I867898,I867500,I867833);
DFFARX1 I_50843 (I867898,I3563,I867474,I867445,);
nor I_50844 (I867929,I867777,I867833);
not I_50845 (I867946,I867929);
nand I_50846 (I867454,I867946,I867802);
not I_50847 (I868001,I3570);
DFFARX1 I_50848 (I1331543,I3563,I868001,I868027,);
not I_50849 (I868035,I868027);
nand I_50850 (I868052,I1331540,I1331549);
and I_50851 (I868069,I868052,I1331528);
DFFARX1 I_50852 (I868069,I3563,I868001,I868095,);
DFFARX1 I_50853 (I868095,I3563,I868001,I867990,);
DFFARX1 I_50854 (I1331531,I3563,I868001,I868126,);
nand I_50855 (I868134,I868126,I1331546);
not I_50856 (I868151,I868134);
DFFARX1 I_50857 (I868151,I3563,I868001,I868177,);
not I_50858 (I868185,I868177);
nor I_50859 (I867993,I868035,I868185);
DFFARX1 I_50860 (I1331552,I3563,I868001,I868225,);
nor I_50861 (I867984,I868225,I868095);
nor I_50862 (I867975,I868225,I868151);
nand I_50863 (I868261,I1331534,I1331555);
and I_50864 (I868278,I868261,I1331537);
DFFARX1 I_50865 (I868278,I3563,I868001,I868304,);
not I_50866 (I868312,I868304);
nand I_50867 (I868329,I868312,I868225);
nand I_50868 (I867978,I868312,I868134);
nor I_50869 (I868360,I1331528,I1331555);
and I_50870 (I868377,I868225,I868360);
nor I_50871 (I868394,I868312,I868377);
DFFARX1 I_50872 (I868394,I3563,I868001,I867987,);
nor I_50873 (I868425,I868027,I868360);
DFFARX1 I_50874 (I868425,I3563,I868001,I867972,);
nor I_50875 (I868456,I868304,I868360);
not I_50876 (I868473,I868456);
nand I_50877 (I867981,I868473,I868329);
not I_50878 (I868528,I3570);
DFFARX1 I_50879 (I1203145,I3563,I868528,I868554,);
not I_50880 (I868562,I868554);
nand I_50881 (I868579,I1203127,I1203127);
and I_50882 (I868596,I868579,I1203133);
DFFARX1 I_50883 (I868596,I3563,I868528,I868622,);
DFFARX1 I_50884 (I868622,I3563,I868528,I868517,);
DFFARX1 I_50885 (I1203130,I3563,I868528,I868653,);
nand I_50886 (I868661,I868653,I1203139);
not I_50887 (I868678,I868661);
DFFARX1 I_50888 (I868678,I3563,I868528,I868704,);
not I_50889 (I868712,I868704);
nor I_50890 (I868520,I868562,I868712);
DFFARX1 I_50891 (I1203151,I3563,I868528,I868752,);
nor I_50892 (I868511,I868752,I868622);
nor I_50893 (I868502,I868752,I868678);
nand I_50894 (I868788,I1203142,I1203136);
and I_50895 (I868805,I868788,I1203130);
DFFARX1 I_50896 (I868805,I3563,I868528,I868831,);
not I_50897 (I868839,I868831);
nand I_50898 (I868856,I868839,I868752);
nand I_50899 (I868505,I868839,I868661);
nor I_50900 (I868887,I1203148,I1203136);
and I_50901 (I868904,I868752,I868887);
nor I_50902 (I868921,I868839,I868904);
DFFARX1 I_50903 (I868921,I3563,I868528,I868514,);
nor I_50904 (I868952,I868554,I868887);
DFFARX1 I_50905 (I868952,I3563,I868528,I868499,);
nor I_50906 (I868983,I868831,I868887);
not I_50907 (I869000,I868983);
nand I_50908 (I868508,I869000,I868856);
not I_50909 (I869055,I3570);
DFFARX1 I_50910 (I480072,I3563,I869055,I869081,);
not I_50911 (I869089,I869081);
nand I_50912 (I869106,I480069,I480078);
and I_50913 (I869123,I869106,I480087);
DFFARX1 I_50914 (I869123,I3563,I869055,I869149,);
DFFARX1 I_50915 (I869149,I3563,I869055,I869044,);
DFFARX1 I_50916 (I480090,I3563,I869055,I869180,);
nand I_50917 (I869188,I869180,I480093);
not I_50918 (I869205,I869188);
DFFARX1 I_50919 (I869205,I3563,I869055,I869231,);
not I_50920 (I869239,I869231);
nor I_50921 (I869047,I869089,I869239);
DFFARX1 I_50922 (I480066,I3563,I869055,I869279,);
nor I_50923 (I869038,I869279,I869149);
nor I_50924 (I869029,I869279,I869205);
nand I_50925 (I869315,I480081,I480084);
and I_50926 (I869332,I869315,I480075);
DFFARX1 I_50927 (I869332,I3563,I869055,I869358,);
not I_50928 (I869366,I869358);
nand I_50929 (I869383,I869366,I869279);
nand I_50930 (I869032,I869366,I869188);
nor I_50931 (I869414,I480066,I480084);
and I_50932 (I869431,I869279,I869414);
nor I_50933 (I869448,I869366,I869431);
DFFARX1 I_50934 (I869448,I3563,I869055,I869041,);
nor I_50935 (I869479,I869081,I869414);
DFFARX1 I_50936 (I869479,I3563,I869055,I869026,);
nor I_50937 (I869510,I869358,I869414);
not I_50938 (I869527,I869510);
nand I_50939 (I869035,I869527,I869383);
not I_50940 (I869582,I3570);
DFFARX1 I_50941 (I442536,I3563,I869582,I869608,);
not I_50942 (I869616,I869608);
nand I_50943 (I869633,I442533,I442542);
and I_50944 (I869650,I869633,I442551);
DFFARX1 I_50945 (I869650,I3563,I869582,I869676,);
DFFARX1 I_50946 (I869676,I3563,I869582,I869571,);
DFFARX1 I_50947 (I442554,I3563,I869582,I869707,);
nand I_50948 (I869715,I869707,I442557);
not I_50949 (I869732,I869715);
DFFARX1 I_50950 (I869732,I3563,I869582,I869758,);
not I_50951 (I869766,I869758);
nor I_50952 (I869574,I869616,I869766);
DFFARX1 I_50953 (I442530,I3563,I869582,I869806,);
nor I_50954 (I869565,I869806,I869676);
nor I_50955 (I869556,I869806,I869732);
nand I_50956 (I869842,I442545,I442548);
and I_50957 (I869859,I869842,I442539);
DFFARX1 I_50958 (I869859,I3563,I869582,I869885,);
not I_50959 (I869893,I869885);
nand I_50960 (I869910,I869893,I869806);
nand I_50961 (I869559,I869893,I869715);
nor I_50962 (I869941,I442530,I442548);
and I_50963 (I869958,I869806,I869941);
nor I_50964 (I869975,I869893,I869958);
DFFARX1 I_50965 (I869975,I3563,I869582,I869568,);
nor I_50966 (I870006,I869608,I869941);
DFFARX1 I_50967 (I870006,I3563,I869582,I869553,);
nor I_50968 (I870037,I869885,I869941);
not I_50969 (I870054,I870037);
nand I_50970 (I869562,I870054,I869910);
not I_50971 (I870109,I3570);
DFFARX1 I_50972 (I701185,I3563,I870109,I870135,);
not I_50973 (I870143,I870135);
nand I_50974 (I870160,I701188,I701185);
and I_50975 (I870177,I870160,I701197);
DFFARX1 I_50976 (I870177,I3563,I870109,I870203,);
DFFARX1 I_50977 (I870203,I3563,I870109,I870098,);
DFFARX1 I_50978 (I701194,I3563,I870109,I870234,);
nand I_50979 (I870242,I870234,I701200);
not I_50980 (I870259,I870242);
DFFARX1 I_50981 (I870259,I3563,I870109,I870285,);
not I_50982 (I870293,I870285);
nor I_50983 (I870101,I870143,I870293);
DFFARX1 I_50984 (I701209,I3563,I870109,I870333,);
nor I_50985 (I870092,I870333,I870203);
nor I_50986 (I870083,I870333,I870259);
nand I_50987 (I870369,I701203,I701191);
and I_50988 (I870386,I870369,I701188);
DFFARX1 I_50989 (I870386,I3563,I870109,I870412,);
not I_50990 (I870420,I870412);
nand I_50991 (I870437,I870420,I870333);
nand I_50992 (I870086,I870420,I870242);
nor I_50993 (I870468,I701206,I701191);
and I_50994 (I870485,I870333,I870468);
nor I_50995 (I870502,I870420,I870485);
DFFARX1 I_50996 (I870502,I3563,I870109,I870095,);
nor I_50997 (I870533,I870135,I870468);
DFFARX1 I_50998 (I870533,I3563,I870109,I870080,);
nor I_50999 (I870564,I870412,I870468);
not I_51000 (I870581,I870564);
nand I_51001 (I870089,I870581,I870437);
not I_51002 (I870636,I3570);
DFFARX1 I_51003 (I1205457,I3563,I870636,I870662,);
not I_51004 (I870670,I870662);
nand I_51005 (I870687,I1205439,I1205439);
and I_51006 (I870704,I870687,I1205445);
DFFARX1 I_51007 (I870704,I3563,I870636,I870730,);
DFFARX1 I_51008 (I870730,I3563,I870636,I870625,);
DFFARX1 I_51009 (I1205442,I3563,I870636,I870761,);
nand I_51010 (I870769,I870761,I1205451);
not I_51011 (I870786,I870769);
DFFARX1 I_51012 (I870786,I3563,I870636,I870812,);
not I_51013 (I870820,I870812);
nor I_51014 (I870628,I870670,I870820);
DFFARX1 I_51015 (I1205463,I3563,I870636,I870860,);
nor I_51016 (I870619,I870860,I870730);
nor I_51017 (I870610,I870860,I870786);
nand I_51018 (I870896,I1205454,I1205448);
and I_51019 (I870913,I870896,I1205442);
DFFARX1 I_51020 (I870913,I3563,I870636,I870939,);
not I_51021 (I870947,I870939);
nand I_51022 (I870964,I870947,I870860);
nand I_51023 (I870613,I870947,I870769);
nor I_51024 (I870995,I1205460,I1205448);
and I_51025 (I871012,I870860,I870995);
nor I_51026 (I871029,I870947,I871012);
DFFARX1 I_51027 (I871029,I3563,I870636,I870622,);
nor I_51028 (I871060,I870662,I870995);
DFFARX1 I_51029 (I871060,I3563,I870636,I870607,);
nor I_51030 (I871091,I870939,I870995);
not I_51031 (I871108,I871091);
nand I_51032 (I870616,I871108,I870964);
not I_51033 (I871163,I3570);
DFFARX1 I_51034 (I173239,I3563,I871163,I871189,);
not I_51035 (I871197,I871189);
nand I_51036 (I871214,I173236,I173254);
and I_51037 (I871231,I871214,I173245);
DFFARX1 I_51038 (I871231,I3563,I871163,I871257,);
DFFARX1 I_51039 (I871257,I3563,I871163,I871152,);
DFFARX1 I_51040 (I173251,I3563,I871163,I871288,);
nand I_51041 (I871296,I871288,I173248);
not I_51042 (I871313,I871296);
DFFARX1 I_51043 (I871313,I3563,I871163,I871339,);
not I_51044 (I871347,I871339);
nor I_51045 (I871155,I871197,I871347);
DFFARX1 I_51046 (I173242,I3563,I871163,I871387,);
nor I_51047 (I871146,I871387,I871257);
nor I_51048 (I871137,I871387,I871313);
nand I_51049 (I871423,I173233,I173257);
and I_51050 (I871440,I871423,I173236);
DFFARX1 I_51051 (I871440,I3563,I871163,I871466,);
not I_51052 (I871474,I871466);
nand I_51053 (I871491,I871474,I871387);
nand I_51054 (I871140,I871474,I871296);
nor I_51055 (I871522,I173233,I173257);
and I_51056 (I871539,I871387,I871522);
nor I_51057 (I871556,I871474,I871539);
DFFARX1 I_51058 (I871556,I3563,I871163,I871149,);
nor I_51059 (I871587,I871189,I871522);
DFFARX1 I_51060 (I871587,I3563,I871163,I871134,);
nor I_51061 (I871618,I871466,I871522);
not I_51062 (I871635,I871618);
nand I_51063 (I871143,I871635,I871491);
not I_51064 (I871690,I3570);
DFFARX1 I_51065 (I273199,I3563,I871690,I871716,);
not I_51066 (I871724,I871716);
nand I_51067 (I871741,I273196,I273214);
and I_51068 (I871758,I871741,I273205);
DFFARX1 I_51069 (I871758,I3563,I871690,I871784,);
DFFARX1 I_51070 (I871784,I3563,I871690,I871679,);
DFFARX1 I_51071 (I273211,I3563,I871690,I871815,);
nand I_51072 (I871823,I871815,I273208);
not I_51073 (I871840,I871823);
DFFARX1 I_51074 (I871840,I3563,I871690,I871866,);
not I_51075 (I871874,I871866);
nor I_51076 (I871682,I871724,I871874);
DFFARX1 I_51077 (I273202,I3563,I871690,I871914,);
nor I_51078 (I871673,I871914,I871784);
nor I_51079 (I871664,I871914,I871840);
nand I_51080 (I871950,I273193,I273217);
and I_51081 (I871967,I871950,I273196);
DFFARX1 I_51082 (I871967,I3563,I871690,I871993,);
not I_51083 (I872001,I871993);
nand I_51084 (I872018,I872001,I871914);
nand I_51085 (I871667,I872001,I871823);
nor I_51086 (I872049,I273193,I273217);
and I_51087 (I872066,I871914,I872049);
nor I_51088 (I872083,I872001,I872066);
DFFARX1 I_51089 (I872083,I3563,I871690,I871676,);
nor I_51090 (I872114,I871716,I872049);
DFFARX1 I_51091 (I872114,I3563,I871690,I871661,);
nor I_51092 (I872145,I871993,I872049);
not I_51093 (I872162,I872145);
nand I_51094 (I871670,I872162,I872018);
not I_51095 (I872217,I3570);
DFFARX1 I_51096 (I1221063,I3563,I872217,I872243,);
not I_51097 (I872251,I872243);
nand I_51098 (I872268,I1221045,I1221045);
and I_51099 (I872285,I872268,I1221051);
DFFARX1 I_51100 (I872285,I3563,I872217,I872311,);
DFFARX1 I_51101 (I872311,I3563,I872217,I872206,);
DFFARX1 I_51102 (I1221048,I3563,I872217,I872342,);
nand I_51103 (I872350,I872342,I1221057);
not I_51104 (I872367,I872350);
DFFARX1 I_51105 (I872367,I3563,I872217,I872393,);
not I_51106 (I872401,I872393);
nor I_51107 (I872209,I872251,I872401);
DFFARX1 I_51108 (I1221069,I3563,I872217,I872441,);
nor I_51109 (I872200,I872441,I872311);
nor I_51110 (I872191,I872441,I872367);
nand I_51111 (I872477,I1221060,I1221054);
and I_51112 (I872494,I872477,I1221048);
DFFARX1 I_51113 (I872494,I3563,I872217,I872520,);
not I_51114 (I872528,I872520);
nand I_51115 (I872545,I872528,I872441);
nand I_51116 (I872194,I872528,I872350);
nor I_51117 (I872576,I1221066,I1221054);
and I_51118 (I872593,I872441,I872576);
nor I_51119 (I872610,I872528,I872593);
DFFARX1 I_51120 (I872610,I3563,I872217,I872203,);
nor I_51121 (I872641,I872243,I872576);
DFFARX1 I_51122 (I872641,I3563,I872217,I872188,);
nor I_51123 (I872672,I872520,I872576);
not I_51124 (I872689,I872672);
nand I_51125 (I872197,I872689,I872545);
not I_51126 (I872744,I3570);
DFFARX1 I_51127 (I693093,I3563,I872744,I872770,);
not I_51128 (I872778,I872770);
nand I_51129 (I872795,I693096,I693093);
and I_51130 (I872812,I872795,I693105);
DFFARX1 I_51131 (I872812,I3563,I872744,I872838,);
DFFARX1 I_51132 (I872838,I3563,I872744,I872733,);
DFFARX1 I_51133 (I693102,I3563,I872744,I872869,);
nand I_51134 (I872877,I872869,I693108);
not I_51135 (I872894,I872877);
DFFARX1 I_51136 (I872894,I3563,I872744,I872920,);
not I_51137 (I872928,I872920);
nor I_51138 (I872736,I872778,I872928);
DFFARX1 I_51139 (I693117,I3563,I872744,I872968,);
nor I_51140 (I872727,I872968,I872838);
nor I_51141 (I872718,I872968,I872894);
nand I_51142 (I873004,I693111,I693099);
and I_51143 (I873021,I873004,I693096);
DFFARX1 I_51144 (I873021,I3563,I872744,I873047,);
not I_51145 (I873055,I873047);
nand I_51146 (I873072,I873055,I872968);
nand I_51147 (I872721,I873055,I872877);
nor I_51148 (I873103,I693114,I693099);
and I_51149 (I873120,I872968,I873103);
nor I_51150 (I873137,I873055,I873120);
DFFARX1 I_51151 (I873137,I3563,I872744,I872730,);
nor I_51152 (I873168,I872770,I873103);
DFFARX1 I_51153 (I873168,I3563,I872744,I872715,);
nor I_51154 (I873199,I873047,I873103);
not I_51155 (I873216,I873199);
nand I_51156 (I872724,I873216,I873072);
not I_51157 (I873271,I3570);
DFFARX1 I_51158 (I366532,I3563,I873271,I873297,);
not I_51159 (I873305,I873297);
nand I_51160 (I873322,I366523,I366523);
and I_51161 (I873339,I873322,I366541);
DFFARX1 I_51162 (I873339,I3563,I873271,I873365,);
DFFARX1 I_51163 (I873365,I3563,I873271,I873260,);
DFFARX1 I_51164 (I366544,I3563,I873271,I873396,);
nand I_51165 (I873404,I873396,I366526);
not I_51166 (I873421,I873404);
DFFARX1 I_51167 (I873421,I3563,I873271,I873447,);
not I_51168 (I873455,I873447);
nor I_51169 (I873263,I873305,I873455);
DFFARX1 I_51170 (I366538,I3563,I873271,I873495,);
nor I_51171 (I873254,I873495,I873365);
nor I_51172 (I873245,I873495,I873421);
nand I_51173 (I873531,I366550,I366529);
and I_51174 (I873548,I873531,I366535);
DFFARX1 I_51175 (I873548,I3563,I873271,I873574,);
not I_51176 (I873582,I873574);
nand I_51177 (I873599,I873582,I873495);
nand I_51178 (I873248,I873582,I873404);
nor I_51179 (I873630,I366547,I366529);
and I_51180 (I873647,I873495,I873630);
nor I_51181 (I873664,I873582,I873647);
DFFARX1 I_51182 (I873664,I3563,I873271,I873257,);
nor I_51183 (I873695,I873297,I873630);
DFFARX1 I_51184 (I873695,I3563,I873271,I873242,);
nor I_51185 (I873726,I873574,I873630);
not I_51186 (I873743,I873726);
nand I_51187 (I873251,I873743,I873599);
not I_51188 (I873798,I3570);
DFFARX1 I_51189 (I786729,I3563,I873798,I873824,);
not I_51190 (I873832,I873824);
nand I_51191 (I873849,I786732,I786729);
and I_51192 (I873866,I873849,I786741);
DFFARX1 I_51193 (I873866,I3563,I873798,I873892,);
DFFARX1 I_51194 (I873892,I3563,I873798,I873787,);
DFFARX1 I_51195 (I786738,I3563,I873798,I873923,);
nand I_51196 (I873931,I873923,I786744);
not I_51197 (I873948,I873931);
DFFARX1 I_51198 (I873948,I3563,I873798,I873974,);
not I_51199 (I873982,I873974);
nor I_51200 (I873790,I873832,I873982);
DFFARX1 I_51201 (I786753,I3563,I873798,I874022,);
nor I_51202 (I873781,I874022,I873892);
nor I_51203 (I873772,I874022,I873948);
nand I_51204 (I874058,I786747,I786735);
and I_51205 (I874075,I874058,I786732);
DFFARX1 I_51206 (I874075,I3563,I873798,I874101,);
not I_51207 (I874109,I874101);
nand I_51208 (I874126,I874109,I874022);
nand I_51209 (I873775,I874109,I873931);
nor I_51210 (I874157,I786750,I786735);
and I_51211 (I874174,I874022,I874157);
nor I_51212 (I874191,I874109,I874174);
DFFARX1 I_51213 (I874191,I3563,I873798,I873784,);
nor I_51214 (I874222,I873824,I874157);
DFFARX1 I_51215 (I874222,I3563,I873798,I873769,);
nor I_51216 (I874253,I874101,I874157);
not I_51217 (I874270,I874253);
nand I_51218 (I873778,I874270,I874126);
not I_51219 (I874325,I3570);
DFFARX1 I_51220 (I106209,I3563,I874325,I874351,);
not I_51221 (I874359,I874351);
nand I_51222 (I874376,I106185,I106194);
and I_51223 (I874393,I874376,I106188);
DFFARX1 I_51224 (I874393,I3563,I874325,I874419,);
DFFARX1 I_51225 (I874419,I3563,I874325,I874314,);
DFFARX1 I_51226 (I106206,I3563,I874325,I874450,);
nand I_51227 (I874458,I874450,I106197);
not I_51228 (I874475,I874458);
DFFARX1 I_51229 (I874475,I3563,I874325,I874501,);
not I_51230 (I874509,I874501);
nor I_51231 (I874317,I874359,I874509);
DFFARX1 I_51232 (I106191,I3563,I874325,I874549,);
nor I_51233 (I874308,I874549,I874419);
nor I_51234 (I874299,I874549,I874475);
nand I_51235 (I874585,I106203,I106200);
and I_51236 (I874602,I874585,I106188);
DFFARX1 I_51237 (I874602,I3563,I874325,I874628,);
not I_51238 (I874636,I874628);
nand I_51239 (I874653,I874636,I874549);
nand I_51240 (I874302,I874636,I874458);
nor I_51241 (I874684,I106185,I106200);
and I_51242 (I874701,I874549,I874684);
nor I_51243 (I874718,I874636,I874701);
DFFARX1 I_51244 (I874718,I3563,I874325,I874311,);
nor I_51245 (I874749,I874351,I874684);
DFFARX1 I_51246 (I874749,I3563,I874325,I874296,);
nor I_51247 (I874780,I874628,I874684);
not I_51248 (I874797,I874780);
nand I_51249 (I874305,I874797,I874653);
not I_51250 (I874852,I3570);
DFFARX1 I_51251 (I468104,I3563,I874852,I874878,);
not I_51252 (I874886,I874878);
nand I_51253 (I874903,I468101,I468110);
and I_51254 (I874920,I874903,I468119);
DFFARX1 I_51255 (I874920,I3563,I874852,I874946,);
DFFARX1 I_51256 (I874946,I3563,I874852,I874841,);
DFFARX1 I_51257 (I468122,I3563,I874852,I874977,);
nand I_51258 (I874985,I874977,I468125);
not I_51259 (I875002,I874985);
DFFARX1 I_51260 (I875002,I3563,I874852,I875028,);
not I_51261 (I875036,I875028);
nor I_51262 (I874844,I874886,I875036);
DFFARX1 I_51263 (I468098,I3563,I874852,I875076,);
nor I_51264 (I874835,I875076,I874946);
nor I_51265 (I874826,I875076,I875002);
nand I_51266 (I875112,I468113,I468116);
and I_51267 (I875129,I875112,I468107);
DFFARX1 I_51268 (I875129,I3563,I874852,I875155,);
not I_51269 (I875163,I875155);
nand I_51270 (I875180,I875163,I875076);
nand I_51271 (I874829,I875163,I874985);
nor I_51272 (I875211,I468098,I468116);
and I_51273 (I875228,I875076,I875211);
nor I_51274 (I875245,I875163,I875228);
DFFARX1 I_51275 (I875245,I3563,I874852,I874838,);
nor I_51276 (I875276,I874878,I875211);
DFFARX1 I_51277 (I875276,I3563,I874852,I874823,);
nor I_51278 (I875307,I875155,I875211);
not I_51279 (I875324,I875307);
nand I_51280 (I874832,I875324,I875180);
not I_51281 (I875379,I3570);
DFFARX1 I_51282 (I925860,I3563,I875379,I875405,);
not I_51283 (I875413,I875405);
nand I_51284 (I875430,I925875,I925857);
and I_51285 (I875447,I875430,I925857);
DFFARX1 I_51286 (I875447,I3563,I875379,I875473,);
DFFARX1 I_51287 (I875473,I3563,I875379,I875368,);
DFFARX1 I_51288 (I925866,I3563,I875379,I875504,);
nand I_51289 (I875512,I875504,I925884);
not I_51290 (I875529,I875512);
DFFARX1 I_51291 (I875529,I3563,I875379,I875555,);
not I_51292 (I875563,I875555);
nor I_51293 (I875371,I875413,I875563);
DFFARX1 I_51294 (I925881,I3563,I875379,I875603,);
nor I_51295 (I875362,I875603,I875473);
nor I_51296 (I875353,I875603,I875529);
nand I_51297 (I875639,I925878,I925869);
and I_51298 (I875656,I875639,I925863);
DFFARX1 I_51299 (I875656,I3563,I875379,I875682,);
not I_51300 (I875690,I875682);
nand I_51301 (I875707,I875690,I875603);
nand I_51302 (I875356,I875690,I875512);
nor I_51303 (I875738,I925872,I925869);
and I_51304 (I875755,I875603,I875738);
nor I_51305 (I875772,I875690,I875755);
DFFARX1 I_51306 (I875772,I3563,I875379,I875365,);
nor I_51307 (I875803,I875405,I875738);
DFFARX1 I_51308 (I875803,I3563,I875379,I875350,);
nor I_51309 (I875834,I875682,I875738);
not I_51310 (I875851,I875834);
nand I_51311 (I875359,I875851,I875707);
not I_51312 (I875906,I3570);
DFFARX1 I_51313 (I545947,I3563,I875906,I875932,);
not I_51314 (I875940,I875932);
nand I_51315 (I875957,I545965,I545956);
and I_51316 (I875974,I875957,I545959);
DFFARX1 I_51317 (I875974,I3563,I875906,I876000,);
DFFARX1 I_51318 (I876000,I3563,I875906,I875895,);
DFFARX1 I_51319 (I545953,I3563,I875906,I876031,);
nand I_51320 (I876039,I876031,I545944);
not I_51321 (I876056,I876039);
DFFARX1 I_51322 (I876056,I3563,I875906,I876082,);
not I_51323 (I876090,I876082);
nor I_51324 (I875898,I875940,I876090);
DFFARX1 I_51325 (I545950,I3563,I875906,I876130,);
nor I_51326 (I875889,I876130,I876000);
nor I_51327 (I875880,I876130,I876056);
nand I_51328 (I876166,I545944,I545941);
and I_51329 (I876183,I876166,I545962);
DFFARX1 I_51330 (I876183,I3563,I875906,I876209,);
not I_51331 (I876217,I876209);
nand I_51332 (I876234,I876217,I876130);
nand I_51333 (I875883,I876217,I876039);
nor I_51334 (I876265,I545941,I545941);
and I_51335 (I876282,I876130,I876265);
nor I_51336 (I876299,I876217,I876282);
DFFARX1 I_51337 (I876299,I3563,I875906,I875892,);
nor I_51338 (I876330,I875932,I876265);
DFFARX1 I_51339 (I876330,I3563,I875906,I875877,);
nor I_51340 (I876361,I876209,I876265);
not I_51341 (I876378,I876361);
nand I_51342 (I875886,I876378,I876234);
not I_51343 (I876433,I3570);
DFFARX1 I_51344 (I1167887,I3563,I876433,I876459,);
not I_51345 (I876467,I876459);
nand I_51346 (I876484,I1167869,I1167869);
and I_51347 (I876501,I876484,I1167875);
DFFARX1 I_51348 (I876501,I3563,I876433,I876527,);
DFFARX1 I_51349 (I876527,I3563,I876433,I876422,);
DFFARX1 I_51350 (I1167872,I3563,I876433,I876558,);
nand I_51351 (I876566,I876558,I1167881);
not I_51352 (I876583,I876566);
DFFARX1 I_51353 (I876583,I3563,I876433,I876609,);
not I_51354 (I876617,I876609);
nor I_51355 (I876425,I876467,I876617);
DFFARX1 I_51356 (I1167893,I3563,I876433,I876657,);
nor I_51357 (I876416,I876657,I876527);
nor I_51358 (I876407,I876657,I876583);
nand I_51359 (I876693,I1167884,I1167878);
and I_51360 (I876710,I876693,I1167872);
DFFARX1 I_51361 (I876710,I3563,I876433,I876736,);
not I_51362 (I876744,I876736);
nand I_51363 (I876761,I876744,I876657);
nand I_51364 (I876410,I876744,I876566);
nor I_51365 (I876792,I1167890,I1167878);
and I_51366 (I876809,I876657,I876792);
nor I_51367 (I876826,I876744,I876809);
DFFARX1 I_51368 (I876826,I3563,I876433,I876419,);
nor I_51369 (I876857,I876459,I876792);
DFFARX1 I_51370 (I876857,I3563,I876433,I876404,);
nor I_51371 (I876888,I876736,I876792);
not I_51372 (I876905,I876888);
nand I_51373 (I876413,I876905,I876761);
not I_51374 (I876960,I3570);
DFFARX1 I_51375 (I473000,I3563,I876960,I876986,);
not I_51376 (I876994,I876986);
nand I_51377 (I877011,I472997,I473006);
and I_51378 (I877028,I877011,I473015);
DFFARX1 I_51379 (I877028,I3563,I876960,I877054,);
DFFARX1 I_51380 (I877054,I3563,I876960,I876949,);
DFFARX1 I_51381 (I473018,I3563,I876960,I877085,);
nand I_51382 (I877093,I877085,I473021);
not I_51383 (I877110,I877093);
DFFARX1 I_51384 (I877110,I3563,I876960,I877136,);
not I_51385 (I877144,I877136);
nor I_51386 (I876952,I876994,I877144);
DFFARX1 I_51387 (I472994,I3563,I876960,I877184,);
nor I_51388 (I876943,I877184,I877054);
nor I_51389 (I876934,I877184,I877110);
nand I_51390 (I877220,I473009,I473012);
and I_51391 (I877237,I877220,I473003);
DFFARX1 I_51392 (I877237,I3563,I876960,I877263,);
not I_51393 (I877271,I877263);
nand I_51394 (I877288,I877271,I877184);
nand I_51395 (I876937,I877271,I877093);
nor I_51396 (I877319,I472994,I473012);
and I_51397 (I877336,I877184,I877319);
nor I_51398 (I877353,I877271,I877336);
DFFARX1 I_51399 (I877353,I3563,I876960,I876946,);
nor I_51400 (I877384,I876986,I877319);
DFFARX1 I_51401 (I877384,I3563,I876960,I876931,);
nor I_51402 (I877415,I877263,I877319);
not I_51403 (I877432,I877415);
nand I_51404 (I876940,I877432,I877288);
not I_51405 (I877487,I3570);
DFFARX1 I_51406 (I274984,I3563,I877487,I877513,);
not I_51407 (I877521,I877513);
nand I_51408 (I877538,I274981,I274999);
and I_51409 (I877555,I877538,I274990);
DFFARX1 I_51410 (I877555,I3563,I877487,I877581,);
DFFARX1 I_51411 (I877581,I3563,I877487,I877476,);
DFFARX1 I_51412 (I274996,I3563,I877487,I877612,);
nand I_51413 (I877620,I877612,I274993);
not I_51414 (I877637,I877620);
DFFARX1 I_51415 (I877637,I3563,I877487,I877663,);
not I_51416 (I877671,I877663);
nor I_51417 (I877479,I877521,I877671);
DFFARX1 I_51418 (I274987,I3563,I877487,I877711,);
nor I_51419 (I877470,I877711,I877581);
nor I_51420 (I877461,I877711,I877637);
nand I_51421 (I877747,I274978,I275002);
and I_51422 (I877764,I877747,I274981);
DFFARX1 I_51423 (I877764,I3563,I877487,I877790,);
not I_51424 (I877798,I877790);
nand I_51425 (I877815,I877798,I877711);
nand I_51426 (I877464,I877798,I877620);
nor I_51427 (I877846,I274978,I275002);
and I_51428 (I877863,I877711,I877846);
nor I_51429 (I877880,I877798,I877863);
DFFARX1 I_51430 (I877880,I3563,I877487,I877473,);
nor I_51431 (I877911,I877513,I877846);
DFFARX1 I_51432 (I877911,I3563,I877487,I877458,);
nor I_51433 (I877942,I877790,I877846);
not I_51434 (I877959,I877942);
nand I_51435 (I877467,I877959,I877815);
not I_51436 (I878014,I3570);
DFFARX1 I_51437 (I1118757,I3563,I878014,I878040,);
not I_51438 (I878048,I878040);
nand I_51439 (I878065,I1118739,I1118739);
and I_51440 (I878082,I878065,I1118745);
DFFARX1 I_51441 (I878082,I3563,I878014,I878108,);
DFFARX1 I_51442 (I878108,I3563,I878014,I878003,);
DFFARX1 I_51443 (I1118742,I3563,I878014,I878139,);
nand I_51444 (I878147,I878139,I1118751);
not I_51445 (I878164,I878147);
DFFARX1 I_51446 (I878164,I3563,I878014,I878190,);
not I_51447 (I878198,I878190);
nor I_51448 (I878006,I878048,I878198);
DFFARX1 I_51449 (I1118763,I3563,I878014,I878238,);
nor I_51450 (I877997,I878238,I878108);
nor I_51451 (I877988,I878238,I878164);
nand I_51452 (I878274,I1118754,I1118748);
and I_51453 (I878291,I878274,I1118742);
DFFARX1 I_51454 (I878291,I3563,I878014,I878317,);
not I_51455 (I878325,I878317);
nand I_51456 (I878342,I878325,I878238);
nand I_51457 (I877991,I878325,I878147);
nor I_51458 (I878373,I1118760,I1118748);
and I_51459 (I878390,I878238,I878373);
nor I_51460 (I878407,I878325,I878390);
DFFARX1 I_51461 (I878407,I3563,I878014,I878000,);
nor I_51462 (I878438,I878040,I878373);
DFFARX1 I_51463 (I878438,I3563,I878014,I877985,);
nor I_51464 (I878469,I878317,I878373);
not I_51465 (I878486,I878469);
nand I_51466 (I877994,I878486,I878342);
not I_51467 (I878541,I3570);
DFFARX1 I_51468 (I708699,I3563,I878541,I878567,);
not I_51469 (I878575,I878567);
nand I_51470 (I878592,I708702,I708699);
and I_51471 (I878609,I878592,I708711);
DFFARX1 I_51472 (I878609,I3563,I878541,I878635,);
DFFARX1 I_51473 (I878635,I3563,I878541,I878530,);
DFFARX1 I_51474 (I708708,I3563,I878541,I878666,);
nand I_51475 (I878674,I878666,I708714);
not I_51476 (I878691,I878674);
DFFARX1 I_51477 (I878691,I3563,I878541,I878717,);
not I_51478 (I878725,I878717);
nor I_51479 (I878533,I878575,I878725);
DFFARX1 I_51480 (I708723,I3563,I878541,I878765,);
nor I_51481 (I878524,I878765,I878635);
nor I_51482 (I878515,I878765,I878691);
nand I_51483 (I878801,I708717,I708705);
and I_51484 (I878818,I878801,I708702);
DFFARX1 I_51485 (I878818,I3563,I878541,I878844,);
not I_51486 (I878852,I878844);
nand I_51487 (I878869,I878852,I878765);
nand I_51488 (I878518,I878852,I878674);
nor I_51489 (I878900,I708720,I708705);
and I_51490 (I878917,I878765,I878900);
nor I_51491 (I878934,I878852,I878917);
DFFARX1 I_51492 (I878934,I3563,I878541,I878527,);
nor I_51493 (I878965,I878567,I878900);
DFFARX1 I_51494 (I878965,I3563,I878541,I878512,);
nor I_51495 (I878996,I878844,I878900);
not I_51496 (I879013,I878996);
nand I_51497 (I878521,I879013,I878869);
not I_51498 (I879068,I3570);
DFFARX1 I_51499 (I623748,I3563,I879068,I879094,);
not I_51500 (I879102,I879094);
nand I_51501 (I879119,I623733,I623754);
and I_51502 (I879136,I879119,I623742);
DFFARX1 I_51503 (I879136,I3563,I879068,I879162,);
DFFARX1 I_51504 (I879162,I3563,I879068,I879057,);
DFFARX1 I_51505 (I623736,I3563,I879068,I879193,);
nand I_51506 (I879201,I879193,I623745);
not I_51507 (I879218,I879201);
DFFARX1 I_51508 (I879218,I3563,I879068,I879244,);
not I_51509 (I879252,I879244);
nor I_51510 (I879060,I879102,I879252);
DFFARX1 I_51511 (I623751,I3563,I879068,I879292,);
nor I_51512 (I879051,I879292,I879162);
nor I_51513 (I879042,I879292,I879218);
nand I_51514 (I879328,I623733,I623736);
and I_51515 (I879345,I879328,I623757);
DFFARX1 I_51516 (I879345,I3563,I879068,I879371,);
not I_51517 (I879379,I879371);
nand I_51518 (I879396,I879379,I879292);
nand I_51519 (I879045,I879379,I879201);
nor I_51520 (I879427,I623739,I623736);
and I_51521 (I879444,I879292,I879427);
nor I_51522 (I879461,I879379,I879444);
DFFARX1 I_51523 (I879461,I3563,I879068,I879054,);
nor I_51524 (I879492,I879094,I879427);
DFFARX1 I_51525 (I879492,I3563,I879068,I879039,);
nor I_51526 (I879523,I879371,I879427);
not I_51527 (I879540,I879523);
nand I_51528 (I879048,I879540,I879396);
not I_51529 (I879595,I3570);
DFFARX1 I_51530 (I721415,I3563,I879595,I879621,);
not I_51531 (I879629,I879621);
nand I_51532 (I879646,I721418,I721415);
and I_51533 (I879663,I879646,I721427);
DFFARX1 I_51534 (I879663,I3563,I879595,I879689,);
DFFARX1 I_51535 (I879689,I3563,I879595,I879584,);
DFFARX1 I_51536 (I721424,I3563,I879595,I879720,);
nand I_51537 (I879728,I879720,I721430);
not I_51538 (I879745,I879728);
DFFARX1 I_51539 (I879745,I3563,I879595,I879771,);
not I_51540 (I879779,I879771);
nor I_51541 (I879587,I879629,I879779);
DFFARX1 I_51542 (I721439,I3563,I879595,I879819,);
nor I_51543 (I879578,I879819,I879689);
nor I_51544 (I879569,I879819,I879745);
nand I_51545 (I879855,I721433,I721421);
and I_51546 (I879872,I879855,I721418);
DFFARX1 I_51547 (I879872,I3563,I879595,I879898,);
not I_51548 (I879906,I879898);
nand I_51549 (I879923,I879906,I879819);
nand I_51550 (I879572,I879906,I879728);
nor I_51551 (I879954,I721436,I721421);
and I_51552 (I879971,I879819,I879954);
nor I_51553 (I879988,I879906,I879971);
DFFARX1 I_51554 (I879988,I3563,I879595,I879581,);
nor I_51555 (I880019,I879621,I879954);
DFFARX1 I_51556 (I880019,I3563,I879595,I879566,);
nor I_51557 (I880050,I879898,I879954);
not I_51558 (I880067,I880050);
nand I_51559 (I879575,I880067,I879923);
not I_51560 (I880122,I3570);
DFFARX1 I_51561 (I1115289,I3563,I880122,I880148,);
not I_51562 (I880156,I880148);
nand I_51563 (I880173,I1115271,I1115271);
and I_51564 (I880190,I880173,I1115277);
DFFARX1 I_51565 (I880190,I3563,I880122,I880216,);
DFFARX1 I_51566 (I880216,I3563,I880122,I880111,);
DFFARX1 I_51567 (I1115274,I3563,I880122,I880247,);
nand I_51568 (I880255,I880247,I1115283);
not I_51569 (I880272,I880255);
DFFARX1 I_51570 (I880272,I3563,I880122,I880298,);
not I_51571 (I880306,I880298);
nor I_51572 (I880114,I880156,I880306);
DFFARX1 I_51573 (I1115295,I3563,I880122,I880346,);
nor I_51574 (I880105,I880346,I880216);
nor I_51575 (I880096,I880346,I880272);
nand I_51576 (I880382,I1115286,I1115280);
and I_51577 (I880399,I880382,I1115274);
DFFARX1 I_51578 (I880399,I3563,I880122,I880425,);
not I_51579 (I880433,I880425);
nand I_51580 (I880450,I880433,I880346);
nand I_51581 (I880099,I880433,I880255);
nor I_51582 (I880481,I1115292,I1115280);
and I_51583 (I880498,I880346,I880481);
nor I_51584 (I880515,I880433,I880498);
DFFARX1 I_51585 (I880515,I3563,I880122,I880108,);
nor I_51586 (I880546,I880148,I880481);
DFFARX1 I_51587 (I880546,I3563,I880122,I880093,);
nor I_51588 (I880577,I880425,I880481);
not I_51589 (I880594,I880577);
nand I_51590 (I880102,I880594,I880450);
not I_51591 (I880649,I3570);
DFFARX1 I_51592 (I790197,I3563,I880649,I880675,);
not I_51593 (I880683,I880675);
nand I_51594 (I880700,I790200,I790197);
and I_51595 (I880717,I880700,I790209);
DFFARX1 I_51596 (I880717,I3563,I880649,I880743,);
DFFARX1 I_51597 (I880743,I3563,I880649,I880638,);
DFFARX1 I_51598 (I790206,I3563,I880649,I880774,);
nand I_51599 (I880782,I880774,I790212);
not I_51600 (I880799,I880782);
DFFARX1 I_51601 (I880799,I3563,I880649,I880825,);
not I_51602 (I880833,I880825);
nor I_51603 (I880641,I880683,I880833);
DFFARX1 I_51604 (I790221,I3563,I880649,I880873,);
nor I_51605 (I880632,I880873,I880743);
nor I_51606 (I880623,I880873,I880799);
nand I_51607 (I880909,I790215,I790203);
and I_51608 (I880926,I880909,I790200);
DFFARX1 I_51609 (I880926,I3563,I880649,I880952,);
not I_51610 (I880960,I880952);
nand I_51611 (I880977,I880960,I880873);
nand I_51612 (I880626,I880960,I880782);
nor I_51613 (I881008,I790218,I790203);
and I_51614 (I881025,I880873,I881008);
nor I_51615 (I881042,I880960,I881025);
DFFARX1 I_51616 (I881042,I3563,I880649,I880635,);
nor I_51617 (I881073,I880675,I881008);
DFFARX1 I_51618 (I881073,I3563,I880649,I880620,);
nor I_51619 (I881104,I880952,I881008);
not I_51620 (I881121,I881104);
nand I_51621 (I880629,I881121,I880977);
not I_51622 (I881176,I3570);
DFFARX1 I_51623 (I791931,I3563,I881176,I881202,);
not I_51624 (I881210,I881202);
nand I_51625 (I881227,I791934,I791931);
and I_51626 (I881244,I881227,I791943);
DFFARX1 I_51627 (I881244,I3563,I881176,I881270,);
DFFARX1 I_51628 (I881270,I3563,I881176,I881165,);
DFFARX1 I_51629 (I791940,I3563,I881176,I881301,);
nand I_51630 (I881309,I881301,I791946);
not I_51631 (I881326,I881309);
DFFARX1 I_51632 (I881326,I3563,I881176,I881352,);
not I_51633 (I881360,I881352);
nor I_51634 (I881168,I881210,I881360);
DFFARX1 I_51635 (I791955,I3563,I881176,I881400,);
nor I_51636 (I881159,I881400,I881270);
nor I_51637 (I881150,I881400,I881326);
nand I_51638 (I881436,I791949,I791937);
and I_51639 (I881453,I881436,I791934);
DFFARX1 I_51640 (I881453,I3563,I881176,I881479,);
not I_51641 (I881487,I881479);
nand I_51642 (I881504,I881487,I881400);
nand I_51643 (I881153,I881487,I881309);
nor I_51644 (I881535,I791952,I791937);
and I_51645 (I881552,I881400,I881535);
nor I_51646 (I881569,I881487,I881552);
DFFARX1 I_51647 (I881569,I3563,I881176,I881162,);
nor I_51648 (I881600,I881202,I881535);
DFFARX1 I_51649 (I881600,I3563,I881176,I881147,);
nor I_51650 (I881631,I881479,I881535);
not I_51651 (I881648,I881631);
nand I_51652 (I881156,I881648,I881504);
not I_51653 (I881703,I3570);
DFFARX1 I_51654 (I245234,I3563,I881703,I881729,);
not I_51655 (I881737,I881729);
nand I_51656 (I881754,I245231,I245249);
and I_51657 (I881771,I881754,I245240);
DFFARX1 I_51658 (I881771,I3563,I881703,I881797,);
DFFARX1 I_51659 (I881797,I3563,I881703,I881692,);
DFFARX1 I_51660 (I245246,I3563,I881703,I881828,);
nand I_51661 (I881836,I881828,I245243);
not I_51662 (I881853,I881836);
DFFARX1 I_51663 (I881853,I3563,I881703,I881879,);
not I_51664 (I881887,I881879);
nor I_51665 (I881695,I881737,I881887);
DFFARX1 I_51666 (I245237,I3563,I881703,I881927,);
nor I_51667 (I881686,I881927,I881797);
nor I_51668 (I881677,I881927,I881853);
nand I_51669 (I881963,I245228,I245252);
and I_51670 (I881980,I881963,I245231);
DFFARX1 I_51671 (I881980,I3563,I881703,I882006,);
not I_51672 (I882014,I882006);
nand I_51673 (I882031,I882014,I881927);
nand I_51674 (I881680,I882014,I881836);
nor I_51675 (I882062,I245228,I245252);
and I_51676 (I882079,I881927,I882062);
nor I_51677 (I882096,I882014,I882079);
DFFARX1 I_51678 (I882096,I3563,I881703,I881689,);
nor I_51679 (I882127,I881729,I882062);
DFFARX1 I_51680 (I882127,I3563,I881703,I881674,);
nor I_51681 (I882158,I882006,I882062);
not I_51682 (I882175,I882158);
nand I_51683 (I881683,I882175,I882031);
not I_51684 (I882230,I3570);
DFFARX1 I_51685 (I1492,I3563,I882230,I882256,);
not I_51686 (I882264,I882256);
nand I_51687 (I882281,I2100,I2724);
and I_51688 (I882298,I882281,I2444);
DFFARX1 I_51689 (I882298,I3563,I882230,I882324,);
DFFARX1 I_51690 (I882324,I3563,I882230,I882219,);
DFFARX1 I_51691 (I3476,I3563,I882230,I882355,);
nand I_51692 (I882363,I882355,I1828);
not I_51693 (I882380,I882363);
DFFARX1 I_51694 (I882380,I3563,I882230,I882406,);
not I_51695 (I882414,I882406);
nor I_51696 (I882222,I882264,I882414);
DFFARX1 I_51697 (I2220,I3563,I882230,I882454,);
nor I_51698 (I882213,I882454,I882324);
nor I_51699 (I882204,I882454,I882380);
nand I_51700 (I882490,I2196,I1380);
and I_51701 (I882507,I882490,I3156);
DFFARX1 I_51702 (I882507,I3563,I882230,I882533,);
not I_51703 (I882541,I882533);
nand I_51704 (I882558,I882541,I882454);
nand I_51705 (I882207,I882541,I882363);
nor I_51706 (I882589,I2364,I1380);
and I_51707 (I882606,I882454,I882589);
nor I_51708 (I882623,I882541,I882606);
DFFARX1 I_51709 (I882623,I3563,I882230,I882216,);
nor I_51710 (I882654,I882256,I882589);
DFFARX1 I_51711 (I882654,I3563,I882230,I882201,);
nor I_51712 (I882685,I882533,I882589);
not I_51713 (I882702,I882685);
nand I_51714 (I882210,I882702,I882558);
not I_51715 (I882757,I3570);
DFFARX1 I_51716 (I295914,I3563,I882757,I882783,);
not I_51717 (I882791,I882783);
nand I_51718 (I882808,I295905,I295905);
and I_51719 (I882825,I882808,I295923);
DFFARX1 I_51720 (I882825,I3563,I882757,I882851,);
DFFARX1 I_51721 (I882851,I3563,I882757,I882746,);
DFFARX1 I_51722 (I295926,I3563,I882757,I882882,);
nand I_51723 (I882890,I882882,I295908);
not I_51724 (I882907,I882890);
DFFARX1 I_51725 (I882907,I3563,I882757,I882933,);
not I_51726 (I882941,I882933);
nor I_51727 (I882749,I882791,I882941);
DFFARX1 I_51728 (I295920,I3563,I882757,I882981,);
nor I_51729 (I882740,I882981,I882851);
nor I_51730 (I882731,I882981,I882907);
nand I_51731 (I883017,I295932,I295911);
and I_51732 (I883034,I883017,I295917);
DFFARX1 I_51733 (I883034,I3563,I882757,I883060,);
not I_51734 (I883068,I883060);
nand I_51735 (I883085,I883068,I882981);
nand I_51736 (I882734,I883068,I882890);
nor I_51737 (I883116,I295929,I295911);
and I_51738 (I883133,I882981,I883116);
nor I_51739 (I883150,I883068,I883133);
DFFARX1 I_51740 (I883150,I3563,I882757,I882743,);
nor I_51741 (I883181,I882783,I883116);
DFFARX1 I_51742 (I883181,I3563,I882757,I882728,);
nor I_51743 (I883212,I883060,I883116);
not I_51744 (I883229,I883212);
nand I_51745 (I882737,I883229,I883085);
not I_51746 (I883284,I3570);
DFFARX1 I_51747 (I1299331,I3563,I883284,I883310,);
not I_51748 (I883318,I883310);
nand I_51749 (I883335,I1299313,I1299316);
and I_51750 (I883352,I883335,I1299328);
DFFARX1 I_51751 (I883352,I3563,I883284,I883378,);
DFFARX1 I_51752 (I883378,I3563,I883284,I883273,);
DFFARX1 I_51753 (I1299337,I3563,I883284,I883409,);
nand I_51754 (I883417,I883409,I1299322);
not I_51755 (I883434,I883417);
DFFARX1 I_51756 (I883434,I3563,I883284,I883460,);
not I_51757 (I883468,I883460);
nor I_51758 (I883276,I883318,I883468);
DFFARX1 I_51759 (I1299334,I3563,I883284,I883508,);
nor I_51760 (I883267,I883508,I883378);
nor I_51761 (I883258,I883508,I883434);
nand I_51762 (I883544,I1299325,I1299319);
and I_51763 (I883561,I883544,I1299313);
DFFARX1 I_51764 (I883561,I3563,I883284,I883587,);
not I_51765 (I883595,I883587);
nand I_51766 (I883612,I883595,I883508);
nand I_51767 (I883261,I883595,I883417);
nor I_51768 (I883643,I1299316,I1299319);
and I_51769 (I883660,I883508,I883643);
nor I_51770 (I883677,I883595,I883660);
DFFARX1 I_51771 (I883677,I3563,I883284,I883270,);
nor I_51772 (I883708,I883310,I883643);
DFFARX1 I_51773 (I883708,I3563,I883284,I883255,);
nor I_51774 (I883739,I883587,I883643);
not I_51775 (I883756,I883739);
nand I_51776 (I883264,I883756,I883612);
not I_51777 (I883811,I3570);
DFFARX1 I_51778 (I13108,I3563,I883811,I883837,);
not I_51779 (I883845,I883837);
nand I_51780 (I883862,I13114,I13096);
and I_51781 (I883879,I883862,I13105);
DFFARX1 I_51782 (I883879,I3563,I883811,I883905,);
DFFARX1 I_51783 (I883905,I3563,I883811,I883800,);
DFFARX1 I_51784 (I13096,I3563,I883811,I883936,);
nand I_51785 (I883944,I883936,I13099);
not I_51786 (I883961,I883944);
DFFARX1 I_51787 (I883961,I3563,I883811,I883987,);
not I_51788 (I883995,I883987);
nor I_51789 (I883803,I883845,I883995);
DFFARX1 I_51790 (I13099,I3563,I883811,I884035,);
nor I_51791 (I883794,I884035,I883905);
nor I_51792 (I883785,I884035,I883961);
nand I_51793 (I884071,I13102,I13111);
and I_51794 (I884088,I884071,I13093);
DFFARX1 I_51795 (I884088,I3563,I883811,I884114,);
not I_51796 (I884122,I884114);
nand I_51797 (I884139,I884122,I884035);
nand I_51798 (I883788,I884122,I883944);
nor I_51799 (I884170,I13093,I13111);
and I_51800 (I884187,I884035,I884170);
nor I_51801 (I884204,I884122,I884187);
DFFARX1 I_51802 (I884204,I3563,I883811,I883797,);
nor I_51803 (I884235,I883837,I884170);
DFFARX1 I_51804 (I884235,I3563,I883811,I883782,);
nor I_51805 (I884266,I884114,I884170);
not I_51806 (I884283,I884266);
nand I_51807 (I883791,I884283,I884139);
not I_51808 (I884338,I3570);
DFFARX1 I_51809 (I76697,I3563,I884338,I884364,);
not I_51810 (I884372,I884364);
nand I_51811 (I884389,I76673,I76682);
and I_51812 (I884406,I884389,I76676);
DFFARX1 I_51813 (I884406,I3563,I884338,I884432,);
DFFARX1 I_51814 (I884432,I3563,I884338,I884327,);
DFFARX1 I_51815 (I76694,I3563,I884338,I884463,);
nand I_51816 (I884471,I884463,I76685);
not I_51817 (I884488,I884471);
DFFARX1 I_51818 (I884488,I3563,I884338,I884514,);
not I_51819 (I884522,I884514);
nor I_51820 (I884330,I884372,I884522);
DFFARX1 I_51821 (I76679,I3563,I884338,I884562,);
nor I_51822 (I884321,I884562,I884432);
nor I_51823 (I884312,I884562,I884488);
nand I_51824 (I884598,I76691,I76688);
and I_51825 (I884615,I884598,I76676);
DFFARX1 I_51826 (I884615,I3563,I884338,I884641,);
not I_51827 (I884649,I884641);
nand I_51828 (I884666,I884649,I884562);
nand I_51829 (I884315,I884649,I884471);
nor I_51830 (I884697,I76673,I76688);
and I_51831 (I884714,I884562,I884697);
nor I_51832 (I884731,I884649,I884714);
DFFARX1 I_51833 (I884731,I3563,I884338,I884324,);
nor I_51834 (I884762,I884364,I884697);
DFFARX1 I_51835 (I884762,I3563,I884338,I884309,);
nor I_51836 (I884793,I884641,I884697);
not I_51837 (I884810,I884793);
nand I_51838 (I884318,I884810,I884666);
not I_51839 (I884865,I3570);
DFFARX1 I_51840 (I683267,I3563,I884865,I884891,);
not I_51841 (I884899,I884891);
nand I_51842 (I884916,I683270,I683267);
and I_51843 (I884933,I884916,I683279);
DFFARX1 I_51844 (I884933,I3563,I884865,I884959,);
DFFARX1 I_51845 (I884959,I3563,I884865,I884854,);
DFFARX1 I_51846 (I683276,I3563,I884865,I884990,);
nand I_51847 (I884998,I884990,I683282);
not I_51848 (I885015,I884998);
DFFARX1 I_51849 (I885015,I3563,I884865,I885041,);
not I_51850 (I885049,I885041);
nor I_51851 (I884857,I884899,I885049);
DFFARX1 I_51852 (I683291,I3563,I884865,I885089,);
nor I_51853 (I884848,I885089,I884959);
nor I_51854 (I884839,I885089,I885015);
nand I_51855 (I885125,I683285,I683273);
and I_51856 (I885142,I885125,I683270);
DFFARX1 I_51857 (I885142,I3563,I884865,I885168,);
not I_51858 (I885176,I885168);
nand I_51859 (I885193,I885176,I885089);
nand I_51860 (I884842,I885176,I884998);
nor I_51861 (I885224,I683288,I683273);
and I_51862 (I885241,I885089,I885224);
nor I_51863 (I885258,I885176,I885241);
DFFARX1 I_51864 (I885258,I3563,I884865,I884851,);
nor I_51865 (I885289,I884891,I885224);
DFFARX1 I_51866 (I885289,I3563,I884865,I884836,);
nor I_51867 (I885320,I885168,I885224);
not I_51868 (I885337,I885320);
nand I_51869 (I884845,I885337,I885193);
not I_51870 (I885392,I3570);
DFFARX1 I_51871 (I214294,I3563,I885392,I885418,);
not I_51872 (I885426,I885418);
nand I_51873 (I885443,I214291,I214309);
and I_51874 (I885460,I885443,I214300);
DFFARX1 I_51875 (I885460,I3563,I885392,I885486,);
DFFARX1 I_51876 (I885486,I3563,I885392,I885381,);
DFFARX1 I_51877 (I214306,I3563,I885392,I885517,);
nand I_51878 (I885525,I885517,I214303);
not I_51879 (I885542,I885525);
DFFARX1 I_51880 (I885542,I3563,I885392,I885568,);
not I_51881 (I885576,I885568);
nor I_51882 (I885384,I885426,I885576);
DFFARX1 I_51883 (I214297,I3563,I885392,I885616,);
nor I_51884 (I885375,I885616,I885486);
nor I_51885 (I885366,I885616,I885542);
nand I_51886 (I885652,I214288,I214312);
and I_51887 (I885669,I885652,I214291);
DFFARX1 I_51888 (I885669,I3563,I885392,I885695,);
not I_51889 (I885703,I885695);
nand I_51890 (I885720,I885703,I885616);
nand I_51891 (I885369,I885703,I885525);
nor I_51892 (I885751,I214288,I214312);
and I_51893 (I885768,I885616,I885751);
nor I_51894 (I885785,I885703,I885768);
DFFARX1 I_51895 (I885785,I3563,I885392,I885378,);
nor I_51896 (I885816,I885418,I885751);
DFFARX1 I_51897 (I885816,I3563,I885392,I885363,);
nor I_51898 (I885847,I885695,I885751);
not I_51899 (I885864,I885847);
nand I_51900 (I885372,I885864,I885720);
not I_51901 (I885919,I3570);
DFFARX1 I_51902 (I393936,I3563,I885919,I885945,);
not I_51903 (I885953,I885945);
nand I_51904 (I885970,I393927,I393927);
and I_51905 (I885987,I885970,I393945);
DFFARX1 I_51906 (I885987,I3563,I885919,I886013,);
DFFARX1 I_51907 (I886013,I3563,I885919,I885908,);
DFFARX1 I_51908 (I393948,I3563,I885919,I886044,);
nand I_51909 (I886052,I886044,I393930);
not I_51910 (I886069,I886052);
DFFARX1 I_51911 (I886069,I3563,I885919,I886095,);
not I_51912 (I886103,I886095);
nor I_51913 (I885911,I885953,I886103);
DFFARX1 I_51914 (I393942,I3563,I885919,I886143,);
nor I_51915 (I885902,I886143,I886013);
nor I_51916 (I885893,I886143,I886069);
nand I_51917 (I886179,I393954,I393933);
and I_51918 (I886196,I886179,I393939);
DFFARX1 I_51919 (I886196,I3563,I885919,I886222,);
not I_51920 (I886230,I886222);
nand I_51921 (I886247,I886230,I886143);
nand I_51922 (I885896,I886230,I886052);
nor I_51923 (I886278,I393951,I393933);
and I_51924 (I886295,I886143,I886278);
nor I_51925 (I886312,I886230,I886295);
DFFARX1 I_51926 (I886312,I3563,I885919,I885905,);
nor I_51927 (I886343,I885945,I886278);
DFFARX1 I_51928 (I886343,I3563,I885919,I885890,);
nor I_51929 (I886374,I886222,I886278);
not I_51930 (I886391,I886374);
nand I_51931 (I885899,I886391,I886247);
not I_51932 (I886446,I3570);
DFFARX1 I_51933 (I266654,I3563,I886446,I886472,);
not I_51934 (I886480,I886472);
nand I_51935 (I886497,I266651,I266669);
and I_51936 (I886514,I886497,I266660);
DFFARX1 I_51937 (I886514,I3563,I886446,I886540,);
DFFARX1 I_51938 (I886540,I3563,I886446,I886435,);
DFFARX1 I_51939 (I266666,I3563,I886446,I886571,);
nand I_51940 (I886579,I886571,I266663);
not I_51941 (I886596,I886579);
DFFARX1 I_51942 (I886596,I3563,I886446,I886622,);
not I_51943 (I886630,I886622);
nor I_51944 (I886438,I886480,I886630);
DFFARX1 I_51945 (I266657,I3563,I886446,I886670,);
nor I_51946 (I886429,I886670,I886540);
nor I_51947 (I886420,I886670,I886596);
nand I_51948 (I886706,I266648,I266672);
and I_51949 (I886723,I886706,I266651);
DFFARX1 I_51950 (I886723,I3563,I886446,I886749,);
not I_51951 (I886757,I886749);
nand I_51952 (I886774,I886757,I886670);
nand I_51953 (I886423,I886757,I886579);
nor I_51954 (I886805,I266648,I266672);
and I_51955 (I886822,I886670,I886805);
nor I_51956 (I886839,I886757,I886822);
DFFARX1 I_51957 (I886839,I3563,I886446,I886432,);
nor I_51958 (I886870,I886472,I886805);
DFFARX1 I_51959 (I886870,I3563,I886446,I886417,);
nor I_51960 (I886901,I886749,I886805);
not I_51961 (I886918,I886901);
nand I_51962 (I886426,I886918,I886774);
not I_51963 (I886973,I3570);
DFFARX1 I_51964 (I717369,I3563,I886973,I886999,);
not I_51965 (I887007,I886999);
nand I_51966 (I887024,I717372,I717369);
and I_51967 (I887041,I887024,I717381);
DFFARX1 I_51968 (I887041,I3563,I886973,I887067,);
DFFARX1 I_51969 (I887067,I3563,I886973,I886962,);
DFFARX1 I_51970 (I717378,I3563,I886973,I887098,);
nand I_51971 (I887106,I887098,I717384);
not I_51972 (I887123,I887106);
DFFARX1 I_51973 (I887123,I3563,I886973,I887149,);
not I_51974 (I887157,I887149);
nor I_51975 (I886965,I887007,I887157);
DFFARX1 I_51976 (I717393,I3563,I886973,I887197,);
nor I_51977 (I886956,I887197,I887067);
nor I_51978 (I886947,I887197,I887123);
nand I_51979 (I887233,I717387,I717375);
and I_51980 (I887250,I887233,I717372);
DFFARX1 I_51981 (I887250,I3563,I886973,I887276,);
not I_51982 (I887284,I887276);
nand I_51983 (I887301,I887284,I887197);
nand I_51984 (I886950,I887284,I887106);
nor I_51985 (I887332,I717390,I717375);
and I_51986 (I887349,I887197,I887332);
nor I_51987 (I887366,I887284,I887349);
DFFARX1 I_51988 (I887366,I3563,I886973,I886959,);
nor I_51989 (I887397,I886999,I887332);
DFFARX1 I_51990 (I887397,I3563,I886973,I886944,);
nor I_51991 (I887428,I887276,I887332);
not I_51992 (I887445,I887428);
nand I_51993 (I886953,I887445,I887301);
not I_51994 (I887500,I3570);
DFFARX1 I_51995 (I28725,I3563,I887500,I887526,);
not I_51996 (I887534,I887526);
nand I_51997 (I887551,I28737,I28740);
and I_51998 (I887568,I887551,I28716);
DFFARX1 I_51999 (I887568,I3563,I887500,I887594,);
DFFARX1 I_52000 (I887594,I3563,I887500,I887489,);
DFFARX1 I_52001 (I28734,I3563,I887500,I887625,);
nand I_52002 (I887633,I887625,I28722);
not I_52003 (I887650,I887633);
DFFARX1 I_52004 (I887650,I3563,I887500,I887676,);
not I_52005 (I887684,I887676);
nor I_52006 (I887492,I887534,I887684);
DFFARX1 I_52007 (I28719,I3563,I887500,I887724,);
nor I_52008 (I887483,I887724,I887594);
nor I_52009 (I887474,I887724,I887650);
nand I_52010 (I887760,I28728,I28719);
and I_52011 (I887777,I887760,I28716);
DFFARX1 I_52012 (I887777,I3563,I887500,I887803,);
not I_52013 (I887811,I887803);
nand I_52014 (I887828,I887811,I887724);
nand I_52015 (I887477,I887811,I887633);
nor I_52016 (I887859,I28731,I28719);
and I_52017 (I887876,I887724,I887859);
nor I_52018 (I887893,I887811,I887876);
DFFARX1 I_52019 (I887893,I3563,I887500,I887486,);
nor I_52020 (I887924,I887526,I887859);
DFFARX1 I_52021 (I887924,I3563,I887500,I887471,);
nor I_52022 (I887955,I887803,I887859);
not I_52023 (I887972,I887955);
nand I_52024 (I887480,I887972,I887828);
not I_52025 (I888027,I3570);
DFFARX1 I_52026 (I144680,I3563,I888027,I888053,);
not I_52027 (I888061,I888053);
nand I_52028 (I888078,I144656,I144665);
and I_52029 (I888095,I888078,I144659);
DFFARX1 I_52030 (I888095,I3563,I888027,I888121,);
DFFARX1 I_52031 (I888121,I3563,I888027,I888016,);
DFFARX1 I_52032 (I144677,I3563,I888027,I888152,);
nand I_52033 (I888160,I888152,I144668);
not I_52034 (I888177,I888160);
DFFARX1 I_52035 (I888177,I3563,I888027,I888203,);
not I_52036 (I888211,I888203);
nor I_52037 (I888019,I888061,I888211);
DFFARX1 I_52038 (I144662,I3563,I888027,I888251,);
nor I_52039 (I888010,I888251,I888121);
nor I_52040 (I888001,I888251,I888177);
nand I_52041 (I888287,I144674,I144671);
and I_52042 (I888304,I888287,I144659);
DFFARX1 I_52043 (I888304,I3563,I888027,I888330,);
not I_52044 (I888338,I888330);
nand I_52045 (I888355,I888338,I888251);
nand I_52046 (I888004,I888338,I888160);
nor I_52047 (I888386,I144656,I144671);
and I_52048 (I888403,I888251,I888386);
nor I_52049 (I888420,I888338,I888403);
DFFARX1 I_52050 (I888420,I3563,I888027,I888013,);
nor I_52051 (I888451,I888053,I888386);
DFFARX1 I_52052 (I888451,I3563,I888027,I887998,);
nor I_52053 (I888482,I888330,I888386);
not I_52054 (I888499,I888482);
nand I_52055 (I888007,I888499,I888355);
not I_52056 (I888554,I3570);
DFFARX1 I_52057 (I758407,I3563,I888554,I888580,);
not I_52058 (I888588,I888580);
nand I_52059 (I888605,I758410,I758407);
and I_52060 (I888622,I888605,I758419);
DFFARX1 I_52061 (I888622,I3563,I888554,I888648,);
DFFARX1 I_52062 (I888648,I3563,I888554,I888543,);
DFFARX1 I_52063 (I758416,I3563,I888554,I888679,);
nand I_52064 (I888687,I888679,I758422);
not I_52065 (I888704,I888687);
DFFARX1 I_52066 (I888704,I3563,I888554,I888730,);
not I_52067 (I888738,I888730);
nor I_52068 (I888546,I888588,I888738);
DFFARX1 I_52069 (I758431,I3563,I888554,I888778,);
nor I_52070 (I888537,I888778,I888648);
nor I_52071 (I888528,I888778,I888704);
nand I_52072 (I888814,I758425,I758413);
and I_52073 (I888831,I888814,I758410);
DFFARX1 I_52074 (I888831,I3563,I888554,I888857,);
not I_52075 (I888865,I888857);
nand I_52076 (I888882,I888865,I888778);
nand I_52077 (I888531,I888865,I888687);
nor I_52078 (I888913,I758428,I758413);
and I_52079 (I888930,I888778,I888913);
nor I_52080 (I888947,I888865,I888930);
DFFARX1 I_52081 (I888947,I3563,I888554,I888540,);
nor I_52082 (I888978,I888580,I888913);
DFFARX1 I_52083 (I888978,I3563,I888554,I888525,);
nor I_52084 (I889009,I888857,I888913);
not I_52085 (I889026,I889009);
nand I_52086 (I888534,I889026,I888882);
not I_52087 (I889081,I3570);
DFFARX1 I_52088 (I465928,I3563,I889081,I889107,);
not I_52089 (I889115,I889107);
nand I_52090 (I889132,I465925,I465934);
and I_52091 (I889149,I889132,I465943);
DFFARX1 I_52092 (I889149,I3563,I889081,I889175,);
DFFARX1 I_52093 (I889175,I3563,I889081,I889070,);
DFFARX1 I_52094 (I465946,I3563,I889081,I889206,);
nand I_52095 (I889214,I889206,I465949);
not I_52096 (I889231,I889214);
DFFARX1 I_52097 (I889231,I3563,I889081,I889257,);
not I_52098 (I889265,I889257);
nor I_52099 (I889073,I889115,I889265);
DFFARX1 I_52100 (I465922,I3563,I889081,I889305,);
nor I_52101 (I889064,I889305,I889175);
nor I_52102 (I889055,I889305,I889231);
nand I_52103 (I889341,I465937,I465940);
and I_52104 (I889358,I889341,I465931);
DFFARX1 I_52105 (I889358,I3563,I889081,I889384,);
not I_52106 (I889392,I889384);
nand I_52107 (I889409,I889392,I889305);
nand I_52108 (I889058,I889392,I889214);
nor I_52109 (I889440,I465922,I465940);
and I_52110 (I889457,I889305,I889440);
nor I_52111 (I889474,I889392,I889457);
DFFARX1 I_52112 (I889474,I3563,I889081,I889067,);
nor I_52113 (I889505,I889107,I889440);
DFFARX1 I_52114 (I889505,I3563,I889081,I889052,);
nor I_52115 (I889536,I889384,I889440);
not I_52116 (I889553,I889536);
nand I_52117 (I889061,I889553,I889409);
not I_52118 (I889608,I3570);
DFFARX1 I_52119 (I238689,I3563,I889608,I889634,);
not I_52120 (I889642,I889634);
nand I_52121 (I889659,I238686,I238704);
and I_52122 (I889676,I889659,I238695);
DFFARX1 I_52123 (I889676,I3563,I889608,I889702,);
DFFARX1 I_52124 (I889702,I3563,I889608,I889597,);
DFFARX1 I_52125 (I238701,I3563,I889608,I889733,);
nand I_52126 (I889741,I889733,I238698);
not I_52127 (I889758,I889741);
DFFARX1 I_52128 (I889758,I3563,I889608,I889784,);
not I_52129 (I889792,I889784);
nor I_52130 (I889600,I889642,I889792);
DFFARX1 I_52131 (I238692,I3563,I889608,I889832,);
nor I_52132 (I889591,I889832,I889702);
nor I_52133 (I889582,I889832,I889758);
nand I_52134 (I889868,I238683,I238707);
and I_52135 (I889885,I889868,I238686);
DFFARX1 I_52136 (I889885,I3563,I889608,I889911,);
not I_52137 (I889919,I889911);
nand I_52138 (I889936,I889919,I889832);
nand I_52139 (I889585,I889919,I889741);
nor I_52140 (I889967,I238683,I238707);
and I_52141 (I889984,I889832,I889967);
nor I_52142 (I890001,I889919,I889984);
DFFARX1 I_52143 (I890001,I3563,I889608,I889594,);
nor I_52144 (I890032,I889634,I889967);
DFFARX1 I_52145 (I890032,I3563,I889608,I889579,);
nor I_52146 (I890063,I889911,I889967);
not I_52147 (I890080,I890063);
nand I_52148 (I889588,I890080,I889936);
not I_52149 (I890135,I3570);
DFFARX1 I_52150 (I431656,I3563,I890135,I890161,);
not I_52151 (I890169,I890161);
nand I_52152 (I890186,I431653,I431662);
and I_52153 (I890203,I890186,I431671);
DFFARX1 I_52154 (I890203,I3563,I890135,I890229,);
DFFARX1 I_52155 (I890229,I3563,I890135,I890124,);
DFFARX1 I_52156 (I431674,I3563,I890135,I890260,);
nand I_52157 (I890268,I890260,I431677);
not I_52158 (I890285,I890268);
DFFARX1 I_52159 (I890285,I3563,I890135,I890311,);
not I_52160 (I890319,I890311);
nor I_52161 (I890127,I890169,I890319);
DFFARX1 I_52162 (I431650,I3563,I890135,I890359,);
nor I_52163 (I890118,I890359,I890229);
nor I_52164 (I890109,I890359,I890285);
nand I_52165 (I890395,I431665,I431668);
and I_52166 (I890412,I890395,I431659);
DFFARX1 I_52167 (I890412,I3563,I890135,I890438,);
not I_52168 (I890446,I890438);
nand I_52169 (I890463,I890446,I890359);
nand I_52170 (I890112,I890446,I890268);
nor I_52171 (I890494,I431650,I431668);
and I_52172 (I890511,I890359,I890494);
nor I_52173 (I890528,I890446,I890511);
DFFARX1 I_52174 (I890528,I3563,I890135,I890121,);
nor I_52175 (I890559,I890161,I890494);
DFFARX1 I_52176 (I890559,I3563,I890135,I890106,);
nor I_52177 (I890590,I890438,I890494);
not I_52178 (I890607,I890590);
nand I_52179 (I890115,I890607,I890463);
not I_52180 (I890662,I3570);
DFFARX1 I_52181 (I147315,I3563,I890662,I890688,);
not I_52182 (I890696,I890688);
nand I_52183 (I890713,I147291,I147300);
and I_52184 (I890730,I890713,I147294);
DFFARX1 I_52185 (I890730,I3563,I890662,I890756,);
DFFARX1 I_52186 (I890756,I3563,I890662,I890651,);
DFFARX1 I_52187 (I147312,I3563,I890662,I890787,);
nand I_52188 (I890795,I890787,I147303);
not I_52189 (I890812,I890795);
DFFARX1 I_52190 (I890812,I3563,I890662,I890838,);
not I_52191 (I890846,I890838);
nor I_52192 (I890654,I890696,I890846);
DFFARX1 I_52193 (I147297,I3563,I890662,I890886,);
nor I_52194 (I890645,I890886,I890756);
nor I_52195 (I890636,I890886,I890812);
nand I_52196 (I890922,I147309,I147306);
and I_52197 (I890939,I890922,I147294);
DFFARX1 I_52198 (I890939,I3563,I890662,I890965,);
not I_52199 (I890973,I890965);
nand I_52200 (I890990,I890973,I890886);
nand I_52201 (I890639,I890973,I890795);
nor I_52202 (I891021,I147291,I147306);
and I_52203 (I891038,I890886,I891021);
nor I_52204 (I891055,I890973,I891038);
DFFARX1 I_52205 (I891055,I3563,I890662,I890648,);
nor I_52206 (I891086,I890688,I891021);
DFFARX1 I_52207 (I891086,I3563,I890662,I890633,);
nor I_52208 (I891117,I890965,I891021);
not I_52209 (I891134,I891117);
nand I_52210 (I890642,I891134,I890990);
not I_52211 (I891189,I3570);
DFFARX1 I_52212 (I480616,I3563,I891189,I891215,);
not I_52213 (I891223,I891215);
nand I_52214 (I891240,I480613,I480622);
and I_52215 (I891257,I891240,I480631);
DFFARX1 I_52216 (I891257,I3563,I891189,I891283,);
DFFARX1 I_52217 (I891283,I3563,I891189,I891178,);
DFFARX1 I_52218 (I480634,I3563,I891189,I891314,);
nand I_52219 (I891322,I891314,I480637);
not I_52220 (I891339,I891322);
DFFARX1 I_52221 (I891339,I3563,I891189,I891365,);
not I_52222 (I891373,I891365);
nor I_52223 (I891181,I891223,I891373);
DFFARX1 I_52224 (I480610,I3563,I891189,I891413,);
nor I_52225 (I891172,I891413,I891283);
nor I_52226 (I891163,I891413,I891339);
nand I_52227 (I891449,I480625,I480628);
and I_52228 (I891466,I891449,I480619);
DFFARX1 I_52229 (I891466,I3563,I891189,I891492,);
not I_52230 (I891500,I891492);
nand I_52231 (I891517,I891500,I891413);
nand I_52232 (I891166,I891500,I891322);
nor I_52233 (I891548,I480610,I480628);
and I_52234 (I891565,I891413,I891548);
nor I_52235 (I891582,I891500,I891565);
DFFARX1 I_52236 (I891582,I3563,I891189,I891175,);
nor I_52237 (I891613,I891215,I891548);
DFFARX1 I_52238 (I891613,I3563,I891189,I891160,);
nor I_52239 (I891644,I891492,I891548);
not I_52240 (I891661,I891644);
nand I_52241 (I891169,I891661,I891517);
not I_52242 (I891716,I3570);
DFFARX1 I_52243 (I1035680,I3563,I891716,I891742,);
not I_52244 (I891750,I891742);
nand I_52245 (I891767,I1035695,I1035677);
and I_52246 (I891784,I891767,I1035677);
DFFARX1 I_52247 (I891784,I3563,I891716,I891810,);
DFFARX1 I_52248 (I891810,I3563,I891716,I891705,);
DFFARX1 I_52249 (I1035686,I3563,I891716,I891841,);
nand I_52250 (I891849,I891841,I1035704);
not I_52251 (I891866,I891849);
DFFARX1 I_52252 (I891866,I3563,I891716,I891892,);
not I_52253 (I891900,I891892);
nor I_52254 (I891708,I891750,I891900);
DFFARX1 I_52255 (I1035701,I3563,I891716,I891940,);
nor I_52256 (I891699,I891940,I891810);
nor I_52257 (I891690,I891940,I891866);
nand I_52258 (I891976,I1035698,I1035689);
and I_52259 (I891993,I891976,I1035683);
DFFARX1 I_52260 (I891993,I3563,I891716,I892019,);
not I_52261 (I892027,I892019);
nand I_52262 (I892044,I892027,I891940);
nand I_52263 (I891693,I892027,I891849);
nor I_52264 (I892075,I1035692,I1035689);
and I_52265 (I892092,I891940,I892075);
nor I_52266 (I892109,I892027,I892092);
DFFARX1 I_52267 (I892109,I3563,I891716,I891702,);
nor I_52268 (I892140,I891742,I892075);
DFFARX1 I_52269 (I892140,I3563,I891716,I891687,);
nor I_52270 (I892171,I892019,I892075);
not I_52271 (I892188,I892171);
nand I_52272 (I891696,I892188,I892044);
not I_52273 (I892243,I3570);
DFFARX1 I_52274 (I797711,I3563,I892243,I892269,);
not I_52275 (I892277,I892269);
nand I_52276 (I892294,I797714,I797711);
and I_52277 (I892311,I892294,I797723);
DFFARX1 I_52278 (I892311,I3563,I892243,I892337,);
DFFARX1 I_52279 (I892337,I3563,I892243,I892232,);
DFFARX1 I_52280 (I797720,I3563,I892243,I892368,);
nand I_52281 (I892376,I892368,I797726);
not I_52282 (I892393,I892376);
DFFARX1 I_52283 (I892393,I3563,I892243,I892419,);
not I_52284 (I892427,I892419);
nor I_52285 (I892235,I892277,I892427);
DFFARX1 I_52286 (I797735,I3563,I892243,I892467,);
nor I_52287 (I892226,I892467,I892337);
nor I_52288 (I892217,I892467,I892393);
nand I_52289 (I892503,I797729,I797717);
and I_52290 (I892520,I892503,I797714);
DFFARX1 I_52291 (I892520,I3563,I892243,I892546,);
not I_52292 (I892554,I892546);
nand I_52293 (I892571,I892554,I892467);
nand I_52294 (I892220,I892554,I892376);
nor I_52295 (I892602,I797732,I797717);
and I_52296 (I892619,I892467,I892602);
nor I_52297 (I892636,I892554,I892619);
DFFARX1 I_52298 (I892636,I3563,I892243,I892229,);
nor I_52299 (I892667,I892269,I892602);
DFFARX1 I_52300 (I892667,I3563,I892243,I892214,);
nor I_52301 (I892698,I892546,I892602);
not I_52302 (I892715,I892698);
nand I_52303 (I892223,I892715,I892571);
not I_52304 (I892770,I3570);
DFFARX1 I_52305 (I21347,I3563,I892770,I892796,);
not I_52306 (I892804,I892796);
nand I_52307 (I892821,I21359,I21362);
and I_52308 (I892838,I892821,I21338);
DFFARX1 I_52309 (I892838,I3563,I892770,I892864,);
DFFARX1 I_52310 (I892864,I3563,I892770,I892759,);
DFFARX1 I_52311 (I21356,I3563,I892770,I892895,);
nand I_52312 (I892903,I892895,I21344);
not I_52313 (I892920,I892903);
DFFARX1 I_52314 (I892920,I3563,I892770,I892946,);
not I_52315 (I892954,I892946);
nor I_52316 (I892762,I892804,I892954);
DFFARX1 I_52317 (I21341,I3563,I892770,I892994,);
nor I_52318 (I892753,I892994,I892864);
nor I_52319 (I892744,I892994,I892920);
nand I_52320 (I893030,I21350,I21341);
and I_52321 (I893047,I893030,I21338);
DFFARX1 I_52322 (I893047,I3563,I892770,I893073,);
not I_52323 (I893081,I893073);
nand I_52324 (I893098,I893081,I892994);
nand I_52325 (I892747,I893081,I892903);
nor I_52326 (I893129,I21353,I21341);
and I_52327 (I893146,I892994,I893129);
nor I_52328 (I893163,I893081,I893146);
DFFARX1 I_52329 (I893163,I3563,I892770,I892756,);
nor I_52330 (I893194,I892796,I893129);
DFFARX1 I_52331 (I893194,I3563,I892770,I892741,);
nor I_52332 (I893225,I893073,I893129);
not I_52333 (I893242,I893225);
nand I_52334 (I892750,I893242,I893098);
not I_52335 (I893297,I3570);
DFFARX1 I_52336 (I1140143,I3563,I893297,I893323,);
not I_52337 (I893331,I893323);
nand I_52338 (I893348,I1140125,I1140125);
and I_52339 (I893365,I893348,I1140131);
DFFARX1 I_52340 (I893365,I3563,I893297,I893391,);
DFFARX1 I_52341 (I893391,I3563,I893297,I893286,);
DFFARX1 I_52342 (I1140128,I3563,I893297,I893422,);
nand I_52343 (I893430,I893422,I1140137);
not I_52344 (I893447,I893430);
DFFARX1 I_52345 (I893447,I3563,I893297,I893473,);
not I_52346 (I893481,I893473);
nor I_52347 (I893289,I893331,I893481);
DFFARX1 I_52348 (I1140149,I3563,I893297,I893521,);
nor I_52349 (I893280,I893521,I893391);
nor I_52350 (I893271,I893521,I893447);
nand I_52351 (I893557,I1140140,I1140134);
and I_52352 (I893574,I893557,I1140128);
DFFARX1 I_52353 (I893574,I3563,I893297,I893600,);
not I_52354 (I893608,I893600);
nand I_52355 (I893625,I893608,I893521);
nand I_52356 (I893274,I893608,I893430);
nor I_52357 (I893656,I1140146,I1140134);
and I_52358 (I893673,I893521,I893656);
nor I_52359 (I893690,I893608,I893673);
DFFARX1 I_52360 (I893690,I3563,I893297,I893283,);
nor I_52361 (I893721,I893323,I893656);
DFFARX1 I_52362 (I893721,I3563,I893297,I893268,);
nor I_52363 (I893752,I893600,I893656);
not I_52364 (I893769,I893752);
nand I_52365 (I893277,I893769,I893625);
not I_52366 (I893824,I3570);
DFFARX1 I_52367 (I1227999,I3563,I893824,I893850,);
not I_52368 (I893858,I893850);
nand I_52369 (I893875,I1227981,I1227981);
and I_52370 (I893892,I893875,I1227987);
DFFARX1 I_52371 (I893892,I3563,I893824,I893918,);
DFFARX1 I_52372 (I893918,I3563,I893824,I893813,);
DFFARX1 I_52373 (I1227984,I3563,I893824,I893949,);
nand I_52374 (I893957,I893949,I1227993);
not I_52375 (I893974,I893957);
DFFARX1 I_52376 (I893974,I3563,I893824,I894000,);
not I_52377 (I894008,I894000);
nor I_52378 (I893816,I893858,I894008);
DFFARX1 I_52379 (I1228005,I3563,I893824,I894048,);
nor I_52380 (I893807,I894048,I893918);
nor I_52381 (I893798,I894048,I893974);
nand I_52382 (I894084,I1227996,I1227990);
and I_52383 (I894101,I894084,I1227984);
DFFARX1 I_52384 (I894101,I3563,I893824,I894127,);
not I_52385 (I894135,I894127);
nand I_52386 (I894152,I894135,I894048);
nand I_52387 (I893801,I894135,I893957);
nor I_52388 (I894183,I1228002,I1227990);
and I_52389 (I894200,I894048,I894183);
nor I_52390 (I894217,I894135,I894200);
DFFARX1 I_52391 (I894217,I3563,I893824,I893810,);
nor I_52392 (I894248,I893850,I894183);
DFFARX1 I_52393 (I894248,I3563,I893824,I893795,);
nor I_52394 (I894279,I894127,I894183);
not I_52395 (I894296,I894279);
nand I_52396 (I893804,I894296,I894152);
not I_52397 (I894351,I3570);
DFFARX1 I_52398 (I775169,I3563,I894351,I894377,);
not I_52399 (I894385,I894377);
nand I_52400 (I894402,I775172,I775169);
and I_52401 (I894419,I894402,I775181);
DFFARX1 I_52402 (I894419,I3563,I894351,I894445,);
DFFARX1 I_52403 (I894445,I3563,I894351,I894340,);
DFFARX1 I_52404 (I775178,I3563,I894351,I894476,);
nand I_52405 (I894484,I894476,I775184);
not I_52406 (I894501,I894484);
DFFARX1 I_52407 (I894501,I3563,I894351,I894527,);
not I_52408 (I894535,I894527);
nor I_52409 (I894343,I894385,I894535);
DFFARX1 I_52410 (I775193,I3563,I894351,I894575,);
nor I_52411 (I894334,I894575,I894445);
nor I_52412 (I894325,I894575,I894501);
nand I_52413 (I894611,I775187,I775175);
and I_52414 (I894628,I894611,I775172);
DFFARX1 I_52415 (I894628,I3563,I894351,I894654,);
not I_52416 (I894662,I894654);
nand I_52417 (I894679,I894662,I894575);
nand I_52418 (I894328,I894662,I894484);
nor I_52419 (I894710,I775190,I775175);
and I_52420 (I894727,I894575,I894710);
nor I_52421 (I894744,I894662,I894727);
DFFARX1 I_52422 (I894744,I3563,I894351,I894337,);
nor I_52423 (I894775,I894377,I894710);
DFFARX1 I_52424 (I894775,I3563,I894351,I894322,);
nor I_52425 (I894806,I894654,I894710);
not I_52426 (I894823,I894806);
nand I_52427 (I894331,I894823,I894679);
not I_52428 (I894878,I3570);
DFFARX1 I_52429 (I63522,I3563,I894878,I894904,);
not I_52430 (I894912,I894904);
nand I_52431 (I894929,I63498,I63507);
and I_52432 (I894946,I894929,I63501);
DFFARX1 I_52433 (I894946,I3563,I894878,I894972,);
DFFARX1 I_52434 (I894972,I3563,I894878,I894867,);
DFFARX1 I_52435 (I63519,I3563,I894878,I895003,);
nand I_52436 (I895011,I895003,I63510);
not I_52437 (I895028,I895011);
DFFARX1 I_52438 (I895028,I3563,I894878,I895054,);
not I_52439 (I895062,I895054);
nor I_52440 (I894870,I894912,I895062);
DFFARX1 I_52441 (I63504,I3563,I894878,I895102,);
nor I_52442 (I894861,I895102,I894972);
nor I_52443 (I894852,I895102,I895028);
nand I_52444 (I895138,I63516,I63513);
and I_52445 (I895155,I895138,I63501);
DFFARX1 I_52446 (I895155,I3563,I894878,I895181,);
not I_52447 (I895189,I895181);
nand I_52448 (I895206,I895189,I895102);
nand I_52449 (I894855,I895189,I895011);
nor I_52450 (I895237,I63498,I63513);
and I_52451 (I895254,I895102,I895237);
nor I_52452 (I895271,I895189,I895254);
DFFARX1 I_52453 (I895271,I3563,I894878,I894864,);
nor I_52454 (I895302,I894904,I895237);
DFFARX1 I_52455 (I895302,I3563,I894878,I894849,);
nor I_52456 (I895333,I895181,I895237);
not I_52457 (I895350,I895333);
nand I_52458 (I894858,I895350,I895206);
not I_52459 (I895405,I3570);
DFFARX1 I_52460 (I432744,I3563,I895405,I895431,);
not I_52461 (I895439,I895431);
nand I_52462 (I895456,I432741,I432750);
and I_52463 (I895473,I895456,I432759);
DFFARX1 I_52464 (I895473,I3563,I895405,I895499,);
DFFARX1 I_52465 (I895499,I3563,I895405,I895394,);
DFFARX1 I_52466 (I432762,I3563,I895405,I895530,);
nand I_52467 (I895538,I895530,I432765);
not I_52468 (I895555,I895538);
DFFARX1 I_52469 (I895555,I3563,I895405,I895581,);
not I_52470 (I895589,I895581);
nor I_52471 (I895397,I895439,I895589);
DFFARX1 I_52472 (I432738,I3563,I895405,I895629,);
nor I_52473 (I895388,I895629,I895499);
nor I_52474 (I895379,I895629,I895555);
nand I_52475 (I895665,I432753,I432756);
and I_52476 (I895682,I895665,I432747);
DFFARX1 I_52477 (I895682,I3563,I895405,I895708,);
not I_52478 (I895716,I895708);
nand I_52479 (I895733,I895716,I895629);
nand I_52480 (I895382,I895716,I895538);
nor I_52481 (I895764,I432738,I432756);
and I_52482 (I895781,I895629,I895764);
nor I_52483 (I895798,I895716,I895781);
DFFARX1 I_52484 (I895798,I3563,I895405,I895391,);
nor I_52485 (I895829,I895431,I895764);
DFFARX1 I_52486 (I895829,I3563,I895405,I895376,);
nor I_52487 (I895860,I895708,I895764);
not I_52488 (I895877,I895860);
nand I_52489 (I895385,I895877,I895733);
not I_52490 (I895932,I3570);
DFFARX1 I_52491 (I294860,I3563,I895932,I895958,);
not I_52492 (I895966,I895958);
nand I_52493 (I895983,I294851,I294851);
and I_52494 (I896000,I895983,I294869);
DFFARX1 I_52495 (I896000,I3563,I895932,I896026,);
DFFARX1 I_52496 (I896026,I3563,I895932,I895921,);
DFFARX1 I_52497 (I294872,I3563,I895932,I896057,);
nand I_52498 (I896065,I896057,I294854);
not I_52499 (I896082,I896065);
DFFARX1 I_52500 (I896082,I3563,I895932,I896108,);
not I_52501 (I896116,I896108);
nor I_52502 (I895924,I895966,I896116);
DFFARX1 I_52503 (I294866,I3563,I895932,I896156,);
nor I_52504 (I895915,I896156,I896026);
nor I_52505 (I895906,I896156,I896082);
nand I_52506 (I896192,I294878,I294857);
and I_52507 (I896209,I896192,I294863);
DFFARX1 I_52508 (I896209,I3563,I895932,I896235,);
not I_52509 (I896243,I896235);
nand I_52510 (I896260,I896243,I896156);
nand I_52511 (I895909,I896243,I896065);
nor I_52512 (I896291,I294875,I294857);
and I_52513 (I896308,I896156,I896291);
nor I_52514 (I896325,I896243,I896308);
DFFARX1 I_52515 (I896325,I3563,I895932,I895918,);
nor I_52516 (I896356,I895958,I896291);
DFFARX1 I_52517 (I896356,I3563,I895932,I895903,);
nor I_52518 (I896387,I896235,I896291);
not I_52519 (I896404,I896387);
nand I_52520 (I895912,I896404,I896260);
not I_52521 (I896459,I3570);
DFFARX1 I_52522 (I990460,I3563,I896459,I896485,);
not I_52523 (I896493,I896485);
nand I_52524 (I896510,I990475,I990457);
and I_52525 (I896527,I896510,I990457);
DFFARX1 I_52526 (I896527,I3563,I896459,I896553,);
DFFARX1 I_52527 (I896553,I3563,I896459,I896448,);
DFFARX1 I_52528 (I990466,I3563,I896459,I896584,);
nand I_52529 (I896592,I896584,I990484);
not I_52530 (I896609,I896592);
DFFARX1 I_52531 (I896609,I3563,I896459,I896635,);
not I_52532 (I896643,I896635);
nor I_52533 (I896451,I896493,I896643);
DFFARX1 I_52534 (I990481,I3563,I896459,I896683,);
nor I_52535 (I896442,I896683,I896553);
nor I_52536 (I896433,I896683,I896609);
nand I_52537 (I896719,I990478,I990469);
and I_52538 (I896736,I896719,I990463);
DFFARX1 I_52539 (I896736,I3563,I896459,I896762,);
not I_52540 (I896770,I896762);
nand I_52541 (I896787,I896770,I896683);
nand I_52542 (I896436,I896770,I896592);
nor I_52543 (I896818,I990472,I990469);
and I_52544 (I896835,I896683,I896818);
nor I_52545 (I896852,I896770,I896835);
DFFARX1 I_52546 (I896852,I3563,I896459,I896445,);
nor I_52547 (I896883,I896485,I896818);
DFFARX1 I_52548 (I896883,I3563,I896459,I896430,);
nor I_52549 (I896914,I896762,I896818);
not I_52550 (I896931,I896914);
nand I_52551 (I896439,I896931,I896787);
not I_52552 (I896986,I3570);
DFFARX1 I_52553 (I1280693,I3563,I896986,I897012,);
not I_52554 (I897020,I897012);
nand I_52555 (I897037,I1280699,I1280681);
and I_52556 (I897054,I897037,I1280690);
DFFARX1 I_52557 (I897054,I3563,I896986,I897080,);
DFFARX1 I_52558 (I897080,I3563,I896986,I896975,);
DFFARX1 I_52559 (I1280696,I3563,I896986,I897111,);
nand I_52560 (I897119,I897111,I1280684);
not I_52561 (I897136,I897119);
DFFARX1 I_52562 (I897136,I3563,I896986,I897162,);
not I_52563 (I897170,I897162);
nor I_52564 (I896978,I897020,I897170);
DFFARX1 I_52565 (I1280702,I3563,I896986,I897210,);
nor I_52566 (I896969,I897210,I897080);
nor I_52567 (I896960,I897210,I897136);
nand I_52568 (I897246,I1280681,I1280687);
and I_52569 (I897263,I897246,I1280705);
DFFARX1 I_52570 (I897263,I3563,I896986,I897289,);
not I_52571 (I897297,I897289);
nand I_52572 (I897314,I897297,I897210);
nand I_52573 (I896963,I897297,I897119);
nor I_52574 (I897345,I1280684,I1280687);
and I_52575 (I897362,I897210,I897345);
nor I_52576 (I897379,I897297,I897362);
DFFARX1 I_52577 (I897379,I3563,I896986,I896972,);
nor I_52578 (I897410,I897012,I897345);
DFFARX1 I_52579 (I897410,I3563,I896986,I896957,);
nor I_52580 (I897441,I897289,I897345);
not I_52581 (I897458,I897441);
nand I_52582 (I896966,I897458,I897314);
not I_52583 (I897513,I3570);
DFFARX1 I_52584 (I1038910,I3563,I897513,I897539,);
not I_52585 (I897547,I897539);
nand I_52586 (I897564,I1038925,I1038907);
and I_52587 (I897581,I897564,I1038907);
DFFARX1 I_52588 (I897581,I3563,I897513,I897607,);
DFFARX1 I_52589 (I897607,I3563,I897513,I897502,);
DFFARX1 I_52590 (I1038916,I3563,I897513,I897638,);
nand I_52591 (I897646,I897638,I1038934);
not I_52592 (I897663,I897646);
DFFARX1 I_52593 (I897663,I3563,I897513,I897689,);
not I_52594 (I897697,I897689);
nor I_52595 (I897505,I897547,I897697);
DFFARX1 I_52596 (I1038931,I3563,I897513,I897737,);
nor I_52597 (I897496,I897737,I897607);
nor I_52598 (I897487,I897737,I897663);
nand I_52599 (I897773,I1038928,I1038919);
and I_52600 (I897790,I897773,I1038913);
DFFARX1 I_52601 (I897790,I3563,I897513,I897816,);
not I_52602 (I897824,I897816);
nand I_52603 (I897841,I897824,I897737);
nand I_52604 (I897490,I897824,I897646);
nor I_52605 (I897872,I1038922,I1038919);
and I_52606 (I897889,I897737,I897872);
nor I_52607 (I897906,I897824,I897889);
DFFARX1 I_52608 (I897906,I3563,I897513,I897499,);
nor I_52609 (I897937,I897539,I897872);
DFFARX1 I_52610 (I897937,I3563,I897513,I897484,);
nor I_52611 (I897968,I897816,I897872);
not I_52612 (I897985,I897968);
nand I_52613 (I897493,I897985,I897841);
not I_52614 (I898040,I3570);
DFFARX1 I_52615 (I422952,I3563,I898040,I898066,);
not I_52616 (I898074,I898066);
nand I_52617 (I898091,I422949,I422958);
and I_52618 (I898108,I898091,I422967);
DFFARX1 I_52619 (I898108,I3563,I898040,I898134,);
DFFARX1 I_52620 (I898134,I3563,I898040,I898029,);
DFFARX1 I_52621 (I422970,I3563,I898040,I898165,);
nand I_52622 (I898173,I898165,I422973);
not I_52623 (I898190,I898173);
DFFARX1 I_52624 (I898190,I3563,I898040,I898216,);
not I_52625 (I898224,I898216);
nor I_52626 (I898032,I898074,I898224);
DFFARX1 I_52627 (I422946,I3563,I898040,I898264,);
nor I_52628 (I898023,I898264,I898134);
nor I_52629 (I898014,I898264,I898190);
nand I_52630 (I898300,I422961,I422964);
and I_52631 (I898317,I898300,I422955);
DFFARX1 I_52632 (I898317,I3563,I898040,I898343,);
not I_52633 (I898351,I898343);
nand I_52634 (I898368,I898351,I898264);
nand I_52635 (I898017,I898351,I898173);
nor I_52636 (I898399,I422946,I422964);
and I_52637 (I898416,I898264,I898399);
nor I_52638 (I898433,I898351,I898416);
DFFARX1 I_52639 (I898433,I3563,I898040,I898026,);
nor I_52640 (I898464,I898066,I898399);
DFFARX1 I_52641 (I898464,I3563,I898040,I898011,);
nor I_52642 (I898495,I898343,I898399);
not I_52643 (I898512,I898495);
nand I_52644 (I898020,I898512,I898368);
not I_52645 (I898567,I3570);
DFFARX1 I_52646 (I1053400,I3563,I898567,I898593,);
not I_52647 (I898601,I898593);
nand I_52648 (I898618,I1053409,I1053397);
and I_52649 (I898635,I898618,I1053394);
DFFARX1 I_52650 (I898635,I3563,I898567,I898661,);
DFFARX1 I_52651 (I898661,I3563,I898567,I898556,);
DFFARX1 I_52652 (I1053394,I3563,I898567,I898692,);
nand I_52653 (I898700,I898692,I1053391);
not I_52654 (I898717,I898700);
DFFARX1 I_52655 (I898717,I3563,I898567,I898743,);
not I_52656 (I898751,I898743);
nor I_52657 (I898559,I898601,I898751);
DFFARX1 I_52658 (I1053397,I3563,I898567,I898791,);
nor I_52659 (I898550,I898791,I898661);
nor I_52660 (I898541,I898791,I898717);
nand I_52661 (I898827,I1053412,I1053403);
and I_52662 (I898844,I898827,I1053406);
DFFARX1 I_52663 (I898844,I3563,I898567,I898870,);
not I_52664 (I898878,I898870);
nand I_52665 (I898895,I898878,I898791);
nand I_52666 (I898544,I898878,I898700);
nor I_52667 (I898926,I1053391,I1053403);
and I_52668 (I898943,I898791,I898926);
nor I_52669 (I898960,I898878,I898943);
DFFARX1 I_52670 (I898960,I3563,I898567,I898553,);
nor I_52671 (I898991,I898593,I898926);
DFFARX1 I_52672 (I898991,I3563,I898567,I898538,);
nor I_52673 (I899022,I898870,I898926);
not I_52674 (I899039,I899022);
nand I_52675 (I898547,I899039,I898895);
not I_52676 (I899094,I3570);
DFFARX1 I_52677 (I56656,I3563,I899094,I899120,);
not I_52678 (I899128,I899120);
nand I_52679 (I899145,I56668,I56671);
and I_52680 (I899162,I899145,I56647);
DFFARX1 I_52681 (I899162,I3563,I899094,I899188,);
DFFARX1 I_52682 (I899188,I3563,I899094,I899083,);
DFFARX1 I_52683 (I56665,I3563,I899094,I899219,);
nand I_52684 (I899227,I899219,I56653);
not I_52685 (I899244,I899227);
DFFARX1 I_52686 (I899244,I3563,I899094,I899270,);
not I_52687 (I899278,I899270);
nor I_52688 (I899086,I899128,I899278);
DFFARX1 I_52689 (I56650,I3563,I899094,I899318,);
nor I_52690 (I899077,I899318,I899188);
nor I_52691 (I899068,I899318,I899244);
nand I_52692 (I899354,I56659,I56650);
and I_52693 (I899371,I899354,I56647);
DFFARX1 I_52694 (I899371,I3563,I899094,I899397,);
not I_52695 (I899405,I899397);
nand I_52696 (I899422,I899405,I899318);
nand I_52697 (I899071,I899405,I899227);
nor I_52698 (I899453,I56662,I56650);
and I_52699 (I899470,I899318,I899453);
nor I_52700 (I899487,I899405,I899470);
DFFARX1 I_52701 (I899487,I3563,I899094,I899080,);
nor I_52702 (I899518,I899120,I899453);
DFFARX1 I_52703 (I899518,I3563,I899094,I899065,);
nor I_52704 (I899549,I899397,I899453);
not I_52705 (I899566,I899549);
nand I_52706 (I899074,I899566,I899422);
not I_52707 (I899621,I3570);
DFFARX1 I_52708 (I128343,I3563,I899621,I899647,);
not I_52709 (I899655,I899647);
nand I_52710 (I899672,I128319,I128328);
and I_52711 (I899689,I899672,I128322);
DFFARX1 I_52712 (I899689,I3563,I899621,I899715,);
DFFARX1 I_52713 (I899715,I3563,I899621,I899610,);
DFFARX1 I_52714 (I128340,I3563,I899621,I899746,);
nand I_52715 (I899754,I899746,I128331);
not I_52716 (I899771,I899754);
DFFARX1 I_52717 (I899771,I3563,I899621,I899797,);
not I_52718 (I899805,I899797);
nor I_52719 (I899613,I899655,I899805);
DFFARX1 I_52720 (I128325,I3563,I899621,I899845,);
nor I_52721 (I899604,I899845,I899715);
nor I_52722 (I899595,I899845,I899771);
nand I_52723 (I899881,I128337,I128334);
and I_52724 (I899898,I899881,I128322);
DFFARX1 I_52725 (I899898,I3563,I899621,I899924,);
not I_52726 (I899932,I899924);
nand I_52727 (I899949,I899932,I899845);
nand I_52728 (I899598,I899932,I899754);
nor I_52729 (I899980,I128319,I128334);
and I_52730 (I899997,I899845,I899980);
nor I_52731 (I900014,I899932,I899997);
DFFARX1 I_52732 (I900014,I3563,I899621,I899607,);
nor I_52733 (I900045,I899647,I899980);
DFFARX1 I_52734 (I900045,I3563,I899621,I899592,);
nor I_52735 (I900076,I899924,I899980);
not I_52736 (I900093,I900076);
nand I_52737 (I899601,I900093,I899949);
not I_52738 (I900148,I3570);
DFFARX1 I_52739 (I232144,I3563,I900148,I900174,);
not I_52740 (I900182,I900174);
nand I_52741 (I900199,I232141,I232159);
and I_52742 (I900216,I900199,I232150);
DFFARX1 I_52743 (I900216,I3563,I900148,I900242,);
DFFARX1 I_52744 (I900242,I3563,I900148,I900137,);
DFFARX1 I_52745 (I232156,I3563,I900148,I900273,);
nand I_52746 (I900281,I900273,I232153);
not I_52747 (I900298,I900281);
DFFARX1 I_52748 (I900298,I3563,I900148,I900324,);
not I_52749 (I900332,I900324);
nor I_52750 (I900140,I900182,I900332);
DFFARX1 I_52751 (I232147,I3563,I900148,I900372,);
nor I_52752 (I900131,I900372,I900242);
nor I_52753 (I900122,I900372,I900298);
nand I_52754 (I900408,I232138,I232162);
and I_52755 (I900425,I900408,I232141);
DFFARX1 I_52756 (I900425,I3563,I900148,I900451,);
not I_52757 (I900459,I900451);
nand I_52758 (I900476,I900459,I900372);
nand I_52759 (I900125,I900459,I900281);
nor I_52760 (I900507,I232138,I232162);
and I_52761 (I900524,I900372,I900507);
nor I_52762 (I900541,I900459,I900524);
DFFARX1 I_52763 (I900541,I3563,I900148,I900134,);
nor I_52764 (I900572,I900174,I900507);
DFFARX1 I_52765 (I900572,I3563,I900148,I900119,);
nor I_52766 (I900603,I900451,I900507);
not I_52767 (I900620,I900603);
nand I_52768 (I900128,I900620,I900476);
not I_52769 (I900675,I3570);
DFFARX1 I_52770 (I667083,I3563,I900675,I900701,);
not I_52771 (I900709,I900701);
nand I_52772 (I900726,I667086,I667083);
and I_52773 (I900743,I900726,I667095);
DFFARX1 I_52774 (I900743,I3563,I900675,I900769,);
DFFARX1 I_52775 (I900769,I3563,I900675,I900664,);
DFFARX1 I_52776 (I667092,I3563,I900675,I900800,);
nand I_52777 (I900808,I900800,I667098);
not I_52778 (I900825,I900808);
DFFARX1 I_52779 (I900825,I3563,I900675,I900851,);
not I_52780 (I900859,I900851);
nor I_52781 (I900667,I900709,I900859);
DFFARX1 I_52782 (I667107,I3563,I900675,I900899,);
nor I_52783 (I900658,I900899,I900769);
nor I_52784 (I900649,I900899,I900825);
nand I_52785 (I900935,I667101,I667089);
and I_52786 (I900952,I900935,I667086);
DFFARX1 I_52787 (I900952,I3563,I900675,I900978,);
not I_52788 (I900986,I900978);
nand I_52789 (I901003,I900986,I900899);
nand I_52790 (I900652,I900986,I900808);
nor I_52791 (I901034,I667104,I667089);
and I_52792 (I901051,I900899,I901034);
nor I_52793 (I901068,I900986,I901051);
DFFARX1 I_52794 (I901068,I3563,I900675,I900661,);
nor I_52795 (I901099,I900701,I901034);
DFFARX1 I_52796 (I901099,I3563,I900675,I900646,);
nor I_52797 (I901130,I900978,I901034);
not I_52798 (I901147,I901130);
nand I_52799 (I900655,I901147,I901003);
not I_52800 (I901202,I3570);
DFFARX1 I_52801 (I420813,I3563,I901202,I901228,);
not I_52802 (I901236,I901228);
nand I_52803 (I901253,I420804,I420804);
and I_52804 (I901270,I901253,I420822);
DFFARX1 I_52805 (I901270,I3563,I901202,I901296,);
DFFARX1 I_52806 (I901296,I3563,I901202,I901191,);
DFFARX1 I_52807 (I420825,I3563,I901202,I901327,);
nand I_52808 (I901335,I901327,I420807);
not I_52809 (I901352,I901335);
DFFARX1 I_52810 (I901352,I3563,I901202,I901378,);
not I_52811 (I901386,I901378);
nor I_52812 (I901194,I901236,I901386);
DFFARX1 I_52813 (I420819,I3563,I901202,I901426,);
nor I_52814 (I901185,I901426,I901296);
nor I_52815 (I901176,I901426,I901352);
nand I_52816 (I901462,I420831,I420810);
and I_52817 (I901479,I901462,I420816);
DFFARX1 I_52818 (I901479,I3563,I901202,I901505,);
not I_52819 (I901513,I901505);
nand I_52820 (I901530,I901513,I901426);
nand I_52821 (I901179,I901513,I901335);
nor I_52822 (I901561,I420828,I420810);
and I_52823 (I901578,I901426,I901561);
nor I_52824 (I901595,I901513,I901578);
DFFARX1 I_52825 (I901595,I3563,I901202,I901188,);
nor I_52826 (I901626,I901228,I901561);
DFFARX1 I_52827 (I901626,I3563,I901202,I901173,);
nor I_52828 (I901657,I901505,I901561);
not I_52829 (I901674,I901657);
nand I_52830 (I901182,I901674,I901530);
not I_52831 (I901729,I3570);
DFFARX1 I_52832 (I208939,I3563,I901729,I901755,);
not I_52833 (I901763,I901755);
nand I_52834 (I901780,I208936,I208954);
and I_52835 (I901797,I901780,I208945);
DFFARX1 I_52836 (I901797,I3563,I901729,I901823,);
DFFARX1 I_52837 (I901823,I3563,I901729,I901718,);
DFFARX1 I_52838 (I208951,I3563,I901729,I901854,);
nand I_52839 (I901862,I901854,I208948);
not I_52840 (I901879,I901862);
DFFARX1 I_52841 (I901879,I3563,I901729,I901905,);
not I_52842 (I901913,I901905);
nor I_52843 (I901721,I901763,I901913);
DFFARX1 I_52844 (I208942,I3563,I901729,I901953,);
nor I_52845 (I901712,I901953,I901823);
nor I_52846 (I901703,I901953,I901879);
nand I_52847 (I901989,I208933,I208957);
and I_52848 (I902006,I901989,I208936);
DFFARX1 I_52849 (I902006,I3563,I901729,I902032,);
not I_52850 (I902040,I902032);
nand I_52851 (I902057,I902040,I901953);
nand I_52852 (I901706,I902040,I901862);
nor I_52853 (I902088,I208933,I208957);
and I_52854 (I902105,I901953,I902088);
nor I_52855 (I902122,I902040,I902105);
DFFARX1 I_52856 (I902122,I3563,I901729,I901715,);
nor I_52857 (I902153,I901755,I902088);
DFFARX1 I_52858 (I902153,I3563,I901729,I901700,);
nor I_52859 (I902184,I902032,I902088);
not I_52860 (I902201,I902184);
nand I_52861 (I901709,I902201,I902057);
not I_52862 (I902256,I3570);
DFFARX1 I_52863 (I1057327,I3563,I902256,I902282,);
not I_52864 (I902290,I902282);
nand I_52865 (I902307,I1057336,I1057324);
and I_52866 (I902324,I902307,I1057321);
DFFARX1 I_52867 (I902324,I3563,I902256,I902350,);
DFFARX1 I_52868 (I902350,I3563,I902256,I902245,);
DFFARX1 I_52869 (I1057321,I3563,I902256,I902381,);
nand I_52870 (I902389,I902381,I1057318);
not I_52871 (I902406,I902389);
DFFARX1 I_52872 (I902406,I3563,I902256,I902432,);
not I_52873 (I902440,I902432);
nor I_52874 (I902248,I902290,I902440);
DFFARX1 I_52875 (I1057324,I3563,I902256,I902480,);
nor I_52876 (I902239,I902480,I902350);
nor I_52877 (I902230,I902480,I902406);
nand I_52878 (I902516,I1057339,I1057330);
and I_52879 (I902533,I902516,I1057333);
DFFARX1 I_52880 (I902533,I3563,I902256,I902559,);
not I_52881 (I902567,I902559);
nand I_52882 (I902584,I902567,I902480);
nand I_52883 (I902233,I902567,I902389);
nor I_52884 (I902615,I1057318,I1057330);
and I_52885 (I902632,I902480,I902615);
nor I_52886 (I902649,I902567,I902632);
DFFARX1 I_52887 (I902649,I3563,I902256,I902242,);
nor I_52888 (I902680,I902282,I902615);
DFFARX1 I_52889 (I902680,I3563,I902256,I902227,);
nor I_52890 (I902711,I902559,I902615);
not I_52891 (I902728,I902711);
nand I_52892 (I902236,I902728,I902584);
not I_52893 (I902783,I3570);
DFFARX1 I_52894 (I665349,I3563,I902783,I902809,);
not I_52895 (I902817,I902809);
nand I_52896 (I902834,I665352,I665349);
and I_52897 (I902851,I902834,I665361);
DFFARX1 I_52898 (I902851,I3563,I902783,I902877,);
DFFARX1 I_52899 (I902877,I3563,I902783,I902772,);
DFFARX1 I_52900 (I665358,I3563,I902783,I902908,);
nand I_52901 (I902916,I902908,I665364);
not I_52902 (I902933,I902916);
DFFARX1 I_52903 (I902933,I3563,I902783,I902959,);
not I_52904 (I902967,I902959);
nor I_52905 (I902775,I902817,I902967);
DFFARX1 I_52906 (I665373,I3563,I902783,I903007,);
nor I_52907 (I902766,I903007,I902877);
nor I_52908 (I902757,I903007,I902933);
nand I_52909 (I903043,I665367,I665355);
and I_52910 (I903060,I903043,I665352);
DFFARX1 I_52911 (I903060,I3563,I902783,I903086,);
not I_52912 (I903094,I903086);
nand I_52913 (I903111,I903094,I903007);
nand I_52914 (I902760,I903094,I902916);
nor I_52915 (I903142,I665370,I665355);
and I_52916 (I903159,I903007,I903142);
nor I_52917 (I903176,I903094,I903159);
DFFARX1 I_52918 (I903176,I3563,I902783,I902769,);
nor I_52919 (I903207,I902809,I903142);
DFFARX1 I_52920 (I903207,I3563,I902783,I902754,);
nor I_52921 (I903238,I903086,I903142);
not I_52922 (I903255,I903238);
nand I_52923 (I902763,I903255,I903111);
not I_52924 (I903310,I3570);
DFFARX1 I_52925 (I185734,I3563,I903310,I903336,);
not I_52926 (I903344,I903336);
nand I_52927 (I903361,I185731,I185749);
and I_52928 (I903378,I903361,I185740);
DFFARX1 I_52929 (I903378,I3563,I903310,I903404,);
DFFARX1 I_52930 (I903404,I3563,I903310,I903299,);
DFFARX1 I_52931 (I185746,I3563,I903310,I903435,);
nand I_52932 (I903443,I903435,I185743);
not I_52933 (I903460,I903443);
DFFARX1 I_52934 (I903460,I3563,I903310,I903486,);
not I_52935 (I903494,I903486);
nor I_52936 (I903302,I903344,I903494);
DFFARX1 I_52937 (I185737,I3563,I903310,I903534,);
nor I_52938 (I903293,I903534,I903404);
nor I_52939 (I903284,I903534,I903460);
nand I_52940 (I903570,I185728,I185752);
and I_52941 (I903587,I903570,I185731);
DFFARX1 I_52942 (I903587,I3563,I903310,I903613,);
not I_52943 (I903621,I903613);
nand I_52944 (I903638,I903621,I903534);
nand I_52945 (I903287,I903621,I903443);
nor I_52946 (I903669,I185728,I185752);
and I_52947 (I903686,I903534,I903669);
nor I_52948 (I903703,I903621,I903686);
DFFARX1 I_52949 (I903703,I3563,I903310,I903296,);
nor I_52950 (I903734,I903336,I903669);
DFFARX1 I_52951 (I903734,I3563,I903310,I903281,);
nor I_52952 (I903765,I903613,I903669);
not I_52953 (I903782,I903765);
nand I_52954 (I903290,I903782,I903638);
not I_52955 (I903837,I3570);
DFFARX1 I_52956 (I467016,I3563,I903837,I903863,);
not I_52957 (I903871,I903863);
nand I_52958 (I903888,I467013,I467022);
and I_52959 (I903905,I903888,I467031);
DFFARX1 I_52960 (I903905,I3563,I903837,I903931,);
DFFARX1 I_52961 (I903931,I3563,I903837,I903826,);
DFFARX1 I_52962 (I467034,I3563,I903837,I903962,);
nand I_52963 (I903970,I903962,I467037);
not I_52964 (I903987,I903970);
DFFARX1 I_52965 (I903987,I3563,I903837,I904013,);
not I_52966 (I904021,I904013);
nor I_52967 (I903829,I903871,I904021);
DFFARX1 I_52968 (I467010,I3563,I903837,I904061,);
nor I_52969 (I903820,I904061,I903931);
nor I_52970 (I903811,I904061,I903987);
nand I_52971 (I904097,I467025,I467028);
and I_52972 (I904114,I904097,I467019);
DFFARX1 I_52973 (I904114,I3563,I903837,I904140,);
not I_52974 (I904148,I904140);
nand I_52975 (I904165,I904148,I904061);
nand I_52976 (I903814,I904148,I903970);
nor I_52977 (I904196,I467010,I467028);
and I_52978 (I904213,I904061,I904196);
nor I_52979 (I904230,I904148,I904213);
DFFARX1 I_52980 (I904230,I3563,I903837,I903823,);
nor I_52981 (I904261,I903863,I904196);
DFFARX1 I_52982 (I904261,I3563,I903837,I903808,);
nor I_52983 (I904292,I904140,I904196);
not I_52984 (I904309,I904292);
nand I_52985 (I903817,I904309,I904165);
not I_52986 (I904364,I3570);
DFFARX1 I_52987 (I477352,I3563,I904364,I904390,);
not I_52988 (I904398,I904390);
nand I_52989 (I904415,I477349,I477358);
and I_52990 (I904432,I904415,I477367);
DFFARX1 I_52991 (I904432,I3563,I904364,I904458,);
DFFARX1 I_52992 (I904458,I3563,I904364,I904353,);
DFFARX1 I_52993 (I477370,I3563,I904364,I904489,);
nand I_52994 (I904497,I904489,I477373);
not I_52995 (I904514,I904497);
DFFARX1 I_52996 (I904514,I3563,I904364,I904540,);
not I_52997 (I904548,I904540);
nor I_52998 (I904356,I904398,I904548);
DFFARX1 I_52999 (I477346,I3563,I904364,I904588,);
nor I_53000 (I904347,I904588,I904458);
nor I_53001 (I904338,I904588,I904514);
nand I_53002 (I904624,I477361,I477364);
and I_53003 (I904641,I904624,I477355);
DFFARX1 I_53004 (I904641,I3563,I904364,I904667,);
not I_53005 (I904675,I904667);
nand I_53006 (I904692,I904675,I904588);
nand I_53007 (I904341,I904675,I904497);
nor I_53008 (I904723,I477346,I477364);
and I_53009 (I904740,I904588,I904723);
nor I_53010 (I904757,I904675,I904740);
DFFARX1 I_53011 (I904757,I3563,I904364,I904350,);
nor I_53012 (I904788,I904390,I904723);
DFFARX1 I_53013 (I904788,I3563,I904364,I904335,);
nor I_53014 (I904819,I904667,I904723);
not I_53015 (I904836,I904819);
nand I_53016 (I904344,I904836,I904692);
not I_53017 (I904891,I3570);
DFFARX1 I_53018 (I580976,I3563,I904891,I904917,);
not I_53019 (I904925,I904917);
nand I_53020 (I904942,I580961,I580982);
and I_53021 (I904959,I904942,I580970);
DFFARX1 I_53022 (I904959,I3563,I904891,I904985,);
DFFARX1 I_53023 (I904985,I3563,I904891,I904880,);
DFFARX1 I_53024 (I580964,I3563,I904891,I905016,);
nand I_53025 (I905024,I905016,I580973);
not I_53026 (I905041,I905024);
DFFARX1 I_53027 (I905041,I3563,I904891,I905067,);
not I_53028 (I905075,I905067);
nor I_53029 (I904883,I904925,I905075);
DFFARX1 I_53030 (I580979,I3563,I904891,I905115,);
nor I_53031 (I904874,I905115,I904985);
nor I_53032 (I904865,I905115,I905041);
nand I_53033 (I905151,I580961,I580964);
and I_53034 (I905168,I905151,I580985);
DFFARX1 I_53035 (I905168,I3563,I904891,I905194,);
not I_53036 (I905202,I905194);
nand I_53037 (I905219,I905202,I905115);
nand I_53038 (I904868,I905202,I905024);
nor I_53039 (I905250,I580967,I580964);
and I_53040 (I905267,I905115,I905250);
nor I_53041 (I905284,I905202,I905267);
DFFARX1 I_53042 (I905284,I3563,I904891,I904877,);
nor I_53043 (I905315,I904917,I905250);
DFFARX1 I_53044 (I905315,I3563,I904891,I904862,);
nor I_53045 (I905346,I905194,I905250);
not I_53046 (I905363,I905346);
nand I_53047 (I904871,I905363,I905219);
not I_53048 (I905418,I3570);
DFFARX1 I_53049 (I24509,I3563,I905418,I905444,);
not I_53050 (I905452,I905444);
nand I_53051 (I905469,I24521,I24524);
and I_53052 (I905486,I905469,I24500);
DFFARX1 I_53053 (I905486,I3563,I905418,I905512,);
DFFARX1 I_53054 (I905512,I3563,I905418,I905407,);
DFFARX1 I_53055 (I24518,I3563,I905418,I905543,);
nand I_53056 (I905551,I905543,I24506);
not I_53057 (I905568,I905551);
DFFARX1 I_53058 (I905568,I3563,I905418,I905594,);
not I_53059 (I905602,I905594);
nor I_53060 (I905410,I905452,I905602);
DFFARX1 I_53061 (I24503,I3563,I905418,I905642,);
nor I_53062 (I905401,I905642,I905512);
nor I_53063 (I905392,I905642,I905568);
nand I_53064 (I905678,I24512,I24503);
and I_53065 (I905695,I905678,I24500);
DFFARX1 I_53066 (I905695,I3563,I905418,I905721,);
not I_53067 (I905729,I905721);
nand I_53068 (I905746,I905729,I905642);
nand I_53069 (I905395,I905729,I905551);
nor I_53070 (I905777,I24515,I24503);
and I_53071 (I905794,I905642,I905777);
nor I_53072 (I905811,I905729,I905794);
DFFARX1 I_53073 (I905811,I3563,I905418,I905404,);
nor I_53074 (I905842,I905444,I905777);
DFFARX1 I_53075 (I905842,I3563,I905418,I905389,);
nor I_53076 (I905873,I905721,I905777);
not I_53077 (I905890,I905873);
nand I_53078 (I905398,I905890,I905746);
not I_53079 (I905945,I3570);
DFFARX1 I_53080 (I427848,I3563,I905945,I905971,);
not I_53081 (I905979,I905971);
nand I_53082 (I905996,I427845,I427854);
and I_53083 (I906013,I905996,I427863);
DFFARX1 I_53084 (I906013,I3563,I905945,I906039,);
DFFARX1 I_53085 (I906039,I3563,I905945,I905934,);
DFFARX1 I_53086 (I427866,I3563,I905945,I906070,);
nand I_53087 (I906078,I906070,I427869);
not I_53088 (I906095,I906078);
DFFARX1 I_53089 (I906095,I3563,I905945,I906121,);
not I_53090 (I906129,I906121);
nor I_53091 (I905937,I905979,I906129);
DFFARX1 I_53092 (I427842,I3563,I905945,I906169,);
nor I_53093 (I905928,I906169,I906039);
nor I_53094 (I905919,I906169,I906095);
nand I_53095 (I906205,I427857,I427860);
and I_53096 (I906222,I906205,I427851);
DFFARX1 I_53097 (I906222,I3563,I905945,I906248,);
not I_53098 (I906256,I906248);
nand I_53099 (I906273,I906256,I906169);
nand I_53100 (I905922,I906256,I906078);
nor I_53101 (I906304,I427842,I427860);
and I_53102 (I906321,I906169,I906304);
nor I_53103 (I906338,I906256,I906321);
DFFARX1 I_53104 (I906338,I3563,I905945,I905931,);
nor I_53105 (I906369,I905971,I906304);
DFFARX1 I_53106 (I906369,I3563,I905945,I905916,);
nor I_53107 (I906400,I906248,I906304);
not I_53108 (I906417,I906400);
nand I_53109 (I905925,I906417,I906273);
not I_53110 (I906472,I3570);
DFFARX1 I_53111 (I355465,I3563,I906472,I906498,);
not I_53112 (I906506,I906498);
nand I_53113 (I906523,I355456,I355456);
and I_53114 (I906540,I906523,I355474);
DFFARX1 I_53115 (I906540,I3563,I906472,I906566,);
DFFARX1 I_53116 (I906566,I3563,I906472,I906461,);
DFFARX1 I_53117 (I355477,I3563,I906472,I906597,);
nand I_53118 (I906605,I906597,I355459);
not I_53119 (I906622,I906605);
DFFARX1 I_53120 (I906622,I3563,I906472,I906648,);
not I_53121 (I906656,I906648);
nor I_53122 (I906464,I906506,I906656);
DFFARX1 I_53123 (I355471,I3563,I906472,I906696,);
nor I_53124 (I906455,I906696,I906566);
nor I_53125 (I906446,I906696,I906622);
nand I_53126 (I906732,I355483,I355462);
and I_53127 (I906749,I906732,I355468);
DFFARX1 I_53128 (I906749,I3563,I906472,I906775,);
not I_53129 (I906783,I906775);
nand I_53130 (I906800,I906783,I906696);
nand I_53131 (I906449,I906783,I906605);
nor I_53132 (I906831,I355480,I355462);
and I_53133 (I906848,I906696,I906831);
nor I_53134 (I906865,I906783,I906848);
DFFARX1 I_53135 (I906865,I3563,I906472,I906458,);
nor I_53136 (I906896,I906498,I906831);
DFFARX1 I_53137 (I906896,I3563,I906472,I906443,);
nor I_53138 (I906927,I906775,I906831);
not I_53139 (I906944,I906927);
nand I_53140 (I906452,I906944,I906800);
not I_53141 (I906999,I3570);
DFFARX1 I_53142 (I734709,I3563,I906999,I907025,);
not I_53143 (I907033,I907025);
nand I_53144 (I907050,I734712,I734709);
and I_53145 (I907067,I907050,I734721);
DFFARX1 I_53146 (I907067,I3563,I906999,I907093,);
DFFARX1 I_53147 (I907093,I3563,I906999,I906988,);
DFFARX1 I_53148 (I734718,I3563,I906999,I907124,);
nand I_53149 (I907132,I907124,I734724);
not I_53150 (I907149,I907132);
DFFARX1 I_53151 (I907149,I3563,I906999,I907175,);
not I_53152 (I907183,I907175);
nor I_53153 (I906991,I907033,I907183);
DFFARX1 I_53154 (I734733,I3563,I906999,I907223,);
nor I_53155 (I906982,I907223,I907093);
nor I_53156 (I906973,I907223,I907149);
nand I_53157 (I907259,I734727,I734715);
and I_53158 (I907276,I907259,I734712);
DFFARX1 I_53159 (I907276,I3563,I906999,I907302,);
not I_53160 (I907310,I907302);
nand I_53161 (I907327,I907310,I907223);
nand I_53162 (I906976,I907310,I907132);
nor I_53163 (I907358,I734730,I734715);
and I_53164 (I907375,I907223,I907358);
nor I_53165 (I907392,I907310,I907375);
DFFARX1 I_53166 (I907392,I3563,I906999,I906985,);
nor I_53167 (I907423,I907025,I907358);
DFFARX1 I_53168 (I907423,I3563,I906999,I906970,);
nor I_53169 (I907454,I907302,I907358);
not I_53170 (I907471,I907454);
nand I_53171 (I906979,I907471,I907327);
not I_53172 (I907526,I3570);
DFFARX1 I_53173 (I983354,I3563,I907526,I907552,);
not I_53174 (I907560,I907552);
nand I_53175 (I907577,I983369,I983351);
and I_53176 (I907594,I907577,I983351);
DFFARX1 I_53177 (I907594,I3563,I907526,I907620,);
DFFARX1 I_53178 (I907620,I3563,I907526,I907515,);
DFFARX1 I_53179 (I983360,I3563,I907526,I907651,);
nand I_53180 (I907659,I907651,I983378);
not I_53181 (I907676,I907659);
DFFARX1 I_53182 (I907676,I3563,I907526,I907702,);
not I_53183 (I907710,I907702);
nor I_53184 (I907518,I907560,I907710);
DFFARX1 I_53185 (I983375,I3563,I907526,I907750,);
nor I_53186 (I907509,I907750,I907620);
nor I_53187 (I907500,I907750,I907676);
nand I_53188 (I907786,I983372,I983363);
and I_53189 (I907803,I907786,I983357);
DFFARX1 I_53190 (I907803,I3563,I907526,I907829,);
not I_53191 (I907837,I907829);
nand I_53192 (I907854,I907837,I907750);
nand I_53193 (I907503,I907837,I907659);
nor I_53194 (I907885,I983366,I983363);
and I_53195 (I907902,I907750,I907885);
nor I_53196 (I907919,I907837,I907902);
DFFARX1 I_53197 (I907919,I3563,I907526,I907512,);
nor I_53198 (I907950,I907552,I907885);
DFFARX1 I_53199 (I907950,I3563,I907526,I907497,);
nor I_53200 (I907981,I907829,I907885);
not I_53201 (I907998,I907981);
nand I_53202 (I907506,I907998,I907854);
not I_53203 (I908053,I3570);
DFFARX1 I_53204 (I52967,I3563,I908053,I908079,);
not I_53205 (I908087,I908079);
nand I_53206 (I908104,I52979,I52982);
and I_53207 (I908121,I908104,I52958);
DFFARX1 I_53208 (I908121,I3563,I908053,I908147,);
DFFARX1 I_53209 (I908147,I3563,I908053,I908042,);
DFFARX1 I_53210 (I52976,I3563,I908053,I908178,);
nand I_53211 (I908186,I908178,I52964);
not I_53212 (I908203,I908186);
DFFARX1 I_53213 (I908203,I3563,I908053,I908229,);
not I_53214 (I908237,I908229);
nor I_53215 (I908045,I908087,I908237);
DFFARX1 I_53216 (I52961,I3563,I908053,I908277,);
nor I_53217 (I908036,I908277,I908147);
nor I_53218 (I908027,I908277,I908203);
nand I_53219 (I908313,I52970,I52961);
and I_53220 (I908330,I908313,I52958);
DFFARX1 I_53221 (I908330,I3563,I908053,I908356,);
not I_53222 (I908364,I908356);
nand I_53223 (I908381,I908364,I908277);
nand I_53224 (I908030,I908364,I908186);
nor I_53225 (I908412,I52973,I52961);
and I_53226 (I908429,I908277,I908412);
nor I_53227 (I908446,I908364,I908429);
DFFARX1 I_53228 (I908446,I3563,I908053,I908039,);
nor I_53229 (I908477,I908079,I908412);
DFFARX1 I_53230 (I908477,I3563,I908053,I908024,);
nor I_53231 (I908508,I908356,I908412);
not I_53232 (I908525,I908508);
nand I_53233 (I908033,I908525,I908381);
not I_53234 (I908580,I3570);
DFFARX1 I_53235 (I731241,I3563,I908580,I908606,);
not I_53236 (I908614,I908606);
nand I_53237 (I908631,I731244,I731241);
and I_53238 (I908648,I908631,I731253);
DFFARX1 I_53239 (I908648,I3563,I908580,I908674,);
DFFARX1 I_53240 (I908674,I3563,I908580,I908569,);
DFFARX1 I_53241 (I731250,I3563,I908580,I908705,);
nand I_53242 (I908713,I908705,I731256);
not I_53243 (I908730,I908713);
DFFARX1 I_53244 (I908730,I3563,I908580,I908756,);
not I_53245 (I908764,I908756);
nor I_53246 (I908572,I908614,I908764);
DFFARX1 I_53247 (I731265,I3563,I908580,I908804,);
nor I_53248 (I908563,I908804,I908674);
nor I_53249 (I908554,I908804,I908730);
nand I_53250 (I908840,I731259,I731247);
and I_53251 (I908857,I908840,I731244);
DFFARX1 I_53252 (I908857,I3563,I908580,I908883,);
not I_53253 (I908891,I908883);
nand I_53254 (I908908,I908891,I908804);
nand I_53255 (I908557,I908891,I908713);
nor I_53256 (I908939,I731262,I731247);
and I_53257 (I908956,I908804,I908939);
nor I_53258 (I908973,I908891,I908956);
DFFARX1 I_53259 (I908973,I3563,I908580,I908566,);
nor I_53260 (I909004,I908606,I908939);
DFFARX1 I_53261 (I909004,I3563,I908580,I908551,);
nor I_53262 (I909035,I908883,I908939);
not I_53263 (I909052,I909035);
nand I_53264 (I908560,I909052,I908908);
not I_53265 (I909107,I3570);
DFFARX1 I_53266 (I409746,I3563,I909107,I909133,);
not I_53267 (I909141,I909133);
nand I_53268 (I909158,I409737,I409737);
and I_53269 (I909175,I909158,I409755);
DFFARX1 I_53270 (I909175,I3563,I909107,I909201,);
DFFARX1 I_53271 (I909201,I3563,I909107,I909096,);
DFFARX1 I_53272 (I409758,I3563,I909107,I909232,);
nand I_53273 (I909240,I909232,I409740);
not I_53274 (I909257,I909240);
DFFARX1 I_53275 (I909257,I3563,I909107,I909283,);
not I_53276 (I909291,I909283);
nor I_53277 (I909099,I909141,I909291);
DFFARX1 I_53278 (I409752,I3563,I909107,I909331,);
nor I_53279 (I909090,I909331,I909201);
nor I_53280 (I909081,I909331,I909257);
nand I_53281 (I909367,I409764,I409743);
and I_53282 (I909384,I909367,I409749);
DFFARX1 I_53283 (I909384,I3563,I909107,I909410,);
not I_53284 (I909418,I909410);
nand I_53285 (I909435,I909418,I909331);
nand I_53286 (I909084,I909418,I909240);
nor I_53287 (I909466,I409761,I409743);
and I_53288 (I909483,I909331,I909466);
nor I_53289 (I909500,I909418,I909483);
DFFARX1 I_53290 (I909500,I3563,I909107,I909093,);
nor I_53291 (I909531,I909133,I909466);
DFFARX1 I_53292 (I909531,I3563,I909107,I909078,);
nor I_53293 (I909562,I909410,I909466);
not I_53294 (I909579,I909562);
nand I_53295 (I909087,I909579,I909435);
not I_53296 (I909634,I3570);
DFFARX1 I_53297 (I101993,I3563,I909634,I909660,);
not I_53298 (I909668,I909660);
nand I_53299 (I909685,I101969,I101978);
and I_53300 (I909702,I909685,I101972);
DFFARX1 I_53301 (I909702,I3563,I909634,I909728,);
DFFARX1 I_53302 (I909728,I3563,I909634,I909623,);
DFFARX1 I_53303 (I101990,I3563,I909634,I909759,);
nand I_53304 (I909767,I909759,I101981);
not I_53305 (I909784,I909767);
DFFARX1 I_53306 (I909784,I3563,I909634,I909810,);
not I_53307 (I909818,I909810);
nor I_53308 (I909626,I909668,I909818);
DFFARX1 I_53309 (I101975,I3563,I909634,I909858,);
nor I_53310 (I909617,I909858,I909728);
nor I_53311 (I909608,I909858,I909784);
nand I_53312 (I909894,I101987,I101984);
and I_53313 (I909911,I909894,I101972);
DFFARX1 I_53314 (I909911,I3563,I909634,I909937,);
not I_53315 (I909945,I909937);
nand I_53316 (I909962,I909945,I909858);
nand I_53317 (I909611,I909945,I909767);
nor I_53318 (I909993,I101969,I101984);
and I_53319 (I910010,I909858,I909993);
nor I_53320 (I910027,I909945,I910010);
DFFARX1 I_53321 (I910027,I3563,I909634,I909620,);
nor I_53322 (I910058,I909660,I909993);
DFFARX1 I_53323 (I910058,I3563,I909634,I909605,);
nor I_53324 (I910089,I909937,I909993);
not I_53325 (I910106,I910089);
nand I_53326 (I909614,I910106,I909962);
not I_53327 (I910161,I3570);
DFFARX1 I_53328 (I989814,I3563,I910161,I910187,);
not I_53329 (I910195,I910187);
nand I_53330 (I910212,I989829,I989811);
and I_53331 (I910229,I910212,I989811);
DFFARX1 I_53332 (I910229,I3563,I910161,I910255,);
DFFARX1 I_53333 (I910255,I3563,I910161,I910150,);
DFFARX1 I_53334 (I989820,I3563,I910161,I910286,);
nand I_53335 (I910294,I910286,I989838);
not I_53336 (I910311,I910294);
DFFARX1 I_53337 (I910311,I3563,I910161,I910337,);
not I_53338 (I910345,I910337);
nor I_53339 (I910153,I910195,I910345);
DFFARX1 I_53340 (I989835,I3563,I910161,I910385,);
nor I_53341 (I910144,I910385,I910255);
nor I_53342 (I910135,I910385,I910311);
nand I_53343 (I910421,I989832,I989823);
and I_53344 (I910438,I910421,I989817);
DFFARX1 I_53345 (I910438,I3563,I910161,I910464,);
not I_53346 (I910472,I910464);
nand I_53347 (I910489,I910472,I910385);
nand I_53348 (I910138,I910472,I910294);
nor I_53349 (I910520,I989826,I989823);
and I_53350 (I910537,I910385,I910520);
nor I_53351 (I910554,I910472,I910537);
DFFARX1 I_53352 (I910554,I3563,I910161,I910147,);
nor I_53353 (I910585,I910187,I910520);
DFFARX1 I_53354 (I910585,I3563,I910161,I910132,);
nor I_53355 (I910616,I910464,I910520);
not I_53356 (I910633,I910616);
nand I_53357 (I910141,I910633,I910489);
not I_53358 (I910688,I3570);
DFFARX1 I_53359 (I1067986,I3563,I910688,I910714,);
not I_53360 (I910722,I910714);
nand I_53361 (I910739,I1067995,I1067983);
and I_53362 (I910756,I910739,I1067980);
DFFARX1 I_53363 (I910756,I3563,I910688,I910782,);
DFFARX1 I_53364 (I910782,I3563,I910688,I910677,);
DFFARX1 I_53365 (I1067980,I3563,I910688,I910813,);
nand I_53366 (I910821,I910813,I1067977);
not I_53367 (I910838,I910821);
DFFARX1 I_53368 (I910838,I3563,I910688,I910864,);
not I_53369 (I910872,I910864);
nor I_53370 (I910680,I910722,I910872);
DFFARX1 I_53371 (I1067983,I3563,I910688,I910912,);
nor I_53372 (I910671,I910912,I910782);
nor I_53373 (I910662,I910912,I910838);
nand I_53374 (I910948,I1067998,I1067989);
and I_53375 (I910965,I910948,I1067992);
DFFARX1 I_53376 (I910965,I3563,I910688,I910991,);
not I_53377 (I910999,I910991);
nand I_53378 (I911016,I910999,I910912);
nand I_53379 (I910665,I910999,I910821);
nor I_53380 (I911047,I1067977,I1067989);
and I_53381 (I911064,I910912,I911047);
nor I_53382 (I911081,I910999,I911064);
DFFARX1 I_53383 (I911081,I3563,I910688,I910674,);
nor I_53384 (I911112,I910714,I911047);
DFFARX1 I_53385 (I911112,I3563,I910688,I910659,);
nor I_53386 (I911143,I910991,I911047);
not I_53387 (I911160,I911143);
nand I_53388 (I910668,I911160,I911016);
not I_53389 (I911215,I3570);
DFFARX1 I_53390 (I398152,I3563,I911215,I911241,);
not I_53391 (I911249,I911241);
nand I_53392 (I911266,I398143,I398143);
and I_53393 (I911283,I911266,I398161);
DFFARX1 I_53394 (I911283,I3563,I911215,I911309,);
DFFARX1 I_53395 (I911309,I3563,I911215,I911204,);
DFFARX1 I_53396 (I398164,I3563,I911215,I911340,);
nand I_53397 (I911348,I911340,I398146);
not I_53398 (I911365,I911348);
DFFARX1 I_53399 (I911365,I3563,I911215,I911391,);
not I_53400 (I911399,I911391);
nor I_53401 (I911207,I911249,I911399);
DFFARX1 I_53402 (I398158,I3563,I911215,I911439,);
nor I_53403 (I911198,I911439,I911309);
nor I_53404 (I911189,I911439,I911365);
nand I_53405 (I911475,I398170,I398149);
and I_53406 (I911492,I911475,I398155);
DFFARX1 I_53407 (I911492,I3563,I911215,I911518,);
not I_53408 (I911526,I911518);
nand I_53409 (I911543,I911526,I911439);
nand I_53410 (I911192,I911526,I911348);
nor I_53411 (I911574,I398167,I398149);
and I_53412 (I911591,I911439,I911574);
nor I_53413 (I911608,I911526,I911591);
DFFARX1 I_53414 (I911608,I3563,I911215,I911201,);
nor I_53415 (I911639,I911241,I911574);
DFFARX1 I_53416 (I911639,I3563,I911215,I911186,);
nor I_53417 (I911670,I911518,I911574);
not I_53418 (I911687,I911670);
nand I_53419 (I911195,I911687,I911543);
not I_53420 (I911742,I3570);
DFFARX1 I_53421 (I611610,I3563,I911742,I911768,);
not I_53422 (I911776,I911768);
nand I_53423 (I911793,I611595,I611616);
and I_53424 (I911810,I911793,I611604);
DFFARX1 I_53425 (I911810,I3563,I911742,I911836,);
DFFARX1 I_53426 (I911836,I3563,I911742,I911731,);
DFFARX1 I_53427 (I611598,I3563,I911742,I911867,);
nand I_53428 (I911875,I911867,I611607);
not I_53429 (I911892,I911875);
DFFARX1 I_53430 (I911892,I3563,I911742,I911918,);
not I_53431 (I911926,I911918);
nor I_53432 (I911734,I911776,I911926);
DFFARX1 I_53433 (I611613,I3563,I911742,I911966,);
nor I_53434 (I911725,I911966,I911836);
nor I_53435 (I911716,I911966,I911892);
nand I_53436 (I912002,I611595,I611598);
and I_53437 (I912019,I912002,I611619);
DFFARX1 I_53438 (I912019,I3563,I911742,I912045,);
not I_53439 (I912053,I912045);
nand I_53440 (I912070,I912053,I911966);
nand I_53441 (I911719,I912053,I911875);
nor I_53442 (I912101,I611601,I611598);
and I_53443 (I912118,I911966,I912101);
nor I_53444 (I912135,I912053,I912118);
DFFARX1 I_53445 (I912135,I3563,I911742,I911728,);
nor I_53446 (I912166,I911768,I912101);
DFFARX1 I_53447 (I912166,I3563,I911742,I911713,);
nor I_53448 (I912197,I912045,I912101);
not I_53449 (I912214,I912197);
nand I_53450 (I911722,I912214,I912070);
not I_53451 (I912269,I3570);
DFFARX1 I_53452 (I1014362,I3563,I912269,I912295,);
not I_53453 (I912303,I912295);
nand I_53454 (I912320,I1014377,I1014359);
and I_53455 (I912337,I912320,I1014359);
DFFARX1 I_53456 (I912337,I3563,I912269,I912363,);
DFFARX1 I_53457 (I912363,I3563,I912269,I912258,);
DFFARX1 I_53458 (I1014368,I3563,I912269,I912394,);
nand I_53459 (I912402,I912394,I1014386);
not I_53460 (I912419,I912402);
DFFARX1 I_53461 (I912419,I3563,I912269,I912445,);
not I_53462 (I912453,I912445);
nor I_53463 (I912261,I912303,I912453);
DFFARX1 I_53464 (I1014383,I3563,I912269,I912493,);
nor I_53465 (I912252,I912493,I912363);
nor I_53466 (I912243,I912493,I912419);
nand I_53467 (I912529,I1014380,I1014371);
and I_53468 (I912546,I912529,I1014365);
DFFARX1 I_53469 (I912546,I3563,I912269,I912572,);
not I_53470 (I912580,I912572);
nand I_53471 (I912597,I912580,I912493);
nand I_53472 (I912246,I912580,I912402);
nor I_53473 (I912628,I1014374,I1014371);
and I_53474 (I912645,I912493,I912628);
nor I_53475 (I912662,I912580,I912645);
DFFARX1 I_53476 (I912662,I3563,I912269,I912255,);
nor I_53477 (I912693,I912295,I912628);
DFFARX1 I_53478 (I912693,I3563,I912269,I912240,);
nor I_53479 (I912724,I912572,I912628);
not I_53480 (I912741,I912724);
nand I_53481 (I912249,I912741,I912597);
not I_53482 (I912796,I3570);
DFFARX1 I_53483 (I532262,I3563,I912796,I912822,);
not I_53484 (I912830,I912822);
nand I_53485 (I912847,I532280,I532271);
and I_53486 (I912864,I912847,I532274);
DFFARX1 I_53487 (I912864,I3563,I912796,I912890,);
DFFARX1 I_53488 (I912890,I3563,I912796,I912785,);
DFFARX1 I_53489 (I532268,I3563,I912796,I912921,);
nand I_53490 (I912929,I912921,I532259);
not I_53491 (I912946,I912929);
DFFARX1 I_53492 (I912946,I3563,I912796,I912972,);
not I_53493 (I912980,I912972);
nor I_53494 (I912788,I912830,I912980);
DFFARX1 I_53495 (I532265,I3563,I912796,I913020,);
nor I_53496 (I912779,I913020,I912890);
nor I_53497 (I912770,I913020,I912946);
nand I_53498 (I913056,I532259,I532256);
and I_53499 (I913073,I913056,I532277);
DFFARX1 I_53500 (I913073,I3563,I912796,I913099,);
not I_53501 (I913107,I913099);
nand I_53502 (I913124,I913107,I913020);
nand I_53503 (I912773,I913107,I912929);
nor I_53504 (I913155,I532256,I532256);
and I_53505 (I913172,I913020,I913155);
nor I_53506 (I913189,I913107,I913172);
DFFARX1 I_53507 (I913189,I3563,I912796,I912782,);
nor I_53508 (I913220,I912822,I913155);
DFFARX1 I_53509 (I913220,I3563,I912796,I912767,);
nor I_53510 (I913251,I913099,I913155);
not I_53511 (I913268,I913251);
nand I_53512 (I912776,I913268,I913124);
not I_53513 (I913323,I3570);
DFFARX1 I_53514 (I560822,I3563,I913323,I913349,);
not I_53515 (I913357,I913349);
nand I_53516 (I913374,I560840,I560831);
and I_53517 (I913391,I913374,I560834);
DFFARX1 I_53518 (I913391,I3563,I913323,I913417,);
DFFARX1 I_53519 (I913417,I3563,I913323,I913312,);
DFFARX1 I_53520 (I560828,I3563,I913323,I913448,);
nand I_53521 (I913456,I913448,I560819);
not I_53522 (I913473,I913456);
DFFARX1 I_53523 (I913473,I3563,I913323,I913499,);
not I_53524 (I913507,I913499);
nor I_53525 (I913315,I913357,I913507);
DFFARX1 I_53526 (I560825,I3563,I913323,I913547,);
nor I_53527 (I913306,I913547,I913417);
nor I_53528 (I913297,I913547,I913473);
nand I_53529 (I913583,I560819,I560816);
and I_53530 (I913600,I913583,I560837);
DFFARX1 I_53531 (I913600,I3563,I913323,I913626,);
not I_53532 (I913634,I913626);
nand I_53533 (I913651,I913634,I913547);
nand I_53534 (I913300,I913634,I913456);
nor I_53535 (I913682,I560816,I560816);
and I_53536 (I913699,I913547,I913682);
nor I_53537 (I913716,I913634,I913699);
DFFARX1 I_53538 (I913716,I3563,I913323,I913309,);
nor I_53539 (I913747,I913349,I913682);
DFFARX1 I_53540 (I913747,I3563,I913323,I913294,);
nor I_53541 (I913778,I913626,I913682);
not I_53542 (I913795,I913778);
nand I_53543 (I913303,I913795,I913651);
not I_53544 (I913850,I3570);
DFFARX1 I_53545 (I1192163,I3563,I913850,I913876,);
not I_53546 (I913884,I913876);
nand I_53547 (I913901,I1192145,I1192145);
and I_53548 (I913918,I913901,I1192151);
DFFARX1 I_53549 (I913918,I3563,I913850,I913944,);
DFFARX1 I_53550 (I913944,I3563,I913850,I913839,);
DFFARX1 I_53551 (I1192148,I3563,I913850,I913975,);
nand I_53552 (I913983,I913975,I1192157);
not I_53553 (I914000,I913983);
DFFARX1 I_53554 (I914000,I3563,I913850,I914026,);
not I_53555 (I914034,I914026);
nor I_53556 (I913842,I913884,I914034);
DFFARX1 I_53557 (I1192169,I3563,I913850,I914074,);
nor I_53558 (I913833,I914074,I913944);
nor I_53559 (I913824,I914074,I914000);
nand I_53560 (I914110,I1192160,I1192154);
and I_53561 (I914127,I914110,I1192148);
DFFARX1 I_53562 (I914127,I3563,I913850,I914153,);
not I_53563 (I914161,I914153);
nand I_53564 (I914178,I914161,I914074);
nand I_53565 (I913827,I914161,I913983);
nor I_53566 (I914209,I1192166,I1192154);
and I_53567 (I914226,I914074,I914209);
nor I_53568 (I914243,I914161,I914226);
DFFARX1 I_53569 (I914243,I3563,I913850,I913836,);
nor I_53570 (I914274,I913876,I914209);
DFFARX1 I_53571 (I914274,I3563,I913850,I913821,);
nor I_53572 (I914305,I914153,I914209);
not I_53573 (I914322,I914305);
nand I_53574 (I913830,I914322,I914178);
not I_53575 (I914377,I3570);
DFFARX1 I_53576 (I675175,I3563,I914377,I914403,);
not I_53577 (I914411,I914403);
nand I_53578 (I914428,I675178,I675175);
and I_53579 (I914445,I914428,I675187);
DFFARX1 I_53580 (I914445,I3563,I914377,I914471,);
DFFARX1 I_53581 (I914471,I3563,I914377,I914366,);
DFFARX1 I_53582 (I675184,I3563,I914377,I914502,);
nand I_53583 (I914510,I914502,I675190);
not I_53584 (I914527,I914510);
DFFARX1 I_53585 (I914527,I3563,I914377,I914553,);
not I_53586 (I914561,I914553);
nor I_53587 (I914369,I914411,I914561);
DFFARX1 I_53588 (I675199,I3563,I914377,I914601,);
nor I_53589 (I914360,I914601,I914471);
nor I_53590 (I914351,I914601,I914527);
nand I_53591 (I914637,I675193,I675181);
and I_53592 (I914654,I914637,I675178);
DFFARX1 I_53593 (I914654,I3563,I914377,I914680,);
not I_53594 (I914688,I914680);
nand I_53595 (I914705,I914688,I914601);
nand I_53596 (I914354,I914688,I914510);
nor I_53597 (I914736,I675196,I675181);
and I_53598 (I914753,I914601,I914736);
nor I_53599 (I914770,I914688,I914753);
DFFARX1 I_53600 (I914770,I3563,I914377,I914363,);
nor I_53601 (I914801,I914403,I914736);
DFFARX1 I_53602 (I914801,I3563,I914377,I914348,);
nor I_53603 (I914832,I914680,I914736);
not I_53604 (I914849,I914832);
nand I_53605 (I914357,I914849,I914705);
not I_53606 (I914910,I3570);
DFFARX1 I_53607 (I1321286,I3563,I914910,I914936,);
DFFARX1 I_53608 (I1321280,I3563,I914910,I914953,);
not I_53609 (I914961,I914953);
not I_53610 (I914978,I1321289);
nor I_53611 (I914995,I914978,I1321301);
not I_53612 (I915012,I1321283);
nor I_53613 (I915029,I914995,I1321280);
nor I_53614 (I915046,I914953,I915029);
DFFARX1 I_53615 (I915046,I3563,I914910,I914896,);
nor I_53616 (I915077,I1321280,I1321301);
nand I_53617 (I915094,I915077,I1321289);
DFFARX1 I_53618 (I915094,I3563,I914910,I914899,);
nor I_53619 (I915125,I915012,I1321280);
nand I_53620 (I915142,I915125,I1321277);
nor I_53621 (I915159,I914936,I915142);
DFFARX1 I_53622 (I915159,I3563,I914910,I914875,);
not I_53623 (I915190,I915142);
nand I_53624 (I914887,I914953,I915190);
DFFARX1 I_53625 (I915142,I3563,I914910,I915230,);
not I_53626 (I915238,I915230);
not I_53627 (I915255,I1321280);
not I_53628 (I915272,I1321298);
nor I_53629 (I915289,I915272,I1321283);
nor I_53630 (I914902,I915238,I915289);
nor I_53631 (I915320,I915272,I1321292);
and I_53632 (I915337,I915320,I1321277);
or I_53633 (I915354,I915337,I1321295);
DFFARX1 I_53634 (I915354,I3563,I914910,I915380,);
nor I_53635 (I914890,I915380,I914936);
not I_53636 (I915402,I915380);
and I_53637 (I915419,I915402,I914936);
nor I_53638 (I914884,I914961,I915419);
nand I_53639 (I915450,I915402,I915012);
nor I_53640 (I914878,I915272,I915450);
nand I_53641 (I914881,I915402,I915190);
nand I_53642 (I915495,I915012,I1321298);
nor I_53643 (I914893,I915255,I915495);
not I_53644 (I915556,I3570);
DFFARX1 I_53645 (I317512,I3563,I915556,I915582,);
DFFARX1 I_53646 (I317518,I3563,I915556,I915599,);
not I_53647 (I915607,I915599);
not I_53648 (I915624,I317539);
nor I_53649 (I915641,I915624,I317527);
not I_53650 (I915658,I317536);
nor I_53651 (I915675,I915641,I317521);
nor I_53652 (I915692,I915599,I915675);
DFFARX1 I_53653 (I915692,I3563,I915556,I915542,);
nor I_53654 (I915723,I317521,I317527);
nand I_53655 (I915740,I915723,I317539);
DFFARX1 I_53656 (I915740,I3563,I915556,I915545,);
nor I_53657 (I915771,I915658,I317521);
nand I_53658 (I915788,I915771,I317512);
nor I_53659 (I915805,I915582,I915788);
DFFARX1 I_53660 (I915805,I3563,I915556,I915521,);
not I_53661 (I915836,I915788);
nand I_53662 (I915533,I915599,I915836);
DFFARX1 I_53663 (I915788,I3563,I915556,I915876,);
not I_53664 (I915884,I915876);
not I_53665 (I915901,I317521);
not I_53666 (I915918,I317524);
nor I_53667 (I915935,I915918,I317536);
nor I_53668 (I915548,I915884,I915935);
nor I_53669 (I915966,I915918,I317533);
and I_53670 (I915983,I915966,I317515);
or I_53671 (I916000,I915983,I317530);
DFFARX1 I_53672 (I916000,I3563,I915556,I916026,);
nor I_53673 (I915536,I916026,I915582);
not I_53674 (I916048,I916026);
and I_53675 (I916065,I916048,I915582);
nor I_53676 (I915530,I915607,I916065);
nand I_53677 (I916096,I916048,I915658);
nor I_53678 (I915524,I915918,I916096);
nand I_53679 (I915527,I916048,I915836);
nand I_53680 (I916141,I915658,I317524);
nor I_53681 (I915539,I915901,I916141);
not I_53682 (I916202,I3570);
DFFARX1 I_53683 (I583854,I3563,I916202,I916228,);
DFFARX1 I_53684 (I583866,I3563,I916202,I916245,);
not I_53685 (I916253,I916245);
not I_53686 (I916270,I583875);
nor I_53687 (I916287,I916270,I583851);
not I_53688 (I916304,I583869);
nor I_53689 (I916321,I916287,I583863);
nor I_53690 (I916338,I916245,I916321);
DFFARX1 I_53691 (I916338,I3563,I916202,I916188,);
nor I_53692 (I916369,I583863,I583851);
nand I_53693 (I916386,I916369,I583875);
DFFARX1 I_53694 (I916386,I3563,I916202,I916191,);
nor I_53695 (I916417,I916304,I583863);
nand I_53696 (I916434,I916417,I583857);
nor I_53697 (I916451,I916228,I916434);
DFFARX1 I_53698 (I916451,I3563,I916202,I916167,);
not I_53699 (I916482,I916434);
nand I_53700 (I916179,I916245,I916482);
DFFARX1 I_53701 (I916434,I3563,I916202,I916522,);
not I_53702 (I916530,I916522);
not I_53703 (I916547,I583863);
not I_53704 (I916564,I583872);
nor I_53705 (I916581,I916564,I583869);
nor I_53706 (I916194,I916530,I916581);
nor I_53707 (I916612,I916564,I583854);
and I_53708 (I916629,I916612,I583851);
or I_53709 (I916646,I916629,I583860);
DFFARX1 I_53710 (I916646,I3563,I916202,I916672,);
nor I_53711 (I916182,I916672,I916228);
not I_53712 (I916694,I916672);
and I_53713 (I916711,I916694,I916228);
nor I_53714 (I916176,I916253,I916711);
nand I_53715 (I916742,I916694,I916304);
nor I_53716 (I916170,I916564,I916742);
nand I_53717 (I916173,I916694,I916482);
nand I_53718 (I916787,I916304,I583872);
nor I_53719 (I916185,I916547,I916787);
not I_53720 (I916848,I3570);
DFFARX1 I_53721 (I760725,I3563,I916848,I916874,);
DFFARX1 I_53722 (I760719,I3563,I916848,I916891,);
not I_53723 (I916899,I916891);
not I_53724 (I916916,I760734);
nor I_53725 (I916933,I916916,I760719);
not I_53726 (I916950,I760728);
nor I_53727 (I916967,I916933,I760737);
nor I_53728 (I916984,I916891,I916967);
DFFARX1 I_53729 (I916984,I3563,I916848,I916834,);
nor I_53730 (I917015,I760737,I760719);
nand I_53731 (I917032,I917015,I760734);
DFFARX1 I_53732 (I917032,I3563,I916848,I916837,);
nor I_53733 (I917063,I916950,I760737);
nand I_53734 (I917080,I917063,I760722);
nor I_53735 (I917097,I916874,I917080);
DFFARX1 I_53736 (I917097,I3563,I916848,I916813,);
not I_53737 (I917128,I917080);
nand I_53738 (I916825,I916891,I917128);
DFFARX1 I_53739 (I917080,I3563,I916848,I917168,);
not I_53740 (I917176,I917168);
not I_53741 (I917193,I760737);
not I_53742 (I917210,I760731);
nor I_53743 (I917227,I917210,I760728);
nor I_53744 (I916840,I917176,I917227);
nor I_53745 (I917258,I917210,I760740);
and I_53746 (I917275,I917258,I760743);
or I_53747 (I917292,I917275,I760722);
DFFARX1 I_53748 (I917292,I3563,I916848,I917318,);
nor I_53749 (I916828,I917318,I916874);
not I_53750 (I917340,I917318);
and I_53751 (I917357,I917340,I916874);
nor I_53752 (I916822,I916899,I917357);
nand I_53753 (I917388,I917340,I916950);
nor I_53754 (I916816,I917210,I917388);
nand I_53755 (I916819,I917340,I917128);
nand I_53756 (I917433,I916950,I760731);
nor I_53757 (I916831,I917193,I917433);
not I_53758 (I917494,I3570);
DFFARX1 I_53759 (I742229,I3563,I917494,I917520,);
DFFARX1 I_53760 (I742223,I3563,I917494,I917537,);
not I_53761 (I917545,I917537);
not I_53762 (I917562,I742238);
nor I_53763 (I917579,I917562,I742223);
not I_53764 (I917596,I742232);
nor I_53765 (I917613,I917579,I742241);
nor I_53766 (I917630,I917537,I917613);
DFFARX1 I_53767 (I917630,I3563,I917494,I917480,);
nor I_53768 (I917661,I742241,I742223);
nand I_53769 (I917678,I917661,I742238);
DFFARX1 I_53770 (I917678,I3563,I917494,I917483,);
nor I_53771 (I917709,I917596,I742241);
nand I_53772 (I917726,I917709,I742226);
nor I_53773 (I917743,I917520,I917726);
DFFARX1 I_53774 (I917743,I3563,I917494,I917459,);
not I_53775 (I917774,I917726);
nand I_53776 (I917471,I917537,I917774);
DFFARX1 I_53777 (I917726,I3563,I917494,I917814,);
not I_53778 (I917822,I917814);
not I_53779 (I917839,I742241);
not I_53780 (I917856,I742235);
nor I_53781 (I917873,I917856,I742232);
nor I_53782 (I917486,I917822,I917873);
nor I_53783 (I917904,I917856,I742244);
and I_53784 (I917921,I917904,I742247);
or I_53785 (I917938,I917921,I742226);
DFFARX1 I_53786 (I917938,I3563,I917494,I917964,);
nor I_53787 (I917474,I917964,I917520);
not I_53788 (I917986,I917964);
and I_53789 (I918003,I917986,I917520);
nor I_53790 (I917468,I917545,I918003);
nand I_53791 (I918034,I917986,I917596);
nor I_53792 (I917462,I917856,I918034);
nand I_53793 (I917465,I917986,I917774);
nand I_53794 (I918079,I917596,I742235);
nor I_53795 (I917477,I917839,I918079);
not I_53796 (I918140,I3570);
DFFARX1 I_53797 (I1407688,I3563,I918140,I918166,);
DFFARX1 I_53798 (I1407712,I3563,I918140,I918183,);
not I_53799 (I918191,I918183);
not I_53800 (I918208,I1407694);
nor I_53801 (I918225,I918208,I1407703);
not I_53802 (I918242,I1407688);
nor I_53803 (I918259,I918225,I1407709);
nor I_53804 (I918276,I918183,I918259);
DFFARX1 I_53805 (I918276,I3563,I918140,I918126,);
nor I_53806 (I918307,I1407709,I1407703);
nand I_53807 (I918324,I918307,I1407694);
DFFARX1 I_53808 (I918324,I3563,I918140,I918129,);
nor I_53809 (I918355,I918242,I1407709);
nand I_53810 (I918372,I918355,I1407706);
nor I_53811 (I918389,I918166,I918372);
DFFARX1 I_53812 (I918389,I3563,I918140,I918105,);
not I_53813 (I918420,I918372);
nand I_53814 (I918117,I918183,I918420);
DFFARX1 I_53815 (I918372,I3563,I918140,I918460,);
not I_53816 (I918468,I918460);
not I_53817 (I918485,I1407709);
not I_53818 (I918502,I1407700);
nor I_53819 (I918519,I918502,I1407688);
nor I_53820 (I918132,I918468,I918519);
nor I_53821 (I918550,I918502,I1407691);
and I_53822 (I918567,I918550,I1407715);
or I_53823 (I918584,I918567,I1407697);
DFFARX1 I_53824 (I918584,I3563,I918140,I918610,);
nor I_53825 (I918120,I918610,I918166);
not I_53826 (I918632,I918610);
and I_53827 (I918649,I918632,I918166);
nor I_53828 (I918114,I918191,I918649);
nand I_53829 (I918680,I918632,I918242);
nor I_53830 (I918108,I918502,I918680);
nand I_53831 (I918111,I918632,I918420);
nand I_53832 (I918725,I918242,I1407700);
nor I_53833 (I918123,I918485,I918725);
not I_53834 (I918786,I3570);
DFFARX1 I_53835 (I1330338,I3563,I918786,I918812,);
DFFARX1 I_53836 (I1330362,I3563,I918786,I918829,);
not I_53837 (I918837,I918829);
not I_53838 (I918854,I1330344);
nor I_53839 (I918871,I918854,I1330353);
not I_53840 (I918888,I1330338);
nor I_53841 (I918905,I918871,I1330359);
nor I_53842 (I918922,I918829,I918905);
DFFARX1 I_53843 (I918922,I3563,I918786,I918772,);
nor I_53844 (I918953,I1330359,I1330353);
nand I_53845 (I918970,I918953,I1330344);
DFFARX1 I_53846 (I918970,I3563,I918786,I918775,);
nor I_53847 (I919001,I918888,I1330359);
nand I_53848 (I919018,I919001,I1330356);
nor I_53849 (I919035,I918812,I919018);
DFFARX1 I_53850 (I919035,I3563,I918786,I918751,);
not I_53851 (I919066,I919018);
nand I_53852 (I918763,I918829,I919066);
DFFARX1 I_53853 (I919018,I3563,I918786,I919106,);
not I_53854 (I919114,I919106);
not I_53855 (I919131,I1330359);
not I_53856 (I919148,I1330350);
nor I_53857 (I919165,I919148,I1330338);
nor I_53858 (I918778,I919114,I919165);
nor I_53859 (I919196,I919148,I1330341);
and I_53860 (I919213,I919196,I1330365);
or I_53861 (I919230,I919213,I1330347);
DFFARX1 I_53862 (I919230,I3563,I918786,I919256,);
nor I_53863 (I918766,I919256,I918812);
not I_53864 (I919278,I919256);
and I_53865 (I919295,I919278,I918812);
nor I_53866 (I918760,I918837,I919295);
nand I_53867 (I919326,I919278,I918888);
nor I_53868 (I918754,I919148,I919326);
nand I_53869 (I918757,I919278,I919066);
nand I_53870 (I919371,I918888,I1330350);
nor I_53871 (I918769,I919131,I919371);
not I_53872 (I919432,I3570);
DFFARX1 I_53873 (I416061,I3563,I919432,I919458,);
DFFARX1 I_53874 (I416067,I3563,I919432,I919475,);
not I_53875 (I919483,I919475);
not I_53876 (I919500,I416088);
nor I_53877 (I919517,I919500,I416076);
not I_53878 (I919534,I416085);
nor I_53879 (I919551,I919517,I416070);
nor I_53880 (I919568,I919475,I919551);
DFFARX1 I_53881 (I919568,I3563,I919432,I919418,);
nor I_53882 (I919599,I416070,I416076);
nand I_53883 (I919616,I919599,I416088);
DFFARX1 I_53884 (I919616,I3563,I919432,I919421,);
nor I_53885 (I919647,I919534,I416070);
nand I_53886 (I919664,I919647,I416061);
nor I_53887 (I919681,I919458,I919664);
DFFARX1 I_53888 (I919681,I3563,I919432,I919397,);
not I_53889 (I919712,I919664);
nand I_53890 (I919409,I919475,I919712);
DFFARX1 I_53891 (I919664,I3563,I919432,I919752,);
not I_53892 (I919760,I919752);
not I_53893 (I919777,I416070);
not I_53894 (I919794,I416073);
nor I_53895 (I919811,I919794,I416085);
nor I_53896 (I919424,I919760,I919811);
nor I_53897 (I919842,I919794,I416082);
and I_53898 (I919859,I919842,I416064);
or I_53899 (I919876,I919859,I416079);
DFFARX1 I_53900 (I919876,I3563,I919432,I919902,);
nor I_53901 (I919412,I919902,I919458);
not I_53902 (I919924,I919902);
and I_53903 (I919941,I919924,I919458);
nor I_53904 (I919406,I919483,I919941);
nand I_53905 (I919972,I919924,I919534);
nor I_53906 (I919400,I919794,I919972);
nand I_53907 (I919403,I919924,I919712);
nand I_53908 (I920017,I919534,I416073);
nor I_53909 (I919415,I919777,I920017);
not I_53910 (I920078,I3570);
DFFARX1 I_53911 (I266059,I3563,I920078,I920104,);
DFFARX1 I_53912 (I266071,I3563,I920078,I920121,);
not I_53913 (I920129,I920121);
not I_53914 (I920146,I266077);
nor I_53915 (I920163,I920146,I266062);
not I_53916 (I920180,I266053);
nor I_53917 (I920197,I920163,I266074);
nor I_53918 (I920214,I920121,I920197);
DFFARX1 I_53919 (I920214,I3563,I920078,I920064,);
nor I_53920 (I920245,I266074,I266062);
nand I_53921 (I920262,I920245,I266077);
DFFARX1 I_53922 (I920262,I3563,I920078,I920067,);
nor I_53923 (I920293,I920180,I266074);
nand I_53924 (I920310,I920293,I266056);
nor I_53925 (I920327,I920104,I920310);
DFFARX1 I_53926 (I920327,I3563,I920078,I920043,);
not I_53927 (I920358,I920310);
nand I_53928 (I920055,I920121,I920358);
DFFARX1 I_53929 (I920310,I3563,I920078,I920398,);
not I_53930 (I920406,I920398);
not I_53931 (I920423,I266074);
not I_53932 (I920440,I266065);
nor I_53933 (I920457,I920440,I266053);
nor I_53934 (I920070,I920406,I920457);
nor I_53935 (I920488,I920440,I266068);
and I_53936 (I920505,I920488,I266056);
or I_53937 (I920522,I920505,I266053);
DFFARX1 I_53938 (I920522,I3563,I920078,I920548,);
nor I_53939 (I920058,I920548,I920104);
not I_53940 (I920570,I920548);
and I_53941 (I920587,I920570,I920104);
nor I_53942 (I920052,I920129,I920587);
nand I_53943 (I920618,I920570,I920180);
nor I_53944 (I920046,I920440,I920618);
nand I_53945 (I920049,I920570,I920358);
nand I_53946 (I920663,I920180,I266065);
nor I_53947 (I920061,I920423,I920663);
not I_53948 (I920724,I3570);
DFFARX1 I_53949 (I668823,I3563,I920724,I920750,);
DFFARX1 I_53950 (I668817,I3563,I920724,I920767,);
not I_53951 (I920775,I920767);
not I_53952 (I920792,I668832);
nor I_53953 (I920809,I920792,I668817);
not I_53954 (I920826,I668826);
nor I_53955 (I920843,I920809,I668835);
nor I_53956 (I920860,I920767,I920843);
DFFARX1 I_53957 (I920860,I3563,I920724,I920710,);
nor I_53958 (I920891,I668835,I668817);
nand I_53959 (I920908,I920891,I668832);
DFFARX1 I_53960 (I920908,I3563,I920724,I920713,);
nor I_53961 (I920939,I920826,I668835);
nand I_53962 (I920956,I920939,I668820);
nor I_53963 (I920973,I920750,I920956);
DFFARX1 I_53964 (I920973,I3563,I920724,I920689,);
not I_53965 (I921004,I920956);
nand I_53966 (I920701,I920767,I921004);
DFFARX1 I_53967 (I920956,I3563,I920724,I921044,);
not I_53968 (I921052,I921044);
not I_53969 (I921069,I668835);
not I_53970 (I921086,I668829);
nor I_53971 (I921103,I921086,I668826);
nor I_53972 (I920716,I921052,I921103);
nor I_53973 (I921134,I921086,I668838);
and I_53974 (I921151,I921134,I668841);
or I_53975 (I921168,I921151,I668820);
DFFARX1 I_53976 (I921168,I3563,I920724,I921194,);
nor I_53977 (I920704,I921194,I920750);
not I_53978 (I921216,I921194);
and I_53979 (I921233,I921216,I920750);
nor I_53980 (I920698,I920775,I921233);
nand I_53981 (I921264,I921216,I920826);
nor I_53982 (I920692,I921086,I921264);
nand I_53983 (I920695,I921216,I921004);
nand I_53984 (I921309,I920826,I668829);
nor I_53985 (I920707,I921069,I921309);
not I_53986 (I921370,I3570);
DFFARX1 I_53987 (I848479,I3563,I921370,I921396,);
DFFARX1 I_53988 (I848476,I3563,I921370,I921413,);
not I_53989 (I921421,I921413);
not I_53990 (I921438,I848476);
nor I_53991 (I921455,I921438,I848479);
not I_53992 (I921472,I848491);
nor I_53993 (I921489,I921455,I848485);
nor I_53994 (I921506,I921413,I921489);
DFFARX1 I_53995 (I921506,I3563,I921370,I921356,);
nor I_53996 (I921537,I848485,I848479);
nand I_53997 (I921554,I921537,I848476);
DFFARX1 I_53998 (I921554,I3563,I921370,I921359,);
nor I_53999 (I921585,I921472,I848485);
nand I_54000 (I921602,I921585,I848473);
nor I_54001 (I921619,I921396,I921602);
DFFARX1 I_54002 (I921619,I3563,I921370,I921335,);
not I_54003 (I921650,I921602);
nand I_54004 (I921347,I921413,I921650);
DFFARX1 I_54005 (I921602,I3563,I921370,I921690,);
not I_54006 (I921698,I921690);
not I_54007 (I921715,I848485);
not I_54008 (I921732,I848482);
nor I_54009 (I921749,I921732,I848491);
nor I_54010 (I921362,I921698,I921749);
nor I_54011 (I921780,I921732,I848488);
and I_54012 (I921797,I921780,I848494);
or I_54013 (I921814,I921797,I848473);
DFFARX1 I_54014 (I921814,I3563,I921370,I921840,);
nor I_54015 (I921350,I921840,I921396);
not I_54016 (I921862,I921840);
and I_54017 (I921879,I921862,I921396);
nor I_54018 (I921344,I921421,I921879);
nand I_54019 (I921910,I921862,I921472);
nor I_54020 (I921338,I921732,I921910);
nand I_54021 (I921341,I921862,I921650);
nand I_54022 (I921955,I921472,I848482);
nor I_54023 (I921353,I921715,I921955);
not I_54024 (I922016,I3570);
DFFARX1 I_54025 (I1254587,I3563,I922016,I922042,);
DFFARX1 I_54026 (I1254593,I3563,I922016,I922059,);
not I_54027 (I922067,I922059);
not I_54028 (I922084,I1254590);
nor I_54029 (I922101,I922084,I1254569);
not I_54030 (I922118,I1254572);
nor I_54031 (I922135,I922101,I1254578);
nor I_54032 (I922152,I922059,I922135);
DFFARX1 I_54033 (I922152,I3563,I922016,I922002,);
nor I_54034 (I922183,I1254578,I1254569);
nand I_54035 (I922200,I922183,I1254590);
DFFARX1 I_54036 (I922200,I3563,I922016,I922005,);
nor I_54037 (I922231,I922118,I1254578);
nand I_54038 (I922248,I922231,I1254572);
nor I_54039 (I922265,I922042,I922248);
DFFARX1 I_54040 (I922265,I3563,I922016,I921981,);
not I_54041 (I922296,I922248);
nand I_54042 (I921993,I922059,I922296);
DFFARX1 I_54043 (I922248,I3563,I922016,I922336,);
not I_54044 (I922344,I922336);
not I_54045 (I922361,I1254578);
not I_54046 (I922378,I1254581);
nor I_54047 (I922395,I922378,I1254572);
nor I_54048 (I922008,I922344,I922395);
nor I_54049 (I922426,I922378,I1254569);
and I_54050 (I922443,I922426,I1254575);
or I_54051 (I922460,I922443,I1254584);
DFFARX1 I_54052 (I922460,I3563,I922016,I922486,);
nor I_54053 (I921996,I922486,I922042);
not I_54054 (I922508,I922486);
and I_54055 (I922525,I922508,I922042);
nor I_54056 (I921990,I922067,I922525);
nand I_54057 (I922556,I922508,I922118);
nor I_54058 (I921984,I922378,I922556);
nand I_54059 (I921987,I922508,I922296);
nand I_54060 (I922601,I922118,I1254581);
nor I_54061 (I921999,I922361,I922601);
not I_54062 (I922662,I3570);
DFFARX1 I_54063 (I514344,I3563,I922662,I922688,);
DFFARX1 I_54064 (I514341,I3563,I922662,I922705,);
not I_54065 (I922713,I922705);
not I_54066 (I922730,I514356);
nor I_54067 (I922747,I922730,I514359);
not I_54068 (I922764,I514347);
nor I_54069 (I922781,I922747,I514353);
nor I_54070 (I922798,I922705,I922781);
DFFARX1 I_54071 (I922798,I3563,I922662,I922648,);
nor I_54072 (I922829,I514353,I514359);
nand I_54073 (I922846,I922829,I514356);
DFFARX1 I_54074 (I922846,I3563,I922662,I922651,);
nor I_54075 (I922877,I922764,I514353);
nand I_54076 (I922894,I922877,I514365);
nor I_54077 (I922911,I922688,I922894);
DFFARX1 I_54078 (I922911,I3563,I922662,I922627,);
not I_54079 (I922942,I922894);
nand I_54080 (I922639,I922705,I922942);
DFFARX1 I_54081 (I922894,I3563,I922662,I922982,);
not I_54082 (I922990,I922982);
not I_54083 (I923007,I514353);
not I_54084 (I923024,I514338);
nor I_54085 (I923041,I923024,I514347);
nor I_54086 (I922654,I922990,I923041);
nor I_54087 (I923072,I923024,I514350);
and I_54088 (I923089,I923072,I514338);
or I_54089 (I923106,I923089,I514362);
DFFARX1 I_54090 (I923106,I3563,I922662,I923132,);
nor I_54091 (I922642,I923132,I922688);
not I_54092 (I923154,I923132);
and I_54093 (I923171,I923154,I922688);
nor I_54094 (I922636,I922713,I923171);
nand I_54095 (I923202,I923154,I922764);
nor I_54096 (I922630,I923024,I923202);
nand I_54097 (I922633,I923154,I922942);
nand I_54098 (I923247,I922764,I514338);
nor I_54099 (I922645,I923007,I923247);
not I_54100 (I923308,I3570);
DFFARX1 I_54101 (I809855,I3563,I923308,I923334,);
DFFARX1 I_54102 (I809849,I3563,I923308,I923351,);
not I_54103 (I923359,I923351);
not I_54104 (I923376,I809864);
nor I_54105 (I923393,I923376,I809849);
not I_54106 (I923410,I809858);
nor I_54107 (I923427,I923393,I809867);
nor I_54108 (I923444,I923351,I923427);
DFFARX1 I_54109 (I923444,I3563,I923308,I923294,);
nor I_54110 (I923475,I809867,I809849);
nand I_54111 (I923492,I923475,I809864);
DFFARX1 I_54112 (I923492,I3563,I923308,I923297,);
nor I_54113 (I923523,I923410,I809867);
nand I_54114 (I923540,I923523,I809852);
nor I_54115 (I923557,I923334,I923540);
DFFARX1 I_54116 (I923557,I3563,I923308,I923273,);
not I_54117 (I923588,I923540);
nand I_54118 (I923285,I923351,I923588);
DFFARX1 I_54119 (I923540,I3563,I923308,I923628,);
not I_54120 (I923636,I923628);
not I_54121 (I923653,I809867);
not I_54122 (I923670,I809861);
nor I_54123 (I923687,I923670,I809858);
nor I_54124 (I923300,I923636,I923687);
nor I_54125 (I923718,I923670,I809870);
and I_54126 (I923735,I923718,I809873);
or I_54127 (I923752,I923735,I809852);
DFFARX1 I_54128 (I923752,I3563,I923308,I923778,);
nor I_54129 (I923288,I923778,I923334);
not I_54130 (I923800,I923778);
and I_54131 (I923817,I923800,I923334);
nor I_54132 (I923282,I923359,I923817);
nand I_54133 (I923848,I923800,I923410);
nor I_54134 (I923276,I923670,I923848);
nand I_54135 (I923279,I923800,I923588);
nand I_54136 (I923893,I923410,I809861);
nor I_54137 (I923291,I923653,I923893);
not I_54138 (I923954,I3570);
DFFARX1 I_54139 (I1099105,I3563,I923954,I923980,);
DFFARX1 I_54140 (I1099087,I3563,I923954,I923997,);
not I_54141 (I924005,I923997);
not I_54142 (I924022,I1099096);
nor I_54143 (I924039,I924022,I1099108);
not I_54144 (I924056,I1099090);
nor I_54145 (I924073,I924039,I1099099);
nor I_54146 (I924090,I923997,I924073);
DFFARX1 I_54147 (I924090,I3563,I923954,I923940,);
nor I_54148 (I924121,I1099099,I1099108);
nand I_54149 (I924138,I924121,I1099096);
DFFARX1 I_54150 (I924138,I3563,I923954,I923943,);
nor I_54151 (I924169,I924056,I1099099);
nand I_54152 (I924186,I924169,I1099111);
nor I_54153 (I924203,I923980,I924186);
DFFARX1 I_54154 (I924203,I3563,I923954,I923919,);
not I_54155 (I924234,I924186);
nand I_54156 (I923931,I923997,I924234);
DFFARX1 I_54157 (I924186,I3563,I923954,I924274,);
not I_54158 (I924282,I924274);
not I_54159 (I924299,I1099099);
not I_54160 (I924316,I1099087);
nor I_54161 (I924333,I924316,I1099090);
nor I_54162 (I923946,I924282,I924333);
nor I_54163 (I924364,I924316,I1099093);
and I_54164 (I924381,I924364,I1099102);
or I_54165 (I924398,I924381,I1099090);
DFFARX1 I_54166 (I924398,I3563,I923954,I924424,);
nor I_54167 (I923934,I924424,I923980);
not I_54168 (I924446,I924424);
and I_54169 (I924463,I924446,I923980);
nor I_54170 (I923928,I924005,I924463);
nand I_54171 (I924494,I924446,I924056);
nor I_54172 (I923922,I924316,I924494);
nand I_54173 (I923925,I924446,I924234);
nand I_54174 (I924539,I924056,I1099087);
nor I_54175 (I923937,I924299,I924539);
not I_54176 (I924600,I3570);
DFFARX1 I_54177 (I830561,I3563,I924600,I924626,);
DFFARX1 I_54178 (I830558,I3563,I924600,I924643,);
not I_54179 (I924651,I924643);
not I_54180 (I924668,I830558);
nor I_54181 (I924685,I924668,I830561);
not I_54182 (I924702,I830573);
nor I_54183 (I924719,I924685,I830567);
nor I_54184 (I924736,I924643,I924719);
DFFARX1 I_54185 (I924736,I3563,I924600,I924586,);
nor I_54186 (I924767,I830567,I830561);
nand I_54187 (I924784,I924767,I830558);
DFFARX1 I_54188 (I924784,I3563,I924600,I924589,);
nor I_54189 (I924815,I924702,I830567);
nand I_54190 (I924832,I924815,I830555);
nor I_54191 (I924849,I924626,I924832);
DFFARX1 I_54192 (I924849,I3563,I924600,I924565,);
not I_54193 (I924880,I924832);
nand I_54194 (I924577,I924643,I924880);
DFFARX1 I_54195 (I924832,I3563,I924600,I924920,);
not I_54196 (I924928,I924920);
not I_54197 (I924945,I830567);
not I_54198 (I924962,I830564);
nor I_54199 (I924979,I924962,I830573);
nor I_54200 (I924592,I924928,I924979);
nor I_54201 (I925010,I924962,I830570);
and I_54202 (I925027,I925010,I830576);
or I_54203 (I925044,I925027,I830555);
DFFARX1 I_54204 (I925044,I3563,I924600,I925070,);
nor I_54205 (I924580,I925070,I924626);
not I_54206 (I925092,I925070);
and I_54207 (I925109,I925092,I924626);
nor I_54208 (I924574,I924651,I925109);
nand I_54209 (I925140,I925092,I924702);
nor I_54210 (I924568,I924962,I925140);
nand I_54211 (I924571,I925092,I924880);
nand I_54212 (I925185,I924702,I830564);
nor I_54213 (I924583,I924945,I925185);
not I_54214 (I925246,I3570);
DFFARX1 I_54215 (I710439,I3563,I925246,I925272,);
DFFARX1 I_54216 (I710433,I3563,I925246,I925289,);
not I_54217 (I925297,I925289);
not I_54218 (I925314,I710448);
nor I_54219 (I925331,I925314,I710433);
not I_54220 (I925348,I710442);
nor I_54221 (I925365,I925331,I710451);
nor I_54222 (I925382,I925289,I925365);
DFFARX1 I_54223 (I925382,I3563,I925246,I925232,);
nor I_54224 (I925413,I710451,I710433);
nand I_54225 (I925430,I925413,I710448);
DFFARX1 I_54226 (I925430,I3563,I925246,I925235,);
nor I_54227 (I925461,I925348,I710451);
nand I_54228 (I925478,I925461,I710436);
nor I_54229 (I925495,I925272,I925478);
DFFARX1 I_54230 (I925495,I3563,I925246,I925211,);
not I_54231 (I925526,I925478);
nand I_54232 (I925223,I925289,I925526);
DFFARX1 I_54233 (I925478,I3563,I925246,I925566,);
not I_54234 (I925574,I925566);
not I_54235 (I925591,I710451);
not I_54236 (I925608,I710445);
nor I_54237 (I925625,I925608,I710442);
nor I_54238 (I925238,I925574,I925625);
nor I_54239 (I925656,I925608,I710454);
and I_54240 (I925673,I925656,I710457);
or I_54241 (I925690,I925673,I710436);
DFFARX1 I_54242 (I925690,I3563,I925246,I925716,);
nor I_54243 (I925226,I925716,I925272);
not I_54244 (I925738,I925716);
and I_54245 (I925755,I925738,I925272);
nor I_54246 (I925220,I925297,I925755);
nand I_54247 (I925786,I925738,I925348);
nor I_54248 (I925214,I925608,I925786);
nand I_54249 (I925217,I925738,I925526);
nand I_54250 (I925831,I925348,I710445);
nor I_54251 (I925229,I925591,I925831);
not I_54252 (I925892,I3570);
DFFARX1 I_54253 (I140967,I3563,I925892,I925918,);
DFFARX1 I_54254 (I140973,I3563,I925892,I925935,);
not I_54255 (I925943,I925935);
not I_54256 (I925960,I140991);
nor I_54257 (I925977,I925960,I140970);
not I_54258 (I925994,I140976);
nor I_54259 (I926011,I925977,I140982);
nor I_54260 (I926028,I925935,I926011);
DFFARX1 I_54261 (I926028,I3563,I925892,I925878,);
nor I_54262 (I926059,I140982,I140970);
nand I_54263 (I926076,I926059,I140991);
DFFARX1 I_54264 (I926076,I3563,I925892,I925881,);
nor I_54265 (I926107,I925994,I140982);
nand I_54266 (I926124,I926107,I140988);
nor I_54267 (I926141,I925918,I926124);
DFFARX1 I_54268 (I926141,I3563,I925892,I925857,);
not I_54269 (I926172,I926124);
nand I_54270 (I925869,I925935,I926172);
DFFARX1 I_54271 (I926124,I3563,I925892,I926212,);
not I_54272 (I926220,I926212);
not I_54273 (I926237,I140982);
not I_54274 (I926254,I140970);
nor I_54275 (I926271,I926254,I140976);
nor I_54276 (I925884,I926220,I926271);
nor I_54277 (I926302,I926254,I140979);
and I_54278 (I926319,I926302,I140967);
or I_54279 (I926336,I926319,I140985);
DFFARX1 I_54280 (I926336,I3563,I925892,I926362,);
nor I_54281 (I925872,I926362,I925918);
not I_54282 (I926384,I926362);
and I_54283 (I926401,I926384,I925918);
nor I_54284 (I925866,I925943,I926401);
nand I_54285 (I926432,I926384,I925994);
nor I_54286 (I925860,I926254,I926432);
nand I_54287 (I925863,I926384,I926172);
nand I_54288 (I926477,I925994,I140970);
nor I_54289 (I925875,I926237,I926477);
not I_54290 (I926538,I3570);
DFFARX1 I_54291 (I50850,I3563,I926538,I926564,);
DFFARX1 I_54292 (I50856,I3563,I926538,I926581,);
not I_54293 (I926589,I926581);
not I_54294 (I926606,I50850);
nor I_54295 (I926623,I926606,I50862);
not I_54296 (I926640,I50874);
nor I_54297 (I926657,I926623,I50868);
nor I_54298 (I926674,I926581,I926657);
DFFARX1 I_54299 (I926674,I3563,I926538,I926524,);
nor I_54300 (I926705,I50868,I50862);
nand I_54301 (I926722,I926705,I50850);
DFFARX1 I_54302 (I926722,I3563,I926538,I926527,);
nor I_54303 (I926753,I926640,I50868);
nand I_54304 (I926770,I926753,I50853);
nor I_54305 (I926787,I926564,I926770);
DFFARX1 I_54306 (I926787,I3563,I926538,I926503,);
not I_54307 (I926818,I926770);
nand I_54308 (I926515,I926581,I926818);
DFFARX1 I_54309 (I926770,I3563,I926538,I926858,);
not I_54310 (I926866,I926858);
not I_54311 (I926883,I50868);
not I_54312 (I926900,I50853);
nor I_54313 (I926917,I926900,I50874);
nor I_54314 (I926530,I926866,I926917);
nor I_54315 (I926948,I926900,I50871);
and I_54316 (I926965,I926948,I50865);
or I_54317 (I926982,I926965,I50859);
DFFARX1 I_54318 (I926982,I3563,I926538,I927008,);
nor I_54319 (I926518,I927008,I926564);
not I_54320 (I927030,I927008);
and I_54321 (I927047,I927030,I926564);
nor I_54322 (I926512,I926589,I927047);
nand I_54323 (I927078,I927030,I926640);
nor I_54324 (I926506,I926900,I927078);
nand I_54325 (I926509,I927030,I926818);
nand I_54326 (I927123,I926640,I50853);
nor I_54327 (I926521,I926883,I927123);
not I_54328 (I927184,I3570);
DFFARX1 I_54329 (I902760,I3563,I927184,I927210,);
DFFARX1 I_54330 (I902757,I3563,I927184,I927227,);
not I_54331 (I927235,I927227);
not I_54332 (I927252,I902757);
nor I_54333 (I927269,I927252,I902760);
not I_54334 (I927286,I902772);
nor I_54335 (I927303,I927269,I902766);
nor I_54336 (I927320,I927227,I927303);
DFFARX1 I_54337 (I927320,I3563,I927184,I927170,);
nor I_54338 (I927351,I902766,I902760);
nand I_54339 (I927368,I927351,I902757);
DFFARX1 I_54340 (I927368,I3563,I927184,I927173,);
nor I_54341 (I927399,I927286,I902766);
nand I_54342 (I927416,I927399,I902754);
nor I_54343 (I927433,I927210,I927416);
DFFARX1 I_54344 (I927433,I3563,I927184,I927149,);
not I_54345 (I927464,I927416);
nand I_54346 (I927161,I927227,I927464);
DFFARX1 I_54347 (I927416,I3563,I927184,I927504,);
not I_54348 (I927512,I927504);
not I_54349 (I927529,I902766);
not I_54350 (I927546,I902763);
nor I_54351 (I927563,I927546,I902772);
nor I_54352 (I927176,I927512,I927563);
nor I_54353 (I927594,I927546,I902769);
and I_54354 (I927611,I927594,I902775);
or I_54355 (I927628,I927611,I902754);
DFFARX1 I_54356 (I927628,I3563,I927184,I927654,);
nor I_54357 (I927164,I927654,I927210);
not I_54358 (I927676,I927654);
and I_54359 (I927693,I927676,I927210);
nor I_54360 (I927158,I927235,I927693);
nand I_54361 (I927724,I927676,I927286);
nor I_54362 (I927152,I927546,I927724);
nand I_54363 (I927155,I927676,I927464);
nand I_54364 (I927769,I927286,I902763);
nor I_54365 (I927167,I927529,I927769);
not I_54366 (I927830,I3570);
DFFARX1 I_54367 (I846898,I3563,I927830,I927856,);
DFFARX1 I_54368 (I846895,I3563,I927830,I927873,);
not I_54369 (I927881,I927873);
not I_54370 (I927898,I846895);
nor I_54371 (I927915,I927898,I846898);
not I_54372 (I927932,I846910);
nor I_54373 (I927949,I927915,I846904);
nor I_54374 (I927966,I927873,I927949);
DFFARX1 I_54375 (I927966,I3563,I927830,I927816,);
nor I_54376 (I927997,I846904,I846898);
nand I_54377 (I928014,I927997,I846895);
DFFARX1 I_54378 (I928014,I3563,I927830,I927819,);
nor I_54379 (I928045,I927932,I846904);
nand I_54380 (I928062,I928045,I846892);
nor I_54381 (I928079,I927856,I928062);
DFFARX1 I_54382 (I928079,I3563,I927830,I927795,);
not I_54383 (I928110,I928062);
nand I_54384 (I927807,I927873,I928110);
DFFARX1 I_54385 (I928062,I3563,I927830,I928150,);
not I_54386 (I928158,I928150);
not I_54387 (I928175,I846904);
not I_54388 (I928192,I846901);
nor I_54389 (I928209,I928192,I846910);
nor I_54390 (I927822,I928158,I928209);
nor I_54391 (I928240,I928192,I846907);
and I_54392 (I928257,I928240,I846913);
or I_54393 (I928274,I928257,I846892);
DFFARX1 I_54394 (I928274,I3563,I927830,I928300,);
nor I_54395 (I927810,I928300,I927856);
not I_54396 (I928322,I928300);
and I_54397 (I928339,I928322,I927856);
nor I_54398 (I927804,I927881,I928339);
nand I_54399 (I928370,I928322,I927932);
nor I_54400 (I927798,I928192,I928370);
nand I_54401 (I927801,I928322,I928110);
nand I_54402 (I928415,I927932,I846901);
nor I_54403 (I927813,I928175,I928415);
not I_54404 (I928476,I3570);
DFFARX1 I_54405 (I828453,I3563,I928476,I928502,);
DFFARX1 I_54406 (I828450,I3563,I928476,I928519,);
not I_54407 (I928527,I928519);
not I_54408 (I928544,I828450);
nor I_54409 (I928561,I928544,I828453);
not I_54410 (I928578,I828465);
nor I_54411 (I928595,I928561,I828459);
nor I_54412 (I928612,I928519,I928595);
DFFARX1 I_54413 (I928612,I3563,I928476,I928462,);
nor I_54414 (I928643,I828459,I828453);
nand I_54415 (I928660,I928643,I828450);
DFFARX1 I_54416 (I928660,I3563,I928476,I928465,);
nor I_54417 (I928691,I928578,I828459);
nand I_54418 (I928708,I928691,I828447);
nor I_54419 (I928725,I928502,I928708);
DFFARX1 I_54420 (I928725,I3563,I928476,I928441,);
not I_54421 (I928756,I928708);
nand I_54422 (I928453,I928519,I928756);
DFFARX1 I_54423 (I928708,I3563,I928476,I928796,);
not I_54424 (I928804,I928796);
not I_54425 (I928821,I828459);
not I_54426 (I928838,I828456);
nor I_54427 (I928855,I928838,I828465);
nor I_54428 (I928468,I928804,I928855);
nor I_54429 (I928886,I928838,I828462);
and I_54430 (I928903,I928886,I828468);
or I_54431 (I928920,I928903,I828447);
DFFARX1 I_54432 (I928920,I3563,I928476,I928946,);
nor I_54433 (I928456,I928946,I928502);
not I_54434 (I928968,I928946);
and I_54435 (I928985,I928968,I928502);
nor I_54436 (I928450,I928527,I928985);
nand I_54437 (I929016,I928968,I928578);
nor I_54438 (I928444,I928838,I929016);
nand I_54439 (I928447,I928968,I928756);
nand I_54440 (I929061,I928578,I828456);
nor I_54441 (I928459,I928821,I929061);
not I_54442 (I929122,I3570);
DFFARX1 I_54443 (I157831,I3563,I929122,I929148,);
DFFARX1 I_54444 (I157837,I3563,I929122,I929165,);
not I_54445 (I929173,I929165);
not I_54446 (I929190,I157855);
nor I_54447 (I929207,I929190,I157834);
not I_54448 (I929224,I157840);
nor I_54449 (I929241,I929207,I157846);
nor I_54450 (I929258,I929165,I929241);
DFFARX1 I_54451 (I929258,I3563,I929122,I929108,);
nor I_54452 (I929289,I157846,I157834);
nand I_54453 (I929306,I929289,I157855);
DFFARX1 I_54454 (I929306,I3563,I929122,I929111,);
nor I_54455 (I929337,I929224,I157846);
nand I_54456 (I929354,I929337,I157852);
nor I_54457 (I929371,I929148,I929354);
DFFARX1 I_54458 (I929371,I3563,I929122,I929087,);
not I_54459 (I929402,I929354);
nand I_54460 (I929099,I929165,I929402);
DFFARX1 I_54461 (I929354,I3563,I929122,I929442,);
not I_54462 (I929450,I929442);
not I_54463 (I929467,I157846);
not I_54464 (I929484,I157834);
nor I_54465 (I929501,I929484,I157840);
nor I_54466 (I929114,I929450,I929501);
nor I_54467 (I929532,I929484,I157843);
and I_54468 (I929549,I929532,I157831);
or I_54469 (I929566,I929549,I157849);
DFFARX1 I_54470 (I929566,I3563,I929122,I929592,);
nor I_54471 (I929102,I929592,I929148);
not I_54472 (I929614,I929592);
and I_54473 (I929631,I929614,I929148);
nor I_54474 (I929096,I929173,I929631);
nand I_54475 (I929662,I929614,I929224);
nor I_54476 (I929090,I929484,I929662);
nand I_54477 (I929093,I929614,I929402);
nand I_54478 (I929707,I929224,I157834);
nor I_54479 (I929105,I929467,I929707);
not I_54480 (I929768,I3570);
DFFARX1 I_54481 (I1230889,I3563,I929768,I929794,);
DFFARX1 I_54482 (I1230871,I3563,I929768,I929811,);
not I_54483 (I929819,I929811);
not I_54484 (I929836,I1230880);
nor I_54485 (I929853,I929836,I1230892);
not I_54486 (I929870,I1230874);
nor I_54487 (I929887,I929853,I1230883);
nor I_54488 (I929904,I929811,I929887);
DFFARX1 I_54489 (I929904,I3563,I929768,I929754,);
nor I_54490 (I929935,I1230883,I1230892);
nand I_54491 (I929952,I929935,I1230880);
DFFARX1 I_54492 (I929952,I3563,I929768,I929757,);
nor I_54493 (I929983,I929870,I1230883);
nand I_54494 (I930000,I929983,I1230895);
nor I_54495 (I930017,I929794,I930000);
DFFARX1 I_54496 (I930017,I3563,I929768,I929733,);
not I_54497 (I930048,I930000);
nand I_54498 (I929745,I929811,I930048);
DFFARX1 I_54499 (I930000,I3563,I929768,I930088,);
not I_54500 (I930096,I930088);
not I_54501 (I930113,I1230883);
not I_54502 (I930130,I1230871);
nor I_54503 (I930147,I930130,I1230874);
nor I_54504 (I929760,I930096,I930147);
nor I_54505 (I930178,I930130,I1230877);
and I_54506 (I930195,I930178,I1230886);
or I_54507 (I930212,I930195,I1230874);
DFFARX1 I_54508 (I930212,I3563,I929768,I930238,);
nor I_54509 (I929748,I930238,I929794);
not I_54510 (I930260,I930238);
and I_54511 (I930277,I930260,I929794);
nor I_54512 (I929742,I929819,I930277);
nand I_54513 (I930308,I930260,I929870);
nor I_54514 (I929736,I930130,I930308);
nand I_54515 (I929739,I930260,I930048);
nand I_54516 (I930353,I929870,I1230871);
nor I_54517 (I929751,I930113,I930353);
not I_54518 (I930414,I3570);
DFFARX1 I_54519 (I780955,I3563,I930414,I930440,);
DFFARX1 I_54520 (I780949,I3563,I930414,I930457,);
not I_54521 (I930465,I930457);
not I_54522 (I930482,I780964);
nor I_54523 (I930499,I930482,I780949);
not I_54524 (I930516,I780958);
nor I_54525 (I930533,I930499,I780967);
nor I_54526 (I930550,I930457,I930533);
DFFARX1 I_54527 (I930550,I3563,I930414,I930400,);
nor I_54528 (I930581,I780967,I780949);
nand I_54529 (I930598,I930581,I780964);
DFFARX1 I_54530 (I930598,I3563,I930414,I930403,);
nor I_54531 (I930629,I930516,I780967);
nand I_54532 (I930646,I930629,I780952);
nor I_54533 (I930663,I930440,I930646);
DFFARX1 I_54534 (I930663,I3563,I930414,I930379,);
not I_54535 (I930694,I930646);
nand I_54536 (I930391,I930457,I930694);
DFFARX1 I_54537 (I930646,I3563,I930414,I930734,);
not I_54538 (I930742,I930734);
not I_54539 (I930759,I780967);
not I_54540 (I930776,I780961);
nor I_54541 (I930793,I930776,I780958);
nor I_54542 (I930406,I930742,I930793);
nor I_54543 (I930824,I930776,I780970);
and I_54544 (I930841,I930824,I780973);
or I_54545 (I930858,I930841,I780952);
DFFARX1 I_54546 (I930858,I3563,I930414,I930884,);
nor I_54547 (I930394,I930884,I930440);
not I_54548 (I930906,I930884);
and I_54549 (I930923,I930906,I930440);
nor I_54550 (I930388,I930465,I930923);
nand I_54551 (I930954,I930906,I930516);
nor I_54552 (I930382,I930776,I930954);
nand I_54553 (I930385,I930906,I930694);
nand I_54554 (I930999,I930516,I780961);
nor I_54555 (I930397,I930759,I930999);
not I_54556 (I931060,I3570);
DFFARX1 I_54557 (I1156327,I3563,I931060,I931086,);
DFFARX1 I_54558 (I1156309,I3563,I931060,I931103,);
not I_54559 (I931111,I931103);
not I_54560 (I931128,I1156318);
nor I_54561 (I931145,I931128,I1156330);
not I_54562 (I931162,I1156312);
nor I_54563 (I931179,I931145,I1156321);
nor I_54564 (I931196,I931103,I931179);
DFFARX1 I_54565 (I931196,I3563,I931060,I931046,);
nor I_54566 (I931227,I1156321,I1156330);
nand I_54567 (I931244,I931227,I1156318);
DFFARX1 I_54568 (I931244,I3563,I931060,I931049,);
nor I_54569 (I931275,I931162,I1156321);
nand I_54570 (I931292,I931275,I1156333);
nor I_54571 (I931309,I931086,I931292);
DFFARX1 I_54572 (I931309,I3563,I931060,I931025,);
not I_54573 (I931340,I931292);
nand I_54574 (I931037,I931103,I931340);
DFFARX1 I_54575 (I931292,I3563,I931060,I931380,);
not I_54576 (I931388,I931380);
not I_54577 (I931405,I1156321);
not I_54578 (I931422,I1156309);
nor I_54579 (I931439,I931422,I1156312);
nor I_54580 (I931052,I931388,I931439);
nor I_54581 (I931470,I931422,I1156315);
and I_54582 (I931487,I931470,I1156324);
or I_54583 (I931504,I931487,I1156312);
DFFARX1 I_54584 (I931504,I3563,I931060,I931530,);
nor I_54585 (I931040,I931530,I931086);
not I_54586 (I931552,I931530);
and I_54587 (I931569,I931552,I931086);
nor I_54588 (I931034,I931111,I931569);
nand I_54589 (I931600,I931552,I931162);
nor I_54590 (I931028,I931422,I931600);
nand I_54591 (I931031,I931552,I931340);
nand I_54592 (I931645,I931162,I1156309);
nor I_54593 (I931043,I931405,I931645);
not I_54594 (I931706,I3570);
DFFARX1 I_54595 (I108820,I3563,I931706,I931732,);
DFFARX1 I_54596 (I108826,I3563,I931706,I931749,);
not I_54597 (I931757,I931749);
not I_54598 (I931774,I108844);
nor I_54599 (I931791,I931774,I108823);
not I_54600 (I931808,I108829);
nor I_54601 (I931825,I931791,I108835);
nor I_54602 (I931842,I931749,I931825);
DFFARX1 I_54603 (I931842,I3563,I931706,I931692,);
nor I_54604 (I931873,I108835,I108823);
nand I_54605 (I931890,I931873,I108844);
DFFARX1 I_54606 (I931890,I3563,I931706,I931695,);
nor I_54607 (I931921,I931808,I108835);
nand I_54608 (I931938,I931921,I108841);
nor I_54609 (I931955,I931732,I931938);
DFFARX1 I_54610 (I931955,I3563,I931706,I931671,);
not I_54611 (I931986,I931938);
nand I_54612 (I931683,I931749,I931986);
DFFARX1 I_54613 (I931938,I3563,I931706,I932026,);
not I_54614 (I932034,I932026);
not I_54615 (I932051,I108835);
not I_54616 (I932068,I108823);
nor I_54617 (I932085,I932068,I108829);
nor I_54618 (I931698,I932034,I932085);
nor I_54619 (I932116,I932068,I108832);
and I_54620 (I932133,I932116,I108820);
or I_54621 (I932150,I932133,I108838);
DFFARX1 I_54622 (I932150,I3563,I931706,I932176,);
nor I_54623 (I931686,I932176,I931732);
not I_54624 (I932198,I932176);
and I_54625 (I932215,I932198,I931732);
nor I_54626 (I931680,I931757,I932215);
nand I_54627 (I932246,I932198,I931808);
nor I_54628 (I931674,I932068,I932246);
nand I_54629 (I931677,I932198,I931986);
nand I_54630 (I932291,I931808,I108823);
nor I_54631 (I931689,I932051,I932291);
not I_54632 (I932352,I3570);
DFFARX1 I_54633 (I1110087,I3563,I932352,I932378,);
DFFARX1 I_54634 (I1110069,I3563,I932352,I932395,);
not I_54635 (I932403,I932395);
not I_54636 (I932420,I1110078);
nor I_54637 (I932437,I932420,I1110090);
not I_54638 (I932454,I1110072);
nor I_54639 (I932471,I932437,I1110081);
nor I_54640 (I932488,I932395,I932471);
DFFARX1 I_54641 (I932488,I3563,I932352,I932338,);
nor I_54642 (I932519,I1110081,I1110090);
nand I_54643 (I932536,I932519,I1110078);
DFFARX1 I_54644 (I932536,I3563,I932352,I932341,);
nor I_54645 (I932567,I932454,I1110081);
nand I_54646 (I932584,I932567,I1110093);
nor I_54647 (I932601,I932378,I932584);
DFFARX1 I_54648 (I932601,I3563,I932352,I932317,);
not I_54649 (I932632,I932584);
nand I_54650 (I932329,I932395,I932632);
DFFARX1 I_54651 (I932584,I3563,I932352,I932672,);
not I_54652 (I932680,I932672);
not I_54653 (I932697,I1110081);
not I_54654 (I932714,I1110069);
nor I_54655 (I932731,I932714,I1110072);
nor I_54656 (I932344,I932680,I932731);
nor I_54657 (I932762,I932714,I1110075);
and I_54658 (I932779,I932762,I1110084);
or I_54659 (I932796,I932779,I1110072);
DFFARX1 I_54660 (I932796,I3563,I932352,I932822,);
nor I_54661 (I932332,I932822,I932378);
not I_54662 (I932844,I932822);
and I_54663 (I932861,I932844,I932378);
nor I_54664 (I932326,I932403,I932861);
nand I_54665 (I932892,I932844,I932454);
nor I_54666 (I932320,I932714,I932892);
nand I_54667 (I932323,I932844,I932632);
nand I_54668 (I932937,I932454,I1110069);
nor I_54669 (I932335,I932697,I932937);
not I_54670 (I932998,I3570);
DFFARX1 I_54671 (I537019,I3563,I932998,I933024,);
DFFARX1 I_54672 (I537031,I3563,I932998,I933041,);
not I_54673 (I933049,I933041);
not I_54674 (I933066,I537016);
nor I_54675 (I933083,I933066,I537034);
not I_54676 (I933100,I537040);
nor I_54677 (I933117,I933083,I537022);
nor I_54678 (I933134,I933041,I933117);
DFFARX1 I_54679 (I933134,I3563,I932998,I932984,);
nor I_54680 (I933165,I537022,I537034);
nand I_54681 (I933182,I933165,I537016);
DFFARX1 I_54682 (I933182,I3563,I932998,I932987,);
nor I_54683 (I933213,I933100,I537022);
nand I_54684 (I933230,I933213,I537025);
nor I_54685 (I933247,I933024,I933230);
DFFARX1 I_54686 (I933247,I3563,I932998,I932963,);
not I_54687 (I933278,I933230);
nand I_54688 (I932975,I933041,I933278);
DFFARX1 I_54689 (I933230,I3563,I932998,I933318,);
not I_54690 (I933326,I933318);
not I_54691 (I933343,I537022);
not I_54692 (I933360,I537028);
nor I_54693 (I933377,I933360,I537040);
nor I_54694 (I932990,I933326,I933377);
nor I_54695 (I933408,I933360,I537037);
and I_54696 (I933425,I933408,I537016);
or I_54697 (I933442,I933425,I537019);
DFFARX1 I_54698 (I933442,I3563,I932998,I933468,);
nor I_54699 (I932978,I933468,I933024);
not I_54700 (I933490,I933468);
and I_54701 (I933507,I933490,I933024);
nor I_54702 (I932972,I933049,I933507);
nand I_54703 (I933538,I933490,I933100);
nor I_54704 (I932966,I933360,I933538);
nand I_54705 (I932969,I933490,I933278);
nand I_54706 (I933583,I933100,I537028);
nor I_54707 (I932981,I933343,I933583);
not I_54708 (I933644,I3570);
DFFARX1 I_54709 (I98807,I3563,I933644,I933670,);
DFFARX1 I_54710 (I98813,I3563,I933644,I933687,);
not I_54711 (I933695,I933687);
not I_54712 (I933712,I98831);
nor I_54713 (I933729,I933712,I98810);
not I_54714 (I933746,I98816);
nor I_54715 (I933763,I933729,I98822);
nor I_54716 (I933780,I933687,I933763);
DFFARX1 I_54717 (I933780,I3563,I933644,I933630,);
nor I_54718 (I933811,I98822,I98810);
nand I_54719 (I933828,I933811,I98831);
DFFARX1 I_54720 (I933828,I3563,I933644,I933633,);
nor I_54721 (I933859,I933746,I98822);
nand I_54722 (I933876,I933859,I98828);
nor I_54723 (I933893,I933670,I933876);
DFFARX1 I_54724 (I933893,I3563,I933644,I933609,);
not I_54725 (I933924,I933876);
nand I_54726 (I933621,I933687,I933924);
DFFARX1 I_54727 (I933876,I3563,I933644,I933964,);
not I_54728 (I933972,I933964);
not I_54729 (I933989,I98822);
not I_54730 (I934006,I98810);
nor I_54731 (I934023,I934006,I98816);
nor I_54732 (I933636,I933972,I934023);
nor I_54733 (I934054,I934006,I98819);
and I_54734 (I934071,I934054,I98807);
or I_54735 (I934088,I934071,I98825);
DFFARX1 I_54736 (I934088,I3563,I933644,I934114,);
nor I_54737 (I933624,I934114,I933670);
not I_54738 (I934136,I934114);
and I_54739 (I934153,I934136,I933670);
nor I_54740 (I933618,I933695,I934153);
nand I_54741 (I934184,I934136,I933746);
nor I_54742 (I933612,I934006,I934184);
nand I_54743 (I933615,I934136,I933924);
nand I_54744 (I934229,I933746,I98810);
nor I_54745 (I933627,I933989,I934229);
not I_54746 (I934290,I3570);
DFFARX1 I_54747 (I41364,I3563,I934290,I934316,);
DFFARX1 I_54748 (I41370,I3563,I934290,I934333,);
not I_54749 (I934341,I934333);
not I_54750 (I934358,I41364);
nor I_54751 (I934375,I934358,I41376);
not I_54752 (I934392,I41388);
nor I_54753 (I934409,I934375,I41382);
nor I_54754 (I934426,I934333,I934409);
DFFARX1 I_54755 (I934426,I3563,I934290,I934276,);
nor I_54756 (I934457,I41382,I41376);
nand I_54757 (I934474,I934457,I41364);
DFFARX1 I_54758 (I934474,I3563,I934290,I934279,);
nor I_54759 (I934505,I934392,I41382);
nand I_54760 (I934522,I934505,I41367);
nor I_54761 (I934539,I934316,I934522);
DFFARX1 I_54762 (I934539,I3563,I934290,I934255,);
not I_54763 (I934570,I934522);
nand I_54764 (I934267,I934333,I934570);
DFFARX1 I_54765 (I934522,I3563,I934290,I934610,);
not I_54766 (I934618,I934610);
not I_54767 (I934635,I41382);
not I_54768 (I934652,I41367);
nor I_54769 (I934669,I934652,I41388);
nor I_54770 (I934282,I934618,I934669);
nor I_54771 (I934700,I934652,I41385);
and I_54772 (I934717,I934700,I41379);
or I_54773 (I934734,I934717,I41373);
DFFARX1 I_54774 (I934734,I3563,I934290,I934760,);
nor I_54775 (I934270,I934760,I934316);
not I_54776 (I934782,I934760);
and I_54777 (I934799,I934782,I934316);
nor I_54778 (I934264,I934341,I934799);
nand I_54779 (I934830,I934782,I934392);
nor I_54780 (I934258,I934652,I934830);
nand I_54781 (I934261,I934782,I934570);
nand I_54782 (I934875,I934392,I41367);
nor I_54783 (I934273,I934635,I934875);
not I_54784 (I934936,I3570);
DFFARX1 I_54785 (I62444,I3563,I934936,I934962,);
DFFARX1 I_54786 (I62450,I3563,I934936,I934979,);
not I_54787 (I934987,I934979);
not I_54788 (I935004,I62468);
nor I_54789 (I935021,I935004,I62447);
not I_54790 (I935038,I62453);
nor I_54791 (I935055,I935021,I62459);
nor I_54792 (I935072,I934979,I935055);
DFFARX1 I_54793 (I935072,I3563,I934936,I934922,);
nor I_54794 (I935103,I62459,I62447);
nand I_54795 (I935120,I935103,I62468);
DFFARX1 I_54796 (I935120,I3563,I934936,I934925,);
nor I_54797 (I935151,I935038,I62459);
nand I_54798 (I935168,I935151,I62465);
nor I_54799 (I935185,I934962,I935168);
DFFARX1 I_54800 (I935185,I3563,I934936,I934901,);
not I_54801 (I935216,I935168);
nand I_54802 (I934913,I934979,I935216);
DFFARX1 I_54803 (I935168,I3563,I934936,I935256,);
not I_54804 (I935264,I935256);
not I_54805 (I935281,I62459);
not I_54806 (I935298,I62447);
nor I_54807 (I935315,I935298,I62453);
nor I_54808 (I934928,I935264,I935315);
nor I_54809 (I935346,I935298,I62456);
and I_54810 (I935363,I935346,I62444);
or I_54811 (I935380,I935363,I62462);
DFFARX1 I_54812 (I935380,I3563,I934936,I935406,);
nor I_54813 (I934916,I935406,I934962);
not I_54814 (I935428,I935406);
and I_54815 (I935445,I935428,I934962);
nor I_54816 (I934910,I934987,I935445);
nand I_54817 (I935476,I935428,I935038);
nor I_54818 (I934904,I935298,I935476);
nand I_54819 (I934907,I935428,I935216);
nand I_54820 (I935521,I935038,I62447);
nor I_54821 (I934919,I935281,I935521);
not I_54822 (I935582,I3570);
DFFARX1 I_54823 (I619112,I3563,I935582,I935608,);
DFFARX1 I_54824 (I619124,I3563,I935582,I935625,);
not I_54825 (I935633,I935625);
not I_54826 (I935650,I619133);
nor I_54827 (I935667,I935650,I619109);
not I_54828 (I935684,I619127);
nor I_54829 (I935701,I935667,I619121);
nor I_54830 (I935718,I935625,I935701);
DFFARX1 I_54831 (I935718,I3563,I935582,I935568,);
nor I_54832 (I935749,I619121,I619109);
nand I_54833 (I935766,I935749,I619133);
DFFARX1 I_54834 (I935766,I3563,I935582,I935571,);
nor I_54835 (I935797,I935684,I619121);
nand I_54836 (I935814,I935797,I619115);
nor I_54837 (I935831,I935608,I935814);
DFFARX1 I_54838 (I935831,I3563,I935582,I935547,);
not I_54839 (I935862,I935814);
nand I_54840 (I935559,I935625,I935862);
DFFARX1 I_54841 (I935814,I3563,I935582,I935902,);
not I_54842 (I935910,I935902);
not I_54843 (I935927,I619121);
not I_54844 (I935944,I619130);
nor I_54845 (I935961,I935944,I619127);
nor I_54846 (I935574,I935910,I935961);
nor I_54847 (I935992,I935944,I619112);
and I_54848 (I936009,I935992,I619109);
or I_54849 (I936026,I936009,I619118);
DFFARX1 I_54850 (I936026,I3563,I935582,I936052,);
nor I_54851 (I935562,I936052,I935608);
not I_54852 (I936074,I936052);
and I_54853 (I936091,I936074,I935608);
nor I_54854 (I935556,I935633,I936091);
nand I_54855 (I936122,I936074,I935684);
nor I_54856 (I935550,I935944,I936122);
nand I_54857 (I935553,I936074,I935862);
nand I_54858 (I936167,I935684,I619130);
nor I_54859 (I935565,I935927,I936167);
not I_54860 (I936228,I3570);
DFFARX1 I_54861 (I457224,I3563,I936228,I936254,);
DFFARX1 I_54862 (I457221,I3563,I936228,I936271,);
not I_54863 (I936279,I936271);
not I_54864 (I936296,I457236);
nor I_54865 (I936313,I936296,I457239);
not I_54866 (I936330,I457227);
nor I_54867 (I936347,I936313,I457233);
nor I_54868 (I936364,I936271,I936347);
DFFARX1 I_54869 (I936364,I3563,I936228,I936214,);
nor I_54870 (I936395,I457233,I457239);
nand I_54871 (I936412,I936395,I457236);
DFFARX1 I_54872 (I936412,I3563,I936228,I936217,);
nor I_54873 (I936443,I936330,I457233);
nand I_54874 (I936460,I936443,I457245);
nor I_54875 (I936477,I936254,I936460);
DFFARX1 I_54876 (I936477,I3563,I936228,I936193,);
not I_54877 (I936508,I936460);
nand I_54878 (I936205,I936271,I936508);
DFFARX1 I_54879 (I936460,I3563,I936228,I936548,);
not I_54880 (I936556,I936548);
not I_54881 (I936573,I457233);
not I_54882 (I936590,I457218);
nor I_54883 (I936607,I936590,I457227);
nor I_54884 (I936220,I936556,I936607);
nor I_54885 (I936638,I936590,I457230);
and I_54886 (I936655,I936638,I457218);
or I_54887 (I936672,I936655,I457242);
DFFARX1 I_54888 (I936672,I3563,I936228,I936698,);
nor I_54889 (I936208,I936698,I936254);
not I_54890 (I936720,I936698);
and I_54891 (I936737,I936720,I936254);
nor I_54892 (I936202,I936279,I936737);
nand I_54893 (I936768,I936720,I936330);
nor I_54894 (I936196,I936590,I936768);
nand I_54895 (I936199,I936720,I936508);
nand I_54896 (I936813,I936330,I457218);
nor I_54897 (I936211,I936573,I936813);
not I_54898 (I936874,I3570);
DFFARX1 I_54899 (I154142,I3563,I936874,I936900,);
DFFARX1 I_54900 (I154148,I3563,I936874,I936917,);
not I_54901 (I936925,I936917);
not I_54902 (I936942,I154166);
nor I_54903 (I936959,I936942,I154145);
not I_54904 (I936976,I154151);
nor I_54905 (I936993,I936959,I154157);
nor I_54906 (I937010,I936917,I936993);
DFFARX1 I_54907 (I937010,I3563,I936874,I936860,);
nor I_54908 (I937041,I154157,I154145);
nand I_54909 (I937058,I937041,I154166);
DFFARX1 I_54910 (I937058,I3563,I936874,I936863,);
nor I_54911 (I937089,I936976,I154157);
nand I_54912 (I937106,I937089,I154163);
nor I_54913 (I937123,I936900,I937106);
DFFARX1 I_54914 (I937123,I3563,I936874,I936839,);
not I_54915 (I937154,I937106);
nand I_54916 (I936851,I936917,I937154);
DFFARX1 I_54917 (I937106,I3563,I936874,I937194,);
not I_54918 (I937202,I937194);
not I_54919 (I937219,I154157);
not I_54920 (I937236,I154145);
nor I_54921 (I937253,I937236,I154151);
nor I_54922 (I936866,I937202,I937253);
nor I_54923 (I937284,I937236,I154154);
and I_54924 (I937301,I937284,I154142);
or I_54925 (I937318,I937301,I154160);
DFFARX1 I_54926 (I937318,I3563,I936874,I937344,);
nor I_54927 (I936854,I937344,I936900);
not I_54928 (I937366,I937344);
and I_54929 (I937383,I937366,I936900);
nor I_54930 (I936848,I936925,I937383);
nand I_54931 (I937414,I937366,I936976);
nor I_54932 (I936842,I937236,I937414);
nand I_54933 (I936845,I937366,I937154);
nand I_54934 (I937459,I936976,I154145);
nor I_54935 (I936857,I937219,I937459);
not I_54936 (I937520,I3570);
DFFARX1 I_54937 (I640498,I3563,I937520,I937546,);
DFFARX1 I_54938 (I640510,I3563,I937520,I937563,);
not I_54939 (I937571,I937563);
not I_54940 (I937588,I640519);
nor I_54941 (I937605,I937588,I640495);
not I_54942 (I937622,I640513);
nor I_54943 (I937639,I937605,I640507);
nor I_54944 (I937656,I937563,I937639);
DFFARX1 I_54945 (I937656,I3563,I937520,I937506,);
nor I_54946 (I937687,I640507,I640495);
nand I_54947 (I937704,I937687,I640519);
DFFARX1 I_54948 (I937704,I3563,I937520,I937509,);
nor I_54949 (I937735,I937622,I640507);
nand I_54950 (I937752,I937735,I640501);
nor I_54951 (I937769,I937546,I937752);
DFFARX1 I_54952 (I937769,I3563,I937520,I937485,);
not I_54953 (I937800,I937752);
nand I_54954 (I937497,I937563,I937800);
DFFARX1 I_54955 (I937752,I3563,I937520,I937840,);
not I_54956 (I937848,I937840);
not I_54957 (I937865,I640507);
not I_54958 (I937882,I640516);
nor I_54959 (I937899,I937882,I640513);
nor I_54960 (I937512,I937848,I937899);
nor I_54961 (I937930,I937882,I640498);
and I_54962 (I937947,I937930,I640495);
or I_54963 (I937964,I937947,I640504);
DFFARX1 I_54964 (I937964,I3563,I937520,I937990,);
nor I_54965 (I937500,I937990,I937546);
not I_54966 (I938012,I937990);
and I_54967 (I938029,I938012,I937546);
nor I_54968 (I937494,I937571,I938029);
nand I_54969 (I938060,I938012,I937622);
nor I_54970 (I937488,I937882,I938060);
nand I_54971 (I937491,I938012,I937800);
nand I_54972 (I938105,I937622,I640516);
nor I_54973 (I937503,I937865,I938105);
not I_54974 (I938166,I3570);
DFFARX1 I_54975 (I1208347,I3563,I938166,I938192,);
DFFARX1 I_54976 (I1208329,I3563,I938166,I938209,);
not I_54977 (I938217,I938209);
not I_54978 (I938234,I1208338);
nor I_54979 (I938251,I938234,I1208350);
not I_54980 (I938268,I1208332);
nor I_54981 (I938285,I938251,I1208341);
nor I_54982 (I938302,I938209,I938285);
DFFARX1 I_54983 (I938302,I3563,I938166,I938152,);
nor I_54984 (I938333,I1208341,I1208350);
nand I_54985 (I938350,I938333,I1208338);
DFFARX1 I_54986 (I938350,I3563,I938166,I938155,);
nor I_54987 (I938381,I938268,I1208341);
nand I_54988 (I938398,I938381,I1208353);
nor I_54989 (I938415,I938192,I938398);
DFFARX1 I_54990 (I938415,I3563,I938166,I938131,);
not I_54991 (I938446,I938398);
nand I_54992 (I938143,I938209,I938446);
DFFARX1 I_54993 (I938398,I3563,I938166,I938486,);
not I_54994 (I938494,I938486);
not I_54995 (I938511,I1208341);
not I_54996 (I938528,I1208329);
nor I_54997 (I938545,I938528,I1208332);
nor I_54998 (I938158,I938494,I938545);
nor I_54999 (I938576,I938528,I1208335);
and I_55000 (I938593,I938576,I1208344);
or I_55001 (I938610,I938593,I1208332);
DFFARX1 I_55002 (I938610,I3563,I938166,I938636,);
nor I_55003 (I938146,I938636,I938192);
not I_55004 (I938658,I938636);
and I_55005 (I938675,I938658,I938192);
nor I_55006 (I938140,I938217,I938675);
nand I_55007 (I938706,I938658,I938268);
nor I_55008 (I938134,I938528,I938706);
nand I_55009 (I938137,I938658,I938446);
nand I_55010 (I938751,I938268,I1208329);
nor I_55011 (I938149,I938511,I938751);
not I_55012 (I938812,I3570);
DFFARX1 I_55013 (I152561,I3563,I938812,I938838,);
DFFARX1 I_55014 (I152567,I3563,I938812,I938855,);
not I_55015 (I938863,I938855);
not I_55016 (I938880,I152585);
nor I_55017 (I938897,I938880,I152564);
not I_55018 (I938914,I152570);
nor I_55019 (I938931,I938897,I152576);
nor I_55020 (I938948,I938855,I938931);
DFFARX1 I_55021 (I938948,I3563,I938812,I938798,);
nor I_55022 (I938979,I152576,I152564);
nand I_55023 (I938996,I938979,I152585);
DFFARX1 I_55024 (I938996,I3563,I938812,I938801,);
nor I_55025 (I939027,I938914,I152576);
nand I_55026 (I939044,I939027,I152582);
nor I_55027 (I939061,I938838,I939044);
DFFARX1 I_55028 (I939061,I3563,I938812,I938777,);
not I_55029 (I939092,I939044);
nand I_55030 (I938789,I938855,I939092);
DFFARX1 I_55031 (I939044,I3563,I938812,I939132,);
not I_55032 (I939140,I939132);
not I_55033 (I939157,I152576);
not I_55034 (I939174,I152564);
nor I_55035 (I939191,I939174,I152570);
nor I_55036 (I938804,I939140,I939191);
nor I_55037 (I939222,I939174,I152573);
and I_55038 (I939239,I939222,I152561);
or I_55039 (I939256,I939239,I152579);
DFFARX1 I_55040 (I939256,I3563,I938812,I939282,);
nor I_55041 (I938792,I939282,I938838);
not I_55042 (I939304,I939282);
and I_55043 (I939321,I939304,I938838);
nor I_55044 (I938786,I938863,I939321);
nand I_55045 (I939352,I939304,I938914);
nor I_55046 (I938780,I939174,I939352);
nand I_55047 (I938783,I939304,I939092);
nand I_55048 (I939397,I938914,I152564);
nor I_55049 (I938795,I939157,I939397);
not I_55050 (I939458,I3570);
DFFARX1 I_55051 (I1335693,I3563,I939458,I939484,);
DFFARX1 I_55052 (I1335717,I3563,I939458,I939501,);
not I_55053 (I939509,I939501);
not I_55054 (I939526,I1335699);
nor I_55055 (I939543,I939526,I1335708);
not I_55056 (I939560,I1335693);
nor I_55057 (I939577,I939543,I1335714);
nor I_55058 (I939594,I939501,I939577);
DFFARX1 I_55059 (I939594,I3563,I939458,I939444,);
nor I_55060 (I939625,I1335714,I1335708);
nand I_55061 (I939642,I939625,I1335699);
DFFARX1 I_55062 (I939642,I3563,I939458,I939447,);
nor I_55063 (I939673,I939560,I1335714);
nand I_55064 (I939690,I939673,I1335711);
nor I_55065 (I939707,I939484,I939690);
DFFARX1 I_55066 (I939707,I3563,I939458,I939423,);
not I_55067 (I939738,I939690);
nand I_55068 (I939435,I939501,I939738);
DFFARX1 I_55069 (I939690,I3563,I939458,I939778,);
not I_55070 (I939786,I939778);
not I_55071 (I939803,I1335714);
not I_55072 (I939820,I1335705);
nor I_55073 (I939837,I939820,I1335693);
nor I_55074 (I939450,I939786,I939837);
nor I_55075 (I939868,I939820,I1335696);
and I_55076 (I939885,I939868,I1335720);
or I_55077 (I939902,I939885,I1335702);
DFFARX1 I_55078 (I939902,I3563,I939458,I939928,);
nor I_55079 (I939438,I939928,I939484);
not I_55080 (I939950,I939928);
and I_55081 (I939967,I939950,I939484);
nor I_55082 (I939432,I939509,I939967);
nand I_55083 (I939998,I939950,I939560);
nor I_55084 (I939426,I939820,I939998);
nand I_55085 (I939429,I939950,I939738);
nand I_55086 (I940043,I939560,I1335705);
nor I_55087 (I939441,I939803,I940043);
not I_55088 (I940104,I3570);
DFFARX1 I_55089 (I441992,I3563,I940104,I940130,);
DFFARX1 I_55090 (I441989,I3563,I940104,I940147,);
not I_55091 (I940155,I940147);
not I_55092 (I940172,I442004);
nor I_55093 (I940189,I940172,I442007);
not I_55094 (I940206,I441995);
nor I_55095 (I940223,I940189,I442001);
nor I_55096 (I940240,I940147,I940223);
DFFARX1 I_55097 (I940240,I3563,I940104,I940090,);
nor I_55098 (I940271,I442001,I442007);
nand I_55099 (I940288,I940271,I442004);
DFFARX1 I_55100 (I940288,I3563,I940104,I940093,);
nor I_55101 (I940319,I940206,I442001);
nand I_55102 (I940336,I940319,I442013);
nor I_55103 (I940353,I940130,I940336);
DFFARX1 I_55104 (I940353,I3563,I940104,I940069,);
not I_55105 (I940384,I940336);
nand I_55106 (I940081,I940147,I940384);
DFFARX1 I_55107 (I940336,I3563,I940104,I940424,);
not I_55108 (I940432,I940424);
not I_55109 (I940449,I442001);
not I_55110 (I940466,I441986);
nor I_55111 (I940483,I940466,I441995);
nor I_55112 (I940096,I940432,I940483);
nor I_55113 (I940514,I940466,I441998);
and I_55114 (I940531,I940514,I441986);
or I_55115 (I940548,I940531,I442010);
DFFARX1 I_55116 (I940548,I3563,I940104,I940574,);
nor I_55117 (I940084,I940574,I940130);
not I_55118 (I940596,I940574);
and I_55119 (I940613,I940596,I940130);
nor I_55120 (I940078,I940155,I940613);
nand I_55121 (I940644,I940596,I940206);
nor I_55122 (I940072,I940466,I940644);
nand I_55123 (I940075,I940596,I940384);
nand I_55124 (I940689,I940206,I441986);
nor I_55125 (I940087,I940449,I940689);
not I_55126 (I940750,I3570);
DFFARX1 I_55127 (I422408,I3563,I940750,I940776,);
DFFARX1 I_55128 (I422405,I3563,I940750,I940793,);
not I_55129 (I940801,I940793);
not I_55130 (I940818,I422420);
nor I_55131 (I940835,I940818,I422423);
not I_55132 (I940852,I422411);
nor I_55133 (I940869,I940835,I422417);
nor I_55134 (I940886,I940793,I940869);
DFFARX1 I_55135 (I940886,I3563,I940750,I940736,);
nor I_55136 (I940917,I422417,I422423);
nand I_55137 (I940934,I940917,I422420);
DFFARX1 I_55138 (I940934,I3563,I940750,I940739,);
nor I_55139 (I940965,I940852,I422417);
nand I_55140 (I940982,I940965,I422429);
nor I_55141 (I940999,I940776,I940982);
DFFARX1 I_55142 (I940999,I3563,I940750,I940715,);
not I_55143 (I941030,I940982);
nand I_55144 (I940727,I940793,I941030);
DFFARX1 I_55145 (I940982,I3563,I940750,I941070,);
not I_55146 (I941078,I941070);
not I_55147 (I941095,I422417);
not I_55148 (I941112,I422402);
nor I_55149 (I941129,I941112,I422411);
nor I_55150 (I940742,I941078,I941129);
nor I_55151 (I941160,I941112,I422414);
and I_55152 (I941177,I941160,I422402);
or I_55153 (I941194,I941177,I422426);
DFFARX1 I_55154 (I941194,I3563,I940750,I941220,);
nor I_55155 (I940730,I941220,I940776);
not I_55156 (I941242,I941220);
and I_55157 (I941259,I941242,I940776);
nor I_55158 (I940724,I940801,I941259);
nand I_55159 (I941290,I941242,I940852);
nor I_55160 (I940718,I941112,I941290);
nand I_55161 (I940721,I941242,I941030);
nand I_55162 (I941335,I940852,I422402);
nor I_55163 (I940733,I941095,I941335);
not I_55164 (I941396,I3570);
DFFARX1 I_55165 (I1341643,I3563,I941396,I941422,);
DFFARX1 I_55166 (I1341667,I3563,I941396,I941439,);
not I_55167 (I941447,I941439);
not I_55168 (I941464,I1341649);
nor I_55169 (I941481,I941464,I1341658);
not I_55170 (I941498,I1341643);
nor I_55171 (I941515,I941481,I1341664);
nor I_55172 (I941532,I941439,I941515);
DFFARX1 I_55173 (I941532,I3563,I941396,I941382,);
nor I_55174 (I941563,I1341664,I1341658);
nand I_55175 (I941580,I941563,I1341649);
DFFARX1 I_55176 (I941580,I3563,I941396,I941385,);
nor I_55177 (I941611,I941498,I1341664);
nand I_55178 (I941628,I941611,I1341661);
nor I_55179 (I941645,I941422,I941628);
DFFARX1 I_55180 (I941645,I3563,I941396,I941361,);
not I_55181 (I941676,I941628);
nand I_55182 (I941373,I941439,I941676);
DFFARX1 I_55183 (I941628,I3563,I941396,I941716,);
not I_55184 (I941724,I941716);
not I_55185 (I941741,I1341664);
not I_55186 (I941758,I1341655);
nor I_55187 (I941775,I941758,I1341643);
nor I_55188 (I941388,I941724,I941775);
nor I_55189 (I941806,I941758,I1341646);
and I_55190 (I941823,I941806,I1341670);
or I_55191 (I941840,I941823,I1341652);
DFFARX1 I_55192 (I941840,I3563,I941396,I941866,);
nor I_55193 (I941376,I941866,I941422);
not I_55194 (I941888,I941866);
and I_55195 (I941905,I941888,I941422);
nor I_55196 (I941370,I941447,I941905);
nand I_55197 (I941936,I941888,I941498);
nor I_55198 (I941364,I941758,I941936);
nand I_55199 (I941367,I941888,I941676);
nand I_55200 (I941981,I941498,I1341655);
nor I_55201 (I941379,I941741,I941981);
not I_55202 (I942042,I3570);
DFFARX1 I_55203 (I155723,I3563,I942042,I942068,);
DFFARX1 I_55204 (I155729,I3563,I942042,I942085,);
not I_55205 (I942093,I942085);
not I_55206 (I942110,I155747);
nor I_55207 (I942127,I942110,I155726);
not I_55208 (I942144,I155732);
nor I_55209 (I942161,I942127,I155738);
nor I_55210 (I942178,I942085,I942161);
DFFARX1 I_55211 (I942178,I3563,I942042,I942028,);
nor I_55212 (I942209,I155738,I155726);
nand I_55213 (I942226,I942209,I155747);
DFFARX1 I_55214 (I942226,I3563,I942042,I942031,);
nor I_55215 (I942257,I942144,I155738);
nand I_55216 (I942274,I942257,I155744);
nor I_55217 (I942291,I942068,I942274);
DFFARX1 I_55218 (I942291,I3563,I942042,I942007,);
not I_55219 (I942322,I942274);
nand I_55220 (I942019,I942085,I942322);
DFFARX1 I_55221 (I942274,I3563,I942042,I942362,);
not I_55222 (I942370,I942362);
not I_55223 (I942387,I155738);
not I_55224 (I942404,I155726);
nor I_55225 (I942421,I942404,I155732);
nor I_55226 (I942034,I942370,I942421);
nor I_55227 (I942452,I942404,I155735);
and I_55228 (I942469,I942452,I155723);
or I_55229 (I942486,I942469,I155741);
DFFARX1 I_55230 (I942486,I3563,I942042,I942512,);
nor I_55231 (I942022,I942512,I942068);
not I_55232 (I942534,I942512);
and I_55233 (I942551,I942534,I942068);
nor I_55234 (I942016,I942093,I942551);
nand I_55235 (I942582,I942534,I942144);
nor I_55236 (I942010,I942404,I942582);
nand I_55237 (I942013,I942534,I942322);
nand I_55238 (I942627,I942144,I155726);
nor I_55239 (I942025,I942387,I942627);
not I_55240 (I942688,I3570);
DFFARX1 I_55241 (I808121,I3563,I942688,I942714,);
DFFARX1 I_55242 (I808115,I3563,I942688,I942731,);
not I_55243 (I942739,I942731);
not I_55244 (I942756,I808130);
nor I_55245 (I942773,I942756,I808115);
not I_55246 (I942790,I808124);
nor I_55247 (I942807,I942773,I808133);
nor I_55248 (I942824,I942731,I942807);
DFFARX1 I_55249 (I942824,I3563,I942688,I942674,);
nor I_55250 (I942855,I808133,I808115);
nand I_55251 (I942872,I942855,I808130);
DFFARX1 I_55252 (I942872,I3563,I942688,I942677,);
nor I_55253 (I942903,I942790,I808133);
nand I_55254 (I942920,I942903,I808118);
nor I_55255 (I942937,I942714,I942920);
DFFARX1 I_55256 (I942937,I3563,I942688,I942653,);
not I_55257 (I942968,I942920);
nand I_55258 (I942665,I942731,I942968);
DFFARX1 I_55259 (I942920,I3563,I942688,I943008,);
not I_55260 (I943016,I943008);
not I_55261 (I943033,I808133);
not I_55262 (I943050,I808127);
nor I_55263 (I943067,I943050,I808124);
nor I_55264 (I942680,I943016,I943067);
nor I_55265 (I943098,I943050,I808136);
and I_55266 (I943115,I943098,I808139);
or I_55267 (I943132,I943115,I808118);
DFFARX1 I_55268 (I943132,I3563,I942688,I943158,);
nor I_55269 (I942668,I943158,I942714);
not I_55270 (I943180,I943158);
and I_55271 (I943197,I943180,I942714);
nor I_55272 (I942662,I942739,I943197);
nand I_55273 (I943228,I943180,I942790);
nor I_55274 (I942656,I943050,I943228);
nand I_55275 (I942659,I943180,I942968);
nand I_55276 (I943273,I942790,I808127);
nor I_55277 (I942671,I943033,I943273);
not I_55278 (I943334,I3570);
DFFARX1 I_55279 (I1071904,I3563,I943334,I943360,);
DFFARX1 I_55280 (I1071907,I3563,I943334,I943377,);
not I_55281 (I943385,I943377);
not I_55282 (I943402,I1071904);
nor I_55283 (I943419,I943402,I1071916);
not I_55284 (I943436,I1071925);
nor I_55285 (I943453,I943419,I1071913);
nor I_55286 (I943470,I943377,I943453);
DFFARX1 I_55287 (I943470,I3563,I943334,I943320,);
nor I_55288 (I943501,I1071913,I1071916);
nand I_55289 (I943518,I943501,I1071904);
DFFARX1 I_55290 (I943518,I3563,I943334,I943323,);
nor I_55291 (I943549,I943436,I1071913);
nand I_55292 (I943566,I943549,I1071919);
nor I_55293 (I943583,I943360,I943566);
DFFARX1 I_55294 (I943583,I3563,I943334,I943299,);
not I_55295 (I943614,I943566);
nand I_55296 (I943311,I943377,I943614);
DFFARX1 I_55297 (I943566,I3563,I943334,I943654,);
not I_55298 (I943662,I943654);
not I_55299 (I943679,I1071913);
not I_55300 (I943696,I1071910);
nor I_55301 (I943713,I943696,I1071925);
nor I_55302 (I943326,I943662,I943713);
nor I_55303 (I943744,I943696,I1071922);
and I_55304 (I943761,I943744,I1071910);
or I_55305 (I943778,I943761,I1071907);
DFFARX1 I_55306 (I943778,I3563,I943334,I943804,);
nor I_55307 (I943314,I943804,I943360);
not I_55308 (I943826,I943804);
and I_55309 (I943843,I943826,I943360);
nor I_55310 (I943308,I943385,I943843);
nand I_55311 (I943874,I943826,I943436);
nor I_55312 (I943302,I943696,I943874);
nand I_55313 (I943305,I943826,I943614);
nand I_55314 (I943919,I943436,I1071910);
nor I_55315 (I943317,I943679,I943919);
not I_55316 (I943980,I3570);
DFFARX1 I_55317 (I86686,I3563,I943980,I944006,);
DFFARX1 I_55318 (I86692,I3563,I943980,I944023,);
not I_55319 (I944031,I944023);
not I_55320 (I944048,I86710);
nor I_55321 (I944065,I944048,I86689);
not I_55322 (I944082,I86695);
nor I_55323 (I944099,I944065,I86701);
nor I_55324 (I944116,I944023,I944099);
DFFARX1 I_55325 (I944116,I3563,I943980,I943966,);
nor I_55326 (I944147,I86701,I86689);
nand I_55327 (I944164,I944147,I86710);
DFFARX1 I_55328 (I944164,I3563,I943980,I943969,);
nor I_55329 (I944195,I944082,I86701);
nand I_55330 (I944212,I944195,I86707);
nor I_55331 (I944229,I944006,I944212);
DFFARX1 I_55332 (I944229,I3563,I943980,I943945,);
not I_55333 (I944260,I944212);
nand I_55334 (I943957,I944023,I944260);
DFFARX1 I_55335 (I944212,I3563,I943980,I944300,);
not I_55336 (I944308,I944300);
not I_55337 (I944325,I86701);
not I_55338 (I944342,I86689);
nor I_55339 (I944359,I944342,I86695);
nor I_55340 (I943972,I944308,I944359);
nor I_55341 (I944390,I944342,I86698);
and I_55342 (I944407,I944390,I86686);
or I_55343 (I944424,I944407,I86704);
DFFARX1 I_55344 (I944424,I3563,I943980,I944450,);
nor I_55345 (I943960,I944450,I944006);
not I_55346 (I944472,I944450);
and I_55347 (I944489,I944472,I944006);
nor I_55348 (I943954,I944031,I944489);
nand I_55349 (I944520,I944472,I944082);
nor I_55350 (I943948,I944342,I944520);
nand I_55351 (I943951,I944472,I944260);
nand I_55352 (I944565,I944082,I86689);
nor I_55353 (I943963,I944325,I944565);
not I_55354 (I944626,I3570);
DFFARX1 I_55355 (I369158,I3563,I944626,I944652,);
DFFARX1 I_55356 (I369164,I3563,I944626,I944669,);
not I_55357 (I944677,I944669);
not I_55358 (I944694,I369185);
nor I_55359 (I944711,I944694,I369173);
not I_55360 (I944728,I369182);
nor I_55361 (I944745,I944711,I369167);
nor I_55362 (I944762,I944669,I944745);
DFFARX1 I_55363 (I944762,I3563,I944626,I944612,);
nor I_55364 (I944793,I369167,I369173);
nand I_55365 (I944810,I944793,I369185);
DFFARX1 I_55366 (I944810,I3563,I944626,I944615,);
nor I_55367 (I944841,I944728,I369167);
nand I_55368 (I944858,I944841,I369158);
nor I_55369 (I944875,I944652,I944858);
DFFARX1 I_55370 (I944875,I3563,I944626,I944591,);
not I_55371 (I944906,I944858);
nand I_55372 (I944603,I944669,I944906);
DFFARX1 I_55373 (I944858,I3563,I944626,I944946,);
not I_55374 (I944954,I944946);
not I_55375 (I944971,I369167);
not I_55376 (I944988,I369170);
nor I_55377 (I945005,I944988,I369182);
nor I_55378 (I944618,I944954,I945005);
nor I_55379 (I945036,I944988,I369179);
and I_55380 (I945053,I945036,I369161);
or I_55381 (I945070,I945053,I369176);
DFFARX1 I_55382 (I945070,I3563,I944626,I945096,);
nor I_55383 (I944606,I945096,I944652);
not I_55384 (I945118,I945096);
and I_55385 (I945135,I945118,I944652);
nor I_55386 (I944600,I944677,I945135);
nand I_55387 (I945166,I945118,I944728);
nor I_55388 (I944594,I944988,I945166);
nand I_55389 (I944597,I945118,I944906);
nand I_55390 (I945211,I944728,I369170);
nor I_55391 (I944609,I944971,I945211);
not I_55392 (I945272,I3570);
DFFARX1 I_55393 (I270819,I3563,I945272,I945298,);
DFFARX1 I_55394 (I270831,I3563,I945272,I945315,);
not I_55395 (I945323,I945315);
not I_55396 (I945340,I270837);
nor I_55397 (I945357,I945340,I270822);
not I_55398 (I945374,I270813);
nor I_55399 (I945391,I945357,I270834);
nor I_55400 (I945408,I945315,I945391);
DFFARX1 I_55401 (I945408,I3563,I945272,I945258,);
nor I_55402 (I945439,I270834,I270822);
nand I_55403 (I945456,I945439,I270837);
DFFARX1 I_55404 (I945456,I3563,I945272,I945261,);
nor I_55405 (I945487,I945374,I270834);
nand I_55406 (I945504,I945487,I270816);
nor I_55407 (I945521,I945298,I945504);
DFFARX1 I_55408 (I945521,I3563,I945272,I945237,);
not I_55409 (I945552,I945504);
nand I_55410 (I945249,I945315,I945552);
DFFARX1 I_55411 (I945504,I3563,I945272,I945592,);
not I_55412 (I945600,I945592);
not I_55413 (I945617,I270834);
not I_55414 (I945634,I270825);
nor I_55415 (I945651,I945634,I270813);
nor I_55416 (I945264,I945600,I945651);
nor I_55417 (I945682,I945634,I270828);
and I_55418 (I945699,I945682,I270816);
or I_55419 (I945716,I945699,I270813);
DFFARX1 I_55420 (I945716,I3563,I945272,I945742,);
nor I_55421 (I945252,I945742,I945298);
not I_55422 (I945764,I945742);
and I_55423 (I945781,I945764,I945298);
nor I_55424 (I945246,I945323,I945781);
nand I_55425 (I945812,I945764,I945374);
nor I_55426 (I945240,I945634,I945812);
nand I_55427 (I945243,I945764,I945552);
nand I_55428 (I945857,I945374,I270825);
nor I_55429 (I945255,I945617,I945857);
not I_55430 (I945918,I3570);
DFFARX1 I_55431 (I672869,I3563,I945918,I945944,);
DFFARX1 I_55432 (I672863,I3563,I945918,I945961,);
not I_55433 (I945969,I945961);
not I_55434 (I945986,I672878);
nor I_55435 (I946003,I945986,I672863);
not I_55436 (I946020,I672872);
nor I_55437 (I946037,I946003,I672881);
nor I_55438 (I946054,I945961,I946037);
DFFARX1 I_55439 (I946054,I3563,I945918,I945904,);
nor I_55440 (I946085,I672881,I672863);
nand I_55441 (I946102,I946085,I672878);
DFFARX1 I_55442 (I946102,I3563,I945918,I945907,);
nor I_55443 (I946133,I946020,I672881);
nand I_55444 (I946150,I946133,I672866);
nor I_55445 (I946167,I945944,I946150);
DFFARX1 I_55446 (I946167,I3563,I945918,I945883,);
not I_55447 (I946198,I946150);
nand I_55448 (I945895,I945961,I946198);
DFFARX1 I_55449 (I946150,I3563,I945918,I946238,);
not I_55450 (I946246,I946238);
not I_55451 (I946263,I672881);
not I_55452 (I946280,I672875);
nor I_55453 (I946297,I946280,I672872);
nor I_55454 (I945910,I946246,I946297);
nor I_55455 (I946328,I946280,I672884);
and I_55456 (I946345,I946328,I672887);
or I_55457 (I946362,I946345,I672866);
DFFARX1 I_55458 (I946362,I3563,I945918,I946388,);
nor I_55459 (I945898,I946388,I945944);
not I_55460 (I946410,I946388);
and I_55461 (I946427,I946410,I945944);
nor I_55462 (I945892,I945969,I946427);
nand I_55463 (I946458,I946410,I946020);
nor I_55464 (I945886,I946280,I946458);
nand I_55465 (I945889,I946410,I946198);
nand I_55466 (I946503,I946020,I672875);
nor I_55467 (I945901,I946263,I946503);
not I_55468 (I946564,I3570);
DFFARX1 I_55469 (I1148813,I3563,I946564,I946590,);
DFFARX1 I_55470 (I1148795,I3563,I946564,I946607,);
not I_55471 (I946615,I946607);
not I_55472 (I946632,I1148804);
nor I_55473 (I946649,I946632,I1148816);
not I_55474 (I946666,I1148798);
nor I_55475 (I946683,I946649,I1148807);
nor I_55476 (I946700,I946607,I946683);
DFFARX1 I_55477 (I946700,I3563,I946564,I946550,);
nor I_55478 (I946731,I1148807,I1148816);
nand I_55479 (I946748,I946731,I1148804);
DFFARX1 I_55480 (I946748,I3563,I946564,I946553,);
nor I_55481 (I946779,I946666,I1148807);
nand I_55482 (I946796,I946779,I1148819);
nor I_55483 (I946813,I946590,I946796);
DFFARX1 I_55484 (I946813,I3563,I946564,I946529,);
not I_55485 (I946844,I946796);
nand I_55486 (I946541,I946607,I946844);
DFFARX1 I_55487 (I946796,I3563,I946564,I946884,);
not I_55488 (I946892,I946884);
not I_55489 (I946909,I1148807);
not I_55490 (I946926,I1148795);
nor I_55491 (I946943,I946926,I1148798);
nor I_55492 (I946556,I946892,I946943);
nor I_55493 (I946974,I946926,I1148801);
and I_55494 (I946991,I946974,I1148810);
or I_55495 (I947008,I946991,I1148798);
DFFARX1 I_55496 (I947008,I3563,I946564,I947034,);
nor I_55497 (I946544,I947034,I946590);
not I_55498 (I947056,I947034);
and I_55499 (I947073,I947056,I946590);
nor I_55500 (I946538,I946615,I947073);
nand I_55501 (I947104,I947056,I946666);
nor I_55502 (I946532,I946926,I947104);
nand I_55503 (I946535,I947056,I946844);
nand I_55504 (I947149,I946666,I1148795);
nor I_55505 (I946547,I946909,I947149);
not I_55506 (I947210,I3570);
DFFARX1 I_55507 (I890639,I3563,I947210,I947236,);
DFFARX1 I_55508 (I890636,I3563,I947210,I947253,);
not I_55509 (I947261,I947253);
not I_55510 (I947278,I890636);
nor I_55511 (I947295,I947278,I890639);
not I_55512 (I947312,I890651);
nor I_55513 (I947329,I947295,I890645);
nor I_55514 (I947346,I947253,I947329);
DFFARX1 I_55515 (I947346,I3563,I947210,I947196,);
nor I_55516 (I947377,I890645,I890639);
nand I_55517 (I947394,I947377,I890636);
DFFARX1 I_55518 (I947394,I3563,I947210,I947199,);
nor I_55519 (I947425,I947312,I890645);
nand I_55520 (I947442,I947425,I890633);
nor I_55521 (I947459,I947236,I947442);
DFFARX1 I_55522 (I947459,I3563,I947210,I947175,);
not I_55523 (I947490,I947442);
nand I_55524 (I947187,I947253,I947490);
DFFARX1 I_55525 (I947442,I3563,I947210,I947530,);
not I_55526 (I947538,I947530);
not I_55527 (I947555,I890645);
not I_55528 (I947572,I890642);
nor I_55529 (I947589,I947572,I890651);
nor I_55530 (I947202,I947538,I947589);
nor I_55531 (I947620,I947572,I890648);
and I_55532 (I947637,I947620,I890654);
or I_55533 (I947654,I947637,I890633);
DFFARX1 I_55534 (I947654,I3563,I947210,I947680,);
nor I_55535 (I947190,I947680,I947236);
not I_55536 (I947702,I947680);
and I_55537 (I947719,I947702,I947236);
nor I_55538 (I947184,I947261,I947719);
nand I_55539 (I947750,I947702,I947312);
nor I_55540 (I947178,I947572,I947750);
nand I_55541 (I947181,I947702,I947490);
nand I_55542 (I947795,I947312,I890642);
nor I_55543 (I947193,I947555,I947795);
not I_55544 (I947856,I3570);
DFFARX1 I_55545 (I496936,I3563,I947856,I947882,);
DFFARX1 I_55546 (I496933,I3563,I947856,I947899,);
not I_55547 (I947907,I947899);
not I_55548 (I947924,I496948);
nor I_55549 (I947941,I947924,I496951);
not I_55550 (I947958,I496939);
nor I_55551 (I947975,I947941,I496945);
nor I_55552 (I947992,I947899,I947975);
DFFARX1 I_55553 (I947992,I3563,I947856,I947842,);
nor I_55554 (I948023,I496945,I496951);
nand I_55555 (I948040,I948023,I496948);
DFFARX1 I_55556 (I948040,I3563,I947856,I947845,);
nor I_55557 (I948071,I947958,I496945);
nand I_55558 (I948088,I948071,I496957);
nor I_55559 (I948105,I947882,I948088);
DFFARX1 I_55560 (I948105,I3563,I947856,I947821,);
not I_55561 (I948136,I948088);
nand I_55562 (I947833,I947899,I948136);
DFFARX1 I_55563 (I948088,I3563,I947856,I948176,);
not I_55564 (I948184,I948176);
not I_55565 (I948201,I496945);
not I_55566 (I948218,I496930);
nor I_55567 (I948235,I948218,I496939);
nor I_55568 (I947848,I948184,I948235);
nor I_55569 (I948266,I948218,I496942);
and I_55570 (I948283,I948266,I496930);
or I_55571 (I948300,I948283,I496954);
DFFARX1 I_55572 (I948300,I3563,I947856,I948326,);
nor I_55573 (I947836,I948326,I947882);
not I_55574 (I948348,I948326);
and I_55575 (I948365,I948348,I947882);
nor I_55576 (I947830,I947907,I948365);
nand I_55577 (I948396,I948348,I947958);
nor I_55578 (I947824,I948218,I948396);
nand I_55579 (I947827,I948348,I948136);
nand I_55580 (I948441,I947958,I496930);
nor I_55581 (I947839,I948201,I948441);
not I_55582 (I948502,I3570);
DFFARX1 I_55583 (I658419,I3563,I948502,I948528,);
DFFARX1 I_55584 (I658413,I3563,I948502,I948545,);
not I_55585 (I948553,I948545);
not I_55586 (I948570,I658428);
nor I_55587 (I948587,I948570,I658413);
not I_55588 (I948604,I658422);
nor I_55589 (I948621,I948587,I658431);
nor I_55590 (I948638,I948545,I948621);
DFFARX1 I_55591 (I948638,I3563,I948502,I948488,);
nor I_55592 (I948669,I658431,I658413);
nand I_55593 (I948686,I948669,I658428);
DFFARX1 I_55594 (I948686,I3563,I948502,I948491,);
nor I_55595 (I948717,I948604,I658431);
nand I_55596 (I948734,I948717,I658416);
nor I_55597 (I948751,I948528,I948734);
DFFARX1 I_55598 (I948751,I3563,I948502,I948467,);
not I_55599 (I948782,I948734);
nand I_55600 (I948479,I948545,I948782);
DFFARX1 I_55601 (I948734,I3563,I948502,I948822,);
not I_55602 (I948830,I948822);
not I_55603 (I948847,I658431);
not I_55604 (I948864,I658425);
nor I_55605 (I948881,I948864,I658422);
nor I_55606 (I948494,I948830,I948881);
nor I_55607 (I948912,I948864,I658434);
and I_55608 (I948929,I948912,I658437);
or I_55609 (I948946,I948929,I658416);
DFFARX1 I_55610 (I948946,I3563,I948502,I948972,);
nor I_55611 (I948482,I948972,I948528);
not I_55612 (I948994,I948972);
and I_55613 (I949011,I948994,I948528);
nor I_55614 (I948476,I948553,I949011);
nand I_55615 (I949042,I948994,I948604);
nor I_55616 (I948470,I948864,I949042);
nand I_55617 (I948473,I948994,I948782);
nand I_55618 (I949087,I948604,I658425);
nor I_55619 (I948485,I948847,I949087);
not I_55620 (I949148,I3570);
DFFARX1 I_55621 (I1369013,I3563,I949148,I949174,);
DFFARX1 I_55622 (I1369037,I3563,I949148,I949191,);
not I_55623 (I949199,I949191);
not I_55624 (I949216,I1369019);
nor I_55625 (I949233,I949216,I1369028);
not I_55626 (I949250,I1369013);
nor I_55627 (I949267,I949233,I1369034);
nor I_55628 (I949284,I949191,I949267);
DFFARX1 I_55629 (I949284,I3563,I949148,I949134,);
nor I_55630 (I949315,I1369034,I1369028);
nand I_55631 (I949332,I949315,I1369019);
DFFARX1 I_55632 (I949332,I3563,I949148,I949137,);
nor I_55633 (I949363,I949250,I1369034);
nand I_55634 (I949380,I949363,I1369031);
nor I_55635 (I949397,I949174,I949380);
DFFARX1 I_55636 (I949397,I3563,I949148,I949113,);
not I_55637 (I949428,I949380);
nand I_55638 (I949125,I949191,I949428);
DFFARX1 I_55639 (I949380,I3563,I949148,I949468,);
not I_55640 (I949476,I949468);
not I_55641 (I949493,I1369034);
not I_55642 (I949510,I1369025);
nor I_55643 (I949527,I949510,I1369013);
nor I_55644 (I949140,I949476,I949527);
nor I_55645 (I949558,I949510,I1369016);
and I_55646 (I949575,I949558,I1369040);
or I_55647 (I949592,I949575,I1369022);
DFFARX1 I_55648 (I949592,I3563,I949148,I949618,);
nor I_55649 (I949128,I949618,I949174);
not I_55650 (I949640,I949618);
and I_55651 (I949657,I949640,I949174);
nor I_55652 (I949122,I949199,I949657);
nand I_55653 (I949688,I949640,I949250);
nor I_55654 (I949116,I949510,I949688);
nand I_55655 (I949119,I949640,I949428);
nand I_55656 (I949733,I949250,I1369025);
nor I_55657 (I949131,I949493,I949733);
not I_55658 (I949794,I3570);
DFFARX1 I_55659 (I282719,I3563,I949794,I949820,);
DFFARX1 I_55660 (I282731,I3563,I949794,I949837,);
not I_55661 (I949845,I949837);
not I_55662 (I949862,I282737);
nor I_55663 (I949879,I949862,I282722);
not I_55664 (I949896,I282713);
nor I_55665 (I949913,I949879,I282734);
nor I_55666 (I949930,I949837,I949913);
DFFARX1 I_55667 (I949930,I3563,I949794,I949780,);
nor I_55668 (I949961,I282734,I282722);
nand I_55669 (I949978,I949961,I282737);
DFFARX1 I_55670 (I949978,I3563,I949794,I949783,);
nor I_55671 (I950009,I949896,I282734);
nand I_55672 (I950026,I950009,I282716);
nor I_55673 (I950043,I949820,I950026);
DFFARX1 I_55674 (I950043,I3563,I949794,I949759,);
not I_55675 (I950074,I950026);
nand I_55676 (I949771,I949837,I950074);
DFFARX1 I_55677 (I950026,I3563,I949794,I950114,);
not I_55678 (I950122,I950114);
not I_55679 (I950139,I282734);
not I_55680 (I950156,I282725);
nor I_55681 (I950173,I950156,I282713);
nor I_55682 (I949786,I950122,I950173);
nor I_55683 (I950204,I950156,I282728);
and I_55684 (I950221,I950204,I282716);
or I_55685 (I950238,I950221,I282713);
DFFARX1 I_55686 (I950238,I3563,I949794,I950264,);
nor I_55687 (I949774,I950264,I949820);
not I_55688 (I950286,I950264);
and I_55689 (I950303,I950286,I949820);
nor I_55690 (I949768,I949845,I950303);
nand I_55691 (I950334,I950286,I949896);
nor I_55692 (I949762,I950156,I950334);
nand I_55693 (I949765,I950286,I950074);
nand I_55694 (I950379,I949896,I282725);
nor I_55695 (I949777,I950139,I950379);
not I_55696 (I950440,I3570);
DFFARX1 I_55697 (I263084,I3563,I950440,I950466,);
DFFARX1 I_55698 (I263096,I3563,I950440,I950483,);
not I_55699 (I950491,I950483);
not I_55700 (I950508,I263102);
nor I_55701 (I950525,I950508,I263087);
not I_55702 (I950542,I263078);
nor I_55703 (I950559,I950525,I263099);
nor I_55704 (I950576,I950483,I950559);
DFFARX1 I_55705 (I950576,I3563,I950440,I950426,);
nor I_55706 (I950607,I263099,I263087);
nand I_55707 (I950624,I950607,I263102);
DFFARX1 I_55708 (I950624,I3563,I950440,I950429,);
nor I_55709 (I950655,I950542,I263099);
nand I_55710 (I950672,I950655,I263081);
nor I_55711 (I950689,I950466,I950672);
DFFARX1 I_55712 (I950689,I3563,I950440,I950405,);
not I_55713 (I950720,I950672);
nand I_55714 (I950417,I950483,I950720);
DFFARX1 I_55715 (I950672,I3563,I950440,I950760,);
not I_55716 (I950768,I950760);
not I_55717 (I950785,I263099);
not I_55718 (I950802,I263090);
nor I_55719 (I950819,I950802,I263078);
nor I_55720 (I950432,I950768,I950819);
nor I_55721 (I950850,I950802,I263093);
and I_55722 (I950867,I950850,I263081);
or I_55723 (I950884,I950867,I263078);
DFFARX1 I_55724 (I950884,I3563,I950440,I950910,);
nor I_55725 (I950420,I950910,I950466);
not I_55726 (I950932,I950910);
and I_55727 (I950949,I950932,I950466);
nor I_55728 (I950414,I950491,I950949);
nand I_55729 (I950980,I950932,I950542);
nor I_55730 (I950408,I950802,I950980);
nand I_55731 (I950411,I950932,I950720);
nand I_55732 (I951025,I950542,I263090);
nor I_55733 (I950423,I950785,I951025);
not I_55734 (I951086,I3570);
DFFARX1 I_55735 (I1255131,I3563,I951086,I951112,);
DFFARX1 I_55736 (I1255137,I3563,I951086,I951129,);
not I_55737 (I951137,I951129);
not I_55738 (I951154,I1255134);
nor I_55739 (I951171,I951154,I1255113);
not I_55740 (I951188,I1255116);
nor I_55741 (I951205,I951171,I1255122);
nor I_55742 (I951222,I951129,I951205);
DFFARX1 I_55743 (I951222,I3563,I951086,I951072,);
nor I_55744 (I951253,I1255122,I1255113);
nand I_55745 (I951270,I951253,I1255134);
DFFARX1 I_55746 (I951270,I3563,I951086,I951075,);
nor I_55747 (I951301,I951188,I1255122);
nand I_55748 (I951318,I951301,I1255116);
nor I_55749 (I951335,I951112,I951318);
DFFARX1 I_55750 (I951335,I3563,I951086,I951051,);
not I_55751 (I951366,I951318);
nand I_55752 (I951063,I951129,I951366);
DFFARX1 I_55753 (I951318,I3563,I951086,I951406,);
not I_55754 (I951414,I951406);
not I_55755 (I951431,I1255122);
not I_55756 (I951448,I1255125);
nor I_55757 (I951465,I951448,I1255116);
nor I_55758 (I951078,I951414,I951465);
nor I_55759 (I951496,I951448,I1255113);
and I_55760 (I951513,I951496,I1255119);
or I_55761 (I951530,I951513,I1255128);
DFFARX1 I_55762 (I951530,I3563,I951086,I951556,);
nor I_55763 (I951066,I951556,I951112);
not I_55764 (I951578,I951556);
and I_55765 (I951595,I951578,I951112);
nor I_55766 (I951060,I951137,I951595);
nand I_55767 (I951626,I951578,I951188);
nor I_55768 (I951054,I951448,I951626);
nand I_55769 (I951057,I951578,I951366);
nand I_55770 (I951671,I951188,I1255125);
nor I_55771 (I951069,I951431,I951671);
not I_55772 (I951732,I3570);
DFFARX1 I_55773 (I55593,I3563,I951732,I951758,);
DFFARX1 I_55774 (I55599,I3563,I951732,I951775,);
not I_55775 (I951783,I951775);
not I_55776 (I951800,I55593);
nor I_55777 (I951817,I951800,I55605);
not I_55778 (I951834,I55617);
nor I_55779 (I951851,I951817,I55611);
nor I_55780 (I951868,I951775,I951851);
DFFARX1 I_55781 (I951868,I3563,I951732,I951718,);
nor I_55782 (I951899,I55611,I55605);
nand I_55783 (I951916,I951899,I55593);
DFFARX1 I_55784 (I951916,I3563,I951732,I951721,);
nor I_55785 (I951947,I951834,I55611);
nand I_55786 (I951964,I951947,I55596);
nor I_55787 (I951981,I951758,I951964);
DFFARX1 I_55788 (I951981,I3563,I951732,I951697,);
not I_55789 (I952012,I951964);
nand I_55790 (I951709,I951775,I952012);
DFFARX1 I_55791 (I951964,I3563,I951732,I952052,);
not I_55792 (I952060,I952052);
not I_55793 (I952077,I55611);
not I_55794 (I952094,I55596);
nor I_55795 (I952111,I952094,I55617);
nor I_55796 (I951724,I952060,I952111);
nor I_55797 (I952142,I952094,I55614);
and I_55798 (I952159,I952142,I55608);
or I_55799 (I952176,I952159,I55602);
DFFARX1 I_55800 (I952176,I3563,I951732,I952202,);
nor I_55801 (I951712,I952202,I951758);
not I_55802 (I952224,I952202);
and I_55803 (I952241,I952224,I951758);
nor I_55804 (I951706,I951783,I952241);
nand I_55805 (I952272,I952224,I951834);
nor I_55806 (I951700,I952094,I952272);
nand I_55807 (I951703,I952224,I952012);
nand I_55808 (I952317,I951834,I55596);
nor I_55809 (I951715,I952077,I952317);
not I_55810 (I952378,I3570);
DFFARX1 I_55811 (I888531,I3563,I952378,I952404,);
DFFARX1 I_55812 (I888528,I3563,I952378,I952421,);
not I_55813 (I952429,I952421);
not I_55814 (I952446,I888528);
nor I_55815 (I952463,I952446,I888531);
not I_55816 (I952480,I888543);
nor I_55817 (I952497,I952463,I888537);
nor I_55818 (I952514,I952421,I952497);
DFFARX1 I_55819 (I952514,I3563,I952378,I952364,);
nor I_55820 (I952545,I888537,I888531);
nand I_55821 (I952562,I952545,I888528);
DFFARX1 I_55822 (I952562,I3563,I952378,I952367,);
nor I_55823 (I952593,I952480,I888537);
nand I_55824 (I952610,I952593,I888525);
nor I_55825 (I952627,I952404,I952610);
DFFARX1 I_55826 (I952627,I3563,I952378,I952343,);
not I_55827 (I952658,I952610);
nand I_55828 (I952355,I952421,I952658);
DFFARX1 I_55829 (I952610,I3563,I952378,I952698,);
not I_55830 (I952706,I952698);
not I_55831 (I952723,I888537);
not I_55832 (I952740,I888534);
nor I_55833 (I952757,I952740,I888543);
nor I_55834 (I952370,I952706,I952757);
nor I_55835 (I952788,I952740,I888540);
and I_55836 (I952805,I952788,I888546);
or I_55837 (I952822,I952805,I888525);
DFFARX1 I_55838 (I952822,I3563,I952378,I952848,);
nor I_55839 (I952358,I952848,I952404);
not I_55840 (I952870,I952848);
and I_55841 (I952887,I952870,I952404);
nor I_55842 (I952352,I952429,I952887);
nand I_55843 (I952918,I952870,I952480);
nor I_55844 (I952346,I952740,I952918);
nand I_55845 (I952349,I952870,I952658);
nand I_55846 (I952963,I952480,I888534);
nor I_55847 (I952361,I952723,I952963);
not I_55848 (I953024,I3570);
DFFARX1 I_55849 (I851114,I3563,I953024,I953050,);
DFFARX1 I_55850 (I851111,I3563,I953024,I953067,);
not I_55851 (I953075,I953067);
not I_55852 (I953092,I851111);
nor I_55853 (I953109,I953092,I851114);
not I_55854 (I953126,I851126);
nor I_55855 (I953143,I953109,I851120);
nor I_55856 (I953160,I953067,I953143);
DFFARX1 I_55857 (I953160,I3563,I953024,I953010,);
nor I_55858 (I953191,I851120,I851114);
nand I_55859 (I953208,I953191,I851111);
DFFARX1 I_55860 (I953208,I3563,I953024,I953013,);
nor I_55861 (I953239,I953126,I851120);
nand I_55862 (I953256,I953239,I851108);
nor I_55863 (I953273,I953050,I953256);
DFFARX1 I_55864 (I953273,I3563,I953024,I952989,);
not I_55865 (I953304,I953256);
nand I_55866 (I953001,I953067,I953304);
DFFARX1 I_55867 (I953256,I3563,I953024,I953344,);
not I_55868 (I953352,I953344);
not I_55869 (I953369,I851120);
not I_55870 (I953386,I851117);
nor I_55871 (I953403,I953386,I851126);
nor I_55872 (I953016,I953352,I953403);
nor I_55873 (I953434,I953386,I851123);
and I_55874 (I953451,I953434,I851129);
or I_55875 (I953468,I953451,I851108);
DFFARX1 I_55876 (I953468,I3563,I953024,I953494,);
nor I_55877 (I953004,I953494,I953050);
not I_55878 (I953516,I953494);
and I_55879 (I953533,I953516,I953050);
nor I_55880 (I952998,I953075,I953533);
nand I_55881 (I953564,I953516,I953126);
nor I_55882 (I952992,I953386,I953564);
nand I_55883 (I952995,I953516,I953304);
nand I_55884 (I953609,I953126,I851117);
nor I_55885 (I953007,I953369,I953609);
not I_55886 (I953670,I3570);
DFFARX1 I_55887 (I494760,I3563,I953670,I953696,);
DFFARX1 I_55888 (I494757,I3563,I953670,I953713,);
not I_55889 (I953721,I953713);
not I_55890 (I953738,I494772);
nor I_55891 (I953755,I953738,I494775);
not I_55892 (I953772,I494763);
nor I_55893 (I953789,I953755,I494769);
nor I_55894 (I953806,I953713,I953789);
DFFARX1 I_55895 (I953806,I3563,I953670,I953656,);
nor I_55896 (I953837,I494769,I494775);
nand I_55897 (I953854,I953837,I494772);
DFFARX1 I_55898 (I953854,I3563,I953670,I953659,);
nor I_55899 (I953885,I953772,I494769);
nand I_55900 (I953902,I953885,I494781);
nor I_55901 (I953919,I953696,I953902);
DFFARX1 I_55902 (I953919,I3563,I953670,I953635,);
not I_55903 (I953950,I953902);
nand I_55904 (I953647,I953713,I953950);
DFFARX1 I_55905 (I953902,I3563,I953670,I953990,);
not I_55906 (I953998,I953990);
not I_55907 (I954015,I494769);
not I_55908 (I954032,I494754);
nor I_55909 (I954049,I954032,I494763);
nor I_55910 (I953662,I953998,I954049);
nor I_55911 (I954080,I954032,I494766);
and I_55912 (I954097,I954080,I494754);
or I_55913 (I954114,I954097,I494778);
DFFARX1 I_55914 (I954114,I3563,I953670,I954140,);
nor I_55915 (I953650,I954140,I953696);
not I_55916 (I954162,I954140);
and I_55917 (I954179,I954162,I953696);
nor I_55918 (I953644,I953721,I954179);
nand I_55919 (I954210,I954162,I953772);
nor I_55920 (I953638,I954032,I954210);
nand I_55921 (I953641,I954162,I953950);
nand I_55922 (I954255,I953772,I494754);
nor I_55923 (I953653,I954015,I954255);
not I_55924 (I954316,I3570);
DFFARX1 I_55925 (I795983,I3563,I954316,I954342,);
DFFARX1 I_55926 (I795977,I3563,I954316,I954359,);
not I_55927 (I954367,I954359);
not I_55928 (I954384,I795992);
nor I_55929 (I954401,I954384,I795977);
not I_55930 (I954418,I795986);
nor I_55931 (I954435,I954401,I795995);
nor I_55932 (I954452,I954359,I954435);
DFFARX1 I_55933 (I954452,I3563,I954316,I954302,);
nor I_55934 (I954483,I795995,I795977);
nand I_55935 (I954500,I954483,I795992);
DFFARX1 I_55936 (I954500,I3563,I954316,I954305,);
nor I_55937 (I954531,I954418,I795995);
nand I_55938 (I954548,I954531,I795980);
nor I_55939 (I954565,I954342,I954548);
DFFARX1 I_55940 (I954565,I3563,I954316,I954281,);
not I_55941 (I954596,I954548);
nand I_55942 (I954293,I954359,I954596);
DFFARX1 I_55943 (I954548,I3563,I954316,I954636,);
not I_55944 (I954644,I954636);
not I_55945 (I954661,I795995);
not I_55946 (I954678,I795989);
nor I_55947 (I954695,I954678,I795986);
nor I_55948 (I954308,I954644,I954695);
nor I_55949 (I954726,I954678,I795998);
and I_55950 (I954743,I954726,I796001);
or I_55951 (I954760,I954743,I795980);
DFFARX1 I_55952 (I954760,I3563,I954316,I954786,);
nor I_55953 (I954296,I954786,I954342);
not I_55954 (I954808,I954786);
and I_55955 (I954825,I954808,I954342);
nor I_55956 (I954290,I954367,I954825);
nand I_55957 (I954856,I954808,I954418);
nor I_55958 (I954284,I954678,I954856);
nand I_55959 (I954287,I954808,I954596);
nand I_55960 (I954901,I954418,I795989);
nor I_55961 (I954299,I954661,I954901);
not I_55962 (I954962,I3570);
DFFARX1 I_55963 (I53485,I3563,I954962,I954988,);
DFFARX1 I_55964 (I53491,I3563,I954962,I955005,);
not I_55965 (I955013,I955005);
not I_55966 (I955030,I53485);
nor I_55967 (I955047,I955030,I53497);
not I_55968 (I955064,I53509);
nor I_55969 (I955081,I955047,I53503);
nor I_55970 (I955098,I955005,I955081);
DFFARX1 I_55971 (I955098,I3563,I954962,I954948,);
nor I_55972 (I955129,I53503,I53497);
nand I_55973 (I955146,I955129,I53485);
DFFARX1 I_55974 (I955146,I3563,I954962,I954951,);
nor I_55975 (I955177,I955064,I53503);
nand I_55976 (I955194,I955177,I53488);
nor I_55977 (I955211,I954988,I955194);
DFFARX1 I_55978 (I955211,I3563,I954962,I954927,);
not I_55979 (I955242,I955194);
nand I_55980 (I954939,I955005,I955242);
DFFARX1 I_55981 (I955194,I3563,I954962,I955282,);
not I_55982 (I955290,I955282);
not I_55983 (I955307,I53503);
not I_55984 (I955324,I53488);
nor I_55985 (I955341,I955324,I53509);
nor I_55986 (I954954,I955290,I955341);
nor I_55987 (I955372,I955324,I53506);
and I_55988 (I955389,I955372,I53500);
or I_55989 (I955406,I955389,I53494);
DFFARX1 I_55990 (I955406,I3563,I954962,I955432,);
nor I_55991 (I954942,I955432,I954988);
not I_55992 (I955454,I955432);
and I_55993 (I955471,I955454,I954988);
nor I_55994 (I954936,I955013,I955471);
nand I_55995 (I955502,I955454,I955064);
nor I_55996 (I954930,I955324,I955502);
nand I_55997 (I954933,I955454,I955242);
nand I_55998 (I955547,I955064,I53488);
nor I_55999 (I954945,I955307,I955547);
not I_56000 (I955608,I3570);
DFFARX1 I_56001 (I1341048,I3563,I955608,I955634,);
DFFARX1 I_56002 (I1341072,I3563,I955608,I955651,);
not I_56003 (I955659,I955651);
not I_56004 (I955676,I1341054);
nor I_56005 (I955693,I955676,I1341063);
not I_56006 (I955710,I1341048);
nor I_56007 (I955727,I955693,I1341069);
nor I_56008 (I955744,I955651,I955727);
DFFARX1 I_56009 (I955744,I3563,I955608,I955594,);
nor I_56010 (I955775,I1341069,I1341063);
nand I_56011 (I955792,I955775,I1341054);
DFFARX1 I_56012 (I955792,I3563,I955608,I955597,);
nor I_56013 (I955823,I955710,I1341069);
nand I_56014 (I955840,I955823,I1341066);
nor I_56015 (I955857,I955634,I955840);
DFFARX1 I_56016 (I955857,I3563,I955608,I955573,);
not I_56017 (I955888,I955840);
nand I_56018 (I955585,I955651,I955888);
DFFARX1 I_56019 (I955840,I3563,I955608,I955928,);
not I_56020 (I955936,I955928);
not I_56021 (I955953,I1341069);
not I_56022 (I955970,I1341060);
nor I_56023 (I955987,I955970,I1341048);
nor I_56024 (I955600,I955936,I955987);
nor I_56025 (I956018,I955970,I1341051);
and I_56026 (I956035,I956018,I1341075);
or I_56027 (I956052,I956035,I1341057);
DFFARX1 I_56028 (I956052,I3563,I955608,I956078,);
nor I_56029 (I955588,I956078,I955634);
not I_56030 (I956100,I956078);
and I_56031 (I956117,I956100,I955634);
nor I_56032 (I955582,I955659,I956117);
nand I_56033 (I956148,I956100,I955710);
nor I_56034 (I955576,I955970,I956148);
nand I_56035 (I955579,I956100,I955888);
nand I_56036 (I956193,I955710,I1341060);
nor I_56037 (I955591,I955953,I956193);
not I_56038 (I956254,I3570);
DFFARX1 I_56039 (I102496,I3563,I956254,I956280,);
DFFARX1 I_56040 (I102502,I3563,I956254,I956297,);
not I_56041 (I956305,I956297);
not I_56042 (I956322,I102520);
nor I_56043 (I956339,I956322,I102499);
not I_56044 (I956356,I102505);
nor I_56045 (I956373,I956339,I102511);
nor I_56046 (I956390,I956297,I956373);
DFFARX1 I_56047 (I956390,I3563,I956254,I956240,);
nor I_56048 (I956421,I102511,I102499);
nand I_56049 (I956438,I956421,I102520);
DFFARX1 I_56050 (I956438,I3563,I956254,I956243,);
nor I_56051 (I956469,I956356,I102511);
nand I_56052 (I956486,I956469,I102517);
nor I_56053 (I956503,I956280,I956486);
DFFARX1 I_56054 (I956503,I3563,I956254,I956219,);
not I_56055 (I956534,I956486);
nand I_56056 (I956231,I956297,I956534);
DFFARX1 I_56057 (I956486,I3563,I956254,I956574,);
not I_56058 (I956582,I956574);
not I_56059 (I956599,I102511);
not I_56060 (I956616,I102499);
nor I_56061 (I956633,I956616,I102505);
nor I_56062 (I956246,I956582,I956633);
nor I_56063 (I956664,I956616,I102508);
and I_56064 (I956681,I956664,I102496);
or I_56065 (I956698,I956681,I102514);
DFFARX1 I_56066 (I956698,I3563,I956254,I956724,);
nor I_56067 (I956234,I956724,I956280);
not I_56068 (I956746,I956724);
and I_56069 (I956763,I956746,I956280);
nor I_56070 (I956228,I956305,I956763);
nand I_56071 (I956794,I956746,I956356);
nor I_56072 (I956222,I956616,I956794);
nand I_56073 (I956225,I956746,I956534);
nand I_56074 (I956839,I956356,I102499);
nor I_56075 (I956237,I956599,I956839);
not I_56076 (I956900,I3570);
DFFARX1 I_56077 (I824764,I3563,I956900,I956926,);
DFFARX1 I_56078 (I824761,I3563,I956900,I956943,);
not I_56079 (I956951,I956943);
not I_56080 (I956968,I824761);
nor I_56081 (I956985,I956968,I824764);
not I_56082 (I957002,I824776);
nor I_56083 (I957019,I956985,I824770);
nor I_56084 (I957036,I956943,I957019);
DFFARX1 I_56085 (I957036,I3563,I956900,I956886,);
nor I_56086 (I957067,I824770,I824764);
nand I_56087 (I957084,I957067,I824761);
DFFARX1 I_56088 (I957084,I3563,I956900,I956889,);
nor I_56089 (I957115,I957002,I824770);
nand I_56090 (I957132,I957115,I824758);
nor I_56091 (I957149,I956926,I957132);
DFFARX1 I_56092 (I957149,I3563,I956900,I956865,);
not I_56093 (I957180,I957132);
nand I_56094 (I956877,I956943,I957180);
DFFARX1 I_56095 (I957132,I3563,I956900,I957220,);
not I_56096 (I957228,I957220);
not I_56097 (I957245,I824770);
not I_56098 (I957262,I824767);
nor I_56099 (I957279,I957262,I824776);
nor I_56100 (I956892,I957228,I957279);
nor I_56101 (I957310,I957262,I824773);
and I_56102 (I957327,I957310,I824779);
or I_56103 (I957344,I957327,I824758);
DFFARX1 I_56104 (I957344,I3563,I956900,I957370,);
nor I_56105 (I956880,I957370,I956926);
not I_56106 (I957392,I957370);
and I_56107 (I957409,I957392,I956926);
nor I_56108 (I956874,I956951,I957409);
nand I_56109 (I957440,I957392,I957002);
nor I_56110 (I956868,I957262,I957440);
nand I_56111 (I956871,I957392,I957180);
nand I_56112 (I957485,I957002,I824767);
nor I_56113 (I956883,I957245,I957485);
not I_56114 (I957546,I3570);
DFFARX1 I_56115 (I707549,I3563,I957546,I957572,);
DFFARX1 I_56116 (I707543,I3563,I957546,I957589,);
not I_56117 (I957597,I957589);
not I_56118 (I957614,I707558);
nor I_56119 (I957631,I957614,I707543);
not I_56120 (I957648,I707552);
nor I_56121 (I957665,I957631,I707561);
nor I_56122 (I957682,I957589,I957665);
DFFARX1 I_56123 (I957682,I3563,I957546,I957532,);
nor I_56124 (I957713,I707561,I707543);
nand I_56125 (I957730,I957713,I707558);
DFFARX1 I_56126 (I957730,I3563,I957546,I957535,);
nor I_56127 (I957761,I957648,I707561);
nand I_56128 (I957778,I957761,I707546);
nor I_56129 (I957795,I957572,I957778);
DFFARX1 I_56130 (I957795,I3563,I957546,I957511,);
not I_56131 (I957826,I957778);
nand I_56132 (I957523,I957589,I957826);
DFFARX1 I_56133 (I957778,I3563,I957546,I957866,);
not I_56134 (I957874,I957866);
not I_56135 (I957891,I707561);
not I_56136 (I957908,I707555);
nor I_56137 (I957925,I957908,I707552);
nor I_56138 (I957538,I957874,I957925);
nor I_56139 (I957956,I957908,I707564);
and I_56140 (I957973,I957956,I707567);
or I_56141 (I957990,I957973,I707546);
DFFARX1 I_56142 (I957990,I3563,I957546,I958016,);
nor I_56143 (I957526,I958016,I957572);
not I_56144 (I958038,I958016);
and I_56145 (I958055,I958038,I957572);
nor I_56146 (I957520,I957597,I958055);
nand I_56147 (I958086,I958038,I957648);
nor I_56148 (I957514,I957908,I958086);
nand I_56149 (I957517,I958038,I957826);
nand I_56150 (I958131,I957648,I707555);
nor I_56151 (I957529,I957891,I958131);
not I_56152 (I958192,I3570);
DFFARX1 I_56153 (I1112977,I3563,I958192,I958218,);
DFFARX1 I_56154 (I1112959,I3563,I958192,I958235,);
not I_56155 (I958243,I958235);
not I_56156 (I958260,I1112968);
nor I_56157 (I958277,I958260,I1112980);
not I_56158 (I958294,I1112962);
nor I_56159 (I958311,I958277,I1112971);
nor I_56160 (I958328,I958235,I958311);
DFFARX1 I_56161 (I958328,I3563,I958192,I958178,);
nor I_56162 (I958359,I1112971,I1112980);
nand I_56163 (I958376,I958359,I1112968);
DFFARX1 I_56164 (I958376,I3563,I958192,I958181,);
nor I_56165 (I958407,I958294,I1112971);
nand I_56166 (I958424,I958407,I1112983);
nor I_56167 (I958441,I958218,I958424);
DFFARX1 I_56168 (I958441,I3563,I958192,I958157,);
not I_56169 (I958472,I958424);
nand I_56170 (I958169,I958235,I958472);
DFFARX1 I_56171 (I958424,I3563,I958192,I958512,);
not I_56172 (I958520,I958512);
not I_56173 (I958537,I1112971);
not I_56174 (I958554,I1112959);
nor I_56175 (I958571,I958554,I1112962);
nor I_56176 (I958184,I958520,I958571);
nor I_56177 (I958602,I958554,I1112965);
and I_56178 (I958619,I958602,I1112974);
or I_56179 (I958636,I958619,I1112962);
DFFARX1 I_56180 (I958636,I3563,I958192,I958662,);
nor I_56181 (I958172,I958662,I958218);
not I_56182 (I958684,I958662);
and I_56183 (I958701,I958684,I958218);
nor I_56184 (I958166,I958243,I958701);
nand I_56185 (I958732,I958684,I958294);
nor I_56186 (I958160,I958554,I958732);
nand I_56187 (I958163,I958684,I958472);
nand I_56188 (I958777,I958294,I1112959);
nor I_56189 (I958175,I958537,I958777);
not I_56190 (I958838,I3570);
DFFARX1 I_56191 (I657260,I3563,I958838,I958864,);
DFFARX1 I_56192 (I657272,I3563,I958838,I958881,);
not I_56193 (I958889,I958881);
not I_56194 (I958906,I657281);
nor I_56195 (I958923,I958906,I657257);
not I_56196 (I958940,I657275);
nor I_56197 (I958957,I958923,I657269);
nor I_56198 (I958974,I958881,I958957);
DFFARX1 I_56199 (I958974,I3563,I958838,I958824,);
nor I_56200 (I959005,I657269,I657257);
nand I_56201 (I959022,I959005,I657281);
DFFARX1 I_56202 (I959022,I3563,I958838,I958827,);
nor I_56203 (I959053,I958940,I657269);
nand I_56204 (I959070,I959053,I657263);
nor I_56205 (I959087,I958864,I959070);
DFFARX1 I_56206 (I959087,I3563,I958838,I958803,);
not I_56207 (I959118,I959070);
nand I_56208 (I958815,I958881,I959118);
DFFARX1 I_56209 (I959070,I3563,I958838,I959158,);
not I_56210 (I959166,I959158);
not I_56211 (I959183,I657269);
not I_56212 (I959200,I657278);
nor I_56213 (I959217,I959200,I657275);
nor I_56214 (I958830,I959166,I959217);
nor I_56215 (I959248,I959200,I657260);
and I_56216 (I959265,I959248,I657257);
or I_56217 (I959282,I959265,I657266);
DFFARX1 I_56218 (I959282,I3563,I958838,I959308,);
nor I_56219 (I958818,I959308,I958864);
not I_56220 (I959330,I959308);
and I_56221 (I959347,I959330,I958864);
nor I_56222 (I958812,I958889,I959347);
nand I_56223 (I959378,I959330,I958940);
nor I_56224 (I958806,I959200,I959378);
nand I_56225 (I958809,I959330,I959118);
nand I_56226 (I959423,I958940,I657278);
nor I_56227 (I958821,I959183,I959423);
not I_56228 (I959484,I3570);
DFFARX1 I_56229 (I66133,I3563,I959484,I959510,);
DFFARX1 I_56230 (I66139,I3563,I959484,I959527,);
not I_56231 (I959535,I959527);
not I_56232 (I959552,I66157);
nor I_56233 (I959569,I959552,I66136);
not I_56234 (I959586,I66142);
nor I_56235 (I959603,I959569,I66148);
nor I_56236 (I959620,I959527,I959603);
DFFARX1 I_56237 (I959620,I3563,I959484,I959470,);
nor I_56238 (I959651,I66148,I66136);
nand I_56239 (I959668,I959651,I66157);
DFFARX1 I_56240 (I959668,I3563,I959484,I959473,);
nor I_56241 (I959699,I959586,I66148);
nand I_56242 (I959716,I959699,I66154);
nor I_56243 (I959733,I959510,I959716);
DFFARX1 I_56244 (I959733,I3563,I959484,I959449,);
not I_56245 (I959764,I959716);
nand I_56246 (I959461,I959527,I959764);
DFFARX1 I_56247 (I959716,I3563,I959484,I959804,);
not I_56248 (I959812,I959804);
not I_56249 (I959829,I66148);
not I_56250 (I959846,I66136);
nor I_56251 (I959863,I959846,I66142);
nor I_56252 (I959476,I959812,I959863);
nor I_56253 (I959894,I959846,I66145);
and I_56254 (I959911,I959894,I66133);
or I_56255 (I959928,I959911,I66151);
DFFARX1 I_56256 (I959928,I3563,I959484,I959954,);
nor I_56257 (I959464,I959954,I959510);
not I_56258 (I959976,I959954);
and I_56259 (I959993,I959976,I959510);
nor I_56260 (I959458,I959535,I959993);
nand I_56261 (I960024,I959976,I959586);
nor I_56262 (I959452,I959846,I960024);
nand I_56263 (I959455,I959976,I959764);
nand I_56264 (I960069,I959586,I66136);
nor I_56265 (I959467,I959829,I960069);
not I_56266 (I960130,I3570);
DFFARX1 I_56267 (I706971,I3563,I960130,I960156,);
DFFARX1 I_56268 (I706965,I3563,I960130,I960173,);
not I_56269 (I960181,I960173);
not I_56270 (I960198,I706980);
nor I_56271 (I960215,I960198,I706965);
not I_56272 (I960232,I706974);
nor I_56273 (I960249,I960215,I706983);
nor I_56274 (I960266,I960173,I960249);
DFFARX1 I_56275 (I960266,I3563,I960130,I960116,);
nor I_56276 (I960297,I706983,I706965);
nand I_56277 (I960314,I960297,I706980);
DFFARX1 I_56278 (I960314,I3563,I960130,I960119,);
nor I_56279 (I960345,I960232,I706983);
nand I_56280 (I960362,I960345,I706968);
nor I_56281 (I960379,I960156,I960362);
DFFARX1 I_56282 (I960379,I3563,I960130,I960095,);
not I_56283 (I960410,I960362);
nand I_56284 (I960107,I960173,I960410);
DFFARX1 I_56285 (I960362,I3563,I960130,I960450,);
not I_56286 (I960458,I960450);
not I_56287 (I960475,I706983);
not I_56288 (I960492,I706977);
nor I_56289 (I960509,I960492,I706974);
nor I_56290 (I960122,I960458,I960509);
nor I_56291 (I960540,I960492,I706986);
and I_56292 (I960557,I960540,I706989);
or I_56293 (I960574,I960557,I706968);
DFFARX1 I_56294 (I960574,I3563,I960130,I960600,);
nor I_56295 (I960110,I960600,I960156);
not I_56296 (I960622,I960600);
and I_56297 (I960639,I960622,I960156);
nor I_56298 (I960104,I960181,I960639);
nand I_56299 (I960670,I960622,I960232);
nor I_56300 (I960098,I960492,I960670);
nand I_56301 (I960101,I960622,I960410);
nand I_56302 (I960715,I960232,I706977);
nor I_56303 (I960113,I960475,I960715);
not I_56304 (I960776,I3570);
DFFARX1 I_56305 (I754367,I3563,I960776,I960802,);
DFFARX1 I_56306 (I754361,I3563,I960776,I960819,);
not I_56307 (I960827,I960819);
not I_56308 (I960844,I754376);
nor I_56309 (I960861,I960844,I754361);
not I_56310 (I960878,I754370);
nor I_56311 (I960895,I960861,I754379);
nor I_56312 (I960912,I960819,I960895);
DFFARX1 I_56313 (I960912,I3563,I960776,I960762,);
nor I_56314 (I960943,I754379,I754361);
nand I_56315 (I960960,I960943,I754376);
DFFARX1 I_56316 (I960960,I3563,I960776,I960765,);
nor I_56317 (I960991,I960878,I754379);
nand I_56318 (I961008,I960991,I754364);
nor I_56319 (I961025,I960802,I961008);
DFFARX1 I_56320 (I961025,I3563,I960776,I960741,);
not I_56321 (I961056,I961008);
nand I_56322 (I960753,I960819,I961056);
DFFARX1 I_56323 (I961008,I3563,I960776,I961096,);
not I_56324 (I961104,I961096);
not I_56325 (I961121,I754379);
not I_56326 (I961138,I754373);
nor I_56327 (I961155,I961138,I754370);
nor I_56328 (I960768,I961104,I961155);
nor I_56329 (I961186,I961138,I754382);
and I_56330 (I961203,I961186,I754385);
or I_56331 (I961220,I961203,I754364);
DFFARX1 I_56332 (I961220,I3563,I960776,I961246,);
nor I_56333 (I960756,I961246,I960802);
not I_56334 (I961268,I961246);
and I_56335 (I961285,I961268,I960802);
nor I_56336 (I960750,I960827,I961285);
nand I_56337 (I961316,I961268,I960878);
nor I_56338 (I960744,I961138,I961316);
nand I_56339 (I960747,I961268,I961056);
nand I_56340 (I961361,I960878,I754373);
nor I_56341 (I960759,I961121,I961361);
not I_56342 (I961422,I3570);
DFFARX1 I_56343 (I1258939,I3563,I961422,I961448,);
DFFARX1 I_56344 (I1258945,I3563,I961422,I961465,);
not I_56345 (I961473,I961465);
not I_56346 (I961490,I1258942);
nor I_56347 (I961507,I961490,I1258921);
not I_56348 (I961524,I1258924);
nor I_56349 (I961541,I961507,I1258930);
nor I_56350 (I961558,I961465,I961541);
DFFARX1 I_56351 (I961558,I3563,I961422,I961408,);
nor I_56352 (I961589,I1258930,I1258921);
nand I_56353 (I961606,I961589,I1258942);
DFFARX1 I_56354 (I961606,I3563,I961422,I961411,);
nor I_56355 (I961637,I961524,I1258930);
nand I_56356 (I961654,I961637,I1258924);
nor I_56357 (I961671,I961448,I961654);
DFFARX1 I_56358 (I961671,I3563,I961422,I961387,);
not I_56359 (I961702,I961654);
nand I_56360 (I961399,I961465,I961702);
DFFARX1 I_56361 (I961654,I3563,I961422,I961742,);
not I_56362 (I961750,I961742);
not I_56363 (I961767,I1258930);
not I_56364 (I961784,I1258933);
nor I_56365 (I961801,I961784,I1258924);
nor I_56366 (I961414,I961750,I961801);
nor I_56367 (I961832,I961784,I1258921);
and I_56368 (I961849,I961832,I1258927);
or I_56369 (I961866,I961849,I1258936);
DFFARX1 I_56370 (I961866,I3563,I961422,I961892,);
nor I_56371 (I961402,I961892,I961448);
not I_56372 (I961914,I961892);
and I_56373 (I961931,I961914,I961448);
nor I_56374 (I961396,I961473,I961931);
nand I_56375 (I961962,I961914,I961524);
nor I_56376 (I961390,I961784,I961962);
nand I_56377 (I961393,I961914,I961702);
nand I_56378 (I962007,I961524,I1258933);
nor I_56379 (I961405,I961767,I962007);
not I_56380 (I962068,I3570);
DFFARX1 I_56381 (I724311,I3563,I962068,I962094,);
DFFARX1 I_56382 (I724305,I3563,I962068,I962111,);
not I_56383 (I962119,I962111);
not I_56384 (I962136,I724320);
nor I_56385 (I962153,I962136,I724305);
not I_56386 (I962170,I724314);
nor I_56387 (I962187,I962153,I724323);
nor I_56388 (I962204,I962111,I962187);
DFFARX1 I_56389 (I962204,I3563,I962068,I962054,);
nor I_56390 (I962235,I724323,I724305);
nand I_56391 (I962252,I962235,I724320);
DFFARX1 I_56392 (I962252,I3563,I962068,I962057,);
nor I_56393 (I962283,I962170,I724323);
nand I_56394 (I962300,I962283,I724308);
nor I_56395 (I962317,I962094,I962300);
DFFARX1 I_56396 (I962317,I3563,I962068,I962033,);
not I_56397 (I962348,I962300);
nand I_56398 (I962045,I962111,I962348);
DFFARX1 I_56399 (I962300,I3563,I962068,I962388,);
not I_56400 (I962396,I962388);
not I_56401 (I962413,I724323);
not I_56402 (I962430,I724317);
nor I_56403 (I962447,I962430,I724314);
nor I_56404 (I962060,I962396,I962447);
nor I_56405 (I962478,I962430,I724326);
and I_56406 (I962495,I962478,I724329);
or I_56407 (I962512,I962495,I724308);
DFFARX1 I_56408 (I962512,I3563,I962068,I962538,);
nor I_56409 (I962048,I962538,I962094);
not I_56410 (I962560,I962538);
and I_56411 (I962577,I962560,I962094);
nor I_56412 (I962042,I962119,I962577);
nand I_56413 (I962608,I962560,I962170);
nor I_56414 (I962036,I962430,I962608);
nand I_56415 (I962039,I962560,I962348);
nand I_56416 (I962653,I962170,I724317);
nor I_56417 (I962051,I962413,I962653);
not I_56418 (I962714,I3570);
DFFARX1 I_56419 (I799451,I3563,I962714,I962740,);
DFFARX1 I_56420 (I799445,I3563,I962714,I962757,);
not I_56421 (I962765,I962757);
not I_56422 (I962782,I799460);
nor I_56423 (I962799,I962782,I799445);
not I_56424 (I962816,I799454);
nor I_56425 (I962833,I962799,I799463);
nor I_56426 (I962850,I962757,I962833);
DFFARX1 I_56427 (I962850,I3563,I962714,I962700,);
nor I_56428 (I962881,I799463,I799445);
nand I_56429 (I962898,I962881,I799460);
DFFARX1 I_56430 (I962898,I3563,I962714,I962703,);
nor I_56431 (I962929,I962816,I799463);
nand I_56432 (I962946,I962929,I799448);
nor I_56433 (I962963,I962740,I962946);
DFFARX1 I_56434 (I962963,I3563,I962714,I962679,);
not I_56435 (I962994,I962946);
nand I_56436 (I962691,I962757,I962994);
DFFARX1 I_56437 (I962946,I3563,I962714,I963034,);
not I_56438 (I963042,I963034);
not I_56439 (I963059,I799463);
not I_56440 (I963076,I799457);
nor I_56441 (I963093,I963076,I799454);
nor I_56442 (I962706,I963042,I963093);
nor I_56443 (I963124,I963076,I799466);
and I_56444 (I963141,I963124,I799469);
or I_56445 (I963158,I963141,I799448);
DFFARX1 I_56446 (I963158,I3563,I962714,I963184,);
nor I_56447 (I962694,I963184,I962740);
not I_56448 (I963206,I963184);
and I_56449 (I963223,I963206,I962740);
nor I_56450 (I962688,I962765,I963223);
nand I_56451 (I963254,I963206,I962816);
nor I_56452 (I962682,I963076,I963254);
nand I_56453 (I962685,I963206,I962994);
nand I_56454 (I963299,I962816,I799457);
nor I_56455 (I962697,I963059,I963299);
not I_56456 (I963360,I3570);
DFFARX1 I_56457 (I1383888,I3563,I963360,I963386,);
DFFARX1 I_56458 (I1383912,I3563,I963360,I963403,);
not I_56459 (I963411,I963403);
not I_56460 (I963428,I1383894);
nor I_56461 (I963445,I963428,I1383903);
not I_56462 (I963462,I1383888);
nor I_56463 (I963479,I963445,I1383909);
nor I_56464 (I963496,I963403,I963479);
DFFARX1 I_56465 (I963496,I3563,I963360,I963346,);
nor I_56466 (I963527,I1383909,I1383903);
nand I_56467 (I963544,I963527,I1383894);
DFFARX1 I_56468 (I963544,I3563,I963360,I963349,);
nor I_56469 (I963575,I963462,I1383909);
nand I_56470 (I963592,I963575,I1383906);
nor I_56471 (I963609,I963386,I963592);
DFFARX1 I_56472 (I963609,I3563,I963360,I963325,);
not I_56473 (I963640,I963592);
nand I_56474 (I963337,I963403,I963640);
DFFARX1 I_56475 (I963592,I3563,I963360,I963680,);
not I_56476 (I963688,I963680);
not I_56477 (I963705,I1383909);
not I_56478 (I963722,I1383900);
nor I_56479 (I963739,I963722,I1383888);
nor I_56480 (I963352,I963688,I963739);
nor I_56481 (I963770,I963722,I1383891);
and I_56482 (I963787,I963770,I1383915);
or I_56483 (I963804,I963787,I1383897);
DFFARX1 I_56484 (I963804,I3563,I963360,I963830,);
nor I_56485 (I963340,I963830,I963386);
not I_56486 (I963852,I963830);
and I_56487 (I963869,I963852,I963386);
nor I_56488 (I963334,I963411,I963869);
nand I_56489 (I963900,I963852,I963462);
nor I_56490 (I963328,I963722,I963900);
nand I_56491 (I963331,I963852,I963640);
nand I_56492 (I963945,I963462,I1383900);
nor I_56493 (I963343,I963705,I963945);
not I_56494 (I964006,I3570);
DFFARX1 I_56495 (I670557,I3563,I964006,I964032,);
DFFARX1 I_56496 (I670551,I3563,I964006,I964049,);
not I_56497 (I964057,I964049);
not I_56498 (I964074,I670566);
nor I_56499 (I964091,I964074,I670551);
not I_56500 (I964108,I670560);
nor I_56501 (I964125,I964091,I670569);
nor I_56502 (I964142,I964049,I964125);
DFFARX1 I_56503 (I964142,I3563,I964006,I963992,);
nor I_56504 (I964173,I670569,I670551);
nand I_56505 (I964190,I964173,I670566);
DFFARX1 I_56506 (I964190,I3563,I964006,I963995,);
nor I_56507 (I964221,I964108,I670569);
nand I_56508 (I964238,I964221,I670554);
nor I_56509 (I964255,I964032,I964238);
DFFARX1 I_56510 (I964255,I3563,I964006,I963971,);
not I_56511 (I964286,I964238);
nand I_56512 (I963983,I964049,I964286);
DFFARX1 I_56513 (I964238,I3563,I964006,I964326,);
not I_56514 (I964334,I964326);
not I_56515 (I964351,I670569);
not I_56516 (I964368,I670563);
nor I_56517 (I964385,I964368,I670560);
nor I_56518 (I963998,I964334,I964385);
nor I_56519 (I964416,I964368,I670572);
and I_56520 (I964433,I964416,I670575);
or I_56521 (I964450,I964433,I670554);
DFFARX1 I_56522 (I964450,I3563,I964006,I964476,);
nor I_56523 (I963986,I964476,I964032);
not I_56524 (I964498,I964476);
and I_56525 (I964515,I964498,I964032);
nor I_56526 (I963980,I964057,I964515);
nand I_56527 (I964546,I964498,I964108);
nor I_56528 (I963974,I964368,I964546);
nand I_56529 (I963977,I964498,I964286);
nand I_56530 (I964591,I964108,I670563);
nor I_56531 (I963989,I964351,I964591);
not I_56532 (I964652,I3570);
DFFARX1 I_56533 (I727779,I3563,I964652,I964678,);
DFFARX1 I_56534 (I727773,I3563,I964652,I964695,);
not I_56535 (I964703,I964695);
not I_56536 (I964720,I727788);
nor I_56537 (I964737,I964720,I727773);
not I_56538 (I964754,I727782);
nor I_56539 (I964771,I964737,I727791);
nor I_56540 (I964788,I964695,I964771);
DFFARX1 I_56541 (I964788,I3563,I964652,I964638,);
nor I_56542 (I964819,I727791,I727773);
nand I_56543 (I964836,I964819,I727788);
DFFARX1 I_56544 (I964836,I3563,I964652,I964641,);
nor I_56545 (I964867,I964754,I727791);
nand I_56546 (I964884,I964867,I727776);
nor I_56547 (I964901,I964678,I964884);
DFFARX1 I_56548 (I964901,I3563,I964652,I964617,);
not I_56549 (I964932,I964884);
nand I_56550 (I964629,I964695,I964932);
DFFARX1 I_56551 (I964884,I3563,I964652,I964972,);
not I_56552 (I964980,I964972);
not I_56553 (I964997,I727791);
not I_56554 (I965014,I727785);
nor I_56555 (I965031,I965014,I727782);
nor I_56556 (I964644,I964980,I965031);
nor I_56557 (I965062,I965014,I727794);
and I_56558 (I965079,I965062,I727797);
or I_56559 (I965096,I965079,I727776);
DFFARX1 I_56560 (I965096,I3563,I964652,I965122,);
nor I_56561 (I964632,I965122,I964678);
not I_56562 (I965144,I965122);
and I_56563 (I965161,I965144,I964678);
nor I_56564 (I964626,I964703,I965161);
nand I_56565 (I965192,I965144,I964754);
nor I_56566 (I964620,I965014,I965192);
nand I_56567 (I964623,I965144,I964932);
nand I_56568 (I965237,I964754,I727785);
nor I_56569 (I964635,I964997,I965237);
not I_56570 (I965298,I3570);
DFFARX1 I_56571 (I1218173,I3563,I965298,I965324,);
DFFARX1 I_56572 (I1218155,I3563,I965298,I965341,);
not I_56573 (I965349,I965341);
not I_56574 (I965366,I1218164);
nor I_56575 (I965383,I965366,I1218176);
not I_56576 (I965400,I1218158);
nor I_56577 (I965417,I965383,I1218167);
nor I_56578 (I965434,I965341,I965417);
DFFARX1 I_56579 (I965434,I3563,I965298,I965284,);
nor I_56580 (I965465,I1218167,I1218176);
nand I_56581 (I965482,I965465,I1218164);
DFFARX1 I_56582 (I965482,I3563,I965298,I965287,);
nor I_56583 (I965513,I965400,I1218167);
nand I_56584 (I965530,I965513,I1218179);
nor I_56585 (I965547,I965324,I965530);
DFFARX1 I_56586 (I965547,I3563,I965298,I965263,);
not I_56587 (I965578,I965530);
nand I_56588 (I965275,I965341,I965578);
DFFARX1 I_56589 (I965530,I3563,I965298,I965618,);
not I_56590 (I965626,I965618);
not I_56591 (I965643,I1218167);
not I_56592 (I965660,I1218155);
nor I_56593 (I965677,I965660,I1218158);
nor I_56594 (I965290,I965626,I965677);
nor I_56595 (I965708,I965660,I1218161);
and I_56596 (I965725,I965708,I1218170);
or I_56597 (I965742,I965725,I1218158);
DFFARX1 I_56598 (I965742,I3563,I965298,I965768,);
nor I_56599 (I965278,I965768,I965324);
not I_56600 (I965790,I965768);
and I_56601 (I965807,I965790,I965324);
nor I_56602 (I965272,I965349,I965807);
nand I_56603 (I965838,I965790,I965400);
nor I_56604 (I965266,I965660,I965838);
nand I_56605 (I965269,I965790,I965578);
nand I_56606 (I965883,I965400,I1218155);
nor I_56607 (I965281,I965643,I965883);
not I_56608 (I965944,I3570);
DFFARX1 I_56609 (I1226265,I3563,I965944,I965970,);
DFFARX1 I_56610 (I1226247,I3563,I965944,I965987,);
not I_56611 (I965995,I965987);
not I_56612 (I966012,I1226256);
nor I_56613 (I966029,I966012,I1226268);
not I_56614 (I966046,I1226250);
nor I_56615 (I966063,I966029,I1226259);
nor I_56616 (I966080,I965987,I966063);
DFFARX1 I_56617 (I966080,I3563,I965944,I965930,);
nor I_56618 (I966111,I1226259,I1226268);
nand I_56619 (I966128,I966111,I1226256);
DFFARX1 I_56620 (I966128,I3563,I965944,I965933,);
nor I_56621 (I966159,I966046,I1226259);
nand I_56622 (I966176,I966159,I1226271);
nor I_56623 (I966193,I965970,I966176);
DFFARX1 I_56624 (I966193,I3563,I965944,I965909,);
not I_56625 (I966224,I966176);
nand I_56626 (I965921,I965987,I966224);
DFFARX1 I_56627 (I966176,I3563,I965944,I966264,);
not I_56628 (I966272,I966264);
not I_56629 (I966289,I1226259);
not I_56630 (I966306,I1226247);
nor I_56631 (I966323,I966306,I1226250);
nor I_56632 (I965936,I966272,I966323);
nor I_56633 (I966354,I966306,I1226253);
and I_56634 (I966371,I966354,I1226262);
or I_56635 (I966388,I966371,I1226250);
DFFARX1 I_56636 (I966388,I3563,I965944,I966414,);
nor I_56637 (I965924,I966414,I965970);
not I_56638 (I966436,I966414);
and I_56639 (I966453,I966436,I965970);
nor I_56640 (I965918,I965995,I966453);
nand I_56641 (I966484,I966436,I966046);
nor I_56642 (I965912,I966306,I966484);
nand I_56643 (I965915,I966436,I966224);
nand I_56644 (I966529,I966046,I1226247);
nor I_56645 (I965927,I966289,I966529);
not I_56646 (I966590,I3570);
DFFARX1 I_56647 (I772863,I3563,I966590,I966616,);
DFFARX1 I_56648 (I772857,I3563,I966590,I966633,);
not I_56649 (I966641,I966633);
not I_56650 (I966658,I772872);
nor I_56651 (I966675,I966658,I772857);
not I_56652 (I966692,I772866);
nor I_56653 (I966709,I966675,I772875);
nor I_56654 (I966726,I966633,I966709);
DFFARX1 I_56655 (I966726,I3563,I966590,I966576,);
nor I_56656 (I966757,I772875,I772857);
nand I_56657 (I966774,I966757,I772872);
DFFARX1 I_56658 (I966774,I3563,I966590,I966579,);
nor I_56659 (I966805,I966692,I772875);
nand I_56660 (I966822,I966805,I772860);
nor I_56661 (I966839,I966616,I966822);
DFFARX1 I_56662 (I966839,I3563,I966590,I966555,);
not I_56663 (I966870,I966822);
nand I_56664 (I966567,I966633,I966870);
DFFARX1 I_56665 (I966822,I3563,I966590,I966910,);
not I_56666 (I966918,I966910);
not I_56667 (I966935,I772875);
not I_56668 (I966952,I772869);
nor I_56669 (I966969,I966952,I772866);
nor I_56670 (I966582,I966918,I966969);
nor I_56671 (I967000,I966952,I772878);
and I_56672 (I967017,I967000,I772881);
or I_56673 (I967034,I967017,I772860);
DFFARX1 I_56674 (I967034,I3563,I966590,I967060,);
nor I_56675 (I966570,I967060,I966616);
not I_56676 (I967082,I967060);
and I_56677 (I967099,I967082,I966616);
nor I_56678 (I966564,I966641,I967099);
nand I_56679 (I967130,I967082,I966692);
nor I_56680 (I966558,I966952,I967130);
nand I_56681 (I966561,I967082,I966870);
nand I_56682 (I967175,I966692,I772869);
nor I_56683 (I966573,I966935,I967175);
not I_56684 (I967236,I3570);
DFFARX1 I_56685 (I1321864,I3563,I967236,I967262,);
DFFARX1 I_56686 (I1321858,I3563,I967236,I967279,);
not I_56687 (I967287,I967279);
not I_56688 (I967304,I1321867);
nor I_56689 (I967321,I967304,I1321879);
not I_56690 (I967338,I1321861);
nor I_56691 (I967355,I967321,I1321858);
nor I_56692 (I967372,I967279,I967355);
DFFARX1 I_56693 (I967372,I3563,I967236,I967222,);
nor I_56694 (I967403,I1321858,I1321879);
nand I_56695 (I967420,I967403,I1321867);
DFFARX1 I_56696 (I967420,I3563,I967236,I967225,);
nor I_56697 (I967451,I967338,I1321858);
nand I_56698 (I967468,I967451,I1321855);
nor I_56699 (I967485,I967262,I967468);
DFFARX1 I_56700 (I967485,I3563,I967236,I967201,);
not I_56701 (I967516,I967468);
nand I_56702 (I967213,I967279,I967516);
DFFARX1 I_56703 (I967468,I3563,I967236,I967556,);
not I_56704 (I967564,I967556);
not I_56705 (I967581,I1321858);
not I_56706 (I967598,I1321876);
nor I_56707 (I967615,I967598,I1321861);
nor I_56708 (I967228,I967564,I967615);
nor I_56709 (I967646,I967598,I1321870);
and I_56710 (I967663,I967646,I1321855);
or I_56711 (I967680,I967663,I1321873);
DFFARX1 I_56712 (I967680,I3563,I967236,I967706,);
nor I_56713 (I967216,I967706,I967262);
not I_56714 (I967728,I967706);
and I_56715 (I967745,I967728,I967262);
nor I_56716 (I967210,I967287,I967745);
nand I_56717 (I967776,I967728,I967338);
nor I_56718 (I967204,I967598,I967776);
nand I_56719 (I967207,I967728,I967516);
nand I_56720 (I967821,I967338,I1321876);
nor I_56721 (I967219,I967581,I967821);
not I_56722 (I967882,I3570);
DFFARX1 I_56723 (I491496,I3563,I967882,I967908,);
DFFARX1 I_56724 (I491493,I3563,I967882,I967925,);
not I_56725 (I967933,I967925);
not I_56726 (I967950,I491508);
nor I_56727 (I967967,I967950,I491511);
not I_56728 (I967984,I491499);
nor I_56729 (I968001,I967967,I491505);
nor I_56730 (I968018,I967925,I968001);
DFFARX1 I_56731 (I968018,I3563,I967882,I967868,);
nor I_56732 (I968049,I491505,I491511);
nand I_56733 (I968066,I968049,I491508);
DFFARX1 I_56734 (I968066,I3563,I967882,I967871,);
nor I_56735 (I968097,I967984,I491505);
nand I_56736 (I968114,I968097,I491517);
nor I_56737 (I968131,I967908,I968114);
DFFARX1 I_56738 (I968131,I3563,I967882,I967847,);
not I_56739 (I968162,I968114);
nand I_56740 (I967859,I967925,I968162);
DFFARX1 I_56741 (I968114,I3563,I967882,I968202,);
not I_56742 (I968210,I968202);
not I_56743 (I968227,I491505);
not I_56744 (I968244,I491490);
nor I_56745 (I968261,I968244,I491499);
nor I_56746 (I967874,I968210,I968261);
nor I_56747 (I968292,I968244,I491502);
and I_56748 (I968309,I968292,I491490);
or I_56749 (I968326,I968309,I491514);
DFFARX1 I_56750 (I968326,I3563,I967882,I968352,);
nor I_56751 (I967862,I968352,I967908);
not I_56752 (I968374,I968352);
and I_56753 (I968391,I968374,I967908);
nor I_56754 (I967856,I967933,I968391);
nand I_56755 (I968422,I968374,I967984);
nor I_56756 (I967850,I968244,I968422);
nand I_56757 (I967853,I968374,I968162);
nand I_56758 (I968467,I967984,I491490);
nor I_56759 (I967865,I968227,I968467);
not I_56760 (I968528,I3570);
DFFARX1 I_56761 (I289581,I3563,I968528,I968554,);
DFFARX1 I_56762 (I289587,I3563,I968528,I968571,);
not I_56763 (I968579,I968571);
not I_56764 (I968596,I289608);
nor I_56765 (I968613,I968596,I289596);
not I_56766 (I968630,I289605);
nor I_56767 (I968647,I968613,I289590);
nor I_56768 (I968664,I968571,I968647);
DFFARX1 I_56769 (I968664,I3563,I968528,I968514,);
nor I_56770 (I968695,I289590,I289596);
nand I_56771 (I968712,I968695,I289608);
DFFARX1 I_56772 (I968712,I3563,I968528,I968517,);
nor I_56773 (I968743,I968630,I289590);
nand I_56774 (I968760,I968743,I289581);
nor I_56775 (I968777,I968554,I968760);
DFFARX1 I_56776 (I968777,I3563,I968528,I968493,);
not I_56777 (I968808,I968760);
nand I_56778 (I968505,I968571,I968808);
DFFARX1 I_56779 (I968760,I3563,I968528,I968848,);
not I_56780 (I968856,I968848);
not I_56781 (I968873,I289590);
not I_56782 (I968890,I289593);
nor I_56783 (I968907,I968890,I289605);
nor I_56784 (I968520,I968856,I968907);
nor I_56785 (I968938,I968890,I289602);
and I_56786 (I968955,I968938,I289584);
or I_56787 (I968972,I968955,I289599);
DFFARX1 I_56788 (I968972,I3563,I968528,I968998,);
nor I_56789 (I968508,I968998,I968554);
not I_56790 (I969020,I968998);
and I_56791 (I969037,I969020,I968554);
nor I_56792 (I968502,I968579,I969037);
nand I_56793 (I969068,I969020,I968630);
nor I_56794 (I968496,I968890,I969068);
nand I_56795 (I968499,I969020,I968808);
nand I_56796 (I969113,I968630,I289593);
nor I_56797 (I968511,I968873,I969113);
not I_56798 (I969174,I3570);
DFFARX1 I_56799 (I2036,I3563,I969174,I969200,);
DFFARX1 I_56800 (I1436,I3563,I969174,I969217,);
not I_56801 (I969225,I969217);
not I_56802 (I969242,I1484);
nor I_56803 (I969259,I969242,I3276);
not I_56804 (I969276,I3076);
nor I_56805 (I969293,I969259,I2172);
nor I_56806 (I969310,I969217,I969293);
DFFARX1 I_56807 (I969310,I3563,I969174,I969160,);
nor I_56808 (I969341,I2172,I3276);
nand I_56809 (I969358,I969341,I1484);
DFFARX1 I_56810 (I969358,I3563,I969174,I969163,);
nor I_56811 (I969389,I969276,I2172);
nand I_56812 (I969406,I969389,I1972);
nor I_56813 (I969423,I969200,I969406);
DFFARX1 I_56814 (I969423,I3563,I969174,I969139,);
not I_56815 (I969454,I969406);
nand I_56816 (I969151,I969217,I969454);
DFFARX1 I_56817 (I969406,I3563,I969174,I969494,);
not I_56818 (I969502,I969494);
not I_56819 (I969519,I2172);
not I_56820 (I969536,I2668);
nor I_56821 (I969553,I969536,I3076);
nor I_56822 (I969166,I969502,I969553);
nor I_56823 (I969584,I969536,I3172);
and I_56824 (I969601,I969584,I2660);
or I_56825 (I969618,I969601,I2348);
DFFARX1 I_56826 (I969618,I3563,I969174,I969644,);
nor I_56827 (I969154,I969644,I969200);
not I_56828 (I969666,I969644);
and I_56829 (I969683,I969666,I969200);
nor I_56830 (I969148,I969225,I969683);
nand I_56831 (I969714,I969666,I969276);
nor I_56832 (I969142,I969536,I969714);
nand I_56833 (I969145,I969666,I969454);
nand I_56834 (I969759,I969276,I2668);
nor I_56835 (I969157,I969519,I969759);
not I_56836 (I969820,I3570);
DFFARX1 I_56837 (I603506,I3563,I969820,I969846,);
DFFARX1 I_56838 (I603518,I3563,I969820,I969863,);
not I_56839 (I969871,I969863);
not I_56840 (I969888,I603527);
nor I_56841 (I969905,I969888,I603503);
not I_56842 (I969922,I603521);
nor I_56843 (I969939,I969905,I603515);
nor I_56844 (I969956,I969863,I969939);
DFFARX1 I_56845 (I969956,I3563,I969820,I969806,);
nor I_56846 (I969987,I603515,I603503);
nand I_56847 (I970004,I969987,I603527);
DFFARX1 I_56848 (I970004,I3563,I969820,I969809,);
nor I_56849 (I970035,I969922,I603515);
nand I_56850 (I970052,I970035,I603509);
nor I_56851 (I970069,I969846,I970052);
DFFARX1 I_56852 (I970069,I3563,I969820,I969785,);
not I_56853 (I970100,I970052);
nand I_56854 (I969797,I969863,I970100);
DFFARX1 I_56855 (I970052,I3563,I969820,I970140,);
not I_56856 (I970148,I970140);
not I_56857 (I970165,I603515);
not I_56858 (I970182,I603524);
nor I_56859 (I970199,I970182,I603521);
nor I_56860 (I969812,I970148,I970199);
nor I_56861 (I970230,I970182,I603506);
and I_56862 (I970247,I970230,I603503);
or I_56863 (I970264,I970247,I603512);
DFFARX1 I_56864 (I970264,I3563,I969820,I970290,);
nor I_56865 (I969800,I970290,I969846);
not I_56866 (I970312,I970290);
and I_56867 (I970329,I970312,I969846);
nor I_56868 (I969794,I969871,I970329);
nand I_56869 (I970360,I970312,I969922);
nor I_56870 (I969788,I970182,I970360);
nand I_56871 (I969791,I970312,I970100);
nand I_56872 (I970405,I969922,I603524);
nor I_56873 (I969803,I970165,I970405);
not I_56874 (I970466,I3570);
DFFARX1 I_56875 (I287473,I3563,I970466,I970492,);
DFFARX1 I_56876 (I287479,I3563,I970466,I970509,);
not I_56877 (I970517,I970509);
not I_56878 (I970534,I287500);
nor I_56879 (I970551,I970534,I287488);
not I_56880 (I970568,I287497);
nor I_56881 (I970585,I970551,I287482);
nor I_56882 (I970602,I970509,I970585);
DFFARX1 I_56883 (I970602,I3563,I970466,I970452,);
nor I_56884 (I970633,I287482,I287488);
nand I_56885 (I970650,I970633,I287500);
DFFARX1 I_56886 (I970650,I3563,I970466,I970455,);
nor I_56887 (I970681,I970568,I287482);
nand I_56888 (I970698,I970681,I287473);
nor I_56889 (I970715,I970492,I970698);
DFFARX1 I_56890 (I970715,I3563,I970466,I970431,);
not I_56891 (I970746,I970698);
nand I_56892 (I970443,I970509,I970746);
DFFARX1 I_56893 (I970698,I3563,I970466,I970786,);
not I_56894 (I970794,I970786);
not I_56895 (I970811,I287482);
not I_56896 (I970828,I287485);
nor I_56897 (I970845,I970828,I287497);
nor I_56898 (I970458,I970794,I970845);
nor I_56899 (I970876,I970828,I287494);
and I_56900 (I970893,I970876,I287476);
or I_56901 (I970910,I970893,I287491);
DFFARX1 I_56902 (I970910,I3563,I970466,I970936,);
nor I_56903 (I970446,I970936,I970492);
not I_56904 (I970958,I970936);
and I_56905 (I970975,I970958,I970492);
nor I_56906 (I970440,I970517,I970975);
nand I_56907 (I971006,I970958,I970568);
nor I_56908 (I970434,I970828,I971006);
nand I_56909 (I970437,I970958,I970746);
nand I_56910 (I971051,I970568,I287485);
nor I_56911 (I970449,I970811,I971051);
not I_56912 (I971112,I3570);
DFFARX1 I_56913 (I589634,I3563,I971112,I971138,);
DFFARX1 I_56914 (I589646,I3563,I971112,I971155,);
not I_56915 (I971163,I971155);
not I_56916 (I971180,I589655);
nor I_56917 (I971197,I971180,I589631);
not I_56918 (I971214,I589649);
nor I_56919 (I971231,I971197,I589643);
nor I_56920 (I971248,I971155,I971231);
DFFARX1 I_56921 (I971248,I3563,I971112,I971098,);
nor I_56922 (I971279,I589643,I589631);
nand I_56923 (I971296,I971279,I589655);
DFFARX1 I_56924 (I971296,I3563,I971112,I971101,);
nor I_56925 (I971327,I971214,I589643);
nand I_56926 (I971344,I971327,I589637);
nor I_56927 (I971361,I971138,I971344);
DFFARX1 I_56928 (I971361,I3563,I971112,I971077,);
not I_56929 (I971392,I971344);
nand I_56930 (I971089,I971155,I971392);
DFFARX1 I_56931 (I971344,I3563,I971112,I971432,);
not I_56932 (I971440,I971432);
not I_56933 (I971457,I589643);
not I_56934 (I971474,I589652);
nor I_56935 (I971491,I971474,I589649);
nor I_56936 (I971104,I971440,I971491);
nor I_56937 (I971522,I971474,I589634);
and I_56938 (I971539,I971522,I589631);
or I_56939 (I971556,I971539,I589640);
DFFARX1 I_56940 (I971556,I3563,I971112,I971582,);
nor I_56941 (I971092,I971582,I971138);
not I_56942 (I971604,I971582);
and I_56943 (I971621,I971604,I971138);
nor I_56944 (I971086,I971163,I971621);
nand I_56945 (I971652,I971604,I971214);
nor I_56946 (I971080,I971474,I971652);
nand I_56947 (I971083,I971604,I971392);
nand I_56948 (I971697,I971214,I589652);
nor I_56949 (I971095,I971457,I971697);
not I_56950 (I971758,I3570);
DFFARX1 I_56951 (I330160,I3563,I971758,I971784,);
DFFARX1 I_56952 (I330166,I3563,I971758,I971801,);
not I_56953 (I971809,I971801);
not I_56954 (I971826,I330187);
nor I_56955 (I971843,I971826,I330175);
not I_56956 (I971860,I330184);
nor I_56957 (I971877,I971843,I330169);
nor I_56958 (I971894,I971801,I971877);
DFFARX1 I_56959 (I971894,I3563,I971758,I971744,);
nor I_56960 (I971925,I330169,I330175);
nand I_56961 (I971942,I971925,I330187);
DFFARX1 I_56962 (I971942,I3563,I971758,I971747,);
nor I_56963 (I971973,I971860,I330169);
nand I_56964 (I971990,I971973,I330160);
nor I_56965 (I972007,I971784,I971990);
DFFARX1 I_56966 (I972007,I3563,I971758,I971723,);
not I_56967 (I972038,I971990);
nand I_56968 (I971735,I971801,I972038);
DFFARX1 I_56969 (I971990,I3563,I971758,I972078,);
not I_56970 (I972086,I972078);
not I_56971 (I972103,I330169);
not I_56972 (I972120,I330172);
nor I_56973 (I972137,I972120,I330184);
nor I_56974 (I971750,I972086,I972137);
nor I_56975 (I972168,I972120,I330181);
and I_56976 (I972185,I972168,I330163);
or I_56977 (I972202,I972185,I330178);
DFFARX1 I_56978 (I972202,I3563,I971758,I972228,);
nor I_56979 (I971738,I972228,I971784);
not I_56980 (I972250,I972228);
and I_56981 (I972267,I972250,I971784);
nor I_56982 (I971732,I971809,I972267);
nand I_56983 (I972298,I972250,I971860);
nor I_56984 (I971726,I972120,I972298);
nand I_56985 (I971729,I972250,I972038);
nand I_56986 (I972343,I971860,I330172);
nor I_56987 (I971741,I972103,I972343);
not I_56988 (I972404,I3570);
DFFARX1 I_56989 (I412899,I3563,I972404,I972430,);
DFFARX1 I_56990 (I412905,I3563,I972404,I972447,);
not I_56991 (I972455,I972447);
not I_56992 (I972472,I412926);
nor I_56993 (I972489,I972472,I412914);
not I_56994 (I972506,I412923);
nor I_56995 (I972523,I972489,I412908);
nor I_56996 (I972540,I972447,I972523);
DFFARX1 I_56997 (I972540,I3563,I972404,I972390,);
nor I_56998 (I972571,I412908,I412914);
nand I_56999 (I972588,I972571,I412926);
DFFARX1 I_57000 (I972588,I3563,I972404,I972393,);
nor I_57001 (I972619,I972506,I412908);
nand I_57002 (I972636,I972619,I412899);
nor I_57003 (I972653,I972430,I972636);
DFFARX1 I_57004 (I972653,I3563,I972404,I972369,);
not I_57005 (I972684,I972636);
nand I_57006 (I972381,I972447,I972684);
DFFARX1 I_57007 (I972636,I3563,I972404,I972724,);
not I_57008 (I972732,I972724);
not I_57009 (I972749,I412908);
not I_57010 (I972766,I412911);
nor I_57011 (I972783,I972766,I412923);
nor I_57012 (I972396,I972732,I972783);
nor I_57013 (I972814,I972766,I412920);
and I_57014 (I972831,I972814,I412902);
or I_57015 (I972848,I972831,I412917);
DFFARX1 I_57016 (I972848,I3563,I972404,I972874,);
nor I_57017 (I972384,I972874,I972430);
not I_57018 (I972896,I972874);
and I_57019 (I972913,I972896,I972430);
nor I_57020 (I972378,I972455,I972913);
nand I_57021 (I972944,I972896,I972506);
nor I_57022 (I972372,I972766,I972944);
nand I_57023 (I972375,I972896,I972684);
nand I_57024 (I972989,I972506,I412911);
nor I_57025 (I972387,I972749,I972989);
not I_57026 (I973050,I3570);
DFFARX1 I_57027 (I227979,I3563,I973050,I973076,);
DFFARX1 I_57028 (I227991,I3563,I973050,I973093,);
not I_57029 (I973101,I973093);
not I_57030 (I973118,I227997);
nor I_57031 (I973135,I973118,I227982);
not I_57032 (I973152,I227973);
nor I_57033 (I973169,I973135,I227994);
nor I_57034 (I973186,I973093,I973169);
DFFARX1 I_57035 (I973186,I3563,I973050,I973036,);
nor I_57036 (I973217,I227994,I227982);
nand I_57037 (I973234,I973217,I227997);
DFFARX1 I_57038 (I973234,I3563,I973050,I973039,);
nor I_57039 (I973265,I973152,I227994);
nand I_57040 (I973282,I973265,I227976);
nor I_57041 (I973299,I973076,I973282);
DFFARX1 I_57042 (I973299,I3563,I973050,I973015,);
not I_57043 (I973330,I973282);
nand I_57044 (I973027,I973093,I973330);
DFFARX1 I_57045 (I973282,I3563,I973050,I973370,);
not I_57046 (I973378,I973370);
not I_57047 (I973395,I227994);
not I_57048 (I973412,I227985);
nor I_57049 (I973429,I973412,I227973);
nor I_57050 (I973042,I973378,I973429);
nor I_57051 (I973460,I973412,I227988);
and I_57052 (I973477,I973460,I227976);
or I_57053 (I973494,I973477,I227973);
DFFARX1 I_57054 (I973494,I3563,I973050,I973520,);
nor I_57055 (I973030,I973520,I973076);
not I_57056 (I973542,I973520);
and I_57057 (I973559,I973542,I973076);
nor I_57058 (I973024,I973101,I973559);
nand I_57059 (I973590,I973542,I973152);
nor I_57060 (I973018,I973412,I973590);
nand I_57061 (I973021,I973542,I973330);
nand I_57062 (I973635,I973152,I227985);
nor I_57063 (I973033,I973395,I973635);
not I_57064 (I973696,I3570);
DFFARX1 I_57065 (I769395,I3563,I973696,I973722,);
DFFARX1 I_57066 (I769389,I3563,I973696,I973739,);
not I_57067 (I973747,I973739);
not I_57068 (I973764,I769404);
nor I_57069 (I973781,I973764,I769389);
not I_57070 (I973798,I769398);
nor I_57071 (I973815,I973781,I769407);
nor I_57072 (I973832,I973739,I973815);
DFFARX1 I_57073 (I973832,I3563,I973696,I973682,);
nor I_57074 (I973863,I769407,I769389);
nand I_57075 (I973880,I973863,I769404);
DFFARX1 I_57076 (I973880,I3563,I973696,I973685,);
nor I_57077 (I973911,I973798,I769407);
nand I_57078 (I973928,I973911,I769392);
nor I_57079 (I973945,I973722,I973928);
DFFARX1 I_57080 (I973945,I3563,I973696,I973661,);
not I_57081 (I973976,I973928);
nand I_57082 (I973673,I973739,I973976);
DFFARX1 I_57083 (I973928,I3563,I973696,I974016,);
not I_57084 (I974024,I974016);
not I_57085 (I974041,I769407);
not I_57086 (I974058,I769401);
nor I_57087 (I974075,I974058,I769398);
nor I_57088 (I973688,I974024,I974075);
nor I_57089 (I974106,I974058,I769410);
and I_57090 (I974123,I974106,I769413);
or I_57091 (I974140,I974123,I769392);
DFFARX1 I_57092 (I974140,I3563,I973696,I974166,);
nor I_57093 (I973676,I974166,I973722);
not I_57094 (I974188,I974166);
and I_57095 (I974205,I974188,I973722);
nor I_57096 (I973670,I973747,I974205);
nand I_57097 (I974236,I974188,I973798);
nor I_57098 (I973664,I974058,I974236);
nand I_57099 (I973667,I974188,I973976);
nand I_57100 (I974281,I973798,I769401);
nor I_57101 (I973679,I974041,I974281);
not I_57102 (I974342,I3570);
DFFARX1 I_57103 (I664199,I3563,I974342,I974368,);
DFFARX1 I_57104 (I664193,I3563,I974342,I974385,);
not I_57105 (I974393,I974385);
not I_57106 (I974410,I664208);
nor I_57107 (I974427,I974410,I664193);
not I_57108 (I974444,I664202);
nor I_57109 (I974461,I974427,I664211);
nor I_57110 (I974478,I974385,I974461);
DFFARX1 I_57111 (I974478,I3563,I974342,I974328,);
nor I_57112 (I974509,I664211,I664193);
nand I_57113 (I974526,I974509,I664208);
DFFARX1 I_57114 (I974526,I3563,I974342,I974331,);
nor I_57115 (I974557,I974444,I664211);
nand I_57116 (I974574,I974557,I664196);
nor I_57117 (I974591,I974368,I974574);
DFFARX1 I_57118 (I974591,I3563,I974342,I974307,);
not I_57119 (I974622,I974574);
nand I_57120 (I974319,I974385,I974622);
DFFARX1 I_57121 (I974574,I3563,I974342,I974662,);
not I_57122 (I974670,I974662);
not I_57123 (I974687,I664211);
not I_57124 (I974704,I664205);
nor I_57125 (I974721,I974704,I664202);
nor I_57126 (I974334,I974670,I974721);
nor I_57127 (I974752,I974704,I664214);
and I_57128 (I974769,I974752,I664217);
or I_57129 (I974786,I974769,I664196);
DFFARX1 I_57130 (I974786,I3563,I974342,I974812,);
nor I_57131 (I974322,I974812,I974368);
not I_57132 (I974834,I974812);
and I_57133 (I974851,I974834,I974368);
nor I_57134 (I974316,I974393,I974851);
nand I_57135 (I974882,I974834,I974444);
nor I_57136 (I974310,I974704,I974882);
nand I_57137 (I974313,I974834,I974622);
nand I_57138 (I974927,I974444,I664205);
nor I_57139 (I974325,I974687,I974927);
not I_57140 (I974988,I3570);
DFFARX1 I_57141 (I385495,I3563,I974988,I975014,);
DFFARX1 I_57142 (I385501,I3563,I974988,I975031,);
not I_57143 (I975039,I975031);
not I_57144 (I975056,I385522);
nor I_57145 (I975073,I975056,I385510);
not I_57146 (I975090,I385519);
nor I_57147 (I975107,I975073,I385504);
nor I_57148 (I975124,I975031,I975107);
DFFARX1 I_57149 (I975124,I3563,I974988,I974974,);
nor I_57150 (I975155,I385504,I385510);
nand I_57151 (I975172,I975155,I385522);
DFFARX1 I_57152 (I975172,I3563,I974988,I974977,);
nor I_57153 (I975203,I975090,I385504);
nand I_57154 (I975220,I975203,I385495);
nor I_57155 (I975237,I975014,I975220);
DFFARX1 I_57156 (I975237,I3563,I974988,I974953,);
not I_57157 (I975268,I975220);
nand I_57158 (I974965,I975031,I975268);
DFFARX1 I_57159 (I975220,I3563,I974988,I975308,);
not I_57160 (I975316,I975308);
not I_57161 (I975333,I385504);
not I_57162 (I975350,I385507);
nor I_57163 (I975367,I975350,I385519);
nor I_57164 (I974980,I975316,I975367);
nor I_57165 (I975398,I975350,I385516);
and I_57166 (I975415,I975398,I385498);
or I_57167 (I975432,I975415,I385513);
DFFARX1 I_57168 (I975432,I3563,I974988,I975458,);
nor I_57169 (I974968,I975458,I975014);
not I_57170 (I975480,I975458);
and I_57171 (I975497,I975480,I975014);
nor I_57172 (I974962,I975039,I975497);
nand I_57173 (I975528,I975480,I975090);
nor I_57174 (I974956,I975350,I975528);
nand I_57175 (I974959,I975480,I975268);
nand I_57176 (I975573,I975090,I385507);
nor I_57177 (I974971,I975333,I975573);
not I_57178 (I975634,I3570);
DFFARX1 I_57179 (I585588,I3563,I975634,I975660,);
DFFARX1 I_57180 (I585600,I3563,I975634,I975677,);
not I_57181 (I975685,I975677);
not I_57182 (I975702,I585609);
nor I_57183 (I975719,I975702,I585585);
not I_57184 (I975736,I585603);
nor I_57185 (I975753,I975719,I585597);
nor I_57186 (I975770,I975677,I975753);
DFFARX1 I_57187 (I975770,I3563,I975634,I975620,);
nor I_57188 (I975801,I585597,I585585);
nand I_57189 (I975818,I975801,I585609);
DFFARX1 I_57190 (I975818,I3563,I975634,I975623,);
nor I_57191 (I975849,I975736,I585597);
nand I_57192 (I975866,I975849,I585591);
nor I_57193 (I975883,I975660,I975866);
DFFARX1 I_57194 (I975883,I3563,I975634,I975599,);
not I_57195 (I975914,I975866);
nand I_57196 (I975611,I975677,I975914);
DFFARX1 I_57197 (I975866,I3563,I975634,I975954,);
not I_57198 (I975962,I975954);
not I_57199 (I975979,I585597);
not I_57200 (I975996,I585606);
nor I_57201 (I976013,I975996,I585603);
nor I_57202 (I975626,I975962,I976013);
nor I_57203 (I976044,I975996,I585588);
and I_57204 (I976061,I976044,I585585);
or I_57205 (I976078,I976061,I585594);
DFFARX1 I_57206 (I976078,I3563,I975634,I976104,);
nor I_57207 (I975614,I976104,I975660);
not I_57208 (I976126,I976104);
and I_57209 (I976143,I976126,I975660);
nor I_57210 (I975608,I975685,I976143);
nand I_57211 (I976174,I976126,I975736);
nor I_57212 (I975602,I975996,I976174);
nand I_57213 (I975605,I976126,I975914);
nand I_57214 (I976219,I975736,I585606);
nor I_57215 (I975617,I975979,I976219);
not I_57216 (I976280,I3570);
DFFARX1 I_57217 (I674603,I3563,I976280,I976306,);
DFFARX1 I_57218 (I674597,I3563,I976280,I976323,);
not I_57219 (I976331,I976323);
not I_57220 (I976348,I674612);
nor I_57221 (I976365,I976348,I674597);
not I_57222 (I976382,I674606);
nor I_57223 (I976399,I976365,I674615);
nor I_57224 (I976416,I976323,I976399);
DFFARX1 I_57225 (I976416,I3563,I976280,I976266,);
nor I_57226 (I976447,I674615,I674597);
nand I_57227 (I976464,I976447,I674612);
DFFARX1 I_57228 (I976464,I3563,I976280,I976269,);
nor I_57229 (I976495,I976382,I674615);
nand I_57230 (I976512,I976495,I674600);
nor I_57231 (I976529,I976306,I976512);
DFFARX1 I_57232 (I976529,I3563,I976280,I976245,);
not I_57233 (I976560,I976512);
nand I_57234 (I976257,I976323,I976560);
DFFARX1 I_57235 (I976512,I3563,I976280,I976600,);
not I_57236 (I976608,I976600);
not I_57237 (I976625,I674615);
not I_57238 (I976642,I674609);
nor I_57239 (I976659,I976642,I674606);
nor I_57240 (I976272,I976608,I976659);
nor I_57241 (I976690,I976642,I674618);
and I_57242 (I976707,I976690,I674621);
or I_57243 (I976724,I976707,I674600);
DFFARX1 I_57244 (I976724,I3563,I976280,I976750,);
nor I_57245 (I976260,I976750,I976306);
not I_57246 (I976772,I976750);
and I_57247 (I976789,I976772,I976306);
nor I_57248 (I976254,I976331,I976789);
nand I_57249 (I976820,I976772,I976382);
nor I_57250 (I976248,I976642,I976820);
nand I_57251 (I976251,I976772,I976560);
nand I_57252 (I976865,I976382,I674609);
nor I_57253 (I976263,I976625,I976865);
not I_57254 (I976926,I3570);
DFFARX1 I_57255 (I677493,I3563,I976926,I976952,);
DFFARX1 I_57256 (I677487,I3563,I976926,I976969,);
not I_57257 (I976977,I976969);
not I_57258 (I976994,I677502);
nor I_57259 (I977011,I976994,I677487);
not I_57260 (I977028,I677496);
nor I_57261 (I977045,I977011,I677505);
nor I_57262 (I977062,I976969,I977045);
DFFARX1 I_57263 (I977062,I3563,I976926,I976912,);
nor I_57264 (I977093,I677505,I677487);
nand I_57265 (I977110,I977093,I677502);
DFFARX1 I_57266 (I977110,I3563,I976926,I976915,);
nor I_57267 (I977141,I977028,I677505);
nand I_57268 (I977158,I977141,I677490);
nor I_57269 (I977175,I976952,I977158);
DFFARX1 I_57270 (I977175,I3563,I976926,I976891,);
not I_57271 (I977206,I977158);
nand I_57272 (I976903,I976969,I977206);
DFFARX1 I_57273 (I977158,I3563,I976926,I977246,);
not I_57274 (I977254,I977246);
not I_57275 (I977271,I677505);
not I_57276 (I977288,I677499);
nor I_57277 (I977305,I977288,I677496);
nor I_57278 (I976918,I977254,I977305);
nor I_57279 (I977336,I977288,I677508);
and I_57280 (I977353,I977336,I677511);
or I_57281 (I977370,I977353,I677490);
DFFARX1 I_57282 (I977370,I3563,I976926,I977396,);
nor I_57283 (I976906,I977396,I976952);
not I_57284 (I977418,I977396);
and I_57285 (I977435,I977418,I976952);
nor I_57286 (I976900,I976977,I977435);
nand I_57287 (I977466,I977418,I977028);
nor I_57288 (I976894,I977288,I977466);
nand I_57289 (I976897,I977418,I977206);
nand I_57290 (I977511,I977028,I677499);
nor I_57291 (I976909,I977271,I977511);
not I_57292 (I977572,I3570);
DFFARX1 I_57293 (I396562,I3563,I977572,I977598,);
DFFARX1 I_57294 (I396568,I3563,I977572,I977615,);
not I_57295 (I977623,I977615);
not I_57296 (I977640,I396589);
nor I_57297 (I977657,I977640,I396577);
not I_57298 (I977674,I396586);
nor I_57299 (I977691,I977657,I396571);
nor I_57300 (I977708,I977615,I977691);
DFFARX1 I_57301 (I977708,I3563,I977572,I977558,);
nor I_57302 (I977739,I396571,I396577);
nand I_57303 (I977756,I977739,I396589);
DFFARX1 I_57304 (I977756,I3563,I977572,I977561,);
nor I_57305 (I977787,I977674,I396571);
nand I_57306 (I977804,I977787,I396562);
nor I_57307 (I977821,I977598,I977804);
DFFARX1 I_57308 (I977821,I3563,I977572,I977537,);
not I_57309 (I977852,I977804);
nand I_57310 (I977549,I977615,I977852);
DFFARX1 I_57311 (I977804,I3563,I977572,I977892,);
not I_57312 (I977900,I977892);
not I_57313 (I977917,I396571);
not I_57314 (I977934,I396574);
nor I_57315 (I977951,I977934,I396586);
nor I_57316 (I977564,I977900,I977951);
nor I_57317 (I977982,I977934,I396583);
and I_57318 (I977999,I977982,I396565);
or I_57319 (I978016,I977999,I396580);
DFFARX1 I_57320 (I978016,I3563,I977572,I978042,);
nor I_57321 (I977552,I978042,I977598);
not I_57322 (I978064,I978042);
and I_57323 (I978081,I978064,I977598);
nor I_57324 (I977546,I977623,I978081);
nand I_57325 (I978112,I978064,I977674);
nor I_57326 (I977540,I977934,I978112);
nand I_57327 (I977543,I978064,I977852);
nand I_57328 (I978157,I977674,I396574);
nor I_57329 (I977555,I977917,I978157);
not I_57330 (I978218,I3570);
DFFARX1 I_57331 (I1225109,I3563,I978218,I978244,);
DFFARX1 I_57332 (I1225091,I3563,I978218,I978261,);
not I_57333 (I978269,I978261);
not I_57334 (I978286,I1225100);
nor I_57335 (I978303,I978286,I1225112);
not I_57336 (I978320,I1225094);
nor I_57337 (I978337,I978303,I1225103);
nor I_57338 (I978354,I978261,I978337);
DFFARX1 I_57339 (I978354,I3563,I978218,I978204,);
nor I_57340 (I978385,I1225103,I1225112);
nand I_57341 (I978402,I978385,I1225100);
DFFARX1 I_57342 (I978402,I3563,I978218,I978207,);
nor I_57343 (I978433,I978320,I1225103);
nand I_57344 (I978450,I978433,I1225115);
nor I_57345 (I978467,I978244,I978450);
DFFARX1 I_57346 (I978467,I3563,I978218,I978183,);
not I_57347 (I978498,I978450);
nand I_57348 (I978195,I978261,I978498);
DFFARX1 I_57349 (I978450,I3563,I978218,I978538,);
not I_57350 (I978546,I978538);
not I_57351 (I978563,I1225103);
not I_57352 (I978580,I1225091);
nor I_57353 (I978597,I978580,I1225094);
nor I_57354 (I978210,I978546,I978597);
nor I_57355 (I978628,I978580,I1225097);
and I_57356 (I978645,I978628,I1225106);
or I_57357 (I978662,I978645,I1225094);
DFFARX1 I_57358 (I978662,I3563,I978218,I978688,);
nor I_57359 (I978198,I978688,I978244);
not I_57360 (I978710,I978688);
and I_57361 (I978727,I978710,I978244);
nor I_57362 (I978192,I978269,I978727);
nand I_57363 (I978758,I978710,I978320);
nor I_57364 (I978186,I978580,I978758);
nand I_57365 (I978189,I978710,I978498);
nand I_57366 (I978803,I978320,I1225091);
nor I_57367 (I978201,I978563,I978803);
not I_57368 (I978864,I3570);
DFFARX1 I_57369 (I522504,I3563,I978864,I978890,);
DFFARX1 I_57370 (I522501,I3563,I978864,I978907,);
not I_57371 (I978915,I978907);
not I_57372 (I978932,I522516);
nor I_57373 (I978949,I978932,I522519);
not I_57374 (I978966,I522507);
nor I_57375 (I978983,I978949,I522513);
nor I_57376 (I979000,I978907,I978983);
DFFARX1 I_57377 (I979000,I3563,I978864,I978850,);
nor I_57378 (I979031,I522513,I522519);
nand I_57379 (I979048,I979031,I522516);
DFFARX1 I_57380 (I979048,I3563,I978864,I978853,);
nor I_57381 (I979079,I978966,I522513);
nand I_57382 (I979096,I979079,I522525);
nor I_57383 (I979113,I978890,I979096);
DFFARX1 I_57384 (I979113,I3563,I978864,I978829,);
not I_57385 (I979144,I979096);
nand I_57386 (I978841,I978907,I979144);
DFFARX1 I_57387 (I979096,I3563,I978864,I979184,);
not I_57388 (I979192,I979184);
not I_57389 (I979209,I522513);
not I_57390 (I979226,I522498);
nor I_57391 (I979243,I979226,I522507);
nor I_57392 (I978856,I979192,I979243);
nor I_57393 (I979274,I979226,I522510);
and I_57394 (I979291,I979274,I522498);
or I_57395 (I979308,I979291,I522522);
DFFARX1 I_57396 (I979308,I3563,I978864,I979334,);
nor I_57397 (I978844,I979334,I978890);
not I_57398 (I979356,I979334);
and I_57399 (I979373,I979356,I978890);
nor I_57400 (I978838,I978915,I979373);
nand I_57401 (I979404,I979356,I978966);
nor I_57402 (I978832,I979226,I979404);
nand I_57403 (I978835,I979356,I979144);
nand I_57404 (I979449,I978966,I522498);
nor I_57405 (I978847,I979209,I979449);
not I_57406 (I979510,I3570);
DFFARX1 I_57407 (I42945,I3563,I979510,I979536,);
DFFARX1 I_57408 (I42951,I3563,I979510,I979553,);
not I_57409 (I979561,I979553);
not I_57410 (I979578,I42945);
nor I_57411 (I979595,I979578,I42957);
not I_57412 (I979612,I42969);
nor I_57413 (I979629,I979595,I42963);
nor I_57414 (I979646,I979553,I979629);
DFFARX1 I_57415 (I979646,I3563,I979510,I979496,);
nor I_57416 (I979677,I42963,I42957);
nand I_57417 (I979694,I979677,I42945);
DFFARX1 I_57418 (I979694,I3563,I979510,I979499,);
nor I_57419 (I979725,I979612,I42963);
nand I_57420 (I979742,I979725,I42948);
nor I_57421 (I979759,I979536,I979742);
DFFARX1 I_57422 (I979759,I3563,I979510,I979475,);
not I_57423 (I979790,I979742);
nand I_57424 (I979487,I979553,I979790);
DFFARX1 I_57425 (I979742,I3563,I979510,I979830,);
not I_57426 (I979838,I979830);
not I_57427 (I979855,I42963);
not I_57428 (I979872,I42948);
nor I_57429 (I979889,I979872,I42969);
nor I_57430 (I979502,I979838,I979889);
nor I_57431 (I979920,I979872,I42966);
and I_57432 (I979937,I979920,I42960);
or I_57433 (I979954,I979937,I42954);
DFFARX1 I_57434 (I979954,I3563,I979510,I979980,);
nor I_57435 (I979490,I979980,I979536);
not I_57436 (I980002,I979980);
and I_57437 (I980019,I980002,I979536);
nor I_57438 (I979484,I979561,I980019);
nand I_57439 (I980050,I980002,I979612);
nor I_57440 (I979478,I979872,I980050);
nand I_57441 (I979481,I980002,I979790);
nand I_57442 (I980095,I979612,I42948);
nor I_57443 (I979493,I979855,I980095);
not I_57444 (I980156,I3570);
DFFARX1 I_57445 (I71930,I3563,I980156,I980182,);
DFFARX1 I_57446 (I71936,I3563,I980156,I980199,);
not I_57447 (I980207,I980199);
not I_57448 (I980224,I71954);
nor I_57449 (I980241,I980224,I71933);
not I_57450 (I980258,I71939);
nor I_57451 (I980275,I980241,I71945);
nor I_57452 (I980292,I980199,I980275);
DFFARX1 I_57453 (I980292,I3563,I980156,I980142,);
nor I_57454 (I980323,I71945,I71933);
nand I_57455 (I980340,I980323,I71954);
DFFARX1 I_57456 (I980340,I3563,I980156,I980145,);
nor I_57457 (I980371,I980258,I71945);
nand I_57458 (I980388,I980371,I71951);
nor I_57459 (I980405,I980182,I980388);
DFFARX1 I_57460 (I980405,I3563,I980156,I980121,);
not I_57461 (I980436,I980388);
nand I_57462 (I980133,I980199,I980436);
DFFARX1 I_57463 (I980388,I3563,I980156,I980476,);
not I_57464 (I980484,I980476);
not I_57465 (I980501,I71945);
not I_57466 (I980518,I71933);
nor I_57467 (I980535,I980518,I71939);
nor I_57468 (I980148,I980484,I980535);
nor I_57469 (I980566,I980518,I71942);
and I_57470 (I980583,I980566,I71930);
or I_57471 (I980600,I980583,I71948);
DFFARX1 I_57472 (I980600,I3563,I980156,I980626,);
nor I_57473 (I980136,I980626,I980182);
not I_57474 (I980648,I980626);
and I_57475 (I980665,I980648,I980182);
nor I_57476 (I980130,I980207,I980665);
nand I_57477 (I980696,I980648,I980258);
nor I_57478 (I980124,I980518,I980696);
nand I_57479 (I980127,I980648,I980436);
nand I_57480 (I980741,I980258,I71933);
nor I_57481 (I980139,I980501,I980741);
not I_57482 (I980802,I3570);
DFFARX1 I_57483 (I65079,I3563,I980802,I980828,);
DFFARX1 I_57484 (I65085,I3563,I980802,I980845,);
not I_57485 (I980853,I980845);
not I_57486 (I980870,I65103);
nor I_57487 (I980887,I980870,I65082);
not I_57488 (I980904,I65088);
nor I_57489 (I980921,I980887,I65094);
nor I_57490 (I980938,I980845,I980921);
DFFARX1 I_57491 (I980938,I3563,I980802,I980788,);
nor I_57492 (I980969,I65094,I65082);
nand I_57493 (I980986,I980969,I65103);
DFFARX1 I_57494 (I980986,I3563,I980802,I980791,);
nor I_57495 (I981017,I980904,I65094);
nand I_57496 (I981034,I981017,I65100);
nor I_57497 (I981051,I980828,I981034);
DFFARX1 I_57498 (I981051,I3563,I980802,I980767,);
not I_57499 (I981082,I981034);
nand I_57500 (I980779,I980845,I981082);
DFFARX1 I_57501 (I981034,I3563,I980802,I981122,);
not I_57502 (I981130,I981122);
not I_57503 (I981147,I65094);
not I_57504 (I981164,I65082);
nor I_57505 (I981181,I981164,I65088);
nor I_57506 (I980794,I981130,I981181);
nor I_57507 (I981212,I981164,I65091);
and I_57508 (I981229,I981212,I65079);
or I_57509 (I981246,I981229,I65097);
DFFARX1 I_57510 (I981246,I3563,I980802,I981272,);
nor I_57511 (I980782,I981272,I980828);
not I_57512 (I981294,I981272);
and I_57513 (I981311,I981294,I980828);
nor I_57514 (I980776,I980853,I981311);
nand I_57515 (I981342,I981294,I980904);
nor I_57516 (I980770,I981164,I981342);
nand I_57517 (I980773,I981294,I981082);
nand I_57518 (I981387,I980904,I65082);
nor I_57519 (I980785,I981147,I981387);
not I_57520 (I981448,I3570);
DFFARX1 I_57521 (I1100839,I3563,I981448,I981474,);
DFFARX1 I_57522 (I1100821,I3563,I981448,I981491,);
not I_57523 (I981499,I981491);
not I_57524 (I981516,I1100830);
nor I_57525 (I981533,I981516,I1100842);
not I_57526 (I981550,I1100824);
nor I_57527 (I981567,I981533,I1100833);
nor I_57528 (I981584,I981491,I981567);
DFFARX1 I_57529 (I981584,I3563,I981448,I981434,);
nor I_57530 (I981615,I1100833,I1100842);
nand I_57531 (I981632,I981615,I1100830);
DFFARX1 I_57532 (I981632,I3563,I981448,I981437,);
nor I_57533 (I981663,I981550,I1100833);
nand I_57534 (I981680,I981663,I1100845);
nor I_57535 (I981697,I981474,I981680);
DFFARX1 I_57536 (I981697,I3563,I981448,I981413,);
not I_57537 (I981728,I981680);
nand I_57538 (I981425,I981491,I981728);
DFFARX1 I_57539 (I981680,I3563,I981448,I981768,);
not I_57540 (I981776,I981768);
not I_57541 (I981793,I1100833);
not I_57542 (I981810,I1100821);
nor I_57543 (I981827,I981810,I1100824);
nor I_57544 (I981440,I981776,I981827);
nor I_57545 (I981858,I981810,I1100827);
and I_57546 (I981875,I981858,I1100836);
or I_57547 (I981892,I981875,I1100824);
DFFARX1 I_57548 (I981892,I3563,I981448,I981918,);
nor I_57549 (I981428,I981918,I981474);
not I_57550 (I981940,I981918);
and I_57551 (I981957,I981940,I981474);
nor I_57552 (I981422,I981499,I981957);
nand I_57553 (I981988,I981940,I981550);
nor I_57554 (I981416,I981810,I981988);
nand I_57555 (I981419,I981940,I981728);
nand I_57556 (I982033,I981550,I1100821);
nor I_57557 (I981431,I981793,I982033);
not I_57558 (I982094,I3570);
DFFARX1 I_57559 (I572719,I3563,I982094,I982120,);
DFFARX1 I_57560 (I572731,I3563,I982094,I982137,);
not I_57561 (I982145,I982137);
not I_57562 (I982162,I572716);
nor I_57563 (I982179,I982162,I572734);
not I_57564 (I982196,I572740);
nor I_57565 (I982213,I982179,I572722);
nor I_57566 (I982230,I982137,I982213);
DFFARX1 I_57567 (I982230,I3563,I982094,I982080,);
nor I_57568 (I982261,I572722,I572734);
nand I_57569 (I982278,I982261,I572716);
DFFARX1 I_57570 (I982278,I3563,I982094,I982083,);
nor I_57571 (I982309,I982196,I572722);
nand I_57572 (I982326,I982309,I572725);
nor I_57573 (I982343,I982120,I982326);
DFFARX1 I_57574 (I982343,I3563,I982094,I982059,);
not I_57575 (I982374,I982326);
nand I_57576 (I982071,I982137,I982374);
DFFARX1 I_57577 (I982326,I3563,I982094,I982414,);
not I_57578 (I982422,I982414);
not I_57579 (I982439,I572722);
not I_57580 (I982456,I572728);
nor I_57581 (I982473,I982456,I572740);
nor I_57582 (I982086,I982422,I982473);
nor I_57583 (I982504,I982456,I572737);
and I_57584 (I982521,I982504,I572716);
or I_57585 (I982538,I982521,I572719);
DFFARX1 I_57586 (I982538,I3563,I982094,I982564,);
nor I_57587 (I982074,I982564,I982120);
not I_57588 (I982586,I982564);
and I_57589 (I982603,I982586,I982120);
nor I_57590 (I982068,I982145,I982603);
nand I_57591 (I982634,I982586,I982196);
nor I_57592 (I982062,I982456,I982634);
nand I_57593 (I982065,I982586,I982374);
nand I_57594 (I982679,I982196,I572728);
nor I_57595 (I982077,I982439,I982679);
not I_57596 (I982740,I3570);
DFFARX1 I_57597 (I315404,I3563,I982740,I982766,);
DFFARX1 I_57598 (I315410,I3563,I982740,I982783,);
not I_57599 (I982791,I982783);
not I_57600 (I982808,I315431);
nor I_57601 (I982825,I982808,I315419);
not I_57602 (I982842,I315428);
nor I_57603 (I982859,I982825,I315413);
nor I_57604 (I982876,I982783,I982859);
DFFARX1 I_57605 (I982876,I3563,I982740,I982726,);
nor I_57606 (I982907,I315413,I315419);
nand I_57607 (I982924,I982907,I315431);
DFFARX1 I_57608 (I982924,I3563,I982740,I982729,);
nor I_57609 (I982955,I982842,I315413);
nand I_57610 (I982972,I982955,I315404);
nor I_57611 (I982989,I982766,I982972);
DFFARX1 I_57612 (I982989,I3563,I982740,I982705,);
not I_57613 (I983020,I982972);
nand I_57614 (I982717,I982783,I983020);
DFFARX1 I_57615 (I982972,I3563,I982740,I983060,);
not I_57616 (I983068,I983060);
not I_57617 (I983085,I315413);
not I_57618 (I983102,I315416);
nor I_57619 (I983119,I983102,I315428);
nor I_57620 (I982732,I983068,I983119);
nor I_57621 (I983150,I983102,I315425);
and I_57622 (I983167,I983150,I315407);
or I_57623 (I983184,I983167,I315422);
DFFARX1 I_57624 (I983184,I3563,I982740,I983210,);
nor I_57625 (I982720,I983210,I982766);
not I_57626 (I983232,I983210);
and I_57627 (I983249,I983232,I982766);
nor I_57628 (I982714,I982791,I983249);
nand I_57629 (I983280,I983232,I982842);
nor I_57630 (I982708,I983102,I983280);
nand I_57631 (I982711,I983232,I983020);
nand I_57632 (I983325,I982842,I315416);
nor I_57633 (I982723,I983085,I983325);
not I_57634 (I983386,I3570);
DFFARX1 I_57635 (I1620,I3563,I983386,I983412,);
DFFARX1 I_57636 (I2020,I3563,I983386,I983429,);
not I_57637 (I983437,I983429);
not I_57638 (I983454,I3284);
nor I_57639 (I983471,I983454,I2428);
not I_57640 (I983488,I3388);
nor I_57641 (I983505,I983471,I2060);
nor I_57642 (I983522,I983429,I983505);
DFFARX1 I_57643 (I983522,I3563,I983386,I983372,);
nor I_57644 (I983553,I2060,I2428);
nand I_57645 (I983570,I983553,I3284);
DFFARX1 I_57646 (I983570,I3563,I983386,I983375,);
nor I_57647 (I983601,I983488,I2060);
nand I_57648 (I983618,I983601,I1564);
nor I_57649 (I983635,I983412,I983618);
DFFARX1 I_57650 (I983635,I3563,I983386,I983351,);
not I_57651 (I983666,I983618);
nand I_57652 (I983363,I983429,I983666);
DFFARX1 I_57653 (I983618,I3563,I983386,I983706,);
not I_57654 (I983714,I983706);
not I_57655 (I983731,I2060);
not I_57656 (I983748,I1852);
nor I_57657 (I983765,I983748,I3388);
nor I_57658 (I983378,I983714,I983765);
nor I_57659 (I983796,I983748,I2276);
and I_57660 (I983813,I983796,I2268);
or I_57661 (I983830,I983813,I1980);
DFFARX1 I_57662 (I983830,I3563,I983386,I983856,);
nor I_57663 (I983366,I983856,I983412);
not I_57664 (I983878,I983856);
and I_57665 (I983895,I983878,I983412);
nor I_57666 (I983360,I983437,I983895);
nand I_57667 (I983926,I983878,I983488);
nor I_57668 (I983354,I983748,I983926);
nand I_57669 (I983357,I983878,I983666);
nand I_57670 (I983971,I983488,I1852);
nor I_57671 (I983369,I983731,I983971);
not I_57672 (I984032,I3570);
DFFARX1 I_57673 (I236309,I3563,I984032,I984058,);
DFFARX1 I_57674 (I236321,I3563,I984032,I984075,);
not I_57675 (I984083,I984075);
not I_57676 (I984100,I236327);
nor I_57677 (I984117,I984100,I236312);
not I_57678 (I984134,I236303);
nor I_57679 (I984151,I984117,I236324);
nor I_57680 (I984168,I984075,I984151);
DFFARX1 I_57681 (I984168,I3563,I984032,I984018,);
nor I_57682 (I984199,I236324,I236312);
nand I_57683 (I984216,I984199,I236327);
DFFARX1 I_57684 (I984216,I3563,I984032,I984021,);
nor I_57685 (I984247,I984134,I236324);
nand I_57686 (I984264,I984247,I236306);
nor I_57687 (I984281,I984058,I984264);
DFFARX1 I_57688 (I984281,I3563,I984032,I983997,);
not I_57689 (I984312,I984264);
nand I_57690 (I984009,I984075,I984312);
DFFARX1 I_57691 (I984264,I3563,I984032,I984352,);
not I_57692 (I984360,I984352);
not I_57693 (I984377,I236324);
not I_57694 (I984394,I236315);
nor I_57695 (I984411,I984394,I236303);
nor I_57696 (I984024,I984360,I984411);
nor I_57697 (I984442,I984394,I236318);
and I_57698 (I984459,I984442,I236306);
or I_57699 (I984476,I984459,I236303);
DFFARX1 I_57700 (I984476,I3563,I984032,I984502,);
nor I_57701 (I984012,I984502,I984058);
not I_57702 (I984524,I984502);
and I_57703 (I984541,I984524,I984058);
nor I_57704 (I984006,I984083,I984541);
nand I_57705 (I984572,I984524,I984134);
nor I_57706 (I984000,I984394,I984572);
nand I_57707 (I984003,I984524,I984312);
nand I_57708 (I984617,I984134,I236315);
nor I_57709 (I984015,I984377,I984617);
not I_57710 (I984678,I3570);
DFFARX1 I_57711 (I1244761,I3563,I984678,I984704,);
DFFARX1 I_57712 (I1244743,I3563,I984678,I984721,);
not I_57713 (I984729,I984721);
not I_57714 (I984746,I1244752);
nor I_57715 (I984763,I984746,I1244764);
not I_57716 (I984780,I1244746);
nor I_57717 (I984797,I984763,I1244755);
nor I_57718 (I984814,I984721,I984797);
DFFARX1 I_57719 (I984814,I3563,I984678,I984664,);
nor I_57720 (I984845,I1244755,I1244764);
nand I_57721 (I984862,I984845,I1244752);
DFFARX1 I_57722 (I984862,I3563,I984678,I984667,);
nor I_57723 (I984893,I984780,I1244755);
nand I_57724 (I984910,I984893,I1244767);
nor I_57725 (I984927,I984704,I984910);
DFFARX1 I_57726 (I984927,I3563,I984678,I984643,);
not I_57727 (I984958,I984910);
nand I_57728 (I984655,I984721,I984958);
DFFARX1 I_57729 (I984910,I3563,I984678,I984998,);
not I_57730 (I985006,I984998);
not I_57731 (I985023,I1244755);
not I_57732 (I985040,I1244743);
nor I_57733 (I985057,I985040,I1244746);
nor I_57734 (I984670,I985006,I985057);
nor I_57735 (I985088,I985040,I1244749);
and I_57736 (I985105,I985088,I1244758);
or I_57737 (I985122,I985105,I1244746);
DFFARX1 I_57738 (I985122,I3563,I984678,I985148,);
nor I_57739 (I984658,I985148,I984704);
not I_57740 (I985170,I985148);
and I_57741 (I985187,I985170,I984704);
nor I_57742 (I984652,I984729,I985187);
nand I_57743 (I985218,I985170,I984780);
nor I_57744 (I984646,I985040,I985218);
nand I_57745 (I984649,I985170,I984958);
nand I_57746 (I985263,I984780,I1244743);
nor I_57747 (I984661,I985023,I985263);
not I_57748 (I985324,I3570);
DFFARX1 I_57749 (I1385673,I3563,I985324,I985350,);
DFFARX1 I_57750 (I1385697,I3563,I985324,I985367,);
not I_57751 (I985375,I985367);
not I_57752 (I985392,I1385679);
nor I_57753 (I985409,I985392,I1385688);
not I_57754 (I985426,I1385673);
nor I_57755 (I985443,I985409,I1385694);
nor I_57756 (I985460,I985367,I985443);
DFFARX1 I_57757 (I985460,I3563,I985324,I985310,);
nor I_57758 (I985491,I1385694,I1385688);
nand I_57759 (I985508,I985491,I1385679);
DFFARX1 I_57760 (I985508,I3563,I985324,I985313,);
nor I_57761 (I985539,I985426,I1385694);
nand I_57762 (I985556,I985539,I1385691);
nor I_57763 (I985573,I985350,I985556);
DFFARX1 I_57764 (I985573,I3563,I985324,I985289,);
not I_57765 (I985604,I985556);
nand I_57766 (I985301,I985367,I985604);
DFFARX1 I_57767 (I985556,I3563,I985324,I985644,);
not I_57768 (I985652,I985644);
not I_57769 (I985669,I1385694);
not I_57770 (I985686,I1385685);
nor I_57771 (I985703,I985686,I1385673);
nor I_57772 (I985316,I985652,I985703);
nor I_57773 (I985734,I985686,I1385676);
and I_57774 (I985751,I985734,I1385700);
or I_57775 (I985768,I985751,I1385682);
DFFARX1 I_57776 (I985768,I3563,I985324,I985794,);
nor I_57777 (I985304,I985794,I985350);
not I_57778 (I985816,I985794);
and I_57779 (I985833,I985816,I985350);
nor I_57780 (I985298,I985375,I985833);
nand I_57781 (I985864,I985816,I985426);
nor I_57782 (I985292,I985686,I985864);
nand I_57783 (I985295,I985816,I985604);
nand I_57784 (I985909,I985426,I1385685);
nor I_57785 (I985307,I985669,I985909);
not I_57786 (I985970,I3570);
DFFARX1 I_57787 (I1398763,I3563,I985970,I985996,);
DFFARX1 I_57788 (I1398787,I3563,I985970,I986013,);
not I_57789 (I986021,I986013);
not I_57790 (I986038,I1398769);
nor I_57791 (I986055,I986038,I1398778);
not I_57792 (I986072,I1398763);
nor I_57793 (I986089,I986055,I1398784);
nor I_57794 (I986106,I986013,I986089);
DFFARX1 I_57795 (I986106,I3563,I985970,I985956,);
nor I_57796 (I986137,I1398784,I1398778);
nand I_57797 (I986154,I986137,I1398769);
DFFARX1 I_57798 (I986154,I3563,I985970,I985959,);
nor I_57799 (I986185,I986072,I1398784);
nand I_57800 (I986202,I986185,I1398781);
nor I_57801 (I986219,I985996,I986202);
DFFARX1 I_57802 (I986219,I3563,I985970,I985935,);
not I_57803 (I986250,I986202);
nand I_57804 (I985947,I986013,I986250);
DFFARX1 I_57805 (I986202,I3563,I985970,I986290,);
not I_57806 (I986298,I986290);
not I_57807 (I986315,I1398784);
not I_57808 (I986332,I1398775);
nor I_57809 (I986349,I986332,I1398763);
nor I_57810 (I985962,I986298,I986349);
nor I_57811 (I986380,I986332,I1398766);
and I_57812 (I986397,I986380,I1398790);
or I_57813 (I986414,I986397,I1398772);
DFFARX1 I_57814 (I986414,I3563,I985970,I986440,);
nor I_57815 (I985950,I986440,I985996);
not I_57816 (I986462,I986440);
and I_57817 (I986479,I986462,I985996);
nor I_57818 (I985944,I986021,I986479);
nand I_57819 (I986510,I986462,I986072);
nor I_57820 (I985938,I986332,I986510);
nand I_57821 (I985941,I986462,I986250);
nand I_57822 (I986555,I986072,I1398775);
nor I_57823 (I985953,I986315,I986555);
not I_57824 (I986616,I3570);
DFFARX1 I_57825 (I612176,I3563,I986616,I986642,);
DFFARX1 I_57826 (I612188,I3563,I986616,I986659,);
not I_57827 (I986667,I986659);
not I_57828 (I986684,I612197);
nor I_57829 (I986701,I986684,I612173);
not I_57830 (I986718,I612191);
nor I_57831 (I986735,I986701,I612185);
nor I_57832 (I986752,I986659,I986735);
DFFARX1 I_57833 (I986752,I3563,I986616,I986602,);
nor I_57834 (I986783,I612185,I612173);
nand I_57835 (I986800,I986783,I612197);
DFFARX1 I_57836 (I986800,I3563,I986616,I986605,);
nor I_57837 (I986831,I986718,I612185);
nand I_57838 (I986848,I986831,I612179);
nor I_57839 (I986865,I986642,I986848);
DFFARX1 I_57840 (I986865,I3563,I986616,I986581,);
not I_57841 (I986896,I986848);
nand I_57842 (I986593,I986659,I986896);
DFFARX1 I_57843 (I986848,I3563,I986616,I986936,);
not I_57844 (I986944,I986936);
not I_57845 (I986961,I612185);
not I_57846 (I986978,I612194);
nor I_57847 (I986995,I986978,I612191);
nor I_57848 (I986608,I986944,I986995);
nor I_57849 (I987026,I986978,I612176);
and I_57850 (I987043,I987026,I612173);
or I_57851 (I987060,I987043,I612182);
DFFARX1 I_57852 (I987060,I3563,I986616,I987086,);
nor I_57853 (I986596,I987086,I986642);
not I_57854 (I987108,I987086);
and I_57855 (I987125,I987108,I986642);
nor I_57856 (I986590,I986667,I987125);
nand I_57857 (I987156,I987108,I986718);
nor I_57858 (I986584,I986978,I987156);
nand I_57859 (I986587,I987108,I986896);
nand I_57860 (I987201,I986718,I612194);
nor I_57861 (I986599,I986961,I987201);
not I_57862 (I987262,I3570);
DFFARX1 I_57863 (I1403523,I3563,I987262,I987288,);
DFFARX1 I_57864 (I1403547,I3563,I987262,I987305,);
not I_57865 (I987313,I987305);
not I_57866 (I987330,I1403529);
nor I_57867 (I987347,I987330,I1403538);
not I_57868 (I987364,I1403523);
nor I_57869 (I987381,I987347,I1403544);
nor I_57870 (I987398,I987305,I987381);
DFFARX1 I_57871 (I987398,I3563,I987262,I987248,);
nor I_57872 (I987429,I1403544,I1403538);
nand I_57873 (I987446,I987429,I1403529);
DFFARX1 I_57874 (I987446,I3563,I987262,I987251,);
nor I_57875 (I987477,I987364,I1403544);
nand I_57876 (I987494,I987477,I1403541);
nor I_57877 (I987511,I987288,I987494);
DFFARX1 I_57878 (I987511,I3563,I987262,I987227,);
not I_57879 (I987542,I987494);
nand I_57880 (I987239,I987305,I987542);
DFFARX1 I_57881 (I987494,I3563,I987262,I987582,);
not I_57882 (I987590,I987582);
not I_57883 (I987607,I1403544);
not I_57884 (I987624,I1403535);
nor I_57885 (I987641,I987624,I1403523);
nor I_57886 (I987254,I987590,I987641);
nor I_57887 (I987672,I987624,I1403526);
and I_57888 (I987689,I987672,I1403550);
or I_57889 (I987706,I987689,I1403532);
DFFARX1 I_57890 (I987706,I3563,I987262,I987732,);
nor I_57891 (I987242,I987732,I987288);
not I_57892 (I987754,I987732);
and I_57893 (I987771,I987754,I987288);
nor I_57894 (I987236,I987313,I987771);
nand I_57895 (I987802,I987754,I987364);
nor I_57896 (I987230,I987624,I987802);
nand I_57897 (I987233,I987754,I987542);
nand I_57898 (I987847,I987364,I1403535);
nor I_57899 (I987245,I987607,I987847);
not I_57900 (I987908,I3570);
DFFARX1 I_57901 (I247614,I3563,I987908,I987934,);
DFFARX1 I_57902 (I247626,I3563,I987908,I987951,);
not I_57903 (I987959,I987951);
not I_57904 (I987976,I247632);
nor I_57905 (I987993,I987976,I247617);
not I_57906 (I988010,I247608);
nor I_57907 (I988027,I987993,I247629);
nor I_57908 (I988044,I987951,I988027);
DFFARX1 I_57909 (I988044,I3563,I987908,I987894,);
nor I_57910 (I988075,I247629,I247617);
nand I_57911 (I988092,I988075,I247632);
DFFARX1 I_57912 (I988092,I3563,I987908,I987897,);
nor I_57913 (I988123,I988010,I247629);
nand I_57914 (I988140,I988123,I247611);
nor I_57915 (I988157,I987934,I988140);
DFFARX1 I_57916 (I988157,I3563,I987908,I987873,);
not I_57917 (I988188,I988140);
nand I_57918 (I987885,I987951,I988188);
DFFARX1 I_57919 (I988140,I3563,I987908,I988228,);
not I_57920 (I988236,I988228);
not I_57921 (I988253,I247629);
not I_57922 (I988270,I247620);
nor I_57923 (I988287,I988270,I247608);
nor I_57924 (I987900,I988236,I988287);
nor I_57925 (I988318,I988270,I247623);
and I_57926 (I988335,I988318,I247611);
or I_57927 (I988352,I988335,I247608);
DFFARX1 I_57928 (I988352,I3563,I987908,I988378,);
nor I_57929 (I987888,I988378,I987934);
not I_57930 (I988400,I988378);
and I_57931 (I988417,I988400,I987934);
nor I_57932 (I987882,I987959,I988417);
nand I_57933 (I988448,I988400,I988010);
nor I_57934 (I987876,I988270,I988448);
nand I_57935 (I987879,I988400,I988188);
nand I_57936 (I988493,I988010,I247620);
nor I_57937 (I987891,I988253,I988493);
not I_57938 (I988554,I3570);
DFFARX1 I_57939 (I1083685,I3563,I988554,I988580,);
DFFARX1 I_57940 (I1083688,I3563,I988554,I988597,);
not I_57941 (I988605,I988597);
not I_57942 (I988622,I1083685);
nor I_57943 (I988639,I988622,I1083697);
not I_57944 (I988656,I1083706);
nor I_57945 (I988673,I988639,I1083694);
nor I_57946 (I988690,I988597,I988673);
DFFARX1 I_57947 (I988690,I3563,I988554,I988540,);
nor I_57948 (I988721,I1083694,I1083697);
nand I_57949 (I988738,I988721,I1083685);
DFFARX1 I_57950 (I988738,I3563,I988554,I988543,);
nor I_57951 (I988769,I988656,I1083694);
nand I_57952 (I988786,I988769,I1083700);
nor I_57953 (I988803,I988580,I988786);
DFFARX1 I_57954 (I988803,I3563,I988554,I988519,);
not I_57955 (I988834,I988786);
nand I_57956 (I988531,I988597,I988834);
DFFARX1 I_57957 (I988786,I3563,I988554,I988874,);
not I_57958 (I988882,I988874);
not I_57959 (I988899,I1083694);
not I_57960 (I988916,I1083691);
nor I_57961 (I988933,I988916,I1083706);
nor I_57962 (I988546,I988882,I988933);
nor I_57963 (I988964,I988916,I1083703);
and I_57964 (I988981,I988964,I1083691);
or I_57965 (I988998,I988981,I1083688);
DFFARX1 I_57966 (I988998,I3563,I988554,I989024,);
nor I_57967 (I988534,I989024,I988580);
not I_57968 (I989046,I989024);
and I_57969 (I989063,I989046,I988580);
nor I_57970 (I988528,I988605,I989063);
nand I_57971 (I989094,I989046,I988656);
nor I_57972 (I988522,I988916,I989094);
nand I_57973 (I988525,I989046,I988834);
nand I_57974 (I989139,I988656,I1083691);
nor I_57975 (I988537,I988899,I989139);
not I_57976 (I989200,I3570);
DFFARX1 I_57977 (I622002,I3563,I989200,I989226,);
DFFARX1 I_57978 (I622014,I3563,I989200,I989243,);
not I_57979 (I989251,I989243);
not I_57980 (I989268,I622023);
nor I_57981 (I989285,I989268,I621999);
not I_57982 (I989302,I622017);
nor I_57983 (I989319,I989285,I622011);
nor I_57984 (I989336,I989243,I989319);
DFFARX1 I_57985 (I989336,I3563,I989200,I989186,);
nor I_57986 (I989367,I622011,I621999);
nand I_57987 (I989384,I989367,I622023);
DFFARX1 I_57988 (I989384,I3563,I989200,I989189,);
nor I_57989 (I989415,I989302,I622011);
nand I_57990 (I989432,I989415,I622005);
nor I_57991 (I989449,I989226,I989432);
DFFARX1 I_57992 (I989449,I3563,I989200,I989165,);
not I_57993 (I989480,I989432);
nand I_57994 (I989177,I989243,I989480);
DFFARX1 I_57995 (I989432,I3563,I989200,I989520,);
not I_57996 (I989528,I989520);
not I_57997 (I989545,I622011);
not I_57998 (I989562,I622020);
nor I_57999 (I989579,I989562,I622017);
nor I_58000 (I989192,I989528,I989579);
nor I_58001 (I989610,I989562,I622002);
and I_58002 (I989627,I989610,I621999);
or I_58003 (I989644,I989627,I622008);
DFFARX1 I_58004 (I989644,I3563,I989200,I989670,);
nor I_58005 (I989180,I989670,I989226);
not I_58006 (I989692,I989670);
and I_58007 (I989709,I989692,I989226);
nor I_58008 (I989174,I989251,I989709);
nand I_58009 (I989740,I989692,I989302);
nor I_58010 (I989168,I989562,I989740);
nand I_58011 (I989171,I989692,I989480);
nand I_58012 (I989785,I989302,I622020);
nor I_58013 (I989183,I989545,I989785);
not I_58014 (I989846,I3570);
DFFARX1 I_58015 (I894328,I3563,I989846,I989872,);
DFFARX1 I_58016 (I894325,I3563,I989846,I989889,);
not I_58017 (I989897,I989889);
not I_58018 (I989914,I894325);
nor I_58019 (I989931,I989914,I894328);
not I_58020 (I989948,I894340);
nor I_58021 (I989965,I989931,I894334);
nor I_58022 (I989982,I989889,I989965);
DFFARX1 I_58023 (I989982,I3563,I989846,I989832,);
nor I_58024 (I990013,I894334,I894328);
nand I_58025 (I990030,I990013,I894325);
DFFARX1 I_58026 (I990030,I3563,I989846,I989835,);
nor I_58027 (I990061,I989948,I894334);
nand I_58028 (I990078,I990061,I894322);
nor I_58029 (I990095,I989872,I990078);
DFFARX1 I_58030 (I990095,I3563,I989846,I989811,);
not I_58031 (I990126,I990078);
nand I_58032 (I989823,I989889,I990126);
DFFARX1 I_58033 (I990078,I3563,I989846,I990166,);
not I_58034 (I990174,I990166);
not I_58035 (I990191,I894334);
not I_58036 (I990208,I894331);
nor I_58037 (I990225,I990208,I894340);
nor I_58038 (I989838,I990174,I990225);
nor I_58039 (I990256,I990208,I894337);
and I_58040 (I990273,I990256,I894343);
or I_58041 (I990290,I990273,I894322);
DFFARX1 I_58042 (I990290,I3563,I989846,I990316,);
nor I_58043 (I989826,I990316,I989872);
not I_58044 (I990338,I990316);
and I_58045 (I990355,I990338,I989872);
nor I_58046 (I989820,I989897,I990355);
nand I_58047 (I990386,I990338,I989948);
nor I_58048 (I989814,I990208,I990386);
nand I_58049 (I989817,I990338,I990126);
nand I_58050 (I990431,I989948,I894331);
nor I_58051 (I989829,I990191,I990431);
not I_58052 (I990492,I3570);
DFFARX1 I_58053 (I489864,I3563,I990492,I990518,);
DFFARX1 I_58054 (I489861,I3563,I990492,I990535,);
not I_58055 (I990543,I990535);
not I_58056 (I990560,I489876);
nor I_58057 (I990577,I990560,I489879);
not I_58058 (I990594,I489867);
nor I_58059 (I990611,I990577,I489873);
nor I_58060 (I990628,I990535,I990611);
DFFARX1 I_58061 (I990628,I3563,I990492,I990478,);
nor I_58062 (I990659,I489873,I489879);
nand I_58063 (I990676,I990659,I489876);
DFFARX1 I_58064 (I990676,I3563,I990492,I990481,);
nor I_58065 (I990707,I990594,I489873);
nand I_58066 (I990724,I990707,I489885);
nor I_58067 (I990741,I990518,I990724);
DFFARX1 I_58068 (I990741,I3563,I990492,I990457,);
not I_58069 (I990772,I990724);
nand I_58070 (I990469,I990535,I990772);
DFFARX1 I_58071 (I990724,I3563,I990492,I990812,);
not I_58072 (I990820,I990812);
not I_58073 (I990837,I489873);
not I_58074 (I990854,I489858);
nor I_58075 (I990871,I990854,I489867);
nor I_58076 (I990484,I990820,I990871);
nor I_58077 (I990902,I990854,I489870);
and I_58078 (I990919,I990902,I489858);
or I_58079 (I990936,I990919,I489882);
DFFARX1 I_58080 (I990936,I3563,I990492,I990962,);
nor I_58081 (I990472,I990962,I990518);
not I_58082 (I990984,I990962);
and I_58083 (I991001,I990984,I990518);
nor I_58084 (I990466,I990543,I991001);
nand I_58085 (I991032,I990984,I990594);
nor I_58086 (I990460,I990854,I991032);
nand I_58087 (I990463,I990984,I990772);
nand I_58088 (I991077,I990594,I489858);
nor I_58089 (I990475,I990837,I991077);
not I_58090 (I991138,I3570);
DFFARX1 I_58091 (I1115867,I3563,I991138,I991164,);
DFFARX1 I_58092 (I1115849,I3563,I991138,I991181,);
not I_58093 (I991189,I991181);
not I_58094 (I991206,I1115858);
nor I_58095 (I991223,I991206,I1115870);
not I_58096 (I991240,I1115852);
nor I_58097 (I991257,I991223,I1115861);
nor I_58098 (I991274,I991181,I991257);
DFFARX1 I_58099 (I991274,I3563,I991138,I991124,);
nor I_58100 (I991305,I1115861,I1115870);
nand I_58101 (I991322,I991305,I1115858);
DFFARX1 I_58102 (I991322,I3563,I991138,I991127,);
nor I_58103 (I991353,I991240,I1115861);
nand I_58104 (I991370,I991353,I1115873);
nor I_58105 (I991387,I991164,I991370);
DFFARX1 I_58106 (I991387,I3563,I991138,I991103,);
not I_58107 (I991418,I991370);
nand I_58108 (I991115,I991181,I991418);
DFFARX1 I_58109 (I991370,I3563,I991138,I991458,);
not I_58110 (I991466,I991458);
not I_58111 (I991483,I1115861);
not I_58112 (I991500,I1115849);
nor I_58113 (I991517,I991500,I1115852);
nor I_58114 (I991130,I991466,I991517);
nor I_58115 (I991548,I991500,I1115855);
and I_58116 (I991565,I991548,I1115864);
or I_58117 (I991582,I991565,I1115852);
DFFARX1 I_58118 (I991582,I3563,I991138,I991608,);
nor I_58119 (I991118,I991608,I991164);
not I_58120 (I991630,I991608);
and I_58121 (I991647,I991630,I991164);
nor I_58122 (I991112,I991189,I991647);
nand I_58123 (I991678,I991630,I991240);
nor I_58124 (I991106,I991500,I991678);
nand I_58125 (I991109,I991630,I991418);
nand I_58126 (I991723,I991240,I1115849);
nor I_58127 (I991121,I991483,I991723);
not I_58128 (I991784,I3570);
DFFARX1 I_58129 (I459944,I3563,I991784,I991810,);
DFFARX1 I_58130 (I459941,I3563,I991784,I991827,);
not I_58131 (I991835,I991827);
not I_58132 (I991852,I459956);
nor I_58133 (I991869,I991852,I459959);
not I_58134 (I991886,I459947);
nor I_58135 (I991903,I991869,I459953);
nor I_58136 (I991920,I991827,I991903);
DFFARX1 I_58137 (I991920,I3563,I991784,I991770,);
nor I_58138 (I991951,I459953,I459959);
nand I_58139 (I991968,I991951,I459956);
DFFARX1 I_58140 (I991968,I3563,I991784,I991773,);
nor I_58141 (I991999,I991886,I459953);
nand I_58142 (I992016,I991999,I459965);
nor I_58143 (I992033,I991810,I992016);
DFFARX1 I_58144 (I992033,I3563,I991784,I991749,);
not I_58145 (I992064,I992016);
nand I_58146 (I991761,I991827,I992064);
DFFARX1 I_58147 (I992016,I3563,I991784,I992104,);
not I_58148 (I992112,I992104);
not I_58149 (I992129,I459953);
not I_58150 (I992146,I459938);
nor I_58151 (I992163,I992146,I459947);
nor I_58152 (I991776,I992112,I992163);
nor I_58153 (I992194,I992146,I459950);
and I_58154 (I992211,I992194,I459938);
or I_58155 (I992228,I992211,I459962);
DFFARX1 I_58156 (I992228,I3563,I991784,I992254,);
nor I_58157 (I991764,I992254,I991810);
not I_58158 (I992276,I992254);
and I_58159 (I992293,I992276,I991810);
nor I_58160 (I991758,I991835,I992293);
nand I_58161 (I992324,I992276,I991886);
nor I_58162 (I991752,I992146,I992324);
nand I_58163 (I991755,I992276,I992064);
nand I_58164 (I992369,I991886,I459938);
nor I_58165 (I991767,I992129,I992369);
not I_58166 (I992430,I3570);
DFFARX1 I_58167 (I449608,I3563,I992430,I992456,);
DFFARX1 I_58168 (I449605,I3563,I992430,I992473,);
not I_58169 (I992481,I992473);
not I_58170 (I992498,I449620);
nor I_58171 (I992515,I992498,I449623);
not I_58172 (I992532,I449611);
nor I_58173 (I992549,I992515,I449617);
nor I_58174 (I992566,I992473,I992549);
DFFARX1 I_58175 (I992566,I3563,I992430,I992416,);
nor I_58176 (I992597,I449617,I449623);
nand I_58177 (I992614,I992597,I449620);
DFFARX1 I_58178 (I992614,I3563,I992430,I992419,);
nor I_58179 (I992645,I992532,I449617);
nand I_58180 (I992662,I992645,I449629);
nor I_58181 (I992679,I992456,I992662);
DFFARX1 I_58182 (I992679,I3563,I992430,I992395,);
not I_58183 (I992710,I992662);
nand I_58184 (I992407,I992473,I992710);
DFFARX1 I_58185 (I992662,I3563,I992430,I992750,);
not I_58186 (I992758,I992750);
not I_58187 (I992775,I449617);
not I_58188 (I992792,I449602);
nor I_58189 (I992809,I992792,I449611);
nor I_58190 (I992422,I992758,I992809);
nor I_58191 (I992840,I992792,I449614);
and I_58192 (I992857,I992840,I449602);
or I_58193 (I992874,I992857,I449626);
DFFARX1 I_58194 (I992874,I3563,I992430,I992900,);
nor I_58195 (I992410,I992900,I992456);
not I_58196 (I992922,I992900);
and I_58197 (I992939,I992922,I992456);
nor I_58198 (I992404,I992481,I992939);
nand I_58199 (I992970,I992922,I992532);
nor I_58200 (I992398,I992792,I992970);
nand I_58201 (I992401,I992922,I992710);
nand I_58202 (I993015,I992532,I449602);
nor I_58203 (I992413,I992775,I993015);
not I_58204 (I993076,I3570);
DFFARX1 I_58205 (I249994,I3563,I993076,I993102,);
DFFARX1 I_58206 (I250006,I3563,I993076,I993119,);
not I_58207 (I993127,I993119);
not I_58208 (I993144,I250012);
nor I_58209 (I993161,I993144,I249997);
not I_58210 (I993178,I249988);
nor I_58211 (I993195,I993161,I250009);
nor I_58212 (I993212,I993119,I993195);
DFFARX1 I_58213 (I993212,I3563,I993076,I993062,);
nor I_58214 (I993243,I250009,I249997);
nand I_58215 (I993260,I993243,I250012);
DFFARX1 I_58216 (I993260,I3563,I993076,I993065,);
nor I_58217 (I993291,I993178,I250009);
nand I_58218 (I993308,I993291,I249991);
nor I_58219 (I993325,I993102,I993308);
DFFARX1 I_58220 (I993325,I3563,I993076,I993041,);
not I_58221 (I993356,I993308);
nand I_58222 (I993053,I993119,I993356);
DFFARX1 I_58223 (I993308,I3563,I993076,I993396,);
not I_58224 (I993404,I993396);
not I_58225 (I993421,I250009);
not I_58226 (I993438,I250000);
nor I_58227 (I993455,I993438,I249988);
nor I_58228 (I993068,I993404,I993455);
nor I_58229 (I993486,I993438,I250003);
and I_58230 (I993503,I993486,I249991);
or I_58231 (I993520,I993503,I249988);
DFFARX1 I_58232 (I993520,I3563,I993076,I993546,);
nor I_58233 (I993056,I993546,I993102);
not I_58234 (I993568,I993546);
and I_58235 (I993585,I993568,I993102);
nor I_58236 (I993050,I993127,I993585);
nand I_58237 (I993616,I993568,I993178);
nor I_58238 (I993044,I993438,I993616);
nand I_58239 (I993047,I993568,I993356);
nand I_58240 (I993661,I993178,I250000);
nor I_58241 (I993059,I993421,I993661);
not I_58242 (I993722,I3570);
DFFARX1 I_58243 (I123049,I3563,I993722,I993748,);
DFFARX1 I_58244 (I123055,I3563,I993722,I993765,);
not I_58245 (I993773,I993765);
not I_58246 (I993790,I123073);
nor I_58247 (I993807,I993790,I123052);
not I_58248 (I993824,I123058);
nor I_58249 (I993841,I993807,I123064);
nor I_58250 (I993858,I993765,I993841);
DFFARX1 I_58251 (I993858,I3563,I993722,I993708,);
nor I_58252 (I993889,I123064,I123052);
nand I_58253 (I993906,I993889,I123073);
DFFARX1 I_58254 (I993906,I3563,I993722,I993711,);
nor I_58255 (I993937,I993824,I123064);
nand I_58256 (I993954,I993937,I123070);
nor I_58257 (I993971,I993748,I993954);
DFFARX1 I_58258 (I993971,I3563,I993722,I993687,);
not I_58259 (I994002,I993954);
nand I_58260 (I993699,I993765,I994002);
DFFARX1 I_58261 (I993954,I3563,I993722,I994042,);
not I_58262 (I994050,I994042);
not I_58263 (I994067,I123064);
not I_58264 (I994084,I123052);
nor I_58265 (I994101,I994084,I123058);
nor I_58266 (I993714,I994050,I994101);
nor I_58267 (I994132,I994084,I123061);
and I_58268 (I994149,I994132,I123049);
or I_58269 (I994166,I994149,I123067);
DFFARX1 I_58270 (I994166,I3563,I993722,I994192,);
nor I_58271 (I993702,I994192,I993748);
not I_58272 (I994214,I994192);
and I_58273 (I994231,I994214,I993748);
nor I_58274 (I993696,I993773,I994231);
nand I_58275 (I994262,I994214,I993824);
nor I_58276 (I993690,I994084,I994262);
nand I_58277 (I993693,I994214,I994002);
nand I_58278 (I994307,I993824,I123052);
nor I_58279 (I993705,I994067,I994307);
not I_58280 (I994368,I3570);
DFFARX1 I_58281 (I1114711,I3563,I994368,I994394,);
DFFARX1 I_58282 (I1114693,I3563,I994368,I994411,);
not I_58283 (I994419,I994411);
not I_58284 (I994436,I1114702);
nor I_58285 (I994453,I994436,I1114714);
not I_58286 (I994470,I1114696);
nor I_58287 (I994487,I994453,I1114705);
nor I_58288 (I994504,I994411,I994487);
DFFARX1 I_58289 (I994504,I3563,I994368,I994354,);
nor I_58290 (I994535,I1114705,I1114714);
nand I_58291 (I994552,I994535,I1114702);
DFFARX1 I_58292 (I994552,I3563,I994368,I994357,);
nor I_58293 (I994583,I994470,I1114705);
nand I_58294 (I994600,I994583,I1114717);
nor I_58295 (I994617,I994394,I994600);
DFFARX1 I_58296 (I994617,I3563,I994368,I994333,);
not I_58297 (I994648,I994600);
nand I_58298 (I994345,I994411,I994648);
DFFARX1 I_58299 (I994600,I3563,I994368,I994688,);
not I_58300 (I994696,I994688);
not I_58301 (I994713,I1114705);
not I_58302 (I994730,I1114693);
nor I_58303 (I994747,I994730,I1114696);
nor I_58304 (I994360,I994696,I994747);
nor I_58305 (I994778,I994730,I1114699);
and I_58306 (I994795,I994778,I1114708);
or I_58307 (I994812,I994795,I1114696);
DFFARX1 I_58308 (I994812,I3563,I994368,I994838,);
nor I_58309 (I994348,I994838,I994394);
not I_58310 (I994860,I994838);
and I_58311 (I994877,I994860,I994394);
nor I_58312 (I994342,I994419,I994877);
nand I_58313 (I994908,I994860,I994470);
nor I_58314 (I994336,I994730,I994908);
nand I_58315 (I994339,I994860,I994648);
nand I_58316 (I994953,I994470,I1114693);
nor I_58317 (I994351,I994713,I994953);
not I_58318 (I995014,I3570);
DFFARX1 I_58319 (I456136,I3563,I995014,I995040,);
DFFARX1 I_58320 (I456133,I3563,I995014,I995057,);
not I_58321 (I995065,I995057);
not I_58322 (I995082,I456148);
nor I_58323 (I995099,I995082,I456151);
not I_58324 (I995116,I456139);
nor I_58325 (I995133,I995099,I456145);
nor I_58326 (I995150,I995057,I995133);
DFFARX1 I_58327 (I995150,I3563,I995014,I995000,);
nor I_58328 (I995181,I456145,I456151);
nand I_58329 (I995198,I995181,I456148);
DFFARX1 I_58330 (I995198,I3563,I995014,I995003,);
nor I_58331 (I995229,I995116,I456145);
nand I_58332 (I995246,I995229,I456157);
nor I_58333 (I995263,I995040,I995246);
DFFARX1 I_58334 (I995263,I3563,I995014,I994979,);
not I_58335 (I995294,I995246);
nand I_58336 (I994991,I995057,I995294);
DFFARX1 I_58337 (I995246,I3563,I995014,I995334,);
not I_58338 (I995342,I995334);
not I_58339 (I995359,I456145);
not I_58340 (I995376,I456130);
nor I_58341 (I995393,I995376,I456139);
nor I_58342 (I995006,I995342,I995393);
nor I_58343 (I995424,I995376,I456142);
and I_58344 (I995441,I995424,I456130);
or I_58345 (I995458,I995441,I456154);
DFFARX1 I_58346 (I995458,I3563,I995014,I995484,);
nor I_58347 (I994994,I995484,I995040);
not I_58348 (I995506,I995484);
and I_58349 (I995523,I995506,I995040);
nor I_58350 (I994988,I995065,I995523);
nand I_58351 (I995554,I995506,I995116);
nor I_58352 (I994982,I995376,I995554);
nand I_58353 (I994985,I995506,I995294);
nand I_58354 (I995599,I995116,I456130);
nor I_58355 (I994997,I995359,I995599);
not I_58356 (I995660,I3570);
DFFARX1 I_58357 (I433832,I3563,I995660,I995686,);
DFFARX1 I_58358 (I433829,I3563,I995660,I995703,);
not I_58359 (I995711,I995703);
not I_58360 (I995728,I433844);
nor I_58361 (I995745,I995728,I433847);
not I_58362 (I995762,I433835);
nor I_58363 (I995779,I995745,I433841);
nor I_58364 (I995796,I995703,I995779);
DFFARX1 I_58365 (I995796,I3563,I995660,I995646,);
nor I_58366 (I995827,I433841,I433847);
nand I_58367 (I995844,I995827,I433844);
DFFARX1 I_58368 (I995844,I3563,I995660,I995649,);
nor I_58369 (I995875,I995762,I433841);
nand I_58370 (I995892,I995875,I433853);
nor I_58371 (I995909,I995686,I995892);
DFFARX1 I_58372 (I995909,I3563,I995660,I995625,);
not I_58373 (I995940,I995892);
nand I_58374 (I995637,I995703,I995940);
DFFARX1 I_58375 (I995892,I3563,I995660,I995980,);
not I_58376 (I995988,I995980);
not I_58377 (I996005,I433841);
not I_58378 (I996022,I433826);
nor I_58379 (I996039,I996022,I433835);
nor I_58380 (I995652,I995988,I996039);
nor I_58381 (I996070,I996022,I433838);
and I_58382 (I996087,I996070,I433826);
or I_58383 (I996104,I996087,I433850);
DFFARX1 I_58384 (I996104,I3563,I995660,I996130,);
nor I_58385 (I995640,I996130,I995686);
not I_58386 (I996152,I996130);
and I_58387 (I996169,I996152,I995686);
nor I_58388 (I995634,I995711,I996169);
nand I_58389 (I996200,I996152,I995762);
nor I_58390 (I995628,I996022,I996200);
nand I_58391 (I995631,I996152,I995940);
nand I_58392 (I996245,I995762,I433826);
nor I_58393 (I995643,I996005,I996245);
not I_58394 (I996306,I3570);
DFFARX1 I_58395 (I777487,I3563,I996306,I996332,);
DFFARX1 I_58396 (I777481,I3563,I996306,I996349,);
not I_58397 (I996357,I996349);
not I_58398 (I996374,I777496);
nor I_58399 (I996391,I996374,I777481);
not I_58400 (I996408,I777490);
nor I_58401 (I996425,I996391,I777499);
nor I_58402 (I996442,I996349,I996425);
DFFARX1 I_58403 (I996442,I3563,I996306,I996292,);
nor I_58404 (I996473,I777499,I777481);
nand I_58405 (I996490,I996473,I777496);
DFFARX1 I_58406 (I996490,I3563,I996306,I996295,);
nor I_58407 (I996521,I996408,I777499);
nand I_58408 (I996538,I996521,I777484);
nor I_58409 (I996555,I996332,I996538);
DFFARX1 I_58410 (I996555,I3563,I996306,I996271,);
not I_58411 (I996586,I996538);
nand I_58412 (I996283,I996349,I996586);
DFFARX1 I_58413 (I996538,I3563,I996306,I996626,);
not I_58414 (I996634,I996626);
not I_58415 (I996651,I777499);
not I_58416 (I996668,I777493);
nor I_58417 (I996685,I996668,I777490);
nor I_58418 (I996298,I996634,I996685);
nor I_58419 (I996716,I996668,I777502);
and I_58420 (I996733,I996716,I777505);
or I_58421 (I996750,I996733,I777484);
DFFARX1 I_58422 (I996750,I3563,I996306,I996776,);
nor I_58423 (I996286,I996776,I996332);
not I_58424 (I996798,I996776);
and I_58425 (I996815,I996798,I996332);
nor I_58426 (I996280,I996357,I996815);
nand I_58427 (I996846,I996798,I996408);
nor I_58428 (I996274,I996668,I996846);
nand I_58429 (I996277,I996798,I996586);
nand I_58430 (I996891,I996408,I777493);
nor I_58431 (I996289,I996651,I996891);
not I_58432 (I996952,I3570);
DFFARX1 I_58433 (I521960,I3563,I996952,I996978,);
DFFARX1 I_58434 (I521957,I3563,I996952,I996995,);
not I_58435 (I997003,I996995);
not I_58436 (I997020,I521972);
nor I_58437 (I997037,I997020,I521975);
not I_58438 (I997054,I521963);
nor I_58439 (I997071,I997037,I521969);
nor I_58440 (I997088,I996995,I997071);
DFFARX1 I_58441 (I997088,I3563,I996952,I996938,);
nor I_58442 (I997119,I521969,I521975);
nand I_58443 (I997136,I997119,I521972);
DFFARX1 I_58444 (I997136,I3563,I996952,I996941,);
nor I_58445 (I997167,I997054,I521969);
nand I_58446 (I997184,I997167,I521981);
nor I_58447 (I997201,I996978,I997184);
DFFARX1 I_58448 (I997201,I3563,I996952,I996917,);
not I_58449 (I997232,I997184);
nand I_58450 (I996929,I996995,I997232);
DFFARX1 I_58451 (I997184,I3563,I996952,I997272,);
not I_58452 (I997280,I997272);
not I_58453 (I997297,I521969);
not I_58454 (I997314,I521954);
nor I_58455 (I997331,I997314,I521963);
nor I_58456 (I996944,I997280,I997331);
nor I_58457 (I997362,I997314,I521966);
and I_58458 (I997379,I997362,I521954);
or I_58459 (I997396,I997379,I521978);
DFFARX1 I_58460 (I997396,I3563,I996952,I997422,);
nor I_58461 (I996932,I997422,I996978);
not I_58462 (I997444,I997422);
and I_58463 (I997461,I997444,I996978);
nor I_58464 (I996926,I997003,I997461);
nand I_58465 (I997492,I997444,I997054);
nor I_58466 (I996920,I997314,I997492);
nand I_58467 (I996923,I997444,I997232);
nand I_58468 (I997537,I997054,I521954);
nor I_58469 (I996935,I997297,I997537);
not I_58470 (I997598,I3570);
DFFARX1 I_58471 (I439272,I3563,I997598,I997624,);
DFFARX1 I_58472 (I439269,I3563,I997598,I997641,);
not I_58473 (I997649,I997641);
not I_58474 (I997666,I439284);
nor I_58475 (I997683,I997666,I439287);
not I_58476 (I997700,I439275);
nor I_58477 (I997717,I997683,I439281);
nor I_58478 (I997734,I997641,I997717);
DFFARX1 I_58479 (I997734,I3563,I997598,I997584,);
nor I_58480 (I997765,I439281,I439287);
nand I_58481 (I997782,I997765,I439284);
DFFARX1 I_58482 (I997782,I3563,I997598,I997587,);
nor I_58483 (I997813,I997700,I439281);
nand I_58484 (I997830,I997813,I439293);
nor I_58485 (I997847,I997624,I997830);
DFFARX1 I_58486 (I997847,I3563,I997598,I997563,);
not I_58487 (I997878,I997830);
nand I_58488 (I997575,I997641,I997878);
DFFARX1 I_58489 (I997830,I3563,I997598,I997918,);
not I_58490 (I997926,I997918);
not I_58491 (I997943,I439281);
not I_58492 (I997960,I439266);
nor I_58493 (I997977,I997960,I439275);
nor I_58494 (I997590,I997926,I997977);
nor I_58495 (I998008,I997960,I439278);
and I_58496 (I998025,I998008,I439266);
or I_58497 (I998042,I998025,I439290);
DFFARX1 I_58498 (I998042,I3563,I997598,I998068,);
nor I_58499 (I997578,I998068,I997624);
not I_58500 (I998090,I998068);
and I_58501 (I998107,I998090,I997624);
nor I_58502 (I997572,I997649,I998107);
nand I_58503 (I998138,I998090,I997700);
nor I_58504 (I997566,I997960,I998138);
nand I_58505 (I997569,I998090,I997878);
nand I_58506 (I998183,I997700,I439266);
nor I_58507 (I997581,I997943,I998183);
not I_58508 (I998244,I3570);
DFFARX1 I_58509 (I617956,I3563,I998244,I998270,);
DFFARX1 I_58510 (I617968,I3563,I998244,I998287,);
not I_58511 (I998295,I998287);
not I_58512 (I998312,I617977);
nor I_58513 (I998329,I998312,I617953);
not I_58514 (I998346,I617971);
nor I_58515 (I998363,I998329,I617965);
nor I_58516 (I998380,I998287,I998363);
DFFARX1 I_58517 (I998380,I3563,I998244,I998230,);
nor I_58518 (I998411,I617965,I617953);
nand I_58519 (I998428,I998411,I617977);
DFFARX1 I_58520 (I998428,I3563,I998244,I998233,);
nor I_58521 (I998459,I998346,I617965);
nand I_58522 (I998476,I998459,I617959);
nor I_58523 (I998493,I998270,I998476);
DFFARX1 I_58524 (I998493,I3563,I998244,I998209,);
not I_58525 (I998524,I998476);
nand I_58526 (I998221,I998287,I998524);
DFFARX1 I_58527 (I998476,I3563,I998244,I998564,);
not I_58528 (I998572,I998564);
not I_58529 (I998589,I617965);
not I_58530 (I998606,I617974);
nor I_58531 (I998623,I998606,I617971);
nor I_58532 (I998236,I998572,I998623);
nor I_58533 (I998654,I998606,I617956);
and I_58534 (I998671,I998654,I617953);
or I_58535 (I998688,I998671,I617962);
DFFARX1 I_58536 (I998688,I3563,I998244,I998714,);
nor I_58537 (I998224,I998714,I998270);
not I_58538 (I998736,I998714);
and I_58539 (I998753,I998736,I998270);
nor I_58540 (I998218,I998295,I998753);
nand I_58541 (I998784,I998736,I998346);
nor I_58542 (I998212,I998606,I998784);
nand I_58543 (I998215,I998736,I998524);
nand I_58544 (I998829,I998346,I617974);
nor I_58545 (I998227,I998589,I998829);
not I_58546 (I998890,I3570);
DFFARX1 I_58547 (I425128,I3563,I998890,I998916,);
DFFARX1 I_58548 (I425125,I3563,I998890,I998933,);
not I_58549 (I998941,I998933);
not I_58550 (I998958,I425140);
nor I_58551 (I998975,I998958,I425143);
not I_58552 (I998992,I425131);
nor I_58553 (I999009,I998975,I425137);
nor I_58554 (I999026,I998933,I999009);
DFFARX1 I_58555 (I999026,I3563,I998890,I998876,);
nor I_58556 (I999057,I425137,I425143);
nand I_58557 (I999074,I999057,I425140);
DFFARX1 I_58558 (I999074,I3563,I998890,I998879,);
nor I_58559 (I999105,I998992,I425137);
nand I_58560 (I999122,I999105,I425149);
nor I_58561 (I999139,I998916,I999122);
DFFARX1 I_58562 (I999139,I3563,I998890,I998855,);
not I_58563 (I999170,I999122);
nand I_58564 (I998867,I998933,I999170);
DFFARX1 I_58565 (I999122,I3563,I998890,I999210,);
not I_58566 (I999218,I999210);
not I_58567 (I999235,I425137);
not I_58568 (I999252,I425122);
nor I_58569 (I999269,I999252,I425131);
nor I_58570 (I998882,I999218,I999269);
nor I_58571 (I999300,I999252,I425134);
and I_58572 (I999317,I999300,I425122);
or I_58573 (I999334,I999317,I425146);
DFFARX1 I_58574 (I999334,I3563,I998890,I999360,);
nor I_58575 (I998870,I999360,I998916);
not I_58576 (I999382,I999360);
and I_58577 (I999399,I999382,I998916);
nor I_58578 (I998864,I998941,I999399);
nand I_58579 (I999430,I999382,I998992);
nor I_58580 (I998858,I999252,I999430);
nand I_58581 (I998861,I999382,I999170);
nand I_58582 (I999475,I998992,I425122);
nor I_58583 (I998873,I999235,I999475);
not I_58584 (I999536,I3570);
DFFARX1 I_58585 (I99861,I3563,I999536,I999562,);
DFFARX1 I_58586 (I99867,I3563,I999536,I999579,);
not I_58587 (I999587,I999579);
not I_58588 (I999604,I99885);
nor I_58589 (I999621,I999604,I99864);
not I_58590 (I999638,I99870);
nor I_58591 (I999655,I999621,I99876);
nor I_58592 (I999672,I999579,I999655);
DFFARX1 I_58593 (I999672,I3563,I999536,I999522,);
nor I_58594 (I999703,I99876,I99864);
nand I_58595 (I999720,I999703,I99885);
DFFARX1 I_58596 (I999720,I3563,I999536,I999525,);
nor I_58597 (I999751,I999638,I99876);
nand I_58598 (I999768,I999751,I99882);
nor I_58599 (I999785,I999562,I999768);
DFFARX1 I_58600 (I999785,I3563,I999536,I999501,);
not I_58601 (I999816,I999768);
nand I_58602 (I999513,I999579,I999816);
DFFARX1 I_58603 (I999768,I3563,I999536,I999856,);
not I_58604 (I999864,I999856);
not I_58605 (I999881,I99876);
not I_58606 (I999898,I99864);
nor I_58607 (I999915,I999898,I99870);
nor I_58608 (I999528,I999864,I999915);
nor I_58609 (I999946,I999898,I99873);
and I_58610 (I999963,I999946,I99861);
or I_58611 (I999980,I999963,I99879);
DFFARX1 I_58612 (I999980,I3563,I999536,I1000006,);
nor I_58613 (I999516,I1000006,I999562);
not I_58614 (I1000028,I1000006);
and I_58615 (I1000045,I1000028,I999562);
nor I_58616 (I999510,I999587,I1000045);
nand I_58617 (I1000076,I1000028,I999638);
nor I_58618 (I999504,I999898,I1000076);
nand I_58619 (I999507,I1000028,I999816);
nand I_58620 (I1000121,I999638,I99864);
nor I_58621 (I999519,I999881,I1000121);
not I_58622 (I1000182,I3570);
DFFARX1 I_58623 (I38202,I3563,I1000182,I1000208,);
DFFARX1 I_58624 (I38208,I3563,I1000182,I1000225,);
not I_58625 (I1000233,I1000225);
not I_58626 (I1000250,I38202);
nor I_58627 (I1000267,I1000250,I38214);
not I_58628 (I1000284,I38226);
nor I_58629 (I1000301,I1000267,I38220);
nor I_58630 (I1000318,I1000225,I1000301);
DFFARX1 I_58631 (I1000318,I3563,I1000182,I1000168,);
nor I_58632 (I1000349,I38220,I38214);
nand I_58633 (I1000366,I1000349,I38202);
DFFARX1 I_58634 (I1000366,I3563,I1000182,I1000171,);
nor I_58635 (I1000397,I1000284,I38220);
nand I_58636 (I1000414,I1000397,I38205);
nor I_58637 (I1000431,I1000208,I1000414);
DFFARX1 I_58638 (I1000431,I3563,I1000182,I1000147,);
not I_58639 (I1000462,I1000414);
nand I_58640 (I1000159,I1000225,I1000462);
DFFARX1 I_58641 (I1000414,I3563,I1000182,I1000502,);
not I_58642 (I1000510,I1000502);
not I_58643 (I1000527,I38220);
not I_58644 (I1000544,I38205);
nor I_58645 (I1000561,I1000544,I38226);
nor I_58646 (I1000174,I1000510,I1000561);
nor I_58647 (I1000592,I1000544,I38223);
and I_58648 (I1000609,I1000592,I38217);
or I_58649 (I1000626,I1000609,I38211);
DFFARX1 I_58650 (I1000626,I3563,I1000182,I1000652,);
nor I_58651 (I1000162,I1000652,I1000208);
not I_58652 (I1000674,I1000652);
and I_58653 (I1000691,I1000674,I1000208);
nor I_58654 (I1000156,I1000233,I1000691);
nand I_58655 (I1000722,I1000674,I1000284);
nor I_58656 (I1000150,I1000544,I1000722);
nand I_58657 (I1000153,I1000674,I1000462);
nand I_58658 (I1000767,I1000284,I38205);
nor I_58659 (I1000165,I1000527,I1000767);
not I_58660 (I1000828,I3570);
DFFARX1 I_58661 (I583276,I3563,I1000828,I1000854,);
DFFARX1 I_58662 (I583288,I3563,I1000828,I1000871,);
not I_58663 (I1000879,I1000871);
not I_58664 (I1000896,I583297);
nor I_58665 (I1000913,I1000896,I583273);
not I_58666 (I1000930,I583291);
nor I_58667 (I1000947,I1000913,I583285);
nor I_58668 (I1000964,I1000871,I1000947);
DFFARX1 I_58669 (I1000964,I3563,I1000828,I1000814,);
nor I_58670 (I1000995,I583285,I583273);
nand I_58671 (I1001012,I1000995,I583297);
DFFARX1 I_58672 (I1001012,I3563,I1000828,I1000817,);
nor I_58673 (I1001043,I1000930,I583285);
nand I_58674 (I1001060,I1001043,I583279);
nor I_58675 (I1001077,I1000854,I1001060);
DFFARX1 I_58676 (I1001077,I3563,I1000828,I1000793,);
not I_58677 (I1001108,I1001060);
nand I_58678 (I1000805,I1000871,I1001108);
DFFARX1 I_58679 (I1001060,I3563,I1000828,I1001148,);
not I_58680 (I1001156,I1001148);
not I_58681 (I1001173,I583285);
not I_58682 (I1001190,I583294);
nor I_58683 (I1001207,I1001190,I583291);
nor I_58684 (I1000820,I1001156,I1001207);
nor I_58685 (I1001238,I1001190,I583276);
and I_58686 (I1001255,I1001238,I583273);
or I_58687 (I1001272,I1001255,I583282);
DFFARX1 I_58688 (I1001272,I3563,I1000828,I1001298,);
nor I_58689 (I1000808,I1001298,I1000854);
not I_58690 (I1001320,I1001298);
and I_58691 (I1001337,I1001320,I1000854);
nor I_58692 (I1000802,I1000879,I1001337);
nand I_58693 (I1001368,I1001320,I1000930);
nor I_58694 (I1000796,I1001190,I1001368);
nand I_58695 (I1000799,I1001320,I1001108);
nand I_58696 (I1001413,I1000930,I583294);
nor I_58697 (I1000811,I1001173,I1001413);
not I_58698 (I1001474,I3570);
DFFARX1 I_58699 (I775753,I3563,I1001474,I1001500,);
DFFARX1 I_58700 (I775747,I3563,I1001474,I1001517,);
not I_58701 (I1001525,I1001517);
not I_58702 (I1001542,I775762);
nor I_58703 (I1001559,I1001542,I775747);
not I_58704 (I1001576,I775756);
nor I_58705 (I1001593,I1001559,I775765);
nor I_58706 (I1001610,I1001517,I1001593);
DFFARX1 I_58707 (I1001610,I3563,I1001474,I1001460,);
nor I_58708 (I1001641,I775765,I775747);
nand I_58709 (I1001658,I1001641,I775762);
DFFARX1 I_58710 (I1001658,I3563,I1001474,I1001463,);
nor I_58711 (I1001689,I1001576,I775765);
nand I_58712 (I1001706,I1001689,I775750);
nor I_58713 (I1001723,I1001500,I1001706);
DFFARX1 I_58714 (I1001723,I3563,I1001474,I1001439,);
not I_58715 (I1001754,I1001706);
nand I_58716 (I1001451,I1001517,I1001754);
DFFARX1 I_58717 (I1001706,I3563,I1001474,I1001794,);
not I_58718 (I1001802,I1001794);
not I_58719 (I1001819,I775765);
not I_58720 (I1001836,I775759);
nor I_58721 (I1001853,I1001836,I775756);
nor I_58722 (I1001466,I1001802,I1001853);
nor I_58723 (I1001884,I1001836,I775768);
and I_58724 (I1001901,I1001884,I775771);
or I_58725 (I1001918,I1001901,I775750);
DFFARX1 I_58726 (I1001918,I3563,I1001474,I1001944,);
nor I_58727 (I1001454,I1001944,I1001500);
not I_58728 (I1001966,I1001944);
and I_58729 (I1001983,I1001966,I1001500);
nor I_58730 (I1001448,I1001525,I1001983);
nand I_58731 (I1002014,I1001966,I1001576);
nor I_58732 (I1001442,I1001836,I1002014);
nand I_58733 (I1001445,I1001966,I1001754);
nand I_58734 (I1002059,I1001576,I775759);
nor I_58735 (I1001457,I1001819,I1002059);
not I_58736 (I1002120,I3570);
DFFARX1 I_58737 (I683851,I3563,I1002120,I1002146,);
DFFARX1 I_58738 (I683845,I3563,I1002120,I1002163,);
not I_58739 (I1002171,I1002163);
not I_58740 (I1002188,I683860);
nor I_58741 (I1002205,I1002188,I683845);
not I_58742 (I1002222,I683854);
nor I_58743 (I1002239,I1002205,I683863);
nor I_58744 (I1002256,I1002163,I1002239);
DFFARX1 I_58745 (I1002256,I3563,I1002120,I1002106,);
nor I_58746 (I1002287,I683863,I683845);
nand I_58747 (I1002304,I1002287,I683860);
DFFARX1 I_58748 (I1002304,I3563,I1002120,I1002109,);
nor I_58749 (I1002335,I1002222,I683863);
nand I_58750 (I1002352,I1002335,I683848);
nor I_58751 (I1002369,I1002146,I1002352);
DFFARX1 I_58752 (I1002369,I3563,I1002120,I1002085,);
not I_58753 (I1002400,I1002352);
nand I_58754 (I1002097,I1002163,I1002400);
DFFARX1 I_58755 (I1002352,I3563,I1002120,I1002440,);
not I_58756 (I1002448,I1002440);
not I_58757 (I1002465,I683863);
not I_58758 (I1002482,I683857);
nor I_58759 (I1002499,I1002482,I683854);
nor I_58760 (I1002112,I1002448,I1002499);
nor I_58761 (I1002530,I1002482,I683866);
and I_58762 (I1002547,I1002530,I683869);
or I_58763 (I1002564,I1002547,I683848);
DFFARX1 I_58764 (I1002564,I3563,I1002120,I1002590,);
nor I_58765 (I1002100,I1002590,I1002146);
not I_58766 (I1002612,I1002590);
and I_58767 (I1002629,I1002612,I1002146);
nor I_58768 (I1002094,I1002171,I1002629);
nand I_58769 (I1002660,I1002612,I1002222);
nor I_58770 (I1002088,I1002482,I1002660);
nand I_58771 (I1002091,I1002612,I1002400);
nand I_58772 (I1002705,I1002222,I683857);
nor I_58773 (I1002103,I1002465,I1002705);
not I_58774 (I1002766,I3570);
DFFARX1 I_58775 (I551299,I3563,I1002766,I1002792,);
DFFARX1 I_58776 (I551311,I3563,I1002766,I1002809,);
not I_58777 (I1002817,I1002809);
not I_58778 (I1002834,I551296);
nor I_58779 (I1002851,I1002834,I551314);
not I_58780 (I1002868,I551320);
nor I_58781 (I1002885,I1002851,I551302);
nor I_58782 (I1002902,I1002809,I1002885);
DFFARX1 I_58783 (I1002902,I3563,I1002766,I1002752,);
nor I_58784 (I1002933,I551302,I551314);
nand I_58785 (I1002950,I1002933,I551296);
DFFARX1 I_58786 (I1002950,I3563,I1002766,I1002755,);
nor I_58787 (I1002981,I1002868,I551302);
nand I_58788 (I1002998,I1002981,I551305);
nor I_58789 (I1003015,I1002792,I1002998);
DFFARX1 I_58790 (I1003015,I3563,I1002766,I1002731,);
not I_58791 (I1003046,I1002998);
nand I_58792 (I1002743,I1002809,I1003046);
DFFARX1 I_58793 (I1002998,I3563,I1002766,I1003086,);
not I_58794 (I1003094,I1003086);
not I_58795 (I1003111,I551302);
not I_58796 (I1003128,I551308);
nor I_58797 (I1003145,I1003128,I551320);
nor I_58798 (I1002758,I1003094,I1003145);
nor I_58799 (I1003176,I1003128,I551317);
and I_58800 (I1003193,I1003176,I551296);
or I_58801 (I1003210,I1003193,I551299);
DFFARX1 I_58802 (I1003210,I3563,I1002766,I1003236,);
nor I_58803 (I1002746,I1003236,I1002792);
not I_58804 (I1003258,I1003236);
and I_58805 (I1003275,I1003258,I1002792);
nor I_58806 (I1002740,I1002817,I1003275);
nand I_58807 (I1003306,I1003258,I1002868);
nor I_58808 (I1002734,I1003128,I1003306);
nand I_58809 (I1002737,I1003258,I1003046);
nand I_58810 (I1003351,I1002868,I551308);
nor I_58811 (I1002749,I1003111,I1003351);
not I_58812 (I1003412,I3570);
DFFARX1 I_58813 (I857965,I3563,I1003412,I1003438,);
DFFARX1 I_58814 (I857962,I3563,I1003412,I1003455,);
not I_58815 (I1003463,I1003455);
not I_58816 (I1003480,I857962);
nor I_58817 (I1003497,I1003480,I857965);
not I_58818 (I1003514,I857977);
nor I_58819 (I1003531,I1003497,I857971);
nor I_58820 (I1003548,I1003455,I1003531);
DFFARX1 I_58821 (I1003548,I3563,I1003412,I1003398,);
nor I_58822 (I1003579,I857971,I857965);
nand I_58823 (I1003596,I1003579,I857962);
DFFARX1 I_58824 (I1003596,I3563,I1003412,I1003401,);
nor I_58825 (I1003627,I1003514,I857971);
nand I_58826 (I1003644,I1003627,I857959);
nor I_58827 (I1003661,I1003438,I1003644);
DFFARX1 I_58828 (I1003661,I3563,I1003412,I1003377,);
not I_58829 (I1003692,I1003644);
nand I_58830 (I1003389,I1003455,I1003692);
DFFARX1 I_58831 (I1003644,I3563,I1003412,I1003732,);
not I_58832 (I1003740,I1003732);
not I_58833 (I1003757,I857971);
not I_58834 (I1003774,I857968);
nor I_58835 (I1003791,I1003774,I857977);
nor I_58836 (I1003404,I1003740,I1003791);
nor I_58837 (I1003822,I1003774,I857974);
and I_58838 (I1003839,I1003822,I857980);
or I_58839 (I1003856,I1003839,I857959);
DFFARX1 I_58840 (I1003856,I3563,I1003412,I1003882,);
nor I_58841 (I1003392,I1003882,I1003438);
not I_58842 (I1003904,I1003882);
and I_58843 (I1003921,I1003904,I1003438);
nor I_58844 (I1003386,I1003463,I1003921);
nand I_58845 (I1003952,I1003904,I1003514);
nor I_58846 (I1003380,I1003774,I1003952);
nand I_58847 (I1003383,I1003904,I1003692);
nand I_58848 (I1003997,I1003514,I857968);
nor I_58849 (I1003395,I1003757,I1003997);
not I_58850 (I1004058,I3570);
DFFARX1 I_58851 (I116725,I3563,I1004058,I1004084,);
DFFARX1 I_58852 (I116731,I3563,I1004058,I1004101,);
not I_58853 (I1004109,I1004101);
not I_58854 (I1004126,I116749);
nor I_58855 (I1004143,I1004126,I116728);
not I_58856 (I1004160,I116734);
nor I_58857 (I1004177,I1004143,I116740);
nor I_58858 (I1004194,I1004101,I1004177);
DFFARX1 I_58859 (I1004194,I3563,I1004058,I1004044,);
nor I_58860 (I1004225,I116740,I116728);
nand I_58861 (I1004242,I1004225,I116749);
DFFARX1 I_58862 (I1004242,I3563,I1004058,I1004047,);
nor I_58863 (I1004273,I1004160,I116740);
nand I_58864 (I1004290,I1004273,I116746);
nor I_58865 (I1004307,I1004084,I1004290);
DFFARX1 I_58866 (I1004307,I3563,I1004058,I1004023,);
not I_58867 (I1004338,I1004290);
nand I_58868 (I1004035,I1004101,I1004338);
DFFARX1 I_58869 (I1004290,I3563,I1004058,I1004378,);
not I_58870 (I1004386,I1004378);
not I_58871 (I1004403,I116740);
not I_58872 (I1004420,I116728);
nor I_58873 (I1004437,I1004420,I116734);
nor I_58874 (I1004050,I1004386,I1004437);
nor I_58875 (I1004468,I1004420,I116737);
and I_58876 (I1004485,I1004468,I116725);
or I_58877 (I1004502,I1004485,I116743);
DFFARX1 I_58878 (I1004502,I3563,I1004058,I1004528,);
nor I_58879 (I1004038,I1004528,I1004084);
not I_58880 (I1004550,I1004528);
and I_58881 (I1004567,I1004550,I1004084);
nor I_58882 (I1004032,I1004109,I1004567);
nand I_58883 (I1004598,I1004550,I1004160);
nor I_58884 (I1004026,I1004420,I1004598);
nand I_58885 (I1004029,I1004550,I1004338);
nand I_58886 (I1004643,I1004160,I116728);
nor I_58887 (I1004041,I1004403,I1004643);
not I_58888 (I1004704,I3570);
DFFARX1 I_58889 (I1307992,I3563,I1004704,I1004730,);
DFFARX1 I_58890 (I1307986,I3563,I1004704,I1004747,);
not I_58891 (I1004755,I1004747);
not I_58892 (I1004772,I1307995);
nor I_58893 (I1004789,I1004772,I1308007);
not I_58894 (I1004806,I1307989);
nor I_58895 (I1004823,I1004789,I1307986);
nor I_58896 (I1004840,I1004747,I1004823);
DFFARX1 I_58897 (I1004840,I3563,I1004704,I1004690,);
nor I_58898 (I1004871,I1307986,I1308007);
nand I_58899 (I1004888,I1004871,I1307995);
DFFARX1 I_58900 (I1004888,I3563,I1004704,I1004693,);
nor I_58901 (I1004919,I1004806,I1307986);
nand I_58902 (I1004936,I1004919,I1307983);
nor I_58903 (I1004953,I1004730,I1004936);
DFFARX1 I_58904 (I1004953,I3563,I1004704,I1004669,);
not I_58905 (I1004984,I1004936);
nand I_58906 (I1004681,I1004747,I1004984);
DFFARX1 I_58907 (I1004936,I3563,I1004704,I1005024,);
not I_58908 (I1005032,I1005024);
not I_58909 (I1005049,I1307986);
not I_58910 (I1005066,I1308004);
nor I_58911 (I1005083,I1005066,I1307989);
nor I_58912 (I1004696,I1005032,I1005083);
nor I_58913 (I1005114,I1005066,I1307998);
and I_58914 (I1005131,I1005114,I1307983);
or I_58915 (I1005148,I1005131,I1308001);
DFFARX1 I_58916 (I1005148,I3563,I1004704,I1005174,);
nor I_58917 (I1004684,I1005174,I1004730);
not I_58918 (I1005196,I1005174);
and I_58919 (I1005213,I1005196,I1004730);
nor I_58920 (I1004678,I1004755,I1005213);
nand I_58921 (I1005244,I1005196,I1004806);
nor I_58922 (I1004672,I1005066,I1005244);
nand I_58923 (I1004675,I1005196,I1004984);
nand I_58924 (I1005289,I1004806,I1308004);
nor I_58925 (I1004687,I1005049,I1005289);
not I_58926 (I1005350,I3570);
DFFARX1 I_58927 (I1202567,I3563,I1005350,I1005376,);
DFFARX1 I_58928 (I1202549,I3563,I1005350,I1005393,);
not I_58929 (I1005401,I1005393);
not I_58930 (I1005418,I1202558);
nor I_58931 (I1005435,I1005418,I1202570);
not I_58932 (I1005452,I1202552);
nor I_58933 (I1005469,I1005435,I1202561);
nor I_58934 (I1005486,I1005393,I1005469);
DFFARX1 I_58935 (I1005486,I3563,I1005350,I1005336,);
nor I_58936 (I1005517,I1202561,I1202570);
nand I_58937 (I1005534,I1005517,I1202558);
DFFARX1 I_58938 (I1005534,I3563,I1005350,I1005339,);
nor I_58939 (I1005565,I1005452,I1202561);
nand I_58940 (I1005582,I1005565,I1202573);
nor I_58941 (I1005599,I1005376,I1005582);
DFFARX1 I_58942 (I1005599,I3563,I1005350,I1005315,);
not I_58943 (I1005630,I1005582);
nand I_58944 (I1005327,I1005393,I1005630);
DFFARX1 I_58945 (I1005582,I3563,I1005350,I1005670,);
not I_58946 (I1005678,I1005670);
not I_58947 (I1005695,I1202561);
not I_58948 (I1005712,I1202549);
nor I_58949 (I1005729,I1005712,I1202552);
nor I_58950 (I1005342,I1005678,I1005729);
nor I_58951 (I1005760,I1005712,I1202555);
and I_58952 (I1005777,I1005760,I1202564);
or I_58953 (I1005794,I1005777,I1202552);
DFFARX1 I_58954 (I1005794,I3563,I1005350,I1005820,);
nor I_58955 (I1005330,I1005820,I1005376);
not I_58956 (I1005842,I1005820);
and I_58957 (I1005859,I1005842,I1005376);
nor I_58958 (I1005324,I1005401,I1005859);
nand I_58959 (I1005890,I1005842,I1005452);
nor I_58960 (I1005318,I1005712,I1005890);
nand I_58961 (I1005321,I1005842,I1005630);
nand I_58962 (I1005935,I1005452,I1202549);
nor I_58963 (I1005333,I1005695,I1005935);
not I_58964 (I1005996,I3570);
DFFARX1 I_58965 (I860600,I3563,I1005996,I1006022,);
DFFARX1 I_58966 (I860597,I3563,I1005996,I1006039,);
not I_58967 (I1006047,I1006039);
not I_58968 (I1006064,I860597);
nor I_58969 (I1006081,I1006064,I860600);
not I_58970 (I1006098,I860612);
nor I_58971 (I1006115,I1006081,I860606);
nor I_58972 (I1006132,I1006039,I1006115);
DFFARX1 I_58973 (I1006132,I3563,I1005996,I1005982,);
nor I_58974 (I1006163,I860606,I860600);
nand I_58975 (I1006180,I1006163,I860597);
DFFARX1 I_58976 (I1006180,I3563,I1005996,I1005985,);
nor I_58977 (I1006211,I1006098,I860606);
nand I_58978 (I1006228,I1006211,I860594);
nor I_58979 (I1006245,I1006022,I1006228);
DFFARX1 I_58980 (I1006245,I3563,I1005996,I1005961,);
not I_58981 (I1006276,I1006228);
nand I_58982 (I1005973,I1006039,I1006276);
DFFARX1 I_58983 (I1006228,I3563,I1005996,I1006316,);
not I_58984 (I1006324,I1006316);
not I_58985 (I1006341,I860606);
not I_58986 (I1006358,I860603);
nor I_58987 (I1006375,I1006358,I860612);
nor I_58988 (I1005988,I1006324,I1006375);
nor I_58989 (I1006406,I1006358,I860609);
and I_58990 (I1006423,I1006406,I860615);
or I_58991 (I1006440,I1006423,I860594);
DFFARX1 I_58992 (I1006440,I3563,I1005996,I1006466,);
nor I_58993 (I1005976,I1006466,I1006022);
not I_58994 (I1006488,I1006466);
and I_58995 (I1006505,I1006488,I1006022);
nor I_58996 (I1005970,I1006047,I1006505);
nand I_58997 (I1006536,I1006488,I1006098);
nor I_58998 (I1005964,I1006358,I1006536);
nand I_58999 (I1005967,I1006488,I1006276);
nand I_59000 (I1006581,I1006098,I860603);
nor I_59001 (I1005979,I1006341,I1006581);
not I_59002 (I1006642,I3570);
DFFARX1 I_59003 (I424584,I3563,I1006642,I1006668,);
DFFARX1 I_59004 (I424581,I3563,I1006642,I1006685,);
not I_59005 (I1006693,I1006685);
not I_59006 (I1006710,I424596);
nor I_59007 (I1006727,I1006710,I424599);
not I_59008 (I1006744,I424587);
nor I_59009 (I1006761,I1006727,I424593);
nor I_59010 (I1006778,I1006685,I1006761);
DFFARX1 I_59011 (I1006778,I3563,I1006642,I1006628,);
nor I_59012 (I1006809,I424593,I424599);
nand I_59013 (I1006826,I1006809,I424596);
DFFARX1 I_59014 (I1006826,I3563,I1006642,I1006631,);
nor I_59015 (I1006857,I1006744,I424593);
nand I_59016 (I1006874,I1006857,I424605);
nor I_59017 (I1006891,I1006668,I1006874);
DFFARX1 I_59018 (I1006891,I3563,I1006642,I1006607,);
not I_59019 (I1006922,I1006874);
nand I_59020 (I1006619,I1006685,I1006922);
DFFARX1 I_59021 (I1006874,I3563,I1006642,I1006962,);
not I_59022 (I1006970,I1006962);
not I_59023 (I1006987,I424593);
not I_59024 (I1007004,I424578);
nor I_59025 (I1007021,I1007004,I424587);
nor I_59026 (I1006634,I1006970,I1007021);
nor I_59027 (I1007052,I1007004,I424590);
and I_59028 (I1007069,I1007052,I424578);
or I_59029 (I1007086,I1007069,I424602);
DFFARX1 I_59030 (I1007086,I3563,I1006642,I1007112,);
nor I_59031 (I1006622,I1007112,I1006668);
not I_59032 (I1007134,I1007112);
and I_59033 (I1007151,I1007134,I1006668);
nor I_59034 (I1006616,I1006693,I1007151);
nand I_59035 (I1007182,I1007134,I1006744);
nor I_59036 (I1006610,I1007004,I1007182);
nand I_59037 (I1006613,I1007134,I1006922);
nand I_59038 (I1007227,I1006744,I424578);
nor I_59039 (I1006625,I1006987,I1007227);
not I_59040 (I1007288,I3570);
DFFARX1 I_59041 (I335957,I3563,I1007288,I1007314,);
DFFARX1 I_59042 (I335963,I3563,I1007288,I1007331,);
not I_59043 (I1007339,I1007331);
not I_59044 (I1007356,I335984);
nor I_59045 (I1007373,I1007356,I335972);
not I_59046 (I1007390,I335981);
nor I_59047 (I1007407,I1007373,I335966);
nor I_59048 (I1007424,I1007331,I1007407);
DFFARX1 I_59049 (I1007424,I3563,I1007288,I1007274,);
nor I_59050 (I1007455,I335966,I335972);
nand I_59051 (I1007472,I1007455,I335984);
DFFARX1 I_59052 (I1007472,I3563,I1007288,I1007277,);
nor I_59053 (I1007503,I1007390,I335966);
nand I_59054 (I1007520,I1007503,I335957);
nor I_59055 (I1007537,I1007314,I1007520);
DFFARX1 I_59056 (I1007537,I3563,I1007288,I1007253,);
not I_59057 (I1007568,I1007520);
nand I_59058 (I1007265,I1007331,I1007568);
DFFARX1 I_59059 (I1007520,I3563,I1007288,I1007608,);
not I_59060 (I1007616,I1007608);
not I_59061 (I1007633,I335966);
not I_59062 (I1007650,I335969);
nor I_59063 (I1007667,I1007650,I335981);
nor I_59064 (I1007280,I1007616,I1007667);
nor I_59065 (I1007698,I1007650,I335978);
and I_59066 (I1007715,I1007698,I335960);
or I_59067 (I1007732,I1007715,I335975);
DFFARX1 I_59068 (I1007732,I3563,I1007288,I1007758,);
nor I_59069 (I1007268,I1007758,I1007314);
not I_59070 (I1007780,I1007758);
and I_59071 (I1007797,I1007780,I1007314);
nor I_59072 (I1007262,I1007339,I1007797);
nand I_59073 (I1007828,I1007780,I1007390);
nor I_59074 (I1007256,I1007650,I1007828);
nand I_59075 (I1007259,I1007780,I1007568);
nand I_59076 (I1007873,I1007390,I335969);
nor I_59077 (I1007271,I1007633,I1007873);
not I_59078 (I1007934,I3570);
DFFARX1 I_59079 (I557249,I3563,I1007934,I1007960,);
DFFARX1 I_59080 (I557261,I3563,I1007934,I1007977,);
not I_59081 (I1007985,I1007977);
not I_59082 (I1008002,I557246);
nor I_59083 (I1008019,I1008002,I557264);
not I_59084 (I1008036,I557270);
nor I_59085 (I1008053,I1008019,I557252);
nor I_59086 (I1008070,I1007977,I1008053);
DFFARX1 I_59087 (I1008070,I3563,I1007934,I1007920,);
nor I_59088 (I1008101,I557252,I557264);
nand I_59089 (I1008118,I1008101,I557246);
DFFARX1 I_59090 (I1008118,I3563,I1007934,I1007923,);
nor I_59091 (I1008149,I1008036,I557252);
nand I_59092 (I1008166,I1008149,I557255);
nor I_59093 (I1008183,I1007960,I1008166);
DFFARX1 I_59094 (I1008183,I3563,I1007934,I1007899,);
not I_59095 (I1008214,I1008166);
nand I_59096 (I1007911,I1007977,I1008214);
DFFARX1 I_59097 (I1008166,I3563,I1007934,I1008254,);
not I_59098 (I1008262,I1008254);
not I_59099 (I1008279,I557252);
not I_59100 (I1008296,I557258);
nor I_59101 (I1008313,I1008296,I557270);
nor I_59102 (I1007926,I1008262,I1008313);
nor I_59103 (I1008344,I1008296,I557267);
and I_59104 (I1008361,I1008344,I557246);
or I_59105 (I1008378,I1008361,I557249);
DFFARX1 I_59106 (I1008378,I3563,I1007934,I1008404,);
nor I_59107 (I1007914,I1008404,I1007960);
not I_59108 (I1008426,I1008404);
and I_59109 (I1008443,I1008426,I1007960);
nor I_59110 (I1007908,I1007985,I1008443);
nand I_59111 (I1008474,I1008426,I1008036);
nor I_59112 (I1007902,I1008296,I1008474);
nand I_59113 (I1007905,I1008426,I1008214);
nand I_59114 (I1008519,I1008036,I557258);
nor I_59115 (I1007917,I1008279,I1008519);
not I_59116 (I1008580,I3570);
DFFARX1 I_59117 (I501288,I3563,I1008580,I1008606,);
DFFARX1 I_59118 (I501285,I3563,I1008580,I1008623,);
not I_59119 (I1008631,I1008623);
not I_59120 (I1008648,I501300);
nor I_59121 (I1008665,I1008648,I501303);
not I_59122 (I1008682,I501291);
nor I_59123 (I1008699,I1008665,I501297);
nor I_59124 (I1008716,I1008623,I1008699);
DFFARX1 I_59125 (I1008716,I3563,I1008580,I1008566,);
nor I_59126 (I1008747,I501297,I501303);
nand I_59127 (I1008764,I1008747,I501300);
DFFARX1 I_59128 (I1008764,I3563,I1008580,I1008569,);
nor I_59129 (I1008795,I1008682,I501297);
nand I_59130 (I1008812,I1008795,I501309);
nor I_59131 (I1008829,I1008606,I1008812);
DFFARX1 I_59132 (I1008829,I3563,I1008580,I1008545,);
not I_59133 (I1008860,I1008812);
nand I_59134 (I1008557,I1008623,I1008860);
DFFARX1 I_59135 (I1008812,I3563,I1008580,I1008900,);
not I_59136 (I1008908,I1008900);
not I_59137 (I1008925,I501297);
not I_59138 (I1008942,I501282);
nor I_59139 (I1008959,I1008942,I501291);
nor I_59140 (I1008572,I1008908,I1008959);
nor I_59141 (I1008990,I1008942,I501294);
and I_59142 (I1009007,I1008990,I501282);
or I_59143 (I1009024,I1009007,I501306);
DFFARX1 I_59144 (I1009024,I3563,I1008580,I1009050,);
nor I_59145 (I1008560,I1009050,I1008606);
not I_59146 (I1009072,I1009050);
and I_59147 (I1009089,I1009072,I1008606);
nor I_59148 (I1008554,I1008631,I1009089);
nand I_59149 (I1009120,I1009072,I1008682);
nor I_59150 (I1008548,I1008942,I1009120);
nand I_59151 (I1008551,I1009072,I1008860);
nand I_59152 (I1009165,I1008682,I501282);
nor I_59153 (I1008563,I1008925,I1009165);
not I_59154 (I1009226,I3570);
DFFARX1 I_59155 (I1078636,I3563,I1009226,I1009252,);
DFFARX1 I_59156 (I1078639,I3563,I1009226,I1009269,);
not I_59157 (I1009277,I1009269);
not I_59158 (I1009294,I1078636);
nor I_59159 (I1009311,I1009294,I1078648);
not I_59160 (I1009328,I1078657);
nor I_59161 (I1009345,I1009311,I1078645);
nor I_59162 (I1009362,I1009269,I1009345);
DFFARX1 I_59163 (I1009362,I3563,I1009226,I1009212,);
nor I_59164 (I1009393,I1078645,I1078648);
nand I_59165 (I1009410,I1009393,I1078636);
DFFARX1 I_59166 (I1009410,I3563,I1009226,I1009215,);
nor I_59167 (I1009441,I1009328,I1078645);
nand I_59168 (I1009458,I1009441,I1078651);
nor I_59169 (I1009475,I1009252,I1009458);
DFFARX1 I_59170 (I1009475,I3563,I1009226,I1009191,);
not I_59171 (I1009506,I1009458);
nand I_59172 (I1009203,I1009269,I1009506);
DFFARX1 I_59173 (I1009458,I3563,I1009226,I1009546,);
not I_59174 (I1009554,I1009546);
not I_59175 (I1009571,I1078645);
not I_59176 (I1009588,I1078642);
nor I_59177 (I1009605,I1009588,I1078657);
nor I_59178 (I1009218,I1009554,I1009605);
nor I_59179 (I1009636,I1009588,I1078654);
and I_59180 (I1009653,I1009636,I1078642);
or I_59181 (I1009670,I1009653,I1078639);
DFFARX1 I_59182 (I1009670,I3563,I1009226,I1009696,);
nor I_59183 (I1009206,I1009696,I1009252);
not I_59184 (I1009718,I1009696);
and I_59185 (I1009735,I1009718,I1009252);
nor I_59186 (I1009200,I1009277,I1009735);
nand I_59187 (I1009766,I1009718,I1009328);
nor I_59188 (I1009194,I1009588,I1009766);
nand I_59189 (I1009197,I1009718,I1009506);
nand I_59190 (I1009811,I1009328,I1078642);
nor I_59191 (I1009209,I1009571,I1009811);
not I_59192 (I1009872,I3570);
DFFARX1 I_59193 (I790781,I3563,I1009872,I1009898,);
DFFARX1 I_59194 (I790775,I3563,I1009872,I1009915,);
not I_59195 (I1009923,I1009915);
not I_59196 (I1009940,I790790);
nor I_59197 (I1009957,I1009940,I790775);
not I_59198 (I1009974,I790784);
nor I_59199 (I1009991,I1009957,I790793);
nor I_59200 (I1010008,I1009915,I1009991);
DFFARX1 I_59201 (I1010008,I3563,I1009872,I1009858,);
nor I_59202 (I1010039,I790793,I790775);
nand I_59203 (I1010056,I1010039,I790790);
DFFARX1 I_59204 (I1010056,I3563,I1009872,I1009861,);
nor I_59205 (I1010087,I1009974,I790793);
nand I_59206 (I1010104,I1010087,I790778);
nor I_59207 (I1010121,I1009898,I1010104);
DFFARX1 I_59208 (I1010121,I3563,I1009872,I1009837,);
not I_59209 (I1010152,I1010104);
nand I_59210 (I1009849,I1009915,I1010152);
DFFARX1 I_59211 (I1010104,I3563,I1009872,I1010192,);
not I_59212 (I1010200,I1010192);
not I_59213 (I1010217,I790793);
not I_59214 (I1010234,I790787);
nor I_59215 (I1010251,I1010234,I790784);
nor I_59216 (I1009864,I1010200,I1010251);
nor I_59217 (I1010282,I1010234,I790796);
and I_59218 (I1010299,I1010282,I790799);
or I_59219 (I1010316,I1010299,I790778);
DFFARX1 I_59220 (I1010316,I3563,I1009872,I1010342,);
nor I_59221 (I1009852,I1010342,I1009898);
not I_59222 (I1010364,I1010342);
and I_59223 (I1010381,I1010364,I1009898);
nor I_59224 (I1009846,I1009923,I1010381);
nand I_59225 (I1010412,I1010364,I1009974);
nor I_59226 (I1009840,I1010234,I1010412);
nand I_59227 (I1009843,I1010364,I1010152);
nand I_59228 (I1010457,I1009974,I790787);
nor I_59229 (I1009855,I1010217,I1010457);
not I_59230 (I1010518,I3570);
DFFARX1 I_59231 (I1085368,I3563,I1010518,I1010544,);
DFFARX1 I_59232 (I1085371,I3563,I1010518,I1010561,);
not I_59233 (I1010569,I1010561);
not I_59234 (I1010586,I1085368);
nor I_59235 (I1010603,I1010586,I1085380);
not I_59236 (I1010620,I1085389);
nor I_59237 (I1010637,I1010603,I1085377);
nor I_59238 (I1010654,I1010561,I1010637);
DFFARX1 I_59239 (I1010654,I3563,I1010518,I1010504,);
nor I_59240 (I1010685,I1085377,I1085380);
nand I_59241 (I1010702,I1010685,I1085368);
DFFARX1 I_59242 (I1010702,I3563,I1010518,I1010507,);
nor I_59243 (I1010733,I1010620,I1085377);
nand I_59244 (I1010750,I1010733,I1085383);
nor I_59245 (I1010767,I1010544,I1010750);
DFFARX1 I_59246 (I1010767,I3563,I1010518,I1010483,);
not I_59247 (I1010798,I1010750);
nand I_59248 (I1010495,I1010561,I1010798);
DFFARX1 I_59249 (I1010750,I3563,I1010518,I1010838,);
not I_59250 (I1010846,I1010838);
not I_59251 (I1010863,I1085377);
not I_59252 (I1010880,I1085374);
nor I_59253 (I1010897,I1010880,I1085389);
nor I_59254 (I1010510,I1010846,I1010897);
nor I_59255 (I1010928,I1010880,I1085386);
and I_59256 (I1010945,I1010928,I1085374);
or I_59257 (I1010962,I1010945,I1085371);
DFFARX1 I_59258 (I1010962,I3563,I1010518,I1010988,);
nor I_59259 (I1010498,I1010988,I1010544);
not I_59260 (I1011010,I1010988);
and I_59261 (I1011027,I1011010,I1010544);
nor I_59262 (I1010492,I1010569,I1011027);
nand I_59263 (I1011058,I1011010,I1010620);
nor I_59264 (I1010486,I1010880,I1011058);
nand I_59265 (I1010489,I1011010,I1010798);
nand I_59266 (I1011103,I1010620,I1085374);
nor I_59267 (I1010501,I1010863,I1011103);
not I_59268 (I1011164,I3570);
DFFARX1 I_59269 (I185139,I3563,I1011164,I1011190,);
DFFARX1 I_59270 (I185151,I3563,I1011164,I1011207,);
not I_59271 (I1011215,I1011207);
not I_59272 (I1011232,I185157);
nor I_59273 (I1011249,I1011232,I185142);
not I_59274 (I1011266,I185133);
nor I_59275 (I1011283,I1011249,I185154);
nor I_59276 (I1011300,I1011207,I1011283);
DFFARX1 I_59277 (I1011300,I3563,I1011164,I1011150,);
nor I_59278 (I1011331,I185154,I185142);
nand I_59279 (I1011348,I1011331,I185157);
DFFARX1 I_59280 (I1011348,I3563,I1011164,I1011153,);
nor I_59281 (I1011379,I1011266,I185154);
nand I_59282 (I1011396,I1011379,I185136);
nor I_59283 (I1011413,I1011190,I1011396);
DFFARX1 I_59284 (I1011413,I3563,I1011164,I1011129,);
not I_59285 (I1011444,I1011396);
nand I_59286 (I1011141,I1011207,I1011444);
DFFARX1 I_59287 (I1011396,I3563,I1011164,I1011484,);
not I_59288 (I1011492,I1011484);
not I_59289 (I1011509,I185154);
not I_59290 (I1011526,I185145);
nor I_59291 (I1011543,I1011526,I185133);
nor I_59292 (I1011156,I1011492,I1011543);
nor I_59293 (I1011574,I1011526,I185148);
and I_59294 (I1011591,I1011574,I185136);
or I_59295 (I1011608,I1011591,I185133);
DFFARX1 I_59296 (I1011608,I3563,I1011164,I1011634,);
nor I_59297 (I1011144,I1011634,I1011190);
not I_59298 (I1011656,I1011634);
and I_59299 (I1011673,I1011656,I1011190);
nor I_59300 (I1011138,I1011215,I1011673);
nand I_59301 (I1011704,I1011656,I1011266);
nor I_59302 (I1011132,I1011526,I1011704);
nand I_59303 (I1011135,I1011656,I1011444);
nand I_59304 (I1011749,I1011266,I185145);
nor I_59305 (I1011147,I1011509,I1011749);
not I_59306 (I1011810,I3570);
DFFARX1 I_59307 (I97753,I3563,I1011810,I1011836,);
DFFARX1 I_59308 (I97759,I3563,I1011810,I1011853,);
not I_59309 (I1011861,I1011853);
not I_59310 (I1011878,I97777);
nor I_59311 (I1011895,I1011878,I97756);
not I_59312 (I1011912,I97762);
nor I_59313 (I1011929,I1011895,I97768);
nor I_59314 (I1011946,I1011853,I1011929);
DFFARX1 I_59315 (I1011946,I3563,I1011810,I1011796,);
nor I_59316 (I1011977,I97768,I97756);
nand I_59317 (I1011994,I1011977,I97777);
DFFARX1 I_59318 (I1011994,I3563,I1011810,I1011799,);
nor I_59319 (I1012025,I1011912,I97768);
nand I_59320 (I1012042,I1012025,I97774);
nor I_59321 (I1012059,I1011836,I1012042);
DFFARX1 I_59322 (I1012059,I3563,I1011810,I1011775,);
not I_59323 (I1012090,I1012042);
nand I_59324 (I1011787,I1011853,I1012090);
DFFARX1 I_59325 (I1012042,I3563,I1011810,I1012130,);
not I_59326 (I1012138,I1012130);
not I_59327 (I1012155,I97768);
not I_59328 (I1012172,I97756);
nor I_59329 (I1012189,I1012172,I97762);
nor I_59330 (I1011802,I1012138,I1012189);
nor I_59331 (I1012220,I1012172,I97765);
and I_59332 (I1012237,I1012220,I97753);
or I_59333 (I1012254,I1012237,I97771);
DFFARX1 I_59334 (I1012254,I3563,I1011810,I1012280,);
nor I_59335 (I1011790,I1012280,I1011836);
not I_59336 (I1012302,I1012280);
and I_59337 (I1012319,I1012302,I1011836);
nor I_59338 (I1011784,I1011861,I1012319);
nand I_59339 (I1012350,I1012302,I1011912);
nor I_59340 (I1011778,I1012172,I1012350);
nand I_59341 (I1011781,I1012302,I1012090);
nand I_59342 (I1012395,I1011912,I97756);
nor I_59343 (I1011793,I1012155,I1012395);
not I_59344 (I1012456,I3570);
DFFARX1 I_59345 (I1108931,I3563,I1012456,I1012482,);
DFFARX1 I_59346 (I1108913,I3563,I1012456,I1012499,);
not I_59347 (I1012507,I1012499);
not I_59348 (I1012524,I1108922);
nor I_59349 (I1012541,I1012524,I1108934);
not I_59350 (I1012558,I1108916);
nor I_59351 (I1012575,I1012541,I1108925);
nor I_59352 (I1012592,I1012499,I1012575);
DFFARX1 I_59353 (I1012592,I3563,I1012456,I1012442,);
nor I_59354 (I1012623,I1108925,I1108934);
nand I_59355 (I1012640,I1012623,I1108922);
DFFARX1 I_59356 (I1012640,I3563,I1012456,I1012445,);
nor I_59357 (I1012671,I1012558,I1108925);
nand I_59358 (I1012688,I1012671,I1108937);
nor I_59359 (I1012705,I1012482,I1012688);
DFFARX1 I_59360 (I1012705,I3563,I1012456,I1012421,);
not I_59361 (I1012736,I1012688);
nand I_59362 (I1012433,I1012499,I1012736);
DFFARX1 I_59363 (I1012688,I3563,I1012456,I1012776,);
not I_59364 (I1012784,I1012776);
not I_59365 (I1012801,I1108925);
not I_59366 (I1012818,I1108913);
nor I_59367 (I1012835,I1012818,I1108916);
nor I_59368 (I1012448,I1012784,I1012835);
nor I_59369 (I1012866,I1012818,I1108919);
and I_59370 (I1012883,I1012866,I1108928);
or I_59371 (I1012900,I1012883,I1108916);
DFFARX1 I_59372 (I1012900,I3563,I1012456,I1012926,);
nor I_59373 (I1012436,I1012926,I1012482);
not I_59374 (I1012948,I1012926);
and I_59375 (I1012965,I1012948,I1012482);
nor I_59376 (I1012430,I1012507,I1012965);
nand I_59377 (I1012996,I1012948,I1012558);
nor I_59378 (I1012424,I1012818,I1012996);
nand I_59379 (I1012427,I1012948,I1012736);
nand I_59380 (I1013041,I1012558,I1108913);
nor I_59381 (I1012439,I1012801,I1013041);
not I_59382 (I1013102,I3570);
DFFARX1 I_59383 (I417642,I3563,I1013102,I1013128,);
DFFARX1 I_59384 (I417648,I3563,I1013102,I1013145,);
not I_59385 (I1013153,I1013145);
not I_59386 (I1013170,I417669);
nor I_59387 (I1013187,I1013170,I417657);
not I_59388 (I1013204,I417666);
nor I_59389 (I1013221,I1013187,I417651);
nor I_59390 (I1013238,I1013145,I1013221);
DFFARX1 I_59391 (I1013238,I3563,I1013102,I1013088,);
nor I_59392 (I1013269,I417651,I417657);
nand I_59393 (I1013286,I1013269,I417669);
DFFARX1 I_59394 (I1013286,I3563,I1013102,I1013091,);
nor I_59395 (I1013317,I1013204,I417651);
nand I_59396 (I1013334,I1013317,I417642);
nor I_59397 (I1013351,I1013128,I1013334);
DFFARX1 I_59398 (I1013351,I3563,I1013102,I1013067,);
not I_59399 (I1013382,I1013334);
nand I_59400 (I1013079,I1013145,I1013382);
DFFARX1 I_59401 (I1013334,I3563,I1013102,I1013422,);
not I_59402 (I1013430,I1013422);
not I_59403 (I1013447,I417651);
not I_59404 (I1013464,I417654);
nor I_59405 (I1013481,I1013464,I417666);
nor I_59406 (I1013094,I1013430,I1013481);
nor I_59407 (I1013512,I1013464,I417663);
and I_59408 (I1013529,I1013512,I417645);
or I_59409 (I1013546,I1013529,I417660);
DFFARX1 I_59410 (I1013546,I3563,I1013102,I1013572,);
nor I_59411 (I1013082,I1013572,I1013128);
not I_59412 (I1013594,I1013572);
and I_59413 (I1013611,I1013594,I1013128);
nor I_59414 (I1013076,I1013153,I1013611);
nand I_59415 (I1013642,I1013594,I1013204);
nor I_59416 (I1013070,I1013464,I1013642);
nand I_59417 (I1013073,I1013594,I1013382);
nand I_59418 (I1013687,I1013204,I417654);
nor I_59419 (I1013085,I1013447,I1013687);
not I_59420 (I1013748,I3570);
DFFARX1 I_59421 (I343862,I3563,I1013748,I1013774,);
DFFARX1 I_59422 (I343868,I3563,I1013748,I1013791,);
not I_59423 (I1013799,I1013791);
not I_59424 (I1013816,I343889);
nor I_59425 (I1013833,I1013816,I343877);
not I_59426 (I1013850,I343886);
nor I_59427 (I1013867,I1013833,I343871);
nor I_59428 (I1013884,I1013791,I1013867);
DFFARX1 I_59429 (I1013884,I3563,I1013748,I1013734,);
nor I_59430 (I1013915,I343871,I343877);
nand I_59431 (I1013932,I1013915,I343889);
DFFARX1 I_59432 (I1013932,I3563,I1013748,I1013737,);
nor I_59433 (I1013963,I1013850,I343871);
nand I_59434 (I1013980,I1013963,I343862);
nor I_59435 (I1013997,I1013774,I1013980);
DFFARX1 I_59436 (I1013997,I3563,I1013748,I1013713,);
not I_59437 (I1014028,I1013980);
nand I_59438 (I1013725,I1013791,I1014028);
DFFARX1 I_59439 (I1013980,I3563,I1013748,I1014068,);
not I_59440 (I1014076,I1014068);
not I_59441 (I1014093,I343871);
not I_59442 (I1014110,I343874);
nor I_59443 (I1014127,I1014110,I343886);
nor I_59444 (I1013740,I1014076,I1014127);
nor I_59445 (I1014158,I1014110,I343883);
and I_59446 (I1014175,I1014158,I343865);
or I_59447 (I1014192,I1014175,I343880);
DFFARX1 I_59448 (I1014192,I3563,I1013748,I1014218,);
nor I_59449 (I1013728,I1014218,I1013774);
not I_59450 (I1014240,I1014218);
and I_59451 (I1014257,I1014240,I1013774);
nor I_59452 (I1013722,I1013799,I1014257);
nand I_59453 (I1014288,I1014240,I1013850);
nor I_59454 (I1013716,I1014110,I1014288);
nand I_59455 (I1013719,I1014240,I1014028);
nand I_59456 (I1014333,I1013850,I343874);
nor I_59457 (I1013731,I1014093,I1014333);
not I_59458 (I1014394,I3570);
DFFARX1 I_59459 (I415534,I3563,I1014394,I1014420,);
DFFARX1 I_59460 (I415540,I3563,I1014394,I1014437,);
not I_59461 (I1014445,I1014437);
not I_59462 (I1014462,I415561);
nor I_59463 (I1014479,I1014462,I415549);
not I_59464 (I1014496,I415558);
nor I_59465 (I1014513,I1014479,I415543);
nor I_59466 (I1014530,I1014437,I1014513);
DFFARX1 I_59467 (I1014530,I3563,I1014394,I1014380,);
nor I_59468 (I1014561,I415543,I415549);
nand I_59469 (I1014578,I1014561,I415561);
DFFARX1 I_59470 (I1014578,I3563,I1014394,I1014383,);
nor I_59471 (I1014609,I1014496,I415543);
nand I_59472 (I1014626,I1014609,I415534);
nor I_59473 (I1014643,I1014420,I1014626);
DFFARX1 I_59474 (I1014643,I3563,I1014394,I1014359,);
not I_59475 (I1014674,I1014626);
nand I_59476 (I1014371,I1014437,I1014674);
DFFARX1 I_59477 (I1014626,I3563,I1014394,I1014714,);
not I_59478 (I1014722,I1014714);
not I_59479 (I1014739,I415543);
not I_59480 (I1014756,I415546);
nor I_59481 (I1014773,I1014756,I415558);
nor I_59482 (I1014386,I1014722,I1014773);
nor I_59483 (I1014804,I1014756,I415555);
and I_59484 (I1014821,I1014804,I415537);
or I_59485 (I1014838,I1014821,I415552);
DFFARX1 I_59486 (I1014838,I3563,I1014394,I1014864,);
nor I_59487 (I1014374,I1014864,I1014420);
not I_59488 (I1014886,I1014864);
and I_59489 (I1014903,I1014886,I1014420);
nor I_59490 (I1014368,I1014445,I1014903);
nand I_59491 (I1014934,I1014886,I1014496);
nor I_59492 (I1014362,I1014756,I1014934);
nand I_59493 (I1014365,I1014886,I1014674);
nand I_59494 (I1014979,I1014496,I415546);
nor I_59495 (I1014377,I1014739,I1014979);
not I_59496 (I1015040,I3570);
DFFARX1 I_59497 (I1229155,I3563,I1015040,I1015066,);
DFFARX1 I_59498 (I1229137,I3563,I1015040,I1015083,);
not I_59499 (I1015091,I1015083);
not I_59500 (I1015108,I1229146);
nor I_59501 (I1015125,I1015108,I1229158);
not I_59502 (I1015142,I1229140);
nor I_59503 (I1015159,I1015125,I1229149);
nor I_59504 (I1015176,I1015083,I1015159);
DFFARX1 I_59505 (I1015176,I3563,I1015040,I1015026,);
nor I_59506 (I1015207,I1229149,I1229158);
nand I_59507 (I1015224,I1015207,I1229146);
DFFARX1 I_59508 (I1015224,I3563,I1015040,I1015029,);
nor I_59509 (I1015255,I1015142,I1229149);
nand I_59510 (I1015272,I1015255,I1229161);
nor I_59511 (I1015289,I1015066,I1015272);
DFFARX1 I_59512 (I1015289,I3563,I1015040,I1015005,);
not I_59513 (I1015320,I1015272);
nand I_59514 (I1015017,I1015083,I1015320);
DFFARX1 I_59515 (I1015272,I3563,I1015040,I1015360,);
not I_59516 (I1015368,I1015360);
not I_59517 (I1015385,I1229149);
not I_59518 (I1015402,I1229137);
nor I_59519 (I1015419,I1015402,I1229140);
nor I_59520 (I1015032,I1015368,I1015419);
nor I_59521 (I1015450,I1015402,I1229143);
and I_59522 (I1015467,I1015450,I1229152);
or I_59523 (I1015484,I1015467,I1229140);
DFFARX1 I_59524 (I1015484,I3563,I1015040,I1015510,);
nor I_59525 (I1015020,I1015510,I1015066);
not I_59526 (I1015532,I1015510);
and I_59527 (I1015549,I1015532,I1015066);
nor I_59528 (I1015014,I1015091,I1015549);
nand I_59529 (I1015580,I1015532,I1015142);
nor I_59530 (I1015008,I1015402,I1015580);
nand I_59531 (I1015011,I1015532,I1015320);
nand I_59532 (I1015625,I1015142,I1229137);
nor I_59533 (I1015023,I1015385,I1015625);
not I_59534 (I1015686,I3570);
DFFARX1 I_59535 (I367577,I3563,I1015686,I1015712,);
DFFARX1 I_59536 (I367583,I3563,I1015686,I1015729,);
not I_59537 (I1015737,I1015729);
not I_59538 (I1015754,I367604);
nor I_59539 (I1015771,I1015754,I367592);
not I_59540 (I1015788,I367601);
nor I_59541 (I1015805,I1015771,I367586);
nor I_59542 (I1015822,I1015729,I1015805);
DFFARX1 I_59543 (I1015822,I3563,I1015686,I1015672,);
nor I_59544 (I1015853,I367586,I367592);
nand I_59545 (I1015870,I1015853,I367604);
DFFARX1 I_59546 (I1015870,I3563,I1015686,I1015675,);
nor I_59547 (I1015901,I1015788,I367586);
nand I_59548 (I1015918,I1015901,I367577);
nor I_59549 (I1015935,I1015712,I1015918);
DFFARX1 I_59550 (I1015935,I3563,I1015686,I1015651,);
not I_59551 (I1015966,I1015918);
nand I_59552 (I1015663,I1015729,I1015966);
DFFARX1 I_59553 (I1015918,I3563,I1015686,I1016006,);
not I_59554 (I1016014,I1016006);
not I_59555 (I1016031,I367586);
not I_59556 (I1016048,I367589);
nor I_59557 (I1016065,I1016048,I367601);
nor I_59558 (I1015678,I1016014,I1016065);
nor I_59559 (I1016096,I1016048,I367598);
and I_59560 (I1016113,I1016096,I367580);
or I_59561 (I1016130,I1016113,I367595);
DFFARX1 I_59562 (I1016130,I3563,I1015686,I1016156,);
nor I_59563 (I1015666,I1016156,I1015712);
not I_59564 (I1016178,I1016156);
and I_59565 (I1016195,I1016178,I1015712);
nor I_59566 (I1015660,I1015737,I1016195);
nand I_59567 (I1016226,I1016178,I1015788);
nor I_59568 (I1015654,I1016048,I1016226);
nand I_59569 (I1015657,I1016178,I1015966);
nand I_59570 (I1016271,I1015788,I367589);
nor I_59571 (I1015669,I1016031,I1016271);
not I_59572 (I1016332,I3570);
DFFARX1 I_59573 (I94064,I3563,I1016332,I1016358,);
DFFARX1 I_59574 (I94070,I3563,I1016332,I1016375,);
not I_59575 (I1016383,I1016375);
not I_59576 (I1016400,I94088);
nor I_59577 (I1016417,I1016400,I94067);
not I_59578 (I1016434,I94073);
nor I_59579 (I1016451,I1016417,I94079);
nor I_59580 (I1016468,I1016375,I1016451);
DFFARX1 I_59581 (I1016468,I3563,I1016332,I1016318,);
nor I_59582 (I1016499,I94079,I94067);
nand I_59583 (I1016516,I1016499,I94088);
DFFARX1 I_59584 (I1016516,I3563,I1016332,I1016321,);
nor I_59585 (I1016547,I1016434,I94079);
nand I_59586 (I1016564,I1016547,I94085);
nor I_59587 (I1016581,I1016358,I1016564);
DFFARX1 I_59588 (I1016581,I3563,I1016332,I1016297,);
not I_59589 (I1016612,I1016564);
nand I_59590 (I1016309,I1016375,I1016612);
DFFARX1 I_59591 (I1016564,I3563,I1016332,I1016652,);
not I_59592 (I1016660,I1016652);
not I_59593 (I1016677,I94079);
not I_59594 (I1016694,I94067);
nor I_59595 (I1016711,I1016694,I94073);
nor I_59596 (I1016324,I1016660,I1016711);
nor I_59597 (I1016742,I1016694,I94076);
and I_59598 (I1016759,I1016742,I94064);
or I_59599 (I1016776,I1016759,I94082);
DFFARX1 I_59600 (I1016776,I3563,I1016332,I1016802,);
nor I_59601 (I1016312,I1016802,I1016358);
not I_59602 (I1016824,I1016802);
and I_59603 (I1016841,I1016824,I1016358);
nor I_59604 (I1016306,I1016383,I1016841);
nand I_59605 (I1016872,I1016824,I1016434);
nor I_59606 (I1016300,I1016694,I1016872);
nand I_59607 (I1016303,I1016824,I1016612);
nand I_59608 (I1016917,I1016434,I94067);
nor I_59609 (I1016315,I1016677,I1016917);
not I_59610 (I1016978,I3570);
DFFARX1 I_59611 (I626048,I3563,I1016978,I1017004,);
DFFARX1 I_59612 (I626060,I3563,I1016978,I1017021,);
not I_59613 (I1017029,I1017021);
not I_59614 (I1017046,I626069);
nor I_59615 (I1017063,I1017046,I626045);
not I_59616 (I1017080,I626063);
nor I_59617 (I1017097,I1017063,I626057);
nor I_59618 (I1017114,I1017021,I1017097);
DFFARX1 I_59619 (I1017114,I3563,I1016978,I1016964,);
nor I_59620 (I1017145,I626057,I626045);
nand I_59621 (I1017162,I1017145,I626069);
DFFARX1 I_59622 (I1017162,I3563,I1016978,I1016967,);
nor I_59623 (I1017193,I1017080,I626057);
nand I_59624 (I1017210,I1017193,I626051);
nor I_59625 (I1017227,I1017004,I1017210);
DFFARX1 I_59626 (I1017227,I3563,I1016978,I1016943,);
not I_59627 (I1017258,I1017210);
nand I_59628 (I1016955,I1017021,I1017258);
DFFARX1 I_59629 (I1017210,I3563,I1016978,I1017298,);
not I_59630 (I1017306,I1017298);
not I_59631 (I1017323,I626057);
not I_59632 (I1017340,I626066);
nor I_59633 (I1017357,I1017340,I626063);
nor I_59634 (I1016970,I1017306,I1017357);
nor I_59635 (I1017388,I1017340,I626048);
and I_59636 (I1017405,I1017388,I626045);
or I_59637 (I1017422,I1017405,I626054);
DFFARX1 I_59638 (I1017422,I3563,I1016978,I1017448,);
nor I_59639 (I1016958,I1017448,I1017004);
not I_59640 (I1017470,I1017448);
and I_59641 (I1017487,I1017470,I1017004);
nor I_59642 (I1016952,I1017029,I1017487);
nand I_59643 (I1017518,I1017470,I1017080);
nor I_59644 (I1016946,I1017340,I1017518);
nand I_59645 (I1016949,I1017470,I1017258);
nand I_59646 (I1017563,I1017080,I626066);
nor I_59647 (I1016961,I1017323,I1017563);
not I_59648 (I1017624,I3570);
DFFARX1 I_59649 (I1147079,I3563,I1017624,I1017650,);
DFFARX1 I_59650 (I1147061,I3563,I1017624,I1017667,);
not I_59651 (I1017675,I1017667);
not I_59652 (I1017692,I1147070);
nor I_59653 (I1017709,I1017692,I1147082);
not I_59654 (I1017726,I1147064);
nor I_59655 (I1017743,I1017709,I1147073);
nor I_59656 (I1017760,I1017667,I1017743);
DFFARX1 I_59657 (I1017760,I3563,I1017624,I1017610,);
nor I_59658 (I1017791,I1147073,I1147082);
nand I_59659 (I1017808,I1017791,I1147070);
DFFARX1 I_59660 (I1017808,I3563,I1017624,I1017613,);
nor I_59661 (I1017839,I1017726,I1147073);
nand I_59662 (I1017856,I1017839,I1147085);
nor I_59663 (I1017873,I1017650,I1017856);
DFFARX1 I_59664 (I1017873,I3563,I1017624,I1017589,);
not I_59665 (I1017904,I1017856);
nand I_59666 (I1017601,I1017667,I1017904);
DFFARX1 I_59667 (I1017856,I3563,I1017624,I1017944,);
not I_59668 (I1017952,I1017944);
not I_59669 (I1017969,I1147073);
not I_59670 (I1017986,I1147061);
nor I_59671 (I1018003,I1017986,I1147064);
nor I_59672 (I1017616,I1017952,I1018003);
nor I_59673 (I1018034,I1017986,I1147067);
and I_59674 (I1018051,I1018034,I1147076);
or I_59675 (I1018068,I1018051,I1147064);
DFFARX1 I_59676 (I1018068,I3563,I1017624,I1018094,);
nor I_59677 (I1017604,I1018094,I1017650);
not I_59678 (I1018116,I1018094);
and I_59679 (I1018133,I1018116,I1017650);
nor I_59680 (I1017598,I1017675,I1018133);
nand I_59681 (I1018164,I1018116,I1017726);
nor I_59682 (I1017592,I1017986,I1018164);
nand I_59683 (I1017595,I1018116,I1017904);
nand I_59684 (I1018209,I1017726,I1147061);
nor I_59685 (I1017607,I1017969,I1018209);
not I_59686 (I1018270,I3570);
DFFARX1 I_59687 (I900125,I3563,I1018270,I1018296,);
DFFARX1 I_59688 (I900122,I3563,I1018270,I1018313,);
not I_59689 (I1018321,I1018313);
not I_59690 (I1018338,I900122);
nor I_59691 (I1018355,I1018338,I900125);
not I_59692 (I1018372,I900137);
nor I_59693 (I1018389,I1018355,I900131);
nor I_59694 (I1018406,I1018313,I1018389);
DFFARX1 I_59695 (I1018406,I3563,I1018270,I1018256,);
nor I_59696 (I1018437,I900131,I900125);
nand I_59697 (I1018454,I1018437,I900122);
DFFARX1 I_59698 (I1018454,I3563,I1018270,I1018259,);
nor I_59699 (I1018485,I1018372,I900131);
nand I_59700 (I1018502,I1018485,I900119);
nor I_59701 (I1018519,I1018296,I1018502);
DFFARX1 I_59702 (I1018519,I3563,I1018270,I1018235,);
not I_59703 (I1018550,I1018502);
nand I_59704 (I1018247,I1018313,I1018550);
DFFARX1 I_59705 (I1018502,I3563,I1018270,I1018590,);
not I_59706 (I1018598,I1018590);
not I_59707 (I1018615,I900131);
not I_59708 (I1018632,I900128);
nor I_59709 (I1018649,I1018632,I900137);
nor I_59710 (I1018262,I1018598,I1018649);
nor I_59711 (I1018680,I1018632,I900134);
and I_59712 (I1018697,I1018680,I900140);
or I_59713 (I1018714,I1018697,I900119);
DFFARX1 I_59714 (I1018714,I3563,I1018270,I1018740,);
nor I_59715 (I1018250,I1018740,I1018296);
not I_59716 (I1018762,I1018740);
and I_59717 (I1018779,I1018762,I1018296);
nor I_59718 (I1018244,I1018321,I1018779);
nand I_59719 (I1018810,I1018762,I1018372);
nor I_59720 (I1018238,I1018632,I1018810);
nand I_59721 (I1018241,I1018762,I1018550);
nand I_59722 (I1018855,I1018372,I900128);
nor I_59723 (I1018253,I1018615,I1018855);
not I_59724 (I1018916,I3570);
DFFARX1 I_59725 (I75619,I3563,I1018916,I1018942,);
DFFARX1 I_59726 (I75625,I3563,I1018916,I1018959,);
not I_59727 (I1018967,I1018959);
not I_59728 (I1018984,I75643);
nor I_59729 (I1019001,I1018984,I75622);
not I_59730 (I1019018,I75628);
nor I_59731 (I1019035,I1019001,I75634);
nor I_59732 (I1019052,I1018959,I1019035);
DFFARX1 I_59733 (I1019052,I3563,I1018916,I1018902,);
nor I_59734 (I1019083,I75634,I75622);
nand I_59735 (I1019100,I1019083,I75643);
DFFARX1 I_59736 (I1019100,I3563,I1018916,I1018905,);
nor I_59737 (I1019131,I1019018,I75634);
nand I_59738 (I1019148,I1019131,I75640);
nor I_59739 (I1019165,I1018942,I1019148);
DFFARX1 I_59740 (I1019165,I3563,I1018916,I1018881,);
not I_59741 (I1019196,I1019148);
nand I_59742 (I1018893,I1018959,I1019196);
DFFARX1 I_59743 (I1019148,I3563,I1018916,I1019236,);
not I_59744 (I1019244,I1019236);
not I_59745 (I1019261,I75634);
not I_59746 (I1019278,I75622);
nor I_59747 (I1019295,I1019278,I75628);
nor I_59748 (I1018908,I1019244,I1019295);
nor I_59749 (I1019326,I1019278,I75631);
and I_59750 (I1019343,I1019326,I75619);
or I_59751 (I1019360,I1019343,I75637);
DFFARX1 I_59752 (I1019360,I3563,I1018916,I1019386,);
nor I_59753 (I1018896,I1019386,I1018942);
not I_59754 (I1019408,I1019386);
and I_59755 (I1019425,I1019408,I1018942);
nor I_59756 (I1018890,I1018967,I1019425);
nand I_59757 (I1019456,I1019408,I1019018);
nor I_59758 (I1018884,I1019278,I1019456);
nand I_59759 (I1018887,I1019408,I1019196);
nand I_59760 (I1019501,I1019018,I75622);
nor I_59761 (I1018899,I1019261,I1019501);
not I_59762 (I1019562,I3570);
DFFARX1 I_59763 (I281529,I3563,I1019562,I1019588,);
DFFARX1 I_59764 (I281541,I3563,I1019562,I1019605,);
not I_59765 (I1019613,I1019605);
not I_59766 (I1019630,I281547);
nor I_59767 (I1019647,I1019630,I281532);
not I_59768 (I1019664,I281523);
nor I_59769 (I1019681,I1019647,I281544);
nor I_59770 (I1019698,I1019605,I1019681);
DFFARX1 I_59771 (I1019698,I3563,I1019562,I1019548,);
nor I_59772 (I1019729,I281544,I281532);
nand I_59773 (I1019746,I1019729,I281547);
DFFARX1 I_59774 (I1019746,I3563,I1019562,I1019551,);
nor I_59775 (I1019777,I1019664,I281544);
nand I_59776 (I1019794,I1019777,I281526);
nor I_59777 (I1019811,I1019588,I1019794);
DFFARX1 I_59778 (I1019811,I3563,I1019562,I1019527,);
not I_59779 (I1019842,I1019794);
nand I_59780 (I1019539,I1019605,I1019842);
DFFARX1 I_59781 (I1019794,I3563,I1019562,I1019882,);
not I_59782 (I1019890,I1019882);
not I_59783 (I1019907,I281544);
not I_59784 (I1019924,I281535);
nor I_59785 (I1019941,I1019924,I281523);
nor I_59786 (I1019554,I1019890,I1019941);
nor I_59787 (I1019972,I1019924,I281538);
and I_59788 (I1019989,I1019972,I281526);
or I_59789 (I1020006,I1019989,I281523);
DFFARX1 I_59790 (I1020006,I3563,I1019562,I1020032,);
nor I_59791 (I1019542,I1020032,I1019588);
not I_59792 (I1020054,I1020032);
and I_59793 (I1020071,I1020054,I1019588);
nor I_59794 (I1019536,I1019613,I1020071);
nand I_59795 (I1020102,I1020054,I1019664);
nor I_59796 (I1019530,I1019924,I1020102);
nand I_59797 (I1019533,I1020054,I1019842);
nand I_59798 (I1020147,I1019664,I281535);
nor I_59799 (I1019545,I1019907,I1020147);
not I_59800 (I1020208,I3570);
DFFARX1 I_59801 (I1217595,I3563,I1020208,I1020234,);
DFFARX1 I_59802 (I1217577,I3563,I1020208,I1020251,);
not I_59803 (I1020259,I1020251);
not I_59804 (I1020276,I1217586);
nor I_59805 (I1020293,I1020276,I1217598);
not I_59806 (I1020310,I1217580);
nor I_59807 (I1020327,I1020293,I1217589);
nor I_59808 (I1020344,I1020251,I1020327);
DFFARX1 I_59809 (I1020344,I3563,I1020208,I1020194,);
nor I_59810 (I1020375,I1217589,I1217598);
nand I_59811 (I1020392,I1020375,I1217586);
DFFARX1 I_59812 (I1020392,I3563,I1020208,I1020197,);
nor I_59813 (I1020423,I1020310,I1217589);
nand I_59814 (I1020440,I1020423,I1217601);
nor I_59815 (I1020457,I1020234,I1020440);
DFFARX1 I_59816 (I1020457,I3563,I1020208,I1020173,);
not I_59817 (I1020488,I1020440);
nand I_59818 (I1020185,I1020251,I1020488);
DFFARX1 I_59819 (I1020440,I3563,I1020208,I1020528,);
not I_59820 (I1020536,I1020528);
not I_59821 (I1020553,I1217589);
not I_59822 (I1020570,I1217577);
nor I_59823 (I1020587,I1020570,I1217580);
nor I_59824 (I1020200,I1020536,I1020587);
nor I_59825 (I1020618,I1020570,I1217583);
and I_59826 (I1020635,I1020618,I1217592);
or I_59827 (I1020652,I1020635,I1217580);
DFFARX1 I_59828 (I1020652,I3563,I1020208,I1020678,);
nor I_59829 (I1020188,I1020678,I1020234);
not I_59830 (I1020700,I1020678);
and I_59831 (I1020717,I1020700,I1020234);
nor I_59832 (I1020182,I1020259,I1020717);
nand I_59833 (I1020748,I1020700,I1020310);
nor I_59834 (I1020176,I1020570,I1020748);
nand I_59835 (I1020179,I1020700,I1020488);
nand I_59836 (I1020793,I1020310,I1217577);
nor I_59837 (I1020191,I1020553,I1020793);
not I_59838 (I1020854,I3570);
DFFARX1 I_59839 (I404467,I3563,I1020854,I1020880,);
DFFARX1 I_59840 (I404473,I3563,I1020854,I1020897,);
not I_59841 (I1020905,I1020897);
not I_59842 (I1020922,I404494);
nor I_59843 (I1020939,I1020922,I404482);
not I_59844 (I1020956,I404491);
nor I_59845 (I1020973,I1020939,I404476);
nor I_59846 (I1020990,I1020897,I1020973);
DFFARX1 I_59847 (I1020990,I3563,I1020854,I1020840,);
nor I_59848 (I1021021,I404476,I404482);
nand I_59849 (I1021038,I1021021,I404494);
DFFARX1 I_59850 (I1021038,I3563,I1020854,I1020843,);
nor I_59851 (I1021069,I1020956,I404476);
nand I_59852 (I1021086,I1021069,I404467);
nor I_59853 (I1021103,I1020880,I1021086);
DFFARX1 I_59854 (I1021103,I3563,I1020854,I1020819,);
not I_59855 (I1021134,I1021086);
nand I_59856 (I1020831,I1020897,I1021134);
DFFARX1 I_59857 (I1021086,I3563,I1020854,I1021174,);
not I_59858 (I1021182,I1021174);
not I_59859 (I1021199,I404476);
not I_59860 (I1021216,I404479);
nor I_59861 (I1021233,I1021216,I404491);
nor I_59862 (I1020846,I1021182,I1021233);
nor I_59863 (I1021264,I1021216,I404488);
and I_59864 (I1021281,I1021264,I404470);
or I_59865 (I1021298,I1021281,I404485);
DFFARX1 I_59866 (I1021298,I3563,I1020854,I1021324,);
nor I_59867 (I1020834,I1021324,I1020880);
not I_59868 (I1021346,I1021324);
and I_59869 (I1021363,I1021346,I1020880);
nor I_59870 (I1020828,I1020905,I1021363);
nand I_59871 (I1021394,I1021346,I1020956);
nor I_59872 (I1020822,I1021216,I1021394);
nand I_59873 (I1020825,I1021346,I1021134);
nand I_59874 (I1021439,I1020956,I404479);
nor I_59875 (I1020837,I1021199,I1021439);
not I_59876 (I1021500,I3570);
DFFARX1 I_59877 (I1061245,I3563,I1021500,I1021526,);
DFFARX1 I_59878 (I1061248,I3563,I1021500,I1021543,);
not I_59879 (I1021551,I1021543);
not I_59880 (I1021568,I1061245);
nor I_59881 (I1021585,I1021568,I1061257);
not I_59882 (I1021602,I1061266);
nor I_59883 (I1021619,I1021585,I1061254);
nor I_59884 (I1021636,I1021543,I1021619);
DFFARX1 I_59885 (I1021636,I3563,I1021500,I1021486,);
nor I_59886 (I1021667,I1061254,I1061257);
nand I_59887 (I1021684,I1021667,I1061245);
DFFARX1 I_59888 (I1021684,I3563,I1021500,I1021489,);
nor I_59889 (I1021715,I1021602,I1061254);
nand I_59890 (I1021732,I1021715,I1061260);
nor I_59891 (I1021749,I1021526,I1021732);
DFFARX1 I_59892 (I1021749,I3563,I1021500,I1021465,);
not I_59893 (I1021780,I1021732);
nand I_59894 (I1021477,I1021543,I1021780);
DFFARX1 I_59895 (I1021732,I3563,I1021500,I1021820,);
not I_59896 (I1021828,I1021820);
not I_59897 (I1021845,I1061254);
not I_59898 (I1021862,I1061251);
nor I_59899 (I1021879,I1021862,I1061266);
nor I_59900 (I1021492,I1021828,I1021879);
nor I_59901 (I1021910,I1021862,I1061263);
and I_59902 (I1021927,I1021910,I1061251);
or I_59903 (I1021944,I1021927,I1061248);
DFFARX1 I_59904 (I1021944,I3563,I1021500,I1021970,);
nor I_59905 (I1021480,I1021970,I1021526);
not I_59906 (I1021992,I1021970);
and I_59907 (I1022009,I1021992,I1021526);
nor I_59908 (I1021474,I1021551,I1022009);
nand I_59909 (I1022040,I1021992,I1021602);
nor I_59910 (I1021468,I1021862,I1022040);
nand I_59911 (I1021471,I1021992,I1021780);
nand I_59912 (I1022085,I1021602,I1061251);
nor I_59913 (I1021483,I1021845,I1022085);
not I_59914 (I1022146,I3570);
DFFARX1 I_59915 (I1114133,I3563,I1022146,I1022172,);
DFFARX1 I_59916 (I1114115,I3563,I1022146,I1022189,);
not I_59917 (I1022197,I1022189);
not I_59918 (I1022214,I1114124);
nor I_59919 (I1022231,I1022214,I1114136);
not I_59920 (I1022248,I1114118);
nor I_59921 (I1022265,I1022231,I1114127);
nor I_59922 (I1022282,I1022189,I1022265);
DFFARX1 I_59923 (I1022282,I3563,I1022146,I1022132,);
nor I_59924 (I1022313,I1114127,I1114136);
nand I_59925 (I1022330,I1022313,I1114124);
DFFARX1 I_59926 (I1022330,I3563,I1022146,I1022135,);
nor I_59927 (I1022361,I1022248,I1114127);
nand I_59928 (I1022378,I1022361,I1114139);
nor I_59929 (I1022395,I1022172,I1022378);
DFFARX1 I_59930 (I1022395,I3563,I1022146,I1022111,);
not I_59931 (I1022426,I1022378);
nand I_59932 (I1022123,I1022189,I1022426);
DFFARX1 I_59933 (I1022378,I3563,I1022146,I1022466,);
not I_59934 (I1022474,I1022466);
not I_59935 (I1022491,I1114127);
not I_59936 (I1022508,I1114115);
nor I_59937 (I1022525,I1022508,I1114118);
nor I_59938 (I1022138,I1022474,I1022525);
nor I_59939 (I1022556,I1022508,I1114121);
and I_59940 (I1022573,I1022556,I1114130);
or I_59941 (I1022590,I1022573,I1114118);
DFFARX1 I_59942 (I1022590,I3563,I1022146,I1022616,);
nor I_59943 (I1022126,I1022616,I1022172);
not I_59944 (I1022638,I1022616);
and I_59945 (I1022655,I1022638,I1022172);
nor I_59946 (I1022120,I1022197,I1022655);
nand I_59947 (I1022686,I1022638,I1022248);
nor I_59948 (I1022114,I1022508,I1022686);
nand I_59949 (I1022117,I1022638,I1022426);
nand I_59950 (I1022731,I1022248,I1114115);
nor I_59951 (I1022129,I1022491,I1022731);
not I_59952 (I1022792,I3570);
DFFARX1 I_59953 (I463752,I3563,I1022792,I1022818,);
DFFARX1 I_59954 (I463749,I3563,I1022792,I1022835,);
not I_59955 (I1022843,I1022835);
not I_59956 (I1022860,I463764);
nor I_59957 (I1022877,I1022860,I463767);
not I_59958 (I1022894,I463755);
nor I_59959 (I1022911,I1022877,I463761);
nor I_59960 (I1022928,I1022835,I1022911);
DFFARX1 I_59961 (I1022928,I3563,I1022792,I1022778,);
nor I_59962 (I1022959,I463761,I463767);
nand I_59963 (I1022976,I1022959,I463764);
DFFARX1 I_59964 (I1022976,I3563,I1022792,I1022781,);
nor I_59965 (I1023007,I1022894,I463761);
nand I_59966 (I1023024,I1023007,I463773);
nor I_59967 (I1023041,I1022818,I1023024);
DFFARX1 I_59968 (I1023041,I3563,I1022792,I1022757,);
not I_59969 (I1023072,I1023024);
nand I_59970 (I1022769,I1022835,I1023072);
DFFARX1 I_59971 (I1023024,I3563,I1022792,I1023112,);
not I_59972 (I1023120,I1023112);
not I_59973 (I1023137,I463761);
not I_59974 (I1023154,I463746);
nor I_59975 (I1023171,I1023154,I463755);
nor I_59976 (I1022784,I1023120,I1023171);
nor I_59977 (I1023202,I1023154,I463758);
and I_59978 (I1023219,I1023202,I463746);
or I_59979 (I1023236,I1023219,I463770);
DFFARX1 I_59980 (I1023236,I3563,I1022792,I1023262,);
nor I_59981 (I1022772,I1023262,I1022818);
not I_59982 (I1023284,I1023262);
and I_59983 (I1023301,I1023284,I1022818);
nor I_59984 (I1022766,I1022843,I1023301);
nand I_59985 (I1023332,I1023284,I1022894);
nor I_59986 (I1022760,I1023154,I1023332);
nand I_59987 (I1022763,I1023284,I1023072);
nand I_59988 (I1023377,I1022894,I463746);
nor I_59989 (I1022775,I1023137,I1023377);
not I_59990 (I1023438,I3570);
DFFARX1 I_59991 (I120414,I3563,I1023438,I1023464,);
DFFARX1 I_59992 (I120420,I3563,I1023438,I1023481,);
not I_59993 (I1023489,I1023481);
not I_59994 (I1023506,I120438);
nor I_59995 (I1023523,I1023506,I120417);
not I_59996 (I1023540,I120423);
nor I_59997 (I1023557,I1023523,I120429);
nor I_59998 (I1023574,I1023481,I1023557);
DFFARX1 I_59999 (I1023574,I3563,I1023438,I1023424,);
nor I_60000 (I1023605,I120429,I120417);
nand I_60001 (I1023622,I1023605,I120438);
DFFARX1 I_60002 (I1023622,I3563,I1023438,I1023427,);
nor I_60003 (I1023653,I1023540,I120429);
nand I_60004 (I1023670,I1023653,I120435);
nor I_60005 (I1023687,I1023464,I1023670);
DFFARX1 I_60006 (I1023687,I3563,I1023438,I1023403,);
not I_60007 (I1023718,I1023670);
nand I_60008 (I1023415,I1023481,I1023718);
DFFARX1 I_60009 (I1023670,I3563,I1023438,I1023758,);
not I_60010 (I1023766,I1023758);
not I_60011 (I1023783,I120429);
not I_60012 (I1023800,I120417);
nor I_60013 (I1023817,I1023800,I120423);
nor I_60014 (I1023430,I1023766,I1023817);
nor I_60015 (I1023848,I1023800,I120426);
and I_60016 (I1023865,I1023848,I120414);
or I_60017 (I1023882,I1023865,I120432);
DFFARX1 I_60018 (I1023882,I3563,I1023438,I1023908,);
nor I_60019 (I1023418,I1023908,I1023464);
not I_60020 (I1023930,I1023908);
and I_60021 (I1023947,I1023930,I1023464);
nor I_60022 (I1023412,I1023489,I1023947);
nand I_60023 (I1023978,I1023930,I1023540);
nor I_60024 (I1023406,I1023800,I1023978);
nand I_60025 (I1023409,I1023930,I1023718);
nand I_60026 (I1024023,I1023540,I120417);
nor I_60027 (I1023421,I1023783,I1024023);
not I_60028 (I1024084,I3570);
DFFARX1 I_60029 (I686741,I3563,I1024084,I1024110,);
DFFARX1 I_60030 (I686735,I3563,I1024084,I1024127,);
not I_60031 (I1024135,I1024127);
not I_60032 (I1024152,I686750);
nor I_60033 (I1024169,I1024152,I686735);
not I_60034 (I1024186,I686744);
nor I_60035 (I1024203,I1024169,I686753);
nor I_60036 (I1024220,I1024127,I1024203);
DFFARX1 I_60037 (I1024220,I3563,I1024084,I1024070,);
nor I_60038 (I1024251,I686753,I686735);
nand I_60039 (I1024268,I1024251,I686750);
DFFARX1 I_60040 (I1024268,I3563,I1024084,I1024073,);
nor I_60041 (I1024299,I1024186,I686753);
nand I_60042 (I1024316,I1024299,I686738);
nor I_60043 (I1024333,I1024110,I1024316);
DFFARX1 I_60044 (I1024333,I3563,I1024084,I1024049,);
not I_60045 (I1024364,I1024316);
nand I_60046 (I1024061,I1024127,I1024364);
DFFARX1 I_60047 (I1024316,I3563,I1024084,I1024404,);
not I_60048 (I1024412,I1024404);
not I_60049 (I1024429,I686753);
not I_60050 (I1024446,I686747);
nor I_60051 (I1024463,I1024446,I686744);
nor I_60052 (I1024076,I1024412,I1024463);
nor I_60053 (I1024494,I1024446,I686756);
and I_60054 (I1024511,I1024494,I686759);
or I_60055 (I1024528,I1024511,I686738);
DFFARX1 I_60056 (I1024528,I3563,I1024084,I1024554,);
nor I_60057 (I1024064,I1024554,I1024110);
not I_60058 (I1024576,I1024554);
and I_60059 (I1024593,I1024576,I1024110);
nor I_60060 (I1024058,I1024135,I1024593);
nand I_60061 (I1024624,I1024576,I1024186);
nor I_60062 (I1024052,I1024446,I1024624);
nand I_60063 (I1024055,I1024576,I1024364);
nand I_60064 (I1024669,I1024186,I686747);
nor I_60065 (I1024067,I1024429,I1024669);
not I_60066 (I1024730,I3570);
DFFARX1 I_60067 (I170859,I3563,I1024730,I1024756,);
DFFARX1 I_60068 (I170871,I3563,I1024730,I1024773,);
not I_60069 (I1024781,I1024773);
not I_60070 (I1024798,I170877);
nor I_60071 (I1024815,I1024798,I170862);
not I_60072 (I1024832,I170853);
nor I_60073 (I1024849,I1024815,I170874);
nor I_60074 (I1024866,I1024773,I1024849);
DFFARX1 I_60075 (I1024866,I3563,I1024730,I1024716,);
nor I_60076 (I1024897,I170874,I170862);
nand I_60077 (I1024914,I1024897,I170877);
DFFARX1 I_60078 (I1024914,I3563,I1024730,I1024719,);
nor I_60079 (I1024945,I1024832,I170874);
nand I_60080 (I1024962,I1024945,I170856);
nor I_60081 (I1024979,I1024756,I1024962);
DFFARX1 I_60082 (I1024979,I3563,I1024730,I1024695,);
not I_60083 (I1025010,I1024962);
nand I_60084 (I1024707,I1024773,I1025010);
DFFARX1 I_60085 (I1024962,I3563,I1024730,I1025050,);
not I_60086 (I1025058,I1025050);
not I_60087 (I1025075,I170874);
not I_60088 (I1025092,I170865);
nor I_60089 (I1025109,I1025092,I170853);
nor I_60090 (I1024722,I1025058,I1025109);
nor I_60091 (I1025140,I1025092,I170868);
and I_60092 (I1025157,I1025140,I170856);
or I_60093 (I1025174,I1025157,I170853);
DFFARX1 I_60094 (I1025174,I3563,I1024730,I1025200,);
nor I_60095 (I1024710,I1025200,I1024756);
not I_60096 (I1025222,I1025200);
and I_60097 (I1025239,I1025222,I1024756);
nor I_60098 (I1024704,I1024781,I1025239);
nand I_60099 (I1025270,I1025222,I1024832);
nor I_60100 (I1024698,I1025092,I1025270);
nand I_60101 (I1024701,I1025222,I1025010);
nand I_60102 (I1025315,I1024832,I170865);
nor I_60103 (I1024713,I1025075,I1025315);
not I_60104 (I1025376,I3570);
DFFARX1 I_60105 (I8931,I3563,I1025376,I1025402,);
DFFARX1 I_60106 (I8928,I3563,I1025376,I1025419,);
not I_60107 (I1025427,I1025419);
not I_60108 (I1025444,I8940);
nor I_60109 (I1025461,I1025444,I8937);
not I_60110 (I1025478,I8946);
nor I_60111 (I1025495,I1025461,I8943);
nor I_60112 (I1025512,I1025419,I1025495);
DFFARX1 I_60113 (I1025512,I3563,I1025376,I1025362,);
nor I_60114 (I1025543,I8943,I8937);
nand I_60115 (I1025560,I1025543,I8940);
DFFARX1 I_60116 (I1025560,I3563,I1025376,I1025365,);
nor I_60117 (I1025591,I1025478,I8943);
nand I_60118 (I1025608,I1025591,I8934);
nor I_60119 (I1025625,I1025402,I1025608);
DFFARX1 I_60120 (I1025625,I3563,I1025376,I1025341,);
not I_60121 (I1025656,I1025608);
nand I_60122 (I1025353,I1025419,I1025656);
DFFARX1 I_60123 (I1025608,I3563,I1025376,I1025696,);
not I_60124 (I1025704,I1025696);
not I_60125 (I1025721,I8943);
not I_60126 (I1025738,I8934);
nor I_60127 (I1025755,I1025738,I8946);
nor I_60128 (I1025368,I1025704,I1025755);
nor I_60129 (I1025786,I1025738,I8928);
and I_60130 (I1025803,I1025786,I8949);
or I_60131 (I1025820,I1025803,I8931);
DFFARX1 I_60132 (I1025820,I3563,I1025376,I1025846,);
nor I_60133 (I1025356,I1025846,I1025402);
not I_60134 (I1025868,I1025846);
and I_60135 (I1025885,I1025868,I1025402);
nor I_60136 (I1025350,I1025427,I1025885);
nand I_60137 (I1025916,I1025868,I1025478);
nor I_60138 (I1025344,I1025738,I1025916);
nand I_60139 (I1025347,I1025868,I1025656);
nand I_60140 (I1025961,I1025478,I8934);
nor I_60141 (I1025359,I1025721,I1025961);
not I_60142 (I1026022,I3570);
DFFARX1 I_60143 (I264869,I3563,I1026022,I1026048,);
DFFARX1 I_60144 (I264881,I3563,I1026022,I1026065,);
not I_60145 (I1026073,I1026065);
not I_60146 (I1026090,I264887);
nor I_60147 (I1026107,I1026090,I264872);
not I_60148 (I1026124,I264863);
nor I_60149 (I1026141,I1026107,I264884);
nor I_60150 (I1026158,I1026065,I1026141);
DFFARX1 I_60151 (I1026158,I3563,I1026022,I1026008,);
nor I_60152 (I1026189,I264884,I264872);
nand I_60153 (I1026206,I1026189,I264887);
DFFARX1 I_60154 (I1026206,I3563,I1026022,I1026011,);
nor I_60155 (I1026237,I1026124,I264884);
nand I_60156 (I1026254,I1026237,I264866);
nor I_60157 (I1026271,I1026048,I1026254);
DFFARX1 I_60158 (I1026271,I3563,I1026022,I1025987,);
not I_60159 (I1026302,I1026254);
nand I_60160 (I1025999,I1026065,I1026302);
DFFARX1 I_60161 (I1026254,I3563,I1026022,I1026342,);
not I_60162 (I1026350,I1026342);
not I_60163 (I1026367,I264884);
not I_60164 (I1026384,I264875);
nor I_60165 (I1026401,I1026384,I264863);
nor I_60166 (I1026014,I1026350,I1026401);
nor I_60167 (I1026432,I1026384,I264878);
and I_60168 (I1026449,I1026432,I264866);
or I_60169 (I1026466,I1026449,I264863);
DFFARX1 I_60170 (I1026466,I3563,I1026022,I1026492,);
nor I_60171 (I1026002,I1026492,I1026048);
not I_60172 (I1026514,I1026492);
and I_60173 (I1026531,I1026514,I1026048);
nor I_60174 (I1025996,I1026073,I1026531);
nand I_60175 (I1026562,I1026514,I1026124);
nor I_60176 (I1025990,I1026384,I1026562);
nand I_60177 (I1025993,I1026514,I1026302);
nand I_60178 (I1026607,I1026124,I264875);
nor I_60179 (I1026005,I1026367,I1026607);
not I_60180 (I1026668,I3570);
DFFARX1 I_60181 (I182759,I3563,I1026668,I1026694,);
DFFARX1 I_60182 (I182771,I3563,I1026668,I1026711,);
not I_60183 (I1026719,I1026711);
not I_60184 (I1026736,I182777);
nor I_60185 (I1026753,I1026736,I182762);
not I_60186 (I1026770,I182753);
nor I_60187 (I1026787,I1026753,I182774);
nor I_60188 (I1026804,I1026711,I1026787);
DFFARX1 I_60189 (I1026804,I3563,I1026668,I1026654,);
nor I_60190 (I1026835,I182774,I182762);
nand I_60191 (I1026852,I1026835,I182777);
DFFARX1 I_60192 (I1026852,I3563,I1026668,I1026657,);
nor I_60193 (I1026883,I1026770,I182774);
nand I_60194 (I1026900,I1026883,I182756);
nor I_60195 (I1026917,I1026694,I1026900);
DFFARX1 I_60196 (I1026917,I3563,I1026668,I1026633,);
not I_60197 (I1026948,I1026900);
nand I_60198 (I1026645,I1026711,I1026948);
DFFARX1 I_60199 (I1026900,I3563,I1026668,I1026988,);
not I_60200 (I1026996,I1026988);
not I_60201 (I1027013,I182774);
not I_60202 (I1027030,I182765);
nor I_60203 (I1027047,I1027030,I182753);
nor I_60204 (I1026660,I1026996,I1027047);
nor I_60205 (I1027078,I1027030,I182768);
and I_60206 (I1027095,I1027078,I182756);
or I_60207 (I1027112,I1027095,I182753);
DFFARX1 I_60208 (I1027112,I3563,I1026668,I1027138,);
nor I_60209 (I1026648,I1027138,I1026694);
not I_60210 (I1027160,I1027138);
and I_60211 (I1027177,I1027160,I1026694);
nor I_60212 (I1026642,I1026719,I1027177);
nand I_60213 (I1027208,I1027160,I1026770);
nor I_60214 (I1026636,I1027030,I1027208);
nand I_60215 (I1026639,I1027160,I1026948);
nand I_60216 (I1027253,I1026770,I182765);
nor I_60217 (I1026651,I1027013,I1027253);
not I_60218 (I1027314,I3570);
DFFARX1 I_60219 (I739339,I3563,I1027314,I1027340,);
DFFARX1 I_60220 (I739333,I3563,I1027314,I1027357,);
not I_60221 (I1027365,I1027357);
not I_60222 (I1027382,I739348);
nor I_60223 (I1027399,I1027382,I739333);
not I_60224 (I1027416,I739342);
nor I_60225 (I1027433,I1027399,I739351);
nor I_60226 (I1027450,I1027357,I1027433);
DFFARX1 I_60227 (I1027450,I3563,I1027314,I1027300,);
nor I_60228 (I1027481,I739351,I739333);
nand I_60229 (I1027498,I1027481,I739348);
DFFARX1 I_60230 (I1027498,I3563,I1027314,I1027303,);
nor I_60231 (I1027529,I1027416,I739351);
nand I_60232 (I1027546,I1027529,I739336);
nor I_60233 (I1027563,I1027340,I1027546);
DFFARX1 I_60234 (I1027563,I3563,I1027314,I1027279,);
not I_60235 (I1027594,I1027546);
nand I_60236 (I1027291,I1027357,I1027594);
DFFARX1 I_60237 (I1027546,I3563,I1027314,I1027634,);
not I_60238 (I1027642,I1027634);
not I_60239 (I1027659,I739351);
not I_60240 (I1027676,I739345);
nor I_60241 (I1027693,I1027676,I739342);
nor I_60242 (I1027306,I1027642,I1027693);
nor I_60243 (I1027724,I1027676,I739354);
and I_60244 (I1027741,I1027724,I739357);
or I_60245 (I1027758,I1027741,I739336);
DFFARX1 I_60246 (I1027758,I3563,I1027314,I1027784,);
nor I_60247 (I1027294,I1027784,I1027340);
not I_60248 (I1027806,I1027784);
and I_60249 (I1027823,I1027806,I1027340);
nor I_60250 (I1027288,I1027365,I1027823);
nand I_60251 (I1027854,I1027806,I1027416);
nor I_60252 (I1027282,I1027676,I1027854);
nand I_60253 (I1027285,I1027806,I1027594);
nand I_60254 (I1027899,I1027416,I739345);
nor I_60255 (I1027297,I1027659,I1027899);
not I_60256 (I1027960,I3570);
DFFARX1 I_60257 (I1362468,I3563,I1027960,I1027986,);
DFFARX1 I_60258 (I1362492,I3563,I1027960,I1028003,);
not I_60259 (I1028011,I1028003);
not I_60260 (I1028028,I1362474);
nor I_60261 (I1028045,I1028028,I1362483);
not I_60262 (I1028062,I1362468);
nor I_60263 (I1028079,I1028045,I1362489);
nor I_60264 (I1028096,I1028003,I1028079);
DFFARX1 I_60265 (I1028096,I3563,I1027960,I1027946,);
nor I_60266 (I1028127,I1362489,I1362483);
nand I_60267 (I1028144,I1028127,I1362474);
DFFARX1 I_60268 (I1028144,I3563,I1027960,I1027949,);
nor I_60269 (I1028175,I1028062,I1362489);
nand I_60270 (I1028192,I1028175,I1362486);
nor I_60271 (I1028209,I1027986,I1028192);
DFFARX1 I_60272 (I1028209,I3563,I1027960,I1027925,);
not I_60273 (I1028240,I1028192);
nand I_60274 (I1027937,I1028003,I1028240);
DFFARX1 I_60275 (I1028192,I3563,I1027960,I1028280,);
not I_60276 (I1028288,I1028280);
not I_60277 (I1028305,I1362489);
not I_60278 (I1028322,I1362480);
nor I_60279 (I1028339,I1028322,I1362468);
nor I_60280 (I1027952,I1028288,I1028339);
nor I_60281 (I1028370,I1028322,I1362471);
and I_60282 (I1028387,I1028370,I1362495);
or I_60283 (I1028404,I1028387,I1362477);
DFFARX1 I_60284 (I1028404,I3563,I1027960,I1028430,);
nor I_60285 (I1027940,I1028430,I1027986);
not I_60286 (I1028452,I1028430);
and I_60287 (I1028469,I1028452,I1027986);
nor I_60288 (I1027934,I1028011,I1028469);
nand I_60289 (I1028500,I1028452,I1028062);
nor I_60290 (I1027928,I1028322,I1028500);
nand I_60291 (I1027931,I1028452,I1028240);
nand I_60292 (I1028545,I1028062,I1362480);
nor I_60293 (I1027943,I1028305,I1028545);
not I_60294 (I1028606,I3570);
DFFARX1 I_60295 (I1177713,I3563,I1028606,I1028632,);
DFFARX1 I_60296 (I1177695,I3563,I1028606,I1028649,);
not I_60297 (I1028657,I1028649);
not I_60298 (I1028674,I1177704);
nor I_60299 (I1028691,I1028674,I1177716);
not I_60300 (I1028708,I1177698);
nor I_60301 (I1028725,I1028691,I1177707);
nor I_60302 (I1028742,I1028649,I1028725);
DFFARX1 I_60303 (I1028742,I3563,I1028606,I1028592,);
nor I_60304 (I1028773,I1177707,I1177716);
nand I_60305 (I1028790,I1028773,I1177704);
DFFARX1 I_60306 (I1028790,I3563,I1028606,I1028595,);
nor I_60307 (I1028821,I1028708,I1177707);
nand I_60308 (I1028838,I1028821,I1177719);
nor I_60309 (I1028855,I1028632,I1028838);
DFFARX1 I_60310 (I1028855,I3563,I1028606,I1028571,);
not I_60311 (I1028886,I1028838);
nand I_60312 (I1028583,I1028649,I1028886);
DFFARX1 I_60313 (I1028838,I3563,I1028606,I1028926,);
not I_60314 (I1028934,I1028926);
not I_60315 (I1028951,I1177707);
not I_60316 (I1028968,I1177695);
nor I_60317 (I1028985,I1028968,I1177698);
nor I_60318 (I1028598,I1028934,I1028985);
nor I_60319 (I1029016,I1028968,I1177701);
and I_60320 (I1029033,I1029016,I1177710);
or I_60321 (I1029050,I1029033,I1177698);
DFFARX1 I_60322 (I1029050,I3563,I1028606,I1029076,);
nor I_60323 (I1028586,I1029076,I1028632);
not I_60324 (I1029098,I1029076);
and I_60325 (I1029115,I1029098,I1028632);
nor I_60326 (I1028580,I1028657,I1029115);
nand I_60327 (I1029146,I1029098,I1028708);
nor I_60328 (I1028574,I1028968,I1029146);
nand I_60329 (I1028577,I1029098,I1028886);
nand I_60330 (I1029191,I1028708,I1177695);
nor I_60331 (I1028589,I1028951,I1029191);
not I_60332 (I1029252,I3570);
DFFARX1 I_60333 (I390238,I3563,I1029252,I1029278,);
DFFARX1 I_60334 (I390244,I3563,I1029252,I1029295,);
not I_60335 (I1029303,I1029295);
not I_60336 (I1029320,I390265);
nor I_60337 (I1029337,I1029320,I390253);
not I_60338 (I1029354,I390262);
nor I_60339 (I1029371,I1029337,I390247);
nor I_60340 (I1029388,I1029295,I1029371);
DFFARX1 I_60341 (I1029388,I3563,I1029252,I1029238,);
nor I_60342 (I1029419,I390247,I390253);
nand I_60343 (I1029436,I1029419,I390265);
DFFARX1 I_60344 (I1029436,I3563,I1029252,I1029241,);
nor I_60345 (I1029467,I1029354,I390247);
nand I_60346 (I1029484,I1029467,I390238);
nor I_60347 (I1029501,I1029278,I1029484);
DFFARX1 I_60348 (I1029501,I3563,I1029252,I1029217,);
not I_60349 (I1029532,I1029484);
nand I_60350 (I1029229,I1029295,I1029532);
DFFARX1 I_60351 (I1029484,I3563,I1029252,I1029572,);
not I_60352 (I1029580,I1029572);
not I_60353 (I1029597,I390247);
not I_60354 (I1029614,I390250);
nor I_60355 (I1029631,I1029614,I390262);
nor I_60356 (I1029244,I1029580,I1029631);
nor I_60357 (I1029662,I1029614,I390259);
and I_60358 (I1029679,I1029662,I390241);
or I_60359 (I1029696,I1029679,I390256);
DFFARX1 I_60360 (I1029696,I3563,I1029252,I1029722,);
nor I_60361 (I1029232,I1029722,I1029278);
not I_60362 (I1029744,I1029722);
and I_60363 (I1029761,I1029744,I1029278);
nor I_60364 (I1029226,I1029303,I1029761);
nand I_60365 (I1029792,I1029744,I1029354);
nor I_60366 (I1029220,I1029614,I1029792);
nand I_60367 (I1029223,I1029744,I1029532);
nand I_60368 (I1029837,I1029354,I390250);
nor I_60369 (I1029235,I1029597,I1029837);
not I_60370 (I1029898,I3570);
DFFARX1 I_60371 (I249399,I3563,I1029898,I1029924,);
DFFARX1 I_60372 (I249411,I3563,I1029898,I1029941,);
not I_60373 (I1029949,I1029941);
not I_60374 (I1029966,I249417);
nor I_60375 (I1029983,I1029966,I249402);
not I_60376 (I1030000,I249393);
nor I_60377 (I1030017,I1029983,I249414);
nor I_60378 (I1030034,I1029941,I1030017);
DFFARX1 I_60379 (I1030034,I3563,I1029898,I1029884,);
nor I_60380 (I1030065,I249414,I249402);
nand I_60381 (I1030082,I1030065,I249417);
DFFARX1 I_60382 (I1030082,I3563,I1029898,I1029887,);
nor I_60383 (I1030113,I1030000,I249414);
nand I_60384 (I1030130,I1030113,I249396);
nor I_60385 (I1030147,I1029924,I1030130);
DFFARX1 I_60386 (I1030147,I3563,I1029898,I1029863,);
not I_60387 (I1030178,I1030130);
nand I_60388 (I1029875,I1029941,I1030178);
DFFARX1 I_60389 (I1030130,I3563,I1029898,I1030218,);
not I_60390 (I1030226,I1030218);
not I_60391 (I1030243,I249414);
not I_60392 (I1030260,I249405);
nor I_60393 (I1030277,I1030260,I249393);
nor I_60394 (I1029890,I1030226,I1030277);
nor I_60395 (I1030308,I1030260,I249408);
and I_60396 (I1030325,I1030308,I249396);
or I_60397 (I1030342,I1030325,I249393);
DFFARX1 I_60398 (I1030342,I3563,I1029898,I1030368,);
nor I_60399 (I1029878,I1030368,I1029924);
not I_60400 (I1030390,I1030368);
and I_60401 (I1030407,I1030390,I1029924);
nor I_60402 (I1029872,I1029949,I1030407);
nand I_60403 (I1030438,I1030390,I1030000);
nor I_60404 (I1029866,I1030260,I1030438);
nand I_60405 (I1029869,I1030390,I1030178);
nand I_60406 (I1030483,I1030000,I249405);
nor I_60407 (I1029881,I1030243,I1030483);
not I_60408 (I1030544,I3570);
DFFARX1 I_60409 (I626626,I3563,I1030544,I1030570,);
DFFARX1 I_60410 (I626638,I3563,I1030544,I1030587,);
not I_60411 (I1030595,I1030587);
not I_60412 (I1030612,I626647);
nor I_60413 (I1030629,I1030612,I626623);
not I_60414 (I1030646,I626641);
nor I_60415 (I1030663,I1030629,I626635);
nor I_60416 (I1030680,I1030587,I1030663);
DFFARX1 I_60417 (I1030680,I3563,I1030544,I1030530,);
nor I_60418 (I1030711,I626635,I626623);
nand I_60419 (I1030728,I1030711,I626647);
DFFARX1 I_60420 (I1030728,I3563,I1030544,I1030533,);
nor I_60421 (I1030759,I1030646,I626635);
nand I_60422 (I1030776,I1030759,I626629);
nor I_60423 (I1030793,I1030570,I1030776);
DFFARX1 I_60424 (I1030793,I3563,I1030544,I1030509,);
not I_60425 (I1030824,I1030776);
nand I_60426 (I1030521,I1030587,I1030824);
DFFARX1 I_60427 (I1030776,I3563,I1030544,I1030864,);
not I_60428 (I1030872,I1030864);
not I_60429 (I1030889,I626635);
not I_60430 (I1030906,I626644);
nor I_60431 (I1030923,I1030906,I626641);
nor I_60432 (I1030536,I1030872,I1030923);
nor I_60433 (I1030954,I1030906,I626626);
and I_60434 (I1030971,I1030954,I626623);
or I_60435 (I1030988,I1030971,I626632);
DFFARX1 I_60436 (I1030988,I3563,I1030544,I1031014,);
nor I_60437 (I1030524,I1031014,I1030570);
not I_60438 (I1031036,I1031014);
and I_60439 (I1031053,I1031036,I1030570);
nor I_60440 (I1030518,I1030595,I1031053);
nand I_60441 (I1031084,I1031036,I1030646);
nor I_60442 (I1030512,I1030906,I1031084);
nand I_60443 (I1030515,I1031036,I1030824);
nand I_60444 (I1031129,I1030646,I626644);
nor I_60445 (I1030527,I1030889,I1031129);
not I_60446 (I1031190,I3570);
DFFARX1 I_60447 (I1395788,I3563,I1031190,I1031216,);
DFFARX1 I_60448 (I1395812,I3563,I1031190,I1031233,);
not I_60449 (I1031241,I1031233);
not I_60450 (I1031258,I1395794);
nor I_60451 (I1031275,I1031258,I1395803);
not I_60452 (I1031292,I1395788);
nor I_60453 (I1031309,I1031275,I1395809);
nor I_60454 (I1031326,I1031233,I1031309);
DFFARX1 I_60455 (I1031326,I3563,I1031190,I1031176,);
nor I_60456 (I1031357,I1395809,I1395803);
nand I_60457 (I1031374,I1031357,I1395794);
DFFARX1 I_60458 (I1031374,I3563,I1031190,I1031179,);
nor I_60459 (I1031405,I1031292,I1395809);
nand I_60460 (I1031422,I1031405,I1395806);
nor I_60461 (I1031439,I1031216,I1031422);
DFFARX1 I_60462 (I1031439,I3563,I1031190,I1031155,);
not I_60463 (I1031470,I1031422);
nand I_60464 (I1031167,I1031233,I1031470);
DFFARX1 I_60465 (I1031422,I3563,I1031190,I1031510,);
not I_60466 (I1031518,I1031510);
not I_60467 (I1031535,I1395809);
not I_60468 (I1031552,I1395800);
nor I_60469 (I1031569,I1031552,I1395788);
nor I_60470 (I1031182,I1031518,I1031569);
nor I_60471 (I1031600,I1031552,I1395791);
and I_60472 (I1031617,I1031600,I1395815);
or I_60473 (I1031634,I1031617,I1395797);
DFFARX1 I_60474 (I1031634,I3563,I1031190,I1031660,);
nor I_60475 (I1031170,I1031660,I1031216);
not I_60476 (I1031682,I1031660);
and I_60477 (I1031699,I1031682,I1031216);
nor I_60478 (I1031164,I1031241,I1031699);
nand I_60479 (I1031730,I1031682,I1031292);
nor I_60480 (I1031158,I1031552,I1031730);
nand I_60481 (I1031161,I1031682,I1031470);
nand I_60482 (I1031775,I1031292,I1395800);
nor I_60483 (I1031173,I1031535,I1031775);
not I_60484 (I1031836,I3570);
DFFARX1 I_60485 (I504008,I3563,I1031836,I1031862,);
DFFARX1 I_60486 (I504005,I3563,I1031836,I1031879,);
not I_60487 (I1031887,I1031879);
not I_60488 (I1031904,I504020);
nor I_60489 (I1031921,I1031904,I504023);
not I_60490 (I1031938,I504011);
nor I_60491 (I1031955,I1031921,I504017);
nor I_60492 (I1031972,I1031879,I1031955);
DFFARX1 I_60493 (I1031972,I3563,I1031836,I1031822,);
nor I_60494 (I1032003,I504017,I504023);
nand I_60495 (I1032020,I1032003,I504020);
DFFARX1 I_60496 (I1032020,I3563,I1031836,I1031825,);
nor I_60497 (I1032051,I1031938,I504017);
nand I_60498 (I1032068,I1032051,I504029);
nor I_60499 (I1032085,I1031862,I1032068);
DFFARX1 I_60500 (I1032085,I3563,I1031836,I1031801,);
not I_60501 (I1032116,I1032068);
nand I_60502 (I1031813,I1031879,I1032116);
DFFARX1 I_60503 (I1032068,I3563,I1031836,I1032156,);
not I_60504 (I1032164,I1032156);
not I_60505 (I1032181,I504017);
not I_60506 (I1032198,I504002);
nor I_60507 (I1032215,I1032198,I504011);
nor I_60508 (I1031828,I1032164,I1032215);
nor I_60509 (I1032246,I1032198,I504014);
and I_60510 (I1032263,I1032246,I504002);
or I_60511 (I1032280,I1032263,I504026);
DFFARX1 I_60512 (I1032280,I3563,I1031836,I1032306,);
nor I_60513 (I1031816,I1032306,I1031862);
not I_60514 (I1032328,I1032306);
and I_60515 (I1032345,I1032328,I1031862);
nor I_60516 (I1031810,I1031887,I1032345);
nand I_60517 (I1032376,I1032328,I1031938);
nor I_60518 (I1031804,I1032198,I1032376);
nand I_60519 (I1031807,I1032328,I1032116);
nand I_60520 (I1032421,I1031938,I504002);
nor I_60521 (I1031819,I1032181,I1032421);
not I_60522 (I1032482,I3570);
DFFARX1 I_60523 (I812643,I3563,I1032482,I1032508,);
DFFARX1 I_60524 (I812640,I3563,I1032482,I1032525,);
not I_60525 (I1032533,I1032525);
not I_60526 (I1032550,I812640);
nor I_60527 (I1032567,I1032550,I812643);
not I_60528 (I1032584,I812655);
nor I_60529 (I1032601,I1032567,I812649);
nor I_60530 (I1032618,I1032525,I1032601);
DFFARX1 I_60531 (I1032618,I3563,I1032482,I1032468,);
nor I_60532 (I1032649,I812649,I812643);
nand I_60533 (I1032666,I1032649,I812640);
DFFARX1 I_60534 (I1032666,I3563,I1032482,I1032471,);
nor I_60535 (I1032697,I1032584,I812649);
nand I_60536 (I1032714,I1032697,I812637);
nor I_60537 (I1032731,I1032508,I1032714);
DFFARX1 I_60538 (I1032731,I3563,I1032482,I1032447,);
not I_60539 (I1032762,I1032714);
nand I_60540 (I1032459,I1032525,I1032762);
DFFARX1 I_60541 (I1032714,I3563,I1032482,I1032802,);
not I_60542 (I1032810,I1032802);
not I_60543 (I1032827,I812649);
not I_60544 (I1032844,I812646);
nor I_60545 (I1032861,I1032844,I812655);
nor I_60546 (I1032474,I1032810,I1032861);
nor I_60547 (I1032892,I1032844,I812652);
and I_60548 (I1032909,I1032892,I812658);
or I_60549 (I1032926,I1032909,I812637);
DFFARX1 I_60550 (I1032926,I3563,I1032482,I1032952,);
nor I_60551 (I1032462,I1032952,I1032508);
not I_60552 (I1032974,I1032952);
and I_60553 (I1032991,I1032974,I1032508);
nor I_60554 (I1032456,I1032533,I1032991);
nand I_60555 (I1033022,I1032974,I1032584);
nor I_60556 (I1032450,I1032844,I1033022);
nand I_60557 (I1032453,I1032974,I1032762);
nand I_60558 (I1033067,I1032584,I812646);
nor I_60559 (I1032465,I1032827,I1033067);
not I_60560 (I1033128,I3570);
DFFARX1 I_60561 (I632406,I3563,I1033128,I1033154,);
DFFARX1 I_60562 (I632418,I3563,I1033128,I1033171,);
not I_60563 (I1033179,I1033171);
not I_60564 (I1033196,I632427);
nor I_60565 (I1033213,I1033196,I632403);
not I_60566 (I1033230,I632421);
nor I_60567 (I1033247,I1033213,I632415);
nor I_60568 (I1033264,I1033171,I1033247);
DFFARX1 I_60569 (I1033264,I3563,I1033128,I1033114,);
nor I_60570 (I1033295,I632415,I632403);
nand I_60571 (I1033312,I1033295,I632427);
DFFARX1 I_60572 (I1033312,I3563,I1033128,I1033117,);
nor I_60573 (I1033343,I1033230,I632415);
nand I_60574 (I1033360,I1033343,I632409);
nor I_60575 (I1033377,I1033154,I1033360);
DFFARX1 I_60576 (I1033377,I3563,I1033128,I1033093,);
not I_60577 (I1033408,I1033360);
nand I_60578 (I1033105,I1033171,I1033408);
DFFARX1 I_60579 (I1033360,I3563,I1033128,I1033448,);
not I_60580 (I1033456,I1033448);
not I_60581 (I1033473,I632415);
not I_60582 (I1033490,I632424);
nor I_60583 (I1033507,I1033490,I632421);
nor I_60584 (I1033120,I1033456,I1033507);
nor I_60585 (I1033538,I1033490,I632406);
and I_60586 (I1033555,I1033538,I632403);
or I_60587 (I1033572,I1033555,I632412);
DFFARX1 I_60588 (I1033572,I3563,I1033128,I1033598,);
nor I_60589 (I1033108,I1033598,I1033154);
not I_60590 (I1033620,I1033598);
and I_60591 (I1033637,I1033620,I1033154);
nor I_60592 (I1033102,I1033179,I1033637);
nand I_60593 (I1033668,I1033620,I1033230);
nor I_60594 (I1033096,I1033490,I1033668);
nand I_60595 (I1033099,I1033620,I1033408);
nand I_60596 (I1033713,I1033230,I632424);
nor I_60597 (I1033111,I1033473,I1033713);
not I_60598 (I1033774,I3570);
DFFARX1 I_60599 (I879572,I3563,I1033774,I1033800,);
DFFARX1 I_60600 (I879569,I3563,I1033774,I1033817,);
not I_60601 (I1033825,I1033817);
not I_60602 (I1033842,I879569);
nor I_60603 (I1033859,I1033842,I879572);
not I_60604 (I1033876,I879584);
nor I_60605 (I1033893,I1033859,I879578);
nor I_60606 (I1033910,I1033817,I1033893);
DFFARX1 I_60607 (I1033910,I3563,I1033774,I1033760,);
nor I_60608 (I1033941,I879578,I879572);
nand I_60609 (I1033958,I1033941,I879569);
DFFARX1 I_60610 (I1033958,I3563,I1033774,I1033763,);
nor I_60611 (I1033989,I1033876,I879578);
nand I_60612 (I1034006,I1033989,I879566);
nor I_60613 (I1034023,I1033800,I1034006);
DFFARX1 I_60614 (I1034023,I3563,I1033774,I1033739,);
not I_60615 (I1034054,I1034006);
nand I_60616 (I1033751,I1033817,I1034054);
DFFARX1 I_60617 (I1034006,I3563,I1033774,I1034094,);
not I_60618 (I1034102,I1034094);
not I_60619 (I1034119,I879578);
not I_60620 (I1034136,I879575);
nor I_60621 (I1034153,I1034136,I879584);
nor I_60622 (I1033766,I1034102,I1034153);
nor I_60623 (I1034184,I1034136,I879581);
and I_60624 (I1034201,I1034184,I879587);
or I_60625 (I1034218,I1034201,I879566);
DFFARX1 I_60626 (I1034218,I3563,I1033774,I1034244,);
nor I_60627 (I1033754,I1034244,I1033800);
not I_60628 (I1034266,I1034244);
and I_60629 (I1034283,I1034266,I1033800);
nor I_60630 (I1033748,I1033825,I1034283);
nand I_60631 (I1034314,I1034266,I1033876);
nor I_60632 (I1033742,I1034136,I1034314);
nand I_60633 (I1033745,I1034266,I1034054);
nand I_60634 (I1034359,I1033876,I879575);
nor I_60635 (I1033757,I1034119,I1034359);
not I_60636 (I1034420,I3570);
DFFARX1 I_60637 (I359145,I3563,I1034420,I1034446,);
DFFARX1 I_60638 (I359151,I3563,I1034420,I1034463,);
not I_60639 (I1034471,I1034463);
not I_60640 (I1034488,I359172);
nor I_60641 (I1034505,I1034488,I359160);
not I_60642 (I1034522,I359169);
nor I_60643 (I1034539,I1034505,I359154);
nor I_60644 (I1034556,I1034463,I1034539);
DFFARX1 I_60645 (I1034556,I3563,I1034420,I1034406,);
nor I_60646 (I1034587,I359154,I359160);
nand I_60647 (I1034604,I1034587,I359172);
DFFARX1 I_60648 (I1034604,I3563,I1034420,I1034409,);
nor I_60649 (I1034635,I1034522,I359154);
nand I_60650 (I1034652,I1034635,I359145);
nor I_60651 (I1034669,I1034446,I1034652);
DFFARX1 I_60652 (I1034669,I3563,I1034420,I1034385,);
not I_60653 (I1034700,I1034652);
nand I_60654 (I1034397,I1034463,I1034700);
DFFARX1 I_60655 (I1034652,I3563,I1034420,I1034740,);
not I_60656 (I1034748,I1034740);
not I_60657 (I1034765,I359154);
not I_60658 (I1034782,I359157);
nor I_60659 (I1034799,I1034782,I359169);
nor I_60660 (I1034412,I1034748,I1034799);
nor I_60661 (I1034830,I1034782,I359166);
and I_60662 (I1034847,I1034830,I359148);
or I_60663 (I1034864,I1034847,I359163);
DFFARX1 I_60664 (I1034864,I3563,I1034420,I1034890,);
nor I_60665 (I1034400,I1034890,I1034446);
not I_60666 (I1034912,I1034890);
and I_60667 (I1034929,I1034912,I1034446);
nor I_60668 (I1034394,I1034471,I1034929);
nand I_60669 (I1034960,I1034912,I1034522);
nor I_60670 (I1034388,I1034782,I1034960);
nand I_60671 (I1034391,I1034912,I1034700);
nand I_60672 (I1035005,I1034522,I359157);
nor I_60673 (I1034403,I1034765,I1035005);
not I_60674 (I1035066,I3570);
DFFARX1 I_60675 (I158971,I3563,I1035066,I1035092,);
DFFARX1 I_60676 (I158974,I3563,I1035066,I1035109,);
not I_60677 (I1035117,I1035109);
not I_60678 (I1035134,I158959);
nor I_60679 (I1035151,I1035134,I158953);
not I_60680 (I1035168,I158962);
nor I_60681 (I1035185,I1035151,I158977);
nor I_60682 (I1035202,I1035109,I1035185);
DFFARX1 I_60683 (I1035202,I3563,I1035066,I1035052,);
nor I_60684 (I1035233,I158977,I158953);
nand I_60685 (I1035250,I1035233,I158959);
DFFARX1 I_60686 (I1035250,I3563,I1035066,I1035055,);
nor I_60687 (I1035281,I1035168,I158977);
nand I_60688 (I1035298,I1035281,I158980);
nor I_60689 (I1035315,I1035092,I1035298);
DFFARX1 I_60690 (I1035315,I3563,I1035066,I1035031,);
not I_60691 (I1035346,I1035298);
nand I_60692 (I1035043,I1035109,I1035346);
DFFARX1 I_60693 (I1035298,I3563,I1035066,I1035386,);
not I_60694 (I1035394,I1035386);
not I_60695 (I1035411,I158977);
not I_60696 (I1035428,I158956);
nor I_60697 (I1035445,I1035428,I158962);
nor I_60698 (I1035058,I1035394,I1035445);
nor I_60699 (I1035476,I1035428,I158965);
and I_60700 (I1035493,I1035476,I158953);
or I_60701 (I1035510,I1035493,I158968);
DFFARX1 I_60702 (I1035510,I3563,I1035066,I1035536,);
nor I_60703 (I1035046,I1035536,I1035092);
not I_60704 (I1035558,I1035536);
and I_60705 (I1035575,I1035558,I1035092);
nor I_60706 (I1035040,I1035117,I1035575);
nand I_60707 (I1035606,I1035558,I1035168);
nor I_60708 (I1035034,I1035428,I1035606);
nand I_60709 (I1035037,I1035558,I1035346);
nand I_60710 (I1035651,I1035168,I158956);
nor I_60711 (I1035049,I1035411,I1035651);
not I_60712 (I1035712,I3570);
DFFARX1 I_60713 (I893801,I3563,I1035712,I1035738,);
DFFARX1 I_60714 (I893798,I3563,I1035712,I1035755,);
not I_60715 (I1035763,I1035755);
not I_60716 (I1035780,I893798);
nor I_60717 (I1035797,I1035780,I893801);
not I_60718 (I1035814,I893813);
nor I_60719 (I1035831,I1035797,I893807);
nor I_60720 (I1035848,I1035755,I1035831);
DFFARX1 I_60721 (I1035848,I3563,I1035712,I1035698,);
nor I_60722 (I1035879,I893807,I893801);
nand I_60723 (I1035896,I1035879,I893798);
DFFARX1 I_60724 (I1035896,I3563,I1035712,I1035701,);
nor I_60725 (I1035927,I1035814,I893807);
nand I_60726 (I1035944,I1035927,I893795);
nor I_60727 (I1035961,I1035738,I1035944);
DFFARX1 I_60728 (I1035961,I3563,I1035712,I1035677,);
not I_60729 (I1035992,I1035944);
nand I_60730 (I1035689,I1035755,I1035992);
DFFARX1 I_60731 (I1035944,I3563,I1035712,I1036032,);
not I_60732 (I1036040,I1036032);
not I_60733 (I1036057,I893807);
not I_60734 (I1036074,I893804);
nor I_60735 (I1036091,I1036074,I893813);
nor I_60736 (I1035704,I1036040,I1036091);
nor I_60737 (I1036122,I1036074,I893810);
and I_60738 (I1036139,I1036122,I893816);
or I_60739 (I1036156,I1036139,I893795);
DFFARX1 I_60740 (I1036156,I3563,I1035712,I1036182,);
nor I_60741 (I1035692,I1036182,I1035738);
not I_60742 (I1036204,I1036182);
and I_60743 (I1036221,I1036204,I1035738);
nor I_60744 (I1035686,I1035763,I1036221);
nand I_60745 (I1036252,I1036204,I1035814);
nor I_60746 (I1035680,I1036074,I1036252);
nand I_60747 (I1035683,I1036204,I1035992);
nand I_60748 (I1036297,I1035814,I893804);
nor I_60749 (I1035695,I1036057,I1036297);
not I_60750 (I1036358,I3570);
DFFARX1 I_60751 (I489320,I3563,I1036358,I1036384,);
DFFARX1 I_60752 (I489317,I3563,I1036358,I1036401,);
not I_60753 (I1036409,I1036401);
not I_60754 (I1036426,I489332);
nor I_60755 (I1036443,I1036426,I489335);
not I_60756 (I1036460,I489323);
nor I_60757 (I1036477,I1036443,I489329);
nor I_60758 (I1036494,I1036401,I1036477);
DFFARX1 I_60759 (I1036494,I3563,I1036358,I1036344,);
nor I_60760 (I1036525,I489329,I489335);
nand I_60761 (I1036542,I1036525,I489332);
DFFARX1 I_60762 (I1036542,I3563,I1036358,I1036347,);
nor I_60763 (I1036573,I1036460,I489329);
nand I_60764 (I1036590,I1036573,I489341);
nor I_60765 (I1036607,I1036384,I1036590);
DFFARX1 I_60766 (I1036607,I3563,I1036358,I1036323,);
not I_60767 (I1036638,I1036590);
nand I_60768 (I1036335,I1036401,I1036638);
DFFARX1 I_60769 (I1036590,I3563,I1036358,I1036678,);
not I_60770 (I1036686,I1036678);
not I_60771 (I1036703,I489329);
not I_60772 (I1036720,I489314);
nor I_60773 (I1036737,I1036720,I489323);
nor I_60774 (I1036350,I1036686,I1036737);
nor I_60775 (I1036768,I1036720,I489326);
and I_60776 (I1036785,I1036768,I489314);
or I_60777 (I1036802,I1036785,I489338);
DFFARX1 I_60778 (I1036802,I3563,I1036358,I1036828,);
nor I_60779 (I1036338,I1036828,I1036384);
not I_60780 (I1036850,I1036828);
and I_60781 (I1036867,I1036850,I1036384);
nor I_60782 (I1036332,I1036409,I1036867);
nand I_60783 (I1036898,I1036850,I1036460);
nor I_60784 (I1036326,I1036720,I1036898);
nand I_60785 (I1036329,I1036850,I1036638);
nand I_60786 (I1036943,I1036460,I489314);
nor I_60787 (I1036341,I1036703,I1036943);
not I_60788 (I1037004,I3570);
DFFARX1 I_60789 (I89848,I3563,I1037004,I1037030,);
DFFARX1 I_60790 (I89854,I3563,I1037004,I1037047,);
not I_60791 (I1037055,I1037047);
not I_60792 (I1037072,I89872);
nor I_60793 (I1037089,I1037072,I89851);
not I_60794 (I1037106,I89857);
nor I_60795 (I1037123,I1037089,I89863);
nor I_60796 (I1037140,I1037047,I1037123);
DFFARX1 I_60797 (I1037140,I3563,I1037004,I1036990,);
nor I_60798 (I1037171,I89863,I89851);
nand I_60799 (I1037188,I1037171,I89872);
DFFARX1 I_60800 (I1037188,I3563,I1037004,I1036993,);
nor I_60801 (I1037219,I1037106,I89863);
nand I_60802 (I1037236,I1037219,I89869);
nor I_60803 (I1037253,I1037030,I1037236);
DFFARX1 I_60804 (I1037253,I3563,I1037004,I1036969,);
not I_60805 (I1037284,I1037236);
nand I_60806 (I1036981,I1037047,I1037284);
DFFARX1 I_60807 (I1037236,I3563,I1037004,I1037324,);
not I_60808 (I1037332,I1037324);
not I_60809 (I1037349,I89863);
not I_60810 (I1037366,I89851);
nor I_60811 (I1037383,I1037366,I89857);
nor I_60812 (I1036996,I1037332,I1037383);
nor I_60813 (I1037414,I1037366,I89860);
and I_60814 (I1037431,I1037414,I89848);
or I_60815 (I1037448,I1037431,I89866);
DFFARX1 I_60816 (I1037448,I3563,I1037004,I1037474,);
nor I_60817 (I1036984,I1037474,I1037030);
not I_60818 (I1037496,I1037474);
and I_60819 (I1037513,I1037496,I1037030);
nor I_60820 (I1036978,I1037055,I1037513);
nand I_60821 (I1037544,I1037496,I1037106);
nor I_60822 (I1036972,I1037366,I1037544);
nand I_60823 (I1036975,I1037496,I1037284);
nand I_60824 (I1037589,I1037106,I89851);
nor I_60825 (I1036987,I1037349,I1037589);
not I_60826 (I1037650,I3570);
DFFARX1 I_60827 (I1214127,I3563,I1037650,I1037676,);
DFFARX1 I_60828 (I1214109,I3563,I1037650,I1037693,);
not I_60829 (I1037701,I1037693);
not I_60830 (I1037718,I1214118);
nor I_60831 (I1037735,I1037718,I1214130);
not I_60832 (I1037752,I1214112);
nor I_60833 (I1037769,I1037735,I1214121);
nor I_60834 (I1037786,I1037693,I1037769);
DFFARX1 I_60835 (I1037786,I3563,I1037650,I1037636,);
nor I_60836 (I1037817,I1214121,I1214130);
nand I_60837 (I1037834,I1037817,I1214118);
DFFARX1 I_60838 (I1037834,I3563,I1037650,I1037639,);
nor I_60839 (I1037865,I1037752,I1214121);
nand I_60840 (I1037882,I1037865,I1214133);
nor I_60841 (I1037899,I1037676,I1037882);
DFFARX1 I_60842 (I1037899,I3563,I1037650,I1037615,);
not I_60843 (I1037930,I1037882);
nand I_60844 (I1037627,I1037693,I1037930);
DFFARX1 I_60845 (I1037882,I3563,I1037650,I1037970,);
not I_60846 (I1037978,I1037970);
not I_60847 (I1037995,I1214121);
not I_60848 (I1038012,I1214109);
nor I_60849 (I1038029,I1038012,I1214112);
nor I_60850 (I1037642,I1037978,I1038029);
nor I_60851 (I1038060,I1038012,I1214115);
and I_60852 (I1038077,I1038060,I1214124);
or I_60853 (I1038094,I1038077,I1214112);
DFFARX1 I_60854 (I1038094,I3563,I1037650,I1038120,);
nor I_60855 (I1037630,I1038120,I1037676);
not I_60856 (I1038142,I1038120);
and I_60857 (I1038159,I1038142,I1037676);
nor I_60858 (I1037624,I1037701,I1038159);
nand I_60859 (I1038190,I1038142,I1037752);
nor I_60860 (I1037618,I1038012,I1038190);
nand I_60861 (I1037621,I1038142,I1037930);
nand I_60862 (I1038235,I1037752,I1214109);
nor I_60863 (I1037633,I1037995,I1038235);
not I_60864 (I1038296,I3570);
DFFARX1 I_60865 (I329633,I3563,I1038296,I1038322,);
DFFARX1 I_60866 (I329639,I3563,I1038296,I1038339,);
not I_60867 (I1038347,I1038339);
not I_60868 (I1038364,I329660);
nor I_60869 (I1038381,I1038364,I329648);
not I_60870 (I1038398,I329657);
nor I_60871 (I1038415,I1038381,I329642);
nor I_60872 (I1038432,I1038339,I1038415);
DFFARX1 I_60873 (I1038432,I3563,I1038296,I1038282,);
nor I_60874 (I1038463,I329642,I329648);
nand I_60875 (I1038480,I1038463,I329660);
DFFARX1 I_60876 (I1038480,I3563,I1038296,I1038285,);
nor I_60877 (I1038511,I1038398,I329642);
nand I_60878 (I1038528,I1038511,I329633);
nor I_60879 (I1038545,I1038322,I1038528);
DFFARX1 I_60880 (I1038545,I3563,I1038296,I1038261,);
not I_60881 (I1038576,I1038528);
nand I_60882 (I1038273,I1038339,I1038576);
DFFARX1 I_60883 (I1038528,I3563,I1038296,I1038616,);
not I_60884 (I1038624,I1038616);
not I_60885 (I1038641,I329642);
not I_60886 (I1038658,I329645);
nor I_60887 (I1038675,I1038658,I329657);
nor I_60888 (I1038288,I1038624,I1038675);
nor I_60889 (I1038706,I1038658,I329654);
and I_60890 (I1038723,I1038706,I329636);
or I_60891 (I1038740,I1038723,I329651);
DFFARX1 I_60892 (I1038740,I3563,I1038296,I1038766,);
nor I_60893 (I1038276,I1038766,I1038322);
not I_60894 (I1038788,I1038766);
and I_60895 (I1038805,I1038788,I1038322);
nor I_60896 (I1038270,I1038347,I1038805);
nand I_60897 (I1038836,I1038788,I1038398);
nor I_60898 (I1038264,I1038658,I1038836);
nand I_60899 (I1038267,I1038788,I1038576);
nand I_60900 (I1038881,I1038398,I329645);
nor I_60901 (I1038279,I1038641,I1038881);
not I_60902 (I1038942,I3570);
DFFARX1 I_60903 (I285694,I3563,I1038942,I1038968,);
DFFARX1 I_60904 (I285706,I3563,I1038942,I1038985,);
not I_60905 (I1038993,I1038985);
not I_60906 (I1039010,I285712);
nor I_60907 (I1039027,I1039010,I285697);
not I_60908 (I1039044,I285688);
nor I_60909 (I1039061,I1039027,I285709);
nor I_60910 (I1039078,I1038985,I1039061);
DFFARX1 I_60911 (I1039078,I3563,I1038942,I1038928,);
nor I_60912 (I1039109,I285709,I285697);
nand I_60913 (I1039126,I1039109,I285712);
DFFARX1 I_60914 (I1039126,I3563,I1038942,I1038931,);
nor I_60915 (I1039157,I1039044,I285709);
nand I_60916 (I1039174,I1039157,I285691);
nor I_60917 (I1039191,I1038968,I1039174);
DFFARX1 I_60918 (I1039191,I3563,I1038942,I1038907,);
not I_60919 (I1039222,I1039174);
nand I_60920 (I1038919,I1038985,I1039222);
DFFARX1 I_60921 (I1039174,I3563,I1038942,I1039262,);
not I_60922 (I1039270,I1039262);
not I_60923 (I1039287,I285709);
not I_60924 (I1039304,I285700);
nor I_60925 (I1039321,I1039304,I285688);
nor I_60926 (I1038934,I1039270,I1039321);
nor I_60927 (I1039352,I1039304,I285703);
and I_60928 (I1039369,I1039352,I285691);
or I_60929 (I1039386,I1039369,I285688);
DFFARX1 I_60930 (I1039386,I3563,I1038942,I1039412,);
nor I_60931 (I1038922,I1039412,I1038968);
not I_60932 (I1039434,I1039412);
and I_60933 (I1039451,I1039434,I1038968);
nor I_60934 (I1038916,I1038993,I1039451);
nand I_60935 (I1039482,I1039434,I1039044);
nor I_60936 (I1038910,I1039304,I1039482);
nand I_60937 (I1038913,I1039434,I1039222);
nand I_60938 (I1039527,I1039044,I285700);
nor I_60939 (I1038925,I1039287,I1039527);
not I_60940 (I1039588,I3570);
DFFARX1 I_60941 (I399724,I3563,I1039588,I1039614,);
DFFARX1 I_60942 (I399730,I3563,I1039588,I1039631,);
not I_60943 (I1039639,I1039631);
not I_60944 (I1039656,I399751);
nor I_60945 (I1039673,I1039656,I399739);
not I_60946 (I1039690,I399748);
nor I_60947 (I1039707,I1039673,I399733);
nor I_60948 (I1039724,I1039631,I1039707);
DFFARX1 I_60949 (I1039724,I3563,I1039588,I1039574,);
nor I_60950 (I1039755,I399733,I399739);
nand I_60951 (I1039772,I1039755,I399751);
DFFARX1 I_60952 (I1039772,I3563,I1039588,I1039577,);
nor I_60953 (I1039803,I1039690,I399733);
nand I_60954 (I1039820,I1039803,I399724);
nor I_60955 (I1039837,I1039614,I1039820);
DFFARX1 I_60956 (I1039837,I3563,I1039588,I1039553,);
not I_60957 (I1039868,I1039820);
nand I_60958 (I1039565,I1039631,I1039868);
DFFARX1 I_60959 (I1039820,I3563,I1039588,I1039908,);
not I_60960 (I1039916,I1039908);
not I_60961 (I1039933,I399733);
not I_60962 (I1039950,I399736);
nor I_60963 (I1039967,I1039950,I399748);
nor I_60964 (I1039580,I1039916,I1039967);
nor I_60965 (I1039998,I1039950,I399745);
and I_60966 (I1040015,I1039998,I399727);
or I_60967 (I1040032,I1040015,I399742);
DFFARX1 I_60968 (I1040032,I3563,I1039588,I1040058,);
nor I_60969 (I1039568,I1040058,I1039614);
not I_60970 (I1040080,I1040058);
and I_60971 (I1040097,I1040080,I1039614);
nor I_60972 (I1039562,I1039639,I1040097);
nand I_60973 (I1040128,I1040080,I1039690);
nor I_60974 (I1039556,I1039950,I1040128);
nand I_60975 (I1039559,I1040080,I1039868);
nand I_60976 (I1040173,I1039690,I399736);
nor I_60977 (I1039571,I1039933,I1040173);
not I_60978 (I1040234,I3570);
DFFARX1 I_60979 (I334376,I3563,I1040234,I1040260,);
DFFARX1 I_60980 (I334382,I3563,I1040234,I1040277,);
not I_60981 (I1040285,I1040277);
not I_60982 (I1040302,I334403);
nor I_60983 (I1040319,I1040302,I334391);
not I_60984 (I1040336,I334400);
nor I_60985 (I1040353,I1040319,I334385);
nor I_60986 (I1040370,I1040277,I1040353);
DFFARX1 I_60987 (I1040370,I3563,I1040234,I1040220,);
nor I_60988 (I1040401,I334385,I334391);
nand I_60989 (I1040418,I1040401,I334403);
DFFARX1 I_60990 (I1040418,I3563,I1040234,I1040223,);
nor I_60991 (I1040449,I1040336,I334385);
nand I_60992 (I1040466,I1040449,I334376);
nor I_60993 (I1040483,I1040260,I1040466);
DFFARX1 I_60994 (I1040483,I3563,I1040234,I1040199,);
not I_60995 (I1040514,I1040466);
nand I_60996 (I1040211,I1040277,I1040514);
DFFARX1 I_60997 (I1040466,I3563,I1040234,I1040554,);
not I_60998 (I1040562,I1040554);
not I_60999 (I1040579,I334385);
not I_61000 (I1040596,I334388);
nor I_61001 (I1040613,I1040596,I334400);
nor I_61002 (I1040226,I1040562,I1040613);
nor I_61003 (I1040644,I1040596,I334397);
and I_61004 (I1040661,I1040644,I334379);
or I_61005 (I1040678,I1040661,I334394);
DFFARX1 I_61006 (I1040678,I3563,I1040234,I1040704,);
nor I_61007 (I1040214,I1040704,I1040260);
not I_61008 (I1040726,I1040704);
and I_61009 (I1040743,I1040726,I1040260);
nor I_61010 (I1040208,I1040285,I1040743);
nand I_61011 (I1040774,I1040726,I1040336);
nor I_61012 (I1040202,I1040596,I1040774);
nand I_61013 (I1040205,I1040726,I1040514);
nand I_61014 (I1040819,I1040336,I334388);
nor I_61015 (I1040217,I1040579,I1040819);
not I_61016 (I1040880,I3570);
DFFARX1 I_61017 (I128846,I3563,I1040880,I1040906,);
DFFARX1 I_61018 (I128852,I3563,I1040880,I1040923,);
not I_61019 (I1040931,I1040923);
not I_61020 (I1040948,I128870);
nor I_61021 (I1040965,I1040948,I128849);
not I_61022 (I1040982,I128855);
nor I_61023 (I1040999,I1040965,I128861);
nor I_61024 (I1041016,I1040923,I1040999);
DFFARX1 I_61025 (I1041016,I3563,I1040880,I1040866,);
nor I_61026 (I1041047,I128861,I128849);
nand I_61027 (I1041064,I1041047,I128870);
DFFARX1 I_61028 (I1041064,I3563,I1040880,I1040869,);
nor I_61029 (I1041095,I1040982,I128861);
nand I_61030 (I1041112,I1041095,I128867);
nor I_61031 (I1041129,I1040906,I1041112);
DFFARX1 I_61032 (I1041129,I3563,I1040880,I1040845,);
not I_61033 (I1041160,I1041112);
nand I_61034 (I1040857,I1040923,I1041160);
DFFARX1 I_61035 (I1041112,I3563,I1040880,I1041200,);
not I_61036 (I1041208,I1041200);
not I_61037 (I1041225,I128861);
not I_61038 (I1041242,I128849);
nor I_61039 (I1041259,I1041242,I128855);
nor I_61040 (I1040872,I1041208,I1041259);
nor I_61041 (I1041290,I1041242,I128858);
and I_61042 (I1041307,I1041290,I128846);
or I_61043 (I1041324,I1041307,I128864);
DFFARX1 I_61044 (I1041324,I3563,I1040880,I1041350,);
nor I_61045 (I1040860,I1041350,I1040906);
not I_61046 (I1041372,I1041350);
and I_61047 (I1041389,I1041372,I1040906);
nor I_61048 (I1040854,I1040931,I1041389);
nand I_61049 (I1041420,I1041372,I1040982);
nor I_61050 (I1040848,I1041242,I1041420);
nand I_61051 (I1040851,I1041372,I1041160);
nand I_61052 (I1041465,I1040982,I128849);
nor I_61053 (I1040863,I1041225,I1041465);
not I_61054 (I1041526,I3570);
DFFARX1 I_61055 (I252374,I3563,I1041526,I1041552,);
DFFARX1 I_61056 (I252386,I3563,I1041526,I1041569,);
not I_61057 (I1041577,I1041569);
not I_61058 (I1041594,I252392);
nor I_61059 (I1041611,I1041594,I252377);
not I_61060 (I1041628,I252368);
nor I_61061 (I1041645,I1041611,I252389);
nor I_61062 (I1041662,I1041569,I1041645);
DFFARX1 I_61063 (I1041662,I3563,I1041526,I1041512,);
nor I_61064 (I1041693,I252389,I252377);
nand I_61065 (I1041710,I1041693,I252392);
DFFARX1 I_61066 (I1041710,I3563,I1041526,I1041515,);
nor I_61067 (I1041741,I1041628,I252389);
nand I_61068 (I1041758,I1041741,I252371);
nor I_61069 (I1041775,I1041552,I1041758);
DFFARX1 I_61070 (I1041775,I3563,I1041526,I1041491,);
not I_61071 (I1041806,I1041758);
nand I_61072 (I1041503,I1041569,I1041806);
DFFARX1 I_61073 (I1041758,I3563,I1041526,I1041846,);
not I_61074 (I1041854,I1041846);
not I_61075 (I1041871,I252389);
not I_61076 (I1041888,I252380);
nor I_61077 (I1041905,I1041888,I252368);
nor I_61078 (I1041518,I1041854,I1041905);
nor I_61079 (I1041936,I1041888,I252383);
and I_61080 (I1041953,I1041936,I252371);
or I_61081 (I1041970,I1041953,I252368);
DFFARX1 I_61082 (I1041970,I3563,I1041526,I1041996,);
nor I_61083 (I1041506,I1041996,I1041552);
not I_61084 (I1042018,I1041996);
and I_61085 (I1042035,I1042018,I1041552);
nor I_61086 (I1041500,I1041577,I1042035);
nand I_61087 (I1042066,I1042018,I1041628);
nor I_61088 (I1041494,I1041888,I1042066);
nand I_61089 (I1041497,I1042018,I1041806);
nand I_61090 (I1042111,I1041628,I252380);
nor I_61091 (I1041509,I1041871,I1042111);
not I_61092 (I1042172,I3570);
DFFARX1 I_61093 (I716219,I3563,I1042172,I1042198,);
DFFARX1 I_61094 (I716213,I3563,I1042172,I1042215,);
not I_61095 (I1042223,I1042215);
not I_61096 (I1042240,I716228);
nor I_61097 (I1042257,I1042240,I716213);
not I_61098 (I1042274,I716222);
nor I_61099 (I1042291,I1042257,I716231);
nor I_61100 (I1042308,I1042215,I1042291);
DFFARX1 I_61101 (I1042308,I3563,I1042172,I1042158,);
nor I_61102 (I1042339,I716231,I716213);
nand I_61103 (I1042356,I1042339,I716228);
DFFARX1 I_61104 (I1042356,I3563,I1042172,I1042161,);
nor I_61105 (I1042387,I1042274,I716231);
nand I_61106 (I1042404,I1042387,I716216);
nor I_61107 (I1042421,I1042198,I1042404);
DFFARX1 I_61108 (I1042421,I3563,I1042172,I1042137,);
not I_61109 (I1042452,I1042404);
nand I_61110 (I1042149,I1042215,I1042452);
DFFARX1 I_61111 (I1042404,I3563,I1042172,I1042492,);
not I_61112 (I1042500,I1042492);
not I_61113 (I1042517,I716231);
not I_61114 (I1042534,I716225);
nor I_61115 (I1042551,I1042534,I716222);
nor I_61116 (I1042164,I1042500,I1042551);
nor I_61117 (I1042582,I1042534,I716234);
and I_61118 (I1042599,I1042582,I716237);
or I_61119 (I1042616,I1042599,I716216);
DFFARX1 I_61120 (I1042616,I3563,I1042172,I1042642,);
nor I_61121 (I1042152,I1042642,I1042198);
not I_61122 (I1042664,I1042642);
and I_61123 (I1042681,I1042664,I1042198);
nor I_61124 (I1042146,I1042223,I1042681);
nand I_61125 (I1042712,I1042664,I1042274);
nor I_61126 (I1042140,I1042534,I1042712);
nand I_61127 (I1042143,I1042664,I1042452);
nand I_61128 (I1042757,I1042274,I716225);
nor I_61129 (I1042155,I1042517,I1042757);
not I_61130 (I1042818,I3570);
DFFARX1 I_61131 (I229169,I3563,I1042818,I1042844,);
DFFARX1 I_61132 (I229181,I3563,I1042818,I1042861,);
not I_61133 (I1042869,I1042861);
not I_61134 (I1042886,I229187);
nor I_61135 (I1042903,I1042886,I229172);
not I_61136 (I1042920,I229163);
nor I_61137 (I1042937,I1042903,I229184);
nor I_61138 (I1042954,I1042861,I1042937);
DFFARX1 I_61139 (I1042954,I3563,I1042818,I1042804,);
nor I_61140 (I1042985,I229184,I229172);
nand I_61141 (I1043002,I1042985,I229187);
DFFARX1 I_61142 (I1043002,I3563,I1042818,I1042807,);
nor I_61143 (I1043033,I1042920,I229184);
nand I_61144 (I1043050,I1043033,I229166);
nor I_61145 (I1043067,I1042844,I1043050);
DFFARX1 I_61146 (I1043067,I3563,I1042818,I1042783,);
not I_61147 (I1043098,I1043050);
nand I_61148 (I1042795,I1042861,I1043098);
DFFARX1 I_61149 (I1043050,I3563,I1042818,I1043138,);
not I_61150 (I1043146,I1043138);
not I_61151 (I1043163,I229184);
not I_61152 (I1043180,I229175);
nor I_61153 (I1043197,I1043180,I229163);
nor I_61154 (I1042810,I1043146,I1043197);
nor I_61155 (I1043228,I1043180,I229178);
and I_61156 (I1043245,I1043228,I229166);
or I_61157 (I1043262,I1043245,I229163);
DFFARX1 I_61158 (I1043262,I3563,I1042818,I1043288,);
nor I_61159 (I1042798,I1043288,I1042844);
not I_61160 (I1043310,I1043288);
and I_61161 (I1043327,I1043310,I1042844);
nor I_61162 (I1042792,I1042869,I1043327);
nand I_61163 (I1043358,I1043310,I1042920);
nor I_61164 (I1042786,I1043180,I1043358);
nand I_61165 (I1042789,I1043310,I1043098);
nand I_61166 (I1043403,I1042920,I229175);
nor I_61167 (I1042801,I1043163,I1043403);
not I_61168 (I1043464,I3570);
DFFARX1 I_61169 (I506184,I3563,I1043464,I1043490,);
DFFARX1 I_61170 (I506181,I3563,I1043464,I1043507,);
not I_61171 (I1043515,I1043507);
not I_61172 (I1043532,I506196);
nor I_61173 (I1043549,I1043532,I506199);
not I_61174 (I1043566,I506187);
nor I_61175 (I1043583,I1043549,I506193);
nor I_61176 (I1043600,I1043507,I1043583);
DFFARX1 I_61177 (I1043600,I3563,I1043464,I1043450,);
nor I_61178 (I1043631,I506193,I506199);
nand I_61179 (I1043648,I1043631,I506196);
DFFARX1 I_61180 (I1043648,I3563,I1043464,I1043453,);
nor I_61181 (I1043679,I1043566,I506193);
nand I_61182 (I1043696,I1043679,I506205);
nor I_61183 (I1043713,I1043490,I1043696);
DFFARX1 I_61184 (I1043713,I3563,I1043464,I1043429,);
not I_61185 (I1043744,I1043696);
nand I_61186 (I1043441,I1043507,I1043744);
DFFARX1 I_61187 (I1043696,I3563,I1043464,I1043784,);
not I_61188 (I1043792,I1043784);
not I_61189 (I1043809,I506193);
not I_61190 (I1043826,I506178);
nor I_61191 (I1043843,I1043826,I506187);
nor I_61192 (I1043456,I1043792,I1043843);
nor I_61193 (I1043874,I1043826,I506190);
and I_61194 (I1043891,I1043874,I506178);
or I_61195 (I1043908,I1043891,I506202);
DFFARX1 I_61196 (I1043908,I3563,I1043464,I1043934,);
nor I_61197 (I1043444,I1043934,I1043490);
not I_61198 (I1043956,I1043934);
and I_61199 (I1043973,I1043956,I1043490);
nor I_61200 (I1043438,I1043515,I1043973);
nand I_61201 (I1044004,I1043956,I1043566);
nor I_61202 (I1043432,I1043826,I1044004);
nand I_61203 (I1043435,I1043956,I1043744);
nand I_61204 (I1044049,I1043566,I506178);
nor I_61205 (I1043447,I1043809,I1044049);
not I_61206 (I1044110,I3570);
DFFARX1 I_61207 (I547729,I3563,I1044110,I1044136,);
DFFARX1 I_61208 (I547741,I3563,I1044110,I1044153,);
not I_61209 (I1044161,I1044153);
not I_61210 (I1044178,I547726);
nor I_61211 (I1044195,I1044178,I547744);
not I_61212 (I1044212,I547750);
nor I_61213 (I1044229,I1044195,I547732);
nor I_61214 (I1044246,I1044153,I1044229);
DFFARX1 I_61215 (I1044246,I3563,I1044110,I1044096,);
nor I_61216 (I1044277,I547732,I547744);
nand I_61217 (I1044294,I1044277,I547726);
DFFARX1 I_61218 (I1044294,I3563,I1044110,I1044099,);
nor I_61219 (I1044325,I1044212,I547732);
nand I_61220 (I1044342,I1044325,I547735);
nor I_61221 (I1044359,I1044136,I1044342);
DFFARX1 I_61222 (I1044359,I3563,I1044110,I1044075,);
not I_61223 (I1044390,I1044342);
nand I_61224 (I1044087,I1044153,I1044390);
DFFARX1 I_61225 (I1044342,I3563,I1044110,I1044430,);
not I_61226 (I1044438,I1044430);
not I_61227 (I1044455,I547732);
not I_61228 (I1044472,I547738);
nor I_61229 (I1044489,I1044472,I547750);
nor I_61230 (I1044102,I1044438,I1044489);
nor I_61231 (I1044520,I1044472,I547747);
and I_61232 (I1044537,I1044520,I547726);
or I_61233 (I1044554,I1044537,I547729);
DFFARX1 I_61234 (I1044554,I3563,I1044110,I1044580,);
nor I_61235 (I1044090,I1044580,I1044136);
not I_61236 (I1044602,I1044580);
and I_61237 (I1044619,I1044602,I1044136);
nor I_61238 (I1044084,I1044161,I1044619);
nand I_61239 (I1044650,I1044602,I1044212);
nor I_61240 (I1044078,I1044472,I1044650);
nand I_61241 (I1044081,I1044602,I1044390);
nand I_61242 (I1044695,I1044212,I547738);
nor I_61243 (I1044093,I1044455,I1044695);
not I_61244 (I1044756,I3570);
DFFARX1 I_61245 (I840574,I3563,I1044756,I1044782,);
DFFARX1 I_61246 (I840571,I3563,I1044756,I1044799,);
not I_61247 (I1044807,I1044799);
not I_61248 (I1044824,I840571);
nor I_61249 (I1044841,I1044824,I840574);
not I_61250 (I1044858,I840586);
nor I_61251 (I1044875,I1044841,I840580);
nor I_61252 (I1044892,I1044799,I1044875);
DFFARX1 I_61253 (I1044892,I3563,I1044756,I1044742,);
nor I_61254 (I1044923,I840580,I840574);
nand I_61255 (I1044940,I1044923,I840571);
DFFARX1 I_61256 (I1044940,I3563,I1044756,I1044745,);
nor I_61257 (I1044971,I1044858,I840580);
nand I_61258 (I1044988,I1044971,I840568);
nor I_61259 (I1045005,I1044782,I1044988);
DFFARX1 I_61260 (I1045005,I3563,I1044756,I1044721,);
not I_61261 (I1045036,I1044988);
nand I_61262 (I1044733,I1044799,I1045036);
DFFARX1 I_61263 (I1044988,I3563,I1044756,I1045076,);
not I_61264 (I1045084,I1045076);
not I_61265 (I1045101,I840580);
not I_61266 (I1045118,I840577);
nor I_61267 (I1045135,I1045118,I840586);
nor I_61268 (I1044748,I1045084,I1045135);
nor I_61269 (I1045166,I1045118,I840583);
and I_61270 (I1045183,I1045166,I840589);
or I_61271 (I1045200,I1045183,I840568);
DFFARX1 I_61272 (I1045200,I3563,I1044756,I1045226,);
nor I_61273 (I1044736,I1045226,I1044782);
not I_61274 (I1045248,I1045226);
and I_61275 (I1045265,I1045248,I1044782);
nor I_61276 (I1044730,I1044807,I1045265);
nand I_61277 (I1045296,I1045248,I1044858);
nor I_61278 (I1044724,I1045118,I1045296);
nand I_61279 (I1044727,I1045248,I1045036);
nand I_61280 (I1045341,I1044858,I840577);
nor I_61281 (I1044739,I1045101,I1045341);
not I_61282 (I1045402,I3570);
DFFARX1 I_61283 (I1116445,I3563,I1045402,I1045428,);
DFFARX1 I_61284 (I1116427,I3563,I1045402,I1045445,);
not I_61285 (I1045453,I1045445);
not I_61286 (I1045470,I1116436);
nor I_61287 (I1045487,I1045470,I1116448);
not I_61288 (I1045504,I1116430);
nor I_61289 (I1045521,I1045487,I1116439);
nor I_61290 (I1045538,I1045445,I1045521);
DFFARX1 I_61291 (I1045538,I3563,I1045402,I1045388,);
nor I_61292 (I1045569,I1116439,I1116448);
nand I_61293 (I1045586,I1045569,I1116436);
DFFARX1 I_61294 (I1045586,I3563,I1045402,I1045391,);
nor I_61295 (I1045617,I1045504,I1116439);
nand I_61296 (I1045634,I1045617,I1116451);
nor I_61297 (I1045651,I1045428,I1045634);
DFFARX1 I_61298 (I1045651,I3563,I1045402,I1045367,);
not I_61299 (I1045682,I1045634);
nand I_61300 (I1045379,I1045445,I1045682);
DFFARX1 I_61301 (I1045634,I3563,I1045402,I1045722,);
not I_61302 (I1045730,I1045722);
not I_61303 (I1045747,I1116439);
not I_61304 (I1045764,I1116427);
nor I_61305 (I1045781,I1045764,I1116430);
nor I_61306 (I1045394,I1045730,I1045781);
nor I_61307 (I1045812,I1045764,I1116433);
and I_61308 (I1045829,I1045812,I1116442);
or I_61309 (I1045846,I1045829,I1116430);
DFFARX1 I_61310 (I1045846,I3563,I1045402,I1045872,);
nor I_61311 (I1045382,I1045872,I1045428);
not I_61312 (I1045894,I1045872);
and I_61313 (I1045911,I1045894,I1045428);
nor I_61314 (I1045376,I1045453,I1045911);
nand I_61315 (I1045942,I1045894,I1045504);
nor I_61316 (I1045370,I1045764,I1045942);
nand I_61317 (I1045373,I1045894,I1045682);
nand I_61318 (I1045987,I1045504,I1116427);
nor I_61319 (I1045385,I1045747,I1045987);
not I_61320 (I1046048,I3570);
DFFARX1 I_61321 (I382333,I3563,I1046048,I1046074,);
DFFARX1 I_61322 (I382339,I3563,I1046048,I1046091,);
not I_61323 (I1046099,I1046091);
not I_61324 (I1046116,I382360);
nor I_61325 (I1046133,I1046116,I382348);
not I_61326 (I1046150,I382357);
nor I_61327 (I1046167,I1046133,I382342);
nor I_61328 (I1046184,I1046091,I1046167);
DFFARX1 I_61329 (I1046184,I3563,I1046048,I1046034,);
nor I_61330 (I1046215,I382342,I382348);
nand I_61331 (I1046232,I1046215,I382360);
DFFARX1 I_61332 (I1046232,I3563,I1046048,I1046037,);
nor I_61333 (I1046263,I1046150,I382342);
nand I_61334 (I1046280,I1046263,I382333);
nor I_61335 (I1046297,I1046074,I1046280);
DFFARX1 I_61336 (I1046297,I3563,I1046048,I1046013,);
not I_61337 (I1046328,I1046280);
nand I_61338 (I1046025,I1046091,I1046328);
DFFARX1 I_61339 (I1046280,I3563,I1046048,I1046368,);
not I_61340 (I1046376,I1046368);
not I_61341 (I1046393,I382342);
not I_61342 (I1046410,I382345);
nor I_61343 (I1046427,I1046410,I382357);
nor I_61344 (I1046040,I1046376,I1046427);
nor I_61345 (I1046458,I1046410,I382354);
and I_61346 (I1046475,I1046458,I382336);
or I_61347 (I1046492,I1046475,I382351);
DFFARX1 I_61348 (I1046492,I3563,I1046048,I1046518,);
nor I_61349 (I1046028,I1046518,I1046074);
not I_61350 (I1046540,I1046518);
and I_61351 (I1046557,I1046540,I1046074);
nor I_61352 (I1046022,I1046099,I1046557);
nand I_61353 (I1046588,I1046540,I1046150);
nor I_61354 (I1046016,I1046410,I1046588);
nand I_61355 (I1046019,I1046540,I1046328);
nand I_61356 (I1046633,I1046150,I382345);
nor I_61357 (I1046031,I1046393,I1046633);
not I_61358 (I1046688,I3570);
DFFARX1 I_61359 (I51395,I3563,I1046688,I1046714,);
DFFARX1 I_61360 (I1046714,I3563,I1046688,I1046731,);
not I_61361 (I1046680,I1046731);
not I_61362 (I1046753,I1046714);
DFFARX1 I_61363 (I51380,I3563,I1046688,I1046779,);
nand I_61364 (I1046787,I1046779,I51392);
not I_61365 (I1046804,I51392);
not I_61366 (I1046821,I51398);
nand I_61367 (I1046838,I51386,I51377);
and I_61368 (I1046855,I51386,I51377);
not I_61369 (I1046872,I51383);
nand I_61370 (I1046889,I1046872,I1046821);
nor I_61371 (I1046662,I1046889,I1046787);
nor I_61372 (I1046920,I1046804,I1046889);
nand I_61373 (I1046665,I1046855,I1046920);
not I_61374 (I1046951,I51389);
nor I_61375 (I1046968,I1046951,I51386);
nor I_61376 (I1046985,I1046968,I51383);
nor I_61377 (I1047002,I1046753,I1046985);
DFFARX1 I_61378 (I1047002,I3563,I1046688,I1046674,);
not I_61379 (I1047033,I1046968);
DFFARX1 I_61380 (I1047033,I3563,I1046688,I1046677,);
and I_61381 (I1046671,I1046779,I1046968);
nor I_61382 (I1047078,I1046951,I51377);
and I_61383 (I1047095,I1047078,I51401);
or I_61384 (I1047112,I1047095,I51380);
DFFARX1 I_61385 (I1047112,I3563,I1046688,I1047138,);
nor I_61386 (I1047146,I1047138,I1046872);
DFFARX1 I_61387 (I1047146,I3563,I1046688,I1046659,);
nand I_61388 (I1047177,I1047138,I1046779);
nand I_61389 (I1047194,I1046872,I1047177);
nor I_61390 (I1046668,I1047194,I1046838);
not I_61391 (I1047249,I3570);
DFFARX1 I_61392 (I766502,I3563,I1047249,I1047275,);
DFFARX1 I_61393 (I1047275,I3563,I1047249,I1047292,);
not I_61394 (I1047241,I1047292);
not I_61395 (I1047314,I1047275);
DFFARX1 I_61396 (I766514,I3563,I1047249,I1047340,);
nand I_61397 (I1047348,I1047340,I766523);
not I_61398 (I1047365,I766523);
not I_61399 (I1047382,I766505);
nand I_61400 (I1047399,I766508,I766499);
and I_61401 (I1047416,I766508,I766499);
not I_61402 (I1047433,I766517);
nand I_61403 (I1047450,I1047433,I1047382);
nor I_61404 (I1047223,I1047450,I1047348);
nor I_61405 (I1047481,I1047365,I1047450);
nand I_61406 (I1047226,I1047416,I1047481);
not I_61407 (I1047512,I766520);
nor I_61408 (I1047529,I1047512,I766508);
nor I_61409 (I1047546,I1047529,I766517);
nor I_61410 (I1047563,I1047314,I1047546);
DFFARX1 I_61411 (I1047563,I3563,I1047249,I1047235,);
not I_61412 (I1047594,I1047529);
DFFARX1 I_61413 (I1047594,I3563,I1047249,I1047238,);
and I_61414 (I1047232,I1047340,I1047529);
nor I_61415 (I1047639,I1047512,I766499);
and I_61416 (I1047656,I1047639,I766511);
or I_61417 (I1047673,I1047656,I766502);
DFFARX1 I_61418 (I1047673,I3563,I1047249,I1047699,);
nor I_61419 (I1047707,I1047699,I1047433);
DFFARX1 I_61420 (I1047707,I3563,I1047249,I1047220,);
nand I_61421 (I1047738,I1047699,I1047340);
nand I_61422 (I1047755,I1047433,I1047738);
nor I_61423 (I1047229,I1047755,I1047399);
not I_61424 (I1047810,I3570);
DFFARX1 I_61425 (I1404728,I3563,I1047810,I1047836,);
DFFARX1 I_61426 (I1047836,I3563,I1047810,I1047853,);
not I_61427 (I1047802,I1047853);
not I_61428 (I1047875,I1047836);
DFFARX1 I_61429 (I1404722,I3563,I1047810,I1047901,);
nand I_61430 (I1047909,I1047901,I1404713);
not I_61431 (I1047926,I1404713);
not I_61432 (I1047943,I1404740);
nand I_61433 (I1047960,I1404725,I1404734);
and I_61434 (I1047977,I1404725,I1404734);
not I_61435 (I1047994,I1404719);
nand I_61436 (I1048011,I1047994,I1047943);
nor I_61437 (I1047784,I1048011,I1047909);
nor I_61438 (I1048042,I1047926,I1048011);
nand I_61439 (I1047787,I1047977,I1048042);
not I_61440 (I1048073,I1404737);
nor I_61441 (I1048090,I1048073,I1404725);
nor I_61442 (I1048107,I1048090,I1404719);
nor I_61443 (I1048124,I1047875,I1048107);
DFFARX1 I_61444 (I1048124,I3563,I1047810,I1047796,);
not I_61445 (I1048155,I1048090);
DFFARX1 I_61446 (I1048155,I3563,I1047810,I1047799,);
and I_61447 (I1047793,I1047901,I1048090);
nor I_61448 (I1048200,I1048073,I1404731);
and I_61449 (I1048217,I1048200,I1404713);
or I_61450 (I1048234,I1048217,I1404716);
DFFARX1 I_61451 (I1048234,I3563,I1047810,I1048260,);
nor I_61452 (I1048268,I1048260,I1047994);
DFFARX1 I_61453 (I1048268,I3563,I1047810,I1047781,);
nand I_61454 (I1048299,I1048260,I1047901);
nand I_61455 (I1048316,I1047994,I1048299);
nor I_61456 (I1047790,I1048316,I1047960);
not I_61457 (I1048371,I3570);
DFFARX1 I_61458 (I899074,I3563,I1048371,I1048397,);
DFFARX1 I_61459 (I1048397,I3563,I1048371,I1048414,);
not I_61460 (I1048363,I1048414);
not I_61461 (I1048436,I1048397);
DFFARX1 I_61462 (I899071,I3563,I1048371,I1048462,);
nand I_61463 (I1048470,I1048462,I899086);
not I_61464 (I1048487,I899086);
not I_61465 (I1048504,I899083);
nand I_61466 (I1048521,I899080,I899068);
and I_61467 (I1048538,I899080,I899068);
not I_61468 (I1048555,I899065);
nand I_61469 (I1048572,I1048555,I1048504);
nor I_61470 (I1048345,I1048572,I1048470);
nor I_61471 (I1048603,I1048487,I1048572);
nand I_61472 (I1048348,I1048538,I1048603);
not I_61473 (I1048634,I899071);
nor I_61474 (I1048651,I1048634,I899080);
nor I_61475 (I1048668,I1048651,I899065);
nor I_61476 (I1048685,I1048436,I1048668);
DFFARX1 I_61477 (I1048685,I3563,I1048371,I1048357,);
not I_61478 (I1048716,I1048651);
DFFARX1 I_61479 (I1048716,I3563,I1048371,I1048360,);
and I_61480 (I1048354,I1048462,I1048651);
nor I_61481 (I1048761,I1048634,I899077);
and I_61482 (I1048778,I1048761,I899065);
or I_61483 (I1048795,I1048778,I899068);
DFFARX1 I_61484 (I1048795,I3563,I1048371,I1048821,);
nor I_61485 (I1048829,I1048821,I1048555);
DFFARX1 I_61486 (I1048829,I3563,I1048371,I1048342,);
nand I_61487 (I1048860,I1048821,I1048462);
nand I_61488 (I1048877,I1048555,I1048860);
nor I_61489 (I1048351,I1048877,I1048521);
not I_61490 (I1048932,I3570);
DFFARX1 I_61491 (I892750,I3563,I1048932,I1048958,);
DFFARX1 I_61492 (I1048958,I3563,I1048932,I1048975,);
not I_61493 (I1048924,I1048975);
not I_61494 (I1048997,I1048958);
DFFARX1 I_61495 (I892747,I3563,I1048932,I1049023,);
nand I_61496 (I1049031,I1049023,I892762);
not I_61497 (I1049048,I892762);
not I_61498 (I1049065,I892759);
nand I_61499 (I1049082,I892756,I892744);
and I_61500 (I1049099,I892756,I892744);
not I_61501 (I1049116,I892741);
nand I_61502 (I1049133,I1049116,I1049065);
nor I_61503 (I1048906,I1049133,I1049031);
nor I_61504 (I1049164,I1049048,I1049133);
nand I_61505 (I1048909,I1049099,I1049164);
not I_61506 (I1049195,I892747);
nor I_61507 (I1049212,I1049195,I892756);
nor I_61508 (I1049229,I1049212,I892741);
nor I_61509 (I1049246,I1048997,I1049229);
DFFARX1 I_61510 (I1049246,I3563,I1048932,I1048918,);
not I_61511 (I1049277,I1049212);
DFFARX1 I_61512 (I1049277,I3563,I1048932,I1048921,);
and I_61513 (I1048915,I1049023,I1049212);
nor I_61514 (I1049322,I1049195,I892753);
and I_61515 (I1049339,I1049322,I892741);
or I_61516 (I1049356,I1049339,I892744);
DFFARX1 I_61517 (I1049356,I3563,I1048932,I1049382,);
nor I_61518 (I1049390,I1049382,I1049116);
DFFARX1 I_61519 (I1049390,I3563,I1048932,I1048903,);
nand I_61520 (I1049421,I1049382,I1049023);
nand I_61521 (I1049438,I1049116,I1049421);
nor I_61522 (I1048912,I1049438,I1049082);
not I_61523 (I1049493,I3570);
DFFARX1 I_61524 (I64037,I3563,I1049493,I1049519,);
DFFARX1 I_61525 (I1049519,I3563,I1049493,I1049536,);
not I_61526 (I1049485,I1049536);
not I_61527 (I1049558,I1049519);
DFFARX1 I_61528 (I64025,I3563,I1049493,I1049584,);
nand I_61529 (I1049592,I1049584,I64040);
not I_61530 (I1049609,I64040);
not I_61531 (I1049626,I64028);
nand I_61532 (I1049643,I64049,I64043);
and I_61533 (I1049660,I64049,I64043);
not I_61534 (I1049677,I64031);
nand I_61535 (I1049694,I1049677,I1049626);
nor I_61536 (I1049467,I1049694,I1049592);
nor I_61537 (I1049725,I1049609,I1049694);
nand I_61538 (I1049470,I1049660,I1049725);
not I_61539 (I1049756,I64034);
nor I_61540 (I1049773,I1049756,I64049);
nor I_61541 (I1049790,I1049773,I64031);
nor I_61542 (I1049807,I1049558,I1049790);
DFFARX1 I_61543 (I1049807,I3563,I1049493,I1049479,);
not I_61544 (I1049838,I1049773);
DFFARX1 I_61545 (I1049838,I3563,I1049493,I1049482,);
and I_61546 (I1049476,I1049584,I1049773);
nor I_61547 (I1049883,I1049756,I64028);
and I_61548 (I1049900,I1049883,I64025);
or I_61549 (I1049917,I1049900,I64046);
DFFARX1 I_61550 (I1049917,I3563,I1049493,I1049943,);
nor I_61551 (I1049951,I1049943,I1049677);
DFFARX1 I_61552 (I1049951,I3563,I1049493,I1049464,);
nand I_61553 (I1049982,I1049943,I1049584);
nand I_61554 (I1049999,I1049677,I1049982);
nor I_61555 (I1049473,I1049999,I1049643);
not I_61556 (I1050054,I3570);
DFFARX1 I_61557 (I93022,I3563,I1050054,I1050080,);
DFFARX1 I_61558 (I1050080,I3563,I1050054,I1050097,);
not I_61559 (I1050046,I1050097);
not I_61560 (I1050119,I1050080);
DFFARX1 I_61561 (I93010,I3563,I1050054,I1050145,);
nand I_61562 (I1050153,I1050145,I93025);
not I_61563 (I1050170,I93025);
not I_61564 (I1050187,I93013);
nand I_61565 (I1050204,I93034,I93028);
and I_61566 (I1050221,I93034,I93028);
not I_61567 (I1050238,I93016);
nand I_61568 (I1050255,I1050238,I1050187);
nor I_61569 (I1050028,I1050255,I1050153);
nor I_61570 (I1050286,I1050170,I1050255);
nand I_61571 (I1050031,I1050221,I1050286);
not I_61572 (I1050317,I93019);
nor I_61573 (I1050334,I1050317,I93034);
nor I_61574 (I1050351,I1050334,I93016);
nor I_61575 (I1050368,I1050119,I1050351);
DFFARX1 I_61576 (I1050368,I3563,I1050054,I1050040,);
not I_61577 (I1050399,I1050334);
DFFARX1 I_61578 (I1050399,I3563,I1050054,I1050043,);
and I_61579 (I1050037,I1050145,I1050334);
nor I_61580 (I1050444,I1050317,I93013);
and I_61581 (I1050461,I1050444,I93010);
or I_61582 (I1050478,I1050461,I93031);
DFFARX1 I_61583 (I1050478,I3563,I1050054,I1050504,);
nor I_61584 (I1050512,I1050504,I1050238);
DFFARX1 I_61585 (I1050512,I3563,I1050054,I1050025,);
nand I_61586 (I1050543,I1050504,I1050145);
nand I_61587 (I1050560,I1050238,I1050543);
nor I_61588 (I1050034,I1050560,I1050204);
not I_61589 (I1050615,I3570);
DFFARX1 I_61590 (I1260015,I3563,I1050615,I1050641,);
DFFARX1 I_61591 (I1050641,I3563,I1050615,I1050658,);
not I_61592 (I1050607,I1050658);
not I_61593 (I1050680,I1050641);
DFFARX1 I_61594 (I1260021,I3563,I1050615,I1050706,);
nand I_61595 (I1050714,I1050706,I1260030);
not I_61596 (I1050731,I1260030);
not I_61597 (I1050748,I1260009);
nand I_61598 (I1050765,I1260012,I1260012);
and I_61599 (I1050782,I1260012,I1260012);
not I_61600 (I1050799,I1260024);
nand I_61601 (I1050816,I1050799,I1050748);
nor I_61602 (I1050589,I1050816,I1050714);
nor I_61603 (I1050847,I1050731,I1050816);
nand I_61604 (I1050592,I1050782,I1050847);
not I_61605 (I1050878,I1260018);
nor I_61606 (I1050895,I1050878,I1260012);
nor I_61607 (I1050912,I1050895,I1260024);
nor I_61608 (I1050929,I1050680,I1050912);
DFFARX1 I_61609 (I1050929,I3563,I1050615,I1050601,);
not I_61610 (I1050960,I1050895);
DFFARX1 I_61611 (I1050960,I3563,I1050615,I1050604,);
and I_61612 (I1050598,I1050706,I1050895);
nor I_61613 (I1051005,I1050878,I1260033);
and I_61614 (I1051022,I1051005,I1260009);
or I_61615 (I1051039,I1051022,I1260027);
DFFARX1 I_61616 (I1051039,I3563,I1050615,I1051065,);
nor I_61617 (I1051073,I1051065,I1050799);
DFFARX1 I_61618 (I1051073,I3563,I1050615,I1050586,);
nand I_61619 (I1051104,I1051065,I1050706);
nand I_61620 (I1051121,I1050799,I1051104);
nor I_61621 (I1050595,I1051121,I1050765);
not I_61622 (I1051176,I3570);
DFFARX1 I_61623 (I146249,I3563,I1051176,I1051202,);
DFFARX1 I_61624 (I1051202,I3563,I1051176,I1051219,);
not I_61625 (I1051168,I1051219);
not I_61626 (I1051241,I1051202);
DFFARX1 I_61627 (I146237,I3563,I1051176,I1051267,);
nand I_61628 (I1051275,I1051267,I146252);
not I_61629 (I1051292,I146252);
not I_61630 (I1051309,I146240);
nand I_61631 (I1051326,I146261,I146255);
and I_61632 (I1051343,I146261,I146255);
not I_61633 (I1051360,I146243);
nand I_61634 (I1051377,I1051360,I1051309);
nor I_61635 (I1051150,I1051377,I1051275);
nor I_61636 (I1051408,I1051292,I1051377);
nand I_61637 (I1051153,I1051343,I1051408);
not I_61638 (I1051439,I146246);
nor I_61639 (I1051456,I1051439,I146261);
nor I_61640 (I1051473,I1051456,I146243);
nor I_61641 (I1051490,I1051241,I1051473);
DFFARX1 I_61642 (I1051490,I3563,I1051176,I1051162,);
not I_61643 (I1051521,I1051456);
DFFARX1 I_61644 (I1051521,I3563,I1051176,I1051165,);
and I_61645 (I1051159,I1051267,I1051456);
nor I_61646 (I1051566,I1051439,I146240);
and I_61647 (I1051583,I1051566,I146237);
or I_61648 (I1051600,I1051583,I146258);
DFFARX1 I_61649 (I1051600,I3563,I1051176,I1051626,);
nor I_61650 (I1051634,I1051626,I1051360);
DFFARX1 I_61651 (I1051634,I3563,I1051176,I1051147,);
nand I_61652 (I1051665,I1051626,I1051267);
nand I_61653 (I1051682,I1051360,I1051665);
nor I_61654 (I1051156,I1051682,I1051326);
not I_61655 (I1051737,I3570);
DFFARX1 I_61656 (I971077,I3563,I1051737,I1051763,);
DFFARX1 I_61657 (I1051763,I3563,I1051737,I1051780,);
not I_61658 (I1051729,I1051780);
not I_61659 (I1051802,I1051763);
DFFARX1 I_61660 (I971104,I3563,I1051737,I1051828,);
nand I_61661 (I1051836,I1051828,I971095);
not I_61662 (I1051853,I971095);
not I_61663 (I1051870,I971077);
nand I_61664 (I1051887,I971089,I971092);
and I_61665 (I1051904,I971089,I971092);
not I_61666 (I1051921,I971101);
nand I_61667 (I1051938,I1051921,I1051870);
nor I_61668 (I1051711,I1051938,I1051836);
nor I_61669 (I1051969,I1051853,I1051938);
nand I_61670 (I1051714,I1051904,I1051969);
not I_61671 (I1052000,I971086);
nor I_61672 (I1052017,I1052000,I971089);
nor I_61673 (I1052034,I1052017,I971101);
nor I_61674 (I1052051,I1051802,I1052034);
DFFARX1 I_61675 (I1052051,I3563,I1051737,I1051723,);
not I_61676 (I1052082,I1052017);
DFFARX1 I_61677 (I1052082,I3563,I1051737,I1051726,);
and I_61678 (I1051720,I1051828,I1052017);
nor I_61679 (I1052127,I1052000,I971080);
and I_61680 (I1052144,I1052127,I971083);
or I_61681 (I1052161,I1052144,I971098);
DFFARX1 I_61682 (I1052161,I3563,I1051737,I1052187,);
nor I_61683 (I1052195,I1052187,I1051921);
DFFARX1 I_61684 (I1052195,I3563,I1051737,I1051708,);
nand I_61685 (I1052226,I1052187,I1051828);
nand I_61686 (I1052243,I1051921,I1052226);
nor I_61687 (I1051717,I1052243,I1051887);
not I_61688 (I1052298,I3570);
DFFARX1 I_61689 (I1286127,I3563,I1052298,I1052324,);
DFFARX1 I_61690 (I1052324,I3563,I1052298,I1052341,);
not I_61691 (I1052290,I1052341);
not I_61692 (I1052363,I1052324);
DFFARX1 I_61693 (I1286133,I3563,I1052298,I1052389,);
nand I_61694 (I1052397,I1052389,I1286142);
not I_61695 (I1052414,I1286142);
not I_61696 (I1052431,I1286121);
nand I_61697 (I1052448,I1286124,I1286124);
and I_61698 (I1052465,I1286124,I1286124);
not I_61699 (I1052482,I1286136);
nand I_61700 (I1052499,I1052482,I1052431);
nor I_61701 (I1052272,I1052499,I1052397);
nor I_61702 (I1052530,I1052414,I1052499);
nand I_61703 (I1052275,I1052465,I1052530);
not I_61704 (I1052561,I1286130);
nor I_61705 (I1052578,I1052561,I1286124);
nor I_61706 (I1052595,I1052578,I1286136);
nor I_61707 (I1052612,I1052363,I1052595);
DFFARX1 I_61708 (I1052612,I3563,I1052298,I1052284,);
not I_61709 (I1052643,I1052578);
DFFARX1 I_61710 (I1052643,I3563,I1052298,I1052287,);
and I_61711 (I1052281,I1052389,I1052578);
nor I_61712 (I1052688,I1052561,I1286145);
and I_61713 (I1052705,I1052688,I1286121);
or I_61714 (I1052722,I1052705,I1286139);
DFFARX1 I_61715 (I1052722,I3563,I1052298,I1052748,);
nor I_61716 (I1052756,I1052748,I1052482);
DFFARX1 I_61717 (I1052756,I3563,I1052298,I1052269,);
nand I_61718 (I1052787,I1052748,I1052389);
nand I_61719 (I1052804,I1052482,I1052787);
nor I_61720 (I1052278,I1052804,I1052448);
not I_61721 (I1052859,I3570);
DFFARX1 I_61722 (I1181756,I3563,I1052859,I1052885,);
DFFARX1 I_61723 (I1052885,I3563,I1052859,I1052902,);
not I_61724 (I1052851,I1052902);
not I_61725 (I1052924,I1052885);
DFFARX1 I_61726 (I1181747,I3563,I1052859,I1052950,);
nand I_61727 (I1052958,I1052950,I1181744);
not I_61728 (I1052975,I1181744);
not I_61729 (I1052992,I1181753);
nand I_61730 (I1053009,I1181762,I1181744);
and I_61731 (I1053026,I1181762,I1181744);
not I_61732 (I1053043,I1181741);
nand I_61733 (I1053060,I1053043,I1052992);
nor I_61734 (I1052833,I1053060,I1052958);
nor I_61735 (I1053091,I1052975,I1053060);
nand I_61736 (I1052836,I1053026,I1053091);
not I_61737 (I1053122,I1181750);
nor I_61738 (I1053139,I1053122,I1181762);
nor I_61739 (I1053156,I1053139,I1181741);
nor I_61740 (I1053173,I1052924,I1053156);
DFFARX1 I_61741 (I1053173,I3563,I1052859,I1052845,);
not I_61742 (I1053204,I1053139);
DFFARX1 I_61743 (I1053204,I3563,I1052859,I1052848,);
and I_61744 (I1052842,I1052950,I1053139);
nor I_61745 (I1053249,I1053122,I1181765);
and I_61746 (I1053266,I1053249,I1181741);
or I_61747 (I1053283,I1053266,I1181759);
DFFARX1 I_61748 (I1053283,I3563,I1052859,I1053309,);
nor I_61749 (I1053317,I1053309,I1053043);
DFFARX1 I_61750 (I1053317,I3563,I1052859,I1052830,);
nand I_61751 (I1053348,I1053309,I1052950);
nand I_61752 (I1053365,I1053043,I1053348);
nor I_61753 (I1052839,I1053365,I1053009);
not I_61754 (I1053420,I3570);
DFFARX1 I_61755 (I1111818,I3563,I1053420,I1053446,);
DFFARX1 I_61756 (I1053446,I3563,I1053420,I1053463,);
not I_61757 (I1053412,I1053463);
not I_61758 (I1053485,I1053446);
DFFARX1 I_61759 (I1111809,I3563,I1053420,I1053511,);
nand I_61760 (I1053519,I1053511,I1111806);
not I_61761 (I1053536,I1111806);
not I_61762 (I1053553,I1111815);
nand I_61763 (I1053570,I1111824,I1111806);
and I_61764 (I1053587,I1111824,I1111806);
not I_61765 (I1053604,I1111803);
nand I_61766 (I1053621,I1053604,I1053553);
nor I_61767 (I1053394,I1053621,I1053519);
nor I_61768 (I1053652,I1053536,I1053621);
nand I_61769 (I1053397,I1053587,I1053652);
not I_61770 (I1053683,I1111812);
nor I_61771 (I1053700,I1053683,I1111824);
nor I_61772 (I1053717,I1053700,I1111803);
nor I_61773 (I1053734,I1053485,I1053717);
DFFARX1 I_61774 (I1053734,I3563,I1053420,I1053406,);
not I_61775 (I1053765,I1053700);
DFFARX1 I_61776 (I1053765,I3563,I1053420,I1053409,);
and I_61777 (I1053403,I1053511,I1053700);
nor I_61778 (I1053810,I1053683,I1111827);
and I_61779 (I1053827,I1053810,I1111803);
or I_61780 (I1053844,I1053827,I1111821);
DFFARX1 I_61781 (I1053844,I3563,I1053420,I1053870,);
nor I_61782 (I1053878,I1053870,I1053604);
DFFARX1 I_61783 (I1053878,I3563,I1053420,I1053391,);
nand I_61784 (I1053909,I1053870,I1053511);
nand I_61785 (I1053926,I1053604,I1053909);
nor I_61786 (I1053400,I1053926,I1053570);
not I_61787 (I1053981,I3570);
DFFARX1 I_61788 (I233926,I3563,I1053981,I1054007,);
DFFARX1 I_61789 (I1054007,I3563,I1053981,I1054024,);
not I_61790 (I1053973,I1054024);
not I_61791 (I1054046,I1054007);
DFFARX1 I_61792 (I233941,I3563,I1053981,I1054072,);
nand I_61793 (I1054080,I1054072,I233923);
not I_61794 (I1054097,I233923);
not I_61795 (I1054114,I233932);
nand I_61796 (I1054131,I233938,I233929);
and I_61797 (I1054148,I233938,I233929);
not I_61798 (I1054165,I233926);
nand I_61799 (I1054182,I1054165,I1054114);
nor I_61800 (I1053955,I1054182,I1054080);
nor I_61801 (I1054213,I1054097,I1054182);
nand I_61802 (I1053958,I1054148,I1054213);
not I_61803 (I1054244,I233923);
nor I_61804 (I1054261,I1054244,I233938);
nor I_61805 (I1054278,I1054261,I233926);
nor I_61806 (I1054295,I1054046,I1054278);
DFFARX1 I_61807 (I1054295,I3563,I1053981,I1053967,);
not I_61808 (I1054326,I1054261);
DFFARX1 I_61809 (I1054326,I3563,I1053981,I1053970,);
and I_61810 (I1053964,I1054072,I1054261);
nor I_61811 (I1054371,I1054244,I233947);
and I_61812 (I1054388,I1054371,I233944);
or I_61813 (I1054405,I1054388,I233935);
DFFARX1 I_61814 (I1054405,I3563,I1053981,I1054431,);
nor I_61815 (I1054439,I1054431,I1054165);
DFFARX1 I_61816 (I1054439,I3563,I1053981,I1053952,);
nand I_61817 (I1054470,I1054431,I1054072);
nand I_61818 (I1054487,I1054165,I1054470);
nor I_61819 (I1053961,I1054487,I1054131);
not I_61820 (I1054542,I3570);
DFFARX1 I_61821 (I556669,I3563,I1054542,I1054568,);
DFFARX1 I_61822 (I1054568,I3563,I1054542,I1054585,);
not I_61823 (I1054534,I1054585);
not I_61824 (I1054607,I1054568);
DFFARX1 I_61825 (I556666,I3563,I1054542,I1054633,);
nand I_61826 (I1054641,I1054633,I556660);
not I_61827 (I1054658,I556660);
not I_61828 (I1054675,I556672);
nand I_61829 (I1054692,I556675,I556654);
and I_61830 (I1054709,I556675,I556654);
not I_61831 (I1054726,I556651);
nand I_61832 (I1054743,I1054726,I1054675);
nor I_61833 (I1054516,I1054743,I1054641);
nor I_61834 (I1054774,I1054658,I1054743);
nand I_61835 (I1054519,I1054709,I1054774);
not I_61836 (I1054805,I556657);
nor I_61837 (I1054822,I1054805,I556675);
nor I_61838 (I1054839,I1054822,I556651);
nor I_61839 (I1054856,I1054607,I1054839);
DFFARX1 I_61840 (I1054856,I3563,I1054542,I1054528,);
not I_61841 (I1054887,I1054822);
DFFARX1 I_61842 (I1054887,I3563,I1054542,I1054531,);
and I_61843 (I1054525,I1054633,I1054822);
nor I_61844 (I1054932,I1054805,I556651);
and I_61845 (I1054949,I1054932,I556663);
or I_61846 (I1054966,I1054949,I556654);
DFFARX1 I_61847 (I1054966,I3563,I1054542,I1054992,);
nor I_61848 (I1055000,I1054992,I1054726);
DFFARX1 I_61849 (I1055000,I3563,I1054542,I1054513,);
nand I_61850 (I1055031,I1054992,I1054633);
nand I_61851 (I1055048,I1054726,I1055031);
nor I_61852 (I1054522,I1055048,I1054692);
not I_61853 (I1055103,I3570);
DFFARX1 I_61854 (I534654,I3563,I1055103,I1055129,);
DFFARX1 I_61855 (I1055129,I3563,I1055103,I1055146,);
not I_61856 (I1055095,I1055146);
not I_61857 (I1055168,I1055129);
DFFARX1 I_61858 (I534651,I3563,I1055103,I1055194,);
nand I_61859 (I1055202,I1055194,I534645);
not I_61860 (I1055219,I534645);
not I_61861 (I1055236,I534657);
nand I_61862 (I1055253,I534660,I534639);
and I_61863 (I1055270,I534660,I534639);
not I_61864 (I1055287,I534636);
nand I_61865 (I1055304,I1055287,I1055236);
nor I_61866 (I1055077,I1055304,I1055202);
nor I_61867 (I1055335,I1055219,I1055304);
nand I_61868 (I1055080,I1055270,I1055335);
not I_61869 (I1055366,I534642);
nor I_61870 (I1055383,I1055366,I534660);
nor I_61871 (I1055400,I1055383,I534636);
nor I_61872 (I1055417,I1055168,I1055400);
DFFARX1 I_61873 (I1055417,I3563,I1055103,I1055089,);
not I_61874 (I1055448,I1055383);
DFFARX1 I_61875 (I1055448,I3563,I1055103,I1055092,);
and I_61876 (I1055086,I1055194,I1055383);
nor I_61877 (I1055493,I1055366,I534636);
and I_61878 (I1055510,I1055493,I534648);
or I_61879 (I1055527,I1055510,I534639);
DFFARX1 I_61880 (I1055527,I3563,I1055103,I1055553,);
nor I_61881 (I1055561,I1055553,I1055287);
DFFARX1 I_61882 (I1055561,I3563,I1055103,I1055074,);
nand I_61883 (I1055592,I1055553,I1055194);
nand I_61884 (I1055609,I1055287,I1055592);
nor I_61885 (I1055083,I1055609,I1055253);
not I_61886 (I1055664,I3570);
DFFARX1 I_61887 (I364963,I3563,I1055664,I1055690,);
DFFARX1 I_61888 (I1055690,I3563,I1055664,I1055707,);
not I_61889 (I1055656,I1055707);
not I_61890 (I1055729,I1055690);
DFFARX1 I_61891 (I364960,I3563,I1055664,I1055755,);
nand I_61892 (I1055763,I1055755,I364954);
not I_61893 (I1055780,I364954);
not I_61894 (I1055797,I364951);
nand I_61895 (I1055814,I364945,I364942);
and I_61896 (I1055831,I364945,I364942);
not I_61897 (I1055848,I364957);
nand I_61898 (I1055865,I1055848,I1055797);
nor I_61899 (I1055638,I1055865,I1055763);
nor I_61900 (I1055896,I1055780,I1055865);
nand I_61901 (I1055641,I1055831,I1055896);
not I_61902 (I1055927,I364969);
nor I_61903 (I1055944,I1055927,I364945);
nor I_61904 (I1055961,I1055944,I364957);
nor I_61905 (I1055978,I1055729,I1055961);
DFFARX1 I_61906 (I1055978,I3563,I1055664,I1055650,);
not I_61907 (I1056009,I1055944);
DFFARX1 I_61908 (I1056009,I3563,I1055664,I1055653,);
and I_61909 (I1055647,I1055755,I1055944);
nor I_61910 (I1056054,I1055927,I364966);
and I_61911 (I1056071,I1056054,I364942);
or I_61912 (I1056088,I1056071,I364948);
DFFARX1 I_61913 (I1056088,I3563,I1055664,I1056114,);
nor I_61914 (I1056122,I1056114,I1055848);
DFFARX1 I_61915 (I1056122,I3563,I1055664,I1055635,);
nand I_61916 (I1056153,I1056114,I1055755);
nand I_61917 (I1056170,I1055848,I1056153);
nor I_61918 (I1055644,I1056170,I1055814);
not I_61919 (I1056225,I3570);
DFFARX1 I_61920 (I440922,I3563,I1056225,I1056251,);
DFFARX1 I_61921 (I1056251,I3563,I1056225,I1056268,);
not I_61922 (I1056217,I1056268);
not I_61923 (I1056290,I1056251);
DFFARX1 I_61924 (I440910,I3563,I1056225,I1056316,);
nand I_61925 (I1056324,I1056316,I440916);
not I_61926 (I1056341,I440916);
not I_61927 (I1056358,I440913);
nand I_61928 (I1056375,I440901,I440898);
and I_61929 (I1056392,I440901,I440898);
not I_61930 (I1056409,I440925);
nand I_61931 (I1056426,I1056409,I1056358);
nor I_61932 (I1056199,I1056426,I1056324);
nor I_61933 (I1056457,I1056341,I1056426);
nand I_61934 (I1056202,I1056392,I1056457);
not I_61935 (I1056488,I440898);
nor I_61936 (I1056505,I1056488,I440901);
nor I_61937 (I1056522,I1056505,I440925);
nor I_61938 (I1056539,I1056290,I1056522);
DFFARX1 I_61939 (I1056539,I3563,I1056225,I1056211,);
not I_61940 (I1056570,I1056505);
DFFARX1 I_61941 (I1056570,I3563,I1056225,I1056214,);
and I_61942 (I1056208,I1056316,I1056505);
nor I_61943 (I1056615,I1056488,I440907);
and I_61944 (I1056632,I1056615,I440904);
or I_61945 (I1056649,I1056632,I440919);
DFFARX1 I_61946 (I1056649,I3563,I1056225,I1056675,);
nor I_61947 (I1056683,I1056675,I1056409);
DFFARX1 I_61948 (I1056683,I3563,I1056225,I1056196,);
nand I_61949 (I1056714,I1056675,I1056316);
nand I_61950 (I1056731,I1056409,I1056714);
nor I_61951 (I1056205,I1056731,I1056375);
not I_61952 (I1056786,I3570);
DFFARX1 I_61953 (I954927,I3563,I1056786,I1056812,);
DFFARX1 I_61954 (I1056812,I3563,I1056786,I1056829,);
not I_61955 (I1056778,I1056829);
not I_61956 (I1056851,I1056812);
DFFARX1 I_61957 (I954954,I3563,I1056786,I1056877,);
nand I_61958 (I1056885,I1056877,I954945);
not I_61959 (I1056902,I954945);
not I_61960 (I1056919,I954927);
nand I_61961 (I1056936,I954939,I954942);
and I_61962 (I1056953,I954939,I954942);
not I_61963 (I1056970,I954951);
nand I_61964 (I1056987,I1056970,I1056919);
nor I_61965 (I1056760,I1056987,I1056885);
nor I_61966 (I1057018,I1056902,I1056987);
nand I_61967 (I1056763,I1056953,I1057018);
not I_61968 (I1057049,I954936);
nor I_61969 (I1057066,I1057049,I954939);
nor I_61970 (I1057083,I1057066,I954951);
nor I_61971 (I1057100,I1056851,I1057083);
DFFARX1 I_61972 (I1057100,I3563,I1056786,I1056772,);
not I_61973 (I1057131,I1057066);
DFFARX1 I_61974 (I1057131,I3563,I1056786,I1056775,);
and I_61975 (I1056769,I1056877,I1057066);
nor I_61976 (I1057176,I1057049,I954930);
and I_61977 (I1057193,I1057176,I954933);
or I_61978 (I1057210,I1057193,I954948);
DFFARX1 I_61979 (I1057210,I3563,I1056786,I1057236,);
nor I_61980 (I1057244,I1057236,I1056970);
DFFARX1 I_61981 (I1057244,I3563,I1056786,I1056757,);
nand I_61982 (I1057275,I1057236,I1056877);
nand I_61983 (I1057292,I1056970,I1057275);
nor I_61984 (I1056766,I1057292,I1056936);
not I_61985 (I1057347,I3570);
DFFARX1 I_61986 (I437114,I3563,I1057347,I1057373,);
DFFARX1 I_61987 (I1057373,I3563,I1057347,I1057390,);
not I_61988 (I1057339,I1057390);
not I_61989 (I1057412,I1057373);
DFFARX1 I_61990 (I437102,I3563,I1057347,I1057438,);
nand I_61991 (I1057446,I1057438,I437108);
not I_61992 (I1057463,I437108);
not I_61993 (I1057480,I437105);
nand I_61994 (I1057497,I437093,I437090);
and I_61995 (I1057514,I437093,I437090);
not I_61996 (I1057531,I437117);
nand I_61997 (I1057548,I1057531,I1057480);
nor I_61998 (I1057321,I1057548,I1057446);
nor I_61999 (I1057579,I1057463,I1057548);
nand I_62000 (I1057324,I1057514,I1057579);
not I_62001 (I1057610,I437090);
nor I_62002 (I1057627,I1057610,I437093);
nor I_62003 (I1057644,I1057627,I437117);
nor I_62004 (I1057661,I1057412,I1057644);
DFFARX1 I_62005 (I1057661,I3563,I1057347,I1057333,);
not I_62006 (I1057692,I1057627);
DFFARX1 I_62007 (I1057692,I3563,I1057347,I1057336,);
and I_62008 (I1057330,I1057438,I1057627);
nor I_62009 (I1057737,I1057610,I437099);
and I_62010 (I1057754,I1057737,I437096);
or I_62011 (I1057771,I1057754,I437111);
DFFARX1 I_62012 (I1057771,I3563,I1057347,I1057797,);
nor I_62013 (I1057805,I1057797,I1057531);
DFFARX1 I_62014 (I1057805,I3563,I1057347,I1057318,);
nand I_62015 (I1057836,I1057797,I1057438);
nand I_62016 (I1057853,I1057531,I1057836);
nor I_62017 (I1057327,I1057853,I1057497);
not I_62018 (I1057908,I3570);
DFFARX1 I_62019 (I48760,I3563,I1057908,I1057934,);
DFFARX1 I_62020 (I1057934,I3563,I1057908,I1057951,);
not I_62021 (I1057900,I1057951);
not I_62022 (I1057973,I1057934);
DFFARX1 I_62023 (I48745,I3563,I1057908,I1057999,);
nand I_62024 (I1058007,I1057999,I48757);
not I_62025 (I1058024,I48757);
not I_62026 (I1058041,I48763);
nand I_62027 (I1058058,I48751,I48742);
and I_62028 (I1058075,I48751,I48742);
not I_62029 (I1058092,I48748);
nand I_62030 (I1058109,I1058092,I1058041);
nor I_62031 (I1057882,I1058109,I1058007);
nor I_62032 (I1058140,I1058024,I1058109);
nand I_62033 (I1057885,I1058075,I1058140);
not I_62034 (I1058171,I48754);
nor I_62035 (I1058188,I1058171,I48751);
nor I_62036 (I1058205,I1058188,I48748);
nor I_62037 (I1058222,I1057973,I1058205);
DFFARX1 I_62038 (I1058222,I3563,I1057908,I1057894,);
not I_62039 (I1058253,I1058188);
DFFARX1 I_62040 (I1058253,I3563,I1057908,I1057897,);
and I_62041 (I1057891,I1057999,I1058188);
nor I_62042 (I1058298,I1058171,I48742);
and I_62043 (I1058315,I1058298,I48766);
or I_62044 (I1058332,I1058315,I48745);
DFFARX1 I_62045 (I1058332,I3563,I1057908,I1058358,);
nor I_62046 (I1058366,I1058358,I1058092);
DFFARX1 I_62047 (I1058366,I3563,I1057908,I1057879,);
nand I_62048 (I1058397,I1058358,I1057999);
nand I_62049 (I1058414,I1058092,I1058397);
nor I_62050 (I1057888,I1058414,I1058058);
not I_62051 (I1058469,I3570);
DFFARX1 I_62052 (I651477,I3563,I1058469,I1058495,);
DFFARX1 I_62053 (I1058495,I3563,I1058469,I1058512,);
not I_62054 (I1058461,I1058512);
not I_62055 (I1058534,I1058495);
DFFARX1 I_62056 (I651492,I3563,I1058469,I1058560,);
nand I_62057 (I1058568,I1058560,I651483);
not I_62058 (I1058585,I651483);
not I_62059 (I1058602,I651489);
nand I_62060 (I1058619,I651486,I651495);
and I_62061 (I1058636,I651486,I651495);
not I_62062 (I1058653,I651480);
nand I_62063 (I1058670,I1058653,I1058602);
nor I_62064 (I1058443,I1058670,I1058568);
nor I_62065 (I1058701,I1058585,I1058670);
nand I_62066 (I1058446,I1058636,I1058701);
not I_62067 (I1058732,I651477);
nor I_62068 (I1058749,I1058732,I651486);
nor I_62069 (I1058766,I1058749,I651480);
nor I_62070 (I1058783,I1058534,I1058766);
DFFARX1 I_62071 (I1058783,I3563,I1058469,I1058455,);
not I_62072 (I1058814,I1058749);
DFFARX1 I_62073 (I1058814,I3563,I1058469,I1058458,);
and I_62074 (I1058452,I1058560,I1058749);
nor I_62075 (I1058859,I1058732,I651501);
and I_62076 (I1058876,I1058859,I651480);
or I_62077 (I1058893,I1058876,I651498);
DFFARX1 I_62078 (I1058893,I3563,I1058469,I1058919,);
nor I_62079 (I1058927,I1058919,I1058653);
DFFARX1 I_62080 (I1058927,I3563,I1058469,I1058440,);
nand I_62081 (I1058958,I1058919,I1058560);
nand I_62082 (I1058975,I1058653,I1058958);
nor I_62083 (I1058449,I1058975,I1058619);
not I_62084 (I1059030,I3570);
DFFARX1 I_62085 (I392894,I3563,I1059030,I1059056,);
DFFARX1 I_62086 (I1059056,I3563,I1059030,I1059073,);
not I_62087 (I1059022,I1059073);
not I_62088 (I1059095,I1059056);
DFFARX1 I_62089 (I392891,I3563,I1059030,I1059121,);
nand I_62090 (I1059129,I1059121,I392885);
not I_62091 (I1059146,I392885);
not I_62092 (I1059163,I392882);
nand I_62093 (I1059180,I392876,I392873);
and I_62094 (I1059197,I392876,I392873);
not I_62095 (I1059214,I392888);
nand I_62096 (I1059231,I1059214,I1059163);
nor I_62097 (I1059004,I1059231,I1059129);
nor I_62098 (I1059262,I1059146,I1059231);
nand I_62099 (I1059007,I1059197,I1059262);
not I_62100 (I1059293,I392900);
nor I_62101 (I1059310,I1059293,I392876);
nor I_62102 (I1059327,I1059310,I392888);
nor I_62103 (I1059344,I1059095,I1059327);
DFFARX1 I_62104 (I1059344,I3563,I1059030,I1059016,);
not I_62105 (I1059375,I1059310);
DFFARX1 I_62106 (I1059375,I3563,I1059030,I1059019,);
and I_62107 (I1059013,I1059121,I1059310);
nor I_62108 (I1059420,I1059293,I392897);
and I_62109 (I1059437,I1059420,I392873);
or I_62110 (I1059454,I1059437,I392879);
DFFARX1 I_62111 (I1059454,I3563,I1059030,I1059480,);
nor I_62112 (I1059488,I1059480,I1059214);
DFFARX1 I_62113 (I1059488,I3563,I1059030,I1059001,);
nand I_62114 (I1059519,I1059480,I1059121);
nand I_62115 (I1059536,I1059214,I1059519);
nor I_62116 (I1059010,I1059536,I1059180);
not I_62117 (I1059591,I3570);
DFFARX1 I_62118 (I1332733,I3563,I1059591,I1059617,);
DFFARX1 I_62119 (I1059617,I3563,I1059591,I1059634,);
not I_62120 (I1059583,I1059634);
not I_62121 (I1059656,I1059617);
DFFARX1 I_62122 (I1332727,I3563,I1059591,I1059682,);
nand I_62123 (I1059690,I1059682,I1332718);
not I_62124 (I1059707,I1332718);
not I_62125 (I1059724,I1332745);
nand I_62126 (I1059741,I1332730,I1332739);
and I_62127 (I1059758,I1332730,I1332739);
not I_62128 (I1059775,I1332724);
nand I_62129 (I1059792,I1059775,I1059724);
nor I_62130 (I1059565,I1059792,I1059690);
nor I_62131 (I1059823,I1059707,I1059792);
nand I_62132 (I1059568,I1059758,I1059823);
not I_62133 (I1059854,I1332742);
nor I_62134 (I1059871,I1059854,I1332730);
nor I_62135 (I1059888,I1059871,I1332724);
nor I_62136 (I1059905,I1059656,I1059888);
DFFARX1 I_62137 (I1059905,I3563,I1059591,I1059577,);
not I_62138 (I1059936,I1059871);
DFFARX1 I_62139 (I1059936,I3563,I1059591,I1059580,);
and I_62140 (I1059574,I1059682,I1059871);
nor I_62141 (I1059981,I1059854,I1332736);
and I_62142 (I1059998,I1059981,I1332718);
or I_62143 (I1060015,I1059998,I1332721);
DFFARX1 I_62144 (I1060015,I3563,I1059591,I1060041,);
nor I_62145 (I1060049,I1060041,I1059775);
DFFARX1 I_62146 (I1060049,I3563,I1059591,I1059562,);
nand I_62147 (I1060080,I1060041,I1059682);
nand I_62148 (I1060097,I1059775,I1060080);
nor I_62149 (I1059571,I1060097,I1059741);
not I_62150 (I1060152,I3570);
DFFARX1 I_62151 (I1342848,I3563,I1060152,I1060178,);
DFFARX1 I_62152 (I1060178,I3563,I1060152,I1060195,);
not I_62153 (I1060144,I1060195);
not I_62154 (I1060217,I1060178);
DFFARX1 I_62155 (I1342842,I3563,I1060152,I1060243,);
nand I_62156 (I1060251,I1060243,I1342833);
not I_62157 (I1060268,I1342833);
not I_62158 (I1060285,I1342860);
nand I_62159 (I1060302,I1342845,I1342854);
and I_62160 (I1060319,I1342845,I1342854);
not I_62161 (I1060336,I1342839);
nand I_62162 (I1060353,I1060336,I1060285);
nor I_62163 (I1060126,I1060353,I1060251);
nor I_62164 (I1060384,I1060268,I1060353);
nand I_62165 (I1060129,I1060319,I1060384);
not I_62166 (I1060415,I1342857);
nor I_62167 (I1060432,I1060415,I1342845);
nor I_62168 (I1060449,I1060432,I1342839);
nor I_62169 (I1060466,I1060217,I1060449);
DFFARX1 I_62170 (I1060466,I3563,I1060152,I1060138,);
not I_62171 (I1060497,I1060432);
DFFARX1 I_62172 (I1060497,I3563,I1060152,I1060141,);
and I_62173 (I1060135,I1060243,I1060432);
nor I_62174 (I1060542,I1060415,I1342851);
and I_62175 (I1060559,I1060542,I1342833);
or I_62176 (I1060576,I1060559,I1342836);
DFFARX1 I_62177 (I1060576,I3563,I1060152,I1060602,);
nor I_62178 (I1060610,I1060602,I1060336);
DFFARX1 I_62179 (I1060610,I3563,I1060152,I1060123,);
nand I_62180 (I1060641,I1060602,I1060243);
nand I_62181 (I1060658,I1060336,I1060641);
nor I_62182 (I1060132,I1060658,I1060302);
not I_62183 (I1060713,I3570);
DFFARX1 I_62184 (I461050,I3563,I1060713,I1060739,);
DFFARX1 I_62185 (I1060739,I3563,I1060713,I1060756,);
not I_62186 (I1060705,I1060756);
not I_62187 (I1060778,I1060739);
DFFARX1 I_62188 (I461038,I3563,I1060713,I1060804,);
nand I_62189 (I1060812,I1060804,I461044);
not I_62190 (I1060829,I461044);
not I_62191 (I1060846,I461041);
nand I_62192 (I1060863,I461029,I461026);
and I_62193 (I1060880,I461029,I461026);
not I_62194 (I1060897,I461053);
nand I_62195 (I1060914,I1060897,I1060846);
nor I_62196 (I1060687,I1060914,I1060812);
nor I_62197 (I1060945,I1060829,I1060914);
nand I_62198 (I1060690,I1060880,I1060945);
not I_62199 (I1060976,I461026);
nor I_62200 (I1060993,I1060976,I461029);
nor I_62201 (I1061010,I1060993,I461053);
nor I_62202 (I1061027,I1060778,I1061010);
DFFARX1 I_62203 (I1061027,I3563,I1060713,I1060699,);
not I_62204 (I1061058,I1060993);
DFFARX1 I_62205 (I1061058,I3563,I1060713,I1060702,);
and I_62206 (I1060696,I1060804,I1060993);
nor I_62207 (I1061103,I1060976,I461035);
and I_62208 (I1061120,I1061103,I461032);
or I_62209 (I1061137,I1061120,I461047);
DFFARX1 I_62210 (I1061137,I3563,I1060713,I1061163,);
nor I_62211 (I1061171,I1061163,I1060897);
DFFARX1 I_62212 (I1061171,I3563,I1060713,I1060684,);
nand I_62213 (I1061202,I1061163,I1060804);
nand I_62214 (I1061219,I1060897,I1061202);
nor I_62215 (I1060693,I1061219,I1060863);
not I_62216 (I1061274,I3570);
DFFARX1 I_62217 (I444730,I3563,I1061274,I1061300,);
DFFARX1 I_62218 (I1061300,I3563,I1061274,I1061317,);
not I_62219 (I1061266,I1061317);
not I_62220 (I1061339,I1061300);
DFFARX1 I_62221 (I444718,I3563,I1061274,I1061365,);
nand I_62222 (I1061373,I1061365,I444724);
not I_62223 (I1061390,I444724);
not I_62224 (I1061407,I444721);
nand I_62225 (I1061424,I444709,I444706);
and I_62226 (I1061441,I444709,I444706);
not I_62227 (I1061458,I444733);
nand I_62228 (I1061475,I1061458,I1061407);
nor I_62229 (I1061248,I1061475,I1061373);
nor I_62230 (I1061506,I1061390,I1061475);
nand I_62231 (I1061251,I1061441,I1061506);
not I_62232 (I1061537,I444706);
nor I_62233 (I1061554,I1061537,I444709);
nor I_62234 (I1061571,I1061554,I444733);
nor I_62235 (I1061588,I1061339,I1061571);
DFFARX1 I_62236 (I1061588,I3563,I1061274,I1061260,);
not I_62237 (I1061619,I1061554);
DFFARX1 I_62238 (I1061619,I3563,I1061274,I1061263,);
and I_62239 (I1061257,I1061365,I1061554);
nor I_62240 (I1061664,I1061537,I444715);
and I_62241 (I1061681,I1061664,I444712);
or I_62242 (I1061698,I1061681,I444727);
DFFARX1 I_62243 (I1061698,I3563,I1061274,I1061724,);
nor I_62244 (I1061732,I1061724,I1061458);
DFFARX1 I_62245 (I1061732,I3563,I1061274,I1061245,);
nand I_62246 (I1061763,I1061724,I1061365);
nand I_62247 (I1061780,I1061458,I1061763);
nor I_62248 (I1061254,I1061780,I1061424);
not I_62249 (I1061835,I3570);
DFFARX1 I_62250 (I10124,I3563,I1061835,I1061861,);
DFFARX1 I_62251 (I1061861,I3563,I1061835,I1061878,);
not I_62252 (I1061827,I1061878);
not I_62253 (I1061900,I1061861);
DFFARX1 I_62254 (I10136,I3563,I1061835,I1061926,);
nand I_62255 (I1061934,I1061926,I10133);
not I_62256 (I1061951,I10133);
not I_62257 (I1061968,I10124);
nand I_62258 (I1061985,I10118,I10118);
and I_62259 (I1062002,I10118,I10118);
not I_62260 (I1062019,I10139);
nand I_62261 (I1062036,I1062019,I1061968);
nor I_62262 (I1061809,I1062036,I1061934);
nor I_62263 (I1062067,I1061951,I1062036);
nand I_62264 (I1061812,I1062002,I1062067);
not I_62265 (I1062098,I10130);
nor I_62266 (I1062115,I1062098,I10118);
nor I_62267 (I1062132,I1062115,I10139);
nor I_62268 (I1062149,I1061900,I1062132);
DFFARX1 I_62269 (I1062149,I3563,I1061835,I1061821,);
not I_62270 (I1062180,I1062115);
DFFARX1 I_62271 (I1062180,I3563,I1061835,I1061824,);
and I_62272 (I1061818,I1061926,I1062115);
nor I_62273 (I1062225,I1062098,I10121);
and I_62274 (I1062242,I1062225,I10121);
or I_62275 (I1062259,I1062242,I10127);
DFFARX1 I_62276 (I1062259,I3563,I1061835,I1062285,);
nor I_62277 (I1062293,I1062285,I1062019);
DFFARX1 I_62278 (I1062293,I3563,I1061835,I1061806,);
nand I_62279 (I1062324,I1062285,I1061926);
nand I_62280 (I1062341,I1062019,I1062324);
nor I_62281 (I1061815,I1062341,I1061985);
not I_62282 (I1062396,I3570);
DFFARX1 I_62283 (I590209,I3563,I1062396,I1062422,);
DFFARX1 I_62284 (I1062422,I3563,I1062396,I1062439,);
not I_62285 (I1062388,I1062439);
not I_62286 (I1062461,I1062422);
DFFARX1 I_62287 (I590224,I3563,I1062396,I1062487,);
nand I_62288 (I1062495,I1062487,I590215);
not I_62289 (I1062512,I590215);
not I_62290 (I1062529,I590221);
nand I_62291 (I1062546,I590218,I590227);
and I_62292 (I1062563,I590218,I590227);
not I_62293 (I1062580,I590212);
nand I_62294 (I1062597,I1062580,I1062529);
nor I_62295 (I1062370,I1062597,I1062495);
nor I_62296 (I1062628,I1062512,I1062597);
nand I_62297 (I1062373,I1062563,I1062628);
not I_62298 (I1062659,I590209);
nor I_62299 (I1062676,I1062659,I590218);
nor I_62300 (I1062693,I1062676,I590212);
nor I_62301 (I1062710,I1062461,I1062693);
DFFARX1 I_62302 (I1062710,I3563,I1062396,I1062382,);
not I_62303 (I1062741,I1062676);
DFFARX1 I_62304 (I1062741,I3563,I1062396,I1062385,);
and I_62305 (I1062379,I1062487,I1062676);
nor I_62306 (I1062786,I1062659,I590233);
and I_62307 (I1062803,I1062786,I590212);
or I_62308 (I1062820,I1062803,I590230);
DFFARX1 I_62309 (I1062820,I3563,I1062396,I1062846,);
nor I_62310 (I1062854,I1062846,I1062580);
DFFARX1 I_62311 (I1062854,I3563,I1062396,I1062367,);
nand I_62312 (I1062885,I1062846,I1062487);
nand I_62313 (I1062902,I1062580,I1062885);
nor I_62314 (I1062376,I1062902,I1062546);
not I_62315 (I1062957,I3570);
DFFARX1 I_62316 (I440378,I3563,I1062957,I1062983,);
DFFARX1 I_62317 (I1062983,I3563,I1062957,I1063000,);
not I_62318 (I1062949,I1063000);
not I_62319 (I1063022,I1062983);
DFFARX1 I_62320 (I440366,I3563,I1062957,I1063048,);
nand I_62321 (I1063056,I1063048,I440372);
not I_62322 (I1063073,I440372);
not I_62323 (I1063090,I440369);
nand I_62324 (I1063107,I440357,I440354);
and I_62325 (I1063124,I440357,I440354);
not I_62326 (I1063141,I440381);
nand I_62327 (I1063158,I1063141,I1063090);
nor I_62328 (I1062931,I1063158,I1063056);
nor I_62329 (I1063189,I1063073,I1063158);
nand I_62330 (I1062934,I1063124,I1063189);
not I_62331 (I1063220,I440354);
nor I_62332 (I1063237,I1063220,I440357);
nor I_62333 (I1063254,I1063237,I440381);
nor I_62334 (I1063271,I1063022,I1063254);
DFFARX1 I_62335 (I1063271,I3563,I1062957,I1062943,);
not I_62336 (I1063302,I1063237);
DFFARX1 I_62337 (I1063302,I3563,I1062957,I1062946,);
and I_62338 (I1062940,I1063048,I1063237);
nor I_62339 (I1063347,I1063220,I440363);
and I_62340 (I1063364,I1063347,I440360);
or I_62341 (I1063381,I1063364,I440375);
DFFARX1 I_62342 (I1063381,I3563,I1062957,I1063407,);
nor I_62343 (I1063415,I1063407,I1063141);
DFFARX1 I_62344 (I1063415,I3563,I1062957,I1062928,);
nand I_62345 (I1063446,I1063407,I1063048);
nand I_62346 (I1063463,I1063141,I1063446);
nor I_62347 (I1062937,I1063463,I1063107);
not I_62348 (I1063518,I3570);
DFFARX1 I_62349 (I169071,I3563,I1063518,I1063544,);
DFFARX1 I_62350 (I1063544,I3563,I1063518,I1063561,);
not I_62351 (I1063510,I1063561);
not I_62352 (I1063583,I1063544);
DFFARX1 I_62353 (I169086,I3563,I1063518,I1063609,);
nand I_62354 (I1063617,I1063609,I169068);
not I_62355 (I1063634,I169068);
not I_62356 (I1063651,I169077);
nand I_62357 (I1063668,I169083,I169074);
and I_62358 (I1063685,I169083,I169074);
not I_62359 (I1063702,I169071);
nand I_62360 (I1063719,I1063702,I1063651);
nor I_62361 (I1063492,I1063719,I1063617);
nor I_62362 (I1063750,I1063634,I1063719);
nand I_62363 (I1063495,I1063685,I1063750);
not I_62364 (I1063781,I169068);
nor I_62365 (I1063798,I1063781,I169083);
nor I_62366 (I1063815,I1063798,I169071);
nor I_62367 (I1063832,I1063583,I1063815);
DFFARX1 I_62368 (I1063832,I3563,I1063518,I1063504,);
not I_62369 (I1063863,I1063798);
DFFARX1 I_62370 (I1063863,I3563,I1063518,I1063507,);
and I_62371 (I1063501,I1063609,I1063798);
nor I_62372 (I1063908,I1063781,I169092);
and I_62373 (I1063925,I1063908,I169089);
or I_62374 (I1063942,I1063925,I169080);
DFFARX1 I_62375 (I1063942,I3563,I1063518,I1063968,);
nor I_62376 (I1063976,I1063968,I1063702);
DFFARX1 I_62377 (I1063976,I3563,I1063518,I1063489,);
nand I_62378 (I1064007,I1063968,I1063609);
nand I_62379 (I1064024,I1063702,I1064007);
nor I_62380 (I1063498,I1064024,I1063668);
not I_62381 (I1064079,I3570);
DFFARX1 I_62382 (I645697,I3563,I1064079,I1064105,);
DFFARX1 I_62383 (I1064105,I3563,I1064079,I1064122,);
not I_62384 (I1064071,I1064122);
not I_62385 (I1064144,I1064105);
DFFARX1 I_62386 (I645712,I3563,I1064079,I1064170,);
nand I_62387 (I1064178,I1064170,I645703);
not I_62388 (I1064195,I645703);
not I_62389 (I1064212,I645709);
nand I_62390 (I1064229,I645706,I645715);
and I_62391 (I1064246,I645706,I645715);
not I_62392 (I1064263,I645700);
nand I_62393 (I1064280,I1064263,I1064212);
nor I_62394 (I1064053,I1064280,I1064178);
nor I_62395 (I1064311,I1064195,I1064280);
nand I_62396 (I1064056,I1064246,I1064311);
not I_62397 (I1064342,I645697);
nor I_62398 (I1064359,I1064342,I645706);
nor I_62399 (I1064376,I1064359,I645700);
nor I_62400 (I1064393,I1064144,I1064376);
DFFARX1 I_62401 (I1064393,I3563,I1064079,I1064065,);
not I_62402 (I1064424,I1064359);
DFFARX1 I_62403 (I1064424,I3563,I1064079,I1064068,);
and I_62404 (I1064062,I1064170,I1064359);
nor I_62405 (I1064469,I1064342,I645721);
and I_62406 (I1064486,I1064469,I645700);
or I_62407 (I1064503,I1064486,I645718);
DFFARX1 I_62408 (I1064503,I3563,I1064079,I1064529,);
nor I_62409 (I1064537,I1064529,I1064263);
DFFARX1 I_62410 (I1064537,I3563,I1064079,I1064050,);
nand I_62411 (I1064568,I1064529,I1064170);
nand I_62412 (I1064585,I1064263,I1064568);
nor I_62413 (I1064059,I1064585,I1064229);
not I_62414 (I1064640,I3570);
DFFARX1 I_62415 (I133074,I3563,I1064640,I1064666,);
DFFARX1 I_62416 (I1064666,I3563,I1064640,I1064683,);
not I_62417 (I1064632,I1064683);
not I_62418 (I1064705,I1064666);
DFFARX1 I_62419 (I133062,I3563,I1064640,I1064731,);
nand I_62420 (I1064739,I1064731,I133077);
not I_62421 (I1064756,I133077);
not I_62422 (I1064773,I133065);
nand I_62423 (I1064790,I133086,I133080);
and I_62424 (I1064807,I133086,I133080);
not I_62425 (I1064824,I133068);
nand I_62426 (I1064841,I1064824,I1064773);
nor I_62427 (I1064614,I1064841,I1064739);
nor I_62428 (I1064872,I1064756,I1064841);
nand I_62429 (I1064617,I1064807,I1064872);
not I_62430 (I1064903,I133071);
nor I_62431 (I1064920,I1064903,I133086);
nor I_62432 (I1064937,I1064920,I133068);
nor I_62433 (I1064954,I1064705,I1064937);
DFFARX1 I_62434 (I1064954,I3563,I1064640,I1064626,);
not I_62435 (I1064985,I1064920);
DFFARX1 I_62436 (I1064985,I3563,I1064640,I1064629,);
and I_62437 (I1064623,I1064731,I1064920);
nor I_62438 (I1065030,I1064903,I133065);
and I_62439 (I1065047,I1065030,I133062);
or I_62440 (I1065064,I1065047,I133083);
DFFARX1 I_62441 (I1065064,I3563,I1064640,I1065090,);
nor I_62442 (I1065098,I1065090,I1064824);
DFFARX1 I_62443 (I1065098,I3563,I1064640,I1064611,);
nand I_62444 (I1065129,I1065090,I1064731);
nand I_62445 (I1065146,I1064824,I1065129);
nor I_62446 (I1064620,I1065146,I1064790);
not I_62447 (I1065201,I3570);
DFFARX1 I_62448 (I352842,I3563,I1065201,I1065227,);
DFFARX1 I_62449 (I1065227,I3563,I1065201,I1065244,);
not I_62450 (I1065193,I1065244);
not I_62451 (I1065266,I1065227);
DFFARX1 I_62452 (I352839,I3563,I1065201,I1065292,);
nand I_62453 (I1065300,I1065292,I352833);
not I_62454 (I1065317,I352833);
not I_62455 (I1065334,I352830);
nand I_62456 (I1065351,I352824,I352821);
and I_62457 (I1065368,I352824,I352821);
not I_62458 (I1065385,I352836);
nand I_62459 (I1065402,I1065385,I1065334);
nor I_62460 (I1065175,I1065402,I1065300);
nor I_62461 (I1065433,I1065317,I1065402);
nand I_62462 (I1065178,I1065368,I1065433);
not I_62463 (I1065464,I352848);
nor I_62464 (I1065481,I1065464,I352824);
nor I_62465 (I1065498,I1065481,I352836);
nor I_62466 (I1065515,I1065266,I1065498);
DFFARX1 I_62467 (I1065515,I3563,I1065201,I1065187,);
not I_62468 (I1065546,I1065481);
DFFARX1 I_62469 (I1065546,I3563,I1065201,I1065190,);
and I_62470 (I1065184,I1065292,I1065481);
nor I_62471 (I1065591,I1065464,I352845);
and I_62472 (I1065608,I1065591,I352821);
or I_62473 (I1065625,I1065608,I352827);
DFFARX1 I_62474 (I1065625,I3563,I1065201,I1065651,);
nor I_62475 (I1065659,I1065651,I1065385);
DFFARX1 I_62476 (I1065659,I3563,I1065201,I1065172,);
nand I_62477 (I1065690,I1065651,I1065292);
nand I_62478 (I1065707,I1065385,I1065690);
nor I_62479 (I1065181,I1065707,I1065351);
not I_62480 (I1065762,I3570);
DFFARX1 I_62481 (I569164,I3563,I1065762,I1065788,);
DFFARX1 I_62482 (I1065788,I3563,I1065762,I1065805,);
not I_62483 (I1065754,I1065805);
not I_62484 (I1065827,I1065788);
DFFARX1 I_62485 (I569161,I3563,I1065762,I1065853,);
nand I_62486 (I1065861,I1065853,I569155);
not I_62487 (I1065878,I569155);
not I_62488 (I1065895,I569167);
nand I_62489 (I1065912,I569170,I569149);
and I_62490 (I1065929,I569170,I569149);
not I_62491 (I1065946,I569146);
nand I_62492 (I1065963,I1065946,I1065895);
nor I_62493 (I1065736,I1065963,I1065861);
nor I_62494 (I1065994,I1065878,I1065963);
nand I_62495 (I1065739,I1065929,I1065994);
not I_62496 (I1066025,I569152);
nor I_62497 (I1066042,I1066025,I569170);
nor I_62498 (I1066059,I1066042,I569146);
nor I_62499 (I1066076,I1065827,I1066059);
DFFARX1 I_62500 (I1066076,I3563,I1065762,I1065748,);
not I_62501 (I1066107,I1066042);
DFFARX1 I_62502 (I1066107,I3563,I1065762,I1065751,);
and I_62503 (I1065745,I1065853,I1066042);
nor I_62504 (I1066152,I1066025,I569146);
and I_62505 (I1066169,I1066152,I569158);
or I_62506 (I1066186,I1066169,I569149);
DFFARX1 I_62507 (I1066186,I3563,I1065762,I1066212,);
nor I_62508 (I1066220,I1066212,I1065946);
DFFARX1 I_62509 (I1066220,I3563,I1065762,I1065733,);
nand I_62510 (I1066251,I1066212,I1065853);
nand I_62511 (I1066268,I1065946,I1066251);
nor I_62512 (I1065742,I1066268,I1065912);
not I_62513 (I1066323,I3570);
DFFARX1 I_62514 (I674022,I3563,I1066323,I1066349,);
DFFARX1 I_62515 (I1066349,I3563,I1066323,I1066366,);
not I_62516 (I1066315,I1066366);
not I_62517 (I1066388,I1066349);
DFFARX1 I_62518 (I674034,I3563,I1066323,I1066414,);
nand I_62519 (I1066422,I1066414,I674043);
not I_62520 (I1066439,I674043);
not I_62521 (I1066456,I674025);
nand I_62522 (I1066473,I674028,I674019);
and I_62523 (I1066490,I674028,I674019);
not I_62524 (I1066507,I674037);
nand I_62525 (I1066524,I1066507,I1066456);
nor I_62526 (I1066297,I1066524,I1066422);
nor I_62527 (I1066555,I1066439,I1066524);
nand I_62528 (I1066300,I1066490,I1066555);
not I_62529 (I1066586,I674040);
nor I_62530 (I1066603,I1066586,I674028);
nor I_62531 (I1066620,I1066603,I674037);
nor I_62532 (I1066637,I1066388,I1066620);
DFFARX1 I_62533 (I1066637,I3563,I1066323,I1066309,);
not I_62534 (I1066668,I1066603);
DFFARX1 I_62535 (I1066668,I3563,I1066323,I1066312,);
and I_62536 (I1066306,I1066414,I1066603);
nor I_62537 (I1066713,I1066586,I674019);
and I_62538 (I1066730,I1066713,I674031);
or I_62539 (I1066747,I1066730,I674022);
DFFARX1 I_62540 (I1066747,I3563,I1066323,I1066773,);
nor I_62541 (I1066781,I1066773,I1066507);
DFFARX1 I_62542 (I1066781,I3563,I1066323,I1066294,);
nand I_62543 (I1066812,I1066773,I1066414);
nand I_62544 (I1066829,I1066507,I1066812);
nor I_62545 (I1066303,I1066829,I1066473);
not I_62546 (I1066884,I3570);
DFFARX1 I_62547 (I84590,I3563,I1066884,I1066910,);
DFFARX1 I_62548 (I1066910,I3563,I1066884,I1066927,);
not I_62549 (I1066876,I1066927);
not I_62550 (I1066949,I1066910);
DFFARX1 I_62551 (I84578,I3563,I1066884,I1066975,);
nand I_62552 (I1066983,I1066975,I84593);
not I_62553 (I1067000,I84593);
not I_62554 (I1067017,I84581);
nand I_62555 (I1067034,I84602,I84596);
and I_62556 (I1067051,I84602,I84596);
not I_62557 (I1067068,I84584);
nand I_62558 (I1067085,I1067068,I1067017);
nor I_62559 (I1066858,I1067085,I1066983);
nor I_62560 (I1067116,I1067000,I1067085);
nand I_62561 (I1066861,I1067051,I1067116);
not I_62562 (I1067147,I84587);
nor I_62563 (I1067164,I1067147,I84602);
nor I_62564 (I1067181,I1067164,I84584);
nor I_62565 (I1067198,I1066949,I1067181);
DFFARX1 I_62566 (I1067198,I3563,I1066884,I1066870,);
not I_62567 (I1067229,I1067164);
DFFARX1 I_62568 (I1067229,I3563,I1066884,I1066873,);
and I_62569 (I1066867,I1066975,I1067164);
nor I_62570 (I1067274,I1067147,I84581);
and I_62571 (I1067291,I1067274,I84578);
or I_62572 (I1067308,I1067291,I84599);
DFFARX1 I_62573 (I1067308,I3563,I1066884,I1067334,);
nor I_62574 (I1067342,I1067334,I1067068);
DFFARX1 I_62575 (I1067342,I3563,I1066884,I1066855,);
nand I_62576 (I1067373,I1067334,I1066975);
nand I_62577 (I1067390,I1067068,I1067373);
nor I_62578 (I1066864,I1067390,I1067034);
not I_62579 (I1067445,I3570);
DFFARX1 I_62580 (I818443,I3563,I1067445,I1067471,);
DFFARX1 I_62581 (I1067471,I3563,I1067445,I1067488,);
not I_62582 (I1067437,I1067488);
not I_62583 (I1067510,I1067471);
DFFARX1 I_62584 (I818440,I3563,I1067445,I1067536,);
nand I_62585 (I1067544,I1067536,I818455);
not I_62586 (I1067561,I818455);
not I_62587 (I1067578,I818452);
nand I_62588 (I1067595,I818449,I818437);
and I_62589 (I1067612,I818449,I818437);
not I_62590 (I1067629,I818434);
nand I_62591 (I1067646,I1067629,I1067578);
nor I_62592 (I1067419,I1067646,I1067544);
nor I_62593 (I1067677,I1067561,I1067646);
nand I_62594 (I1067422,I1067612,I1067677);
not I_62595 (I1067708,I818440);
nor I_62596 (I1067725,I1067708,I818449);
nor I_62597 (I1067742,I1067725,I818434);
nor I_62598 (I1067759,I1067510,I1067742);
DFFARX1 I_62599 (I1067759,I3563,I1067445,I1067431,);
not I_62600 (I1067790,I1067725);
DFFARX1 I_62601 (I1067790,I3563,I1067445,I1067434,);
and I_62602 (I1067428,I1067536,I1067725);
nor I_62603 (I1067835,I1067708,I818446);
and I_62604 (I1067852,I1067835,I818434);
or I_62605 (I1067869,I1067852,I818437);
DFFARX1 I_62606 (I1067869,I3563,I1067445,I1067895,);
nor I_62607 (I1067903,I1067895,I1067629);
DFFARX1 I_62608 (I1067903,I3563,I1067445,I1067416,);
nand I_62609 (I1067934,I1067895,I1067536);
nand I_62610 (I1067951,I1067629,I1067934);
nor I_62611 (I1067425,I1067951,I1067595);
not I_62612 (I1068006,I3570);
DFFARX1 I_62613 (I134655,I3563,I1068006,I1068032,);
DFFARX1 I_62614 (I1068032,I3563,I1068006,I1068049,);
not I_62615 (I1067998,I1068049);
not I_62616 (I1068071,I1068032);
DFFARX1 I_62617 (I134643,I3563,I1068006,I1068097,);
nand I_62618 (I1068105,I1068097,I134658);
not I_62619 (I1068122,I134658);
not I_62620 (I1068139,I134646);
nand I_62621 (I1068156,I134667,I134661);
and I_62622 (I1068173,I134667,I134661);
not I_62623 (I1068190,I134649);
nand I_62624 (I1068207,I1068190,I1068139);
nor I_62625 (I1067980,I1068207,I1068105);
nor I_62626 (I1068238,I1068122,I1068207);
nand I_62627 (I1067983,I1068173,I1068238);
not I_62628 (I1068269,I134652);
nor I_62629 (I1068286,I1068269,I134667);
nor I_62630 (I1068303,I1068286,I134649);
nor I_62631 (I1068320,I1068071,I1068303);
DFFARX1 I_62632 (I1068320,I3563,I1068006,I1067992,);
not I_62633 (I1068351,I1068286);
DFFARX1 I_62634 (I1068351,I3563,I1068006,I1067995,);
and I_62635 (I1067989,I1068097,I1068286);
nor I_62636 (I1068396,I1068269,I134646);
and I_62637 (I1068413,I1068396,I134643);
or I_62638 (I1068430,I1068413,I134664);
DFFARX1 I_62639 (I1068430,I3563,I1068006,I1068456,);
nor I_62640 (I1068464,I1068456,I1068190);
DFFARX1 I_62641 (I1068464,I3563,I1068006,I1067977,);
nand I_62642 (I1068495,I1068456,I1068097);
nand I_62643 (I1068512,I1068190,I1068495);
nor I_62644 (I1067986,I1068512,I1068156);
not I_62645 (I1068567,I3570);
DFFARX1 I_62646 (I148884,I3563,I1068567,I1068593,);
DFFARX1 I_62647 (I1068593,I3563,I1068567,I1068610,);
not I_62648 (I1068559,I1068610);
not I_62649 (I1068632,I1068593);
DFFARX1 I_62650 (I148872,I3563,I1068567,I1068658,);
nand I_62651 (I1068666,I1068658,I148887);
not I_62652 (I1068683,I148887);
not I_62653 (I1068700,I148875);
nand I_62654 (I1068717,I148896,I148890);
and I_62655 (I1068734,I148896,I148890);
not I_62656 (I1068751,I148878);
nand I_62657 (I1068768,I1068751,I1068700);
nor I_62658 (I1068541,I1068768,I1068666);
nor I_62659 (I1068799,I1068683,I1068768);
nand I_62660 (I1068544,I1068734,I1068799);
not I_62661 (I1068830,I148881);
nor I_62662 (I1068847,I1068830,I148896);
nor I_62663 (I1068864,I1068847,I148878);
nor I_62664 (I1068881,I1068632,I1068864);
DFFARX1 I_62665 (I1068881,I3563,I1068567,I1068553,);
not I_62666 (I1068912,I1068847);
DFFARX1 I_62667 (I1068912,I3563,I1068567,I1068556,);
and I_62668 (I1068550,I1068658,I1068847);
nor I_62669 (I1068957,I1068830,I148875);
and I_62670 (I1068974,I1068957,I148872);
or I_62671 (I1068991,I1068974,I148893);
DFFARX1 I_62672 (I1068991,I3563,I1068567,I1069017,);
nor I_62673 (I1069025,I1069017,I1068751);
DFFARX1 I_62674 (I1069025,I3563,I1068567,I1068538,);
nand I_62675 (I1069056,I1069017,I1068658);
nand I_62676 (I1069073,I1068751,I1069056);
nor I_62677 (I1068547,I1069073,I1068717);
not I_62678 (I1069128,I3570);
DFFARX1 I_62679 (I998855,I3563,I1069128,I1069154,);
DFFARX1 I_62680 (I1069154,I3563,I1069128,I1069171,);
not I_62681 (I1069120,I1069171);
not I_62682 (I1069193,I1069154);
DFFARX1 I_62683 (I998882,I3563,I1069128,I1069219,);
nand I_62684 (I1069227,I1069219,I998873);
not I_62685 (I1069244,I998873);
not I_62686 (I1069261,I998855);
nand I_62687 (I1069278,I998867,I998870);
and I_62688 (I1069295,I998867,I998870);
not I_62689 (I1069312,I998879);
nand I_62690 (I1069329,I1069312,I1069261);
nor I_62691 (I1069102,I1069329,I1069227);
nor I_62692 (I1069360,I1069244,I1069329);
nand I_62693 (I1069105,I1069295,I1069360);
not I_62694 (I1069391,I998864);
nor I_62695 (I1069408,I1069391,I998867);
nor I_62696 (I1069425,I1069408,I998879);
nor I_62697 (I1069442,I1069193,I1069425);
DFFARX1 I_62698 (I1069442,I3563,I1069128,I1069114,);
not I_62699 (I1069473,I1069408);
DFFARX1 I_62700 (I1069473,I3563,I1069128,I1069117,);
and I_62701 (I1069111,I1069219,I1069408);
nor I_62702 (I1069518,I1069391,I998858);
and I_62703 (I1069535,I1069518,I998861);
or I_62704 (I1069552,I1069535,I998876);
DFFARX1 I_62705 (I1069552,I3563,I1069128,I1069578,);
nor I_62706 (I1069586,I1069578,I1069312);
DFFARX1 I_62707 (I1069586,I3563,I1069128,I1069099,);
nand I_62708 (I1069617,I1069578,I1069219);
nand I_62709 (I1069634,I1069312,I1069617);
nor I_62710 (I1069108,I1069634,I1069278);
not I_62711 (I1069689,I3570);
DFFARX1 I_62712 (I1221638,I3563,I1069689,I1069715,);
DFFARX1 I_62713 (I1069715,I3563,I1069689,I1069732,);
not I_62714 (I1069681,I1069732);
not I_62715 (I1069754,I1069715);
DFFARX1 I_62716 (I1221629,I3563,I1069689,I1069780,);
nand I_62717 (I1069788,I1069780,I1221626);
not I_62718 (I1069805,I1221626);
not I_62719 (I1069822,I1221635);
nand I_62720 (I1069839,I1221644,I1221626);
and I_62721 (I1069856,I1221644,I1221626);
not I_62722 (I1069873,I1221623);
nand I_62723 (I1069890,I1069873,I1069822);
nor I_62724 (I1069663,I1069890,I1069788);
nor I_62725 (I1069921,I1069805,I1069890);
nand I_62726 (I1069666,I1069856,I1069921);
not I_62727 (I1069952,I1221632);
nor I_62728 (I1069969,I1069952,I1221644);
nor I_62729 (I1069986,I1069969,I1221623);
nor I_62730 (I1070003,I1069754,I1069986);
DFFARX1 I_62731 (I1070003,I3563,I1069689,I1069675,);
not I_62732 (I1070034,I1069969);
DFFARX1 I_62733 (I1070034,I3563,I1069689,I1069678,);
and I_62734 (I1069672,I1069780,I1069969);
nor I_62735 (I1070079,I1069952,I1221647);
and I_62736 (I1070096,I1070079,I1221623);
or I_62737 (I1070113,I1070096,I1221641);
DFFARX1 I_62738 (I1070113,I3563,I1069689,I1070139,);
nor I_62739 (I1070147,I1070139,I1069873);
DFFARX1 I_62740 (I1070147,I3563,I1069689,I1069660,);
nand I_62741 (I1070178,I1070139,I1069780);
nand I_62742 (I1070195,I1069873,I1070178);
nor I_62743 (I1069669,I1070195,I1069839);
not I_62744 (I1070250,I3570);
DFFARX1 I_62745 (I719684,I3563,I1070250,I1070276,);
DFFARX1 I_62746 (I1070276,I3563,I1070250,I1070293,);
not I_62747 (I1070242,I1070293);
not I_62748 (I1070315,I1070276);
DFFARX1 I_62749 (I719696,I3563,I1070250,I1070341,);
nand I_62750 (I1070349,I1070341,I719705);
not I_62751 (I1070366,I719705);
not I_62752 (I1070383,I719687);
nand I_62753 (I1070400,I719690,I719681);
and I_62754 (I1070417,I719690,I719681);
not I_62755 (I1070434,I719699);
nand I_62756 (I1070451,I1070434,I1070383);
nor I_62757 (I1070224,I1070451,I1070349);
nor I_62758 (I1070482,I1070366,I1070451);
nand I_62759 (I1070227,I1070417,I1070482);
not I_62760 (I1070513,I719702);
nor I_62761 (I1070530,I1070513,I719690);
nor I_62762 (I1070547,I1070530,I719699);
nor I_62763 (I1070564,I1070315,I1070547);
DFFARX1 I_62764 (I1070564,I3563,I1070250,I1070236,);
not I_62765 (I1070595,I1070530);
DFFARX1 I_62766 (I1070595,I3563,I1070250,I1070239,);
and I_62767 (I1070233,I1070341,I1070530);
nor I_62768 (I1070640,I1070513,I719681);
and I_62769 (I1070657,I1070640,I719693);
or I_62770 (I1070674,I1070657,I719684);
DFFARX1 I_62771 (I1070674,I3563,I1070250,I1070700,);
nor I_62772 (I1070708,I1070700,I1070434);
DFFARX1 I_62773 (I1070708,I3563,I1070250,I1070221,);
nand I_62774 (I1070739,I1070700,I1070341);
nand I_62775 (I1070756,I1070434,I1070739);
nor I_62776 (I1070230,I1070756,I1070400);
not I_62777 (I1070811,I3570);
DFFARX1 I_62778 (I771704,I3563,I1070811,I1070837,);
DFFARX1 I_62779 (I1070837,I3563,I1070811,I1070854,);
not I_62780 (I1070803,I1070854);
not I_62781 (I1070876,I1070837);
DFFARX1 I_62782 (I771716,I3563,I1070811,I1070902,);
nand I_62783 (I1070910,I1070902,I771725);
not I_62784 (I1070927,I771725);
not I_62785 (I1070944,I771707);
nand I_62786 (I1070961,I771710,I771701);
and I_62787 (I1070978,I771710,I771701);
not I_62788 (I1070995,I771719);
nand I_62789 (I1071012,I1070995,I1070944);
nor I_62790 (I1070785,I1071012,I1070910);
nor I_62791 (I1071043,I1070927,I1071012);
nand I_62792 (I1070788,I1070978,I1071043);
not I_62793 (I1071074,I771722);
nor I_62794 (I1071091,I1071074,I771710);
nor I_62795 (I1071108,I1071091,I771719);
nor I_62796 (I1071125,I1070876,I1071108);
DFFARX1 I_62797 (I1071125,I3563,I1070811,I1070797,);
not I_62798 (I1071156,I1071091);
DFFARX1 I_62799 (I1071156,I3563,I1070811,I1070800,);
and I_62800 (I1070794,I1070902,I1071091);
nor I_62801 (I1071201,I1071074,I771701);
and I_62802 (I1071218,I1071201,I771713);
or I_62803 (I1071235,I1071218,I771704);
DFFARX1 I_62804 (I1071235,I3563,I1070811,I1071261,);
nor I_62805 (I1071269,I1071261,I1070995);
DFFARX1 I_62806 (I1071269,I3563,I1070811,I1070782,);
nand I_62807 (I1071300,I1071261,I1070902);
nand I_62808 (I1071317,I1070995,I1071300);
nor I_62809 (I1070791,I1071317,I1070961);
not I_62810 (I1071372,I3570);
DFFARX1 I_62811 (I1237244,I3563,I1071372,I1071398,);
DFFARX1 I_62812 (I1071398,I3563,I1071372,I1071415,);
not I_62813 (I1071364,I1071415);
not I_62814 (I1071437,I1071398);
DFFARX1 I_62815 (I1237235,I3563,I1071372,I1071463,);
nand I_62816 (I1071471,I1071463,I1237232);
not I_62817 (I1071488,I1237232);
not I_62818 (I1071505,I1237241);
nand I_62819 (I1071522,I1237250,I1237232);
and I_62820 (I1071539,I1237250,I1237232);
not I_62821 (I1071556,I1237229);
nand I_62822 (I1071573,I1071556,I1071505);
nor I_62823 (I1071346,I1071573,I1071471);
nor I_62824 (I1071604,I1071488,I1071573);
nand I_62825 (I1071349,I1071539,I1071604);
not I_62826 (I1071635,I1237238);
nor I_62827 (I1071652,I1071635,I1237250);
nor I_62828 (I1071669,I1071652,I1237229);
nor I_62829 (I1071686,I1071437,I1071669);
DFFARX1 I_62830 (I1071686,I3563,I1071372,I1071358,);
not I_62831 (I1071717,I1071652);
DFFARX1 I_62832 (I1071717,I3563,I1071372,I1071361,);
and I_62833 (I1071355,I1071463,I1071652);
nor I_62834 (I1071762,I1071635,I1237253);
and I_62835 (I1071779,I1071762,I1237229);
or I_62836 (I1071796,I1071779,I1237247);
DFFARX1 I_62837 (I1071796,I3563,I1071372,I1071822,);
nor I_62838 (I1071830,I1071822,I1071556);
DFFARX1 I_62839 (I1071830,I3563,I1071372,I1071343,);
nand I_62840 (I1071861,I1071822,I1071463);
nand I_62841 (I1071878,I1071556,I1071861);
nor I_62842 (I1071352,I1071878,I1071522);
not I_62843 (I1071933,I3570);
DFFARX1 I_62844 (I214886,I3563,I1071933,I1071959,);
DFFARX1 I_62845 (I1071959,I3563,I1071933,I1071976,);
not I_62846 (I1071925,I1071976);
not I_62847 (I1071998,I1071959);
DFFARX1 I_62848 (I214901,I3563,I1071933,I1072024,);
nand I_62849 (I1072032,I1072024,I214883);
not I_62850 (I1072049,I214883);
not I_62851 (I1072066,I214892);
nand I_62852 (I1072083,I214898,I214889);
and I_62853 (I1072100,I214898,I214889);
not I_62854 (I1072117,I214886);
nand I_62855 (I1072134,I1072117,I1072066);
nor I_62856 (I1071907,I1072134,I1072032);
nor I_62857 (I1072165,I1072049,I1072134);
nand I_62858 (I1071910,I1072100,I1072165);
not I_62859 (I1072196,I214883);
nor I_62860 (I1072213,I1072196,I214898);
nor I_62861 (I1072230,I1072213,I214886);
nor I_62862 (I1072247,I1071998,I1072230);
DFFARX1 I_62863 (I1072247,I3563,I1071933,I1071919,);
not I_62864 (I1072278,I1072213);
DFFARX1 I_62865 (I1072278,I3563,I1071933,I1071922,);
and I_62866 (I1071916,I1072024,I1072213);
nor I_62867 (I1072323,I1072196,I214907);
and I_62868 (I1072340,I1072323,I214904);
or I_62869 (I1072357,I1072340,I214895);
DFFARX1 I_62870 (I1072357,I3563,I1071933,I1072383,);
nor I_62871 (I1072391,I1072383,I1072117);
DFFARX1 I_62872 (I1072391,I3563,I1071933,I1071904,);
nand I_62873 (I1072422,I1072383,I1072024);
nand I_62874 (I1072439,I1072117,I1072422);
nor I_62875 (I1071913,I1072439,I1072083);
not I_62876 (I1072494,I3570);
DFFARX1 I_62877 (I798292,I3563,I1072494,I1072520,);
DFFARX1 I_62878 (I1072520,I3563,I1072494,I1072537,);
not I_62879 (I1072486,I1072537);
not I_62880 (I1072559,I1072520);
DFFARX1 I_62881 (I798304,I3563,I1072494,I1072585,);
nand I_62882 (I1072593,I1072585,I798313);
not I_62883 (I1072610,I798313);
not I_62884 (I1072627,I798295);
nand I_62885 (I1072644,I798298,I798289);
and I_62886 (I1072661,I798298,I798289);
not I_62887 (I1072678,I798307);
nand I_62888 (I1072695,I1072678,I1072627);
nor I_62889 (I1072468,I1072695,I1072593);
nor I_62890 (I1072726,I1072610,I1072695);
nand I_62891 (I1072471,I1072661,I1072726);
not I_62892 (I1072757,I798310);
nor I_62893 (I1072774,I1072757,I798298);
nor I_62894 (I1072791,I1072774,I798307);
nor I_62895 (I1072808,I1072559,I1072791);
DFFARX1 I_62896 (I1072808,I3563,I1072494,I1072480,);
not I_62897 (I1072839,I1072774);
DFFARX1 I_62898 (I1072839,I3563,I1072494,I1072483,);
and I_62899 (I1072477,I1072585,I1072774);
nor I_62900 (I1072884,I1072757,I798289);
and I_62901 (I1072901,I1072884,I798301);
or I_62902 (I1072918,I1072901,I798292);
DFFARX1 I_62903 (I1072918,I3563,I1072494,I1072944,);
nor I_62904 (I1072952,I1072944,I1072678);
DFFARX1 I_62905 (I1072952,I3563,I1072494,I1072465,);
nand I_62906 (I1072983,I1072944,I1072585);
nand I_62907 (I1073000,I1072678,I1072983);
nor I_62908 (I1072474,I1073000,I1072644);
not I_62909 (I1073055,I3570);
DFFARX1 I_62910 (I841631,I3563,I1073055,I1073081,);
DFFARX1 I_62911 (I1073081,I3563,I1073055,I1073098,);
not I_62912 (I1073047,I1073098);
not I_62913 (I1073120,I1073081);
DFFARX1 I_62914 (I841628,I3563,I1073055,I1073146,);
nand I_62915 (I1073154,I1073146,I841643);
not I_62916 (I1073171,I841643);
not I_62917 (I1073188,I841640);
nand I_62918 (I1073205,I841637,I841625);
and I_62919 (I1073222,I841637,I841625);
not I_62920 (I1073239,I841622);
nand I_62921 (I1073256,I1073239,I1073188);
nor I_62922 (I1073029,I1073256,I1073154);
nor I_62923 (I1073287,I1073171,I1073256);
nand I_62924 (I1073032,I1073222,I1073287);
not I_62925 (I1073318,I841628);
nor I_62926 (I1073335,I1073318,I841637);
nor I_62927 (I1073352,I1073335,I841622);
nor I_62928 (I1073369,I1073120,I1073352);
DFFARX1 I_62929 (I1073369,I3563,I1073055,I1073041,);
not I_62930 (I1073400,I1073335);
DFFARX1 I_62931 (I1073400,I3563,I1073055,I1073044,);
and I_62932 (I1073038,I1073146,I1073335);
nor I_62933 (I1073445,I1073318,I841634);
and I_62934 (I1073462,I1073445,I841622);
or I_62935 (I1073479,I1073462,I841625);
DFFARX1 I_62936 (I1073479,I3563,I1073055,I1073505,);
nor I_62937 (I1073513,I1073505,I1073239);
DFFARX1 I_62938 (I1073513,I3563,I1073055,I1073026,);
nand I_62939 (I1073544,I1073505,I1073146);
nand I_62940 (I1073561,I1073239,I1073544);
nor I_62941 (I1073035,I1073561,I1073205);
not I_62942 (I1073616,I3570);
DFFARX1 I_62943 (I1044721,I3563,I1073616,I1073642,);
DFFARX1 I_62944 (I1073642,I3563,I1073616,I1073659,);
not I_62945 (I1073608,I1073659);
not I_62946 (I1073681,I1073642);
DFFARX1 I_62947 (I1044748,I3563,I1073616,I1073707,);
nand I_62948 (I1073715,I1073707,I1044739);
not I_62949 (I1073732,I1044739);
not I_62950 (I1073749,I1044721);
nand I_62951 (I1073766,I1044733,I1044736);
and I_62952 (I1073783,I1044733,I1044736);
not I_62953 (I1073800,I1044745);
nand I_62954 (I1073817,I1073800,I1073749);
nor I_62955 (I1073590,I1073817,I1073715);
nor I_62956 (I1073848,I1073732,I1073817);
nand I_62957 (I1073593,I1073783,I1073848);
not I_62958 (I1073879,I1044730);
nor I_62959 (I1073896,I1073879,I1044733);
nor I_62960 (I1073913,I1073896,I1044745);
nor I_62961 (I1073930,I1073681,I1073913);
DFFARX1 I_62962 (I1073930,I3563,I1073616,I1073602,);
not I_62963 (I1073961,I1073896);
DFFARX1 I_62964 (I1073961,I3563,I1073616,I1073605,);
and I_62965 (I1073599,I1073707,I1073896);
nor I_62966 (I1074006,I1073879,I1044724);
and I_62967 (I1074023,I1074006,I1044727);
or I_62968 (I1074040,I1074023,I1044742);
DFFARX1 I_62969 (I1074040,I3563,I1073616,I1074066,);
nor I_62970 (I1074074,I1074066,I1073800);
DFFARX1 I_62971 (I1074074,I3563,I1073616,I1073587,);
nand I_62972 (I1074105,I1074066,I1073707);
nand I_62973 (I1074122,I1073800,I1074105);
nor I_62974 (I1073596,I1074122,I1073766);
not I_62975 (I1074177,I3570);
DFFARX1 I_62976 (I1360698,I3563,I1074177,I1074203,);
DFFARX1 I_62977 (I1074203,I3563,I1074177,I1074220,);
not I_62978 (I1074169,I1074220);
not I_62979 (I1074242,I1074203);
DFFARX1 I_62980 (I1360692,I3563,I1074177,I1074268,);
nand I_62981 (I1074276,I1074268,I1360683);
not I_62982 (I1074293,I1360683);
not I_62983 (I1074310,I1360710);
nand I_62984 (I1074327,I1360695,I1360704);
and I_62985 (I1074344,I1360695,I1360704);
not I_62986 (I1074361,I1360689);
nand I_62987 (I1074378,I1074361,I1074310);
nor I_62988 (I1074151,I1074378,I1074276);
nor I_62989 (I1074409,I1074293,I1074378);
nand I_62990 (I1074154,I1074344,I1074409);
not I_62991 (I1074440,I1360707);
nor I_62992 (I1074457,I1074440,I1360695);
nor I_62993 (I1074474,I1074457,I1360689);
nor I_62994 (I1074491,I1074242,I1074474);
DFFARX1 I_62995 (I1074491,I3563,I1074177,I1074163,);
not I_62996 (I1074522,I1074457);
DFFARX1 I_62997 (I1074522,I3563,I1074177,I1074166,);
and I_62998 (I1074160,I1074268,I1074457);
nor I_62999 (I1074567,I1074440,I1360701);
and I_63000 (I1074584,I1074567,I1360683);
or I_63001 (I1074601,I1074584,I1360686);
DFFARX1 I_63002 (I1074601,I3563,I1074177,I1074627,);
nor I_63003 (I1074635,I1074627,I1074361);
DFFARX1 I_63004 (I1074635,I3563,I1074177,I1074148,);
nand I_63005 (I1074666,I1074627,I1074268);
nand I_63006 (I1074683,I1074361,I1074666);
nor I_63007 (I1074157,I1074683,I1074327);
not I_63008 (I1074738,I3570);
DFFARX1 I_63009 (I566784,I3563,I1074738,I1074764,);
DFFARX1 I_63010 (I1074764,I3563,I1074738,I1074781,);
not I_63011 (I1074730,I1074781);
not I_63012 (I1074803,I1074764);
DFFARX1 I_63013 (I566781,I3563,I1074738,I1074829,);
nand I_63014 (I1074837,I1074829,I566775);
not I_63015 (I1074854,I566775);
not I_63016 (I1074871,I566787);
nand I_63017 (I1074888,I566790,I566769);
and I_63018 (I1074905,I566790,I566769);
not I_63019 (I1074922,I566766);
nand I_63020 (I1074939,I1074922,I1074871);
nor I_63021 (I1074712,I1074939,I1074837);
nor I_63022 (I1074970,I1074854,I1074939);
nand I_63023 (I1074715,I1074905,I1074970);
not I_63024 (I1075001,I566772);
nor I_63025 (I1075018,I1075001,I566790);
nor I_63026 (I1075035,I1075018,I566766);
nor I_63027 (I1075052,I1074803,I1075035);
DFFARX1 I_63028 (I1075052,I3563,I1074738,I1074724,);
not I_63029 (I1075083,I1075018);
DFFARX1 I_63030 (I1075083,I3563,I1074738,I1074727,);
and I_63031 (I1074721,I1074829,I1075018);
nor I_63032 (I1075128,I1075001,I566766);
and I_63033 (I1075145,I1075128,I566778);
or I_63034 (I1075162,I1075145,I566769);
DFFARX1 I_63035 (I1075162,I3563,I1074738,I1075188,);
nor I_63036 (I1075196,I1075188,I1074922);
DFFARX1 I_63037 (I1075196,I3563,I1074738,I1074709,);
nand I_63038 (I1075227,I1075188,I1074829);
nand I_63039 (I1075244,I1074922,I1075227);
nor I_63040 (I1074718,I1075244,I1074888);
not I_63041 (I1075299,I3570);
DFFARX1 I_63042 (I519258,I3563,I1075299,I1075325,);
DFFARX1 I_63043 (I1075325,I3563,I1075299,I1075342,);
not I_63044 (I1075291,I1075342);
not I_63045 (I1075364,I1075325);
DFFARX1 I_63046 (I519246,I3563,I1075299,I1075390,);
nand I_63047 (I1075398,I1075390,I519252);
not I_63048 (I1075415,I519252);
not I_63049 (I1075432,I519249);
nand I_63050 (I1075449,I519237,I519234);
and I_63051 (I1075466,I519237,I519234);
not I_63052 (I1075483,I519261);
nand I_63053 (I1075500,I1075483,I1075432);
nor I_63054 (I1075273,I1075500,I1075398);
nor I_63055 (I1075531,I1075415,I1075500);
nand I_63056 (I1075276,I1075466,I1075531);
not I_63057 (I1075562,I519234);
nor I_63058 (I1075579,I1075562,I519237);
nor I_63059 (I1075596,I1075579,I519261);
nor I_63060 (I1075613,I1075364,I1075596);
DFFARX1 I_63061 (I1075613,I3563,I1075299,I1075285,);
not I_63062 (I1075644,I1075579);
DFFARX1 I_63063 (I1075644,I3563,I1075299,I1075288,);
and I_63064 (I1075282,I1075390,I1075579);
nor I_63065 (I1075689,I1075562,I519243);
and I_63066 (I1075706,I1075689,I519240);
or I_63067 (I1075723,I1075706,I519255);
DFFARX1 I_63068 (I1075723,I3563,I1075299,I1075749,);
nor I_63069 (I1075757,I1075749,I1075483);
DFFARX1 I_63070 (I1075757,I3563,I1075299,I1075270,);
nand I_63071 (I1075788,I1075749,I1075390);
nand I_63072 (I1075805,I1075483,I1075788);
nor I_63073 (I1075279,I1075805,I1075449);
not I_63074 (I1075860,I3570);
DFFARX1 I_63075 (I166096,I3563,I1075860,I1075886,);
DFFARX1 I_63076 (I1075886,I3563,I1075860,I1075903,);
not I_63077 (I1075852,I1075903);
not I_63078 (I1075925,I1075886);
DFFARX1 I_63079 (I166111,I3563,I1075860,I1075951,);
nand I_63080 (I1075959,I1075951,I166093);
not I_63081 (I1075976,I166093);
not I_63082 (I1075993,I166102);
nand I_63083 (I1076010,I166108,I166099);
and I_63084 (I1076027,I166108,I166099);
not I_63085 (I1076044,I166096);
nand I_63086 (I1076061,I1076044,I1075993);
nor I_63087 (I1075834,I1076061,I1075959);
nor I_63088 (I1076092,I1075976,I1076061);
nand I_63089 (I1075837,I1076027,I1076092);
not I_63090 (I1076123,I166093);
nor I_63091 (I1076140,I1076123,I166108);
nor I_63092 (I1076157,I1076140,I166096);
nor I_63093 (I1076174,I1075925,I1076157);
DFFARX1 I_63094 (I1076174,I3563,I1075860,I1075846,);
not I_63095 (I1076205,I1076140);
DFFARX1 I_63096 (I1076205,I3563,I1075860,I1075849,);
and I_63097 (I1075843,I1075951,I1076140);
nor I_63098 (I1076250,I1076123,I166117);
and I_63099 (I1076267,I1076250,I166114);
or I_63100 (I1076284,I1076267,I166105);
DFFARX1 I_63101 (I1076284,I3563,I1075860,I1076310,);
nor I_63102 (I1076318,I1076310,I1076044);
DFFARX1 I_63103 (I1076318,I3563,I1075860,I1075831,);
nand I_63104 (I1076349,I1076310,I1075951);
nand I_63105 (I1076366,I1076044,I1076349);
nor I_63106 (I1075840,I1076366,I1076010);
not I_63107 (I1076421,I3570);
DFFARX1 I_63108 (I226191,I3563,I1076421,I1076447,);
DFFARX1 I_63109 (I1076447,I3563,I1076421,I1076464,);
not I_63110 (I1076413,I1076464);
not I_63111 (I1076486,I1076447);
DFFARX1 I_63112 (I226206,I3563,I1076421,I1076512,);
nand I_63113 (I1076520,I1076512,I226188);
not I_63114 (I1076537,I226188);
not I_63115 (I1076554,I226197);
nand I_63116 (I1076571,I226203,I226194);
and I_63117 (I1076588,I226203,I226194);
not I_63118 (I1076605,I226191);
nand I_63119 (I1076622,I1076605,I1076554);
nor I_63120 (I1076395,I1076622,I1076520);
nor I_63121 (I1076653,I1076537,I1076622);
nand I_63122 (I1076398,I1076588,I1076653);
not I_63123 (I1076684,I226188);
nor I_63124 (I1076701,I1076684,I226203);
nor I_63125 (I1076718,I1076701,I226191);
nor I_63126 (I1076735,I1076486,I1076718);
DFFARX1 I_63127 (I1076735,I3563,I1076421,I1076407,);
not I_63128 (I1076766,I1076701);
DFFARX1 I_63129 (I1076766,I3563,I1076421,I1076410,);
and I_63130 (I1076404,I1076512,I1076701);
nor I_63131 (I1076811,I1076684,I226212);
and I_63132 (I1076828,I1076811,I226209);
or I_63133 (I1076845,I1076828,I226200);
DFFARX1 I_63134 (I1076845,I3563,I1076421,I1076871,);
nor I_63135 (I1076879,I1076871,I1076605);
DFFARX1 I_63136 (I1076879,I3563,I1076421,I1076392,);
nand I_63137 (I1076910,I1076871,I1076512);
nand I_63138 (I1076927,I1076605,I1076910);
nor I_63139 (I1076401,I1076927,I1076571);
not I_63140 (I1076982,I3570);
DFFARX1 I_63141 (I143614,I3563,I1076982,I1077008,);
DFFARX1 I_63142 (I1077008,I3563,I1076982,I1077025,);
not I_63143 (I1076974,I1077025);
not I_63144 (I1077047,I1077008);
DFFARX1 I_63145 (I143602,I3563,I1076982,I1077073,);
nand I_63146 (I1077081,I1077073,I143617);
not I_63147 (I1077098,I143617);
not I_63148 (I1077115,I143605);
nand I_63149 (I1077132,I143626,I143620);
and I_63150 (I1077149,I143626,I143620);
not I_63151 (I1077166,I143608);
nand I_63152 (I1077183,I1077166,I1077115);
nor I_63153 (I1076956,I1077183,I1077081);
nor I_63154 (I1077214,I1077098,I1077183);
nand I_63155 (I1076959,I1077149,I1077214);
not I_63156 (I1077245,I143611);
nor I_63157 (I1077262,I1077245,I143626);
nor I_63158 (I1077279,I1077262,I143608);
nor I_63159 (I1077296,I1077047,I1077279);
DFFARX1 I_63160 (I1077296,I3563,I1076982,I1076968,);
not I_63161 (I1077327,I1077262);
DFFARX1 I_63162 (I1077327,I3563,I1076982,I1076971,);
and I_63163 (I1076965,I1077073,I1077262);
nor I_63164 (I1077372,I1077245,I143605);
and I_63165 (I1077389,I1077372,I143602);
or I_63166 (I1077406,I1077389,I143623);
DFFARX1 I_63167 (I1077406,I3563,I1076982,I1077432,);
nor I_63168 (I1077440,I1077432,I1077166);
DFFARX1 I_63169 (I1077440,I3563,I1076982,I1076953,);
nand I_63170 (I1077471,I1077432,I1077073);
nand I_63171 (I1077488,I1077166,I1077471);
nor I_63172 (I1076962,I1077488,I1077132);
not I_63173 (I1077543,I3570);
DFFARX1 I_63174 (I424058,I3563,I1077543,I1077569,);
DFFARX1 I_63175 (I1077569,I3563,I1077543,I1077586,);
not I_63176 (I1077535,I1077586);
not I_63177 (I1077608,I1077569);
DFFARX1 I_63178 (I424046,I3563,I1077543,I1077634,);
nand I_63179 (I1077642,I1077634,I424052);
not I_63180 (I1077659,I424052);
not I_63181 (I1077676,I424049);
nand I_63182 (I1077693,I424037,I424034);
and I_63183 (I1077710,I424037,I424034);
not I_63184 (I1077727,I424061);
nand I_63185 (I1077744,I1077727,I1077676);
nor I_63186 (I1077517,I1077744,I1077642);
nor I_63187 (I1077775,I1077659,I1077744);
nand I_63188 (I1077520,I1077710,I1077775);
not I_63189 (I1077806,I424034);
nor I_63190 (I1077823,I1077806,I424037);
nor I_63191 (I1077840,I1077823,I424061);
nor I_63192 (I1077857,I1077608,I1077840);
DFFARX1 I_63193 (I1077857,I3563,I1077543,I1077529,);
not I_63194 (I1077888,I1077823);
DFFARX1 I_63195 (I1077888,I3563,I1077543,I1077532,);
and I_63196 (I1077526,I1077634,I1077823);
nor I_63197 (I1077933,I1077806,I424043);
and I_63198 (I1077950,I1077933,I424040);
or I_63199 (I1077967,I1077950,I424055);
DFFARX1 I_63200 (I1077967,I3563,I1077543,I1077993,);
nor I_63201 (I1078001,I1077993,I1077727);
DFFARX1 I_63202 (I1078001,I3563,I1077543,I1077514,);
nand I_63203 (I1078032,I1077993,I1077634);
nand I_63204 (I1078049,I1077727,I1078032);
nor I_63205 (I1077523,I1078049,I1077693);
not I_63206 (I1078104,I3570);
DFFARX1 I_63207 (I535844,I3563,I1078104,I1078130,);
DFFARX1 I_63208 (I1078130,I3563,I1078104,I1078147,);
not I_63209 (I1078096,I1078147);
not I_63210 (I1078169,I1078130);
DFFARX1 I_63211 (I535841,I3563,I1078104,I1078195,);
nand I_63212 (I1078203,I1078195,I535835);
not I_63213 (I1078220,I535835);
not I_63214 (I1078237,I535847);
nand I_63215 (I1078254,I535850,I535829);
and I_63216 (I1078271,I535850,I535829);
not I_63217 (I1078288,I535826);
nand I_63218 (I1078305,I1078288,I1078237);
nor I_63219 (I1078078,I1078305,I1078203);
nor I_63220 (I1078336,I1078220,I1078305);
nand I_63221 (I1078081,I1078271,I1078336);
not I_63222 (I1078367,I535832);
nor I_63223 (I1078384,I1078367,I535850);
nor I_63224 (I1078401,I1078384,I535826);
nor I_63225 (I1078418,I1078169,I1078401);
DFFARX1 I_63226 (I1078418,I3563,I1078104,I1078090,);
not I_63227 (I1078449,I1078384);
DFFARX1 I_63228 (I1078449,I3563,I1078104,I1078093,);
and I_63229 (I1078087,I1078195,I1078384);
nor I_63230 (I1078494,I1078367,I535826);
and I_63231 (I1078511,I1078494,I535838);
or I_63232 (I1078528,I1078511,I535829);
DFFARX1 I_63233 (I1078528,I3563,I1078104,I1078554,);
nor I_63234 (I1078562,I1078554,I1078288);
DFFARX1 I_63235 (I1078562,I3563,I1078104,I1078075,);
nand I_63236 (I1078593,I1078554,I1078195);
nand I_63237 (I1078610,I1078288,I1078593);
nor I_63238 (I1078084,I1078610,I1078254);
not I_63239 (I1078665,I3570);
DFFARX1 I_63240 (I339667,I3563,I1078665,I1078691,);
DFFARX1 I_63241 (I1078691,I3563,I1078665,I1078708,);
not I_63242 (I1078657,I1078708);
not I_63243 (I1078730,I1078691);
DFFARX1 I_63244 (I339664,I3563,I1078665,I1078756,);
nand I_63245 (I1078764,I1078756,I339658);
not I_63246 (I1078781,I339658);
not I_63247 (I1078798,I339655);
nand I_63248 (I1078815,I339649,I339646);
and I_63249 (I1078832,I339649,I339646);
not I_63250 (I1078849,I339661);
nand I_63251 (I1078866,I1078849,I1078798);
nor I_63252 (I1078639,I1078866,I1078764);
nor I_63253 (I1078897,I1078781,I1078866);
nand I_63254 (I1078642,I1078832,I1078897);
not I_63255 (I1078928,I339673);
nor I_63256 (I1078945,I1078928,I339649);
nor I_63257 (I1078962,I1078945,I339661);
nor I_63258 (I1078979,I1078730,I1078962);
DFFARX1 I_63259 (I1078979,I3563,I1078665,I1078651,);
not I_63260 (I1079010,I1078945);
DFFARX1 I_63261 (I1079010,I3563,I1078665,I1078654,);
and I_63262 (I1078648,I1078756,I1078945);
nor I_63263 (I1079055,I1078928,I339670);
and I_63264 (I1079072,I1079055,I339646);
or I_63265 (I1079089,I1079072,I339652);
DFFARX1 I_63266 (I1079089,I3563,I1078665,I1079115,);
nor I_63267 (I1079123,I1079115,I1078849);
DFFARX1 I_63268 (I1079123,I3563,I1078665,I1078636,);
nand I_63269 (I1079154,I1079115,I1078756);
nand I_63270 (I1079171,I1078849,I1079154);
nor I_63271 (I1078645,I1079171,I1078815);
not I_63272 (I1079226,I3570);
DFFARX1 I_63273 (I1277423,I3563,I1079226,I1079252,);
DFFARX1 I_63274 (I1079252,I3563,I1079226,I1079269,);
not I_63275 (I1079218,I1079269);
not I_63276 (I1079291,I1079252);
DFFARX1 I_63277 (I1277429,I3563,I1079226,I1079317,);
nand I_63278 (I1079325,I1079317,I1277438);
not I_63279 (I1079342,I1277438);
not I_63280 (I1079359,I1277417);
nand I_63281 (I1079376,I1277420,I1277420);
and I_63282 (I1079393,I1277420,I1277420);
not I_63283 (I1079410,I1277432);
nand I_63284 (I1079427,I1079410,I1079359);
nor I_63285 (I1079200,I1079427,I1079325);
nor I_63286 (I1079458,I1079342,I1079427);
nand I_63287 (I1079203,I1079393,I1079458);
not I_63288 (I1079489,I1277426);
nor I_63289 (I1079506,I1079489,I1277420);
nor I_63290 (I1079523,I1079506,I1277432);
nor I_63291 (I1079540,I1079291,I1079523);
DFFARX1 I_63292 (I1079540,I3563,I1079226,I1079212,);
not I_63293 (I1079571,I1079506);
DFFARX1 I_63294 (I1079571,I3563,I1079226,I1079215,);
and I_63295 (I1079209,I1079317,I1079506);
nor I_63296 (I1079616,I1079489,I1277441);
and I_63297 (I1079633,I1079616,I1277417);
or I_63298 (I1079650,I1079633,I1277435);
DFFARX1 I_63299 (I1079650,I3563,I1079226,I1079676,);
nor I_63300 (I1079684,I1079676,I1079410);
DFFARX1 I_63301 (I1079684,I3563,I1079226,I1079197,);
nand I_63302 (I1079715,I1079676,I1079317);
nand I_63303 (I1079732,I1079410,I1079715);
nor I_63304 (I1079206,I1079732,I1079376);
not I_63305 (I1079787,I3570);
DFFARX1 I_63306 (I1092744,I3563,I1079787,I1079813,);
DFFARX1 I_63307 (I1079813,I3563,I1079787,I1079830,);
not I_63308 (I1079779,I1079830);
not I_63309 (I1079852,I1079813);
DFFARX1 I_63310 (I1092735,I3563,I1079787,I1079878,);
nand I_63311 (I1079886,I1079878,I1092732);
not I_63312 (I1079903,I1092732);
not I_63313 (I1079920,I1092741);
nand I_63314 (I1079937,I1092750,I1092732);
and I_63315 (I1079954,I1092750,I1092732);
not I_63316 (I1079971,I1092729);
nand I_63317 (I1079988,I1079971,I1079920);
nor I_63318 (I1079761,I1079988,I1079886);
nor I_63319 (I1080019,I1079903,I1079988);
nand I_63320 (I1079764,I1079954,I1080019);
not I_63321 (I1080050,I1092738);
nor I_63322 (I1080067,I1080050,I1092750);
nor I_63323 (I1080084,I1080067,I1092729);
nor I_63324 (I1080101,I1079852,I1080084);
DFFARX1 I_63325 (I1080101,I3563,I1079787,I1079773,);
not I_63326 (I1080132,I1080067);
DFFARX1 I_63327 (I1080132,I3563,I1079787,I1079776,);
and I_63328 (I1079770,I1079878,I1080067);
nor I_63329 (I1080177,I1080050,I1092753);
and I_63330 (I1080194,I1080177,I1092729);
or I_63331 (I1080211,I1080194,I1092747);
DFFARX1 I_63332 (I1080211,I3563,I1079787,I1080237,);
nor I_63333 (I1080245,I1080237,I1079971);
DFFARX1 I_63334 (I1080245,I3563,I1079787,I1079758,);
nand I_63335 (I1080276,I1080237,I1079878);
nand I_63336 (I1080293,I1079971,I1080276);
nor I_63337 (I1079767,I1080293,I1079937);
not I_63338 (I1080348,I3570);
DFFARX1 I_63339 (I890115,I3563,I1080348,I1080374,);
DFFARX1 I_63340 (I1080374,I3563,I1080348,I1080391,);
not I_63341 (I1080340,I1080391);
not I_63342 (I1080413,I1080374);
DFFARX1 I_63343 (I890112,I3563,I1080348,I1080439,);
nand I_63344 (I1080447,I1080439,I890127);
not I_63345 (I1080464,I890127);
not I_63346 (I1080481,I890124);
nand I_63347 (I1080498,I890121,I890109);
and I_63348 (I1080515,I890121,I890109);
not I_63349 (I1080532,I890106);
nand I_63350 (I1080549,I1080532,I1080481);
nor I_63351 (I1080322,I1080549,I1080447);
nor I_63352 (I1080580,I1080464,I1080549);
nand I_63353 (I1080325,I1080515,I1080580);
not I_63354 (I1080611,I890112);
nor I_63355 (I1080628,I1080611,I890121);
nor I_63356 (I1080645,I1080628,I890106);
nor I_63357 (I1080662,I1080413,I1080645);
DFFARX1 I_63358 (I1080662,I3563,I1080348,I1080334,);
not I_63359 (I1080693,I1080628);
DFFARX1 I_63360 (I1080693,I3563,I1080348,I1080337,);
and I_63361 (I1080331,I1080439,I1080628);
nor I_63362 (I1080738,I1080611,I890118);
and I_63363 (I1080755,I1080738,I890106);
or I_63364 (I1080772,I1080755,I890109);
DFFARX1 I_63365 (I1080772,I3563,I1080348,I1080798,);
nor I_63366 (I1080806,I1080798,I1080532);
DFFARX1 I_63367 (I1080806,I3563,I1080348,I1080319,);
nand I_63368 (I1080837,I1080798,I1080439);
nand I_63369 (I1080854,I1080532,I1080837);
nor I_63370 (I1080328,I1080854,I1080498);
not I_63371 (I1080909,I3570);
DFFARX1 I_63372 (I987873,I3563,I1080909,I1080935,);
DFFARX1 I_63373 (I1080935,I3563,I1080909,I1080952,);
not I_63374 (I1080901,I1080952);
not I_63375 (I1080974,I1080935);
DFFARX1 I_63376 (I987900,I3563,I1080909,I1081000,);
nand I_63377 (I1081008,I1081000,I987891);
not I_63378 (I1081025,I987891);
not I_63379 (I1081042,I987873);
nand I_63380 (I1081059,I987885,I987888);
and I_63381 (I1081076,I987885,I987888);
not I_63382 (I1081093,I987897);
nand I_63383 (I1081110,I1081093,I1081042);
nor I_63384 (I1080883,I1081110,I1081008);
nor I_63385 (I1081141,I1081025,I1081110);
nand I_63386 (I1080886,I1081076,I1081141);
not I_63387 (I1081172,I987882);
nor I_63388 (I1081189,I1081172,I987885);
nor I_63389 (I1081206,I1081189,I987897);
nor I_63390 (I1081223,I1080974,I1081206);
DFFARX1 I_63391 (I1081223,I3563,I1080909,I1080895,);
not I_63392 (I1081254,I1081189);
DFFARX1 I_63393 (I1081254,I3563,I1080909,I1080898,);
and I_63394 (I1080892,I1081000,I1081189);
nor I_63395 (I1081299,I1081172,I987876);
and I_63396 (I1081316,I1081299,I987879);
or I_63397 (I1081333,I1081316,I987894);
DFFARX1 I_63398 (I1081333,I3563,I1080909,I1081359,);
nor I_63399 (I1081367,I1081359,I1081093);
DFFARX1 I_63400 (I1081367,I3563,I1080909,I1080880,);
nand I_63401 (I1081398,I1081359,I1081000);
nand I_63402 (I1081415,I1081093,I1081398);
nor I_63403 (I1080889,I1081415,I1081059);
not I_63404 (I1081470,I3570);
DFFARX1 I_63405 (I235711,I3563,I1081470,I1081496,);
DFFARX1 I_63406 (I1081496,I3563,I1081470,I1081513,);
not I_63407 (I1081462,I1081513);
not I_63408 (I1081535,I1081496);
DFFARX1 I_63409 (I235726,I3563,I1081470,I1081561,);
nand I_63410 (I1081569,I1081561,I235708);
not I_63411 (I1081586,I235708);
not I_63412 (I1081603,I235717);
nand I_63413 (I1081620,I235723,I235714);
and I_63414 (I1081637,I235723,I235714);
not I_63415 (I1081654,I235711);
nand I_63416 (I1081671,I1081654,I1081603);
nor I_63417 (I1081444,I1081671,I1081569);
nor I_63418 (I1081702,I1081586,I1081671);
nand I_63419 (I1081447,I1081637,I1081702);
not I_63420 (I1081733,I235708);
nor I_63421 (I1081750,I1081733,I235723);
nor I_63422 (I1081767,I1081750,I235711);
nor I_63423 (I1081784,I1081535,I1081767);
DFFARX1 I_63424 (I1081784,I3563,I1081470,I1081456,);
not I_63425 (I1081815,I1081750);
DFFARX1 I_63426 (I1081815,I3563,I1081470,I1081459,);
and I_63427 (I1081453,I1081561,I1081750);
nor I_63428 (I1081860,I1081733,I235732);
and I_63429 (I1081877,I1081860,I235729);
or I_63430 (I1081894,I1081877,I235720);
DFFARX1 I_63431 (I1081894,I3563,I1081470,I1081920,);
nor I_63432 (I1081928,I1081920,I1081654);
DFFARX1 I_63433 (I1081928,I3563,I1081470,I1081441,);
nand I_63434 (I1081959,I1081920,I1081561);
nand I_63435 (I1081976,I1081654,I1081959);
nor I_63436 (I1081450,I1081976,I1081620);
not I_63437 (I1082031,I3570);
DFFARX1 I_63438 (I1328115,I3563,I1082031,I1082057,);
DFFARX1 I_63439 (I1082057,I3563,I1082031,I1082074,);
not I_63440 (I1082023,I1082074);
not I_63441 (I1082096,I1082057);
DFFARX1 I_63442 (I1328100,I3563,I1082031,I1082122,);
nand I_63443 (I1082130,I1082122,I1328109);
not I_63444 (I1082147,I1328109);
not I_63445 (I1082164,I1328103);
nand I_63446 (I1082181,I1328121,I1328118);
and I_63447 (I1082198,I1328121,I1328118);
not I_63448 (I1082215,I1328094);
nand I_63449 (I1082232,I1082215,I1082164);
nor I_63450 (I1082005,I1082232,I1082130);
nor I_63451 (I1082263,I1082147,I1082232);
nand I_63452 (I1082008,I1082198,I1082263);
not I_63453 (I1082294,I1328097);
nor I_63454 (I1082311,I1082294,I1328121);
nor I_63455 (I1082328,I1082311,I1328094);
nor I_63456 (I1082345,I1082096,I1082328);
DFFARX1 I_63457 (I1082345,I3563,I1082031,I1082017,);
not I_63458 (I1082376,I1082311);
DFFARX1 I_63459 (I1082376,I3563,I1082031,I1082020,);
and I_63460 (I1082014,I1082122,I1082311);
nor I_63461 (I1082421,I1082294,I1328094);
and I_63462 (I1082438,I1082421,I1328112);
or I_63463 (I1082455,I1082438,I1328106);
DFFARX1 I_63464 (I1082455,I3563,I1082031,I1082481,);
nor I_63465 (I1082489,I1082481,I1082215);
DFFARX1 I_63466 (I1082489,I3563,I1082031,I1082002,);
nand I_63467 (I1082520,I1082481,I1082122);
nand I_63468 (I1082537,I1082215,I1082520);
nor I_63469 (I1082011,I1082537,I1082181);
not I_63470 (I1082592,I3570);
DFFARX1 I_63471 (I867454,I3563,I1082592,I1082618,);
DFFARX1 I_63472 (I1082618,I3563,I1082592,I1082635,);
not I_63473 (I1082584,I1082635);
not I_63474 (I1082657,I1082618);
DFFARX1 I_63475 (I867451,I3563,I1082592,I1082683,);
nand I_63476 (I1082691,I1082683,I867466);
not I_63477 (I1082708,I867466);
not I_63478 (I1082725,I867463);
nand I_63479 (I1082742,I867460,I867448);
and I_63480 (I1082759,I867460,I867448);
not I_63481 (I1082776,I867445);
nand I_63482 (I1082793,I1082776,I1082725);
nor I_63483 (I1082566,I1082793,I1082691);
nor I_63484 (I1082824,I1082708,I1082793);
nand I_63485 (I1082569,I1082759,I1082824);
not I_63486 (I1082855,I867451);
nor I_63487 (I1082872,I1082855,I867460);
nor I_63488 (I1082889,I1082872,I867445);
nor I_63489 (I1082906,I1082657,I1082889);
DFFARX1 I_63490 (I1082906,I3563,I1082592,I1082578,);
not I_63491 (I1082937,I1082872);
DFFARX1 I_63492 (I1082937,I3563,I1082592,I1082581,);
and I_63493 (I1082575,I1082683,I1082872);
nor I_63494 (I1082982,I1082855,I867457);
and I_63495 (I1082999,I1082982,I867445);
or I_63496 (I1083016,I1082999,I867448);
DFFARX1 I_63497 (I1083016,I3563,I1082592,I1083042,);
nor I_63498 (I1083050,I1083042,I1082776);
DFFARX1 I_63499 (I1083050,I3563,I1082592,I1082563,);
nand I_63500 (I1083081,I1083042,I1082683);
nand I_63501 (I1083098,I1082776,I1083081);
nor I_63502 (I1082572,I1083098,I1082742);
not I_63503 (I1083153,I3570);
DFFARX1 I_63504 (I590787,I3563,I1083153,I1083179,);
DFFARX1 I_63505 (I1083179,I3563,I1083153,I1083196,);
not I_63506 (I1083145,I1083196);
not I_63507 (I1083218,I1083179);
DFFARX1 I_63508 (I590802,I3563,I1083153,I1083244,);
nand I_63509 (I1083252,I1083244,I590793);
not I_63510 (I1083269,I590793);
not I_63511 (I1083286,I590799);
nand I_63512 (I1083303,I590796,I590805);
and I_63513 (I1083320,I590796,I590805);
not I_63514 (I1083337,I590790);
nand I_63515 (I1083354,I1083337,I1083286);
nor I_63516 (I1083127,I1083354,I1083252);
nor I_63517 (I1083385,I1083269,I1083354);
nand I_63518 (I1083130,I1083320,I1083385);
not I_63519 (I1083416,I590787);
nor I_63520 (I1083433,I1083416,I590796);
nor I_63521 (I1083450,I1083433,I590790);
nor I_63522 (I1083467,I1083218,I1083450);
DFFARX1 I_63523 (I1083467,I3563,I1083153,I1083139,);
not I_63524 (I1083498,I1083433);
DFFARX1 I_63525 (I1083498,I3563,I1083153,I1083142,);
and I_63526 (I1083136,I1083244,I1083433);
nor I_63527 (I1083543,I1083416,I590811);
and I_63528 (I1083560,I1083543,I590790);
or I_63529 (I1083577,I1083560,I590808);
DFFARX1 I_63530 (I1083577,I3563,I1083153,I1083603,);
nor I_63531 (I1083611,I1083603,I1083337);
DFFARX1 I_63532 (I1083611,I3563,I1083153,I1083124,);
nand I_63533 (I1083642,I1083603,I1083244);
nand I_63534 (I1083659,I1083337,I1083642);
nor I_63535 (I1083133,I1083659,I1083303);
not I_63536 (I1083714,I3570);
DFFARX1 I_63537 (I39274,I3563,I1083714,I1083740,);
DFFARX1 I_63538 (I1083740,I3563,I1083714,I1083757,);
not I_63539 (I1083706,I1083757);
not I_63540 (I1083779,I1083740);
DFFARX1 I_63541 (I39259,I3563,I1083714,I1083805,);
nand I_63542 (I1083813,I1083805,I39271);
not I_63543 (I1083830,I39271);
not I_63544 (I1083847,I39277);
nand I_63545 (I1083864,I39265,I39256);
and I_63546 (I1083881,I39265,I39256);
not I_63547 (I1083898,I39262);
nand I_63548 (I1083915,I1083898,I1083847);
nor I_63549 (I1083688,I1083915,I1083813);
nor I_63550 (I1083946,I1083830,I1083915);
nand I_63551 (I1083691,I1083881,I1083946);
not I_63552 (I1083977,I39268);
nor I_63553 (I1083994,I1083977,I39265);
nor I_63554 (I1084011,I1083994,I39262);
nor I_63555 (I1084028,I1083779,I1084011);
DFFARX1 I_63556 (I1084028,I3563,I1083714,I1083700,);
not I_63557 (I1084059,I1083994);
DFFARX1 I_63558 (I1084059,I3563,I1083714,I1083703,);
and I_63559 (I1083697,I1083805,I1083994);
nor I_63560 (I1084104,I1083977,I39256);
and I_63561 (I1084121,I1084104,I39280);
or I_63562 (I1084138,I1084121,I39259);
DFFARX1 I_63563 (I1084138,I3563,I1083714,I1084164,);
nor I_63564 (I1084172,I1084164,I1083898);
DFFARX1 I_63565 (I1084172,I3563,I1083714,I1083685,);
nand I_63566 (I1084203,I1084164,I1083805);
nand I_63567 (I1084220,I1083898,I1084203);
nor I_63568 (I1083694,I1084220,I1083864);
not I_63569 (I1084275,I3570);
DFFARX1 I_63570 (I117264,I3563,I1084275,I1084301,);
DFFARX1 I_63571 (I1084301,I3563,I1084275,I1084318,);
not I_63572 (I1084267,I1084318);
not I_63573 (I1084340,I1084301);
DFFARX1 I_63574 (I117252,I3563,I1084275,I1084366,);
nand I_63575 (I1084374,I1084366,I117267);
not I_63576 (I1084391,I117267);
not I_63577 (I1084408,I117255);
nand I_63578 (I1084425,I117276,I117270);
and I_63579 (I1084442,I117276,I117270);
not I_63580 (I1084459,I117258);
nand I_63581 (I1084476,I1084459,I1084408);
nor I_63582 (I1084249,I1084476,I1084374);
nor I_63583 (I1084507,I1084391,I1084476);
nand I_63584 (I1084252,I1084442,I1084507);
not I_63585 (I1084538,I117261);
nor I_63586 (I1084555,I1084538,I117276);
nor I_63587 (I1084572,I1084555,I117258);
nor I_63588 (I1084589,I1084340,I1084572);
DFFARX1 I_63589 (I1084589,I3563,I1084275,I1084261,);
not I_63590 (I1084620,I1084555);
DFFARX1 I_63591 (I1084620,I3563,I1084275,I1084264,);
and I_63592 (I1084258,I1084366,I1084555);
nor I_63593 (I1084665,I1084538,I117255);
and I_63594 (I1084682,I1084665,I117252);
or I_63595 (I1084699,I1084682,I117273);
DFFARX1 I_63596 (I1084699,I3563,I1084275,I1084725,);
nor I_63597 (I1084733,I1084725,I1084459);
DFFARX1 I_63598 (I1084733,I3563,I1084275,I1084246,);
nand I_63599 (I1084764,I1084725,I1084366);
nand I_63600 (I1084781,I1084459,I1084764);
nor I_63601 (I1084255,I1084781,I1084425);
not I_63602 (I1084836,I3570);
DFFARX1 I_63603 (I243446,I3563,I1084836,I1084862,);
DFFARX1 I_63604 (I1084862,I3563,I1084836,I1084879,);
not I_63605 (I1084828,I1084879);
not I_63606 (I1084901,I1084862);
DFFARX1 I_63607 (I243461,I3563,I1084836,I1084927,);
nand I_63608 (I1084935,I1084927,I243443);
not I_63609 (I1084952,I243443);
not I_63610 (I1084969,I243452);
nand I_63611 (I1084986,I243458,I243449);
and I_63612 (I1085003,I243458,I243449);
not I_63613 (I1085020,I243446);
nand I_63614 (I1085037,I1085020,I1084969);
nor I_63615 (I1084810,I1085037,I1084935);
nor I_63616 (I1085068,I1084952,I1085037);
nand I_63617 (I1084813,I1085003,I1085068);
not I_63618 (I1085099,I243443);
nor I_63619 (I1085116,I1085099,I243458);
nor I_63620 (I1085133,I1085116,I243446);
nor I_63621 (I1085150,I1084901,I1085133);
DFFARX1 I_63622 (I1085150,I3563,I1084836,I1084822,);
not I_63623 (I1085181,I1085116);
DFFARX1 I_63624 (I1085181,I3563,I1084836,I1084825,);
and I_63625 (I1084819,I1084927,I1085116);
nor I_63626 (I1085226,I1085099,I243467);
and I_63627 (I1085243,I1085226,I243464);
or I_63628 (I1085260,I1085243,I243455);
DFFARX1 I_63629 (I1085260,I3563,I1084836,I1085286,);
nor I_63630 (I1085294,I1085286,I1085020);
DFFARX1 I_63631 (I1085294,I3563,I1084836,I1084807,);
nand I_63632 (I1085325,I1085286,I1084927);
nand I_63633 (I1085342,I1085020,I1085325);
nor I_63634 (I1084816,I1085342,I1084986);
not I_63635 (I1085397,I3570);
DFFARX1 I_63636 (I376030,I3563,I1085397,I1085423,);
DFFARX1 I_63637 (I1085423,I3563,I1085397,I1085440,);
not I_63638 (I1085389,I1085440);
not I_63639 (I1085462,I1085423);
DFFARX1 I_63640 (I376027,I3563,I1085397,I1085488,);
nand I_63641 (I1085496,I1085488,I376021);
not I_63642 (I1085513,I376021);
not I_63643 (I1085530,I376018);
nand I_63644 (I1085547,I376012,I376009);
and I_63645 (I1085564,I376012,I376009);
not I_63646 (I1085581,I376024);
nand I_63647 (I1085598,I1085581,I1085530);
nor I_63648 (I1085371,I1085598,I1085496);
nor I_63649 (I1085629,I1085513,I1085598);
nand I_63650 (I1085374,I1085564,I1085629);
not I_63651 (I1085660,I376036);
nor I_63652 (I1085677,I1085660,I376012);
nor I_63653 (I1085694,I1085677,I376024);
nor I_63654 (I1085711,I1085462,I1085694);
DFFARX1 I_63655 (I1085711,I3563,I1085397,I1085383,);
not I_63656 (I1085742,I1085677);
DFFARX1 I_63657 (I1085742,I3563,I1085397,I1085386,);
and I_63658 (I1085380,I1085488,I1085677);
nor I_63659 (I1085787,I1085660,I376033);
and I_63660 (I1085804,I1085787,I376009);
or I_63661 (I1085821,I1085804,I376015);
DFFARX1 I_63662 (I1085821,I3563,I1085397,I1085847,);
nor I_63663 (I1085855,I1085847,I1085581);
DFFARX1 I_63664 (I1085855,I3563,I1085397,I1085368,);
nand I_63665 (I1085886,I1085847,I1085488);
nand I_63666 (I1085903,I1085581,I1085886);
nor I_63667 (I1085377,I1085903,I1085547);
not I_63668 (I1085958,I3570);
DFFARX1 I_63669 (I1117598,I3563,I1085958,I1085984,);
DFFARX1 I_63670 (I1085984,I3563,I1085958,I1086001,);
not I_63671 (I1085950,I1086001);
not I_63672 (I1086023,I1085984);
DFFARX1 I_63673 (I1117589,I3563,I1085958,I1086049,);
nand I_63674 (I1086057,I1086049,I1117586);
not I_63675 (I1086074,I1117586);
not I_63676 (I1086091,I1117595);
nand I_63677 (I1086108,I1117604,I1117586);
and I_63678 (I1086125,I1117604,I1117586);
not I_63679 (I1086142,I1117583);
nand I_63680 (I1086159,I1086142,I1086091);
nor I_63681 (I1085932,I1086159,I1086057);
nor I_63682 (I1086190,I1086074,I1086159);
nand I_63683 (I1085935,I1086125,I1086190);
not I_63684 (I1086221,I1117592);
nor I_63685 (I1086238,I1086221,I1117604);
nor I_63686 (I1086255,I1086238,I1117583);
nor I_63687 (I1086272,I1086023,I1086255);
DFFARX1 I_63688 (I1086272,I3563,I1085958,I1085944,);
not I_63689 (I1086303,I1086238);
DFFARX1 I_63690 (I1086303,I3563,I1085958,I1085947,);
and I_63691 (I1085941,I1086049,I1086238);
nor I_63692 (I1086348,I1086221,I1117607);
and I_63693 (I1086365,I1086348,I1117583);
or I_63694 (I1086382,I1086365,I1117601);
DFFARX1 I_63695 (I1086382,I3563,I1085958,I1086408,);
nor I_63696 (I1086416,I1086408,I1086142);
DFFARX1 I_63697 (I1086416,I3563,I1085958,I1085929,);
nand I_63698 (I1086447,I1086408,I1086049);
nand I_63699 (I1086464,I1086142,I1086447);
nor I_63700 (I1085938,I1086464,I1086108);
not I_63701 (I1086519,I3570);
DFFARX1 I_63702 (I3020,I3563,I1086519,I1086545,);
DFFARX1 I_63703 (I1086545,I3563,I1086519,I1086562,);
not I_63704 (I1086511,I1086562);
not I_63705 (I1086584,I1086545);
DFFARX1 I_63706 (I3124,I3563,I1086519,I1086610,);
nand I_63707 (I1086618,I1086610,I1580);
not I_63708 (I1086635,I1580);
not I_63709 (I1086652,I2748);
nand I_63710 (I1086669,I3444,I2740);
and I_63711 (I1086686,I3444,I2740);
not I_63712 (I1086703,I1740);
nand I_63713 (I1086720,I1086703,I1086652);
nor I_63714 (I1086493,I1086720,I1086618);
nor I_63715 (I1086751,I1086635,I1086720);
nand I_63716 (I1086496,I1086686,I1086751);
not I_63717 (I1086782,I3460);
nor I_63718 (I1086799,I1086782,I3444);
nor I_63719 (I1086816,I1086799,I1740);
nor I_63720 (I1086833,I1086584,I1086816);
DFFARX1 I_63721 (I1086833,I3563,I1086519,I1086505,);
not I_63722 (I1086864,I1086799);
DFFARX1 I_63723 (I1086864,I3563,I1086519,I1086508,);
and I_63724 (I1086502,I1086610,I1086799);
nor I_63725 (I1086909,I1086782,I3132);
and I_63726 (I1086926,I1086909,I2972);
or I_63727 (I1086943,I1086926,I1788);
DFFARX1 I_63728 (I1086943,I3563,I1086519,I1086969,);
nor I_63729 (I1086977,I1086969,I1086703);
DFFARX1 I_63730 (I1086977,I3563,I1086519,I1086490,);
nand I_63731 (I1087008,I1086969,I1086610);
nand I_63732 (I1087025,I1086703,I1087008);
nor I_63733 (I1086499,I1087025,I1086669);
not I_63734 (I1087080,I3570);
DFFARX1 I_63735 (I1215280,I3563,I1087080,I1087106,);
DFFARX1 I_63736 (I1087106,I3563,I1087080,I1087123,);
not I_63737 (I1087072,I1087123);
not I_63738 (I1087145,I1087106);
DFFARX1 I_63739 (I1215271,I3563,I1087080,I1087171,);
nand I_63740 (I1087179,I1087171,I1215268);
not I_63741 (I1087196,I1215268);
not I_63742 (I1087213,I1215277);
nand I_63743 (I1087230,I1215286,I1215268);
and I_63744 (I1087247,I1215286,I1215268);
not I_63745 (I1087264,I1215265);
nand I_63746 (I1087281,I1087264,I1087213);
nor I_63747 (I1087054,I1087281,I1087179);
nor I_63748 (I1087312,I1087196,I1087281);
nand I_63749 (I1087057,I1087247,I1087312);
not I_63750 (I1087343,I1215274);
nor I_63751 (I1087360,I1087343,I1215286);
nor I_63752 (I1087377,I1087360,I1215265);
nor I_63753 (I1087394,I1087145,I1087377);
DFFARX1 I_63754 (I1087394,I3563,I1087080,I1087066,);
not I_63755 (I1087425,I1087360);
DFFARX1 I_63756 (I1087425,I3563,I1087080,I1087069,);
and I_63757 (I1087063,I1087171,I1087360);
nor I_63758 (I1087470,I1087343,I1215289);
and I_63759 (I1087487,I1087470,I1215265);
or I_63760 (I1087504,I1087487,I1215283);
DFFARX1 I_63761 (I1087504,I3563,I1087080,I1087530,);
nor I_63762 (I1087538,I1087530,I1087264);
DFFARX1 I_63763 (I1087538,I3563,I1087080,I1087051,);
nand I_63764 (I1087569,I1087530,I1087171);
nand I_63765 (I1087586,I1087264,I1087569);
nor I_63766 (I1087060,I1087586,I1087230);
not I_63767 (I1087641,I3570);
DFFARX1 I_63768 (I574519,I3563,I1087641,I1087667,);
DFFARX1 I_63769 (I1087667,I3563,I1087641,I1087684,);
not I_63770 (I1087633,I1087684);
not I_63771 (I1087706,I1087667);
DFFARX1 I_63772 (I574516,I3563,I1087641,I1087732,);
nand I_63773 (I1087740,I1087732,I574510);
not I_63774 (I1087757,I574510);
not I_63775 (I1087774,I574522);
nand I_63776 (I1087791,I574525,I574504);
and I_63777 (I1087808,I574525,I574504);
not I_63778 (I1087825,I574501);
nand I_63779 (I1087842,I1087825,I1087774);
nor I_63780 (I1087615,I1087842,I1087740);
nor I_63781 (I1087873,I1087757,I1087842);
nand I_63782 (I1087618,I1087808,I1087873);
not I_63783 (I1087904,I574507);
nor I_63784 (I1087921,I1087904,I574525);
nor I_63785 (I1087938,I1087921,I574501);
nor I_63786 (I1087955,I1087706,I1087938);
DFFARX1 I_63787 (I1087955,I3563,I1087641,I1087627,);
not I_63788 (I1087986,I1087921);
DFFARX1 I_63789 (I1087986,I3563,I1087641,I1087630,);
and I_63790 (I1087624,I1087732,I1087921);
nor I_63791 (I1088031,I1087904,I574501);
and I_63792 (I1088048,I1088031,I574513);
or I_63793 (I1088065,I1088048,I574504);
DFFARX1 I_63794 (I1088065,I3563,I1087641,I1088091,);
nor I_63795 (I1088099,I1088091,I1087825);
DFFARX1 I_63796 (I1088099,I3563,I1087641,I1087612,);
nand I_63797 (I1088130,I1088091,I1087732);
nand I_63798 (I1088147,I1087825,I1088130);
nor I_63799 (I1087621,I1088147,I1087791);
not I_63800 (I1088202,I3570);
DFFARX1 I_63801 (I628935,I3563,I1088202,I1088228,);
DFFARX1 I_63802 (I1088228,I3563,I1088202,I1088245,);
not I_63803 (I1088194,I1088245);
not I_63804 (I1088267,I1088228);
DFFARX1 I_63805 (I628950,I3563,I1088202,I1088293,);
nand I_63806 (I1088301,I1088293,I628941);
not I_63807 (I1088318,I628941);
not I_63808 (I1088335,I628947);
nand I_63809 (I1088352,I628944,I628953);
and I_63810 (I1088369,I628944,I628953);
not I_63811 (I1088386,I628938);
nand I_63812 (I1088403,I1088386,I1088335);
nor I_63813 (I1088176,I1088403,I1088301);
nor I_63814 (I1088434,I1088318,I1088403);
nand I_63815 (I1088179,I1088369,I1088434);
not I_63816 (I1088465,I628935);
nor I_63817 (I1088482,I1088465,I628944);
nor I_63818 (I1088499,I1088482,I628938);
nor I_63819 (I1088516,I1088267,I1088499);
DFFARX1 I_63820 (I1088516,I3563,I1088202,I1088188,);
not I_63821 (I1088547,I1088482);
DFFARX1 I_63822 (I1088547,I3563,I1088202,I1088191,);
and I_63823 (I1088185,I1088293,I1088482);
nor I_63824 (I1088592,I1088465,I628959);
and I_63825 (I1088609,I1088592,I628938);
or I_63826 (I1088626,I1088609,I628956);
DFFARX1 I_63827 (I1088626,I3563,I1088202,I1088652,);
nor I_63828 (I1088660,I1088652,I1088386);
DFFARX1 I_63829 (I1088660,I3563,I1088202,I1088173,);
nand I_63830 (I1088691,I1088652,I1088293);
nand I_63831 (I1088708,I1088386,I1088691);
nor I_63832 (I1088182,I1088708,I1088352);
not I_63833 (I1088763,I3570);
DFFARX1 I_63834 (I484442,I3563,I1088763,I1088789,);
DFFARX1 I_63835 (I1088789,I3563,I1088763,I1088806,);
not I_63836 (I1088755,I1088806);
not I_63837 (I1088828,I1088789);
DFFARX1 I_63838 (I484430,I3563,I1088763,I1088854,);
nand I_63839 (I1088862,I1088854,I484436);
not I_63840 (I1088879,I484436);
not I_63841 (I1088896,I484433);
nand I_63842 (I1088913,I484421,I484418);
and I_63843 (I1088930,I484421,I484418);
not I_63844 (I1088947,I484445);
nand I_63845 (I1088964,I1088947,I1088896);
nor I_63846 (I1088737,I1088964,I1088862);
nor I_63847 (I1088995,I1088879,I1088964);
nand I_63848 (I1088740,I1088930,I1088995);
not I_63849 (I1089026,I484418);
nor I_63850 (I1089043,I1089026,I484421);
nor I_63851 (I1089060,I1089043,I484445);
nor I_63852 (I1089077,I1088828,I1089060);
DFFARX1 I_63853 (I1089077,I3563,I1088763,I1088749,);
not I_63854 (I1089108,I1089043);
DFFARX1 I_63855 (I1089108,I3563,I1088763,I1088752,);
and I_63856 (I1088746,I1088854,I1089043);
nor I_63857 (I1089153,I1089026,I484427);
and I_63858 (I1089170,I1089153,I484424);
or I_63859 (I1089187,I1089170,I484439);
DFFARX1 I_63860 (I1089187,I3563,I1088763,I1089213,);
nor I_63861 (I1089221,I1089213,I1088947);
DFFARX1 I_63862 (I1089221,I3563,I1088763,I1088734,);
nand I_63863 (I1089252,I1089213,I1088854);
nand I_63864 (I1089269,I1088947,I1089252);
nor I_63865 (I1088743,I1089269,I1088913);
not I_63866 (I1089324,I3570);
DFFARX1 I_63867 (I318587,I3563,I1089324,I1089350,);
DFFARX1 I_63868 (I1089350,I3563,I1089324,I1089367,);
not I_63869 (I1089316,I1089367);
not I_63870 (I1089389,I1089350);
DFFARX1 I_63871 (I318584,I3563,I1089324,I1089415,);
nand I_63872 (I1089423,I1089415,I318578);
not I_63873 (I1089440,I318578);
not I_63874 (I1089457,I318575);
nand I_63875 (I1089474,I318569,I318566);
and I_63876 (I1089491,I318569,I318566);
not I_63877 (I1089508,I318581);
nand I_63878 (I1089525,I1089508,I1089457);
nor I_63879 (I1089298,I1089525,I1089423);
nor I_63880 (I1089556,I1089440,I1089525);
nand I_63881 (I1089301,I1089491,I1089556);
not I_63882 (I1089587,I318593);
nor I_63883 (I1089604,I1089587,I318569);
nor I_63884 (I1089621,I1089604,I318581);
nor I_63885 (I1089638,I1089389,I1089621);
DFFARX1 I_63886 (I1089638,I3563,I1089324,I1089310,);
not I_63887 (I1089669,I1089604);
DFFARX1 I_63888 (I1089669,I3563,I1089324,I1089313,);
and I_63889 (I1089307,I1089415,I1089604);
nor I_63890 (I1089714,I1089587,I318590);
and I_63891 (I1089731,I1089714,I318566);
or I_63892 (I1089748,I1089731,I318572);
DFFARX1 I_63893 (I1089748,I3563,I1089324,I1089774,);
nor I_63894 (I1089782,I1089774,I1089508);
DFFARX1 I_63895 (I1089782,I3563,I1089324,I1089295,);
nand I_63896 (I1089813,I1089774,I1089415);
nand I_63897 (I1089830,I1089508,I1089813);
nor I_63898 (I1089304,I1089830,I1089474);
not I_63899 (I1089885,I3570);
DFFARX1 I_63900 (I184541,I3563,I1089885,I1089911,);
DFFARX1 I_63901 (I1089911,I3563,I1089885,I1089928,);
not I_63902 (I1089877,I1089928);
not I_63903 (I1089950,I1089911);
DFFARX1 I_63904 (I184556,I3563,I1089885,I1089976,);
nand I_63905 (I1089984,I1089976,I184538);
not I_63906 (I1090001,I184538);
not I_63907 (I1090018,I184547);
nand I_63908 (I1090035,I184553,I184544);
and I_63909 (I1090052,I184553,I184544);
not I_63910 (I1090069,I184541);
nand I_63911 (I1090086,I1090069,I1090018);
nor I_63912 (I1089859,I1090086,I1089984);
nor I_63913 (I1090117,I1090001,I1090086);
nand I_63914 (I1089862,I1090052,I1090117);
not I_63915 (I1090148,I184538);
nor I_63916 (I1090165,I1090148,I184553);
nor I_63917 (I1090182,I1090165,I184541);
nor I_63918 (I1090199,I1089950,I1090182);
DFFARX1 I_63919 (I1090199,I3563,I1089885,I1089871,);
not I_63920 (I1090230,I1090165);
DFFARX1 I_63921 (I1090230,I3563,I1089885,I1089874,);
and I_63922 (I1089868,I1089976,I1090165);
nor I_63923 (I1090275,I1090148,I184562);
and I_63924 (I1090292,I1090275,I184559);
or I_63925 (I1090309,I1090292,I184550);
DFFARX1 I_63926 (I1090309,I3563,I1089885,I1090335,);
nor I_63927 (I1090343,I1090335,I1090069);
DFFARX1 I_63928 (I1090343,I3563,I1089885,I1089856,);
nand I_63929 (I1090374,I1090335,I1089976);
nand I_63930 (I1090391,I1090069,I1090374);
nor I_63931 (I1089865,I1090391,I1090035);
not I_63932 (I1090449,I3570);
DFFARX1 I_63933 (I961393,I3563,I1090449,I1090475,);
and I_63934 (I1090483,I1090475,I961387);
DFFARX1 I_63935 (I1090483,I3563,I1090449,I1090432,);
DFFARX1 I_63936 (I961405,I3563,I1090449,I1090523,);
not I_63937 (I1090531,I961396);
not I_63938 (I1090548,I961408);
nand I_63939 (I1090565,I1090548,I1090531);
nor I_63940 (I1090420,I1090523,I1090565);
DFFARX1 I_63941 (I1090565,I3563,I1090449,I1090605,);
not I_63942 (I1090441,I1090605);
not I_63943 (I1090627,I961414);
nand I_63944 (I1090644,I1090548,I1090627);
DFFARX1 I_63945 (I1090644,I3563,I1090449,I1090670,);
not I_63946 (I1090678,I1090670);
not I_63947 (I1090695,I961390);
nand I_63948 (I1090712,I1090695,I961411);
and I_63949 (I1090729,I1090531,I1090712);
nor I_63950 (I1090746,I1090644,I1090729);
DFFARX1 I_63951 (I1090746,I3563,I1090449,I1090417,);
DFFARX1 I_63952 (I1090729,I3563,I1090449,I1090438,);
nor I_63953 (I1090791,I961390,I961402);
nor I_63954 (I1090429,I1090644,I1090791);
or I_63955 (I1090822,I961390,I961402);
nor I_63956 (I1090839,I961387,I961399);
DFFARX1 I_63957 (I1090839,I3563,I1090449,I1090865,);
not I_63958 (I1090873,I1090865);
nor I_63959 (I1090435,I1090873,I1090678);
nand I_63960 (I1090904,I1090873,I1090523);
not I_63961 (I1090921,I961387);
nand I_63962 (I1090938,I1090921,I1090627);
nand I_63963 (I1090955,I1090873,I1090938);
nand I_63964 (I1090426,I1090955,I1090904);
nand I_63965 (I1090423,I1090938,I1090822);
not I_63966 (I1091027,I3570);
DFFARX1 I_63967 (I1015657,I3563,I1091027,I1091053,);
and I_63968 (I1091061,I1091053,I1015651);
DFFARX1 I_63969 (I1091061,I3563,I1091027,I1091010,);
DFFARX1 I_63970 (I1015669,I3563,I1091027,I1091101,);
not I_63971 (I1091109,I1015660);
not I_63972 (I1091126,I1015672);
nand I_63973 (I1091143,I1091126,I1091109);
nor I_63974 (I1090998,I1091101,I1091143);
DFFARX1 I_63975 (I1091143,I3563,I1091027,I1091183,);
not I_63976 (I1091019,I1091183);
not I_63977 (I1091205,I1015678);
nand I_63978 (I1091222,I1091126,I1091205);
DFFARX1 I_63979 (I1091222,I3563,I1091027,I1091248,);
not I_63980 (I1091256,I1091248);
not I_63981 (I1091273,I1015654);
nand I_63982 (I1091290,I1091273,I1015675);
and I_63983 (I1091307,I1091109,I1091290);
nor I_63984 (I1091324,I1091222,I1091307);
DFFARX1 I_63985 (I1091324,I3563,I1091027,I1090995,);
DFFARX1 I_63986 (I1091307,I3563,I1091027,I1091016,);
nor I_63987 (I1091369,I1015654,I1015666);
nor I_63988 (I1091007,I1091222,I1091369);
or I_63989 (I1091400,I1015654,I1015666);
nor I_63990 (I1091417,I1015651,I1015663);
DFFARX1 I_63991 (I1091417,I3563,I1091027,I1091443,);
not I_63992 (I1091451,I1091443);
nor I_63993 (I1091013,I1091451,I1091256);
nand I_63994 (I1091482,I1091451,I1091101);
not I_63995 (I1091499,I1015651);
nand I_63996 (I1091516,I1091499,I1091205);
nand I_63997 (I1091533,I1091451,I1091516);
nand I_63998 (I1091004,I1091533,I1091482);
nand I_63999 (I1091001,I1091516,I1091400);
not I_64000 (I1091605,I3570);
DFFARX1 I_64001 (I367077,I3563,I1091605,I1091631,);
and I_64002 (I1091639,I1091631,I367062);
DFFARX1 I_64003 (I1091639,I3563,I1091605,I1091588,);
DFFARX1 I_64004 (I367068,I3563,I1091605,I1091679,);
not I_64005 (I1091687,I367050);
not I_64006 (I1091704,I367071);
nand I_64007 (I1091721,I1091704,I1091687);
nor I_64008 (I1091576,I1091679,I1091721);
DFFARX1 I_64009 (I1091721,I3563,I1091605,I1091761,);
not I_64010 (I1091597,I1091761);
not I_64011 (I1091783,I367074);
nand I_64012 (I1091800,I1091704,I1091783);
DFFARX1 I_64013 (I1091800,I3563,I1091605,I1091826,);
not I_64014 (I1091834,I1091826);
not I_64015 (I1091851,I367065);
nand I_64016 (I1091868,I1091851,I367053);
and I_64017 (I1091885,I1091687,I1091868);
nor I_64018 (I1091902,I1091800,I1091885);
DFFARX1 I_64019 (I1091902,I3563,I1091605,I1091573,);
DFFARX1 I_64020 (I1091885,I3563,I1091605,I1091594,);
nor I_64021 (I1091947,I367065,I367059);
nor I_64022 (I1091585,I1091800,I1091947);
or I_64023 (I1091978,I367065,I367059);
nor I_64024 (I1091995,I367056,I367050);
DFFARX1 I_64025 (I1091995,I3563,I1091605,I1092021,);
not I_64026 (I1092029,I1092021);
nor I_64027 (I1091591,I1092029,I1091834);
nand I_64028 (I1092060,I1092029,I1091679);
not I_64029 (I1092077,I367056);
nand I_64030 (I1092094,I1092077,I1091783);
nand I_64031 (I1092111,I1092029,I1092094);
nand I_64032 (I1091582,I1092111,I1092060);
nand I_64033 (I1091579,I1092094,I1091978);
not I_64034 (I1092183,I3570);
DFFARX1 I_64035 (I35567,I3563,I1092183,I1092209,);
and I_64036 (I1092217,I1092209,I35570);
DFFARX1 I_64037 (I1092217,I3563,I1092183,I1092166,);
DFFARX1 I_64038 (I35570,I3563,I1092183,I1092257,);
not I_64039 (I1092265,I35573);
not I_64040 (I1092282,I35588);
nand I_64041 (I1092299,I1092282,I1092265);
nor I_64042 (I1092154,I1092257,I1092299);
DFFARX1 I_64043 (I1092299,I3563,I1092183,I1092339,);
not I_64044 (I1092175,I1092339);
not I_64045 (I1092361,I35582);
nand I_64046 (I1092378,I1092282,I1092361);
DFFARX1 I_64047 (I1092378,I3563,I1092183,I1092404,);
not I_64048 (I1092412,I1092404);
not I_64049 (I1092429,I35585);
nand I_64050 (I1092446,I1092429,I35567);
and I_64051 (I1092463,I1092265,I1092446);
nor I_64052 (I1092480,I1092378,I1092463);
DFFARX1 I_64053 (I1092480,I3563,I1092183,I1092151,);
DFFARX1 I_64054 (I1092463,I3563,I1092183,I1092172,);
nor I_64055 (I1092525,I35585,I35579);
nor I_64056 (I1092163,I1092378,I1092525);
or I_64057 (I1092556,I35585,I35579);
nor I_64058 (I1092573,I35576,I35591);
DFFARX1 I_64059 (I1092573,I3563,I1092183,I1092599,);
not I_64060 (I1092607,I1092599);
nor I_64061 (I1092169,I1092607,I1092412);
nand I_64062 (I1092638,I1092607,I1092257);
not I_64063 (I1092655,I35576);
nand I_64064 (I1092672,I1092655,I1092361);
nand I_64065 (I1092689,I1092607,I1092672);
nand I_64066 (I1092160,I1092689,I1092638);
nand I_64067 (I1092157,I1092672,I1092556);
not I_64068 (I1092761,I3570);
DFFARX1 I_64069 (I792524,I3563,I1092761,I1092787,);
and I_64070 (I1092795,I1092787,I792512);
DFFARX1 I_64071 (I1092795,I3563,I1092761,I1092744,);
DFFARX1 I_64072 (I792515,I3563,I1092761,I1092835,);
not I_64073 (I1092843,I792509);
not I_64074 (I1092860,I792533);
nand I_64075 (I1092877,I1092860,I1092843);
nor I_64076 (I1092732,I1092835,I1092877);
DFFARX1 I_64077 (I1092877,I3563,I1092761,I1092917,);
not I_64078 (I1092753,I1092917);
not I_64079 (I1092939,I792521);
nand I_64080 (I1092956,I1092860,I1092939);
DFFARX1 I_64081 (I1092956,I3563,I1092761,I1092982,);
not I_64082 (I1092990,I1092982);
not I_64083 (I1093007,I792530);
nand I_64084 (I1093024,I1093007,I792527);
and I_64085 (I1093041,I1092843,I1093024);
nor I_64086 (I1093058,I1092956,I1093041);
DFFARX1 I_64087 (I1093058,I3563,I1092761,I1092729,);
DFFARX1 I_64088 (I1093041,I3563,I1092761,I1092750,);
nor I_64089 (I1093103,I792530,I792518);
nor I_64090 (I1092741,I1092956,I1093103);
or I_64091 (I1093134,I792530,I792518);
nor I_64092 (I1093151,I792509,I792512);
DFFARX1 I_64093 (I1093151,I3563,I1092761,I1093177,);
not I_64094 (I1093185,I1093177);
nor I_64095 (I1092747,I1093185,I1092990);
nand I_64096 (I1093216,I1093185,I1092835);
not I_64097 (I1093233,I792509);
nand I_64098 (I1093250,I1093233,I1092939);
nand I_64099 (I1093267,I1093185,I1093250);
nand I_64100 (I1092738,I1093267,I1093216);
nand I_64101 (I1092735,I1093250,I1093134);
not I_64102 (I1093339,I3570);
DFFARX1 I_64103 (I805240,I3563,I1093339,I1093365,);
and I_64104 (I1093373,I1093365,I805228);
DFFARX1 I_64105 (I1093373,I3563,I1093339,I1093322,);
DFFARX1 I_64106 (I805231,I3563,I1093339,I1093413,);
not I_64107 (I1093421,I805225);
not I_64108 (I1093438,I805249);
nand I_64109 (I1093455,I1093438,I1093421);
nor I_64110 (I1093310,I1093413,I1093455);
DFFARX1 I_64111 (I1093455,I3563,I1093339,I1093495,);
not I_64112 (I1093331,I1093495);
not I_64113 (I1093517,I805237);
nand I_64114 (I1093534,I1093438,I1093517);
DFFARX1 I_64115 (I1093534,I3563,I1093339,I1093560,);
not I_64116 (I1093568,I1093560);
not I_64117 (I1093585,I805246);
nand I_64118 (I1093602,I1093585,I805243);
and I_64119 (I1093619,I1093421,I1093602);
nor I_64120 (I1093636,I1093534,I1093619);
DFFARX1 I_64121 (I1093636,I3563,I1093339,I1093307,);
DFFARX1 I_64122 (I1093619,I3563,I1093339,I1093328,);
nor I_64123 (I1093681,I805246,I805234);
nor I_64124 (I1093319,I1093534,I1093681);
or I_64125 (I1093712,I805246,I805234);
nor I_64126 (I1093729,I805225,I805228);
DFFARX1 I_64127 (I1093729,I3563,I1093339,I1093755,);
not I_64128 (I1093763,I1093755);
nor I_64129 (I1093325,I1093763,I1093568);
nand I_64130 (I1093794,I1093763,I1093413);
not I_64131 (I1093811,I805225);
nand I_64132 (I1093828,I1093811,I1093517);
nand I_64133 (I1093845,I1093763,I1093828);
nand I_64134 (I1093316,I1093845,I1093794);
nand I_64135 (I1093313,I1093828,I1093712);
not I_64136 (I1093917,I3570);
DFFARX1 I_64137 (I351794,I3563,I1093917,I1093943,);
and I_64138 (I1093951,I1093943,I351779);
DFFARX1 I_64139 (I1093951,I3563,I1093917,I1093900,);
DFFARX1 I_64140 (I351785,I3563,I1093917,I1093991,);
not I_64141 (I1093999,I351767);
not I_64142 (I1094016,I351788);
nand I_64143 (I1094033,I1094016,I1093999);
nor I_64144 (I1093888,I1093991,I1094033);
DFFARX1 I_64145 (I1094033,I3563,I1093917,I1094073,);
not I_64146 (I1093909,I1094073);
not I_64147 (I1094095,I351791);
nand I_64148 (I1094112,I1094016,I1094095);
DFFARX1 I_64149 (I1094112,I3563,I1093917,I1094138,);
not I_64150 (I1094146,I1094138);
not I_64151 (I1094163,I351782);
nand I_64152 (I1094180,I1094163,I351770);
and I_64153 (I1094197,I1093999,I1094180);
nor I_64154 (I1094214,I1094112,I1094197);
DFFARX1 I_64155 (I1094214,I3563,I1093917,I1093885,);
DFFARX1 I_64156 (I1094197,I3563,I1093917,I1093906,);
nor I_64157 (I1094259,I351782,I351776);
nor I_64158 (I1093897,I1094112,I1094259);
or I_64159 (I1094290,I351782,I351776);
nor I_64160 (I1094307,I351773,I351767);
DFFARX1 I_64161 (I1094307,I3563,I1093917,I1094333,);
not I_64162 (I1094341,I1094333);
nor I_64163 (I1093903,I1094341,I1094146);
nand I_64164 (I1094372,I1094341,I1093991);
not I_64165 (I1094389,I351773);
nand I_64166 (I1094406,I1094389,I1094095);
nand I_64167 (I1094423,I1094341,I1094406);
nand I_64168 (I1093894,I1094423,I1094372);
nand I_64169 (I1093891,I1094406,I1094290);
not I_64170 (I1094495,I3570);
DFFARX1 I_64171 (I772294,I3563,I1094495,I1094521,);
and I_64172 (I1094529,I1094521,I772282);
DFFARX1 I_64173 (I1094529,I3563,I1094495,I1094478,);
DFFARX1 I_64174 (I772285,I3563,I1094495,I1094569,);
not I_64175 (I1094577,I772279);
not I_64176 (I1094594,I772303);
nand I_64177 (I1094611,I1094594,I1094577);
nor I_64178 (I1094466,I1094569,I1094611);
DFFARX1 I_64179 (I1094611,I3563,I1094495,I1094651,);
not I_64180 (I1094487,I1094651);
not I_64181 (I1094673,I772291);
nand I_64182 (I1094690,I1094594,I1094673);
DFFARX1 I_64183 (I1094690,I3563,I1094495,I1094716,);
not I_64184 (I1094724,I1094716);
not I_64185 (I1094741,I772300);
nand I_64186 (I1094758,I1094741,I772297);
and I_64187 (I1094775,I1094577,I1094758);
nor I_64188 (I1094792,I1094690,I1094775);
DFFARX1 I_64189 (I1094792,I3563,I1094495,I1094463,);
DFFARX1 I_64190 (I1094775,I3563,I1094495,I1094484,);
nor I_64191 (I1094837,I772300,I772288);
nor I_64192 (I1094475,I1094690,I1094837);
or I_64193 (I1094868,I772300,I772288);
nor I_64194 (I1094885,I772279,I772282);
DFFARX1 I_64195 (I1094885,I3563,I1094495,I1094911,);
not I_64196 (I1094919,I1094911);
nor I_64197 (I1094481,I1094919,I1094724);
nand I_64198 (I1094950,I1094919,I1094569);
not I_64199 (I1094967,I772279);
nand I_64200 (I1094984,I1094967,I1094673);
nand I_64201 (I1095001,I1094919,I1094984);
nand I_64202 (I1094472,I1095001,I1094950);
nand I_64203 (I1094469,I1094984,I1094868);
not I_64204 (I1095073,I3570);
DFFARX1 I_64205 (I1328655,I3563,I1095073,I1095099,);
and I_64206 (I1095107,I1095099,I1328682);
DFFARX1 I_64207 (I1095107,I3563,I1095073,I1095056,);
DFFARX1 I_64208 (I1328664,I3563,I1095073,I1095147,);
not I_64209 (I1095155,I1328673);
not I_64210 (I1095172,I1328676);
nand I_64211 (I1095189,I1095172,I1095155);
nor I_64212 (I1095044,I1095147,I1095189);
DFFARX1 I_64213 (I1095189,I3563,I1095073,I1095229,);
not I_64214 (I1095065,I1095229);
not I_64215 (I1095251,I1328670);
nand I_64216 (I1095268,I1095172,I1095251);
DFFARX1 I_64217 (I1095268,I3563,I1095073,I1095294,);
not I_64218 (I1095302,I1095294);
not I_64219 (I1095319,I1328658);
nand I_64220 (I1095336,I1095319,I1328661);
and I_64221 (I1095353,I1095155,I1095336);
nor I_64222 (I1095370,I1095268,I1095353);
DFFARX1 I_64223 (I1095370,I3563,I1095073,I1095041,);
DFFARX1 I_64224 (I1095353,I3563,I1095073,I1095062,);
nor I_64225 (I1095415,I1328658,I1328679);
nor I_64226 (I1095053,I1095268,I1095415);
or I_64227 (I1095446,I1328658,I1328679);
nor I_64228 (I1095463,I1328667,I1328655);
DFFARX1 I_64229 (I1095463,I3563,I1095073,I1095489,);
not I_64230 (I1095497,I1095489);
nor I_64231 (I1095059,I1095497,I1095302);
nand I_64232 (I1095528,I1095497,I1095147);
not I_64233 (I1095545,I1328667);
nand I_64234 (I1095562,I1095545,I1095251);
nand I_64235 (I1095579,I1095497,I1095562);
nand I_64236 (I1095050,I1095579,I1095528);
nand I_64237 (I1095047,I1095562,I1095446);
not I_64238 (I1095651,I3570);
DFFARX1 I_64239 (I45580,I3563,I1095651,I1095677,);
and I_64240 (I1095685,I1095677,I45583);
DFFARX1 I_64241 (I1095685,I3563,I1095651,I1095634,);
DFFARX1 I_64242 (I45583,I3563,I1095651,I1095725,);
not I_64243 (I1095733,I45586);
not I_64244 (I1095750,I45601);
nand I_64245 (I1095767,I1095750,I1095733);
nor I_64246 (I1095622,I1095725,I1095767);
DFFARX1 I_64247 (I1095767,I3563,I1095651,I1095807,);
not I_64248 (I1095643,I1095807);
not I_64249 (I1095829,I45595);
nand I_64250 (I1095846,I1095750,I1095829);
DFFARX1 I_64251 (I1095846,I3563,I1095651,I1095872,);
not I_64252 (I1095880,I1095872);
not I_64253 (I1095897,I45598);
nand I_64254 (I1095914,I1095897,I45580);
and I_64255 (I1095931,I1095733,I1095914);
nor I_64256 (I1095948,I1095846,I1095931);
DFFARX1 I_64257 (I1095948,I3563,I1095651,I1095619,);
DFFARX1 I_64258 (I1095931,I3563,I1095651,I1095640,);
nor I_64259 (I1095993,I45598,I45592);
nor I_64260 (I1095631,I1095846,I1095993);
or I_64261 (I1096024,I45598,I45592);
nor I_64262 (I1096041,I45589,I45604);
DFFARX1 I_64263 (I1096041,I3563,I1095651,I1096067,);
not I_64264 (I1096075,I1096067);
nor I_64265 (I1095637,I1096075,I1095880);
nand I_64266 (I1096106,I1096075,I1095725);
not I_64267 (I1096123,I45589);
nand I_64268 (I1096140,I1096123,I1095829);
nand I_64269 (I1096157,I1096075,I1096140);
nand I_64270 (I1095628,I1096157,I1096106);
nand I_64271 (I1095625,I1096140,I1096024);
not I_64272 (I1096229,I3570);
DFFARX1 I_64273 (I1324167,I3563,I1096229,I1096255,);
and I_64274 (I1096263,I1096255,I1324194);
DFFARX1 I_64275 (I1096263,I3563,I1096229,I1096212,);
DFFARX1 I_64276 (I1324176,I3563,I1096229,I1096303,);
not I_64277 (I1096311,I1324185);
not I_64278 (I1096328,I1324188);
nand I_64279 (I1096345,I1096328,I1096311);
nor I_64280 (I1096200,I1096303,I1096345);
DFFARX1 I_64281 (I1096345,I3563,I1096229,I1096385,);
not I_64282 (I1096221,I1096385);
not I_64283 (I1096407,I1324182);
nand I_64284 (I1096424,I1096328,I1096407);
DFFARX1 I_64285 (I1096424,I3563,I1096229,I1096450,);
not I_64286 (I1096458,I1096450);
not I_64287 (I1096475,I1324170);
nand I_64288 (I1096492,I1096475,I1324173);
and I_64289 (I1096509,I1096311,I1096492);
nor I_64290 (I1096526,I1096424,I1096509);
DFFARX1 I_64291 (I1096526,I3563,I1096229,I1096197,);
DFFARX1 I_64292 (I1096509,I3563,I1096229,I1096218,);
nor I_64293 (I1096571,I1324170,I1324191);
nor I_64294 (I1096209,I1096424,I1096571);
or I_64295 (I1096602,I1324170,I1324191);
nor I_64296 (I1096619,I1324179,I1324167);
DFFARX1 I_64297 (I1096619,I3563,I1096229,I1096645,);
not I_64298 (I1096653,I1096645);
nor I_64299 (I1096215,I1096653,I1096458);
nand I_64300 (I1096684,I1096653,I1096303);
not I_64301 (I1096701,I1324179);
nand I_64302 (I1096718,I1096701,I1096407);
nand I_64303 (I1096735,I1096653,I1096718);
nand I_64304 (I1096206,I1096735,I1096684);
nand I_64305 (I1096203,I1096718,I1096602);
not I_64306 (I1096807,I3570);
DFFARX1 I_64307 (I639354,I3563,I1096807,I1096833,);
and I_64308 (I1096841,I1096833,I639342);
DFFARX1 I_64309 (I1096841,I3563,I1096807,I1096790,);
DFFARX1 I_64310 (I639357,I3563,I1096807,I1096881,);
not I_64311 (I1096889,I639348);
not I_64312 (I1096906,I639339);
nand I_64313 (I1096923,I1096906,I1096889);
nor I_64314 (I1096778,I1096881,I1096923);
DFFARX1 I_64315 (I1096923,I3563,I1096807,I1096963,);
not I_64316 (I1096799,I1096963);
not I_64317 (I1096985,I639345);
nand I_64318 (I1097002,I1096906,I1096985);
DFFARX1 I_64319 (I1097002,I3563,I1096807,I1097028,);
not I_64320 (I1097036,I1097028);
not I_64321 (I1097053,I639360);
nand I_64322 (I1097070,I1097053,I639363);
and I_64323 (I1097087,I1096889,I1097070);
nor I_64324 (I1097104,I1097002,I1097087);
DFFARX1 I_64325 (I1097104,I3563,I1096807,I1096775,);
DFFARX1 I_64326 (I1097087,I3563,I1096807,I1096796,);
nor I_64327 (I1097149,I639360,I639339);
nor I_64328 (I1096787,I1097002,I1097149);
or I_64329 (I1097180,I639360,I639339);
nor I_64330 (I1097197,I639351,I639342);
DFFARX1 I_64331 (I1097197,I3563,I1096807,I1097223,);
not I_64332 (I1097231,I1097223);
nor I_64333 (I1096793,I1097231,I1097036);
nand I_64334 (I1097262,I1097231,I1096881);
not I_64335 (I1097279,I639351);
nand I_64336 (I1097296,I1097279,I1096985);
nand I_64337 (I1097313,I1097231,I1097296);
nand I_64338 (I1096784,I1097313,I1097262);
nand I_64339 (I1096781,I1097296,I1097180);
not I_64340 (I1097385,I3570);
DFFARX1 I_64341 (I1269278,I3563,I1097385,I1097411,);
and I_64342 (I1097419,I1097411,I1269272);
DFFARX1 I_64343 (I1097419,I3563,I1097385,I1097368,);
DFFARX1 I_64344 (I1269257,I3563,I1097385,I1097459,);
not I_64345 (I1097467,I1269263);
not I_64346 (I1097484,I1269275);
nand I_64347 (I1097501,I1097484,I1097467);
nor I_64348 (I1097356,I1097459,I1097501);
DFFARX1 I_64349 (I1097501,I3563,I1097385,I1097541,);
not I_64350 (I1097377,I1097541);
not I_64351 (I1097563,I1269257);
nand I_64352 (I1097580,I1097484,I1097563);
DFFARX1 I_64353 (I1097580,I3563,I1097385,I1097606,);
not I_64354 (I1097614,I1097606);
not I_64355 (I1097631,I1269281);
nand I_64356 (I1097648,I1097631,I1269269);
and I_64357 (I1097665,I1097467,I1097648);
nor I_64358 (I1097682,I1097580,I1097665);
DFFARX1 I_64359 (I1097682,I3563,I1097385,I1097353,);
DFFARX1 I_64360 (I1097665,I3563,I1097385,I1097374,);
nor I_64361 (I1097727,I1269281,I1269260);
nor I_64362 (I1097365,I1097580,I1097727);
or I_64363 (I1097758,I1269281,I1269260);
nor I_64364 (I1097775,I1269266,I1269260);
DFFARX1 I_64365 (I1097775,I3563,I1097385,I1097801,);
not I_64366 (I1097809,I1097801);
nor I_64367 (I1097371,I1097809,I1097614);
nand I_64368 (I1097840,I1097809,I1097459);
not I_64369 (I1097857,I1269266);
nand I_64370 (I1097874,I1097857,I1097563);
nand I_64371 (I1097891,I1097809,I1097874);
nand I_64372 (I1097362,I1097891,I1097840);
nand I_64373 (I1097359,I1097874,I1097758);
not I_64374 (I1097963,I3570);
DFFARX1 I_64375 (I233328,I3563,I1097963,I1097989,);
and I_64376 (I1097997,I1097989,I233331);
DFFARX1 I_64377 (I1097997,I3563,I1097963,I1097946,);
DFFARX1 I_64378 (I233331,I3563,I1097963,I1098037,);
not I_64379 (I1098045,I233346);
not I_64380 (I1098062,I233352);
nand I_64381 (I1098079,I1098062,I1098045);
nor I_64382 (I1097934,I1098037,I1098079);
DFFARX1 I_64383 (I1098079,I3563,I1097963,I1098119,);
not I_64384 (I1097955,I1098119);
not I_64385 (I1098141,I233340);
nand I_64386 (I1098158,I1098062,I1098141);
DFFARX1 I_64387 (I1098158,I3563,I1097963,I1098184,);
not I_64388 (I1098192,I1098184);
not I_64389 (I1098209,I233337);
nand I_64390 (I1098226,I1098209,I233334);
and I_64391 (I1098243,I1098045,I1098226);
nor I_64392 (I1098260,I1098158,I1098243);
DFFARX1 I_64393 (I1098260,I3563,I1097963,I1097931,);
DFFARX1 I_64394 (I1098243,I3563,I1097963,I1097952,);
nor I_64395 (I1098305,I233337,I233328);
nor I_64396 (I1097943,I1098158,I1098305);
or I_64397 (I1098336,I233337,I233328);
nor I_64398 (I1098353,I233343,I233349);
DFFARX1 I_64399 (I1098353,I3563,I1097963,I1098379,);
not I_64400 (I1098387,I1098379);
nor I_64401 (I1097949,I1098387,I1098192);
nand I_64402 (I1098418,I1098387,I1098037);
not I_64403 (I1098435,I233343);
nand I_64404 (I1098452,I1098435,I1098141);
nand I_64405 (I1098469,I1098387,I1098452);
nand I_64406 (I1097940,I1098469,I1098418);
nand I_64407 (I1097937,I1098452,I1098336);
not I_64408 (I1098541,I3570);
DFFARX1 I_64409 (I1016303,I3563,I1098541,I1098567,);
and I_64410 (I1098575,I1098567,I1016297);
DFFARX1 I_64411 (I1098575,I3563,I1098541,I1098524,);
DFFARX1 I_64412 (I1016315,I3563,I1098541,I1098615,);
not I_64413 (I1098623,I1016306);
not I_64414 (I1098640,I1016318);
nand I_64415 (I1098657,I1098640,I1098623);
nor I_64416 (I1098512,I1098615,I1098657);
DFFARX1 I_64417 (I1098657,I3563,I1098541,I1098697,);
not I_64418 (I1098533,I1098697);
not I_64419 (I1098719,I1016324);
nand I_64420 (I1098736,I1098640,I1098719);
DFFARX1 I_64421 (I1098736,I3563,I1098541,I1098762,);
not I_64422 (I1098770,I1098762);
not I_64423 (I1098787,I1016300);
nand I_64424 (I1098804,I1098787,I1016321);
and I_64425 (I1098821,I1098623,I1098804);
nor I_64426 (I1098838,I1098736,I1098821);
DFFARX1 I_64427 (I1098838,I3563,I1098541,I1098509,);
DFFARX1 I_64428 (I1098821,I3563,I1098541,I1098530,);
nor I_64429 (I1098883,I1016300,I1016312);
nor I_64430 (I1098521,I1098736,I1098883);
or I_64431 (I1098914,I1016300,I1016312);
nor I_64432 (I1098931,I1016297,I1016309);
DFFARX1 I_64433 (I1098931,I3563,I1098541,I1098957,);
not I_64434 (I1098965,I1098957);
nor I_64435 (I1098527,I1098965,I1098770);
nand I_64436 (I1098996,I1098965,I1098615);
not I_64437 (I1099013,I1016297);
nand I_64438 (I1099030,I1099013,I1098719);
nand I_64439 (I1099047,I1098965,I1099030);
nand I_64440 (I1098518,I1099047,I1098996);
nand I_64441 (I1098515,I1099030,I1098914);
not I_64442 (I1099119,I3570);
DFFARX1 I_64443 (I763624,I3563,I1099119,I1099145,);
and I_64444 (I1099153,I1099145,I763612);
DFFARX1 I_64445 (I1099153,I3563,I1099119,I1099102,);
DFFARX1 I_64446 (I763615,I3563,I1099119,I1099193,);
not I_64447 (I1099201,I763609);
not I_64448 (I1099218,I763633);
nand I_64449 (I1099235,I1099218,I1099201);
nor I_64450 (I1099090,I1099193,I1099235);
DFFARX1 I_64451 (I1099235,I3563,I1099119,I1099275,);
not I_64452 (I1099111,I1099275);
not I_64453 (I1099297,I763621);
nand I_64454 (I1099314,I1099218,I1099297);
DFFARX1 I_64455 (I1099314,I3563,I1099119,I1099340,);
not I_64456 (I1099348,I1099340);
not I_64457 (I1099365,I763630);
nand I_64458 (I1099382,I1099365,I763627);
and I_64459 (I1099399,I1099201,I1099382);
nor I_64460 (I1099416,I1099314,I1099399);
DFFARX1 I_64461 (I1099416,I3563,I1099119,I1099087,);
DFFARX1 I_64462 (I1099399,I3563,I1099119,I1099108,);
nor I_64463 (I1099461,I763630,I763618);
nor I_64464 (I1099099,I1099314,I1099461);
or I_64465 (I1099492,I763630,I763618);
nor I_64466 (I1099509,I763609,I763612);
DFFARX1 I_64467 (I1099509,I3563,I1099119,I1099535,);
not I_64468 (I1099543,I1099535);
nor I_64469 (I1099105,I1099543,I1099348);
nand I_64470 (I1099574,I1099543,I1099193);
not I_64471 (I1099591,I763609);
nand I_64472 (I1099608,I1099591,I1099297);
nand I_64473 (I1099625,I1099543,I1099608);
nand I_64474 (I1099096,I1099625,I1099574);
nand I_64475 (I1099093,I1099608,I1099492);
not I_64476 (I1099697,I3570);
DFFARX1 I_64477 (I260698,I3563,I1099697,I1099723,);
and I_64478 (I1099731,I1099723,I260701);
DFFARX1 I_64479 (I1099731,I3563,I1099697,I1099680,);
DFFARX1 I_64480 (I260701,I3563,I1099697,I1099771,);
not I_64481 (I1099779,I260716);
not I_64482 (I1099796,I260722);
nand I_64483 (I1099813,I1099796,I1099779);
nor I_64484 (I1099668,I1099771,I1099813);
DFFARX1 I_64485 (I1099813,I3563,I1099697,I1099853,);
not I_64486 (I1099689,I1099853);
not I_64487 (I1099875,I260710);
nand I_64488 (I1099892,I1099796,I1099875);
DFFARX1 I_64489 (I1099892,I3563,I1099697,I1099918,);
not I_64490 (I1099926,I1099918);
not I_64491 (I1099943,I260707);
nand I_64492 (I1099960,I1099943,I260704);
and I_64493 (I1099977,I1099779,I1099960);
nor I_64494 (I1099994,I1099892,I1099977);
DFFARX1 I_64495 (I1099994,I3563,I1099697,I1099665,);
DFFARX1 I_64496 (I1099977,I3563,I1099697,I1099686,);
nor I_64497 (I1100039,I260707,I260698);
nor I_64498 (I1099677,I1099892,I1100039);
or I_64499 (I1100070,I260707,I260698);
nor I_64500 (I1100087,I260713,I260719);
DFFARX1 I_64501 (I1100087,I3563,I1099697,I1100113,);
not I_64502 (I1100121,I1100113);
nor I_64503 (I1099683,I1100121,I1099926);
nand I_64504 (I1100152,I1100121,I1099771);
not I_64505 (I1100169,I260713);
nand I_64506 (I1100186,I1100169,I1099875);
nand I_64507 (I1100203,I1100121,I1100186);
nand I_64508 (I1099674,I1100203,I1100152);
nand I_64509 (I1099671,I1100186,I1100070);
not I_64510 (I1100275,I3570);
DFFARX1 I_64511 (I288554,I3563,I1100275,I1100301,);
and I_64512 (I1100309,I1100301,I288539);
DFFARX1 I_64513 (I1100309,I3563,I1100275,I1100258,);
DFFARX1 I_64514 (I288545,I3563,I1100275,I1100349,);
not I_64515 (I1100357,I288527);
not I_64516 (I1100374,I288548);
nand I_64517 (I1100391,I1100374,I1100357);
nor I_64518 (I1100246,I1100349,I1100391);
DFFARX1 I_64519 (I1100391,I3563,I1100275,I1100431,);
not I_64520 (I1100267,I1100431);
not I_64521 (I1100453,I288551);
nand I_64522 (I1100470,I1100374,I1100453);
DFFARX1 I_64523 (I1100470,I3563,I1100275,I1100496,);
not I_64524 (I1100504,I1100496);
not I_64525 (I1100521,I288542);
nand I_64526 (I1100538,I1100521,I288530);
and I_64527 (I1100555,I1100357,I1100538);
nor I_64528 (I1100572,I1100470,I1100555);
DFFARX1 I_64529 (I1100572,I3563,I1100275,I1100243,);
DFFARX1 I_64530 (I1100555,I3563,I1100275,I1100264,);
nor I_64531 (I1100617,I288542,I288536);
nor I_64532 (I1100255,I1100470,I1100617);
or I_64533 (I1100648,I288542,I288536);
nor I_64534 (I1100665,I288533,I288527);
DFFARX1 I_64535 (I1100665,I3563,I1100275,I1100691,);
not I_64536 (I1100699,I1100691);
nor I_64537 (I1100261,I1100699,I1100504);
nand I_64538 (I1100730,I1100699,I1100349);
not I_64539 (I1100747,I288533);
nand I_64540 (I1100764,I1100747,I1100453);
nand I_64541 (I1100781,I1100699,I1100764);
nand I_64542 (I1100252,I1100781,I1100730);
nand I_64543 (I1100249,I1100764,I1100648);
not I_64544 (I1100853,I3570);
DFFARX1 I_64545 (I74589,I3563,I1100853,I1100879,);
and I_64546 (I1100887,I1100879,I74565);
DFFARX1 I_64547 (I1100887,I3563,I1100853,I1100836,);
DFFARX1 I_64548 (I74583,I3563,I1100853,I1100927,);
not I_64549 (I1100935,I74571);
not I_64550 (I1100952,I74568);
nand I_64551 (I1100969,I1100952,I1100935);
nor I_64552 (I1100824,I1100927,I1100969);
DFFARX1 I_64553 (I1100969,I3563,I1100853,I1101009,);
not I_64554 (I1100845,I1101009);
not I_64555 (I1101031,I74577);
nand I_64556 (I1101048,I1100952,I1101031);
DFFARX1 I_64557 (I1101048,I3563,I1100853,I1101074,);
not I_64558 (I1101082,I1101074);
not I_64559 (I1101099,I74568);
nand I_64560 (I1101116,I1101099,I74586);
and I_64561 (I1101133,I1100935,I1101116);
nor I_64562 (I1101150,I1101048,I1101133);
DFFARX1 I_64563 (I1101150,I3563,I1100853,I1100821,);
DFFARX1 I_64564 (I1101133,I3563,I1100853,I1100842,);
nor I_64565 (I1101195,I74568,I74580);
nor I_64566 (I1100833,I1101048,I1101195);
or I_64567 (I1101226,I74568,I74580);
nor I_64568 (I1101243,I74574,I74565);
DFFARX1 I_64569 (I1101243,I3563,I1100853,I1101269,);
not I_64570 (I1101277,I1101269);
nor I_64571 (I1100839,I1101277,I1101082);
nand I_64572 (I1101308,I1101277,I1100927);
not I_64573 (I1101325,I74574);
nand I_64574 (I1101342,I1101325,I1101031);
nand I_64575 (I1101359,I1101277,I1101342);
nand I_64576 (I1100830,I1101359,I1101308);
nand I_64577 (I1100827,I1101342,I1101226);
not I_64578 (I1101431,I3570);
DFFARX1 I_64579 (I347578,I3563,I1101431,I1101457,);
and I_64580 (I1101465,I1101457,I347563);
DFFARX1 I_64581 (I1101465,I3563,I1101431,I1101414,);
DFFARX1 I_64582 (I347569,I3563,I1101431,I1101505,);
not I_64583 (I1101513,I347551);
not I_64584 (I1101530,I347572);
nand I_64585 (I1101547,I1101530,I1101513);
nor I_64586 (I1101402,I1101505,I1101547);
DFFARX1 I_64587 (I1101547,I3563,I1101431,I1101587,);
not I_64588 (I1101423,I1101587);
not I_64589 (I1101609,I347575);
nand I_64590 (I1101626,I1101530,I1101609);
DFFARX1 I_64591 (I1101626,I3563,I1101431,I1101652,);
not I_64592 (I1101660,I1101652);
not I_64593 (I1101677,I347566);
nand I_64594 (I1101694,I1101677,I347554);
and I_64595 (I1101711,I1101513,I1101694);
nor I_64596 (I1101728,I1101626,I1101711);
DFFARX1 I_64597 (I1101728,I3563,I1101431,I1101399,);
DFFARX1 I_64598 (I1101711,I3563,I1101431,I1101420,);
nor I_64599 (I1101773,I347566,I347560);
nor I_64600 (I1101411,I1101626,I1101773);
or I_64601 (I1101804,I347566,I347560);
nor I_64602 (I1101821,I347557,I347551);
DFFARX1 I_64603 (I1101821,I3563,I1101431,I1101847,);
not I_64604 (I1101855,I1101847);
nor I_64605 (I1101417,I1101855,I1101660);
nand I_64606 (I1101886,I1101855,I1101505);
not I_64607 (I1101903,I347557);
nand I_64608 (I1101920,I1101903,I1101609);
nand I_64609 (I1101937,I1101855,I1101920);
nand I_64610 (I1101408,I1101937,I1101886);
nand I_64611 (I1101405,I1101920,I1101804);
not I_64612 (I1102009,I3570);
DFFARX1 I_64613 (I528689,I3563,I1102009,I1102035,);
and I_64614 (I1102043,I1102035,I528704);
DFFARX1 I_64615 (I1102043,I3563,I1102009,I1101992,);
DFFARX1 I_64616 (I528695,I3563,I1102009,I1102083,);
not I_64617 (I1102091,I528689);
not I_64618 (I1102108,I528707);
nand I_64619 (I1102125,I1102108,I1102091);
nor I_64620 (I1101980,I1102083,I1102125);
DFFARX1 I_64621 (I1102125,I3563,I1102009,I1102165,);
not I_64622 (I1102001,I1102165);
not I_64623 (I1102187,I528698);
nand I_64624 (I1102204,I1102108,I1102187);
DFFARX1 I_64625 (I1102204,I3563,I1102009,I1102230,);
not I_64626 (I1102238,I1102230);
not I_64627 (I1102255,I528710);
nand I_64628 (I1102272,I1102255,I528686);
and I_64629 (I1102289,I1102091,I1102272);
nor I_64630 (I1102306,I1102204,I1102289);
DFFARX1 I_64631 (I1102306,I3563,I1102009,I1101977,);
DFFARX1 I_64632 (I1102289,I3563,I1102009,I1101998,);
nor I_64633 (I1102351,I528710,I528686);
nor I_64634 (I1101989,I1102204,I1102351);
or I_64635 (I1102382,I528710,I528686);
nor I_64636 (I1102399,I528692,I528701);
DFFARX1 I_64637 (I1102399,I3563,I1102009,I1102425,);
not I_64638 (I1102433,I1102425);
nor I_64639 (I1101995,I1102433,I1102238);
nand I_64640 (I1102464,I1102433,I1102083);
not I_64641 (I1102481,I528692);
nand I_64642 (I1102498,I1102481,I1102187);
nand I_64643 (I1102515,I1102433,I1102498);
nand I_64644 (I1101986,I1102515,I1102464);
nand I_64645 (I1101983,I1102498,I1102382);
not I_64646 (I1102587,I3570);
DFFARX1 I_64647 (I815275,I3563,I1102587,I1102613,);
and I_64648 (I1102621,I1102613,I815281);
DFFARX1 I_64649 (I1102621,I3563,I1102587,I1102570,);
DFFARX1 I_64650 (I815287,I3563,I1102587,I1102661,);
not I_64651 (I1102669,I815272);
not I_64652 (I1102686,I815272);
nand I_64653 (I1102703,I1102686,I1102669);
nor I_64654 (I1102558,I1102661,I1102703);
DFFARX1 I_64655 (I1102703,I3563,I1102587,I1102743,);
not I_64656 (I1102579,I1102743);
not I_64657 (I1102765,I815290);
nand I_64658 (I1102782,I1102686,I1102765);
DFFARX1 I_64659 (I1102782,I3563,I1102587,I1102808,);
not I_64660 (I1102816,I1102808);
not I_64661 (I1102833,I815284);
nand I_64662 (I1102850,I1102833,I815275);
and I_64663 (I1102867,I1102669,I1102850);
nor I_64664 (I1102884,I1102782,I1102867);
DFFARX1 I_64665 (I1102884,I3563,I1102587,I1102555,);
DFFARX1 I_64666 (I1102867,I3563,I1102587,I1102576,);
nor I_64667 (I1102929,I815284,I815293);
nor I_64668 (I1102567,I1102782,I1102929);
or I_64669 (I1102960,I815284,I815293);
nor I_64670 (I1102977,I815278,I815278);
DFFARX1 I_64671 (I1102977,I3563,I1102587,I1103003,);
not I_64672 (I1103011,I1103003);
nor I_64673 (I1102573,I1103011,I1102816);
nand I_64674 (I1103042,I1103011,I1102661);
not I_64675 (I1103059,I815278);
nand I_64676 (I1103076,I1103059,I1102765);
nand I_64677 (I1103093,I1103011,I1103076);
nand I_64678 (I1102564,I1103093,I1103042);
nand I_64679 (I1102561,I1103076,I1102960);
not I_64680 (I1103165,I3570);
DFFARX1 I_64681 (I606408,I3563,I1103165,I1103191,);
and I_64682 (I1103199,I1103191,I606396);
DFFARX1 I_64683 (I1103199,I3563,I1103165,I1103148,);
DFFARX1 I_64684 (I606411,I3563,I1103165,I1103239,);
not I_64685 (I1103247,I606402);
not I_64686 (I1103264,I606393);
nand I_64687 (I1103281,I1103264,I1103247);
nor I_64688 (I1103136,I1103239,I1103281);
DFFARX1 I_64689 (I1103281,I3563,I1103165,I1103321,);
not I_64690 (I1103157,I1103321);
not I_64691 (I1103343,I606399);
nand I_64692 (I1103360,I1103264,I1103343);
DFFARX1 I_64693 (I1103360,I3563,I1103165,I1103386,);
not I_64694 (I1103394,I1103386);
not I_64695 (I1103411,I606414);
nand I_64696 (I1103428,I1103411,I606417);
and I_64697 (I1103445,I1103247,I1103428);
nor I_64698 (I1103462,I1103360,I1103445);
DFFARX1 I_64699 (I1103462,I3563,I1103165,I1103133,);
DFFARX1 I_64700 (I1103445,I3563,I1103165,I1103154,);
nor I_64701 (I1103507,I606414,I606393);
nor I_64702 (I1103145,I1103360,I1103507);
or I_64703 (I1103538,I606414,I606393);
nor I_64704 (I1103555,I606405,I606396);
DFFARX1 I_64705 (I1103555,I3563,I1103165,I1103581,);
not I_64706 (I1103589,I1103581);
nor I_64707 (I1103151,I1103589,I1103394);
nand I_64708 (I1103620,I1103589,I1103239);
not I_64709 (I1103637,I606405);
nand I_64710 (I1103654,I1103637,I1103343);
nand I_64711 (I1103671,I1103589,I1103654);
nand I_64712 (I1103142,I1103671,I1103620);
nand I_64713 (I1103139,I1103654,I1103538);
not I_64714 (I1103743,I3570);
DFFARX1 I_64715 (I579242,I3563,I1103743,I1103769,);
and I_64716 (I1103777,I1103769,I579230);
DFFARX1 I_64717 (I1103777,I3563,I1103743,I1103726,);
DFFARX1 I_64718 (I579245,I3563,I1103743,I1103817,);
not I_64719 (I1103825,I579236);
not I_64720 (I1103842,I579227);
nand I_64721 (I1103859,I1103842,I1103825);
nor I_64722 (I1103714,I1103817,I1103859);
DFFARX1 I_64723 (I1103859,I3563,I1103743,I1103899,);
not I_64724 (I1103735,I1103899);
not I_64725 (I1103921,I579233);
nand I_64726 (I1103938,I1103842,I1103921);
DFFARX1 I_64727 (I1103938,I3563,I1103743,I1103964,);
not I_64728 (I1103972,I1103964);
not I_64729 (I1103989,I579248);
nand I_64730 (I1104006,I1103989,I579251);
and I_64731 (I1104023,I1103825,I1104006);
nor I_64732 (I1104040,I1103938,I1104023);
DFFARX1 I_64733 (I1104040,I3563,I1103743,I1103711,);
DFFARX1 I_64734 (I1104023,I3563,I1103743,I1103732,);
nor I_64735 (I1104085,I579248,I579227);
nor I_64736 (I1103723,I1103938,I1104085);
or I_64737 (I1104116,I579248,I579227);
nor I_64738 (I1104133,I579239,I579230);
DFFARX1 I_64739 (I1104133,I3563,I1103743,I1104159,);
not I_64740 (I1104167,I1104159);
nor I_64741 (I1103729,I1104167,I1103972);
nand I_64742 (I1104198,I1104167,I1103817);
not I_64743 (I1104215,I579239);
nand I_64744 (I1104232,I1104215,I1103921);
nand I_64745 (I1104249,I1104167,I1104232);
nand I_64746 (I1103720,I1104249,I1104198);
nand I_64747 (I1103717,I1104232,I1104116);
not I_64748 (I1104321,I3570);
DFFARX1 I_64749 (I682704,I3563,I1104321,I1104347,);
and I_64750 (I1104355,I1104347,I682692);
DFFARX1 I_64751 (I1104355,I3563,I1104321,I1104304,);
DFFARX1 I_64752 (I682695,I3563,I1104321,I1104395,);
not I_64753 (I1104403,I682689);
not I_64754 (I1104420,I682713);
nand I_64755 (I1104437,I1104420,I1104403);
nor I_64756 (I1104292,I1104395,I1104437);
DFFARX1 I_64757 (I1104437,I3563,I1104321,I1104477,);
not I_64758 (I1104313,I1104477);
not I_64759 (I1104499,I682701);
nand I_64760 (I1104516,I1104420,I1104499);
DFFARX1 I_64761 (I1104516,I3563,I1104321,I1104542,);
not I_64762 (I1104550,I1104542);
not I_64763 (I1104567,I682710);
nand I_64764 (I1104584,I1104567,I682707);
and I_64765 (I1104601,I1104403,I1104584);
nor I_64766 (I1104618,I1104516,I1104601);
DFFARX1 I_64767 (I1104618,I3563,I1104321,I1104289,);
DFFARX1 I_64768 (I1104601,I3563,I1104321,I1104310,);
nor I_64769 (I1104663,I682710,I682698);
nor I_64770 (I1104301,I1104516,I1104663);
or I_64771 (I1104694,I682710,I682698);
nor I_64772 (I1104711,I682689,I682692);
DFFARX1 I_64773 (I1104711,I3563,I1104321,I1104737,);
not I_64774 (I1104745,I1104737);
nor I_64775 (I1104307,I1104745,I1104550);
nand I_64776 (I1104776,I1104745,I1104395);
not I_64777 (I1104793,I682689);
nand I_64778 (I1104810,I1104793,I1104499);
nand I_64779 (I1104827,I1104745,I1104810);
nand I_64780 (I1104298,I1104827,I1104776);
nand I_64781 (I1104295,I1104810,I1104694);
not I_64782 (I1104899,I3570);
DFFARX1 I_64783 (I1030515,I3563,I1104899,I1104925,);
and I_64784 (I1104933,I1104925,I1030509);
DFFARX1 I_64785 (I1104933,I3563,I1104899,I1104882,);
DFFARX1 I_64786 (I1030527,I3563,I1104899,I1104973,);
not I_64787 (I1104981,I1030518);
not I_64788 (I1104998,I1030530);
nand I_64789 (I1105015,I1104998,I1104981);
nor I_64790 (I1104870,I1104973,I1105015);
DFFARX1 I_64791 (I1105015,I3563,I1104899,I1105055,);
not I_64792 (I1104891,I1105055);
not I_64793 (I1105077,I1030536);
nand I_64794 (I1105094,I1104998,I1105077);
DFFARX1 I_64795 (I1105094,I3563,I1104899,I1105120,);
not I_64796 (I1105128,I1105120);
not I_64797 (I1105145,I1030512);
nand I_64798 (I1105162,I1105145,I1030533);
and I_64799 (I1105179,I1104981,I1105162);
nor I_64800 (I1105196,I1105094,I1105179);
DFFARX1 I_64801 (I1105196,I3563,I1104899,I1104867,);
DFFARX1 I_64802 (I1105179,I3563,I1104899,I1104888,);
nor I_64803 (I1105241,I1030512,I1030524);
nor I_64804 (I1104879,I1105094,I1105241);
or I_64805 (I1105272,I1030512,I1030524);
nor I_64806 (I1105289,I1030509,I1030521);
DFFARX1 I_64807 (I1105289,I3563,I1104899,I1105315,);
not I_64808 (I1105323,I1105315);
nor I_64809 (I1104885,I1105323,I1105128);
nand I_64810 (I1105354,I1105323,I1104973);
not I_64811 (I1105371,I1030509);
nand I_64812 (I1105388,I1105371,I1105077);
nand I_64813 (I1105405,I1105323,I1105388);
nand I_64814 (I1104876,I1105405,I1105354);
nand I_64815 (I1104873,I1105388,I1105272);
not I_64816 (I1105477,I3570);
DFFARX1 I_64817 (I222618,I3563,I1105477,I1105503,);
and I_64818 (I1105511,I1105503,I222621);
DFFARX1 I_64819 (I1105511,I3563,I1105477,I1105460,);
DFFARX1 I_64820 (I222621,I3563,I1105477,I1105551,);
not I_64821 (I1105559,I222636);
not I_64822 (I1105576,I222642);
nand I_64823 (I1105593,I1105576,I1105559);
nor I_64824 (I1105448,I1105551,I1105593);
DFFARX1 I_64825 (I1105593,I3563,I1105477,I1105633,);
not I_64826 (I1105469,I1105633);
not I_64827 (I1105655,I222630);
nand I_64828 (I1105672,I1105576,I1105655);
DFFARX1 I_64829 (I1105672,I3563,I1105477,I1105698,);
not I_64830 (I1105706,I1105698);
not I_64831 (I1105723,I222627);
nand I_64832 (I1105740,I1105723,I222624);
and I_64833 (I1105757,I1105559,I1105740);
nor I_64834 (I1105774,I1105672,I1105757);
DFFARX1 I_64835 (I1105774,I3563,I1105477,I1105445,);
DFFARX1 I_64836 (I1105757,I3563,I1105477,I1105466,);
nor I_64837 (I1105819,I222627,I222618);
nor I_64838 (I1105457,I1105672,I1105819);
or I_64839 (I1105850,I222627,I222618);
nor I_64840 (I1105867,I222633,I222639);
DFFARX1 I_64841 (I1105867,I3563,I1105477,I1105893,);
not I_64842 (I1105901,I1105893);
nor I_64843 (I1105463,I1105901,I1105706);
nand I_64844 (I1105932,I1105901,I1105551);
not I_64845 (I1105949,I222633);
nand I_64846 (I1105966,I1105949,I1105655);
nand I_64847 (I1105983,I1105901,I1105966);
nand I_64848 (I1105454,I1105983,I1105932);
nand I_64849 (I1105451,I1105966,I1105850);
not I_64850 (I1106055,I3570);
DFFARX1 I_64851 (I1335125,I3563,I1106055,I1106081,);
and I_64852 (I1106089,I1106081,I1335107);
DFFARX1 I_64853 (I1106089,I3563,I1106055,I1106038,);
DFFARX1 I_64854 (I1335098,I3563,I1106055,I1106129,);
not I_64855 (I1106137,I1335113);
not I_64856 (I1106154,I1335101);
nand I_64857 (I1106171,I1106154,I1106137);
nor I_64858 (I1106026,I1106129,I1106171);
DFFARX1 I_64859 (I1106171,I3563,I1106055,I1106211,);
not I_64860 (I1106047,I1106211);
not I_64861 (I1106233,I1335110);
nand I_64862 (I1106250,I1106154,I1106233);
DFFARX1 I_64863 (I1106250,I3563,I1106055,I1106276,);
not I_64864 (I1106284,I1106276);
not I_64865 (I1106301,I1335119);
nand I_64866 (I1106318,I1106301,I1335098);
and I_64867 (I1106335,I1106137,I1106318);
nor I_64868 (I1106352,I1106250,I1106335);
DFFARX1 I_64869 (I1106352,I3563,I1106055,I1106023,);
DFFARX1 I_64870 (I1106335,I3563,I1106055,I1106044,);
nor I_64871 (I1106397,I1335119,I1335122);
nor I_64872 (I1106035,I1106250,I1106397);
or I_64873 (I1106428,I1335119,I1335122);
nor I_64874 (I1106445,I1335116,I1335104);
DFFARX1 I_64875 (I1106445,I3563,I1106055,I1106471,);
not I_64876 (I1106479,I1106471);
nor I_64877 (I1106041,I1106479,I1106284);
nand I_64878 (I1106510,I1106479,I1106129);
not I_64879 (I1106527,I1335116);
nand I_64880 (I1106544,I1106527,I1106233);
nand I_64881 (I1106561,I1106479,I1106544);
nand I_64882 (I1106032,I1106561,I1106510);
nand I_64883 (I1106029,I1106544,I1106428);
not I_64884 (I1106633,I3570);
DFFARX1 I_64885 (I481154,I3563,I1106633,I1106659,);
and I_64886 (I1106667,I1106659,I481169);
DFFARX1 I_64887 (I1106667,I3563,I1106633,I1106616,);
DFFARX1 I_64888 (I481172,I3563,I1106633,I1106707,);
not I_64889 (I1106715,I481166);
not I_64890 (I1106732,I481181);
nand I_64891 (I1106749,I1106732,I1106715);
nor I_64892 (I1106604,I1106707,I1106749);
DFFARX1 I_64893 (I1106749,I3563,I1106633,I1106789,);
not I_64894 (I1106625,I1106789);
not I_64895 (I1106811,I481157);
nand I_64896 (I1106828,I1106732,I1106811);
DFFARX1 I_64897 (I1106828,I3563,I1106633,I1106854,);
not I_64898 (I1106862,I1106854);
not I_64899 (I1106879,I481160);
nand I_64900 (I1106896,I1106879,I481154);
and I_64901 (I1106913,I1106715,I1106896);
nor I_64902 (I1106930,I1106828,I1106913);
DFFARX1 I_64903 (I1106930,I3563,I1106633,I1106601,);
DFFARX1 I_64904 (I1106913,I3563,I1106633,I1106622,);
nor I_64905 (I1106975,I481160,I481163);
nor I_64906 (I1106613,I1106828,I1106975);
or I_64907 (I1107006,I481160,I481163);
nor I_64908 (I1107023,I481178,I481175);
DFFARX1 I_64909 (I1107023,I3563,I1106633,I1107049,);
not I_64910 (I1107057,I1107049);
nor I_64911 (I1106619,I1107057,I1106862);
nand I_64912 (I1107088,I1107057,I1106707);
not I_64913 (I1107105,I481178);
nand I_64914 (I1107122,I1107105,I1106811);
nand I_64915 (I1107139,I1107057,I1107122);
nand I_64916 (I1106610,I1107139,I1107088);
nand I_64917 (I1106607,I1107122,I1107006);
not I_64918 (I1107211,I3570);
DFFARX1 I_64919 (I89345,I3563,I1107211,I1107237,);
and I_64920 (I1107245,I1107237,I89321);
DFFARX1 I_64921 (I1107245,I3563,I1107211,I1107194,);
DFFARX1 I_64922 (I89339,I3563,I1107211,I1107285,);
not I_64923 (I1107293,I89327);
not I_64924 (I1107310,I89324);
nand I_64925 (I1107327,I1107310,I1107293);
nor I_64926 (I1107182,I1107285,I1107327);
DFFARX1 I_64927 (I1107327,I3563,I1107211,I1107367,);
not I_64928 (I1107203,I1107367);
not I_64929 (I1107389,I89333);
nand I_64930 (I1107406,I1107310,I1107389);
DFFARX1 I_64931 (I1107406,I3563,I1107211,I1107432,);
not I_64932 (I1107440,I1107432);
not I_64933 (I1107457,I89324);
nand I_64934 (I1107474,I1107457,I89342);
and I_64935 (I1107491,I1107293,I1107474);
nor I_64936 (I1107508,I1107406,I1107491);
DFFARX1 I_64937 (I1107508,I3563,I1107211,I1107179,);
DFFARX1 I_64938 (I1107491,I3563,I1107211,I1107200,);
nor I_64939 (I1107553,I89324,I89336);
nor I_64940 (I1107191,I1107406,I1107553);
or I_64941 (I1107584,I89324,I89336);
nor I_64942 (I1107601,I89330,I89321);
DFFARX1 I_64943 (I1107601,I3563,I1107211,I1107627,);
not I_64944 (I1107635,I1107627);
nor I_64945 (I1107197,I1107635,I1107440);
nand I_64946 (I1107666,I1107635,I1107285);
not I_64947 (I1107683,I89330);
nand I_64948 (I1107700,I1107683,I1107389);
nand I_64949 (I1107717,I1107635,I1107700);
nand I_64950 (I1107188,I1107717,I1107666);
nand I_64951 (I1107185,I1107700,I1107584);
not I_64952 (I1107789,I3570);
DFFARX1 I_64953 (I1393435,I3563,I1107789,I1107815,);
and I_64954 (I1107823,I1107815,I1393417);
DFFARX1 I_64955 (I1107823,I3563,I1107789,I1107772,);
DFFARX1 I_64956 (I1393408,I3563,I1107789,I1107863,);
not I_64957 (I1107871,I1393423);
not I_64958 (I1107888,I1393411);
nand I_64959 (I1107905,I1107888,I1107871);
nor I_64960 (I1107760,I1107863,I1107905);
DFFARX1 I_64961 (I1107905,I3563,I1107789,I1107945,);
not I_64962 (I1107781,I1107945);
not I_64963 (I1107967,I1393420);
nand I_64964 (I1107984,I1107888,I1107967);
DFFARX1 I_64965 (I1107984,I3563,I1107789,I1108010,);
not I_64966 (I1108018,I1108010);
not I_64967 (I1108035,I1393429);
nand I_64968 (I1108052,I1108035,I1393408);
and I_64969 (I1108069,I1107871,I1108052);
nor I_64970 (I1108086,I1107984,I1108069);
DFFARX1 I_64971 (I1108086,I3563,I1107789,I1107757,);
DFFARX1 I_64972 (I1108069,I3563,I1107789,I1107778,);
nor I_64973 (I1108131,I1393429,I1393432);
nor I_64974 (I1107769,I1107984,I1108131);
or I_64975 (I1108162,I1393429,I1393432);
nor I_64976 (I1108179,I1393426,I1393414);
DFFARX1 I_64977 (I1108179,I3563,I1107789,I1108205,);
not I_64978 (I1108213,I1108205);
nor I_64979 (I1107775,I1108213,I1108018);
nand I_64980 (I1108244,I1108213,I1107863);
not I_64981 (I1108261,I1393426);
nand I_64982 (I1108278,I1108261,I1107967);
nand I_64983 (I1108295,I1108213,I1108278);
nand I_64984 (I1107766,I1108295,I1108244);
nand I_64985 (I1107763,I1108278,I1108162);
not I_64986 (I1108367,I3570);
DFFARX1 I_64987 (I397643,I3563,I1108367,I1108393,);
and I_64988 (I1108401,I1108393,I397628);
DFFARX1 I_64989 (I1108401,I3563,I1108367,I1108350,);
DFFARX1 I_64990 (I397634,I3563,I1108367,I1108441,);
not I_64991 (I1108449,I397616);
not I_64992 (I1108466,I397637);
nand I_64993 (I1108483,I1108466,I1108449);
nor I_64994 (I1108338,I1108441,I1108483);
DFFARX1 I_64995 (I1108483,I3563,I1108367,I1108523,);
not I_64996 (I1108359,I1108523);
not I_64997 (I1108545,I397640);
nand I_64998 (I1108562,I1108466,I1108545);
DFFARX1 I_64999 (I1108562,I3563,I1108367,I1108588,);
not I_65000 (I1108596,I1108588);
not I_65001 (I1108613,I397631);
nand I_65002 (I1108630,I1108613,I397619);
and I_65003 (I1108647,I1108449,I1108630);
nor I_65004 (I1108664,I1108562,I1108647);
DFFARX1 I_65005 (I1108664,I3563,I1108367,I1108335,);
DFFARX1 I_65006 (I1108647,I3563,I1108367,I1108356,);
nor I_65007 (I1108709,I397631,I397625);
nor I_65008 (I1108347,I1108562,I1108709);
or I_65009 (I1108740,I397631,I397625);
nor I_65010 (I1108757,I397622,I397616);
DFFARX1 I_65011 (I1108757,I3563,I1108367,I1108783,);
not I_65012 (I1108791,I1108783);
nor I_65013 (I1108353,I1108791,I1108596);
nand I_65014 (I1108822,I1108791,I1108441);
not I_65015 (I1108839,I397622);
nand I_65016 (I1108856,I1108839,I1108545);
nand I_65017 (I1108873,I1108791,I1108856);
nand I_65018 (I1108344,I1108873,I1108822);
nand I_65019 (I1108341,I1108856,I1108740);
not I_65020 (I1108945,I3570);
DFFARX1 I_65021 (I160738,I3563,I1108945,I1108971,);
and I_65022 (I1108979,I1108971,I160762);
DFFARX1 I_65023 (I1108979,I3563,I1108945,I1108928,);
DFFARX1 I_65024 (I160738,I3563,I1108945,I1109019,);
not I_65025 (I1109027,I160756);
not I_65026 (I1109044,I160741);
nand I_65027 (I1109061,I1109044,I1109027);
nor I_65028 (I1108916,I1109019,I1109061);
DFFARX1 I_65029 (I1109061,I3563,I1108945,I1109101,);
not I_65030 (I1108937,I1109101);
not I_65031 (I1109123,I160750);
nand I_65032 (I1109140,I1109044,I1109123);
DFFARX1 I_65033 (I1109140,I3563,I1108945,I1109166,);
not I_65034 (I1109174,I1109166);
not I_65035 (I1109191,I160747);
nand I_65036 (I1109208,I1109191,I160744);
and I_65037 (I1109225,I1109027,I1109208);
nor I_65038 (I1109242,I1109140,I1109225);
DFFARX1 I_65039 (I1109242,I3563,I1108945,I1108913,);
DFFARX1 I_65040 (I1109225,I3563,I1108945,I1108934,);
nor I_65041 (I1109287,I160747,I160753);
nor I_65042 (I1108925,I1109140,I1109287);
or I_65043 (I1109318,I160747,I160753);
nor I_65044 (I1109335,I160759,I160765);
DFFARX1 I_65045 (I1109335,I3563,I1108945,I1109361,);
not I_65046 (I1109369,I1109361);
nor I_65047 (I1108931,I1109369,I1109174);
nand I_65048 (I1109400,I1109369,I1109019);
not I_65049 (I1109417,I160759);
nand I_65050 (I1109434,I1109417,I1109123);
nand I_65051 (I1109451,I1109369,I1109434);
nand I_65052 (I1108922,I1109451,I1109400);
nand I_65053 (I1108919,I1109434,I1109318);
not I_65054 (I1109523,I3570);
DFFARX1 I_65055 (I996923,I3563,I1109523,I1109549,);
and I_65056 (I1109557,I1109549,I996917);
DFFARX1 I_65057 (I1109557,I3563,I1109523,I1109506,);
DFFARX1 I_65058 (I996935,I3563,I1109523,I1109597,);
not I_65059 (I1109605,I996926);
not I_65060 (I1109622,I996938);
nand I_65061 (I1109639,I1109622,I1109605);
nor I_65062 (I1109494,I1109597,I1109639);
DFFARX1 I_65063 (I1109639,I3563,I1109523,I1109679,);
not I_65064 (I1109515,I1109679);
not I_65065 (I1109701,I996944);
nand I_65066 (I1109718,I1109622,I1109701);
DFFARX1 I_65067 (I1109718,I3563,I1109523,I1109744,);
not I_65068 (I1109752,I1109744);
not I_65069 (I1109769,I996920);
nand I_65070 (I1109786,I1109769,I996941);
and I_65071 (I1109803,I1109605,I1109786);
nor I_65072 (I1109820,I1109718,I1109803);
DFFARX1 I_65073 (I1109820,I3563,I1109523,I1109491,);
DFFARX1 I_65074 (I1109803,I3563,I1109523,I1109512,);
nor I_65075 (I1109865,I996920,I996932);
nor I_65076 (I1109503,I1109718,I1109865);
or I_65077 (I1109896,I996920,I996932);
nor I_65078 (I1109913,I996917,I996929);
DFFARX1 I_65079 (I1109913,I3563,I1109523,I1109939,);
not I_65080 (I1109947,I1109939);
nor I_65081 (I1109509,I1109947,I1109752);
nand I_65082 (I1109978,I1109947,I1109597);
not I_65083 (I1109995,I996917);
nand I_65084 (I1110012,I1109995,I1109701);
nand I_65085 (I1110029,I1109947,I1110012);
nand I_65086 (I1109500,I1110029,I1109978);
nand I_65087 (I1109497,I1110012,I1109896);
not I_65088 (I1110101,I3570);
DFFARX1 I_65089 (I92507,I3563,I1110101,I1110127,);
and I_65090 (I1110135,I1110127,I92483);
DFFARX1 I_65091 (I1110135,I3563,I1110101,I1110084,);
DFFARX1 I_65092 (I92501,I3563,I1110101,I1110175,);
not I_65093 (I1110183,I92489);
not I_65094 (I1110200,I92486);
nand I_65095 (I1110217,I1110200,I1110183);
nor I_65096 (I1110072,I1110175,I1110217);
DFFARX1 I_65097 (I1110217,I3563,I1110101,I1110257,);
not I_65098 (I1110093,I1110257);
not I_65099 (I1110279,I92495);
nand I_65100 (I1110296,I1110200,I1110279);
DFFARX1 I_65101 (I1110296,I3563,I1110101,I1110322,);
not I_65102 (I1110330,I1110322);
not I_65103 (I1110347,I92486);
nand I_65104 (I1110364,I1110347,I92504);
and I_65105 (I1110381,I1110183,I1110364);
nor I_65106 (I1110398,I1110296,I1110381);
DFFARX1 I_65107 (I1110398,I3563,I1110101,I1110069,);
DFFARX1 I_65108 (I1110381,I3563,I1110101,I1110090,);
nor I_65109 (I1110443,I92486,I92498);
nor I_65110 (I1110081,I1110296,I1110443);
or I_65111 (I1110474,I92486,I92498);
nor I_65112 (I1110491,I92492,I92483);
DFFARX1 I_65113 (I1110491,I3563,I1110101,I1110517,);
not I_65114 (I1110525,I1110517);
nor I_65115 (I1110087,I1110525,I1110330);
nand I_65116 (I1110556,I1110525,I1110175);
not I_65117 (I1110573,I92492);
nand I_65118 (I1110590,I1110573,I1110279);
nand I_65119 (I1110607,I1110525,I1110590);
nand I_65120 (I1110078,I1110607,I1110556);
nand I_65121 (I1110075,I1110590,I1110474);
not I_65122 (I1110679,I3570);
DFFARX1 I_65123 (I227378,I3563,I1110679,I1110705,);
and I_65124 (I1110713,I1110705,I227381);
DFFARX1 I_65125 (I1110713,I3563,I1110679,I1110662,);
DFFARX1 I_65126 (I227381,I3563,I1110679,I1110753,);
not I_65127 (I1110761,I227396);
not I_65128 (I1110778,I227402);
nand I_65129 (I1110795,I1110778,I1110761);
nor I_65130 (I1110650,I1110753,I1110795);
DFFARX1 I_65131 (I1110795,I3563,I1110679,I1110835,);
not I_65132 (I1110671,I1110835);
not I_65133 (I1110857,I227390);
nand I_65134 (I1110874,I1110778,I1110857);
DFFARX1 I_65135 (I1110874,I3563,I1110679,I1110900,);
not I_65136 (I1110908,I1110900);
not I_65137 (I1110925,I227387);
nand I_65138 (I1110942,I1110925,I227384);
and I_65139 (I1110959,I1110761,I1110942);
nor I_65140 (I1110976,I1110874,I1110959);
DFFARX1 I_65141 (I1110976,I3563,I1110679,I1110647,);
DFFARX1 I_65142 (I1110959,I3563,I1110679,I1110668,);
nor I_65143 (I1111021,I227387,I227378);
nor I_65144 (I1110659,I1110874,I1111021);
or I_65145 (I1111052,I227387,I227378);
nor I_65146 (I1111069,I227393,I227399);
DFFARX1 I_65147 (I1111069,I3563,I1110679,I1111095,);
not I_65148 (I1111103,I1111095);
nor I_65149 (I1110665,I1111103,I1110908);
nand I_65150 (I1111134,I1111103,I1110753);
not I_65151 (I1111151,I227393);
nand I_65152 (I1111168,I1111151,I1110857);
nand I_65153 (I1111185,I1111103,I1111168);
nand I_65154 (I1110656,I1111185,I1111134);
nand I_65155 (I1110653,I1111168,I1111052);
not I_65156 (I1111257,I3570);
DFFARX1 I_65157 (I693686,I3563,I1111257,I1111283,);
and I_65158 (I1111291,I1111283,I693674);
DFFARX1 I_65159 (I1111291,I3563,I1111257,I1111240,);
DFFARX1 I_65160 (I693677,I3563,I1111257,I1111331,);
not I_65161 (I1111339,I693671);
not I_65162 (I1111356,I693695);
nand I_65163 (I1111373,I1111356,I1111339);
nor I_65164 (I1111228,I1111331,I1111373);
DFFARX1 I_65165 (I1111373,I3563,I1111257,I1111413,);
not I_65166 (I1111249,I1111413);
not I_65167 (I1111435,I693683);
nand I_65168 (I1111452,I1111356,I1111435);
DFFARX1 I_65169 (I1111452,I3563,I1111257,I1111478,);
not I_65170 (I1111486,I1111478);
not I_65171 (I1111503,I693692);
nand I_65172 (I1111520,I1111503,I693689);
and I_65173 (I1111537,I1111339,I1111520);
nor I_65174 (I1111554,I1111452,I1111537);
DFFARX1 I_65175 (I1111554,I3563,I1111257,I1111225,);
DFFARX1 I_65176 (I1111537,I3563,I1111257,I1111246,);
nor I_65177 (I1111599,I693692,I693680);
nor I_65178 (I1111237,I1111452,I1111599);
or I_65179 (I1111630,I693692,I693680);
nor I_65180 (I1111647,I693671,I693674);
DFFARX1 I_65181 (I1111647,I3563,I1111257,I1111673,);
not I_65182 (I1111681,I1111673);
nor I_65183 (I1111243,I1111681,I1111486);
nand I_65184 (I1111712,I1111681,I1111331);
not I_65185 (I1111729,I693671);
nand I_65186 (I1111746,I1111729,I1111435);
nand I_65187 (I1111763,I1111681,I1111746);
nand I_65188 (I1111234,I1111763,I1111712);
nand I_65189 (I1111231,I1111746,I1111630);
not I_65190 (I1111835,I3570);
DFFARX1 I_65191 (I372347,I3563,I1111835,I1111861,);
and I_65192 (I1111869,I1111861,I372332);
DFFARX1 I_65193 (I1111869,I3563,I1111835,I1111818,);
DFFARX1 I_65194 (I372338,I3563,I1111835,I1111909,);
not I_65195 (I1111917,I372320);
not I_65196 (I1111934,I372341);
nand I_65197 (I1111951,I1111934,I1111917);
nor I_65198 (I1111806,I1111909,I1111951);
DFFARX1 I_65199 (I1111951,I3563,I1111835,I1111991,);
not I_65200 (I1111827,I1111991);
not I_65201 (I1112013,I372344);
nand I_65202 (I1112030,I1111934,I1112013);
DFFARX1 I_65203 (I1112030,I3563,I1111835,I1112056,);
not I_65204 (I1112064,I1112056);
not I_65205 (I1112081,I372335);
nand I_65206 (I1112098,I1112081,I372323);
and I_65207 (I1112115,I1111917,I1112098);
nor I_65208 (I1112132,I1112030,I1112115);
DFFARX1 I_65209 (I1112132,I3563,I1111835,I1111803,);
DFFARX1 I_65210 (I1112115,I3563,I1111835,I1111824,);
nor I_65211 (I1112177,I372335,I372329);
nor I_65212 (I1111815,I1112030,I1112177);
or I_65213 (I1112208,I372335,I372329);
nor I_65214 (I1112225,I372326,I372320);
DFFARX1 I_65215 (I1112225,I3563,I1111835,I1112251,);
not I_65216 (I1112259,I1112251);
nor I_65217 (I1111821,I1112259,I1112064);
nand I_65218 (I1112290,I1112259,I1111909);
not I_65219 (I1112307,I372326);
nand I_65220 (I1112324,I1112307,I1112013);
nand I_65221 (I1112341,I1112259,I1112324);
nand I_65222 (I1111812,I1112341,I1112290);
nand I_65223 (I1111809,I1112324,I1112208);
not I_65224 (I1112413,I3570);
DFFARX1 I_65225 (I1347620,I3563,I1112413,I1112439,);
and I_65226 (I1112447,I1112439,I1347602);
DFFARX1 I_65227 (I1112447,I3563,I1112413,I1112396,);
DFFARX1 I_65228 (I1347593,I3563,I1112413,I1112487,);
not I_65229 (I1112495,I1347608);
not I_65230 (I1112512,I1347596);
nand I_65231 (I1112529,I1112512,I1112495);
nor I_65232 (I1112384,I1112487,I1112529);
DFFARX1 I_65233 (I1112529,I3563,I1112413,I1112569,);
not I_65234 (I1112405,I1112569);
not I_65235 (I1112591,I1347605);
nand I_65236 (I1112608,I1112512,I1112591);
DFFARX1 I_65237 (I1112608,I3563,I1112413,I1112634,);
not I_65238 (I1112642,I1112634);
not I_65239 (I1112659,I1347614);
nand I_65240 (I1112676,I1112659,I1347593);
and I_65241 (I1112693,I1112495,I1112676);
nor I_65242 (I1112710,I1112608,I1112693);
DFFARX1 I_65243 (I1112710,I3563,I1112413,I1112381,);
DFFARX1 I_65244 (I1112693,I3563,I1112413,I1112402,);
nor I_65245 (I1112755,I1347614,I1347617);
nor I_65246 (I1112393,I1112608,I1112755);
or I_65247 (I1112786,I1347614,I1347617);
nor I_65248 (I1112803,I1347611,I1347599);
DFFARX1 I_65249 (I1112803,I3563,I1112413,I1112829,);
not I_65250 (I1112837,I1112829);
nor I_65251 (I1112399,I1112837,I1112642);
nand I_65252 (I1112868,I1112837,I1112487);
not I_65253 (I1112885,I1347611);
nand I_65254 (I1112902,I1112885,I1112591);
nand I_65255 (I1112919,I1112837,I1112902);
nand I_65256 (I1112390,I1112919,I1112868);
nand I_65257 (I1112387,I1112902,I1112786);
not I_65258 (I1112991,I3570);
DFFARX1 I_65259 (I492034,I3563,I1112991,I1113017,);
and I_65260 (I1113025,I1113017,I492049);
DFFARX1 I_65261 (I1113025,I3563,I1112991,I1112974,);
DFFARX1 I_65262 (I492052,I3563,I1112991,I1113065,);
not I_65263 (I1113073,I492046);
not I_65264 (I1113090,I492061);
nand I_65265 (I1113107,I1113090,I1113073);
nor I_65266 (I1112962,I1113065,I1113107);
DFFARX1 I_65267 (I1113107,I3563,I1112991,I1113147,);
not I_65268 (I1112983,I1113147);
not I_65269 (I1113169,I492037);
nand I_65270 (I1113186,I1113090,I1113169);
DFFARX1 I_65271 (I1113186,I3563,I1112991,I1113212,);
not I_65272 (I1113220,I1113212);
not I_65273 (I1113237,I492040);
nand I_65274 (I1113254,I1113237,I492034);
and I_65275 (I1113271,I1113073,I1113254);
nor I_65276 (I1113288,I1113186,I1113271);
DFFARX1 I_65277 (I1113288,I3563,I1112991,I1112959,);
DFFARX1 I_65278 (I1113271,I3563,I1112991,I1112980,);
nor I_65279 (I1113333,I492040,I492043);
nor I_65280 (I1112971,I1113186,I1113333);
or I_65281 (I1113364,I492040,I492043);
nor I_65282 (I1113381,I492058,I492055);
DFFARX1 I_65283 (I1113381,I3563,I1112991,I1113407,);
not I_65284 (I1113415,I1113407);
nor I_65285 (I1112977,I1113415,I1113220);
nand I_65286 (I1113446,I1113415,I1113065);
not I_65287 (I1113463,I492058);
nand I_65288 (I1113480,I1113463,I1113169);
nand I_65289 (I1113497,I1113415,I1113480);
nand I_65290 (I1112968,I1113497,I1113446);
nand I_65291 (I1112965,I1113480,I1113364);
not I_65292 (I1113569,I3570);
DFFARX1 I_65293 (I595426,I3563,I1113569,I1113595,);
and I_65294 (I1113603,I1113595,I595414);
DFFARX1 I_65295 (I1113603,I3563,I1113569,I1113552,);
DFFARX1 I_65296 (I595429,I3563,I1113569,I1113643,);
not I_65297 (I1113651,I595420);
not I_65298 (I1113668,I595411);
nand I_65299 (I1113685,I1113668,I1113651);
nor I_65300 (I1113540,I1113643,I1113685);
DFFARX1 I_65301 (I1113685,I3563,I1113569,I1113725,);
not I_65302 (I1113561,I1113725);
not I_65303 (I1113747,I595417);
nand I_65304 (I1113764,I1113668,I1113747);
DFFARX1 I_65305 (I1113764,I3563,I1113569,I1113790,);
not I_65306 (I1113798,I1113790);
not I_65307 (I1113815,I595432);
nand I_65308 (I1113832,I1113815,I595435);
and I_65309 (I1113849,I1113651,I1113832);
nor I_65310 (I1113866,I1113764,I1113849);
DFFARX1 I_65311 (I1113866,I3563,I1113569,I1113537,);
DFFARX1 I_65312 (I1113849,I3563,I1113569,I1113558,);
nor I_65313 (I1113911,I595432,I595411);
nor I_65314 (I1113549,I1113764,I1113911);
or I_65315 (I1113942,I595432,I595411);
nor I_65316 (I1113959,I595423,I595414);
DFFARX1 I_65317 (I1113959,I3563,I1113569,I1113985,);
not I_65318 (I1113993,I1113985);
nor I_65319 (I1113555,I1113993,I1113798);
nand I_65320 (I1114024,I1113993,I1113643);
not I_65321 (I1114041,I595423);
nand I_65322 (I1114058,I1114041,I1113747);
nand I_65323 (I1114075,I1113993,I1114058);
nand I_65324 (I1113546,I1114075,I1114024);
nand I_65325 (I1113543,I1114058,I1113942);
not I_65326 (I1114147,I3570);
DFFARX1 I_65327 (I488226,I3563,I1114147,I1114173,);
and I_65328 (I1114181,I1114173,I488241);
DFFARX1 I_65329 (I1114181,I3563,I1114147,I1114130,);
DFFARX1 I_65330 (I488244,I3563,I1114147,I1114221,);
not I_65331 (I1114229,I488238);
not I_65332 (I1114246,I488253);
nand I_65333 (I1114263,I1114246,I1114229);
nor I_65334 (I1114118,I1114221,I1114263);
DFFARX1 I_65335 (I1114263,I3563,I1114147,I1114303,);
not I_65336 (I1114139,I1114303);
not I_65337 (I1114325,I488229);
nand I_65338 (I1114342,I1114246,I1114325);
DFFARX1 I_65339 (I1114342,I3563,I1114147,I1114368,);
not I_65340 (I1114376,I1114368);
not I_65341 (I1114393,I488232);
nand I_65342 (I1114410,I1114393,I488226);
and I_65343 (I1114427,I1114229,I1114410);
nor I_65344 (I1114444,I1114342,I1114427);
DFFARX1 I_65345 (I1114444,I3563,I1114147,I1114115,);
DFFARX1 I_65346 (I1114427,I3563,I1114147,I1114136,);
nor I_65347 (I1114489,I488232,I488235);
nor I_65348 (I1114127,I1114342,I1114489);
or I_65349 (I1114520,I488232,I488235);
nor I_65350 (I1114537,I488250,I488247);
DFFARX1 I_65351 (I1114537,I3563,I1114147,I1114563,);
not I_65352 (I1114571,I1114563);
nor I_65353 (I1114133,I1114571,I1114376);
nand I_65354 (I1114602,I1114571,I1114221);
not I_65355 (I1114619,I488250);
nand I_65356 (I1114636,I1114619,I1114325);
nand I_65357 (I1114653,I1114571,I1114636);
nand I_65358 (I1114124,I1114653,I1114602);
nand I_65359 (I1114121,I1114636,I1114520);
not I_65360 (I1114725,I3570);
DFFARX1 I_65361 (I91980,I3563,I1114725,I1114751,);
and I_65362 (I1114759,I1114751,I91956);
DFFARX1 I_65363 (I1114759,I3563,I1114725,I1114708,);
DFFARX1 I_65364 (I91974,I3563,I1114725,I1114799,);
not I_65365 (I1114807,I91962);
not I_65366 (I1114824,I91959);
nand I_65367 (I1114841,I1114824,I1114807);
nor I_65368 (I1114696,I1114799,I1114841);
DFFARX1 I_65369 (I1114841,I3563,I1114725,I1114881,);
not I_65370 (I1114717,I1114881);
not I_65371 (I1114903,I91968);
nand I_65372 (I1114920,I1114824,I1114903);
DFFARX1 I_65373 (I1114920,I3563,I1114725,I1114946,);
not I_65374 (I1114954,I1114946);
not I_65375 (I1114971,I91959);
nand I_65376 (I1114988,I1114971,I91977);
and I_65377 (I1115005,I1114807,I1114988);
nor I_65378 (I1115022,I1114920,I1115005);
DFFARX1 I_65379 (I1115022,I3563,I1114725,I1114693,);
DFFARX1 I_65380 (I1115005,I3563,I1114725,I1114714,);
nor I_65381 (I1115067,I91959,I91971);
nor I_65382 (I1114705,I1114920,I1115067);
or I_65383 (I1115098,I91959,I91971);
nor I_65384 (I1115115,I91965,I91956);
DFFARX1 I_65385 (I1115115,I3563,I1114725,I1115141,);
not I_65386 (I1115149,I1115141);
nor I_65387 (I1114711,I1115149,I1114954);
nand I_65388 (I1115180,I1115149,I1114799);
not I_65389 (I1115197,I91965);
nand I_65390 (I1115214,I1115197,I1114903);
nand I_65391 (I1115231,I1115149,I1115214);
nand I_65392 (I1114702,I1115231,I1115180);
nand I_65393 (I1114699,I1115214,I1115098);
not I_65394 (I1115303,I3570);
DFFARX1 I_65395 (I731834,I3563,I1115303,I1115329,);
and I_65396 (I1115337,I1115329,I731822);
DFFARX1 I_65397 (I1115337,I3563,I1115303,I1115286,);
DFFARX1 I_65398 (I731825,I3563,I1115303,I1115377,);
not I_65399 (I1115385,I731819);
not I_65400 (I1115402,I731843);
nand I_65401 (I1115419,I1115402,I1115385);
nor I_65402 (I1115274,I1115377,I1115419);
DFFARX1 I_65403 (I1115419,I3563,I1115303,I1115459,);
not I_65404 (I1115295,I1115459);
not I_65405 (I1115481,I731831);
nand I_65406 (I1115498,I1115402,I1115481);
DFFARX1 I_65407 (I1115498,I3563,I1115303,I1115524,);
not I_65408 (I1115532,I1115524);
not I_65409 (I1115549,I731840);
nand I_65410 (I1115566,I1115549,I731837);
and I_65411 (I1115583,I1115385,I1115566);
nor I_65412 (I1115600,I1115498,I1115583);
DFFARX1 I_65413 (I1115600,I3563,I1115303,I1115271,);
DFFARX1 I_65414 (I1115583,I3563,I1115303,I1115292,);
nor I_65415 (I1115645,I731840,I731828);
nor I_65416 (I1115283,I1115498,I1115645);
or I_65417 (I1115676,I731840,I731828);
nor I_65418 (I1115693,I731819,I731822);
DFFARX1 I_65419 (I1115693,I3563,I1115303,I1115719,);
not I_65420 (I1115727,I1115719);
nor I_65421 (I1115289,I1115727,I1115532);
nand I_65422 (I1115758,I1115727,I1115377);
not I_65423 (I1115775,I731819);
nand I_65424 (I1115792,I1115775,I1115481);
nand I_65425 (I1115809,I1115727,I1115792);
nand I_65426 (I1115280,I1115809,I1115758);
nand I_65427 (I1115277,I1115792,I1115676);
not I_65428 (I1115881,I3570);
DFFARX1 I_65429 (I337038,I3563,I1115881,I1115907,);
and I_65430 (I1115915,I1115907,I337023);
DFFARX1 I_65431 (I1115915,I3563,I1115881,I1115864,);
DFFARX1 I_65432 (I337029,I3563,I1115881,I1115955,);
not I_65433 (I1115963,I337011);
not I_65434 (I1115980,I337032);
nand I_65435 (I1115997,I1115980,I1115963);
nor I_65436 (I1115852,I1115955,I1115997);
DFFARX1 I_65437 (I1115997,I3563,I1115881,I1116037,);
not I_65438 (I1115873,I1116037);
not I_65439 (I1116059,I337035);
nand I_65440 (I1116076,I1115980,I1116059);
DFFARX1 I_65441 (I1116076,I3563,I1115881,I1116102,);
not I_65442 (I1116110,I1116102);
not I_65443 (I1116127,I337026);
nand I_65444 (I1116144,I1116127,I337014);
and I_65445 (I1116161,I1115963,I1116144);
nor I_65446 (I1116178,I1116076,I1116161);
DFFARX1 I_65447 (I1116178,I3563,I1115881,I1115849,);
DFFARX1 I_65448 (I1116161,I3563,I1115881,I1115870,);
nor I_65449 (I1116223,I337026,I337020);
nor I_65450 (I1115861,I1116076,I1116223);
or I_65451 (I1116254,I337026,I337020);
nor I_65452 (I1116271,I337017,I337011);
DFFARX1 I_65453 (I1116271,I3563,I1115881,I1116297,);
not I_65454 (I1116305,I1116297);
nor I_65455 (I1115867,I1116305,I1116110);
nand I_65456 (I1116336,I1116305,I1115955);
not I_65457 (I1116353,I337017);
nand I_65458 (I1116370,I1116353,I1116059);
nand I_65459 (I1116387,I1116305,I1116370);
nand I_65460 (I1115858,I1116387,I1116336);
nand I_65461 (I1115855,I1116370,I1116254);
not I_65462 (I1116459,I3570);
DFFARX1 I_65463 (I878515,I3563,I1116459,I1116485,);
and I_65464 (I1116493,I1116485,I878521);
DFFARX1 I_65465 (I1116493,I3563,I1116459,I1116442,);
DFFARX1 I_65466 (I878527,I3563,I1116459,I1116533,);
not I_65467 (I1116541,I878512);
not I_65468 (I1116558,I878512);
nand I_65469 (I1116575,I1116558,I1116541);
nor I_65470 (I1116430,I1116533,I1116575);
DFFARX1 I_65471 (I1116575,I3563,I1116459,I1116615,);
not I_65472 (I1116451,I1116615);
not I_65473 (I1116637,I878530);
nand I_65474 (I1116654,I1116558,I1116637);
DFFARX1 I_65475 (I1116654,I3563,I1116459,I1116680,);
not I_65476 (I1116688,I1116680);
not I_65477 (I1116705,I878524);
nand I_65478 (I1116722,I1116705,I878515);
and I_65479 (I1116739,I1116541,I1116722);
nor I_65480 (I1116756,I1116654,I1116739);
DFFARX1 I_65481 (I1116756,I3563,I1116459,I1116427,);
DFFARX1 I_65482 (I1116739,I3563,I1116459,I1116448,);
nor I_65483 (I1116801,I878524,I878533);
nor I_65484 (I1116439,I1116654,I1116801);
or I_65485 (I1116832,I878524,I878533);
nor I_65486 (I1116849,I878518,I878518);
DFFARX1 I_65487 (I1116849,I3563,I1116459,I1116875,);
not I_65488 (I1116883,I1116875);
nor I_65489 (I1116445,I1116883,I1116688);
nand I_65490 (I1116914,I1116883,I1116533);
not I_65491 (I1116931,I878518);
nand I_65492 (I1116948,I1116931,I1116637);
nand I_65493 (I1116965,I1116883,I1116948);
nand I_65494 (I1116436,I1116965,I1116914);
nand I_65495 (I1116433,I1116948,I1116832);
not I_65496 (I1117037,I3570);
DFFARX1 I_65497 (I1016949,I3563,I1117037,I1117063,);
and I_65498 (I1117071,I1117063,I1016943);
DFFARX1 I_65499 (I1117071,I3563,I1117037,I1117020,);
DFFARX1 I_65500 (I1016961,I3563,I1117037,I1117111,);
not I_65501 (I1117119,I1016952);
not I_65502 (I1117136,I1016964);
nand I_65503 (I1117153,I1117136,I1117119);
nor I_65504 (I1117008,I1117111,I1117153);
DFFARX1 I_65505 (I1117153,I3563,I1117037,I1117193,);
not I_65506 (I1117029,I1117193);
not I_65507 (I1117215,I1016970);
nand I_65508 (I1117232,I1117136,I1117215);
DFFARX1 I_65509 (I1117232,I3563,I1117037,I1117258,);
not I_65510 (I1117266,I1117258);
not I_65511 (I1117283,I1016946);
nand I_65512 (I1117300,I1117283,I1016967);
and I_65513 (I1117317,I1117119,I1117300);
nor I_65514 (I1117334,I1117232,I1117317);
DFFARX1 I_65515 (I1117334,I3563,I1117037,I1117005,);
DFFARX1 I_65516 (I1117317,I3563,I1117037,I1117026,);
nor I_65517 (I1117379,I1016946,I1016958);
nor I_65518 (I1117017,I1117232,I1117379);
or I_65519 (I1117410,I1016946,I1016958);
nor I_65520 (I1117427,I1016943,I1016955);
DFFARX1 I_65521 (I1117427,I3563,I1117037,I1117453,);
not I_65522 (I1117461,I1117453);
nor I_65523 (I1117023,I1117461,I1117266);
nand I_65524 (I1117492,I1117461,I1117111);
not I_65525 (I1117509,I1016943);
nand I_65526 (I1117526,I1117509,I1117215);
nand I_65527 (I1117543,I1117461,I1117526);
nand I_65528 (I1117014,I1117543,I1117492);
nand I_65529 (I1117011,I1117526,I1117410);
not I_65530 (I1117615,I3570);
DFFARX1 I_65531 (I1345240,I3563,I1117615,I1117641,);
and I_65532 (I1117649,I1117641,I1345222);
DFFARX1 I_65533 (I1117649,I3563,I1117615,I1117598,);
DFFARX1 I_65534 (I1345213,I3563,I1117615,I1117689,);
not I_65535 (I1117697,I1345228);
not I_65536 (I1117714,I1345216);
nand I_65537 (I1117731,I1117714,I1117697);
nor I_65538 (I1117586,I1117689,I1117731);
DFFARX1 I_65539 (I1117731,I3563,I1117615,I1117771,);
not I_65540 (I1117607,I1117771);
not I_65541 (I1117793,I1345225);
nand I_65542 (I1117810,I1117714,I1117793);
DFFARX1 I_65543 (I1117810,I3563,I1117615,I1117836,);
not I_65544 (I1117844,I1117836);
not I_65545 (I1117861,I1345234);
nand I_65546 (I1117878,I1117861,I1345213);
and I_65547 (I1117895,I1117697,I1117878);
nor I_65548 (I1117912,I1117810,I1117895);
DFFARX1 I_65549 (I1117912,I3563,I1117615,I1117583,);
DFFARX1 I_65550 (I1117895,I3563,I1117615,I1117604,);
nor I_65551 (I1117957,I1345234,I1345237);
nor I_65552 (I1117595,I1117810,I1117957);
or I_65553 (I1117988,I1345234,I1345237);
nor I_65554 (I1118005,I1345231,I1345219);
DFFARX1 I_65555 (I1118005,I3563,I1117615,I1118031,);
not I_65556 (I1118039,I1118031);
nor I_65557 (I1117601,I1118039,I1117844);
nand I_65558 (I1118070,I1118039,I1117689);
not I_65559 (I1118087,I1345231);
nand I_65560 (I1118104,I1118087,I1117793);
nand I_65561 (I1118121,I1118039,I1118104);
nand I_65562 (I1117592,I1118121,I1118070);
nand I_65563 (I1117589,I1118104,I1117988);
not I_65564 (I1118193,I3570);
DFFARX1 I_65565 (I968499,I3563,I1118193,I1118219,);
and I_65566 (I1118227,I1118219,I968493);
DFFARX1 I_65567 (I1118227,I3563,I1118193,I1118176,);
DFFARX1 I_65568 (I968511,I3563,I1118193,I1118267,);
not I_65569 (I1118275,I968502);
not I_65570 (I1118292,I968514);
nand I_65571 (I1118309,I1118292,I1118275);
nor I_65572 (I1118164,I1118267,I1118309);
DFFARX1 I_65573 (I1118309,I3563,I1118193,I1118349,);
not I_65574 (I1118185,I1118349);
not I_65575 (I1118371,I968520);
nand I_65576 (I1118388,I1118292,I1118371);
DFFARX1 I_65577 (I1118388,I3563,I1118193,I1118414,);
not I_65578 (I1118422,I1118414);
not I_65579 (I1118439,I968496);
nand I_65580 (I1118456,I1118439,I968517);
and I_65581 (I1118473,I1118275,I1118456);
nor I_65582 (I1118490,I1118388,I1118473);
DFFARX1 I_65583 (I1118490,I3563,I1118193,I1118161,);
DFFARX1 I_65584 (I1118473,I3563,I1118193,I1118182,);
nor I_65585 (I1118535,I968496,I968508);
nor I_65586 (I1118173,I1118388,I1118535);
or I_65587 (I1118566,I968496,I968508);
nor I_65588 (I1118583,I968493,I968505);
DFFARX1 I_65589 (I1118583,I3563,I1118193,I1118609,);
not I_65590 (I1118617,I1118609);
nor I_65591 (I1118179,I1118617,I1118422);
nand I_65592 (I1118648,I1118617,I1118267);
not I_65593 (I1118665,I968493);
nand I_65594 (I1118682,I1118665,I1118371);
nand I_65595 (I1118699,I1118617,I1118682);
nand I_65596 (I1118170,I1118699,I1118648);
nand I_65597 (I1118167,I1118682,I1118566);
not I_65598 (I1118771,I3570);
DFFARX1 I_65599 (I539399,I3563,I1118771,I1118797,);
and I_65600 (I1118805,I1118797,I539414);
DFFARX1 I_65601 (I1118805,I3563,I1118771,I1118754,);
DFFARX1 I_65602 (I539405,I3563,I1118771,I1118845,);
not I_65603 (I1118853,I539399);
not I_65604 (I1118870,I539417);
nand I_65605 (I1118887,I1118870,I1118853);
nor I_65606 (I1118742,I1118845,I1118887);
DFFARX1 I_65607 (I1118887,I3563,I1118771,I1118927,);
not I_65608 (I1118763,I1118927);
not I_65609 (I1118949,I539408);
nand I_65610 (I1118966,I1118870,I1118949);
DFFARX1 I_65611 (I1118966,I3563,I1118771,I1118992,);
not I_65612 (I1119000,I1118992);
not I_65613 (I1119017,I539420);
nand I_65614 (I1119034,I1119017,I539396);
and I_65615 (I1119051,I1118853,I1119034);
nor I_65616 (I1119068,I1118966,I1119051);
DFFARX1 I_65617 (I1119068,I3563,I1118771,I1118739,);
DFFARX1 I_65618 (I1119051,I3563,I1118771,I1118760,);
nor I_65619 (I1119113,I539420,I539396);
nor I_65620 (I1118751,I1118966,I1119113);
or I_65621 (I1119144,I539420,I539396);
nor I_65622 (I1119161,I539402,I539411);
DFFARX1 I_65623 (I1119161,I3563,I1118771,I1119187,);
not I_65624 (I1119195,I1119187);
nor I_65625 (I1118757,I1119195,I1119000);
nand I_65626 (I1119226,I1119195,I1118845);
not I_65627 (I1119243,I539402);
nand I_65628 (I1119260,I1119243,I1118949);
nand I_65629 (I1119277,I1119195,I1119260);
nand I_65630 (I1118748,I1119277,I1119226);
nand I_65631 (I1118745,I1119260,I1119144);
not I_65632 (I1119349,I3570);
DFFARX1 I_65633 (I538804,I3563,I1119349,I1119375,);
and I_65634 (I1119383,I1119375,I538819);
DFFARX1 I_65635 (I1119383,I3563,I1119349,I1119332,);
DFFARX1 I_65636 (I538810,I3563,I1119349,I1119423,);
not I_65637 (I1119431,I538804);
not I_65638 (I1119448,I538822);
nand I_65639 (I1119465,I1119448,I1119431);
nor I_65640 (I1119320,I1119423,I1119465);
DFFARX1 I_65641 (I1119465,I3563,I1119349,I1119505,);
not I_65642 (I1119341,I1119505);
not I_65643 (I1119527,I538813);
nand I_65644 (I1119544,I1119448,I1119527);
DFFARX1 I_65645 (I1119544,I3563,I1119349,I1119570,);
not I_65646 (I1119578,I1119570);
not I_65647 (I1119595,I538825);
nand I_65648 (I1119612,I1119595,I538801);
and I_65649 (I1119629,I1119431,I1119612);
nor I_65650 (I1119646,I1119544,I1119629);
DFFARX1 I_65651 (I1119646,I3563,I1119349,I1119317,);
DFFARX1 I_65652 (I1119629,I3563,I1119349,I1119338,);
nor I_65653 (I1119691,I538825,I538801);
nor I_65654 (I1119329,I1119544,I1119691);
or I_65655 (I1119722,I538825,I538801);
nor I_65656 (I1119739,I538807,I538816);
DFFARX1 I_65657 (I1119739,I3563,I1119349,I1119765,);
not I_65658 (I1119773,I1119765);
nor I_65659 (I1119335,I1119773,I1119578);
nand I_65660 (I1119804,I1119773,I1119423);
not I_65661 (I1119821,I538807);
nand I_65662 (I1119838,I1119821,I1119527);
nand I_65663 (I1119855,I1119773,I1119838);
nand I_65664 (I1119326,I1119855,I1119804);
nand I_65665 (I1119323,I1119838,I1119722);
not I_65666 (I1119927,I3570);
DFFARX1 I_65667 (I1256766,I3563,I1119927,I1119953,);
and I_65668 (I1119961,I1119953,I1256760);
DFFARX1 I_65669 (I1119961,I3563,I1119927,I1119910,);
DFFARX1 I_65670 (I1256745,I3563,I1119927,I1120001,);
not I_65671 (I1120009,I1256751);
not I_65672 (I1120026,I1256763);
nand I_65673 (I1120043,I1120026,I1120009);
nor I_65674 (I1119898,I1120001,I1120043);
DFFARX1 I_65675 (I1120043,I3563,I1119927,I1120083,);
not I_65676 (I1119919,I1120083);
not I_65677 (I1120105,I1256745);
nand I_65678 (I1120122,I1120026,I1120105);
DFFARX1 I_65679 (I1120122,I3563,I1119927,I1120148,);
not I_65680 (I1120156,I1120148);
not I_65681 (I1120173,I1256769);
nand I_65682 (I1120190,I1120173,I1256757);
and I_65683 (I1120207,I1120009,I1120190);
nor I_65684 (I1120224,I1120122,I1120207);
DFFARX1 I_65685 (I1120224,I3563,I1119927,I1119895,);
DFFARX1 I_65686 (I1120207,I3563,I1119927,I1119916,);
nor I_65687 (I1120269,I1256769,I1256748);
nor I_65688 (I1119907,I1120122,I1120269);
or I_65689 (I1120300,I1256769,I1256748);
nor I_65690 (I1120317,I1256754,I1256748);
DFFARX1 I_65691 (I1120317,I3563,I1119927,I1120343,);
not I_65692 (I1120351,I1120343);
nor I_65693 (I1119913,I1120351,I1120156);
nand I_65694 (I1120382,I1120351,I1120001);
not I_65695 (I1120399,I1256754);
nand I_65696 (I1120416,I1120399,I1120105);
nand I_65697 (I1120433,I1120351,I1120416);
nand I_65698 (I1119904,I1120433,I1120382);
nand I_65699 (I1119901,I1120416,I1120300);
not I_65700 (I1120505,I3570);
DFFARX1 I_65701 (I1348215,I3563,I1120505,I1120531,);
and I_65702 (I1120539,I1120531,I1348197);
DFFARX1 I_65703 (I1120539,I3563,I1120505,I1120488,);
DFFARX1 I_65704 (I1348188,I3563,I1120505,I1120579,);
not I_65705 (I1120587,I1348203);
not I_65706 (I1120604,I1348191);
nand I_65707 (I1120621,I1120604,I1120587);
nor I_65708 (I1120476,I1120579,I1120621);
DFFARX1 I_65709 (I1120621,I3563,I1120505,I1120661,);
not I_65710 (I1120497,I1120661);
not I_65711 (I1120683,I1348200);
nand I_65712 (I1120700,I1120604,I1120683);
DFFARX1 I_65713 (I1120700,I3563,I1120505,I1120726,);
not I_65714 (I1120734,I1120726);
not I_65715 (I1120751,I1348209);
nand I_65716 (I1120768,I1120751,I1348188);
and I_65717 (I1120785,I1120587,I1120768);
nor I_65718 (I1120802,I1120700,I1120785);
DFFARX1 I_65719 (I1120802,I3563,I1120505,I1120473,);
DFFARX1 I_65720 (I1120785,I3563,I1120505,I1120494,);
nor I_65721 (I1120847,I1348209,I1348212);
nor I_65722 (I1120485,I1120700,I1120847);
or I_65723 (I1120878,I1348209,I1348212);
nor I_65724 (I1120895,I1348206,I1348194);
DFFARX1 I_65725 (I1120895,I3563,I1120505,I1120921,);
not I_65726 (I1120929,I1120921);
nor I_65727 (I1120491,I1120929,I1120734);
nand I_65728 (I1120960,I1120929,I1120579);
not I_65729 (I1120977,I1348206);
nand I_65730 (I1120994,I1120977,I1120683);
nand I_65731 (I1121011,I1120929,I1120994);
nand I_65732 (I1120482,I1121011,I1120960);
nand I_65733 (I1120479,I1120994,I1120878);
not I_65734 (I1121083,I3570);
DFFARX1 I_65735 (I715072,I3563,I1121083,I1121109,);
and I_65736 (I1121117,I1121109,I715060);
DFFARX1 I_65737 (I1121117,I3563,I1121083,I1121066,);
DFFARX1 I_65738 (I715063,I3563,I1121083,I1121157,);
not I_65739 (I1121165,I715057);
not I_65740 (I1121182,I715081);
nand I_65741 (I1121199,I1121182,I1121165);
nor I_65742 (I1121054,I1121157,I1121199);
DFFARX1 I_65743 (I1121199,I3563,I1121083,I1121239,);
not I_65744 (I1121075,I1121239);
not I_65745 (I1121261,I715069);
nand I_65746 (I1121278,I1121182,I1121261);
DFFARX1 I_65747 (I1121278,I3563,I1121083,I1121304,);
not I_65748 (I1121312,I1121304);
not I_65749 (I1121329,I715078);
nand I_65750 (I1121346,I1121329,I715075);
and I_65751 (I1121363,I1121165,I1121346);
nor I_65752 (I1121380,I1121278,I1121363);
DFFARX1 I_65753 (I1121380,I3563,I1121083,I1121051,);
DFFARX1 I_65754 (I1121363,I3563,I1121083,I1121072,);
nor I_65755 (I1121425,I715078,I715066);
nor I_65756 (I1121063,I1121278,I1121425);
or I_65757 (I1121456,I715078,I715066);
nor I_65758 (I1121473,I715057,I715060);
DFFARX1 I_65759 (I1121473,I3563,I1121083,I1121499,);
not I_65760 (I1121507,I1121499);
nor I_65761 (I1121069,I1121507,I1121312);
nand I_65762 (I1121538,I1121507,I1121157);
not I_65763 (I1121555,I715057);
nand I_65764 (I1121572,I1121555,I1121261);
nand I_65765 (I1121589,I1121507,I1121572);
nand I_65766 (I1121060,I1121589,I1121538);
nand I_65767 (I1121057,I1121572,I1121456);
not I_65768 (I1121661,I3570);
DFFARX1 I_65769 (I407656,I3563,I1121661,I1121687,);
and I_65770 (I1121695,I1121687,I407641);
DFFARX1 I_65771 (I1121695,I3563,I1121661,I1121644,);
DFFARX1 I_65772 (I407647,I3563,I1121661,I1121735,);
not I_65773 (I1121743,I407629);
not I_65774 (I1121760,I407650);
nand I_65775 (I1121777,I1121760,I1121743);
nor I_65776 (I1121632,I1121735,I1121777);
DFFARX1 I_65777 (I1121777,I3563,I1121661,I1121817,);
not I_65778 (I1121653,I1121817);
not I_65779 (I1121839,I407653);
nand I_65780 (I1121856,I1121760,I1121839);
DFFARX1 I_65781 (I1121856,I3563,I1121661,I1121882,);
not I_65782 (I1121890,I1121882);
not I_65783 (I1121907,I407644);
nand I_65784 (I1121924,I1121907,I407632);
and I_65785 (I1121941,I1121743,I1121924);
nor I_65786 (I1121958,I1121856,I1121941);
DFFARX1 I_65787 (I1121958,I3563,I1121661,I1121629,);
DFFARX1 I_65788 (I1121941,I3563,I1121661,I1121650,);
nor I_65789 (I1122003,I407644,I407638);
nor I_65790 (I1121641,I1121856,I1122003);
or I_65791 (I1122034,I407644,I407638);
nor I_65792 (I1122051,I407635,I407629);
DFFARX1 I_65793 (I1122051,I3563,I1121661,I1122077,);
not I_65794 (I1122085,I1122077);
nor I_65795 (I1121647,I1122085,I1121890);
nand I_65796 (I1122116,I1122085,I1121735);
not I_65797 (I1122133,I407635);
nand I_65798 (I1122150,I1122133,I1121839);
nand I_65799 (I1122167,I1122085,I1122150);
nand I_65800 (I1121638,I1122167,I1122116);
nand I_65801 (I1121635,I1122150,I1122034);
not I_65802 (I1122239,I3570);
DFFARX1 I_65803 (I9538,I3563,I1122239,I1122265,);
and I_65804 (I1122273,I1122265,I9544);
DFFARX1 I_65805 (I1122273,I3563,I1122239,I1122222,);
DFFARX1 I_65806 (I9523,I3563,I1122239,I1122313,);
not I_65807 (I1122321,I9529);
not I_65808 (I1122338,I9535);
nand I_65809 (I1122355,I1122338,I1122321);
nor I_65810 (I1122210,I1122313,I1122355);
DFFARX1 I_65811 (I1122355,I3563,I1122239,I1122395,);
not I_65812 (I1122231,I1122395);
not I_65813 (I1122417,I9526);
nand I_65814 (I1122434,I1122338,I1122417);
DFFARX1 I_65815 (I1122434,I3563,I1122239,I1122460,);
not I_65816 (I1122468,I1122460);
not I_65817 (I1122485,I9541);
nand I_65818 (I1122502,I1122485,I9526);
and I_65819 (I1122519,I1122321,I1122502);
nor I_65820 (I1122536,I1122434,I1122519);
DFFARX1 I_65821 (I1122536,I3563,I1122239,I1122207,);
DFFARX1 I_65822 (I1122519,I3563,I1122239,I1122228,);
nor I_65823 (I1122581,I9541,I9529);
nor I_65824 (I1122219,I1122434,I1122581);
or I_65825 (I1122612,I9541,I9529);
nor I_65826 (I1122629,I9532,I9523);
DFFARX1 I_65827 (I1122629,I3563,I1122239,I1122655,);
not I_65828 (I1122663,I1122655);
nor I_65829 (I1122225,I1122663,I1122468);
nand I_65830 (I1122694,I1122663,I1122313);
not I_65831 (I1122711,I9532);
nand I_65832 (I1122728,I1122711,I1122417);
nand I_65833 (I1122745,I1122663,I1122728);
nand I_65834 (I1122216,I1122745,I1122694);
nand I_65835 (I1122213,I1122728,I1122612);
not I_65836 (I1122817,I3570);
DFFARX1 I_65837 (I1377965,I3563,I1122817,I1122843,);
and I_65838 (I1122851,I1122843,I1377947);
DFFARX1 I_65839 (I1122851,I3563,I1122817,I1122800,);
DFFARX1 I_65840 (I1377938,I3563,I1122817,I1122891,);
not I_65841 (I1122899,I1377953);
not I_65842 (I1122916,I1377941);
nand I_65843 (I1122933,I1122916,I1122899);
nor I_65844 (I1122788,I1122891,I1122933);
DFFARX1 I_65845 (I1122933,I3563,I1122817,I1122973,);
not I_65846 (I1122809,I1122973);
not I_65847 (I1122995,I1377950);
nand I_65848 (I1123012,I1122916,I1122995);
DFFARX1 I_65849 (I1123012,I3563,I1122817,I1123038,);
not I_65850 (I1123046,I1123038);
not I_65851 (I1123063,I1377959);
nand I_65852 (I1123080,I1123063,I1377938);
and I_65853 (I1123097,I1122899,I1123080);
nor I_65854 (I1123114,I1123012,I1123097);
DFFARX1 I_65855 (I1123114,I3563,I1122817,I1122785,);
DFFARX1 I_65856 (I1123097,I3563,I1122817,I1122806,);
nor I_65857 (I1123159,I1377959,I1377962);
nor I_65858 (I1122797,I1123012,I1123159);
or I_65859 (I1123190,I1377959,I1377962);
nor I_65860 (I1123207,I1377956,I1377944);
DFFARX1 I_65861 (I1123207,I3563,I1122817,I1123233,);
not I_65862 (I1123241,I1123233);
nor I_65863 (I1122803,I1123241,I1123046);
nand I_65864 (I1123272,I1123241,I1122891);
not I_65865 (I1123289,I1377956);
nand I_65866 (I1123306,I1123289,I1122995);
nand I_65867 (I1123323,I1123241,I1123306);
nand I_65868 (I1122794,I1123323,I1123272);
nand I_65869 (I1122791,I1123306,I1123190);
not I_65870 (I1123395,I3570);
DFFARX1 I_65871 (I903284,I3563,I1123395,I1123421,);
and I_65872 (I1123429,I1123421,I903290);
DFFARX1 I_65873 (I1123429,I3563,I1123395,I1123378,);
DFFARX1 I_65874 (I903296,I3563,I1123395,I1123469,);
not I_65875 (I1123477,I903281);
not I_65876 (I1123494,I903281);
nand I_65877 (I1123511,I1123494,I1123477);
nor I_65878 (I1123366,I1123469,I1123511);
DFFARX1 I_65879 (I1123511,I3563,I1123395,I1123551,);
not I_65880 (I1123387,I1123551);
not I_65881 (I1123573,I903299);
nand I_65882 (I1123590,I1123494,I1123573);
DFFARX1 I_65883 (I1123590,I3563,I1123395,I1123616,);
not I_65884 (I1123624,I1123616);
not I_65885 (I1123641,I903293);
nand I_65886 (I1123658,I1123641,I903284);
and I_65887 (I1123675,I1123477,I1123658);
nor I_65888 (I1123692,I1123590,I1123675);
DFFARX1 I_65889 (I1123692,I3563,I1123395,I1123363,);
DFFARX1 I_65890 (I1123675,I3563,I1123395,I1123384,);
nor I_65891 (I1123737,I903293,I903302);
nor I_65892 (I1123375,I1123590,I1123737);
or I_65893 (I1123768,I903293,I903302);
nor I_65894 (I1123785,I903287,I903287);
DFFARX1 I_65895 (I1123785,I3563,I1123395,I1123811,);
not I_65896 (I1123819,I1123811);
nor I_65897 (I1123381,I1123819,I1123624);
nand I_65898 (I1123850,I1123819,I1123469);
not I_65899 (I1123867,I903287);
nand I_65900 (I1123884,I1123867,I1123573);
nand I_65901 (I1123901,I1123819,I1123884);
nand I_65902 (I1123372,I1123901,I1123850);
nand I_65903 (I1123369,I1123884,I1123768);
not I_65904 (I1123973,I3570);
DFFARX1 I_65905 (I77751,I3563,I1123973,I1123999,);
and I_65906 (I1124007,I1123999,I77727);
DFFARX1 I_65907 (I1124007,I3563,I1123973,I1123956,);
DFFARX1 I_65908 (I77745,I3563,I1123973,I1124047,);
not I_65909 (I1124055,I77733);
not I_65910 (I1124072,I77730);
nand I_65911 (I1124089,I1124072,I1124055);
nor I_65912 (I1123944,I1124047,I1124089);
DFFARX1 I_65913 (I1124089,I3563,I1123973,I1124129,);
not I_65914 (I1123965,I1124129);
not I_65915 (I1124151,I77739);
nand I_65916 (I1124168,I1124072,I1124151);
DFFARX1 I_65917 (I1124168,I3563,I1123973,I1124194,);
not I_65918 (I1124202,I1124194);
not I_65919 (I1124219,I77730);
nand I_65920 (I1124236,I1124219,I77748);
and I_65921 (I1124253,I1124055,I1124236);
nor I_65922 (I1124270,I1124168,I1124253);
DFFARX1 I_65923 (I1124270,I3563,I1123973,I1123941,);
DFFARX1 I_65924 (I1124253,I3563,I1123973,I1123962,);
nor I_65925 (I1124315,I77730,I77742);
nor I_65926 (I1123953,I1124168,I1124315);
or I_65927 (I1124346,I77730,I77742);
nor I_65928 (I1124363,I77736,I77727);
DFFARX1 I_65929 (I1124363,I3563,I1123973,I1124389,);
not I_65930 (I1124397,I1124389);
nor I_65931 (I1123959,I1124397,I1124202);
nand I_65932 (I1124428,I1124397,I1124047);
not I_65933 (I1124445,I77736);
nand I_65934 (I1124462,I1124445,I1124151);
nand I_65935 (I1124479,I1124397,I1124462);
nand I_65936 (I1123950,I1124479,I1124428);
nand I_65937 (I1123947,I1124462,I1124346);
not I_65938 (I1124551,I3570);
DFFARX1 I_65939 (I783276,I3563,I1124551,I1124577,);
and I_65940 (I1124585,I1124577,I783264);
DFFARX1 I_65941 (I1124585,I3563,I1124551,I1124534,);
DFFARX1 I_65942 (I783267,I3563,I1124551,I1124625,);
not I_65943 (I1124633,I783261);
not I_65944 (I1124650,I783285);
nand I_65945 (I1124667,I1124650,I1124633);
nor I_65946 (I1124522,I1124625,I1124667);
DFFARX1 I_65947 (I1124667,I3563,I1124551,I1124707,);
not I_65948 (I1124543,I1124707);
not I_65949 (I1124729,I783273);
nand I_65950 (I1124746,I1124650,I1124729);
DFFARX1 I_65951 (I1124746,I3563,I1124551,I1124772,);
not I_65952 (I1124780,I1124772);
not I_65953 (I1124797,I783282);
nand I_65954 (I1124814,I1124797,I783279);
and I_65955 (I1124831,I1124633,I1124814);
nor I_65956 (I1124848,I1124746,I1124831);
DFFARX1 I_65957 (I1124848,I3563,I1124551,I1124519,);
DFFARX1 I_65958 (I1124831,I3563,I1124551,I1124540,);
nor I_65959 (I1124893,I783282,I783270);
nor I_65960 (I1124531,I1124746,I1124893);
or I_65961 (I1124924,I783282,I783270);
nor I_65962 (I1124941,I783261,I783264);
DFFARX1 I_65963 (I1124941,I3563,I1124551,I1124967,);
not I_65964 (I1124975,I1124967);
nor I_65965 (I1124537,I1124975,I1124780);
nand I_65966 (I1125006,I1124975,I1124625);
not I_65967 (I1125023,I783261);
nand I_65968 (I1125040,I1125023,I1124729);
nand I_65969 (I1125057,I1124975,I1125040);
nand I_65970 (I1124528,I1125057,I1125006);
nand I_65971 (I1124525,I1125040,I1124924);
not I_65972 (I1125129,I3570);
DFFARX1 I_65973 (I229758,I3563,I1125129,I1125155,);
and I_65974 (I1125163,I1125155,I229761);
DFFARX1 I_65975 (I1125163,I3563,I1125129,I1125112,);
DFFARX1 I_65976 (I229761,I3563,I1125129,I1125203,);
not I_65977 (I1125211,I229776);
not I_65978 (I1125228,I229782);
nand I_65979 (I1125245,I1125228,I1125211);
nor I_65980 (I1125100,I1125203,I1125245);
DFFARX1 I_65981 (I1125245,I3563,I1125129,I1125285,);
not I_65982 (I1125121,I1125285);
not I_65983 (I1125307,I229770);
nand I_65984 (I1125324,I1125228,I1125307);
DFFARX1 I_65985 (I1125324,I3563,I1125129,I1125350,);
not I_65986 (I1125358,I1125350);
not I_65987 (I1125375,I229767);
nand I_65988 (I1125392,I1125375,I229764);
and I_65989 (I1125409,I1125211,I1125392);
nor I_65990 (I1125426,I1125324,I1125409);
DFFARX1 I_65991 (I1125426,I3563,I1125129,I1125097,);
DFFARX1 I_65992 (I1125409,I3563,I1125129,I1125118,);
nor I_65993 (I1125471,I229767,I229758);
nor I_65994 (I1125109,I1125324,I1125471);
or I_65995 (I1125502,I229767,I229758);
nor I_65996 (I1125519,I229773,I229779);
DFFARX1 I_65997 (I1125519,I3563,I1125129,I1125545,);
not I_65998 (I1125553,I1125545);
nor I_65999 (I1125115,I1125553,I1125358);
nand I_66000 (I1125584,I1125553,I1125203);
not I_66001 (I1125601,I229773);
nand I_66002 (I1125618,I1125601,I1125307);
nand I_66003 (I1125635,I1125553,I1125618);
nand I_66004 (I1125106,I1125635,I1125584);
nand I_66005 (I1125103,I1125618,I1125502);
not I_66006 (I1125707,I3570);
DFFARX1 I_66007 (I1292401,I3563,I1125707,I1125733,);
and I_66008 (I1125741,I1125733,I1292383);
DFFARX1 I_66009 (I1125741,I3563,I1125707,I1125690,);
DFFARX1 I_66010 (I1292392,I3563,I1125707,I1125781,);
not I_66011 (I1125789,I1292377);
not I_66012 (I1125806,I1292389);
nand I_66013 (I1125823,I1125806,I1125789);
nor I_66014 (I1125678,I1125781,I1125823);
DFFARX1 I_66015 (I1125823,I3563,I1125707,I1125863,);
not I_66016 (I1125699,I1125863);
not I_66017 (I1125885,I1292380);
nand I_66018 (I1125902,I1125806,I1125885);
DFFARX1 I_66019 (I1125902,I3563,I1125707,I1125928,);
not I_66020 (I1125936,I1125928);
not I_66021 (I1125953,I1292377);
nand I_66022 (I1125970,I1125953,I1292380);
and I_66023 (I1125987,I1125789,I1125970);
nor I_66024 (I1126004,I1125902,I1125987);
DFFARX1 I_66025 (I1126004,I3563,I1125707,I1125675,);
DFFARX1 I_66026 (I1125987,I3563,I1125707,I1125696,);
nor I_66027 (I1126049,I1292377,I1292398);
nor I_66028 (I1125687,I1125902,I1126049);
or I_66029 (I1126080,I1292377,I1292398);
nor I_66030 (I1126097,I1292386,I1292395);
DFFARX1 I_66031 (I1126097,I3563,I1125707,I1126123,);
not I_66032 (I1126131,I1126123);
nor I_66033 (I1125693,I1126131,I1125936);
nand I_66034 (I1126162,I1126131,I1125781);
not I_66035 (I1126179,I1292386);
nand I_66036 (I1126196,I1126179,I1125885);
nand I_66037 (I1126213,I1126131,I1126196);
nand I_66038 (I1125684,I1126213,I1126162);
nand I_66039 (I1125681,I1126196,I1126080);
not I_66040 (I1126285,I3570);
DFFARX1 I_66041 (I991109,I3563,I1126285,I1126311,);
and I_66042 (I1126319,I1126311,I991103);
DFFARX1 I_66043 (I1126319,I3563,I1126285,I1126268,);
DFFARX1 I_66044 (I991121,I3563,I1126285,I1126359,);
not I_66045 (I1126367,I991112);
not I_66046 (I1126384,I991124);
nand I_66047 (I1126401,I1126384,I1126367);
nor I_66048 (I1126256,I1126359,I1126401);
DFFARX1 I_66049 (I1126401,I3563,I1126285,I1126441,);
not I_66050 (I1126277,I1126441);
not I_66051 (I1126463,I991130);
nand I_66052 (I1126480,I1126384,I1126463);
DFFARX1 I_66053 (I1126480,I3563,I1126285,I1126506,);
not I_66054 (I1126514,I1126506);
not I_66055 (I1126531,I991106);
nand I_66056 (I1126548,I1126531,I991127);
and I_66057 (I1126565,I1126367,I1126548);
nor I_66058 (I1126582,I1126480,I1126565);
DFFARX1 I_66059 (I1126582,I3563,I1126285,I1126253,);
DFFARX1 I_66060 (I1126565,I3563,I1126285,I1126274,);
nor I_66061 (I1126627,I991106,I991118);
nor I_66062 (I1126265,I1126480,I1126627);
or I_66063 (I1126658,I991106,I991118);
nor I_66064 (I1126675,I991103,I991115);
DFFARX1 I_66065 (I1126675,I3563,I1126285,I1126701,);
not I_66066 (I1126709,I1126701);
nor I_66067 (I1126271,I1126709,I1126514);
nand I_66068 (I1126740,I1126709,I1126359);
not I_66069 (I1126757,I991103);
nand I_66070 (I1126774,I1126757,I1126463);
nand I_66071 (I1126791,I1126709,I1126774);
nand I_66072 (I1126262,I1126791,I1126740);
nand I_66073 (I1126259,I1126774,I1126658);
not I_66074 (I1126863,I3570);
DFFARX1 I_66075 (I61414,I3563,I1126863,I1126889,);
and I_66076 (I1126897,I1126889,I61390);
DFFARX1 I_66077 (I1126897,I3563,I1126863,I1126846,);
DFFARX1 I_66078 (I61408,I3563,I1126863,I1126937,);
not I_66079 (I1126945,I61396);
not I_66080 (I1126962,I61393);
nand I_66081 (I1126979,I1126962,I1126945);
nor I_66082 (I1126834,I1126937,I1126979);
DFFARX1 I_66083 (I1126979,I3563,I1126863,I1127019,);
not I_66084 (I1126855,I1127019);
not I_66085 (I1127041,I61402);
nand I_66086 (I1127058,I1126962,I1127041);
DFFARX1 I_66087 (I1127058,I3563,I1126863,I1127084,);
not I_66088 (I1127092,I1127084);
not I_66089 (I1127109,I61393);
nand I_66090 (I1127126,I1127109,I61411);
and I_66091 (I1127143,I1126945,I1127126);
nor I_66092 (I1127160,I1127058,I1127143);
DFFARX1 I_66093 (I1127160,I3563,I1126863,I1126831,);
DFFARX1 I_66094 (I1127143,I3563,I1126863,I1126852,);
nor I_66095 (I1127205,I61393,I61405);
nor I_66096 (I1126843,I1127058,I1127205);
or I_66097 (I1127236,I61393,I61405);
nor I_66098 (I1127253,I61399,I61390);
DFFARX1 I_66099 (I1127253,I3563,I1126863,I1127279,);
not I_66100 (I1127287,I1127279);
nor I_66101 (I1126849,I1127287,I1127092);
nand I_66102 (I1127318,I1127287,I1126937);
not I_66103 (I1127335,I61399);
nand I_66104 (I1127352,I1127335,I1127041);
nand I_66105 (I1127369,I1127287,I1127352);
nand I_66106 (I1126840,I1127369,I1127318);
nand I_66107 (I1126837,I1127352,I1127236);
not I_66108 (I1127441,I3570);
DFFARX1 I_66109 (I620280,I3563,I1127441,I1127467,);
and I_66110 (I1127475,I1127467,I620268);
DFFARX1 I_66111 (I1127475,I3563,I1127441,I1127424,);
DFFARX1 I_66112 (I620283,I3563,I1127441,I1127515,);
not I_66113 (I1127523,I620274);
not I_66114 (I1127540,I620265);
nand I_66115 (I1127557,I1127540,I1127523);
nor I_66116 (I1127412,I1127515,I1127557);
DFFARX1 I_66117 (I1127557,I3563,I1127441,I1127597,);
not I_66118 (I1127433,I1127597);
not I_66119 (I1127619,I620271);
nand I_66120 (I1127636,I1127540,I1127619);
DFFARX1 I_66121 (I1127636,I3563,I1127441,I1127662,);
not I_66122 (I1127670,I1127662);
not I_66123 (I1127687,I620286);
nand I_66124 (I1127704,I1127687,I620289);
and I_66125 (I1127721,I1127523,I1127704);
nor I_66126 (I1127738,I1127636,I1127721);
DFFARX1 I_66127 (I1127738,I3563,I1127441,I1127409,);
DFFARX1 I_66128 (I1127721,I3563,I1127441,I1127430,);
nor I_66129 (I1127783,I620286,I620265);
nor I_66130 (I1127421,I1127636,I1127783);
or I_66131 (I1127814,I620286,I620265);
nor I_66132 (I1127831,I620277,I620268);
DFFARX1 I_66133 (I1127831,I3563,I1127441,I1127857,);
not I_66134 (I1127865,I1127857);
nor I_66135 (I1127427,I1127865,I1127670);
nand I_66136 (I1127896,I1127865,I1127515);
not I_66137 (I1127913,I620277);
nand I_66138 (I1127930,I1127913,I1127619);
nand I_66139 (I1127947,I1127865,I1127930);
nand I_66140 (I1127418,I1127947,I1127896);
nand I_66141 (I1127415,I1127930,I1127814);
not I_66142 (I1128019,I3570);
DFFARX1 I_66143 (I105682,I3563,I1128019,I1128045,);
and I_66144 (I1128053,I1128045,I105658);
DFFARX1 I_66145 (I1128053,I3563,I1128019,I1128002,);
DFFARX1 I_66146 (I105676,I3563,I1128019,I1128093,);
not I_66147 (I1128101,I105664);
not I_66148 (I1128118,I105661);
nand I_66149 (I1128135,I1128118,I1128101);
nor I_66150 (I1127990,I1128093,I1128135);
DFFARX1 I_66151 (I1128135,I3563,I1128019,I1128175,);
not I_66152 (I1128011,I1128175);
not I_66153 (I1128197,I105670);
nand I_66154 (I1128214,I1128118,I1128197);
DFFARX1 I_66155 (I1128214,I3563,I1128019,I1128240,);
not I_66156 (I1128248,I1128240);
not I_66157 (I1128265,I105661);
nand I_66158 (I1128282,I1128265,I105679);
and I_66159 (I1128299,I1128101,I1128282);
nor I_66160 (I1128316,I1128214,I1128299);
DFFARX1 I_66161 (I1128316,I3563,I1128019,I1127987,);
DFFARX1 I_66162 (I1128299,I3563,I1128019,I1128008,);
nor I_66163 (I1128361,I105661,I105673);
nor I_66164 (I1127999,I1128214,I1128361);
or I_66165 (I1128392,I105661,I105673);
nor I_66166 (I1128409,I105667,I105658);
DFFARX1 I_66167 (I1128409,I3563,I1128019,I1128435,);
not I_66168 (I1128443,I1128435);
nor I_66169 (I1128005,I1128443,I1128248);
nand I_66170 (I1128474,I1128443,I1128093);
not I_66171 (I1128491,I105667);
nand I_66172 (I1128508,I1128491,I1128197);
nand I_66173 (I1128525,I1128443,I1128508);
nand I_66174 (I1127996,I1128525,I1128474);
nand I_66175 (I1127993,I1128508,I1128392);
not I_66176 (I1128597,I3570);
DFFARX1 I_66177 (I475170,I3563,I1128597,I1128623,);
and I_66178 (I1128631,I1128623,I475185);
DFFARX1 I_66179 (I1128631,I3563,I1128597,I1128580,);
DFFARX1 I_66180 (I475188,I3563,I1128597,I1128671,);
not I_66181 (I1128679,I475182);
not I_66182 (I1128696,I475197);
nand I_66183 (I1128713,I1128696,I1128679);
nor I_66184 (I1128568,I1128671,I1128713);
DFFARX1 I_66185 (I1128713,I3563,I1128597,I1128753,);
not I_66186 (I1128589,I1128753);
not I_66187 (I1128775,I475173);
nand I_66188 (I1128792,I1128696,I1128775);
DFFARX1 I_66189 (I1128792,I3563,I1128597,I1128818,);
not I_66190 (I1128826,I1128818);
not I_66191 (I1128843,I475176);
nand I_66192 (I1128860,I1128843,I475170);
and I_66193 (I1128877,I1128679,I1128860);
nor I_66194 (I1128894,I1128792,I1128877);
DFFARX1 I_66195 (I1128894,I3563,I1128597,I1128565,);
DFFARX1 I_66196 (I1128877,I3563,I1128597,I1128586,);
nor I_66197 (I1128939,I475176,I475179);
nor I_66198 (I1128577,I1128792,I1128939);
or I_66199 (I1128970,I475176,I475179);
nor I_66200 (I1128987,I475194,I475191);
DFFARX1 I_66201 (I1128987,I3563,I1128597,I1129013,);
not I_66202 (I1129021,I1129013);
nor I_66203 (I1128583,I1129021,I1128826);
nand I_66204 (I1129052,I1129021,I1128671);
not I_66205 (I1129069,I475194);
nand I_66206 (I1129086,I1129069,I1128775);
nand I_66207 (I1129103,I1129021,I1129086);
nand I_66208 (I1128574,I1129103,I1129052);
nand I_66209 (I1128571,I1129086,I1128970);
not I_66210 (I1129175,I3570);
DFFARX1 I_66211 (I873245,I3563,I1129175,I1129201,);
and I_66212 (I1129209,I1129201,I873251);
DFFARX1 I_66213 (I1129209,I3563,I1129175,I1129158,);
DFFARX1 I_66214 (I873257,I3563,I1129175,I1129249,);
not I_66215 (I1129257,I873242);
not I_66216 (I1129274,I873242);
nand I_66217 (I1129291,I1129274,I1129257);
nor I_66218 (I1129146,I1129249,I1129291);
DFFARX1 I_66219 (I1129291,I3563,I1129175,I1129331,);
not I_66220 (I1129167,I1129331);
not I_66221 (I1129353,I873260);
nand I_66222 (I1129370,I1129274,I1129353);
DFFARX1 I_66223 (I1129370,I3563,I1129175,I1129396,);
not I_66224 (I1129404,I1129396);
not I_66225 (I1129421,I873254);
nand I_66226 (I1129438,I1129421,I873245);
and I_66227 (I1129455,I1129257,I1129438);
nor I_66228 (I1129472,I1129370,I1129455);
DFFARX1 I_66229 (I1129472,I3563,I1129175,I1129143,);
DFFARX1 I_66230 (I1129455,I3563,I1129175,I1129164,);
nor I_66231 (I1129517,I873254,I873263);
nor I_66232 (I1129155,I1129370,I1129517);
or I_66233 (I1129548,I873254,I873263);
nor I_66234 (I1129565,I873248,I873248);
DFFARX1 I_66235 (I1129565,I3563,I1129175,I1129591,);
not I_66236 (I1129599,I1129591);
nor I_66237 (I1129161,I1129599,I1129404);
nand I_66238 (I1129630,I1129599,I1129249);
not I_66239 (I1129647,I873248);
nand I_66240 (I1129664,I1129647,I1129353);
nand I_66241 (I1129681,I1129599,I1129664);
nand I_66242 (I1129152,I1129681,I1129630);
nand I_66243 (I1129149,I1129664,I1129548);
not I_66244 (I1129753,I3570);
DFFARX1 I_66245 (I512162,I3563,I1129753,I1129779,);
and I_66246 (I1129787,I1129779,I512177);
DFFARX1 I_66247 (I1129787,I3563,I1129753,I1129736,);
DFFARX1 I_66248 (I512180,I3563,I1129753,I1129827,);
not I_66249 (I1129835,I512174);
not I_66250 (I1129852,I512189);
nand I_66251 (I1129869,I1129852,I1129835);
nor I_66252 (I1129724,I1129827,I1129869);
DFFARX1 I_66253 (I1129869,I3563,I1129753,I1129909,);
not I_66254 (I1129745,I1129909);
not I_66255 (I1129931,I512165);
nand I_66256 (I1129948,I1129852,I1129931);
DFFARX1 I_66257 (I1129948,I3563,I1129753,I1129974,);
not I_66258 (I1129982,I1129974);
not I_66259 (I1129999,I512168);
nand I_66260 (I1130016,I1129999,I512162);
and I_66261 (I1130033,I1129835,I1130016);
nor I_66262 (I1130050,I1129948,I1130033);
DFFARX1 I_66263 (I1130050,I3563,I1129753,I1129721,);
DFFARX1 I_66264 (I1130033,I3563,I1129753,I1129742,);
nor I_66265 (I1130095,I512168,I512171);
nor I_66266 (I1129733,I1129948,I1130095);
or I_66267 (I1130126,I512168,I512171);
nor I_66268 (I1130143,I512186,I512183);
DFFARX1 I_66269 (I1130143,I3563,I1129753,I1130169,);
not I_66270 (I1130177,I1130169);
nor I_66271 (I1129739,I1130177,I1129982);
nand I_66272 (I1130208,I1130177,I1129827);
not I_66273 (I1130225,I512186);
nand I_66274 (I1130242,I1130225,I1129931);
nand I_66275 (I1130259,I1130177,I1130242);
nand I_66276 (I1129730,I1130259,I1130208);
nand I_66277 (I1129727,I1130242,I1130126);
not I_66278 (I1130331,I3570);
DFFARX1 I_66279 (I646290,I3563,I1130331,I1130357,);
and I_66280 (I1130365,I1130357,I646278);
DFFARX1 I_66281 (I1130365,I3563,I1130331,I1130314,);
DFFARX1 I_66282 (I646293,I3563,I1130331,I1130405,);
not I_66283 (I1130413,I646284);
not I_66284 (I1130430,I646275);
nand I_66285 (I1130447,I1130430,I1130413);
nor I_66286 (I1130302,I1130405,I1130447);
DFFARX1 I_66287 (I1130447,I3563,I1130331,I1130487,);
not I_66288 (I1130323,I1130487);
not I_66289 (I1130509,I646281);
nand I_66290 (I1130526,I1130430,I1130509);
DFFARX1 I_66291 (I1130526,I3563,I1130331,I1130552,);
not I_66292 (I1130560,I1130552);
not I_66293 (I1130577,I646296);
nand I_66294 (I1130594,I1130577,I646299);
and I_66295 (I1130611,I1130413,I1130594);
nor I_66296 (I1130628,I1130526,I1130611);
DFFARX1 I_66297 (I1130628,I3563,I1130331,I1130299,);
DFFARX1 I_66298 (I1130611,I3563,I1130331,I1130320,);
nor I_66299 (I1130673,I646296,I646275);
nor I_66300 (I1130311,I1130526,I1130673);
or I_66301 (I1130704,I646296,I646275);
nor I_66302 (I1130721,I646287,I646278);
DFFARX1 I_66303 (I1130721,I3563,I1130331,I1130747,);
not I_66304 (I1130755,I1130747);
nor I_66305 (I1130317,I1130755,I1130560);
nand I_66306 (I1130786,I1130755,I1130405);
not I_66307 (I1130803,I646287);
nand I_66308 (I1130820,I1130803,I1130509);
nand I_66309 (I1130837,I1130755,I1130820);
nand I_66310 (I1130308,I1130837,I1130786);
nand I_66311 (I1130305,I1130820,I1130704);
not I_66312 (I1130909,I3570);
DFFARX1 I_66313 (I593114,I3563,I1130909,I1130935,);
and I_66314 (I1130943,I1130935,I593102);
DFFARX1 I_66315 (I1130943,I3563,I1130909,I1130892,);
DFFARX1 I_66316 (I593117,I3563,I1130909,I1130983,);
not I_66317 (I1130991,I593108);
not I_66318 (I1131008,I593099);
nand I_66319 (I1131025,I1131008,I1130991);
nor I_66320 (I1130880,I1130983,I1131025);
DFFARX1 I_66321 (I1131025,I3563,I1130909,I1131065,);
not I_66322 (I1130901,I1131065);
not I_66323 (I1131087,I593105);
nand I_66324 (I1131104,I1131008,I1131087);
DFFARX1 I_66325 (I1131104,I3563,I1130909,I1131130,);
not I_66326 (I1131138,I1131130);
not I_66327 (I1131155,I593120);
nand I_66328 (I1131172,I1131155,I593123);
and I_66329 (I1131189,I1130991,I1131172);
nor I_66330 (I1131206,I1131104,I1131189);
DFFARX1 I_66331 (I1131206,I3563,I1130909,I1130877,);
DFFARX1 I_66332 (I1131189,I3563,I1130909,I1130898,);
nor I_66333 (I1131251,I593120,I593099);
nor I_66334 (I1130889,I1131104,I1131251);
or I_66335 (I1131282,I593120,I593099);
nor I_66336 (I1131299,I593111,I593102);
DFFARX1 I_66337 (I1131299,I3563,I1130909,I1131325,);
not I_66338 (I1131333,I1131325);
nor I_66339 (I1130895,I1131333,I1131138);
nand I_66340 (I1131364,I1131333,I1130983);
not I_66341 (I1131381,I593111);
nand I_66342 (I1131398,I1131381,I1131087);
nand I_66343 (I1131415,I1131333,I1131398);
nand I_66344 (I1130886,I1131415,I1131364);
nand I_66345 (I1130883,I1131398,I1131282);
not I_66346 (I1131487,I3570);
DFFARX1 I_66347 (I436002,I3563,I1131487,I1131513,);
and I_66348 (I1131521,I1131513,I436017);
DFFARX1 I_66349 (I1131521,I3563,I1131487,I1131470,);
DFFARX1 I_66350 (I436020,I3563,I1131487,I1131561,);
not I_66351 (I1131569,I436014);
not I_66352 (I1131586,I436029);
nand I_66353 (I1131603,I1131586,I1131569);
nor I_66354 (I1131458,I1131561,I1131603);
DFFARX1 I_66355 (I1131603,I3563,I1131487,I1131643,);
not I_66356 (I1131479,I1131643);
not I_66357 (I1131665,I436005);
nand I_66358 (I1131682,I1131586,I1131665);
DFFARX1 I_66359 (I1131682,I3563,I1131487,I1131708,);
not I_66360 (I1131716,I1131708);
not I_66361 (I1131733,I436008);
nand I_66362 (I1131750,I1131733,I436002);
and I_66363 (I1131767,I1131569,I1131750);
nor I_66364 (I1131784,I1131682,I1131767);
DFFARX1 I_66365 (I1131784,I3563,I1131487,I1131455,);
DFFARX1 I_66366 (I1131767,I3563,I1131487,I1131476,);
nor I_66367 (I1131829,I436008,I436011);
nor I_66368 (I1131467,I1131682,I1131829);
or I_66369 (I1131860,I436008,I436011);
nor I_66370 (I1131877,I436026,I436023);
DFFARX1 I_66371 (I1131877,I3563,I1131487,I1131903,);
not I_66372 (I1131911,I1131903);
nor I_66373 (I1131473,I1131911,I1131716);
nand I_66374 (I1131942,I1131911,I1131561);
not I_66375 (I1131959,I436026);
nand I_66376 (I1131976,I1131959,I1131665);
nand I_66377 (I1131993,I1131911,I1131976);
nand I_66378 (I1131464,I1131993,I1131942);
nand I_66379 (I1131461,I1131976,I1131860);
not I_66380 (I1132065,I3570);
DFFARX1 I_66381 (I573909,I3563,I1132065,I1132091,);
and I_66382 (I1132099,I1132091,I573924);
DFFARX1 I_66383 (I1132099,I3563,I1132065,I1132048,);
DFFARX1 I_66384 (I573915,I3563,I1132065,I1132139,);
not I_66385 (I1132147,I573909);
not I_66386 (I1132164,I573927);
nand I_66387 (I1132181,I1132164,I1132147);
nor I_66388 (I1132036,I1132139,I1132181);
DFFARX1 I_66389 (I1132181,I3563,I1132065,I1132221,);
not I_66390 (I1132057,I1132221);
not I_66391 (I1132243,I573918);
nand I_66392 (I1132260,I1132164,I1132243);
DFFARX1 I_66393 (I1132260,I3563,I1132065,I1132286,);
not I_66394 (I1132294,I1132286);
not I_66395 (I1132311,I573930);
nand I_66396 (I1132328,I1132311,I573906);
and I_66397 (I1132345,I1132147,I1132328);
nor I_66398 (I1132362,I1132260,I1132345);
DFFARX1 I_66399 (I1132362,I3563,I1132065,I1132033,);
DFFARX1 I_66400 (I1132345,I3563,I1132065,I1132054,);
nor I_66401 (I1132407,I573930,I573906);
nor I_66402 (I1132045,I1132260,I1132407);
or I_66403 (I1132438,I573930,I573906);
nor I_66404 (I1132455,I573912,I573921);
DFFARX1 I_66405 (I1132455,I3563,I1132065,I1132481,);
not I_66406 (I1132489,I1132481);
nor I_66407 (I1132051,I1132489,I1132294);
nand I_66408 (I1132520,I1132489,I1132139);
not I_66409 (I1132537,I573912);
nand I_66410 (I1132554,I1132537,I1132243);
nand I_66411 (I1132571,I1132489,I1132554);
nand I_66412 (I1132042,I1132571,I1132520);
nand I_66413 (I1132039,I1132554,I1132438);
not I_66414 (I1132643,I3570);
DFFARX1 I_66415 (I621436,I3563,I1132643,I1132669,);
and I_66416 (I1132677,I1132669,I621424);
DFFARX1 I_66417 (I1132677,I3563,I1132643,I1132626,);
DFFARX1 I_66418 (I621439,I3563,I1132643,I1132717,);
not I_66419 (I1132725,I621430);
not I_66420 (I1132742,I621421);
nand I_66421 (I1132759,I1132742,I1132725);
nor I_66422 (I1132614,I1132717,I1132759);
DFFARX1 I_66423 (I1132759,I3563,I1132643,I1132799,);
not I_66424 (I1132635,I1132799);
not I_66425 (I1132821,I621427);
nand I_66426 (I1132838,I1132742,I1132821);
DFFARX1 I_66427 (I1132838,I3563,I1132643,I1132864,);
not I_66428 (I1132872,I1132864);
not I_66429 (I1132889,I621442);
nand I_66430 (I1132906,I1132889,I621445);
and I_66431 (I1132923,I1132725,I1132906);
nor I_66432 (I1132940,I1132838,I1132923);
DFFARX1 I_66433 (I1132940,I3563,I1132643,I1132611,);
DFFARX1 I_66434 (I1132923,I3563,I1132643,I1132632,);
nor I_66435 (I1132985,I621442,I621421);
nor I_66436 (I1132623,I1132838,I1132985);
or I_66437 (I1133016,I621442,I621421);
nor I_66438 (I1133033,I621433,I621424);
DFFARX1 I_66439 (I1133033,I3563,I1132643,I1133059,);
not I_66440 (I1133067,I1133059);
nor I_66441 (I1132629,I1133067,I1132872);
nand I_66442 (I1133098,I1133067,I1132717);
not I_66443 (I1133115,I621433);
nand I_66444 (I1133132,I1133115,I1132821);
nand I_66445 (I1133149,I1133067,I1133132);
nand I_66446 (I1132620,I1133149,I1133098);
nand I_66447 (I1132617,I1133132,I1133016);
not I_66448 (I1133221,I3570);
DFFARX1 I_66449 (I123600,I3563,I1133221,I1133247,);
and I_66450 (I1133255,I1133247,I123576);
DFFARX1 I_66451 (I1133255,I3563,I1133221,I1133204,);
DFFARX1 I_66452 (I123594,I3563,I1133221,I1133295,);
not I_66453 (I1133303,I123582);
not I_66454 (I1133320,I123579);
nand I_66455 (I1133337,I1133320,I1133303);
nor I_66456 (I1133192,I1133295,I1133337);
DFFARX1 I_66457 (I1133337,I3563,I1133221,I1133377,);
not I_66458 (I1133213,I1133377);
not I_66459 (I1133399,I123588);
nand I_66460 (I1133416,I1133320,I1133399);
DFFARX1 I_66461 (I1133416,I3563,I1133221,I1133442,);
not I_66462 (I1133450,I1133442);
not I_66463 (I1133467,I123579);
nand I_66464 (I1133484,I1133467,I123597);
and I_66465 (I1133501,I1133303,I1133484);
nor I_66466 (I1133518,I1133416,I1133501);
DFFARX1 I_66467 (I1133518,I3563,I1133221,I1133189,);
DFFARX1 I_66468 (I1133501,I3563,I1133221,I1133210,);
nor I_66469 (I1133563,I123579,I123591);
nor I_66470 (I1133201,I1133416,I1133563);
or I_66471 (I1133594,I123579,I123591);
nor I_66472 (I1133611,I123585,I123576);
DFFARX1 I_66473 (I1133611,I3563,I1133221,I1133637,);
not I_66474 (I1133645,I1133637);
nor I_66475 (I1133207,I1133645,I1133450);
nand I_66476 (I1133676,I1133645,I1133295);
not I_66477 (I1133693,I123585);
nand I_66478 (I1133710,I1133693,I1133399);
nand I_66479 (I1133727,I1133645,I1133710);
nand I_66480 (I1133198,I1133727,I1133676);
nand I_66481 (I1133195,I1133710,I1133594);
not I_66482 (I1133799,I3570);
DFFARX1 I_66483 (I737036,I3563,I1133799,I1133825,);
and I_66484 (I1133833,I1133825,I737024);
DFFARX1 I_66485 (I1133833,I3563,I1133799,I1133782,);
DFFARX1 I_66486 (I737027,I3563,I1133799,I1133873,);
not I_66487 (I1133881,I737021);
not I_66488 (I1133898,I737045);
nand I_66489 (I1133915,I1133898,I1133881);
nor I_66490 (I1133770,I1133873,I1133915);
DFFARX1 I_66491 (I1133915,I3563,I1133799,I1133955,);
not I_66492 (I1133791,I1133955);
not I_66493 (I1133977,I737033);
nand I_66494 (I1133994,I1133898,I1133977);
DFFARX1 I_66495 (I1133994,I3563,I1133799,I1134020,);
not I_66496 (I1134028,I1134020);
not I_66497 (I1134045,I737042);
nand I_66498 (I1134062,I1134045,I737039);
and I_66499 (I1134079,I1133881,I1134062);
nor I_66500 (I1134096,I1133994,I1134079);
DFFARX1 I_66501 (I1134096,I3563,I1133799,I1133767,);
DFFARX1 I_66502 (I1134079,I3563,I1133799,I1133788,);
nor I_66503 (I1134141,I737042,I737030);
nor I_66504 (I1133779,I1133994,I1134141);
or I_66505 (I1134172,I737042,I737030);
nor I_66506 (I1134189,I737021,I737024);
DFFARX1 I_66507 (I1134189,I3563,I1133799,I1134215,);
not I_66508 (I1134223,I1134215);
nor I_66509 (I1133785,I1134223,I1134028);
nand I_66510 (I1134254,I1134223,I1133873);
not I_66511 (I1134271,I737021);
nand I_66512 (I1134288,I1134271,I1133977);
nand I_66513 (I1134305,I1134223,I1134288);
nand I_66514 (I1133776,I1134305,I1134254);
nand I_66515 (I1133773,I1134288,I1134172);
not I_66516 (I1134377,I3570);
DFFARX1 I_66517 (I169663,I3563,I1134377,I1134403,);
and I_66518 (I1134411,I1134403,I169666);
DFFARX1 I_66519 (I1134411,I3563,I1134377,I1134360,);
DFFARX1 I_66520 (I169666,I3563,I1134377,I1134451,);
not I_66521 (I1134459,I169681);
not I_66522 (I1134476,I169687);
nand I_66523 (I1134493,I1134476,I1134459);
nor I_66524 (I1134348,I1134451,I1134493);
DFFARX1 I_66525 (I1134493,I3563,I1134377,I1134533,);
not I_66526 (I1134369,I1134533);
not I_66527 (I1134555,I169675);
nand I_66528 (I1134572,I1134476,I1134555);
DFFARX1 I_66529 (I1134572,I3563,I1134377,I1134598,);
not I_66530 (I1134606,I1134598);
not I_66531 (I1134623,I169672);
nand I_66532 (I1134640,I1134623,I169669);
and I_66533 (I1134657,I1134459,I1134640);
nor I_66534 (I1134674,I1134572,I1134657);
DFFARX1 I_66535 (I1134674,I3563,I1134377,I1134345,);
DFFARX1 I_66536 (I1134657,I3563,I1134377,I1134366,);
nor I_66537 (I1134719,I169672,I169663);
nor I_66538 (I1134357,I1134572,I1134719);
or I_66539 (I1134750,I169672,I169663);
nor I_66540 (I1134767,I169678,I169684);
DFFARX1 I_66541 (I1134767,I3563,I1134377,I1134793,);
not I_66542 (I1134801,I1134793);
nor I_66543 (I1134363,I1134801,I1134606);
nand I_66544 (I1134832,I1134801,I1134451);
not I_66545 (I1134849,I169678);
nand I_66546 (I1134866,I1134849,I1134555);
nand I_66547 (I1134883,I1134801,I1134866);
nand I_66548 (I1134354,I1134883,I1134832);
nand I_66549 (I1134351,I1134866,I1134750);
not I_66550 (I1134955,I3570);
DFFARX1 I_66551 (I816329,I3563,I1134955,I1134981,);
and I_66552 (I1134989,I1134981,I816335);
DFFARX1 I_66553 (I1134989,I3563,I1134955,I1134938,);
DFFARX1 I_66554 (I816341,I3563,I1134955,I1135029,);
not I_66555 (I1135037,I816326);
not I_66556 (I1135054,I816326);
nand I_66557 (I1135071,I1135054,I1135037);
nor I_66558 (I1134926,I1135029,I1135071);
DFFARX1 I_66559 (I1135071,I3563,I1134955,I1135111,);
not I_66560 (I1134947,I1135111);
not I_66561 (I1135133,I816344);
nand I_66562 (I1135150,I1135054,I1135133);
DFFARX1 I_66563 (I1135150,I3563,I1134955,I1135176,);
not I_66564 (I1135184,I1135176);
not I_66565 (I1135201,I816338);
nand I_66566 (I1135218,I1135201,I816329);
and I_66567 (I1135235,I1135037,I1135218);
nor I_66568 (I1135252,I1135150,I1135235);
DFFARX1 I_66569 (I1135252,I3563,I1134955,I1134923,);
DFFARX1 I_66570 (I1135235,I3563,I1134955,I1134944,);
nor I_66571 (I1135297,I816338,I816347);
nor I_66572 (I1134935,I1135150,I1135297);
or I_66573 (I1135328,I816338,I816347);
nor I_66574 (I1135345,I816332,I816332);
DFFARX1 I_66575 (I1135345,I3563,I1134955,I1135371,);
not I_66576 (I1135379,I1135371);
nor I_66577 (I1134941,I1135379,I1135184);
nand I_66578 (I1135410,I1135379,I1135029);
not I_66579 (I1135427,I816332);
nand I_66580 (I1135444,I1135427,I1135133);
nand I_66581 (I1135461,I1135379,I1135444);
nand I_66582 (I1134932,I1135461,I1135410);
nand I_66583 (I1134929,I1135444,I1135328);
not I_66584 (I1135533,I3570);
DFFARX1 I_66585 (I194653,I3563,I1135533,I1135559,);
and I_66586 (I1135567,I1135559,I194656);
DFFARX1 I_66587 (I1135567,I3563,I1135533,I1135516,);
DFFARX1 I_66588 (I194656,I3563,I1135533,I1135607,);
not I_66589 (I1135615,I194671);
not I_66590 (I1135632,I194677);
nand I_66591 (I1135649,I1135632,I1135615);
nor I_66592 (I1135504,I1135607,I1135649);
DFFARX1 I_66593 (I1135649,I3563,I1135533,I1135689,);
not I_66594 (I1135525,I1135689);
not I_66595 (I1135711,I194665);
nand I_66596 (I1135728,I1135632,I1135711);
DFFARX1 I_66597 (I1135728,I3563,I1135533,I1135754,);
not I_66598 (I1135762,I1135754);
not I_66599 (I1135779,I194662);
nand I_66600 (I1135796,I1135779,I194659);
and I_66601 (I1135813,I1135615,I1135796);
nor I_66602 (I1135830,I1135728,I1135813);
DFFARX1 I_66603 (I1135830,I3563,I1135533,I1135501,);
DFFARX1 I_66604 (I1135813,I3563,I1135533,I1135522,);
nor I_66605 (I1135875,I194662,I194653);
nor I_66606 (I1135513,I1135728,I1135875);
or I_66607 (I1135906,I194662,I194653);
nor I_66608 (I1135923,I194668,I194674);
DFFARX1 I_66609 (I1135923,I3563,I1135533,I1135949,);
not I_66610 (I1135957,I1135949);
nor I_66611 (I1135519,I1135957,I1135762);
nand I_66612 (I1135988,I1135957,I1135607);
not I_66613 (I1136005,I194668);
nand I_66614 (I1136022,I1136005,I1135711);
nand I_66615 (I1136039,I1135957,I1136022);
nand I_66616 (I1135510,I1136039,I1135988);
nand I_66617 (I1135507,I1136022,I1135906);
not I_66618 (I1136111,I3570);
DFFARX1 I_66619 (I630684,I3563,I1136111,I1136137,);
and I_66620 (I1136145,I1136137,I630672);
DFFARX1 I_66621 (I1136145,I3563,I1136111,I1136094,);
DFFARX1 I_66622 (I630687,I3563,I1136111,I1136185,);
not I_66623 (I1136193,I630678);
not I_66624 (I1136210,I630669);
nand I_66625 (I1136227,I1136210,I1136193);
nor I_66626 (I1136082,I1136185,I1136227);
DFFARX1 I_66627 (I1136227,I3563,I1136111,I1136267,);
not I_66628 (I1136103,I1136267);
not I_66629 (I1136289,I630675);
nand I_66630 (I1136306,I1136210,I1136289);
DFFARX1 I_66631 (I1136306,I3563,I1136111,I1136332,);
not I_66632 (I1136340,I1136332);
not I_66633 (I1136357,I630690);
nand I_66634 (I1136374,I1136357,I630693);
and I_66635 (I1136391,I1136193,I1136374);
nor I_66636 (I1136408,I1136306,I1136391);
DFFARX1 I_66637 (I1136408,I3563,I1136111,I1136079,);
DFFARX1 I_66638 (I1136391,I3563,I1136111,I1136100,);
nor I_66639 (I1136453,I630690,I630669);
nor I_66640 (I1136091,I1136306,I1136453);
or I_66641 (I1136484,I630690,I630669);
nor I_66642 (I1136501,I630681,I630672);
DFFARX1 I_66643 (I1136501,I3563,I1136111,I1136527,);
not I_66644 (I1136535,I1136527);
nor I_66645 (I1136097,I1136535,I1136340);
nand I_66646 (I1136566,I1136535,I1136185);
not I_66647 (I1136583,I630681);
nand I_66648 (I1136600,I1136583,I1136289);
nand I_66649 (I1136617,I1136535,I1136600);
nand I_66650 (I1136088,I1136617,I1136566);
nand I_66651 (I1136085,I1136600,I1136484);
not I_66652 (I1136689,I3570);
DFFARX1 I_66653 (I115168,I3563,I1136689,I1136715,);
and I_66654 (I1136723,I1136715,I115144);
DFFARX1 I_66655 (I1136723,I3563,I1136689,I1136672,);
DFFARX1 I_66656 (I115162,I3563,I1136689,I1136763,);
not I_66657 (I1136771,I115150);
not I_66658 (I1136788,I115147);
nand I_66659 (I1136805,I1136788,I1136771);
nor I_66660 (I1136660,I1136763,I1136805);
DFFARX1 I_66661 (I1136805,I3563,I1136689,I1136845,);
not I_66662 (I1136681,I1136845);
not I_66663 (I1136867,I115156);
nand I_66664 (I1136884,I1136788,I1136867);
DFFARX1 I_66665 (I1136884,I3563,I1136689,I1136910,);
not I_66666 (I1136918,I1136910);
not I_66667 (I1136935,I115147);
nand I_66668 (I1136952,I1136935,I115165);
and I_66669 (I1136969,I1136771,I1136952);
nor I_66670 (I1136986,I1136884,I1136969);
DFFARX1 I_66671 (I1136986,I3563,I1136689,I1136657,);
DFFARX1 I_66672 (I1136969,I3563,I1136689,I1136678,);
nor I_66673 (I1137031,I115147,I115159);
nor I_66674 (I1136669,I1136884,I1137031);
or I_66675 (I1137062,I115147,I115159);
nor I_66676 (I1137079,I115153,I115144);
DFFARX1 I_66677 (I1137079,I3563,I1136689,I1137105,);
not I_66678 (I1137113,I1137105);
nor I_66679 (I1136675,I1137113,I1136918);
nand I_66680 (I1137144,I1137113,I1136763);
not I_66681 (I1137161,I115153);
nand I_66682 (I1137178,I1137161,I1136867);
nand I_66683 (I1137195,I1137113,I1137178);
nand I_66684 (I1136666,I1137195,I1137144);
nand I_66685 (I1136663,I1137178,I1137062);
not I_66686 (I1137267,I3570);
DFFARX1 I_66687 (I557844,I3563,I1137267,I1137293,);
and I_66688 (I1137301,I1137293,I557859);
DFFARX1 I_66689 (I1137301,I3563,I1137267,I1137250,);
DFFARX1 I_66690 (I557850,I3563,I1137267,I1137341,);
not I_66691 (I1137349,I557844);
not I_66692 (I1137366,I557862);
nand I_66693 (I1137383,I1137366,I1137349);
nor I_66694 (I1137238,I1137341,I1137383);
DFFARX1 I_66695 (I1137383,I3563,I1137267,I1137423,);
not I_66696 (I1137259,I1137423);
not I_66697 (I1137445,I557853);
nand I_66698 (I1137462,I1137366,I1137445);
DFFARX1 I_66699 (I1137462,I3563,I1137267,I1137488,);
not I_66700 (I1137496,I1137488);
not I_66701 (I1137513,I557865);
nand I_66702 (I1137530,I1137513,I557841);
and I_66703 (I1137547,I1137349,I1137530);
nor I_66704 (I1137564,I1137462,I1137547);
DFFARX1 I_66705 (I1137564,I3563,I1137267,I1137235,);
DFFARX1 I_66706 (I1137547,I3563,I1137267,I1137256,);
nor I_66707 (I1137609,I557865,I557841);
nor I_66708 (I1137247,I1137462,I1137609);
or I_66709 (I1137640,I557865,I557841);
nor I_66710 (I1137657,I557847,I557856);
DFFARX1 I_66711 (I1137657,I3563,I1137267,I1137683,);
not I_66712 (I1137691,I1137683);
nor I_66713 (I1137253,I1137691,I1137496);
nand I_66714 (I1137722,I1137691,I1137341);
not I_66715 (I1137739,I557847);
nand I_66716 (I1137756,I1137739,I1137445);
nand I_66717 (I1137773,I1137691,I1137756);
nand I_66718 (I1137244,I1137773,I1137722);
nand I_66719 (I1137241,I1137756,I1137640);
not I_66720 (I1137845,I3570);
DFFARX1 I_66721 (I251178,I3563,I1137845,I1137871,);
and I_66722 (I1137879,I1137871,I251181);
DFFARX1 I_66723 (I1137879,I3563,I1137845,I1137828,);
DFFARX1 I_66724 (I251181,I3563,I1137845,I1137919,);
not I_66725 (I1137927,I251196);
not I_66726 (I1137944,I251202);
nand I_66727 (I1137961,I1137944,I1137927);
nor I_66728 (I1137816,I1137919,I1137961);
DFFARX1 I_66729 (I1137961,I3563,I1137845,I1138001,);
not I_66730 (I1137837,I1138001);
not I_66731 (I1138023,I251190);
nand I_66732 (I1138040,I1137944,I1138023);
DFFARX1 I_66733 (I1138040,I3563,I1137845,I1138066,);
not I_66734 (I1138074,I1138066);
not I_66735 (I1138091,I251187);
nand I_66736 (I1138108,I1138091,I251184);
and I_66737 (I1138125,I1137927,I1138108);
nor I_66738 (I1138142,I1138040,I1138125);
DFFARX1 I_66739 (I1138142,I3563,I1137845,I1137813,);
DFFARX1 I_66740 (I1138125,I3563,I1137845,I1137834,);
nor I_66741 (I1138187,I251187,I251178);
nor I_66742 (I1137825,I1138040,I1138187);
or I_66743 (I1138218,I251187,I251178);
nor I_66744 (I1138235,I251193,I251199);
DFFARX1 I_66745 (I1138235,I3563,I1137845,I1138261,);
not I_66746 (I1138269,I1138261);
nor I_66747 (I1137831,I1138269,I1138074);
nand I_66748 (I1138300,I1138269,I1137919);
not I_66749 (I1138317,I251193);
nand I_66750 (I1138334,I1138317,I1138023);
nand I_66751 (I1138351,I1138269,I1138334);
nand I_66752 (I1137822,I1138351,I1138300);
nand I_66753 (I1137819,I1138334,I1138218);
not I_66754 (I1138423,I3570);
DFFARX1 I_66755 (I882731,I3563,I1138423,I1138449,);
and I_66756 (I1138457,I1138449,I882737);
DFFARX1 I_66757 (I1138457,I3563,I1138423,I1138406,);
DFFARX1 I_66758 (I882743,I3563,I1138423,I1138497,);
not I_66759 (I1138505,I882728);
not I_66760 (I1138522,I882728);
nand I_66761 (I1138539,I1138522,I1138505);
nor I_66762 (I1138394,I1138497,I1138539);
DFFARX1 I_66763 (I1138539,I3563,I1138423,I1138579,);
not I_66764 (I1138415,I1138579);
not I_66765 (I1138601,I882746);
nand I_66766 (I1138618,I1138522,I1138601);
DFFARX1 I_66767 (I1138618,I3563,I1138423,I1138644,);
not I_66768 (I1138652,I1138644);
not I_66769 (I1138669,I882740);
nand I_66770 (I1138686,I1138669,I882731);
and I_66771 (I1138703,I1138505,I1138686);
nor I_66772 (I1138720,I1138618,I1138703);
DFFARX1 I_66773 (I1138720,I3563,I1138423,I1138391,);
DFFARX1 I_66774 (I1138703,I3563,I1138423,I1138412,);
nor I_66775 (I1138765,I882740,I882749);
nor I_66776 (I1138403,I1138618,I1138765);
or I_66777 (I1138796,I882740,I882749);
nor I_66778 (I1138813,I882734,I882734);
DFFARX1 I_66779 (I1138813,I3563,I1138423,I1138839,);
not I_66780 (I1138847,I1138839);
nor I_66781 (I1138409,I1138847,I1138652);
nand I_66782 (I1138878,I1138847,I1138497);
not I_66783 (I1138895,I882734);
nand I_66784 (I1138912,I1138895,I1138601);
nand I_66785 (I1138929,I1138847,I1138912);
nand I_66786 (I1138400,I1138929,I1138878);
nand I_66787 (I1138397,I1138912,I1138796);
not I_66788 (I1139001,I3570);
DFFARX1 I_66789 (I446338,I3563,I1139001,I1139027,);
and I_66790 (I1139035,I1139027,I446353);
DFFARX1 I_66791 (I1139035,I3563,I1139001,I1138984,);
DFFARX1 I_66792 (I446356,I3563,I1139001,I1139075,);
not I_66793 (I1139083,I446350);
not I_66794 (I1139100,I446365);
nand I_66795 (I1139117,I1139100,I1139083);
nor I_66796 (I1138972,I1139075,I1139117);
DFFARX1 I_66797 (I1139117,I3563,I1139001,I1139157,);
not I_66798 (I1138993,I1139157);
not I_66799 (I1139179,I446341);
nand I_66800 (I1139196,I1139100,I1139179);
DFFARX1 I_66801 (I1139196,I3563,I1139001,I1139222,);
not I_66802 (I1139230,I1139222);
not I_66803 (I1139247,I446344);
nand I_66804 (I1139264,I1139247,I446338);
and I_66805 (I1139281,I1139083,I1139264);
nor I_66806 (I1139298,I1139196,I1139281);
DFFARX1 I_66807 (I1139298,I3563,I1139001,I1138969,);
DFFARX1 I_66808 (I1139281,I3563,I1139001,I1138990,);
nor I_66809 (I1139343,I446344,I446347);
nor I_66810 (I1138981,I1139196,I1139343);
or I_66811 (I1139374,I446344,I446347);
nor I_66812 (I1139391,I446362,I446359);
DFFARX1 I_66813 (I1139391,I3563,I1139001,I1139417,);
not I_66814 (I1139425,I1139417);
nor I_66815 (I1138987,I1139425,I1139230);
nand I_66816 (I1139456,I1139425,I1139075);
not I_66817 (I1139473,I446362);
nand I_66818 (I1139490,I1139473,I1139179);
nand I_66819 (I1139507,I1139425,I1139490);
nand I_66820 (I1138978,I1139507,I1139456);
nand I_66821 (I1138975,I1139490,I1139374);
not I_66822 (I1139579,I3570);
DFFARX1 I_66823 (I1407120,I3563,I1139579,I1139605,);
and I_66824 (I1139613,I1139605,I1407102);
DFFARX1 I_66825 (I1139613,I3563,I1139579,I1139562,);
DFFARX1 I_66826 (I1407093,I3563,I1139579,I1139653,);
not I_66827 (I1139661,I1407108);
not I_66828 (I1139678,I1407096);
nand I_66829 (I1139695,I1139678,I1139661);
nor I_66830 (I1139550,I1139653,I1139695);
DFFARX1 I_66831 (I1139695,I3563,I1139579,I1139735,);
not I_66832 (I1139571,I1139735);
not I_66833 (I1139757,I1407105);
nand I_66834 (I1139774,I1139678,I1139757);
DFFARX1 I_66835 (I1139774,I3563,I1139579,I1139800,);
not I_66836 (I1139808,I1139800);
not I_66837 (I1139825,I1407114);
nand I_66838 (I1139842,I1139825,I1407093);
and I_66839 (I1139859,I1139661,I1139842);
nor I_66840 (I1139876,I1139774,I1139859);
DFFARX1 I_66841 (I1139876,I3563,I1139579,I1139547,);
DFFARX1 I_66842 (I1139859,I3563,I1139579,I1139568,);
nor I_66843 (I1139921,I1407114,I1407117);
nor I_66844 (I1139559,I1139774,I1139921);
or I_66845 (I1139952,I1407114,I1407117);
nor I_66846 (I1139969,I1407111,I1407099);
DFFARX1 I_66847 (I1139969,I3563,I1139579,I1139995,);
not I_66848 (I1140003,I1139995);
nor I_66849 (I1139565,I1140003,I1139808);
nand I_66850 (I1140034,I1140003,I1139653);
not I_66851 (I1140051,I1407111);
nand I_66852 (I1140068,I1140051,I1139757);
nand I_66853 (I1140085,I1140003,I1140068);
nand I_66854 (I1139556,I1140085,I1140034);
nand I_66855 (I1139553,I1140068,I1139952);
not I_66856 (I1140157,I3570);
DFFARX1 I_66857 (I378671,I3563,I1140157,I1140183,);
and I_66858 (I1140191,I1140183,I378656);
DFFARX1 I_66859 (I1140191,I3563,I1140157,I1140140,);
DFFARX1 I_66860 (I378662,I3563,I1140157,I1140231,);
not I_66861 (I1140239,I378644);
not I_66862 (I1140256,I378665);
nand I_66863 (I1140273,I1140256,I1140239);
nor I_66864 (I1140128,I1140231,I1140273);
DFFARX1 I_66865 (I1140273,I3563,I1140157,I1140313,);
not I_66866 (I1140149,I1140313);
not I_66867 (I1140335,I378668);
nand I_66868 (I1140352,I1140256,I1140335);
DFFARX1 I_66869 (I1140352,I3563,I1140157,I1140378,);
not I_66870 (I1140386,I1140378);
not I_66871 (I1140403,I378659);
nand I_66872 (I1140420,I1140403,I378647);
and I_66873 (I1140437,I1140239,I1140420);
nor I_66874 (I1140454,I1140352,I1140437);
DFFARX1 I_66875 (I1140454,I3563,I1140157,I1140125,);
DFFARX1 I_66876 (I1140437,I3563,I1140157,I1140146,);
nor I_66877 (I1140499,I378659,I378653);
nor I_66878 (I1140137,I1140352,I1140499);
or I_66879 (I1140530,I378659,I378653);
nor I_66880 (I1140547,I378650,I378644);
DFFARX1 I_66881 (I1140547,I3563,I1140157,I1140573,);
not I_66882 (I1140581,I1140573);
nor I_66883 (I1140143,I1140581,I1140386);
nand I_66884 (I1140612,I1140581,I1140231);
not I_66885 (I1140629,I378650);
nand I_66886 (I1140646,I1140629,I1140335);
nand I_66887 (I1140663,I1140581,I1140646);
nand I_66888 (I1140134,I1140663,I1140612);
nand I_66889 (I1140131,I1140646,I1140530);
not I_66890 (I1140735,I3570);
DFFARX1 I_66891 (I654382,I3563,I1140735,I1140761,);
and I_66892 (I1140769,I1140761,I654370);
DFFARX1 I_66893 (I1140769,I3563,I1140735,I1140718,);
DFFARX1 I_66894 (I654385,I3563,I1140735,I1140809,);
not I_66895 (I1140817,I654376);
not I_66896 (I1140834,I654367);
nand I_66897 (I1140851,I1140834,I1140817);
nor I_66898 (I1140706,I1140809,I1140851);
DFFARX1 I_66899 (I1140851,I3563,I1140735,I1140891,);
not I_66900 (I1140727,I1140891);
not I_66901 (I1140913,I654373);
nand I_66902 (I1140930,I1140834,I1140913);
DFFARX1 I_66903 (I1140930,I3563,I1140735,I1140956,);
not I_66904 (I1140964,I1140956);
not I_66905 (I1140981,I654388);
nand I_66906 (I1140998,I1140981,I654391);
and I_66907 (I1141015,I1140817,I1140998);
nor I_66908 (I1141032,I1140930,I1141015);
DFFARX1 I_66909 (I1141032,I3563,I1140735,I1140703,);
DFFARX1 I_66910 (I1141015,I3563,I1140735,I1140724,);
nor I_66911 (I1141077,I654388,I654367);
nor I_66912 (I1140715,I1140930,I1141077);
or I_66913 (I1141108,I654388,I654367);
nor I_66914 (I1141125,I654379,I654370);
DFFARX1 I_66915 (I1141125,I3563,I1140735,I1141151,);
not I_66916 (I1141159,I1141151);
nor I_66917 (I1140721,I1141159,I1140964);
nand I_66918 (I1141190,I1141159,I1140809);
not I_66919 (I1141207,I654379);
nand I_66920 (I1141224,I1141207,I1140913);
nand I_66921 (I1141241,I1141159,I1141224);
nand I_66922 (I1140712,I1141241,I1141190);
nand I_66923 (I1140709,I1141224,I1141108);
not I_66924 (I1141313,I3570);
DFFARX1 I_66925 (I191083,I3563,I1141313,I1141339,);
and I_66926 (I1141347,I1141339,I191086);
DFFARX1 I_66927 (I1141347,I3563,I1141313,I1141296,);
DFFARX1 I_66928 (I191086,I3563,I1141313,I1141387,);
not I_66929 (I1141395,I191101);
not I_66930 (I1141412,I191107);
nand I_66931 (I1141429,I1141412,I1141395);
nor I_66932 (I1141284,I1141387,I1141429);
DFFARX1 I_66933 (I1141429,I3563,I1141313,I1141469,);
not I_66934 (I1141305,I1141469);
not I_66935 (I1141491,I191095);
nand I_66936 (I1141508,I1141412,I1141491);
DFFARX1 I_66937 (I1141508,I3563,I1141313,I1141534,);
not I_66938 (I1141542,I1141534);
not I_66939 (I1141559,I191092);
nand I_66940 (I1141576,I1141559,I191089);
and I_66941 (I1141593,I1141395,I1141576);
nor I_66942 (I1141610,I1141508,I1141593);
DFFARX1 I_66943 (I1141610,I3563,I1141313,I1141281,);
DFFARX1 I_66944 (I1141593,I3563,I1141313,I1141302,);
nor I_66945 (I1141655,I191092,I191083);
nor I_66946 (I1141293,I1141508,I1141655);
or I_66947 (I1141686,I191092,I191083);
nor I_66948 (I1141703,I191098,I191104);
DFFARX1 I_66949 (I1141703,I3563,I1141313,I1141729,);
not I_66950 (I1141737,I1141729);
nor I_66951 (I1141299,I1141737,I1141542);
nand I_66952 (I1141768,I1141737,I1141387);
not I_66953 (I1141785,I191098);
nand I_66954 (I1141802,I1141785,I1141491);
nand I_66955 (I1141819,I1141737,I1141802);
nand I_66956 (I1141290,I1141819,I1141768);
nand I_66957 (I1141287,I1141802,I1141686);
not I_66958 (I1141891,I3570);
DFFARX1 I_66959 (I852165,I3563,I1141891,I1141917,);
and I_66960 (I1141925,I1141917,I852171);
DFFARX1 I_66961 (I1141925,I3563,I1141891,I1141874,);
DFFARX1 I_66962 (I852177,I3563,I1141891,I1141965,);
not I_66963 (I1141973,I852162);
not I_66964 (I1141990,I852162);
nand I_66965 (I1142007,I1141990,I1141973);
nor I_66966 (I1141862,I1141965,I1142007);
DFFARX1 I_66967 (I1142007,I3563,I1141891,I1142047,);
not I_66968 (I1141883,I1142047);
not I_66969 (I1142069,I852180);
nand I_66970 (I1142086,I1141990,I1142069);
DFFARX1 I_66971 (I1142086,I3563,I1141891,I1142112,);
not I_66972 (I1142120,I1142112);
not I_66973 (I1142137,I852174);
nand I_66974 (I1142154,I1142137,I852165);
and I_66975 (I1142171,I1141973,I1142154);
nor I_66976 (I1142188,I1142086,I1142171);
DFFARX1 I_66977 (I1142188,I3563,I1141891,I1141859,);
DFFARX1 I_66978 (I1142171,I3563,I1141891,I1141880,);
nor I_66979 (I1142233,I852174,I852183);
nor I_66980 (I1141871,I1142086,I1142233);
or I_66981 (I1142264,I852174,I852183);
nor I_66982 (I1142281,I852168,I852168);
DFFARX1 I_66983 (I1142281,I3563,I1141891,I1142307,);
not I_66984 (I1142315,I1142307);
nor I_66985 (I1141877,I1142315,I1142120);
nand I_66986 (I1142346,I1142315,I1141965);
not I_66987 (I1142363,I852168);
nand I_66988 (I1142380,I1142363,I1142069);
nand I_66989 (I1142397,I1142315,I1142380);
nand I_66990 (I1141868,I1142397,I1142346);
nand I_66991 (I1141865,I1142380,I1142264);
not I_66992 (I1142469,I3570);
DFFARX1 I_66993 (I703512,I3563,I1142469,I1142495,);
and I_66994 (I1142503,I1142495,I703500);
DFFARX1 I_66995 (I1142503,I3563,I1142469,I1142452,);
DFFARX1 I_66996 (I703503,I3563,I1142469,I1142543,);
not I_66997 (I1142551,I703497);
not I_66998 (I1142568,I703521);
nand I_66999 (I1142585,I1142568,I1142551);
nor I_67000 (I1142440,I1142543,I1142585);
DFFARX1 I_67001 (I1142585,I3563,I1142469,I1142625,);
not I_67002 (I1142461,I1142625);
not I_67003 (I1142647,I703509);
nand I_67004 (I1142664,I1142568,I1142647);
DFFARX1 I_67005 (I1142664,I3563,I1142469,I1142690,);
not I_67006 (I1142698,I1142690);
not I_67007 (I1142715,I703518);
nand I_67008 (I1142732,I1142715,I703515);
and I_67009 (I1142749,I1142551,I1142732);
nor I_67010 (I1142766,I1142664,I1142749);
DFFARX1 I_67011 (I1142766,I3563,I1142469,I1142437,);
DFFARX1 I_67012 (I1142749,I3563,I1142469,I1142458,);
nor I_67013 (I1142811,I703518,I703506);
nor I_67014 (I1142449,I1142664,I1142811);
or I_67015 (I1142842,I703518,I703506);
nor I_67016 (I1142859,I703497,I703500);
DFFARX1 I_67017 (I1142859,I3563,I1142469,I1142885,);
not I_67018 (I1142893,I1142885);
nor I_67019 (I1142455,I1142893,I1142698);
nand I_67020 (I1142924,I1142893,I1142543);
not I_67021 (I1142941,I703497);
nand I_67022 (I1142958,I1142941,I1142647);
nand I_67023 (I1142975,I1142893,I1142958);
nand I_67024 (I1142446,I1142975,I1142924);
nand I_67025 (I1142443,I1142958,I1142842);
not I_67026 (I1143047,I3570);
DFFARX1 I_67027 (I238088,I3563,I1143047,I1143073,);
and I_67028 (I1143081,I1143073,I238091);
DFFARX1 I_67029 (I1143081,I3563,I1143047,I1143030,);
DFFARX1 I_67030 (I238091,I3563,I1143047,I1143121,);
not I_67031 (I1143129,I238106);
not I_67032 (I1143146,I238112);
nand I_67033 (I1143163,I1143146,I1143129);
nor I_67034 (I1143018,I1143121,I1143163);
DFFARX1 I_67035 (I1143163,I3563,I1143047,I1143203,);
not I_67036 (I1143039,I1143203);
not I_67037 (I1143225,I238100);
nand I_67038 (I1143242,I1143146,I1143225);
DFFARX1 I_67039 (I1143242,I3563,I1143047,I1143268,);
not I_67040 (I1143276,I1143268);
not I_67041 (I1143293,I238097);
nand I_67042 (I1143310,I1143293,I238094);
and I_67043 (I1143327,I1143129,I1143310);
nor I_67044 (I1143344,I1143242,I1143327);
DFFARX1 I_67045 (I1143344,I3563,I1143047,I1143015,);
DFFARX1 I_67046 (I1143327,I3563,I1143047,I1143036,);
nor I_67047 (I1143389,I238097,I238088);
nor I_67048 (I1143027,I1143242,I1143389);
or I_67049 (I1143420,I238097,I238088);
nor I_67050 (I1143437,I238103,I238109);
DFFARX1 I_67051 (I1143437,I3563,I1143047,I1143463,);
not I_67052 (I1143471,I1143463);
nor I_67053 (I1143033,I1143471,I1143276);
nand I_67054 (I1143502,I1143471,I1143121);
not I_67055 (I1143519,I238103);
nand I_67056 (I1143536,I1143519,I1143225);
nand I_67057 (I1143553,I1143471,I1143536);
nand I_67058 (I1143024,I1143553,I1143502);
nand I_67059 (I1143021,I1143536,I1143420);
not I_67060 (I1143625,I3570);
DFFARX1 I_67061 (I929739,I3563,I1143625,I1143651,);
and I_67062 (I1143659,I1143651,I929733);
DFFARX1 I_67063 (I1143659,I3563,I1143625,I1143608,);
DFFARX1 I_67064 (I929751,I3563,I1143625,I1143699,);
not I_67065 (I1143707,I929742);
not I_67066 (I1143724,I929754);
nand I_67067 (I1143741,I1143724,I1143707);
nor I_67068 (I1143596,I1143699,I1143741);
DFFARX1 I_67069 (I1143741,I3563,I1143625,I1143781,);
not I_67070 (I1143617,I1143781);
not I_67071 (I1143803,I929760);
nand I_67072 (I1143820,I1143724,I1143803);
DFFARX1 I_67073 (I1143820,I3563,I1143625,I1143846,);
not I_67074 (I1143854,I1143846);
not I_67075 (I1143871,I929736);
nand I_67076 (I1143888,I1143871,I929757);
and I_67077 (I1143905,I1143707,I1143888);
nor I_67078 (I1143922,I1143820,I1143905);
DFFARX1 I_67079 (I1143922,I3563,I1143625,I1143593,);
DFFARX1 I_67080 (I1143905,I3563,I1143625,I1143614,);
nor I_67081 (I1143967,I929736,I929748);
nor I_67082 (I1143605,I1143820,I1143967);
or I_67083 (I1143998,I929736,I929748);
nor I_67084 (I1144015,I929733,I929745);
DFFARX1 I_67085 (I1144015,I3563,I1143625,I1144041,);
not I_67086 (I1144049,I1144041);
nor I_67087 (I1143611,I1144049,I1143854);
nand I_67088 (I1144080,I1144049,I1143699);
not I_67089 (I1144097,I929733);
nand I_67090 (I1144114,I1144097,I1143803);
nand I_67091 (I1144131,I1144049,I1144114);
nand I_67092 (I1143602,I1144131,I1144080);
nand I_67093 (I1143599,I1144114,I1143998);
not I_67094 (I1144203,I3570);
DFFARX1 I_67095 (I627794,I3563,I1144203,I1144229,);
and I_67096 (I1144237,I1144229,I627782);
DFFARX1 I_67097 (I1144237,I3563,I1144203,I1144186,);
DFFARX1 I_67098 (I627797,I3563,I1144203,I1144277,);
not I_67099 (I1144285,I627788);
not I_67100 (I1144302,I627779);
nand I_67101 (I1144319,I1144302,I1144285);
nor I_67102 (I1144174,I1144277,I1144319);
DFFARX1 I_67103 (I1144319,I3563,I1144203,I1144359,);
not I_67104 (I1144195,I1144359);
not I_67105 (I1144381,I627785);
nand I_67106 (I1144398,I1144302,I1144381);
DFFARX1 I_67107 (I1144398,I3563,I1144203,I1144424,);
not I_67108 (I1144432,I1144424);
not I_67109 (I1144449,I627800);
nand I_67110 (I1144466,I1144449,I627803);
and I_67111 (I1144483,I1144285,I1144466);
nor I_67112 (I1144500,I1144398,I1144483);
DFFARX1 I_67113 (I1144500,I3563,I1144203,I1144171,);
DFFARX1 I_67114 (I1144483,I3563,I1144203,I1144192,);
nor I_67115 (I1144545,I627800,I627779);
nor I_67116 (I1144183,I1144398,I1144545);
or I_67117 (I1144576,I627800,I627779);
nor I_67118 (I1144593,I627791,I627782);
DFFARX1 I_67119 (I1144593,I3563,I1144203,I1144619,);
not I_67120 (I1144627,I1144619);
nor I_67121 (I1144189,I1144627,I1144432);
nand I_67122 (I1144658,I1144627,I1144277);
not I_67123 (I1144675,I627791);
nand I_67124 (I1144692,I1144675,I1144381);
nand I_67125 (I1144709,I1144627,I1144692);
nand I_67126 (I1144180,I1144709,I1144658);
nand I_67127 (I1144177,I1144692,I1144576);
not I_67128 (I1144781,I3570);
DFFARX1 I_67129 (I699466,I3563,I1144781,I1144807,);
and I_67130 (I1144815,I1144807,I699454);
DFFARX1 I_67131 (I1144815,I3563,I1144781,I1144764,);
DFFARX1 I_67132 (I699457,I3563,I1144781,I1144855,);
not I_67133 (I1144863,I699451);
not I_67134 (I1144880,I699475);
nand I_67135 (I1144897,I1144880,I1144863);
nor I_67136 (I1144752,I1144855,I1144897);
DFFARX1 I_67137 (I1144897,I3563,I1144781,I1144937,);
not I_67138 (I1144773,I1144937);
not I_67139 (I1144959,I699463);
nand I_67140 (I1144976,I1144880,I1144959);
DFFARX1 I_67141 (I1144976,I3563,I1144781,I1145002,);
not I_67142 (I1145010,I1145002);
not I_67143 (I1145027,I699472);
nand I_67144 (I1145044,I1145027,I699469);
and I_67145 (I1145061,I1144863,I1145044);
nor I_67146 (I1145078,I1144976,I1145061);
DFFARX1 I_67147 (I1145078,I3563,I1144781,I1144749,);
DFFARX1 I_67148 (I1145061,I3563,I1144781,I1144770,);
nor I_67149 (I1145123,I699472,I699460);
nor I_67150 (I1144761,I1144976,I1145123);
or I_67151 (I1145154,I699472,I699460);
nor I_67152 (I1145171,I699451,I699454);
DFFARX1 I_67153 (I1145171,I3563,I1144781,I1145197,);
not I_67154 (I1145205,I1145197);
nor I_67155 (I1144767,I1145205,I1145010);
nand I_67156 (I1145236,I1145205,I1144855);
not I_67157 (I1145253,I699451);
nand I_67158 (I1145270,I1145253,I1144959);
nand I_67159 (I1145287,I1145205,I1145270);
nand I_67160 (I1144758,I1145287,I1145236);
nand I_67161 (I1144755,I1145270,I1145154);
not I_67162 (I1145359,I3570);
DFFARX1 I_67163 (I210718,I3563,I1145359,I1145385,);
and I_67164 (I1145393,I1145385,I210721);
DFFARX1 I_67165 (I1145393,I3563,I1145359,I1145342,);
DFFARX1 I_67166 (I210721,I3563,I1145359,I1145433,);
not I_67167 (I1145441,I210736);
not I_67168 (I1145458,I210742);
nand I_67169 (I1145475,I1145458,I1145441);
nor I_67170 (I1145330,I1145433,I1145475);
DFFARX1 I_67171 (I1145475,I3563,I1145359,I1145515,);
not I_67172 (I1145351,I1145515);
not I_67173 (I1145537,I210730);
nand I_67174 (I1145554,I1145458,I1145537);
DFFARX1 I_67175 (I1145554,I3563,I1145359,I1145580,);
not I_67176 (I1145588,I1145580);
not I_67177 (I1145605,I210727);
nand I_67178 (I1145622,I1145605,I210724);
and I_67179 (I1145639,I1145441,I1145622);
nor I_67180 (I1145656,I1145554,I1145639);
DFFARX1 I_67181 (I1145656,I3563,I1145359,I1145327,);
DFFARX1 I_67182 (I1145639,I3563,I1145359,I1145348,);
nor I_67183 (I1145701,I210727,I210718);
nor I_67184 (I1145339,I1145554,I1145701);
or I_67185 (I1145732,I210727,I210718);
nor I_67186 (I1145749,I210733,I210739);
DFFARX1 I_67187 (I1145749,I3563,I1145359,I1145775,);
not I_67188 (I1145783,I1145775);
nor I_67189 (I1145345,I1145783,I1145588);
nand I_67190 (I1145814,I1145783,I1145433);
not I_67191 (I1145831,I210733);
nand I_67192 (I1145848,I1145831,I1145537);
nand I_67193 (I1145865,I1145783,I1145848);
nand I_67194 (I1145336,I1145865,I1145814);
nand I_67195 (I1145333,I1145848,I1145732);
not I_67196 (I1145937,I3570);
DFFARX1 I_67197 (I1369635,I3563,I1145937,I1145963,);
and I_67198 (I1145971,I1145963,I1369617);
DFFARX1 I_67199 (I1145971,I3563,I1145937,I1145920,);
DFFARX1 I_67200 (I1369608,I3563,I1145937,I1146011,);
not I_67201 (I1146019,I1369623);
not I_67202 (I1146036,I1369611);
nand I_67203 (I1146053,I1146036,I1146019);
nor I_67204 (I1145908,I1146011,I1146053);
DFFARX1 I_67205 (I1146053,I3563,I1145937,I1146093,);
not I_67206 (I1145929,I1146093);
not I_67207 (I1146115,I1369620);
nand I_67208 (I1146132,I1146036,I1146115);
DFFARX1 I_67209 (I1146132,I3563,I1145937,I1146158,);
not I_67210 (I1146166,I1146158);
not I_67211 (I1146183,I1369629);
nand I_67212 (I1146200,I1146183,I1369608);
and I_67213 (I1146217,I1146019,I1146200);
nor I_67214 (I1146234,I1146132,I1146217);
DFFARX1 I_67215 (I1146234,I3563,I1145937,I1145905,);
DFFARX1 I_67216 (I1146217,I3563,I1145937,I1145926,);
nor I_67217 (I1146279,I1369629,I1369632);
nor I_67218 (I1145917,I1146132,I1146279);
or I_67219 (I1146310,I1369629,I1369632);
nor I_67220 (I1146327,I1369626,I1369614);
DFFARX1 I_67221 (I1146327,I3563,I1145937,I1146353,);
not I_67222 (I1146361,I1146353);
nor I_67223 (I1145923,I1146361,I1146166);
nand I_67224 (I1146392,I1146361,I1146011);
not I_67225 (I1146409,I1369626);
nand I_67226 (I1146426,I1146409,I1146115);
nand I_67227 (I1146443,I1146361,I1146426);
nand I_67228 (I1145914,I1146443,I1146392);
nand I_67229 (I1145911,I1146426,I1146310);
not I_67230 (I1146515,I3570);
DFFARX1 I_67231 (I765936,I3563,I1146515,I1146541,);
and I_67232 (I1146549,I1146541,I765924);
DFFARX1 I_67233 (I1146549,I3563,I1146515,I1146498,);
DFFARX1 I_67234 (I765927,I3563,I1146515,I1146589,);
not I_67235 (I1146597,I765921);
not I_67236 (I1146614,I765945);
nand I_67237 (I1146631,I1146614,I1146597);
nor I_67238 (I1146486,I1146589,I1146631);
DFFARX1 I_67239 (I1146631,I3563,I1146515,I1146671,);
not I_67240 (I1146507,I1146671);
not I_67241 (I1146693,I765933);
nand I_67242 (I1146710,I1146614,I1146693);
DFFARX1 I_67243 (I1146710,I3563,I1146515,I1146736,);
not I_67244 (I1146744,I1146736);
not I_67245 (I1146761,I765942);
nand I_67246 (I1146778,I1146761,I765939);
and I_67247 (I1146795,I1146597,I1146778);
nor I_67248 (I1146812,I1146710,I1146795);
DFFARX1 I_67249 (I1146812,I3563,I1146515,I1146483,);
DFFARX1 I_67250 (I1146795,I3563,I1146515,I1146504,);
nor I_67251 (I1146857,I765942,I765930);
nor I_67252 (I1146495,I1146710,I1146857);
or I_67253 (I1146888,I765942,I765930);
nor I_67254 (I1146905,I765921,I765924);
DFFARX1 I_67255 (I1146905,I3563,I1146515,I1146931,);
not I_67256 (I1146939,I1146931);
nor I_67257 (I1146501,I1146939,I1146744);
nand I_67258 (I1146970,I1146939,I1146589);
not I_67259 (I1146987,I765921);
nand I_67260 (I1147004,I1146987,I1146693);
nand I_67261 (I1147021,I1146939,I1147004);
nand I_67262 (I1146492,I1147021,I1146970);
nand I_67263 (I1146489,I1147004,I1146888);
not I_67264 (I1147093,I3570);
DFFARX1 I_67265 (I130451,I3563,I1147093,I1147119,);
and I_67266 (I1147127,I1147119,I130427);
DFFARX1 I_67267 (I1147127,I3563,I1147093,I1147076,);
DFFARX1 I_67268 (I130445,I3563,I1147093,I1147167,);
not I_67269 (I1147175,I130433);
not I_67270 (I1147192,I130430);
nand I_67271 (I1147209,I1147192,I1147175);
nor I_67272 (I1147064,I1147167,I1147209);
DFFARX1 I_67273 (I1147209,I3563,I1147093,I1147249,);
not I_67274 (I1147085,I1147249);
not I_67275 (I1147271,I130439);
nand I_67276 (I1147288,I1147192,I1147271);
DFFARX1 I_67277 (I1147288,I3563,I1147093,I1147314,);
not I_67278 (I1147322,I1147314);
not I_67279 (I1147339,I130430);
nand I_67280 (I1147356,I1147339,I130448);
and I_67281 (I1147373,I1147175,I1147356);
nor I_67282 (I1147390,I1147288,I1147373);
DFFARX1 I_67283 (I1147390,I3563,I1147093,I1147061,);
DFFARX1 I_67284 (I1147373,I3563,I1147093,I1147082,);
nor I_67285 (I1147435,I130430,I130442);
nor I_67286 (I1147073,I1147288,I1147435);
or I_67287 (I1147466,I130430,I130442);
nor I_67288 (I1147483,I130436,I130427);
DFFARX1 I_67289 (I1147483,I3563,I1147093,I1147509,);
not I_67290 (I1147517,I1147509);
nor I_67291 (I1147079,I1147517,I1147322);
nand I_67292 (I1147548,I1147517,I1147167);
not I_67293 (I1147565,I130436);
nand I_67294 (I1147582,I1147565,I1147271);
nand I_67295 (I1147599,I1147517,I1147582);
nand I_67296 (I1147070,I1147599,I1147548);
nand I_67297 (I1147067,I1147582,I1147466);
not I_67298 (I1147671,I3570);
DFFARX1 I_67299 (I1008551,I3563,I1147671,I1147697,);
and I_67300 (I1147705,I1147697,I1008545);
DFFARX1 I_67301 (I1147705,I3563,I1147671,I1147654,);
DFFARX1 I_67302 (I1008563,I3563,I1147671,I1147745,);
not I_67303 (I1147753,I1008554);
not I_67304 (I1147770,I1008566);
nand I_67305 (I1147787,I1147770,I1147753);
nor I_67306 (I1147642,I1147745,I1147787);
DFFARX1 I_67307 (I1147787,I3563,I1147671,I1147827,);
not I_67308 (I1147663,I1147827);
not I_67309 (I1147849,I1008572);
nand I_67310 (I1147866,I1147770,I1147849);
DFFARX1 I_67311 (I1147866,I3563,I1147671,I1147892,);
not I_67312 (I1147900,I1147892);
not I_67313 (I1147917,I1008548);
nand I_67314 (I1147934,I1147917,I1008569);
and I_67315 (I1147951,I1147753,I1147934);
nor I_67316 (I1147968,I1147866,I1147951);
DFFARX1 I_67317 (I1147968,I3563,I1147671,I1147639,);
DFFARX1 I_67318 (I1147951,I3563,I1147671,I1147660,);
nor I_67319 (I1148013,I1008548,I1008560);
nor I_67320 (I1147651,I1147866,I1148013);
or I_67321 (I1148044,I1008548,I1008560);
nor I_67322 (I1148061,I1008545,I1008557);
DFFARX1 I_67323 (I1148061,I3563,I1147671,I1148087,);
not I_67324 (I1148095,I1148087);
nor I_67325 (I1147657,I1148095,I1147900);
nand I_67326 (I1148126,I1148095,I1147745);
not I_67327 (I1148143,I1008545);
nand I_67328 (I1148160,I1148143,I1147849);
nand I_67329 (I1148177,I1148095,I1148160);
nand I_67330 (I1147648,I1148177,I1148126);
nand I_67331 (I1147645,I1148160,I1148044);
not I_67332 (I1148249,I3570);
DFFARX1 I_67333 (I205363,I3563,I1148249,I1148275,);
and I_67334 (I1148283,I1148275,I205366);
DFFARX1 I_67335 (I1148283,I3563,I1148249,I1148232,);
DFFARX1 I_67336 (I205366,I3563,I1148249,I1148323,);
not I_67337 (I1148331,I205381);
not I_67338 (I1148348,I205387);
nand I_67339 (I1148365,I1148348,I1148331);
nor I_67340 (I1148220,I1148323,I1148365);
DFFARX1 I_67341 (I1148365,I3563,I1148249,I1148405,);
not I_67342 (I1148241,I1148405);
not I_67343 (I1148427,I205375);
nand I_67344 (I1148444,I1148348,I1148427);
DFFARX1 I_67345 (I1148444,I3563,I1148249,I1148470,);
not I_67346 (I1148478,I1148470);
not I_67347 (I1148495,I205372);
nand I_67348 (I1148512,I1148495,I205369);
and I_67349 (I1148529,I1148331,I1148512);
nor I_67350 (I1148546,I1148444,I1148529);
DFFARX1 I_67351 (I1148546,I3563,I1148249,I1148217,);
DFFARX1 I_67352 (I1148529,I3563,I1148249,I1148238,);
nor I_67353 (I1148591,I205372,I205363);
nor I_67354 (I1148229,I1148444,I1148591);
or I_67355 (I1148622,I205372,I205363);
nor I_67356 (I1148639,I205378,I205384);
DFFARX1 I_67357 (I1148639,I3563,I1148249,I1148665,);
not I_67358 (I1148673,I1148665);
nor I_67359 (I1148235,I1148673,I1148478);
nand I_67360 (I1148704,I1148673,I1148323);
not I_67361 (I1148721,I205378);
nand I_67362 (I1148738,I1148721,I1148427);
nand I_67363 (I1148755,I1148673,I1148738);
nand I_67364 (I1148226,I1148755,I1148704);
nand I_67365 (I1148223,I1148738,I1148622);
not I_67366 (I1148827,I3570);
DFFARX1 I_67367 (I412399,I3563,I1148827,I1148853,);
and I_67368 (I1148861,I1148853,I412384);
DFFARX1 I_67369 (I1148861,I3563,I1148827,I1148810,);
DFFARX1 I_67370 (I412390,I3563,I1148827,I1148901,);
not I_67371 (I1148909,I412372);
not I_67372 (I1148926,I412393);
nand I_67373 (I1148943,I1148926,I1148909);
nor I_67374 (I1148798,I1148901,I1148943);
DFFARX1 I_67375 (I1148943,I3563,I1148827,I1148983,);
not I_67376 (I1148819,I1148983);
not I_67377 (I1149005,I412396);
nand I_67378 (I1149022,I1148926,I1149005);
DFFARX1 I_67379 (I1149022,I3563,I1148827,I1149048,);
not I_67380 (I1149056,I1149048);
not I_67381 (I1149073,I412387);
nand I_67382 (I1149090,I1149073,I412375);
and I_67383 (I1149107,I1148909,I1149090);
nor I_67384 (I1149124,I1149022,I1149107);
DFFARX1 I_67385 (I1149124,I3563,I1148827,I1148795,);
DFFARX1 I_67386 (I1149107,I3563,I1148827,I1148816,);
nor I_67387 (I1149169,I412387,I412381);
nor I_67388 (I1148807,I1149022,I1149169);
or I_67389 (I1149200,I412387,I412381);
nor I_67390 (I1149217,I412378,I412372);
DFFARX1 I_67391 (I1149217,I3563,I1148827,I1149243,);
not I_67392 (I1149251,I1149243);
nor I_67393 (I1148813,I1149251,I1149056);
nand I_67394 (I1149282,I1149251,I1148901);
not I_67395 (I1149299,I412378);
nand I_67396 (I1149316,I1149299,I1149005);
nand I_67397 (I1149333,I1149251,I1149316);
nand I_67398 (I1148804,I1149333,I1149282);
nand I_67399 (I1148801,I1149316,I1149200);
not I_67400 (I1149405,I3570);
DFFARX1 I_67401 (I1381535,I3563,I1149405,I1149431,);
and I_67402 (I1149439,I1149431,I1381517);
DFFARX1 I_67403 (I1149439,I3563,I1149405,I1149388,);
DFFARX1 I_67404 (I1381508,I3563,I1149405,I1149479,);
not I_67405 (I1149487,I1381523);
not I_67406 (I1149504,I1381511);
nand I_67407 (I1149521,I1149504,I1149487);
nor I_67408 (I1149376,I1149479,I1149521);
DFFARX1 I_67409 (I1149521,I3563,I1149405,I1149561,);
not I_67410 (I1149397,I1149561);
not I_67411 (I1149583,I1381520);
nand I_67412 (I1149600,I1149504,I1149583);
DFFARX1 I_67413 (I1149600,I3563,I1149405,I1149626,);
not I_67414 (I1149634,I1149626);
not I_67415 (I1149651,I1381529);
nand I_67416 (I1149668,I1149651,I1381508);
and I_67417 (I1149685,I1149487,I1149668);
nor I_67418 (I1149702,I1149600,I1149685);
DFFARX1 I_67419 (I1149702,I3563,I1149405,I1149373,);
DFFARX1 I_67420 (I1149685,I3563,I1149405,I1149394,);
nor I_67421 (I1149747,I1381529,I1381532);
nor I_67422 (I1149385,I1149600,I1149747);
or I_67423 (I1149778,I1381529,I1381532);
nor I_67424 (I1149795,I1381526,I1381514);
DFFARX1 I_67425 (I1149795,I3563,I1149405,I1149821,);
not I_67426 (I1149829,I1149821);
nor I_67427 (I1149391,I1149829,I1149634);
nand I_67428 (I1149860,I1149829,I1149479);
not I_67429 (I1149877,I1381526);
nand I_67430 (I1149894,I1149877,I1149583);
nand I_67431 (I1149911,I1149829,I1149894);
nand I_67432 (I1149382,I1149911,I1149860);
nand I_67433 (I1149379,I1149894,I1149778);
not I_67434 (I1149983,I3570);
DFFARX1 I_67435 (I1363090,I3563,I1149983,I1150009,);
and I_67436 (I1150017,I1150009,I1363072);
DFFARX1 I_67437 (I1150017,I3563,I1149983,I1149966,);
DFFARX1 I_67438 (I1363063,I3563,I1149983,I1150057,);
not I_67439 (I1150065,I1363078);
not I_67440 (I1150082,I1363066);
nand I_67441 (I1150099,I1150082,I1150065);
nor I_67442 (I1149954,I1150057,I1150099);
DFFARX1 I_67443 (I1150099,I3563,I1149983,I1150139,);
not I_67444 (I1149975,I1150139);
not I_67445 (I1150161,I1363075);
nand I_67446 (I1150178,I1150082,I1150161);
DFFARX1 I_67447 (I1150178,I3563,I1149983,I1150204,);
not I_67448 (I1150212,I1150204);
not I_67449 (I1150229,I1363084);
nand I_67450 (I1150246,I1150229,I1363063);
and I_67451 (I1150263,I1150065,I1150246);
nor I_67452 (I1150280,I1150178,I1150263);
DFFARX1 I_67453 (I1150280,I3563,I1149983,I1149951,);
DFFARX1 I_67454 (I1150263,I3563,I1149983,I1149972,);
nor I_67455 (I1150325,I1363084,I1363087);
nor I_67456 (I1149963,I1150178,I1150325);
or I_67457 (I1150356,I1363084,I1363087);
nor I_67458 (I1150373,I1363081,I1363069);
DFFARX1 I_67459 (I1150373,I3563,I1149983,I1150399,);
not I_67460 (I1150407,I1150399);
nor I_67461 (I1149969,I1150407,I1150212);
nand I_67462 (I1150438,I1150407,I1150057);
not I_67463 (I1150455,I1363081);
nand I_67464 (I1150472,I1150455,I1150161);
nand I_67465 (I1150489,I1150407,I1150472);
nand I_67466 (I1149960,I1150489,I1150438);
nand I_67467 (I1149957,I1150472,I1150356);
not I_67468 (I1150561,I3570);
DFFARX1 I_67469 (I472450,I3563,I1150561,I1150587,);
and I_67470 (I1150595,I1150587,I472465);
DFFARX1 I_67471 (I1150595,I3563,I1150561,I1150544,);
DFFARX1 I_67472 (I472468,I3563,I1150561,I1150635,);
not I_67473 (I1150643,I472462);
not I_67474 (I1150660,I472477);
nand I_67475 (I1150677,I1150660,I1150643);
nor I_67476 (I1150532,I1150635,I1150677);
DFFARX1 I_67477 (I1150677,I3563,I1150561,I1150717,);
not I_67478 (I1150553,I1150717);
not I_67479 (I1150739,I472453);
nand I_67480 (I1150756,I1150660,I1150739);
DFFARX1 I_67481 (I1150756,I3563,I1150561,I1150782,);
not I_67482 (I1150790,I1150782);
not I_67483 (I1150807,I472456);
nand I_67484 (I1150824,I1150807,I472450);
and I_67485 (I1150841,I1150643,I1150824);
nor I_67486 (I1150858,I1150756,I1150841);
DFFARX1 I_67487 (I1150858,I3563,I1150561,I1150529,);
DFFARX1 I_67488 (I1150841,I3563,I1150561,I1150550,);
nor I_67489 (I1150903,I472456,I472459);
nor I_67490 (I1150541,I1150756,I1150903);
or I_67491 (I1150934,I472456,I472459);
nor I_67492 (I1150951,I472474,I472471);
DFFARX1 I_67493 (I1150951,I3563,I1150561,I1150977,);
not I_67494 (I1150985,I1150977);
nor I_67495 (I1150547,I1150985,I1150790);
nand I_67496 (I1151016,I1150985,I1150635);
not I_67497 (I1151033,I472474);
nand I_67498 (I1151050,I1151033,I1150739);
nand I_67499 (I1151067,I1150985,I1151050);
nand I_67500 (I1150538,I1151067,I1151016);
nand I_67501 (I1150535,I1151050,I1150934);
not I_67502 (I1151139,I3570);
DFFARX1 I_67503 (I352321,I3563,I1151139,I1151165,);
and I_67504 (I1151173,I1151165,I352306);
DFFARX1 I_67505 (I1151173,I3563,I1151139,I1151122,);
DFFARX1 I_67506 (I352312,I3563,I1151139,I1151213,);
not I_67507 (I1151221,I352294);
not I_67508 (I1151238,I352315);
nand I_67509 (I1151255,I1151238,I1151221);
nor I_67510 (I1151110,I1151213,I1151255);
DFFARX1 I_67511 (I1151255,I3563,I1151139,I1151295,);
not I_67512 (I1151131,I1151295);
not I_67513 (I1151317,I352318);
nand I_67514 (I1151334,I1151238,I1151317);
DFFARX1 I_67515 (I1151334,I3563,I1151139,I1151360,);
not I_67516 (I1151368,I1151360);
not I_67517 (I1151385,I352309);
nand I_67518 (I1151402,I1151385,I352297);
and I_67519 (I1151419,I1151221,I1151402);
nor I_67520 (I1151436,I1151334,I1151419);
DFFARX1 I_67521 (I1151436,I3563,I1151139,I1151107,);
DFFARX1 I_67522 (I1151419,I3563,I1151139,I1151128,);
nor I_67523 (I1151481,I352309,I352303);
nor I_67524 (I1151119,I1151334,I1151481);
or I_67525 (I1151512,I352309,I352303);
nor I_67526 (I1151529,I352300,I352294);
DFFARX1 I_67527 (I1151529,I3563,I1151139,I1151555,);
not I_67528 (I1151563,I1151555);
nor I_67529 (I1151125,I1151563,I1151368);
nand I_67530 (I1151594,I1151563,I1151213);
not I_67531 (I1151611,I352300);
nand I_67532 (I1151628,I1151611,I1151317);
nand I_67533 (I1151645,I1151563,I1151628);
nand I_67534 (I1151116,I1151645,I1151594);
nand I_67535 (I1151113,I1151628,I1151512);
not I_67536 (I1151717,I3570);
DFFARX1 I_67537 (I314377,I3563,I1151717,I1151743,);
and I_67538 (I1151751,I1151743,I314362);
DFFARX1 I_67539 (I1151751,I3563,I1151717,I1151700,);
DFFARX1 I_67540 (I314368,I3563,I1151717,I1151791,);
not I_67541 (I1151799,I314350);
not I_67542 (I1151816,I314371);
nand I_67543 (I1151833,I1151816,I1151799);
nor I_67544 (I1151688,I1151791,I1151833);
DFFARX1 I_67545 (I1151833,I3563,I1151717,I1151873,);
not I_67546 (I1151709,I1151873);
not I_67547 (I1151895,I314374);
nand I_67548 (I1151912,I1151816,I1151895);
DFFARX1 I_67549 (I1151912,I3563,I1151717,I1151938,);
not I_67550 (I1151946,I1151938);
not I_67551 (I1151963,I314365);
nand I_67552 (I1151980,I1151963,I314353);
and I_67553 (I1151997,I1151799,I1151980);
nor I_67554 (I1152014,I1151912,I1151997);
DFFARX1 I_67555 (I1152014,I3563,I1151717,I1151685,);
DFFARX1 I_67556 (I1151997,I3563,I1151717,I1151706,);
nor I_67557 (I1152059,I314365,I314359);
nor I_67558 (I1151697,I1151912,I1152059);
or I_67559 (I1152090,I314365,I314359);
nor I_67560 (I1152107,I314356,I314350);
DFFARX1 I_67561 (I1152107,I3563,I1151717,I1152133,);
not I_67562 (I1152141,I1152133);
nor I_67563 (I1151703,I1152141,I1151946);
nand I_67564 (I1152172,I1152141,I1151791);
not I_67565 (I1152189,I314356);
nand I_67566 (I1152206,I1152189,I1151895);
nand I_67567 (I1152223,I1152141,I1152206);
nand I_67568 (I1151694,I1152223,I1152172);
nand I_67569 (I1151691,I1152206,I1152090);
not I_67570 (I1152295,I3570);
DFFARX1 I_67571 (I1266014,I3563,I1152295,I1152321,);
and I_67572 (I1152329,I1152321,I1266008);
DFFARX1 I_67573 (I1152329,I3563,I1152295,I1152278,);
DFFARX1 I_67574 (I1265993,I3563,I1152295,I1152369,);
not I_67575 (I1152377,I1265999);
not I_67576 (I1152394,I1266011);
nand I_67577 (I1152411,I1152394,I1152377);
nor I_67578 (I1152266,I1152369,I1152411);
DFFARX1 I_67579 (I1152411,I3563,I1152295,I1152451,);
not I_67580 (I1152287,I1152451);
not I_67581 (I1152473,I1265993);
nand I_67582 (I1152490,I1152394,I1152473);
DFFARX1 I_67583 (I1152490,I3563,I1152295,I1152516,);
not I_67584 (I1152524,I1152516);
not I_67585 (I1152541,I1266017);
nand I_67586 (I1152558,I1152541,I1266005);
and I_67587 (I1152575,I1152377,I1152558);
nor I_67588 (I1152592,I1152490,I1152575);
DFFARX1 I_67589 (I1152592,I3563,I1152295,I1152263,);
DFFARX1 I_67590 (I1152575,I3563,I1152295,I1152284,);
nor I_67591 (I1152637,I1266017,I1265996);
nor I_67592 (I1152275,I1152490,I1152637);
or I_67593 (I1152668,I1266017,I1265996);
nor I_67594 (I1152685,I1266002,I1265996);
DFFARX1 I_67595 (I1152685,I3563,I1152295,I1152711,);
not I_67596 (I1152719,I1152711);
nor I_67597 (I1152281,I1152719,I1152524);
nand I_67598 (I1152750,I1152719,I1152369);
not I_67599 (I1152767,I1266002);
nand I_67600 (I1152784,I1152767,I1152473);
nand I_67601 (I1152801,I1152719,I1152784);
nand I_67602 (I1152272,I1152801,I1152750);
nand I_67603 (I1152269,I1152784,I1152668);
not I_67604 (I1152873,I3570);
DFFARX1 I_67605 (I744550,I3563,I1152873,I1152899,);
and I_67606 (I1152907,I1152899,I744538);
DFFARX1 I_67607 (I1152907,I3563,I1152873,I1152856,);
DFFARX1 I_67608 (I744541,I3563,I1152873,I1152947,);
not I_67609 (I1152955,I744535);
not I_67610 (I1152972,I744559);
nand I_67611 (I1152989,I1152972,I1152955);
nor I_67612 (I1152844,I1152947,I1152989);
DFFARX1 I_67613 (I1152989,I3563,I1152873,I1153029,);
not I_67614 (I1152865,I1153029);
not I_67615 (I1153051,I744547);
nand I_67616 (I1153068,I1152972,I1153051);
DFFARX1 I_67617 (I1153068,I3563,I1152873,I1153094,);
not I_67618 (I1153102,I1153094);
not I_67619 (I1153119,I744556);
nand I_67620 (I1153136,I1153119,I744553);
and I_67621 (I1153153,I1152955,I1153136);
nor I_67622 (I1153170,I1153068,I1153153);
DFFARX1 I_67623 (I1153170,I3563,I1152873,I1152841,);
DFFARX1 I_67624 (I1153153,I3563,I1152873,I1152862,);
nor I_67625 (I1153215,I744556,I744544);
nor I_67626 (I1152853,I1153068,I1153215);
or I_67627 (I1153246,I744556,I744544);
nor I_67628 (I1153263,I744535,I744538);
DFFARX1 I_67629 (I1153263,I3563,I1152873,I1153289,);
not I_67630 (I1153297,I1153289);
nor I_67631 (I1152859,I1153297,I1153102);
nand I_67632 (I1153328,I1153297,I1152947);
not I_67633 (I1153345,I744535);
nand I_67634 (I1153362,I1153345,I1153051);
nand I_67635 (I1153379,I1153297,I1153362);
nand I_67636 (I1152850,I1153379,I1153328);
nand I_67637 (I1152847,I1153362,I1153246);
not I_67638 (I1153451,I3570);
DFFARX1 I_67639 (I794836,I3563,I1153451,I1153477,);
and I_67640 (I1153485,I1153477,I794824);
DFFARX1 I_67641 (I1153485,I3563,I1153451,I1153434,);
DFFARX1 I_67642 (I794827,I3563,I1153451,I1153525,);
not I_67643 (I1153533,I794821);
not I_67644 (I1153550,I794845);
nand I_67645 (I1153567,I1153550,I1153533);
nor I_67646 (I1153422,I1153525,I1153567);
DFFARX1 I_67647 (I1153567,I3563,I1153451,I1153607,);
not I_67648 (I1153443,I1153607);
not I_67649 (I1153629,I794833);
nand I_67650 (I1153646,I1153550,I1153629);
DFFARX1 I_67651 (I1153646,I3563,I1153451,I1153672,);
not I_67652 (I1153680,I1153672);
not I_67653 (I1153697,I794842);
nand I_67654 (I1153714,I1153697,I794839);
and I_67655 (I1153731,I1153533,I1153714);
nor I_67656 (I1153748,I1153646,I1153731);
DFFARX1 I_67657 (I1153748,I3563,I1153451,I1153419,);
DFFARX1 I_67658 (I1153731,I3563,I1153451,I1153440,);
nor I_67659 (I1153793,I794842,I794830);
nor I_67660 (I1153431,I1153646,I1153793);
or I_67661 (I1153824,I794842,I794830);
nor I_67662 (I1153841,I794821,I794824);
DFFARX1 I_67663 (I1153841,I3563,I1153451,I1153867,);
not I_67664 (I1153875,I1153867);
nor I_67665 (I1153437,I1153875,I1153680);
nand I_67666 (I1153906,I1153875,I1153525);
not I_67667 (I1153923,I794821);
nand I_67668 (I1153940,I1153923,I1153629);
nand I_67669 (I1153957,I1153875,I1153940);
nand I_67670 (I1153428,I1153957,I1153906);
nand I_67671 (I1153425,I1153940,I1153824);
not I_67672 (I1154029,I3570);
DFFARX1 I_67673 (I20284,I3563,I1154029,I1154055,);
and I_67674 (I1154063,I1154055,I20287);
DFFARX1 I_67675 (I1154063,I3563,I1154029,I1154012,);
DFFARX1 I_67676 (I20287,I3563,I1154029,I1154103,);
not I_67677 (I1154111,I20290);
not I_67678 (I1154128,I20305);
nand I_67679 (I1154145,I1154128,I1154111);
nor I_67680 (I1154000,I1154103,I1154145);
DFFARX1 I_67681 (I1154145,I3563,I1154029,I1154185,);
not I_67682 (I1154021,I1154185);
not I_67683 (I1154207,I20299);
nand I_67684 (I1154224,I1154128,I1154207);
DFFARX1 I_67685 (I1154224,I3563,I1154029,I1154250,);
not I_67686 (I1154258,I1154250);
not I_67687 (I1154275,I20302);
nand I_67688 (I1154292,I1154275,I20284);
and I_67689 (I1154309,I1154111,I1154292);
nor I_67690 (I1154326,I1154224,I1154309);
DFFARX1 I_67691 (I1154326,I3563,I1154029,I1153997,);
DFFARX1 I_67692 (I1154309,I3563,I1154029,I1154018,);
nor I_67693 (I1154371,I20302,I20296);
nor I_67694 (I1154009,I1154224,I1154371);
or I_67695 (I1154402,I20302,I20296);
nor I_67696 (I1154419,I20293,I20308);
DFFARX1 I_67697 (I1154419,I3563,I1154029,I1154445,);
not I_67698 (I1154453,I1154445);
nor I_67699 (I1154015,I1154453,I1154258);
nand I_67700 (I1154484,I1154453,I1154103);
not I_67701 (I1154501,I20293);
nand I_67702 (I1154518,I1154501,I1154207);
nand I_67703 (I1154535,I1154453,I1154518);
nand I_67704 (I1154006,I1154535,I1154484);
nand I_67705 (I1154003,I1154518,I1154402);
not I_67706 (I1154607,I3570);
DFFARX1 I_67707 (I942013,I3563,I1154607,I1154633,);
and I_67708 (I1154641,I1154633,I942007);
DFFARX1 I_67709 (I1154641,I3563,I1154607,I1154590,);
DFFARX1 I_67710 (I942025,I3563,I1154607,I1154681,);
not I_67711 (I1154689,I942016);
not I_67712 (I1154706,I942028);
nand I_67713 (I1154723,I1154706,I1154689);
nor I_67714 (I1154578,I1154681,I1154723);
DFFARX1 I_67715 (I1154723,I3563,I1154607,I1154763,);
not I_67716 (I1154599,I1154763);
not I_67717 (I1154785,I942034);
nand I_67718 (I1154802,I1154706,I1154785);
DFFARX1 I_67719 (I1154802,I3563,I1154607,I1154828,);
not I_67720 (I1154836,I1154828);
not I_67721 (I1154853,I942010);
nand I_67722 (I1154870,I1154853,I942031);
and I_67723 (I1154887,I1154689,I1154870);
nor I_67724 (I1154904,I1154802,I1154887);
DFFARX1 I_67725 (I1154904,I3563,I1154607,I1154575,);
DFFARX1 I_67726 (I1154887,I3563,I1154607,I1154596,);
nor I_67727 (I1154949,I942010,I942022);
nor I_67728 (I1154587,I1154802,I1154949);
or I_67729 (I1154980,I942010,I942022);
nor I_67730 (I1154997,I942007,I942019);
DFFARX1 I_67731 (I1154997,I3563,I1154607,I1155023,);
not I_67732 (I1155031,I1155023);
nor I_67733 (I1154593,I1155031,I1154836);
nand I_67734 (I1155062,I1155031,I1154681);
not I_67735 (I1155079,I942007);
nand I_67736 (I1155096,I1155079,I1154785);
nand I_67737 (I1155113,I1155031,I1155096);
nand I_67738 (I1154584,I1155113,I1155062);
nand I_67739 (I1154581,I1155096,I1154980);
not I_67740 (I1155185,I3570);
DFFARX1 I_67741 (I37675,I3563,I1155185,I1155211,);
and I_67742 (I1155219,I1155211,I37678);
DFFARX1 I_67743 (I1155219,I3563,I1155185,I1155168,);
DFFARX1 I_67744 (I37678,I3563,I1155185,I1155259,);
not I_67745 (I1155267,I37681);
not I_67746 (I1155284,I37696);
nand I_67747 (I1155301,I1155284,I1155267);
nor I_67748 (I1155156,I1155259,I1155301);
DFFARX1 I_67749 (I1155301,I3563,I1155185,I1155341,);
not I_67750 (I1155177,I1155341);
not I_67751 (I1155363,I37690);
nand I_67752 (I1155380,I1155284,I1155363);
DFFARX1 I_67753 (I1155380,I3563,I1155185,I1155406,);
not I_67754 (I1155414,I1155406);
not I_67755 (I1155431,I37693);
nand I_67756 (I1155448,I1155431,I37675);
and I_67757 (I1155465,I1155267,I1155448);
nor I_67758 (I1155482,I1155380,I1155465);
DFFARX1 I_67759 (I1155482,I3563,I1155185,I1155153,);
DFFARX1 I_67760 (I1155465,I3563,I1155185,I1155174,);
nor I_67761 (I1155527,I37693,I37687);
nor I_67762 (I1155165,I1155380,I1155527);
or I_67763 (I1155558,I37693,I37687);
nor I_67764 (I1155575,I37684,I37699);
DFFARX1 I_67765 (I1155575,I3563,I1155185,I1155601,);
not I_67766 (I1155609,I1155601);
nor I_67767 (I1155171,I1155609,I1155414);
nand I_67768 (I1155640,I1155609,I1155259);
not I_67769 (I1155657,I37684);
nand I_67770 (I1155674,I1155657,I1155363);
nand I_67771 (I1155691,I1155609,I1155674);
nand I_67772 (I1155162,I1155691,I1155640);
nand I_67773 (I1155159,I1155674,I1155558);
not I_67774 (I1155763,I3570);
DFFARX1 I_67775 (I1343455,I3563,I1155763,I1155789,);
and I_67776 (I1155797,I1155789,I1343437);
DFFARX1 I_67777 (I1155797,I3563,I1155763,I1155746,);
DFFARX1 I_67778 (I1343428,I3563,I1155763,I1155837,);
not I_67779 (I1155845,I1343443);
not I_67780 (I1155862,I1343431);
nand I_67781 (I1155879,I1155862,I1155845);
nor I_67782 (I1155734,I1155837,I1155879);
DFFARX1 I_67783 (I1155879,I3563,I1155763,I1155919,);
not I_67784 (I1155755,I1155919);
not I_67785 (I1155941,I1343440);
nand I_67786 (I1155958,I1155862,I1155941);
DFFARX1 I_67787 (I1155958,I3563,I1155763,I1155984,);
not I_67788 (I1155992,I1155984);
not I_67789 (I1156009,I1343449);
nand I_67790 (I1156026,I1156009,I1343428);
and I_67791 (I1156043,I1155845,I1156026);
nor I_67792 (I1156060,I1155958,I1156043);
DFFARX1 I_67793 (I1156060,I3563,I1155763,I1155731,);
DFFARX1 I_67794 (I1156043,I3563,I1155763,I1155752,);
nor I_67795 (I1156105,I1343449,I1343452);
nor I_67796 (I1155743,I1155958,I1156105);
or I_67797 (I1156136,I1343449,I1343452);
nor I_67798 (I1156153,I1343446,I1343434);
DFFARX1 I_67799 (I1156153,I3563,I1155763,I1156179,);
not I_67800 (I1156187,I1156179);
nor I_67801 (I1155749,I1156187,I1155992);
nand I_67802 (I1156218,I1156187,I1155837);
not I_67803 (I1156235,I1343446);
nand I_67804 (I1156252,I1156235,I1155941);
nand I_67805 (I1156269,I1156187,I1156252);
nand I_67806 (I1155740,I1156269,I1156218);
nand I_67807 (I1155737,I1156252,I1156136);
not I_67808 (I1156341,I3570);
DFFARX1 I_67809 (I615656,I3563,I1156341,I1156367,);
and I_67810 (I1156375,I1156367,I615644);
DFFARX1 I_67811 (I1156375,I3563,I1156341,I1156324,);
DFFARX1 I_67812 (I615659,I3563,I1156341,I1156415,);
not I_67813 (I1156423,I615650);
not I_67814 (I1156440,I615641);
nand I_67815 (I1156457,I1156440,I1156423);
nor I_67816 (I1156312,I1156415,I1156457);
DFFARX1 I_67817 (I1156457,I3563,I1156341,I1156497,);
not I_67818 (I1156333,I1156497);
not I_67819 (I1156519,I615647);
nand I_67820 (I1156536,I1156440,I1156519);
DFFARX1 I_67821 (I1156536,I3563,I1156341,I1156562,);
not I_67822 (I1156570,I1156562);
not I_67823 (I1156587,I615662);
nand I_67824 (I1156604,I1156587,I615665);
and I_67825 (I1156621,I1156423,I1156604);
nor I_67826 (I1156638,I1156536,I1156621);
DFFARX1 I_67827 (I1156638,I3563,I1156341,I1156309,);
DFFARX1 I_67828 (I1156621,I3563,I1156341,I1156330,);
nor I_67829 (I1156683,I615662,I615641);
nor I_67830 (I1156321,I1156536,I1156683);
or I_67831 (I1156714,I615662,I615641);
nor I_67832 (I1156731,I615653,I615644);
DFFARX1 I_67833 (I1156731,I3563,I1156341,I1156757,);
not I_67834 (I1156765,I1156757);
nor I_67835 (I1156327,I1156765,I1156570);
nand I_67836 (I1156796,I1156765,I1156415);
not I_67837 (I1156813,I615653);
nand I_67838 (I1156830,I1156813,I1156519);
nand I_67839 (I1156847,I1156765,I1156830);
nand I_67840 (I1156318,I1156847,I1156796);
nand I_67841 (I1156315,I1156830,I1156714);
not I_67842 (I1156919,I3570);
DFFARX1 I_67843 (I321228,I3563,I1156919,I1156945,);
and I_67844 (I1156953,I1156945,I321213);
DFFARX1 I_67845 (I1156953,I3563,I1156919,I1156902,);
DFFARX1 I_67846 (I321219,I3563,I1156919,I1156993,);
not I_67847 (I1157001,I321201);
not I_67848 (I1157018,I321222);
nand I_67849 (I1157035,I1157018,I1157001);
nor I_67850 (I1156890,I1156993,I1157035);
DFFARX1 I_67851 (I1157035,I3563,I1156919,I1157075,);
not I_67852 (I1156911,I1157075);
not I_67853 (I1157097,I321225);
nand I_67854 (I1157114,I1157018,I1157097);
DFFARX1 I_67855 (I1157114,I3563,I1156919,I1157140,);
not I_67856 (I1157148,I1157140);
not I_67857 (I1157165,I321216);
nand I_67858 (I1157182,I1157165,I321204);
and I_67859 (I1157199,I1157001,I1157182);
nor I_67860 (I1157216,I1157114,I1157199);
DFFARX1 I_67861 (I1157216,I3563,I1156919,I1156887,);
DFFARX1 I_67862 (I1157199,I3563,I1156919,I1156908,);
nor I_67863 (I1157261,I321216,I321210);
nor I_67864 (I1156899,I1157114,I1157261);
or I_67865 (I1157292,I321216,I321210);
nor I_67866 (I1157309,I321207,I321201);
DFFARX1 I_67867 (I1157309,I3563,I1156919,I1157335,);
not I_67868 (I1157343,I1157335);
nor I_67869 (I1156905,I1157343,I1157148);
nand I_67870 (I1157374,I1157343,I1156993);
not I_67871 (I1157391,I321207);
nand I_67872 (I1157408,I1157391,I1157097);
nand I_67873 (I1157425,I1157343,I1157408);
nand I_67874 (I1156896,I1157425,I1157374);
nand I_67875 (I1156893,I1157408,I1157292);
not I_67876 (I1157497,I3570);
DFFARX1 I_67877 (I938137,I3563,I1157497,I1157523,);
and I_67878 (I1157531,I1157523,I938131);
DFFARX1 I_67879 (I1157531,I3563,I1157497,I1157480,);
DFFARX1 I_67880 (I938149,I3563,I1157497,I1157571,);
not I_67881 (I1157579,I938140);
not I_67882 (I1157596,I938152);
nand I_67883 (I1157613,I1157596,I1157579);
nor I_67884 (I1157468,I1157571,I1157613);
DFFARX1 I_67885 (I1157613,I3563,I1157497,I1157653,);
not I_67886 (I1157489,I1157653);
not I_67887 (I1157675,I938158);
nand I_67888 (I1157692,I1157596,I1157675);
DFFARX1 I_67889 (I1157692,I3563,I1157497,I1157718,);
not I_67890 (I1157726,I1157718);
not I_67891 (I1157743,I938134);
nand I_67892 (I1157760,I1157743,I938155);
and I_67893 (I1157777,I1157579,I1157760);
nor I_67894 (I1157794,I1157692,I1157777);
DFFARX1 I_67895 (I1157794,I3563,I1157497,I1157465,);
DFFARX1 I_67896 (I1157777,I3563,I1157497,I1157486,);
nor I_67897 (I1157839,I938134,I938146);
nor I_67898 (I1157477,I1157692,I1157839);
or I_67899 (I1157870,I938134,I938146);
nor I_67900 (I1157887,I938131,I938143);
DFFARX1 I_67901 (I1157887,I3563,I1157497,I1157913,);
not I_67902 (I1157921,I1157913);
nor I_67903 (I1157483,I1157921,I1157726);
nand I_67904 (I1157952,I1157921,I1157571);
not I_67905 (I1157969,I938131);
nand I_67906 (I1157986,I1157969,I1157675);
nand I_67907 (I1158003,I1157921,I1157986);
nand I_67908 (I1157474,I1158003,I1157952);
nand I_67909 (I1157471,I1157986,I1157870);
not I_67910 (I1158075,I3570);
DFFARX1 I_67911 (I154693,I3563,I1158075,I1158101,);
and I_67912 (I1158109,I1158101,I154669);
DFFARX1 I_67913 (I1158109,I3563,I1158075,I1158058,);
DFFARX1 I_67914 (I154687,I3563,I1158075,I1158149,);
not I_67915 (I1158157,I154675);
not I_67916 (I1158174,I154672);
nand I_67917 (I1158191,I1158174,I1158157);
nor I_67918 (I1158046,I1158149,I1158191);
DFFARX1 I_67919 (I1158191,I3563,I1158075,I1158231,);
not I_67920 (I1158067,I1158231);
not I_67921 (I1158253,I154681);
nand I_67922 (I1158270,I1158174,I1158253);
DFFARX1 I_67923 (I1158270,I3563,I1158075,I1158296,);
not I_67924 (I1158304,I1158296);
not I_67925 (I1158321,I154672);
nand I_67926 (I1158338,I1158321,I154690);
and I_67927 (I1158355,I1158157,I1158338);
nor I_67928 (I1158372,I1158270,I1158355);
DFFARX1 I_67929 (I1158372,I3563,I1158075,I1158043,);
DFFARX1 I_67930 (I1158355,I3563,I1158075,I1158064,);
nor I_67931 (I1158417,I154672,I154684);
nor I_67932 (I1158055,I1158270,I1158417);
or I_67933 (I1158448,I154672,I154684);
nor I_67934 (I1158465,I154678,I154669);
DFFARX1 I_67935 (I1158465,I3563,I1158075,I1158491,);
not I_67936 (I1158499,I1158491);
nor I_67937 (I1158061,I1158499,I1158304);
nand I_67938 (I1158530,I1158499,I1158149);
not I_67939 (I1158547,I154678);
nand I_67940 (I1158564,I1158547,I1158253);
nand I_67941 (I1158581,I1158499,I1158564);
nand I_67942 (I1158052,I1158581,I1158530);
nand I_67943 (I1158049,I1158564,I1158448);
not I_67944 (I1158653,I3570);
DFFARX1 I_67945 (I791368,I3563,I1158653,I1158679,);
and I_67946 (I1158687,I1158679,I791356);
DFFARX1 I_67947 (I1158687,I3563,I1158653,I1158636,);
DFFARX1 I_67948 (I791359,I3563,I1158653,I1158727,);
not I_67949 (I1158735,I791353);
not I_67950 (I1158752,I791377);
nand I_67951 (I1158769,I1158752,I1158735);
nor I_67952 (I1158624,I1158727,I1158769);
DFFARX1 I_67953 (I1158769,I3563,I1158653,I1158809,);
not I_67954 (I1158645,I1158809);
not I_67955 (I1158831,I791365);
nand I_67956 (I1158848,I1158752,I1158831);
DFFARX1 I_67957 (I1158848,I3563,I1158653,I1158874,);
not I_67958 (I1158882,I1158874);
not I_67959 (I1158899,I791374);
nand I_67960 (I1158916,I1158899,I791371);
and I_67961 (I1158933,I1158735,I1158916);
nor I_67962 (I1158950,I1158848,I1158933);
DFFARX1 I_67963 (I1158950,I3563,I1158653,I1158621,);
DFFARX1 I_67964 (I1158933,I3563,I1158653,I1158642,);
nor I_67965 (I1158995,I791374,I791362);
nor I_67966 (I1158633,I1158848,I1158995);
or I_67967 (I1159026,I791374,I791362);
nor I_67968 (I1159043,I791353,I791356);
DFFARX1 I_67969 (I1159043,I3563,I1158653,I1159069,);
not I_67970 (I1159077,I1159069);
nor I_67971 (I1158639,I1159077,I1158882);
nand I_67972 (I1159108,I1159077,I1158727);
not I_67973 (I1159125,I791353);
nand I_67974 (I1159142,I1159125,I1158831);
nand I_67975 (I1159159,I1159077,I1159142);
nand I_67976 (I1158630,I1159159,I1159108);
nand I_67977 (I1158627,I1159142,I1159026);
not I_67978 (I1159231,I3570);
DFFARX1 I_67979 (I602362,I3563,I1159231,I1159257,);
and I_67980 (I1159265,I1159257,I602350);
DFFARX1 I_67981 (I1159265,I3563,I1159231,I1159214,);
DFFARX1 I_67982 (I602365,I3563,I1159231,I1159305,);
not I_67983 (I1159313,I602356);
not I_67984 (I1159330,I602347);
nand I_67985 (I1159347,I1159330,I1159313);
nor I_67986 (I1159202,I1159305,I1159347);
DFFARX1 I_67987 (I1159347,I3563,I1159231,I1159387,);
not I_67988 (I1159223,I1159387);
not I_67989 (I1159409,I602353);
nand I_67990 (I1159426,I1159330,I1159409);
DFFARX1 I_67991 (I1159426,I3563,I1159231,I1159452,);
not I_67992 (I1159460,I1159452);
not I_67993 (I1159477,I602368);
nand I_67994 (I1159494,I1159477,I602371);
and I_67995 (I1159511,I1159313,I1159494);
nor I_67996 (I1159528,I1159426,I1159511);
DFFARX1 I_67997 (I1159528,I3563,I1159231,I1159199,);
DFFARX1 I_67998 (I1159511,I3563,I1159231,I1159220,);
nor I_67999 (I1159573,I602368,I602347);
nor I_68000 (I1159211,I1159426,I1159573);
or I_68001 (I1159604,I602368,I602347);
nor I_68002 (I1159621,I602359,I602350);
DFFARX1 I_68003 (I1159621,I3563,I1159231,I1159647,);
not I_68004 (I1159655,I1159647);
nor I_68005 (I1159217,I1159655,I1159460);
nand I_68006 (I1159686,I1159655,I1159305);
not I_68007 (I1159703,I602359);
nand I_68008 (I1159720,I1159703,I1159409);
nand I_68009 (I1159737,I1159655,I1159720);
nand I_68010 (I1159208,I1159737,I1159686);
nand I_68011 (I1159205,I1159720,I1159604);
not I_68012 (I1159809,I3570);
DFFARX1 I_68013 (I54539,I3563,I1159809,I1159835,);
and I_68014 (I1159843,I1159835,I54542);
DFFARX1 I_68015 (I1159843,I3563,I1159809,I1159792,);
DFFARX1 I_68016 (I54542,I3563,I1159809,I1159883,);
not I_68017 (I1159891,I54545);
not I_68018 (I1159908,I54560);
nand I_68019 (I1159925,I1159908,I1159891);
nor I_68020 (I1159780,I1159883,I1159925);
DFFARX1 I_68021 (I1159925,I3563,I1159809,I1159965,);
not I_68022 (I1159801,I1159965);
not I_68023 (I1159987,I54554);
nand I_68024 (I1160004,I1159908,I1159987);
DFFARX1 I_68025 (I1160004,I3563,I1159809,I1160030,);
not I_68026 (I1160038,I1160030);
not I_68027 (I1160055,I54557);
nand I_68028 (I1160072,I1160055,I54539);
and I_68029 (I1160089,I1159891,I1160072);
nor I_68030 (I1160106,I1160004,I1160089);
DFFARX1 I_68031 (I1160106,I3563,I1159809,I1159777,);
DFFARX1 I_68032 (I1160089,I3563,I1159809,I1159798,);
nor I_68033 (I1160151,I54557,I54551);
nor I_68034 (I1159789,I1160004,I1160151);
or I_68035 (I1160182,I54557,I54551);
nor I_68036 (I1160199,I54548,I54563);
DFFARX1 I_68037 (I1160199,I3563,I1159809,I1160225,);
not I_68038 (I1160233,I1160225);
nor I_68039 (I1159795,I1160233,I1160038);
nand I_68040 (I1160264,I1160233,I1159883);
not I_68041 (I1160281,I54548);
nand I_68042 (I1160298,I1160281,I1159987);
nand I_68043 (I1160315,I1160233,I1160298);
nand I_68044 (I1159786,I1160315,I1160264);
nand I_68045 (I1159783,I1160298,I1160182);
not I_68046 (I1160387,I3570);
DFFARX1 I_68047 (I911189,I3563,I1160387,I1160413,);
and I_68048 (I1160421,I1160413,I911195);
DFFARX1 I_68049 (I1160421,I3563,I1160387,I1160370,);
DFFARX1 I_68050 (I911201,I3563,I1160387,I1160461,);
not I_68051 (I1160469,I911186);
not I_68052 (I1160486,I911186);
nand I_68053 (I1160503,I1160486,I1160469);
nor I_68054 (I1160358,I1160461,I1160503);
DFFARX1 I_68055 (I1160503,I3563,I1160387,I1160543,);
not I_68056 (I1160379,I1160543);
not I_68057 (I1160565,I911204);
nand I_68058 (I1160582,I1160486,I1160565);
DFFARX1 I_68059 (I1160582,I3563,I1160387,I1160608,);
not I_68060 (I1160616,I1160608);
not I_68061 (I1160633,I911198);
nand I_68062 (I1160650,I1160633,I911189);
and I_68063 (I1160667,I1160469,I1160650);
nor I_68064 (I1160684,I1160582,I1160667);
DFFARX1 I_68065 (I1160684,I3563,I1160387,I1160355,);
DFFARX1 I_68066 (I1160667,I3563,I1160387,I1160376,);
nor I_68067 (I1160729,I911198,I911207);
nor I_68068 (I1160367,I1160582,I1160729);
or I_68069 (I1160760,I911198,I911207);
nor I_68070 (I1160777,I911192,I911192);
DFFARX1 I_68071 (I1160777,I3563,I1160387,I1160803,);
not I_68072 (I1160811,I1160803);
nor I_68073 (I1160373,I1160811,I1160616);
nand I_68074 (I1160842,I1160811,I1160461);
not I_68075 (I1160859,I911192);
nand I_68076 (I1160876,I1160859,I1160565);
nand I_68077 (I1160893,I1160811,I1160876);
nand I_68078 (I1160364,I1160893,I1160842);
nand I_68079 (I1160361,I1160876,I1160760);
not I_68080 (I1160965,I3570);
DFFARX1 I_68081 (I1276894,I3563,I1160965,I1160991,);
and I_68082 (I1160999,I1160991,I1276888);
DFFARX1 I_68083 (I1160999,I3563,I1160965,I1160948,);
DFFARX1 I_68084 (I1276873,I3563,I1160965,I1161039,);
not I_68085 (I1161047,I1276879);
not I_68086 (I1161064,I1276891);
nand I_68087 (I1161081,I1161064,I1161047);
nor I_68088 (I1160936,I1161039,I1161081);
DFFARX1 I_68089 (I1161081,I3563,I1160965,I1161121,);
not I_68090 (I1160957,I1161121);
not I_68091 (I1161143,I1276873);
nand I_68092 (I1161160,I1161064,I1161143);
DFFARX1 I_68093 (I1161160,I3563,I1160965,I1161186,);
not I_68094 (I1161194,I1161186);
not I_68095 (I1161211,I1276897);
nand I_68096 (I1161228,I1161211,I1276885);
and I_68097 (I1161245,I1161047,I1161228);
nor I_68098 (I1161262,I1161160,I1161245);
DFFARX1 I_68099 (I1161262,I3563,I1160965,I1160933,);
DFFARX1 I_68100 (I1161245,I3563,I1160965,I1160954,);
nor I_68101 (I1161307,I1276897,I1276876);
nor I_68102 (I1160945,I1161160,I1161307);
or I_68103 (I1161338,I1276897,I1276876);
nor I_68104 (I1161355,I1276882,I1276876);
DFFARX1 I_68105 (I1161355,I3563,I1160965,I1161381,);
not I_68106 (I1161389,I1161381);
nor I_68107 (I1160951,I1161389,I1161194);
nand I_68108 (I1161420,I1161389,I1161039);
not I_68109 (I1161437,I1276882);
nand I_68110 (I1161454,I1161437,I1161143);
nand I_68111 (I1161471,I1161389,I1161454);
nand I_68112 (I1160942,I1161471,I1161420);
nand I_68113 (I1160939,I1161454,I1161338);
not I_68114 (I1161543,I3570);
DFFARX1 I_68115 (I273788,I3563,I1161543,I1161569,);
and I_68116 (I1161577,I1161569,I273791);
DFFARX1 I_68117 (I1161577,I3563,I1161543,I1161526,);
DFFARX1 I_68118 (I273791,I3563,I1161543,I1161617,);
not I_68119 (I1161625,I273806);
not I_68120 (I1161642,I273812);
nand I_68121 (I1161659,I1161642,I1161625);
nor I_68122 (I1161514,I1161617,I1161659);
DFFARX1 I_68123 (I1161659,I3563,I1161543,I1161699,);
not I_68124 (I1161535,I1161699);
not I_68125 (I1161721,I273800);
nand I_68126 (I1161738,I1161642,I1161721);
DFFARX1 I_68127 (I1161738,I3563,I1161543,I1161764,);
not I_68128 (I1161772,I1161764);
not I_68129 (I1161789,I273797);
nand I_68130 (I1161806,I1161789,I273794);
and I_68131 (I1161823,I1161625,I1161806);
nor I_68132 (I1161840,I1161738,I1161823);
DFFARX1 I_68133 (I1161840,I3563,I1161543,I1161511,);
DFFARX1 I_68134 (I1161823,I3563,I1161543,I1161532,);
nor I_68135 (I1161885,I273797,I273788);
nor I_68136 (I1161523,I1161738,I1161885);
or I_68137 (I1161916,I273797,I273788);
nor I_68138 (I1161933,I273803,I273809);
DFFARX1 I_68139 (I1161933,I3563,I1161543,I1161959,);
not I_68140 (I1161967,I1161959);
nor I_68141 (I1161529,I1161967,I1161772);
nand I_68142 (I1161998,I1161967,I1161617);
not I_68143 (I1162015,I273803);
nand I_68144 (I1162032,I1162015,I1161721);
nand I_68145 (I1162049,I1161967,I1162032);
nand I_68146 (I1161520,I1162049,I1161998);
nand I_68147 (I1161517,I1162032,I1161916);
not I_68148 (I1162121,I3570);
DFFARX1 I_68149 (I164903,I3563,I1162121,I1162147,);
and I_68150 (I1162155,I1162147,I164927);
DFFARX1 I_68151 (I1162155,I3563,I1162121,I1162104,);
DFFARX1 I_68152 (I164903,I3563,I1162121,I1162195,);
not I_68153 (I1162203,I164921);
not I_68154 (I1162220,I164906);
nand I_68155 (I1162237,I1162220,I1162203);
nor I_68156 (I1162092,I1162195,I1162237);
DFFARX1 I_68157 (I1162237,I3563,I1162121,I1162277,);
not I_68158 (I1162113,I1162277);
not I_68159 (I1162299,I164915);
nand I_68160 (I1162316,I1162220,I1162299);
DFFARX1 I_68161 (I1162316,I3563,I1162121,I1162342,);
not I_68162 (I1162350,I1162342);
not I_68163 (I1162367,I164912);
nand I_68164 (I1162384,I1162367,I164909);
and I_68165 (I1162401,I1162203,I1162384);
nor I_68166 (I1162418,I1162316,I1162401);
DFFARX1 I_68167 (I1162418,I3563,I1162121,I1162089,);
DFFARX1 I_68168 (I1162401,I3563,I1162121,I1162110,);
nor I_68169 (I1162463,I164912,I164918);
nor I_68170 (I1162101,I1162316,I1162463);
or I_68171 (I1162494,I164912,I164918);
nor I_68172 (I1162511,I164924,I164930);
DFFARX1 I_68173 (I1162511,I3563,I1162121,I1162537,);
not I_68174 (I1162545,I1162537);
nor I_68175 (I1162107,I1162545,I1162350);
nand I_68176 (I1162576,I1162545,I1162195);
not I_68177 (I1162593,I164924);
nand I_68178 (I1162610,I1162593,I1162299);
nand I_68179 (I1162627,I1162545,I1162610);
nand I_68180 (I1162098,I1162627,I1162576);
nand I_68181 (I1162095,I1162610,I1162494);
not I_68182 (I1162699,I3570);
DFFARX1 I_68183 (I817910,I3563,I1162699,I1162725,);
and I_68184 (I1162733,I1162725,I817916);
DFFARX1 I_68185 (I1162733,I3563,I1162699,I1162682,);
DFFARX1 I_68186 (I817922,I3563,I1162699,I1162773,);
not I_68187 (I1162781,I817907);
not I_68188 (I1162798,I817907);
nand I_68189 (I1162815,I1162798,I1162781);
nor I_68190 (I1162670,I1162773,I1162815);
DFFARX1 I_68191 (I1162815,I3563,I1162699,I1162855,);
not I_68192 (I1162691,I1162855);
not I_68193 (I1162877,I817925);
nand I_68194 (I1162894,I1162798,I1162877);
DFFARX1 I_68195 (I1162894,I3563,I1162699,I1162920,);
not I_68196 (I1162928,I1162920);
not I_68197 (I1162945,I817919);
nand I_68198 (I1162962,I1162945,I817910);
and I_68199 (I1162979,I1162781,I1162962);
nor I_68200 (I1162996,I1162894,I1162979);
DFFARX1 I_68201 (I1162996,I3563,I1162699,I1162667,);
DFFARX1 I_68202 (I1162979,I3563,I1162699,I1162688,);
nor I_68203 (I1163041,I817919,I817928);
nor I_68204 (I1162679,I1162894,I1163041);
or I_68205 (I1163072,I817919,I817928);
nor I_68206 (I1163089,I817913,I817913);
DFFARX1 I_68207 (I1163089,I3563,I1162699,I1163115,);
not I_68208 (I1163123,I1163115);
nor I_68209 (I1162685,I1163123,I1162928);
nand I_68210 (I1163154,I1163123,I1162773);
not I_68211 (I1163171,I817913);
nand I_68212 (I1163188,I1163171,I1162877);
nand I_68213 (I1163205,I1163123,I1163188);
nand I_68214 (I1162676,I1163205,I1163154);
nand I_68215 (I1162673,I1163188,I1163072);
not I_68216 (I1163277,I3570);
DFFARX1 I_68217 (I262483,I3563,I1163277,I1163303,);
and I_68218 (I1163311,I1163303,I262486);
DFFARX1 I_68219 (I1163311,I3563,I1163277,I1163260,);
DFFARX1 I_68220 (I262486,I3563,I1163277,I1163351,);
not I_68221 (I1163359,I262501);
not I_68222 (I1163376,I262507);
nand I_68223 (I1163393,I1163376,I1163359);
nor I_68224 (I1163248,I1163351,I1163393);
DFFARX1 I_68225 (I1163393,I3563,I1163277,I1163433,);
not I_68226 (I1163269,I1163433);
not I_68227 (I1163455,I262495);
nand I_68228 (I1163472,I1163376,I1163455);
DFFARX1 I_68229 (I1163472,I3563,I1163277,I1163498,);
not I_68230 (I1163506,I1163498);
not I_68231 (I1163523,I262492);
nand I_68232 (I1163540,I1163523,I262489);
and I_68233 (I1163557,I1163359,I1163540);
nor I_68234 (I1163574,I1163472,I1163557);
DFFARX1 I_68235 (I1163574,I3563,I1163277,I1163245,);
DFFARX1 I_68236 (I1163557,I3563,I1163277,I1163266,);
nor I_68237 (I1163619,I262492,I262483);
nor I_68238 (I1163257,I1163472,I1163619);
or I_68239 (I1163650,I262492,I262483);
nor I_68240 (I1163667,I262498,I262504);
DFFARX1 I_68241 (I1163667,I3563,I1163277,I1163693,);
not I_68242 (I1163701,I1163693);
nor I_68243 (I1163263,I1163701,I1163506);
nand I_68244 (I1163732,I1163701,I1163351);
not I_68245 (I1163749,I262498);
nand I_68246 (I1163766,I1163749,I1163455);
nand I_68247 (I1163783,I1163701,I1163766);
nand I_68248 (I1163254,I1163783,I1163732);
nand I_68249 (I1163251,I1163766,I1163650);
not I_68250 (I1163855,I3570);
DFFARX1 I_68251 (I1388675,I3563,I1163855,I1163881,);
and I_68252 (I1163889,I1163881,I1388657);
DFFARX1 I_68253 (I1163889,I3563,I1163855,I1163838,);
DFFARX1 I_68254 (I1388648,I3563,I1163855,I1163929,);
not I_68255 (I1163937,I1388663);
not I_68256 (I1163954,I1388651);
nand I_68257 (I1163971,I1163954,I1163937);
nor I_68258 (I1163826,I1163929,I1163971);
DFFARX1 I_68259 (I1163971,I3563,I1163855,I1164011,);
not I_68260 (I1163847,I1164011);
not I_68261 (I1164033,I1388660);
nand I_68262 (I1164050,I1163954,I1164033);
DFFARX1 I_68263 (I1164050,I3563,I1163855,I1164076,);
not I_68264 (I1164084,I1164076);
not I_68265 (I1164101,I1388669);
nand I_68266 (I1164118,I1164101,I1388648);
and I_68267 (I1164135,I1163937,I1164118);
nor I_68268 (I1164152,I1164050,I1164135);
DFFARX1 I_68269 (I1164152,I3563,I1163855,I1163823,);
DFFARX1 I_68270 (I1164135,I3563,I1163855,I1163844,);
nor I_68271 (I1164197,I1388669,I1388672);
nor I_68272 (I1163835,I1164050,I1164197);
or I_68273 (I1164228,I1388669,I1388672);
nor I_68274 (I1164245,I1388666,I1388654);
DFFARX1 I_68275 (I1164245,I3563,I1163855,I1164271,);
not I_68276 (I1164279,I1164271);
nor I_68277 (I1163841,I1164279,I1164084);
nand I_68278 (I1164310,I1164279,I1163929);
not I_68279 (I1164327,I1388666);
nand I_68280 (I1164344,I1164327,I1164033);
nand I_68281 (I1164361,I1164279,I1164344);
nand I_68282 (I1163832,I1164361,I1164310);
nand I_68283 (I1163829,I1164344,I1164228);
not I_68284 (I1164433,I3570);
DFFARX1 I_68285 (I1255678,I3563,I1164433,I1164459,);
and I_68286 (I1164467,I1164459,I1255672);
DFFARX1 I_68287 (I1164467,I3563,I1164433,I1164416,);
DFFARX1 I_68288 (I1255657,I3563,I1164433,I1164507,);
not I_68289 (I1164515,I1255663);
not I_68290 (I1164532,I1255675);
nand I_68291 (I1164549,I1164532,I1164515);
nor I_68292 (I1164404,I1164507,I1164549);
DFFARX1 I_68293 (I1164549,I3563,I1164433,I1164589,);
not I_68294 (I1164425,I1164589);
not I_68295 (I1164611,I1255657);
nand I_68296 (I1164628,I1164532,I1164611);
DFFARX1 I_68297 (I1164628,I3563,I1164433,I1164654,);
not I_68298 (I1164662,I1164654);
not I_68299 (I1164679,I1255681);
nand I_68300 (I1164696,I1164679,I1255669);
and I_68301 (I1164713,I1164515,I1164696);
nor I_68302 (I1164730,I1164628,I1164713);
DFFARX1 I_68303 (I1164730,I3563,I1164433,I1164401,);
DFFARX1 I_68304 (I1164713,I3563,I1164433,I1164422,);
nor I_68305 (I1164775,I1255681,I1255660);
nor I_68306 (I1164413,I1164628,I1164775);
or I_68307 (I1164806,I1255681,I1255660);
nor I_68308 (I1164823,I1255666,I1255660);
DFFARX1 I_68309 (I1164823,I3563,I1164433,I1164849,);
not I_68310 (I1164857,I1164849);
nor I_68311 (I1164419,I1164857,I1164662);
nand I_68312 (I1164888,I1164857,I1164507);
not I_68313 (I1164905,I1255666);
nand I_68314 (I1164922,I1164905,I1164611);
nand I_68315 (I1164939,I1164857,I1164922);
nand I_68316 (I1164410,I1164939,I1164888);
nand I_68317 (I1164407,I1164922,I1164806);
not I_68318 (I1165011,I3570);
DFFARX1 I_68319 (I706402,I3563,I1165011,I1165037,);
and I_68320 (I1165045,I1165037,I706390);
DFFARX1 I_68321 (I1165045,I3563,I1165011,I1164994,);
DFFARX1 I_68322 (I706393,I3563,I1165011,I1165085,);
not I_68323 (I1165093,I706387);
not I_68324 (I1165110,I706411);
nand I_68325 (I1165127,I1165110,I1165093);
nor I_68326 (I1164982,I1165085,I1165127);
DFFARX1 I_68327 (I1165127,I3563,I1165011,I1165167,);
not I_68328 (I1165003,I1165167);
not I_68329 (I1165189,I706399);
nand I_68330 (I1165206,I1165110,I1165189);
DFFARX1 I_68331 (I1165206,I3563,I1165011,I1165232,);
not I_68332 (I1165240,I1165232);
not I_68333 (I1165257,I706408);
nand I_68334 (I1165274,I1165257,I706405);
and I_68335 (I1165291,I1165093,I1165274);
nor I_68336 (I1165308,I1165206,I1165291);
DFFARX1 I_68337 (I1165308,I3563,I1165011,I1164979,);
DFFARX1 I_68338 (I1165291,I3563,I1165011,I1165000,);
nor I_68339 (I1165353,I706408,I706396);
nor I_68340 (I1164991,I1165206,I1165353);
or I_68341 (I1165384,I706408,I706396);
nor I_68342 (I1165401,I706387,I706390);
DFFARX1 I_68343 (I1165401,I3563,I1165011,I1165427,);
not I_68344 (I1165435,I1165427);
nor I_68345 (I1164997,I1165435,I1165240);
nand I_68346 (I1165466,I1165435,I1165085);
not I_68347 (I1165483,I706387);
nand I_68348 (I1165500,I1165483,I1165189);
nand I_68349 (I1165517,I1165435,I1165500);
nand I_68350 (I1164988,I1165517,I1165466);
nand I_68351 (I1164985,I1165500,I1165384);
not I_68352 (I1165589,I3570);
DFFARX1 I_68353 (I885366,I3563,I1165589,I1165615,);
and I_68354 (I1165623,I1165615,I885372);
DFFARX1 I_68355 (I1165623,I3563,I1165589,I1165572,);
DFFARX1 I_68356 (I885378,I3563,I1165589,I1165663,);
not I_68357 (I1165671,I885363);
not I_68358 (I1165688,I885363);
nand I_68359 (I1165705,I1165688,I1165671);
nor I_68360 (I1165560,I1165663,I1165705);
DFFARX1 I_68361 (I1165705,I3563,I1165589,I1165745,);
not I_68362 (I1165581,I1165745);
not I_68363 (I1165767,I885381);
nand I_68364 (I1165784,I1165688,I1165767);
DFFARX1 I_68365 (I1165784,I3563,I1165589,I1165810,);
not I_68366 (I1165818,I1165810);
not I_68367 (I1165835,I885375);
nand I_68368 (I1165852,I1165835,I885366);
and I_68369 (I1165869,I1165671,I1165852);
nor I_68370 (I1165886,I1165784,I1165869);
DFFARX1 I_68371 (I1165886,I3563,I1165589,I1165557,);
DFFARX1 I_68372 (I1165869,I3563,I1165589,I1165578,);
nor I_68373 (I1165931,I885375,I885384);
nor I_68374 (I1165569,I1165784,I1165931);
or I_68375 (I1165962,I885375,I885384);
nor I_68376 (I1165979,I885369,I885369);
DFFARX1 I_68377 (I1165979,I3563,I1165589,I1166005,);
not I_68378 (I1166013,I1166005);
nor I_68379 (I1165575,I1166013,I1165818);
nand I_68380 (I1166044,I1166013,I1165663);
not I_68381 (I1166061,I885369);
nand I_68382 (I1166078,I1166061,I1165767);
nand I_68383 (I1166095,I1166013,I1166078);
nand I_68384 (I1165566,I1166095,I1166044);
nand I_68385 (I1165563,I1166078,I1165962);
not I_68386 (I1166167,I3570);
DFFARX1 I_68387 (I550704,I3563,I1166167,I1166193,);
and I_68388 (I1166201,I1166193,I550719);
DFFARX1 I_68389 (I1166201,I3563,I1166167,I1166150,);
DFFARX1 I_68390 (I550710,I3563,I1166167,I1166241,);
not I_68391 (I1166249,I550704);
not I_68392 (I1166266,I550722);
nand I_68393 (I1166283,I1166266,I1166249);
nor I_68394 (I1166138,I1166241,I1166283);
DFFARX1 I_68395 (I1166283,I3563,I1166167,I1166323,);
not I_68396 (I1166159,I1166323);
not I_68397 (I1166345,I550713);
nand I_68398 (I1166362,I1166266,I1166345);
DFFARX1 I_68399 (I1166362,I3563,I1166167,I1166388,);
not I_68400 (I1166396,I1166388);
not I_68401 (I1166413,I550725);
nand I_68402 (I1166430,I1166413,I550701);
and I_68403 (I1166447,I1166249,I1166430);
nor I_68404 (I1166464,I1166362,I1166447);
DFFARX1 I_68405 (I1166464,I3563,I1166167,I1166135,);
DFFARX1 I_68406 (I1166447,I3563,I1166167,I1166156,);
nor I_68407 (I1166509,I550725,I550701);
nor I_68408 (I1166147,I1166362,I1166509);
or I_68409 (I1166540,I550725,I550701);
nor I_68410 (I1166557,I550707,I550716);
DFFARX1 I_68411 (I1166557,I3563,I1166167,I1166583,);
not I_68412 (I1166591,I1166583);
nor I_68413 (I1166153,I1166591,I1166396);
nand I_68414 (I1166622,I1166591,I1166241);
not I_68415 (I1166639,I550707);
nand I_68416 (I1166656,I1166639,I1166345);
nand I_68417 (I1166673,I1166591,I1166656);
nand I_68418 (I1166144,I1166673,I1166622);
nand I_68419 (I1166141,I1166656,I1166540);
not I_68420 (I1166745,I3570);
DFFARX1 I_68421 (I871664,I3563,I1166745,I1166771,);
and I_68422 (I1166779,I1166771,I871670);
DFFARX1 I_68423 (I1166779,I3563,I1166745,I1166728,);
DFFARX1 I_68424 (I871676,I3563,I1166745,I1166819,);
not I_68425 (I1166827,I871661);
not I_68426 (I1166844,I871661);
nand I_68427 (I1166861,I1166844,I1166827);
nor I_68428 (I1166716,I1166819,I1166861);
DFFARX1 I_68429 (I1166861,I3563,I1166745,I1166901,);
not I_68430 (I1166737,I1166901);
not I_68431 (I1166923,I871679);
nand I_68432 (I1166940,I1166844,I1166923);
DFFARX1 I_68433 (I1166940,I3563,I1166745,I1166966,);
not I_68434 (I1166974,I1166966);
not I_68435 (I1166991,I871673);
nand I_68436 (I1167008,I1166991,I871664);
and I_68437 (I1167025,I1166827,I1167008);
nor I_68438 (I1167042,I1166940,I1167025);
DFFARX1 I_68439 (I1167042,I3563,I1166745,I1166713,);
DFFARX1 I_68440 (I1167025,I3563,I1166745,I1166734,);
nor I_68441 (I1167087,I871673,I871682);
nor I_68442 (I1166725,I1166940,I1167087);
or I_68443 (I1167118,I871673,I871682);
nor I_68444 (I1167135,I871667,I871667);
DFFARX1 I_68445 (I1167135,I3563,I1166745,I1167161,);
not I_68446 (I1167169,I1167161);
nor I_68447 (I1166731,I1167169,I1166974);
nand I_68448 (I1167200,I1167169,I1166819);
not I_68449 (I1167217,I871667);
nand I_68450 (I1167234,I1167217,I1166923);
nand I_68451 (I1167251,I1167169,I1167234);
nand I_68452 (I1166722,I1167251,I1167200);
nand I_68453 (I1166719,I1167234,I1167118);
not I_68454 (I1167323,I3570);
DFFARX1 I_68455 (I855327,I3563,I1167323,I1167349,);
and I_68456 (I1167357,I1167349,I855333);
DFFARX1 I_68457 (I1167357,I3563,I1167323,I1167306,);
DFFARX1 I_68458 (I855339,I3563,I1167323,I1167397,);
not I_68459 (I1167405,I855324);
not I_68460 (I1167422,I855324);
nand I_68461 (I1167439,I1167422,I1167405);
nor I_68462 (I1167294,I1167397,I1167439);
DFFARX1 I_68463 (I1167439,I3563,I1167323,I1167479,);
not I_68464 (I1167315,I1167479);
not I_68465 (I1167501,I855342);
nand I_68466 (I1167518,I1167422,I1167501);
DFFARX1 I_68467 (I1167518,I3563,I1167323,I1167544,);
not I_68468 (I1167552,I1167544);
not I_68469 (I1167569,I855336);
nand I_68470 (I1167586,I1167569,I855327);
and I_68471 (I1167603,I1167405,I1167586);
nor I_68472 (I1167620,I1167518,I1167603);
DFFARX1 I_68473 (I1167620,I3563,I1167323,I1167291,);
DFFARX1 I_68474 (I1167603,I3563,I1167323,I1167312,);
nor I_68475 (I1167665,I855336,I855345);
nor I_68476 (I1167303,I1167518,I1167665);
or I_68477 (I1167696,I855336,I855345);
nor I_68478 (I1167713,I855330,I855330);
DFFARX1 I_68479 (I1167713,I3563,I1167323,I1167739,);
not I_68480 (I1167747,I1167739);
nor I_68481 (I1167309,I1167747,I1167552);
nand I_68482 (I1167778,I1167747,I1167397);
not I_68483 (I1167795,I855330);
nand I_68484 (I1167812,I1167795,I1167501);
nand I_68485 (I1167829,I1167747,I1167812);
nand I_68486 (I1167300,I1167829,I1167778);
nand I_68487 (I1167297,I1167812,I1167696);
not I_68488 (I1167901,I3570);
DFFARX1 I_68489 (I500738,I3563,I1167901,I1167927,);
and I_68490 (I1167935,I1167927,I500753);
DFFARX1 I_68491 (I1167935,I3563,I1167901,I1167884,);
DFFARX1 I_68492 (I500756,I3563,I1167901,I1167975,);
not I_68493 (I1167983,I500750);
not I_68494 (I1168000,I500765);
nand I_68495 (I1168017,I1168000,I1167983);
nor I_68496 (I1167872,I1167975,I1168017);
DFFARX1 I_68497 (I1168017,I3563,I1167901,I1168057,);
not I_68498 (I1167893,I1168057);
not I_68499 (I1168079,I500741);
nand I_68500 (I1168096,I1168000,I1168079);
DFFARX1 I_68501 (I1168096,I3563,I1167901,I1168122,);
not I_68502 (I1168130,I1168122);
not I_68503 (I1168147,I500744);
nand I_68504 (I1168164,I1168147,I500738);
and I_68505 (I1168181,I1167983,I1168164);
nor I_68506 (I1168198,I1168096,I1168181);
DFFARX1 I_68507 (I1168198,I3563,I1167901,I1167869,);
DFFARX1 I_68508 (I1168181,I3563,I1167901,I1167890,);
nor I_68509 (I1168243,I500744,I500747);
nor I_68510 (I1167881,I1168096,I1168243);
or I_68511 (I1168274,I500744,I500747);
nor I_68512 (I1168291,I500762,I500759);
DFFARX1 I_68513 (I1168291,I3563,I1167901,I1168317,);
not I_68514 (I1168325,I1168317);
nor I_68515 (I1167887,I1168325,I1168130);
nand I_68516 (I1168356,I1168325,I1167975);
not I_68517 (I1168373,I500762);
nand I_68518 (I1168390,I1168373,I1168079);
nand I_68519 (I1168407,I1168325,I1168390);
nand I_68520 (I1167878,I1168407,I1168356);
nand I_68521 (I1167875,I1168390,I1168274);
not I_68522 (I1168479,I3570);
DFFARX1 I_68523 (I808708,I3563,I1168479,I1168505,);
and I_68524 (I1168513,I1168505,I808696);
DFFARX1 I_68525 (I1168513,I3563,I1168479,I1168462,);
DFFARX1 I_68526 (I808699,I3563,I1168479,I1168553,);
not I_68527 (I1168561,I808693);
not I_68528 (I1168578,I808717);
nand I_68529 (I1168595,I1168578,I1168561);
nor I_68530 (I1168450,I1168553,I1168595);
DFFARX1 I_68531 (I1168595,I3563,I1168479,I1168635,);
not I_68532 (I1168471,I1168635);
not I_68533 (I1168657,I808705);
nand I_68534 (I1168674,I1168578,I1168657);
DFFARX1 I_68535 (I1168674,I3563,I1168479,I1168700,);
not I_68536 (I1168708,I1168700);
not I_68537 (I1168725,I808714);
nand I_68538 (I1168742,I1168725,I808711);
and I_68539 (I1168759,I1168561,I1168742);
nor I_68540 (I1168776,I1168674,I1168759);
DFFARX1 I_68541 (I1168776,I3563,I1168479,I1168447,);
DFFARX1 I_68542 (I1168759,I3563,I1168479,I1168468,);
nor I_68543 (I1168821,I808714,I808702);
nor I_68544 (I1168459,I1168674,I1168821);
or I_68545 (I1168852,I808714,I808702);
nor I_68546 (I1168869,I808693,I808696);
DFFARX1 I_68547 (I1168869,I3563,I1168479,I1168895,);
not I_68548 (I1168903,I1168895);
nor I_68549 (I1168465,I1168903,I1168708);
nand I_68550 (I1168934,I1168903,I1168553);
not I_68551 (I1168951,I808693);
nand I_68552 (I1168968,I1168951,I1168657);
nand I_68553 (I1168985,I1168903,I1168968);
nand I_68554 (I1168456,I1168985,I1168934);
nand I_68555 (I1168453,I1168968,I1168852);
not I_68556 (I1169057,I3570);
DFFARX1 I_68557 (I757266,I3563,I1169057,I1169083,);
and I_68558 (I1169091,I1169083,I757254);
DFFARX1 I_68559 (I1169091,I3563,I1169057,I1169040,);
DFFARX1 I_68560 (I757257,I3563,I1169057,I1169131,);
not I_68561 (I1169139,I757251);
not I_68562 (I1169156,I757275);
nand I_68563 (I1169173,I1169156,I1169139);
nor I_68564 (I1169028,I1169131,I1169173);
DFFARX1 I_68565 (I1169173,I3563,I1169057,I1169213,);
not I_68566 (I1169049,I1169213);
not I_68567 (I1169235,I757263);
nand I_68568 (I1169252,I1169156,I1169235);
DFFARX1 I_68569 (I1169252,I3563,I1169057,I1169278,);
not I_68570 (I1169286,I1169278);
not I_68571 (I1169303,I757272);
nand I_68572 (I1169320,I1169303,I757269);
and I_68573 (I1169337,I1169139,I1169320);
nor I_68574 (I1169354,I1169252,I1169337);
DFFARX1 I_68575 (I1169354,I3563,I1169057,I1169025,);
DFFARX1 I_68576 (I1169337,I3563,I1169057,I1169046,);
nor I_68577 (I1169399,I757272,I757260);
nor I_68578 (I1169037,I1169252,I1169399);
or I_68579 (I1169430,I757272,I757260);
nor I_68580 (I1169447,I757251,I757254);
DFFARX1 I_68581 (I1169447,I3563,I1169057,I1169473,);
not I_68582 (I1169481,I1169473);
nor I_68583 (I1169043,I1169481,I1169286);
nand I_68584 (I1169512,I1169481,I1169131);
not I_68585 (I1169529,I757251);
nand I_68586 (I1169546,I1169529,I1169235);
nand I_68587 (I1169563,I1169481,I1169546);
nand I_68588 (I1169034,I1169563,I1169512);
nand I_68589 (I1169031,I1169546,I1169430);
not I_68590 (I1169635,I3570);
DFFARX1 I_68591 (I1245886,I3563,I1169635,I1169661,);
and I_68592 (I1169669,I1169661,I1245880);
DFFARX1 I_68593 (I1169669,I3563,I1169635,I1169618,);
DFFARX1 I_68594 (I1245865,I3563,I1169635,I1169709,);
not I_68595 (I1169717,I1245871);
not I_68596 (I1169734,I1245883);
nand I_68597 (I1169751,I1169734,I1169717);
nor I_68598 (I1169606,I1169709,I1169751);
DFFARX1 I_68599 (I1169751,I3563,I1169635,I1169791,);
not I_68600 (I1169627,I1169791);
not I_68601 (I1169813,I1245865);
nand I_68602 (I1169830,I1169734,I1169813);
DFFARX1 I_68603 (I1169830,I3563,I1169635,I1169856,);
not I_68604 (I1169864,I1169856);
not I_68605 (I1169881,I1245889);
nand I_68606 (I1169898,I1169881,I1245877);
and I_68607 (I1169915,I1169717,I1169898);
nor I_68608 (I1169932,I1169830,I1169915);
DFFARX1 I_68609 (I1169932,I3563,I1169635,I1169603,);
DFFARX1 I_68610 (I1169915,I3563,I1169635,I1169624,);
nor I_68611 (I1169977,I1245889,I1245868);
nor I_68612 (I1169615,I1169830,I1169977);
or I_68613 (I1170008,I1245889,I1245868);
nor I_68614 (I1170025,I1245874,I1245868);
DFFARX1 I_68615 (I1170025,I3563,I1169635,I1170051,);
not I_68616 (I1170059,I1170051);
nor I_68617 (I1169621,I1170059,I1169864);
nand I_68618 (I1170090,I1170059,I1169709);
not I_68619 (I1170107,I1245874);
nand I_68620 (I1170124,I1170107,I1169813);
nand I_68621 (I1170141,I1170059,I1170124);
nand I_68622 (I1169612,I1170141,I1170090);
nand I_68623 (I1169609,I1170124,I1170008);
not I_68624 (I1170213,I3570);
DFFARX1 I_68625 (I454498,I3563,I1170213,I1170239,);
and I_68626 (I1170247,I1170239,I454513);
DFFARX1 I_68627 (I1170247,I3563,I1170213,I1170196,);
DFFARX1 I_68628 (I454516,I3563,I1170213,I1170287,);
not I_68629 (I1170295,I454510);
not I_68630 (I1170312,I454525);
nand I_68631 (I1170329,I1170312,I1170295);
nor I_68632 (I1170184,I1170287,I1170329);
DFFARX1 I_68633 (I1170329,I3563,I1170213,I1170369,);
not I_68634 (I1170205,I1170369);
not I_68635 (I1170391,I454501);
nand I_68636 (I1170408,I1170312,I1170391);
DFFARX1 I_68637 (I1170408,I3563,I1170213,I1170434,);
not I_68638 (I1170442,I1170434);
not I_68639 (I1170459,I454504);
nand I_68640 (I1170476,I1170459,I454498);
and I_68641 (I1170493,I1170295,I1170476);
nor I_68642 (I1170510,I1170408,I1170493);
DFFARX1 I_68643 (I1170510,I3563,I1170213,I1170181,);
DFFARX1 I_68644 (I1170493,I3563,I1170213,I1170202,);
nor I_68645 (I1170555,I454504,I454507);
nor I_68646 (I1170193,I1170408,I1170555);
or I_68647 (I1170586,I454504,I454507);
nor I_68648 (I1170603,I454522,I454519);
DFFARX1 I_68649 (I1170603,I3563,I1170213,I1170629,);
not I_68650 (I1170637,I1170629);
nor I_68651 (I1170199,I1170637,I1170442);
nand I_68652 (I1170668,I1170637,I1170287);
not I_68653 (I1170685,I454522);
nand I_68654 (I1170702,I1170685,I1170391);
nand I_68655 (I1170719,I1170637,I1170702);
nand I_68656 (I1170190,I1170719,I1170668);
nand I_68657 (I1170187,I1170702,I1170586);
not I_68658 (I1170791,I3570);
DFFARX1 I_68659 (I344416,I3563,I1170791,I1170817,);
and I_68660 (I1170825,I1170817,I344401);
DFFARX1 I_68661 (I1170825,I3563,I1170791,I1170774,);
DFFARX1 I_68662 (I344407,I3563,I1170791,I1170865,);
not I_68663 (I1170873,I344389);
not I_68664 (I1170890,I344410);
nand I_68665 (I1170907,I1170890,I1170873);
nor I_68666 (I1170762,I1170865,I1170907);
DFFARX1 I_68667 (I1170907,I3563,I1170791,I1170947,);
not I_68668 (I1170783,I1170947);
not I_68669 (I1170969,I344413);
nand I_68670 (I1170986,I1170890,I1170969);
DFFARX1 I_68671 (I1170986,I3563,I1170791,I1171012,);
not I_68672 (I1171020,I1171012);
not I_68673 (I1171037,I344404);
nand I_68674 (I1171054,I1171037,I344392);
and I_68675 (I1171071,I1170873,I1171054);
nor I_68676 (I1171088,I1170986,I1171071);
DFFARX1 I_68677 (I1171088,I3563,I1170791,I1170759,);
DFFARX1 I_68678 (I1171071,I3563,I1170791,I1170780,);
nor I_68679 (I1171133,I344404,I344398);
nor I_68680 (I1170771,I1170986,I1171133);
or I_68681 (I1171164,I344404,I344398);
nor I_68682 (I1171181,I344395,I344389);
DFFARX1 I_68683 (I1171181,I3563,I1170791,I1171207,);
not I_68684 (I1171215,I1171207);
nor I_68685 (I1170777,I1171215,I1171020);
nand I_68686 (I1171246,I1171215,I1170865);
not I_68687 (I1171263,I344395);
nand I_68688 (I1171280,I1171263,I1170969);
nand I_68689 (I1171297,I1171215,I1171280);
nand I_68690 (I1170768,I1171297,I1171246);
nand I_68691 (I1170765,I1171280,I1171164);
not I_68692 (I1171369,I3570);
DFFARX1 I_68693 (I402386,I3563,I1171369,I1171395,);
and I_68694 (I1171403,I1171395,I402371);
DFFARX1 I_68695 (I1171403,I3563,I1171369,I1171352,);
DFFARX1 I_68696 (I402377,I3563,I1171369,I1171443,);
not I_68697 (I1171451,I402359);
not I_68698 (I1171468,I402380);
nand I_68699 (I1171485,I1171468,I1171451);
nor I_68700 (I1171340,I1171443,I1171485);
DFFARX1 I_68701 (I1171485,I3563,I1171369,I1171525,);
not I_68702 (I1171361,I1171525);
not I_68703 (I1171547,I402383);
nand I_68704 (I1171564,I1171468,I1171547);
DFFARX1 I_68705 (I1171564,I3563,I1171369,I1171590,);
not I_68706 (I1171598,I1171590);
not I_68707 (I1171615,I402374);
nand I_68708 (I1171632,I1171615,I402362);
and I_68709 (I1171649,I1171451,I1171632);
nor I_68710 (I1171666,I1171564,I1171649);
DFFARX1 I_68711 (I1171666,I3563,I1171369,I1171337,);
DFFARX1 I_68712 (I1171649,I3563,I1171369,I1171358,);
nor I_68713 (I1171711,I402374,I402368);
nor I_68714 (I1171349,I1171564,I1171711);
or I_68715 (I1171742,I402374,I402368);
nor I_68716 (I1171759,I402365,I402359);
DFFARX1 I_68717 (I1171759,I3563,I1171369,I1171785,);
not I_68718 (I1171793,I1171785);
nor I_68719 (I1171355,I1171793,I1171598);
nand I_68720 (I1171824,I1171793,I1171443);
not I_68721 (I1171841,I402365);
nand I_68722 (I1171858,I1171841,I1171547);
nand I_68723 (I1171875,I1171793,I1171858);
nand I_68724 (I1171346,I1171875,I1171824);
nand I_68725 (I1171343,I1171858,I1171742);
not I_68726 (I1171947,I3570);
DFFARX1 I_68727 (I2644,I3563,I1171947,I1171973,);
and I_68728 (I1171981,I1171973,I3420);
DFFARX1 I_68729 (I1171981,I3563,I1171947,I1171930,);
DFFARX1 I_68730 (I2708,I3563,I1171947,I1172021,);
not I_68731 (I1172029,I2860);
not I_68732 (I1172046,I2700);
nand I_68733 (I1172063,I1172046,I1172029);
nor I_68734 (I1171918,I1172021,I1172063);
DFFARX1 I_68735 (I1172063,I3563,I1171947,I1172103,);
not I_68736 (I1171939,I1172103);
not I_68737 (I1172125,I3380);
nand I_68738 (I1172142,I1172046,I1172125);
DFFARX1 I_68739 (I1172142,I3563,I1171947,I1172168,);
not I_68740 (I1172176,I1172168);
not I_68741 (I1172193,I2940);
nand I_68742 (I1172210,I1172193,I1756);
and I_68743 (I1172227,I1172029,I1172210);
nor I_68744 (I1172244,I1172142,I1172227);
DFFARX1 I_68745 (I1172244,I3563,I1171947,I1171915,);
DFFARX1 I_68746 (I1172227,I3563,I1171947,I1171936,);
nor I_68747 (I1172289,I2940,I1988);
nor I_68748 (I1171927,I1172142,I1172289);
or I_68749 (I1172320,I2940,I1988);
nor I_68750 (I1172337,I2876,I2124);
DFFARX1 I_68751 (I1172337,I3563,I1171947,I1172363,);
not I_68752 (I1172371,I1172363);
nor I_68753 (I1171933,I1172371,I1172176);
nand I_68754 (I1172402,I1172371,I1172021);
not I_68755 (I1172419,I2876);
nand I_68756 (I1172436,I1172419,I1172125);
nand I_68757 (I1172453,I1172371,I1172436);
nand I_68758 (I1171924,I1172453,I1172402);
nand I_68759 (I1171921,I1172436,I1172320);
not I_68760 (I1172525,I3570);
DFFARX1 I_68761 (I136248,I3563,I1172525,I1172551,);
and I_68762 (I1172559,I1172551,I136224);
DFFARX1 I_68763 (I1172559,I3563,I1172525,I1172508,);
DFFARX1 I_68764 (I136242,I3563,I1172525,I1172599,);
not I_68765 (I1172607,I136230);
not I_68766 (I1172624,I136227);
nand I_68767 (I1172641,I1172624,I1172607);
nor I_68768 (I1172496,I1172599,I1172641);
DFFARX1 I_68769 (I1172641,I3563,I1172525,I1172681,);
not I_68770 (I1172517,I1172681);
not I_68771 (I1172703,I136236);
nand I_68772 (I1172720,I1172624,I1172703);
DFFARX1 I_68773 (I1172720,I3563,I1172525,I1172746,);
not I_68774 (I1172754,I1172746);
not I_68775 (I1172771,I136227);
nand I_68776 (I1172788,I1172771,I136245);
and I_68777 (I1172805,I1172607,I1172788);
nor I_68778 (I1172822,I1172720,I1172805);
DFFARX1 I_68779 (I1172822,I3563,I1172525,I1172493,);
DFFARX1 I_68780 (I1172805,I3563,I1172525,I1172514,);
nor I_68781 (I1172867,I136227,I136239);
nor I_68782 (I1172505,I1172720,I1172867);
or I_68783 (I1172898,I136227,I136239);
nor I_68784 (I1172915,I136233,I136224);
DFFARX1 I_68785 (I1172915,I3563,I1172525,I1172941,);
not I_68786 (I1172949,I1172941);
nor I_68787 (I1172511,I1172949,I1172754);
nand I_68788 (I1172980,I1172949,I1172599);
not I_68789 (I1172997,I136233);
nand I_68790 (I1173014,I1172997,I1172703);
nand I_68791 (I1173031,I1172949,I1173014);
nand I_68792 (I1172502,I1173031,I1172980);
nand I_68793 (I1172499,I1173014,I1172898);
not I_68794 (I1173103,I3570);
DFFARX1 I_68795 (I864813,I3563,I1173103,I1173129,);
and I_68796 (I1173137,I1173129,I864819);
DFFARX1 I_68797 (I1173137,I3563,I1173103,I1173086,);
DFFARX1 I_68798 (I864825,I3563,I1173103,I1173177,);
not I_68799 (I1173185,I864810);
not I_68800 (I1173202,I864810);
nand I_68801 (I1173219,I1173202,I1173185);
nor I_68802 (I1173074,I1173177,I1173219);
DFFARX1 I_68803 (I1173219,I3563,I1173103,I1173259,);
not I_68804 (I1173095,I1173259);
not I_68805 (I1173281,I864828);
nand I_68806 (I1173298,I1173202,I1173281);
DFFARX1 I_68807 (I1173298,I3563,I1173103,I1173324,);
not I_68808 (I1173332,I1173324);
not I_68809 (I1173349,I864822);
nand I_68810 (I1173366,I1173349,I864813);
and I_68811 (I1173383,I1173185,I1173366);
nor I_68812 (I1173400,I1173298,I1173383);
DFFARX1 I_68813 (I1173400,I3563,I1173103,I1173071,);
DFFARX1 I_68814 (I1173383,I3563,I1173103,I1173092,);
nor I_68815 (I1173445,I864822,I864831);
nor I_68816 (I1173083,I1173298,I1173445);
or I_68817 (I1173476,I864822,I864831);
nor I_68818 (I1173493,I864816,I864816);
DFFARX1 I_68819 (I1173493,I3563,I1173103,I1173519,);
not I_68820 (I1173527,I1173519);
nor I_68821 (I1173089,I1173527,I1173332);
nand I_68822 (I1173558,I1173527,I1173177);
not I_68823 (I1173575,I864816);
nand I_68824 (I1173592,I1173575,I1173281);
nand I_68825 (I1173609,I1173527,I1173592);
nand I_68826 (I1173080,I1173609,I1173558);
nand I_68827 (I1173077,I1173592,I1173476);
not I_68828 (I1173681,I3570);
DFFARX1 I_68829 (I1089859,I3563,I1173681,I1173707,);
and I_68830 (I1173715,I1173707,I1089856);
DFFARX1 I_68831 (I1173715,I3563,I1173681,I1173664,);
DFFARX1 I_68832 (I1089862,I3563,I1173681,I1173755,);
not I_68833 (I1173763,I1089865);
not I_68834 (I1173780,I1089859);
nand I_68835 (I1173797,I1173780,I1173763);
nor I_68836 (I1173652,I1173755,I1173797);
DFFARX1 I_68837 (I1173797,I3563,I1173681,I1173837,);
not I_68838 (I1173673,I1173837);
not I_68839 (I1173859,I1089874);
nand I_68840 (I1173876,I1173780,I1173859);
DFFARX1 I_68841 (I1173876,I3563,I1173681,I1173902,);
not I_68842 (I1173910,I1173902);
not I_68843 (I1173927,I1089871);
nand I_68844 (I1173944,I1173927,I1089877);
and I_68845 (I1173961,I1173763,I1173944);
nor I_68846 (I1173978,I1173876,I1173961);
DFFARX1 I_68847 (I1173978,I3563,I1173681,I1173649,);
DFFARX1 I_68848 (I1173961,I3563,I1173681,I1173670,);
nor I_68849 (I1174023,I1089871,I1089856);
nor I_68850 (I1173661,I1173876,I1174023);
or I_68851 (I1174054,I1089871,I1089856);
nor I_68852 (I1174071,I1089868,I1089862);
DFFARX1 I_68853 (I1174071,I3563,I1173681,I1174097,);
not I_68854 (I1174105,I1174097);
nor I_68855 (I1173667,I1174105,I1173910);
nand I_68856 (I1174136,I1174105,I1173755);
not I_68857 (I1174153,I1089868);
nand I_68858 (I1174170,I1174153,I1173859);
nand I_68859 (I1174187,I1174105,I1174170);
nand I_68860 (I1173658,I1174187,I1174136);
nand I_68861 (I1173655,I1174170,I1174054);
not I_68862 (I1174259,I3570);
DFFARX1 I_68863 (I48215,I3563,I1174259,I1174285,);
and I_68864 (I1174293,I1174285,I48218);
DFFARX1 I_68865 (I1174293,I3563,I1174259,I1174242,);
DFFARX1 I_68866 (I48218,I3563,I1174259,I1174333,);
not I_68867 (I1174341,I48221);
not I_68868 (I1174358,I48236);
nand I_68869 (I1174375,I1174358,I1174341);
nor I_68870 (I1174230,I1174333,I1174375);
DFFARX1 I_68871 (I1174375,I3563,I1174259,I1174415,);
not I_68872 (I1174251,I1174415);
not I_68873 (I1174437,I48230);
nand I_68874 (I1174454,I1174358,I1174437);
DFFARX1 I_68875 (I1174454,I3563,I1174259,I1174480,);
not I_68876 (I1174488,I1174480);
not I_68877 (I1174505,I48233);
nand I_68878 (I1174522,I1174505,I48215);
and I_68879 (I1174539,I1174341,I1174522);
nor I_68880 (I1174556,I1174454,I1174539);
DFFARX1 I_68881 (I1174556,I3563,I1174259,I1174227,);
DFFARX1 I_68882 (I1174539,I3563,I1174259,I1174248,);
nor I_68883 (I1174601,I48233,I48227);
nor I_68884 (I1174239,I1174454,I1174601);
or I_68885 (I1174632,I48233,I48227);
nor I_68886 (I1174649,I48224,I48239);
DFFARX1 I_68887 (I1174649,I3563,I1174259,I1174675,);
not I_68888 (I1174683,I1174675);
nor I_68889 (I1174245,I1174683,I1174488);
nand I_68890 (I1174714,I1174683,I1174333);
not I_68891 (I1174731,I48224);
nand I_68892 (I1174748,I1174731,I1174437);
nand I_68893 (I1174765,I1174683,I1174748);
nand I_68894 (I1174236,I1174765,I1174714);
nand I_68895 (I1174233,I1174748,I1174632);
not I_68896 (I1174837,I3570);
DFFARX1 I_68897 (I267838,I3563,I1174837,I1174863,);
and I_68898 (I1174871,I1174863,I267841);
DFFARX1 I_68899 (I1174871,I3563,I1174837,I1174820,);
DFFARX1 I_68900 (I267841,I3563,I1174837,I1174911,);
not I_68901 (I1174919,I267856);
not I_68902 (I1174936,I267862);
nand I_68903 (I1174953,I1174936,I1174919);
nor I_68904 (I1174808,I1174911,I1174953);
DFFARX1 I_68905 (I1174953,I3563,I1174837,I1174993,);
not I_68906 (I1174829,I1174993);
not I_68907 (I1175015,I267850);
nand I_68908 (I1175032,I1174936,I1175015);
DFFARX1 I_68909 (I1175032,I3563,I1174837,I1175058,);
not I_68910 (I1175066,I1175058);
not I_68911 (I1175083,I267847);
nand I_68912 (I1175100,I1175083,I267844);
and I_68913 (I1175117,I1174919,I1175100);
nor I_68914 (I1175134,I1175032,I1175117);
DFFARX1 I_68915 (I1175134,I3563,I1174837,I1174805,);
DFFARX1 I_68916 (I1175117,I3563,I1174837,I1174826,);
nor I_68917 (I1175179,I267847,I267838);
nor I_68918 (I1174817,I1175032,I1175179);
or I_68919 (I1175210,I267847,I267838);
nor I_68920 (I1175227,I267853,I267859);
DFFARX1 I_68921 (I1175227,I3563,I1174837,I1175253,);
not I_68922 (I1175261,I1175253);
nor I_68923 (I1174823,I1175261,I1175066);
nand I_68924 (I1175292,I1175261,I1174911);
not I_68925 (I1175309,I267853);
nand I_68926 (I1175326,I1175309,I1175015);
nand I_68927 (I1175343,I1175261,I1175326);
nand I_68928 (I1174814,I1175343,I1175292);
nand I_68929 (I1174811,I1175326,I1175210);
not I_68930 (I1175415,I3570);
DFFARX1 I_68931 (I1010489,I3563,I1175415,I1175441,);
and I_68932 (I1175449,I1175441,I1010483);
DFFARX1 I_68933 (I1175449,I3563,I1175415,I1175398,);
DFFARX1 I_68934 (I1010501,I3563,I1175415,I1175489,);
not I_68935 (I1175497,I1010492);
not I_68936 (I1175514,I1010504);
nand I_68937 (I1175531,I1175514,I1175497);
nor I_68938 (I1175386,I1175489,I1175531);
DFFARX1 I_68939 (I1175531,I3563,I1175415,I1175571,);
not I_68940 (I1175407,I1175571);
not I_68941 (I1175593,I1010510);
nand I_68942 (I1175610,I1175514,I1175593);
DFFARX1 I_68943 (I1175610,I3563,I1175415,I1175636,);
not I_68944 (I1175644,I1175636);
not I_68945 (I1175661,I1010486);
nand I_68946 (I1175678,I1175661,I1010507);
and I_68947 (I1175695,I1175497,I1175678);
nor I_68948 (I1175712,I1175610,I1175695);
DFFARX1 I_68949 (I1175712,I3563,I1175415,I1175383,);
DFFARX1 I_68950 (I1175695,I3563,I1175415,I1175404,);
nor I_68951 (I1175757,I1010486,I1010498);
nor I_68952 (I1175395,I1175610,I1175757);
or I_68953 (I1175788,I1010486,I1010498);
nor I_68954 (I1175805,I1010483,I1010495);
DFFARX1 I_68955 (I1175805,I3563,I1175415,I1175831,);
not I_68956 (I1175839,I1175831);
nor I_68957 (I1175401,I1175839,I1175644);
nand I_68958 (I1175870,I1175839,I1175489);
not I_68959 (I1175887,I1010483);
nand I_68960 (I1175904,I1175887,I1175593);
nand I_68961 (I1175921,I1175839,I1175904);
nand I_68962 (I1175392,I1175921,I1175870);
nand I_68963 (I1175389,I1175904,I1175788);
not I_68964 (I1175993,I3570);
DFFARX1 I_68965 (I270218,I3563,I1175993,I1176019,);
and I_68966 (I1176027,I1176019,I270221);
DFFARX1 I_68967 (I1176027,I3563,I1175993,I1175976,);
DFFARX1 I_68968 (I270221,I3563,I1175993,I1176067,);
not I_68969 (I1176075,I270236);
not I_68970 (I1176092,I270242);
nand I_68971 (I1176109,I1176092,I1176075);
nor I_68972 (I1175964,I1176067,I1176109);
DFFARX1 I_68973 (I1176109,I3563,I1175993,I1176149,);
not I_68974 (I1175985,I1176149);
not I_68975 (I1176171,I270230);
nand I_68976 (I1176188,I1176092,I1176171);
DFFARX1 I_68977 (I1176188,I3563,I1175993,I1176214,);
not I_68978 (I1176222,I1176214);
not I_68979 (I1176239,I270227);
nand I_68980 (I1176256,I1176239,I270224);
and I_68981 (I1176273,I1176075,I1176256);
nor I_68982 (I1176290,I1176188,I1176273);
DFFARX1 I_68983 (I1176290,I3563,I1175993,I1175961,);
DFFARX1 I_68984 (I1176273,I3563,I1175993,I1175982,);
nor I_68985 (I1176335,I270227,I270218);
nor I_68986 (I1175973,I1176188,I1176335);
or I_68987 (I1176366,I270227,I270218);
nor I_68988 (I1176383,I270233,I270239);
DFFARX1 I_68989 (I1176383,I3563,I1175993,I1176409,);
not I_68990 (I1176417,I1176409);
nor I_68991 (I1175979,I1176417,I1176222);
nand I_68992 (I1176448,I1176417,I1176067);
not I_68993 (I1176465,I270233);
nand I_68994 (I1176482,I1176465,I1176171);
nand I_68995 (I1176499,I1176417,I1176482);
nand I_68996 (I1175970,I1176499,I1176448);
nand I_68997 (I1175967,I1176482,I1176366);
not I_68998 (I1176571,I3570);
DFFARX1 I_68999 (I250583,I3563,I1176571,I1176597,);
and I_69000 (I1176605,I1176597,I250586);
DFFARX1 I_69001 (I1176605,I3563,I1176571,I1176554,);
DFFARX1 I_69002 (I250586,I3563,I1176571,I1176645,);
not I_69003 (I1176653,I250601);
not I_69004 (I1176670,I250607);
nand I_69005 (I1176687,I1176670,I1176653);
nor I_69006 (I1176542,I1176645,I1176687);
DFFARX1 I_69007 (I1176687,I3563,I1176571,I1176727,);
not I_69008 (I1176563,I1176727);
not I_69009 (I1176749,I250595);
nand I_69010 (I1176766,I1176670,I1176749);
DFFARX1 I_69011 (I1176766,I3563,I1176571,I1176792,);
not I_69012 (I1176800,I1176792);
not I_69013 (I1176817,I250592);
nand I_69014 (I1176834,I1176817,I250589);
and I_69015 (I1176851,I1176653,I1176834);
nor I_69016 (I1176868,I1176766,I1176851);
DFFARX1 I_69017 (I1176868,I3563,I1176571,I1176539,);
DFFARX1 I_69018 (I1176851,I3563,I1176571,I1176560,);
nor I_69019 (I1176913,I250592,I250583);
nor I_69020 (I1176551,I1176766,I1176913);
or I_69021 (I1176944,I250592,I250583);
nor I_69022 (I1176961,I250598,I250604);
DFFARX1 I_69023 (I1176961,I3563,I1176571,I1176987,);
not I_69024 (I1176995,I1176987);
nor I_69025 (I1176557,I1176995,I1176800);
nand I_69026 (I1177026,I1176995,I1176645);
not I_69027 (I1177043,I250598);
nand I_69028 (I1177060,I1177043,I1176749);
nand I_69029 (I1177077,I1176995,I1177060);
nand I_69030 (I1176548,I1177077,I1177026);
nand I_69031 (I1176545,I1177060,I1176944);
not I_69032 (I1177149,I3570);
DFFARX1 I_69033 (I910135,I3563,I1177149,I1177175,);
and I_69034 (I1177183,I1177175,I910141);
DFFARX1 I_69035 (I1177183,I3563,I1177149,I1177132,);
DFFARX1 I_69036 (I910147,I3563,I1177149,I1177223,);
not I_69037 (I1177231,I910132);
not I_69038 (I1177248,I910132);
nand I_69039 (I1177265,I1177248,I1177231);
nor I_69040 (I1177120,I1177223,I1177265);
DFFARX1 I_69041 (I1177265,I3563,I1177149,I1177305,);
not I_69042 (I1177141,I1177305);
not I_69043 (I1177327,I910150);
nand I_69044 (I1177344,I1177248,I1177327);
DFFARX1 I_69045 (I1177344,I3563,I1177149,I1177370,);
not I_69046 (I1177378,I1177370);
not I_69047 (I1177395,I910144);
nand I_69048 (I1177412,I1177395,I910135);
and I_69049 (I1177429,I1177231,I1177412);
nor I_69050 (I1177446,I1177344,I1177429);
DFFARX1 I_69051 (I1177446,I3563,I1177149,I1177117,);
DFFARX1 I_69052 (I1177429,I3563,I1177149,I1177138,);
nor I_69053 (I1177491,I910144,I910153);
nor I_69054 (I1177129,I1177344,I1177491);
or I_69055 (I1177522,I910144,I910153);
nor I_69056 (I1177539,I910138,I910138);
DFFARX1 I_69057 (I1177539,I3563,I1177149,I1177565,);
not I_69058 (I1177573,I1177565);
nor I_69059 (I1177135,I1177573,I1177378);
nand I_69060 (I1177604,I1177573,I1177223);
not I_69061 (I1177621,I910138);
nand I_69062 (I1177638,I1177621,I1177327);
nand I_69063 (I1177655,I1177573,I1177638);
nand I_69064 (I1177126,I1177655,I1177604);
nand I_69065 (I1177123,I1177638,I1177522);
not I_69066 (I1177727,I3570);
DFFARX1 I_69067 (I963977,I3563,I1177727,I1177753,);
and I_69068 (I1177761,I1177753,I963971);
DFFARX1 I_69069 (I1177761,I3563,I1177727,I1177710,);
DFFARX1 I_69070 (I963989,I3563,I1177727,I1177801,);
not I_69071 (I1177809,I963980);
not I_69072 (I1177826,I963992);
nand I_69073 (I1177843,I1177826,I1177809);
nor I_69074 (I1177698,I1177801,I1177843);
DFFARX1 I_69075 (I1177843,I3563,I1177727,I1177883,);
not I_69076 (I1177719,I1177883);
not I_69077 (I1177905,I963998);
nand I_69078 (I1177922,I1177826,I1177905);
DFFARX1 I_69079 (I1177922,I3563,I1177727,I1177948,);
not I_69080 (I1177956,I1177948);
not I_69081 (I1177973,I963974);
nand I_69082 (I1177990,I1177973,I963995);
and I_69083 (I1178007,I1177809,I1177990);
nor I_69084 (I1178024,I1177922,I1178007);
DFFARX1 I_69085 (I1178024,I3563,I1177727,I1177695,);
DFFARX1 I_69086 (I1178007,I3563,I1177727,I1177716,);
nor I_69087 (I1178069,I963974,I963986);
nor I_69088 (I1177707,I1177922,I1178069);
or I_69089 (I1178100,I963974,I963986);
nor I_69090 (I1178117,I963971,I963983);
DFFARX1 I_69091 (I1178117,I3563,I1177727,I1178143,);
not I_69092 (I1178151,I1178143);
nor I_69093 (I1177713,I1178151,I1177956);
nand I_69094 (I1178182,I1178151,I1177801);
not I_69095 (I1178199,I963971);
nand I_69096 (I1178216,I1178199,I1177905);
nand I_69097 (I1178233,I1178151,I1178216);
nand I_69098 (I1177704,I1178233,I1178182);
nand I_69099 (I1177701,I1178216,I1178100);
not I_69100 (I1178305,I3570);
DFFARX1 I_69101 (I198818,I3563,I1178305,I1178331,);
and I_69102 (I1178339,I1178331,I198821);
DFFARX1 I_69103 (I1178339,I3563,I1178305,I1178288,);
DFFARX1 I_69104 (I198821,I3563,I1178305,I1178379,);
not I_69105 (I1178387,I198836);
not I_69106 (I1178404,I198842);
nand I_69107 (I1178421,I1178404,I1178387);
nor I_69108 (I1178276,I1178379,I1178421);
DFFARX1 I_69109 (I1178421,I3563,I1178305,I1178461,);
not I_69110 (I1178297,I1178461);
not I_69111 (I1178483,I198830);
nand I_69112 (I1178500,I1178404,I1178483);
DFFARX1 I_69113 (I1178500,I3563,I1178305,I1178526,);
not I_69114 (I1178534,I1178526);
not I_69115 (I1178551,I198827);
nand I_69116 (I1178568,I1178551,I198824);
and I_69117 (I1178585,I1178387,I1178568);
nor I_69118 (I1178602,I1178500,I1178585);
DFFARX1 I_69119 (I1178602,I3563,I1178305,I1178273,);
DFFARX1 I_69120 (I1178585,I3563,I1178305,I1178294,);
nor I_69121 (I1178647,I198827,I198818);
nor I_69122 (I1178285,I1178500,I1178647);
or I_69123 (I1178678,I198827,I198818);
nor I_69124 (I1178695,I198833,I198839);
DFFARX1 I_69125 (I1178695,I3563,I1178305,I1178721,);
not I_69126 (I1178729,I1178721);
nor I_69127 (I1178291,I1178729,I1178534);
nand I_69128 (I1178760,I1178729,I1178379);
not I_69129 (I1178777,I198833);
nand I_69130 (I1178794,I1178777,I1178483);
nand I_69131 (I1178811,I1178729,I1178794);
nand I_69132 (I1178282,I1178811,I1178760);
nand I_69133 (I1178279,I1178794,I1178678);
not I_69134 (I1178883,I3570);
DFFARX1 I_69135 (I905919,I3563,I1178883,I1178909,);
and I_69136 (I1178917,I1178909,I905925);
DFFARX1 I_69137 (I1178917,I3563,I1178883,I1178866,);
DFFARX1 I_69138 (I905931,I3563,I1178883,I1178957,);
not I_69139 (I1178965,I905916);
not I_69140 (I1178982,I905916);
nand I_69141 (I1178999,I1178982,I1178965);
nor I_69142 (I1178854,I1178957,I1178999);
DFFARX1 I_69143 (I1178999,I3563,I1178883,I1179039,);
not I_69144 (I1178875,I1179039);
not I_69145 (I1179061,I905934);
nand I_69146 (I1179078,I1178982,I1179061);
DFFARX1 I_69147 (I1179078,I3563,I1178883,I1179104,);
not I_69148 (I1179112,I1179104);
not I_69149 (I1179129,I905928);
nand I_69150 (I1179146,I1179129,I905919);
and I_69151 (I1179163,I1178965,I1179146);
nor I_69152 (I1179180,I1179078,I1179163);
DFFARX1 I_69153 (I1179180,I3563,I1178883,I1178851,);
DFFARX1 I_69154 (I1179163,I3563,I1178883,I1178872,);
nor I_69155 (I1179225,I905928,I905937);
nor I_69156 (I1178863,I1179078,I1179225);
or I_69157 (I1179256,I905928,I905937);
nor I_69158 (I1179273,I905922,I905922);
DFFARX1 I_69159 (I1179273,I3563,I1178883,I1179299,);
not I_69160 (I1179307,I1179299);
nor I_69161 (I1178869,I1179307,I1179112);
nand I_69162 (I1179338,I1179307,I1178957);
not I_69163 (I1179355,I905922);
nand I_69164 (I1179372,I1179355,I1179061);
nand I_69165 (I1179389,I1179307,I1179372);
nand I_69166 (I1178860,I1179389,I1179338);
nand I_69167 (I1178857,I1179372,I1179256);
not I_69168 (I1179461,I3570);
DFFARX1 I_69169 (I631840,I3563,I1179461,I1179487,);
and I_69170 (I1179495,I1179487,I631828);
DFFARX1 I_69171 (I1179495,I3563,I1179461,I1179444,);
DFFARX1 I_69172 (I631843,I3563,I1179461,I1179535,);
not I_69173 (I1179543,I631834);
not I_69174 (I1179560,I631825);
nand I_69175 (I1179577,I1179560,I1179543);
nor I_69176 (I1179432,I1179535,I1179577);
DFFARX1 I_69177 (I1179577,I3563,I1179461,I1179617,);
not I_69178 (I1179453,I1179617);
not I_69179 (I1179639,I631831);
nand I_69180 (I1179656,I1179560,I1179639);
DFFARX1 I_69181 (I1179656,I3563,I1179461,I1179682,);
not I_69182 (I1179690,I1179682);
not I_69183 (I1179707,I631846);
nand I_69184 (I1179724,I1179707,I631849);
and I_69185 (I1179741,I1179543,I1179724);
nor I_69186 (I1179758,I1179656,I1179741);
DFFARX1 I_69187 (I1179758,I3563,I1179461,I1179429,);
DFFARX1 I_69188 (I1179741,I3563,I1179461,I1179450,);
nor I_69189 (I1179803,I631846,I631825);
nor I_69190 (I1179441,I1179656,I1179803);
or I_69191 (I1179834,I631846,I631825);
nor I_69192 (I1179851,I631837,I631828);
DFFARX1 I_69193 (I1179851,I3563,I1179461,I1179877,);
not I_69194 (I1179885,I1179877);
nor I_69195 (I1179447,I1179885,I1179690);
nand I_69196 (I1179916,I1179885,I1179535);
not I_69197 (I1179933,I631837);
nand I_69198 (I1179950,I1179933,I1179639);
nand I_69199 (I1179967,I1179885,I1179950);
nand I_69200 (I1179438,I1179967,I1179916);
nand I_69201 (I1179435,I1179950,I1179834);
not I_69202 (I1180039,I3570);
DFFARX1 I_69203 (I1376775,I3563,I1180039,I1180065,);
and I_69204 (I1180073,I1180065,I1376757);
DFFARX1 I_69205 (I1180073,I3563,I1180039,I1180022,);
DFFARX1 I_69206 (I1376748,I3563,I1180039,I1180113,);
not I_69207 (I1180121,I1376763);
not I_69208 (I1180138,I1376751);
nand I_69209 (I1180155,I1180138,I1180121);
nor I_69210 (I1180010,I1180113,I1180155);
DFFARX1 I_69211 (I1180155,I3563,I1180039,I1180195,);
not I_69212 (I1180031,I1180195);
not I_69213 (I1180217,I1376760);
nand I_69214 (I1180234,I1180138,I1180217);
DFFARX1 I_69215 (I1180234,I3563,I1180039,I1180260,);
not I_69216 (I1180268,I1180260);
not I_69217 (I1180285,I1376769);
nand I_69218 (I1180302,I1180285,I1376748);
and I_69219 (I1180319,I1180121,I1180302);
nor I_69220 (I1180336,I1180234,I1180319);
DFFARX1 I_69221 (I1180336,I3563,I1180039,I1180007,);
DFFARX1 I_69222 (I1180319,I3563,I1180039,I1180028,);
nor I_69223 (I1180381,I1376769,I1376772);
nor I_69224 (I1180019,I1180234,I1180381);
or I_69225 (I1180412,I1376769,I1376772);
nor I_69226 (I1180429,I1376766,I1376754);
DFFARX1 I_69227 (I1180429,I3563,I1180039,I1180455,);
not I_69228 (I1180463,I1180455);
nor I_69229 (I1180025,I1180463,I1180268);
nand I_69230 (I1180494,I1180463,I1180113);
not I_69231 (I1180511,I1376766);
nand I_69232 (I1180528,I1180511,I1180217);
nand I_69233 (I1180545,I1180463,I1180528);
nand I_69234 (I1180016,I1180545,I1180494);
nand I_69235 (I1180013,I1180528,I1180412);
not I_69236 (I1180617,I3570);
DFFARX1 I_69237 (I459394,I3563,I1180617,I1180643,);
and I_69238 (I1180651,I1180643,I459409);
DFFARX1 I_69239 (I1180651,I3563,I1180617,I1180600,);
DFFARX1 I_69240 (I459412,I3563,I1180617,I1180691,);
not I_69241 (I1180699,I459406);
not I_69242 (I1180716,I459421);
nand I_69243 (I1180733,I1180716,I1180699);
nor I_69244 (I1180588,I1180691,I1180733);
DFFARX1 I_69245 (I1180733,I3563,I1180617,I1180773,);
not I_69246 (I1180609,I1180773);
not I_69247 (I1180795,I459397);
nand I_69248 (I1180812,I1180716,I1180795);
DFFARX1 I_69249 (I1180812,I3563,I1180617,I1180838,);
not I_69250 (I1180846,I1180838);
not I_69251 (I1180863,I459400);
nand I_69252 (I1180880,I1180863,I459394);
and I_69253 (I1180897,I1180699,I1180880);
nor I_69254 (I1180914,I1180812,I1180897);
DFFARX1 I_69255 (I1180914,I3563,I1180617,I1180585,);
DFFARX1 I_69256 (I1180897,I3563,I1180617,I1180606,);
nor I_69257 (I1180959,I459400,I459403);
nor I_69258 (I1180597,I1180812,I1180959);
or I_69259 (I1180990,I459400,I459403);
nor I_69260 (I1181007,I459418,I459415);
DFFARX1 I_69261 (I1181007,I3563,I1180617,I1181033,);
not I_69262 (I1181041,I1181033);
nor I_69263 (I1180603,I1181041,I1180846);
nand I_69264 (I1181072,I1181041,I1180691);
not I_69265 (I1181089,I459418);
nand I_69266 (I1181106,I1181089,I1180795);
nand I_69267 (I1181123,I1181041,I1181106);
nand I_69268 (I1180594,I1181123,I1181072);
nand I_69269 (I1180591,I1181106,I1180990);
not I_69270 (I1181195,I3570);
DFFARX1 I_69271 (I1318411,I3563,I1181195,I1181221,);
and I_69272 (I1181229,I1181221,I1318393);
DFFARX1 I_69273 (I1181229,I3563,I1181195,I1181178,);
DFFARX1 I_69274 (I1318402,I3563,I1181195,I1181269,);
not I_69275 (I1181277,I1318387);
not I_69276 (I1181294,I1318399);
nand I_69277 (I1181311,I1181294,I1181277);
nor I_69278 (I1181166,I1181269,I1181311);
DFFARX1 I_69279 (I1181311,I3563,I1181195,I1181351,);
not I_69280 (I1181187,I1181351);
not I_69281 (I1181373,I1318390);
nand I_69282 (I1181390,I1181294,I1181373);
DFFARX1 I_69283 (I1181390,I3563,I1181195,I1181416,);
not I_69284 (I1181424,I1181416);
not I_69285 (I1181441,I1318387);
nand I_69286 (I1181458,I1181441,I1318390);
and I_69287 (I1181475,I1181277,I1181458);
nor I_69288 (I1181492,I1181390,I1181475);
DFFARX1 I_69289 (I1181492,I3563,I1181195,I1181163,);
DFFARX1 I_69290 (I1181475,I3563,I1181195,I1181184,);
nor I_69291 (I1181537,I1318387,I1318408);
nor I_69292 (I1181175,I1181390,I1181537);
or I_69293 (I1181568,I1318387,I1318408);
nor I_69294 (I1181585,I1318396,I1318405);
DFFARX1 I_69295 (I1181585,I3563,I1181195,I1181611,);
not I_69296 (I1181619,I1181611);
nor I_69297 (I1181181,I1181619,I1181424);
nand I_69298 (I1181650,I1181619,I1181269);
not I_69299 (I1181667,I1318396);
nand I_69300 (I1181684,I1181667,I1181373);
nand I_69301 (I1181701,I1181619,I1181684);
nand I_69302 (I1181172,I1181701,I1181650);
nand I_69303 (I1181169,I1181684,I1181568);
not I_69304 (I1181773,I3570);
DFFARX1 I_69305 (I525762,I3563,I1181773,I1181799,);
and I_69306 (I1181807,I1181799,I525777);
DFFARX1 I_69307 (I1181807,I3563,I1181773,I1181756,);
DFFARX1 I_69308 (I525780,I3563,I1181773,I1181847,);
not I_69309 (I1181855,I525774);
not I_69310 (I1181872,I525789);
nand I_69311 (I1181889,I1181872,I1181855);
nor I_69312 (I1181744,I1181847,I1181889);
DFFARX1 I_69313 (I1181889,I3563,I1181773,I1181929,);
not I_69314 (I1181765,I1181929);
not I_69315 (I1181951,I525765);
nand I_69316 (I1181968,I1181872,I1181951);
DFFARX1 I_69317 (I1181968,I3563,I1181773,I1181994,);
not I_69318 (I1182002,I1181994);
not I_69319 (I1182019,I525768);
nand I_69320 (I1182036,I1182019,I525762);
and I_69321 (I1182053,I1181855,I1182036);
nor I_69322 (I1182070,I1181968,I1182053);
DFFARX1 I_69323 (I1182070,I3563,I1181773,I1181741,);
DFFARX1 I_69324 (I1182053,I3563,I1181773,I1181762,);
nor I_69325 (I1182115,I525768,I525771);
nor I_69326 (I1181753,I1181968,I1182115);
or I_69327 (I1182146,I525768,I525771);
nor I_69328 (I1182163,I525786,I525783);
DFFARX1 I_69329 (I1182163,I3563,I1181773,I1182189,);
not I_69330 (I1182197,I1182189);
nor I_69331 (I1181759,I1182197,I1182002);
nand I_69332 (I1182228,I1182197,I1181847);
not I_69333 (I1182245,I525786);
nand I_69334 (I1182262,I1182245,I1181951);
nand I_69335 (I1182279,I1182197,I1182262);
nand I_69336 (I1181750,I1182279,I1182228);
nand I_69337 (I1181747,I1182262,I1182146);
not I_69338 (I1182351,I3570);
DFFARX1 I_69339 (I1285054,I3563,I1182351,I1182377,);
and I_69340 (I1182385,I1182377,I1285048);
DFFARX1 I_69341 (I1182385,I3563,I1182351,I1182334,);
DFFARX1 I_69342 (I1285033,I3563,I1182351,I1182425,);
not I_69343 (I1182433,I1285039);
not I_69344 (I1182450,I1285051);
nand I_69345 (I1182467,I1182450,I1182433);
nor I_69346 (I1182322,I1182425,I1182467);
DFFARX1 I_69347 (I1182467,I3563,I1182351,I1182507,);
not I_69348 (I1182343,I1182507);
not I_69349 (I1182529,I1285033);
nand I_69350 (I1182546,I1182450,I1182529);
DFFARX1 I_69351 (I1182546,I3563,I1182351,I1182572,);
not I_69352 (I1182580,I1182572);
not I_69353 (I1182597,I1285057);
nand I_69354 (I1182614,I1182597,I1285045);
and I_69355 (I1182631,I1182433,I1182614);
nor I_69356 (I1182648,I1182546,I1182631);
DFFARX1 I_69357 (I1182648,I3563,I1182351,I1182319,);
DFFARX1 I_69358 (I1182631,I3563,I1182351,I1182340,);
nor I_69359 (I1182693,I1285057,I1285036);
nor I_69360 (I1182331,I1182546,I1182693);
or I_69361 (I1182724,I1285057,I1285036);
nor I_69362 (I1182741,I1285042,I1285036);
DFFARX1 I_69363 (I1182741,I3563,I1182351,I1182767,);
not I_69364 (I1182775,I1182767);
nor I_69365 (I1182337,I1182775,I1182580);
nand I_69366 (I1182806,I1182775,I1182425);
not I_69367 (I1182823,I1285042);
nand I_69368 (I1182840,I1182823,I1182529);
nand I_69369 (I1182857,I1182775,I1182840);
nand I_69370 (I1182328,I1182857,I1182806);
nand I_69371 (I1182325,I1182840,I1182724);
not I_69372 (I1182929,I3570);
DFFARX1 I_69373 (I223213,I3563,I1182929,I1182955,);
and I_69374 (I1182963,I1182955,I223216);
DFFARX1 I_69375 (I1182963,I3563,I1182929,I1182912,);
DFFARX1 I_69376 (I223216,I3563,I1182929,I1183003,);
not I_69377 (I1183011,I223231);
not I_69378 (I1183028,I223237);
nand I_69379 (I1183045,I1183028,I1183011);
nor I_69380 (I1182900,I1183003,I1183045);
DFFARX1 I_69381 (I1183045,I3563,I1182929,I1183085,);
not I_69382 (I1182921,I1183085);
not I_69383 (I1183107,I223225);
nand I_69384 (I1183124,I1183028,I1183107);
DFFARX1 I_69385 (I1183124,I3563,I1182929,I1183150,);
not I_69386 (I1183158,I1183150);
not I_69387 (I1183175,I223222);
nand I_69388 (I1183192,I1183175,I223219);
and I_69389 (I1183209,I1183011,I1183192);
nor I_69390 (I1183226,I1183124,I1183209);
DFFARX1 I_69391 (I1183226,I3563,I1182929,I1182897,);
DFFARX1 I_69392 (I1183209,I3563,I1182929,I1182918,);
nor I_69393 (I1183271,I223222,I223213);
nor I_69394 (I1182909,I1183124,I1183271);
or I_69395 (I1183302,I223222,I223213);
nor I_69396 (I1183319,I223228,I223234);
DFFARX1 I_69397 (I1183319,I3563,I1182929,I1183345,);
not I_69398 (I1183353,I1183345);
nor I_69399 (I1182915,I1183353,I1183158);
nand I_69400 (I1183384,I1183353,I1183003);
not I_69401 (I1183401,I223228);
nand I_69402 (I1183418,I1183401,I1183107);
nand I_69403 (I1183435,I1183353,I1183418);
nand I_69404 (I1182906,I1183435,I1183384);
nand I_69405 (I1182903,I1183418,I1183302);
not I_69406 (I1183507,I3570);
DFFARX1 I_69407 (I911716,I3563,I1183507,I1183533,);
and I_69408 (I1183541,I1183533,I911722);
DFFARX1 I_69409 (I1183541,I3563,I1183507,I1183490,);
DFFARX1 I_69410 (I911728,I3563,I1183507,I1183581,);
not I_69411 (I1183589,I911713);
not I_69412 (I1183606,I911713);
nand I_69413 (I1183623,I1183606,I1183589);
nor I_69414 (I1183478,I1183581,I1183623);
DFFARX1 I_69415 (I1183623,I3563,I1183507,I1183663,);
not I_69416 (I1183499,I1183663);
not I_69417 (I1183685,I911731);
nand I_69418 (I1183702,I1183606,I1183685);
DFFARX1 I_69419 (I1183702,I3563,I1183507,I1183728,);
not I_69420 (I1183736,I1183728);
not I_69421 (I1183753,I911725);
nand I_69422 (I1183770,I1183753,I911716);
and I_69423 (I1183787,I1183589,I1183770);
nor I_69424 (I1183804,I1183702,I1183787);
DFFARX1 I_69425 (I1183804,I3563,I1183507,I1183475,);
DFFARX1 I_69426 (I1183787,I3563,I1183507,I1183496,);
nor I_69427 (I1183849,I911725,I911734);
nor I_69428 (I1183487,I1183702,I1183849);
or I_69429 (I1183880,I911725,I911734);
nor I_69430 (I1183897,I911719,I911719);
DFFARX1 I_69431 (I1183897,I3563,I1183507,I1183923,);
not I_69432 (I1183931,I1183923);
nor I_69433 (I1183493,I1183931,I1183736);
nand I_69434 (I1183962,I1183931,I1183581);
not I_69435 (I1183979,I911719);
nand I_69436 (I1183996,I1183979,I1183685);
nand I_69437 (I1184013,I1183931,I1183996);
nand I_69438 (I1183484,I1184013,I1183962);
nand I_69439 (I1183481,I1183996,I1183880);
not I_69440 (I1184085,I3570);
DFFARX1 I_69441 (I94615,I3563,I1184085,I1184111,);
and I_69442 (I1184119,I1184111,I94591);
DFFARX1 I_69443 (I1184119,I3563,I1184085,I1184068,);
DFFARX1 I_69444 (I94609,I3563,I1184085,I1184159,);
not I_69445 (I1184167,I94597);
not I_69446 (I1184184,I94594);
nand I_69447 (I1184201,I1184184,I1184167);
nor I_69448 (I1184056,I1184159,I1184201);
DFFARX1 I_69449 (I1184201,I3563,I1184085,I1184241,);
not I_69450 (I1184077,I1184241);
not I_69451 (I1184263,I94603);
nand I_69452 (I1184280,I1184184,I1184263);
DFFARX1 I_69453 (I1184280,I3563,I1184085,I1184306,);
not I_69454 (I1184314,I1184306);
not I_69455 (I1184331,I94594);
nand I_69456 (I1184348,I1184331,I94612);
and I_69457 (I1184365,I1184167,I1184348);
nor I_69458 (I1184382,I1184280,I1184365);
DFFARX1 I_69459 (I1184382,I3563,I1184085,I1184053,);
DFFARX1 I_69460 (I1184365,I3563,I1184085,I1184074,);
nor I_69461 (I1184427,I94594,I94606);
nor I_69462 (I1184065,I1184280,I1184427);
or I_69463 (I1184458,I94594,I94606);
nor I_69464 (I1184475,I94600,I94591);
DFFARX1 I_69465 (I1184475,I3563,I1184085,I1184501,);
not I_69466 (I1184509,I1184501);
nor I_69467 (I1184071,I1184509,I1184314);
nand I_69468 (I1184540,I1184509,I1184159);
not I_69469 (I1184557,I94600);
nand I_69470 (I1184574,I1184557,I1184263);
nand I_69471 (I1184591,I1184509,I1184574);
nand I_69472 (I1184062,I1184591,I1184540);
nand I_69473 (I1184059,I1184574,I1184458);
not I_69474 (I1184663,I3570);
DFFARX1 I_69475 (I138883,I3563,I1184663,I1184689,);
and I_69476 (I1184697,I1184689,I138859);
DFFARX1 I_69477 (I1184697,I3563,I1184663,I1184646,);
DFFARX1 I_69478 (I138877,I3563,I1184663,I1184737,);
not I_69479 (I1184745,I138865);
not I_69480 (I1184762,I138862);
nand I_69481 (I1184779,I1184762,I1184745);
nor I_69482 (I1184634,I1184737,I1184779);
DFFARX1 I_69483 (I1184779,I3563,I1184663,I1184819,);
not I_69484 (I1184655,I1184819);
not I_69485 (I1184841,I138871);
nand I_69486 (I1184858,I1184762,I1184841);
DFFARX1 I_69487 (I1184858,I3563,I1184663,I1184884,);
not I_69488 (I1184892,I1184884);
not I_69489 (I1184909,I138862);
nand I_69490 (I1184926,I1184909,I138880);
and I_69491 (I1184943,I1184745,I1184926);
nor I_69492 (I1184960,I1184858,I1184943);
DFFARX1 I_69493 (I1184960,I3563,I1184663,I1184631,);
DFFARX1 I_69494 (I1184943,I3563,I1184663,I1184652,);
nor I_69495 (I1185005,I138862,I138874);
nor I_69496 (I1184643,I1184858,I1185005);
or I_69497 (I1185036,I138862,I138874);
nor I_69498 (I1185053,I138868,I138859);
DFFARX1 I_69499 (I1185053,I3563,I1184663,I1185079,);
not I_69500 (I1185087,I1185079);
nor I_69501 (I1184649,I1185087,I1184892);
nand I_69502 (I1185118,I1185087,I1184737);
not I_69503 (I1185135,I138868);
nand I_69504 (I1185152,I1185135,I1184841);
nand I_69505 (I1185169,I1185087,I1185152);
nand I_69506 (I1184640,I1185169,I1185118);
nand I_69507 (I1184637,I1185152,I1185036);
not I_69508 (I1185241,I3570);
DFFARX1 I_69509 (I1075273,I3563,I1185241,I1185267,);
and I_69510 (I1185275,I1185267,I1075270);
DFFARX1 I_69511 (I1185275,I3563,I1185241,I1185224,);
DFFARX1 I_69512 (I1075276,I3563,I1185241,I1185315,);
not I_69513 (I1185323,I1075279);
not I_69514 (I1185340,I1075273);
nand I_69515 (I1185357,I1185340,I1185323);
nor I_69516 (I1185212,I1185315,I1185357);
DFFARX1 I_69517 (I1185357,I3563,I1185241,I1185397,);
not I_69518 (I1185233,I1185397);
not I_69519 (I1185419,I1075288);
nand I_69520 (I1185436,I1185340,I1185419);
DFFARX1 I_69521 (I1185436,I3563,I1185241,I1185462,);
not I_69522 (I1185470,I1185462);
not I_69523 (I1185487,I1075285);
nand I_69524 (I1185504,I1185487,I1075291);
and I_69525 (I1185521,I1185323,I1185504);
nor I_69526 (I1185538,I1185436,I1185521);
DFFARX1 I_69527 (I1185538,I3563,I1185241,I1185209,);
DFFARX1 I_69528 (I1185521,I3563,I1185241,I1185230,);
nor I_69529 (I1185583,I1075285,I1075270);
nor I_69530 (I1185221,I1185436,I1185583);
or I_69531 (I1185614,I1075285,I1075270);
nor I_69532 (I1185631,I1075282,I1075276);
DFFARX1 I_69533 (I1185631,I3563,I1185241,I1185657,);
not I_69534 (I1185665,I1185657);
nor I_69535 (I1185227,I1185665,I1185470);
nand I_69536 (I1185696,I1185665,I1185315);
not I_69537 (I1185713,I1075282);
nand I_69538 (I1185730,I1185713,I1185419);
nand I_69539 (I1185747,I1185665,I1185730);
nand I_69540 (I1185218,I1185747,I1185696);
nand I_69541 (I1185215,I1185730,I1185614);
not I_69542 (I1185819,I3570);
DFFARX1 I_69543 (I1402360,I3563,I1185819,I1185845,);
and I_69544 (I1185853,I1185845,I1402342);
DFFARX1 I_69545 (I1185853,I3563,I1185819,I1185802,);
DFFARX1 I_69546 (I1402333,I3563,I1185819,I1185893,);
not I_69547 (I1185901,I1402348);
not I_69548 (I1185918,I1402336);
nand I_69549 (I1185935,I1185918,I1185901);
nor I_69550 (I1185790,I1185893,I1185935);
DFFARX1 I_69551 (I1185935,I3563,I1185819,I1185975,);
not I_69552 (I1185811,I1185975);
not I_69553 (I1185997,I1402345);
nand I_69554 (I1186014,I1185918,I1185997);
DFFARX1 I_69555 (I1186014,I3563,I1185819,I1186040,);
not I_69556 (I1186048,I1186040);
not I_69557 (I1186065,I1402354);
nand I_69558 (I1186082,I1186065,I1402333);
and I_69559 (I1186099,I1185901,I1186082);
nor I_69560 (I1186116,I1186014,I1186099);
DFFARX1 I_69561 (I1186116,I3563,I1185819,I1185787,);
DFFARX1 I_69562 (I1186099,I3563,I1185819,I1185808,);
nor I_69563 (I1186161,I1402354,I1402357);
nor I_69564 (I1185799,I1186014,I1186161);
or I_69565 (I1186192,I1402354,I1402357);
nor I_69566 (I1186209,I1402351,I1402339);
DFFARX1 I_69567 (I1186209,I3563,I1185819,I1186235,);
not I_69568 (I1186243,I1186235);
nor I_69569 (I1185805,I1186243,I1186048);
nand I_69570 (I1186274,I1186243,I1185893);
not I_69571 (I1186291,I1402351);
nand I_69572 (I1186308,I1186291,I1185997);
nand I_69573 (I1186325,I1186243,I1186308);
nand I_69574 (I1185796,I1186325,I1186274);
nand I_69575 (I1185793,I1186308,I1186192);
not I_69576 (I1186397,I3570);
DFFARX1 I_69577 (I382887,I3563,I1186397,I1186423,);
and I_69578 (I1186431,I1186423,I382872);
DFFARX1 I_69579 (I1186431,I3563,I1186397,I1186380,);
DFFARX1 I_69580 (I382878,I3563,I1186397,I1186471,);
not I_69581 (I1186479,I382860);
not I_69582 (I1186496,I382881);
nand I_69583 (I1186513,I1186496,I1186479);
nor I_69584 (I1186368,I1186471,I1186513);
DFFARX1 I_69585 (I1186513,I3563,I1186397,I1186553,);
not I_69586 (I1186389,I1186553);
not I_69587 (I1186575,I382884);
nand I_69588 (I1186592,I1186496,I1186575);
DFFARX1 I_69589 (I1186592,I3563,I1186397,I1186618,);
not I_69590 (I1186626,I1186618);
not I_69591 (I1186643,I382875);
nand I_69592 (I1186660,I1186643,I382863);
and I_69593 (I1186677,I1186479,I1186660);
nor I_69594 (I1186694,I1186592,I1186677);
DFFARX1 I_69595 (I1186694,I3563,I1186397,I1186365,);
DFFARX1 I_69596 (I1186677,I3563,I1186397,I1186386,);
nor I_69597 (I1186739,I382875,I382869);
nor I_69598 (I1186377,I1186592,I1186739);
or I_69599 (I1186770,I382875,I382869);
nor I_69600 (I1186787,I382866,I382860);
DFFARX1 I_69601 (I1186787,I3563,I1186397,I1186813,);
not I_69602 (I1186821,I1186813);
nor I_69603 (I1186383,I1186821,I1186626);
nand I_69604 (I1186852,I1186821,I1186471);
not I_69605 (I1186869,I382866);
nand I_69606 (I1186886,I1186869,I1186575);
nand I_69607 (I1186903,I1186821,I1186886);
nand I_69608 (I1186374,I1186903,I1186852);
nand I_69609 (I1186371,I1186886,I1186770);
not I_69610 (I1186975,I3570);
DFFARX1 I_69611 (I318066,I3563,I1186975,I1187001,);
and I_69612 (I1187009,I1187001,I318051);
DFFARX1 I_69613 (I1187009,I3563,I1186975,I1186958,);
DFFARX1 I_69614 (I318057,I3563,I1186975,I1187049,);
not I_69615 (I1187057,I318039);
not I_69616 (I1187074,I318060);
nand I_69617 (I1187091,I1187074,I1187057);
nor I_69618 (I1186946,I1187049,I1187091);
DFFARX1 I_69619 (I1187091,I3563,I1186975,I1187131,);
not I_69620 (I1186967,I1187131);
not I_69621 (I1187153,I318063);
nand I_69622 (I1187170,I1187074,I1187153);
DFFARX1 I_69623 (I1187170,I3563,I1186975,I1187196,);
not I_69624 (I1187204,I1187196);
not I_69625 (I1187221,I318054);
nand I_69626 (I1187238,I1187221,I318042);
and I_69627 (I1187255,I1187057,I1187238);
nor I_69628 (I1187272,I1187170,I1187255);
DFFARX1 I_69629 (I1187272,I3563,I1186975,I1186943,);
DFFARX1 I_69630 (I1187255,I3563,I1186975,I1186964,);
nor I_69631 (I1187317,I318054,I318048);
nor I_69632 (I1186955,I1187170,I1187317);
or I_69633 (I1187348,I318054,I318048);
nor I_69634 (I1187365,I318045,I318039);
DFFARX1 I_69635 (I1187365,I3563,I1186975,I1187391,);
not I_69636 (I1187399,I1187391);
nor I_69637 (I1186961,I1187399,I1187204);
nand I_69638 (I1187430,I1187399,I1187049);
not I_69639 (I1187447,I318045);
nand I_69640 (I1187464,I1187447,I1187153);
nand I_69641 (I1187481,I1187399,I1187464);
nand I_69642 (I1186952,I1187481,I1187430);
nand I_69643 (I1186949,I1187464,I1187348);
not I_69644 (I1187553,I3570);
DFFARX1 I_69645 (I1018241,I3563,I1187553,I1187579,);
and I_69646 (I1187587,I1187579,I1018235);
DFFARX1 I_69647 (I1187587,I3563,I1187553,I1187536,);
DFFARX1 I_69648 (I1018253,I3563,I1187553,I1187627,);
not I_69649 (I1187635,I1018244);
not I_69650 (I1187652,I1018256);
nand I_69651 (I1187669,I1187652,I1187635);
nor I_69652 (I1187524,I1187627,I1187669);
DFFARX1 I_69653 (I1187669,I3563,I1187553,I1187709,);
not I_69654 (I1187545,I1187709);
not I_69655 (I1187731,I1018262);
nand I_69656 (I1187748,I1187652,I1187731);
DFFARX1 I_69657 (I1187748,I3563,I1187553,I1187774,);
not I_69658 (I1187782,I1187774);
not I_69659 (I1187799,I1018238);
nand I_69660 (I1187816,I1187799,I1018259);
and I_69661 (I1187833,I1187635,I1187816);
nor I_69662 (I1187850,I1187748,I1187833);
DFFARX1 I_69663 (I1187850,I3563,I1187553,I1187521,);
DFFARX1 I_69664 (I1187833,I3563,I1187553,I1187542,);
nor I_69665 (I1187895,I1018238,I1018250);
nor I_69666 (I1187533,I1187748,I1187895);
or I_69667 (I1187926,I1018238,I1018250);
nor I_69668 (I1187943,I1018235,I1018247);
DFFARX1 I_69669 (I1187943,I3563,I1187553,I1187969,);
not I_69670 (I1187977,I1187969);
nor I_69671 (I1187539,I1187977,I1187782);
nand I_69672 (I1188008,I1187977,I1187627);
not I_69673 (I1188025,I1018235);
nand I_69674 (I1188042,I1188025,I1187731);
nand I_69675 (I1188059,I1187977,I1188042);
nand I_69676 (I1187530,I1188059,I1188008);
nand I_69677 (I1187527,I1188042,I1187926);
not I_69678 (I1188131,I3570);
DFFARX1 I_69679 (I415034,I3563,I1188131,I1188157,);
and I_69680 (I1188165,I1188157,I415019);
DFFARX1 I_69681 (I1188165,I3563,I1188131,I1188114,);
DFFARX1 I_69682 (I415025,I3563,I1188131,I1188205,);
not I_69683 (I1188213,I415007);
not I_69684 (I1188230,I415028);
nand I_69685 (I1188247,I1188230,I1188213);
nor I_69686 (I1188102,I1188205,I1188247);
DFFARX1 I_69687 (I1188247,I3563,I1188131,I1188287,);
not I_69688 (I1188123,I1188287);
not I_69689 (I1188309,I415031);
nand I_69690 (I1188326,I1188230,I1188309);
DFFARX1 I_69691 (I1188326,I3563,I1188131,I1188352,);
not I_69692 (I1188360,I1188352);
not I_69693 (I1188377,I415022);
nand I_69694 (I1188394,I1188377,I415010);
and I_69695 (I1188411,I1188213,I1188394);
nor I_69696 (I1188428,I1188326,I1188411);
DFFARX1 I_69697 (I1188428,I3563,I1188131,I1188099,);
DFFARX1 I_69698 (I1188411,I3563,I1188131,I1188120,);
nor I_69699 (I1188473,I415022,I415016);
nor I_69700 (I1188111,I1188326,I1188473);
or I_69701 (I1188504,I415022,I415016);
nor I_69702 (I1188521,I415013,I415007);
DFFARX1 I_69703 (I1188521,I3563,I1188131,I1188547,);
not I_69704 (I1188555,I1188547);
nor I_69705 (I1188117,I1188555,I1188360);
nand I_69706 (I1188586,I1188555,I1188205);
not I_69707 (I1188603,I415013);
nand I_69708 (I1188620,I1188603,I1188309);
nand I_69709 (I1188637,I1188555,I1188620);
nand I_69710 (I1188108,I1188637,I1188586);
nand I_69711 (I1188105,I1188620,I1188504);
not I_69712 (I1188709,I3570);
DFFARX1 I_69713 (I753220,I3563,I1188709,I1188735,);
and I_69714 (I1188743,I1188735,I753208);
DFFARX1 I_69715 (I1188743,I3563,I1188709,I1188692,);
DFFARX1 I_69716 (I753211,I3563,I1188709,I1188783,);
not I_69717 (I1188791,I753205);
not I_69718 (I1188808,I753229);
nand I_69719 (I1188825,I1188808,I1188791);
nor I_69720 (I1188680,I1188783,I1188825);
DFFARX1 I_69721 (I1188825,I3563,I1188709,I1188865,);
not I_69722 (I1188701,I1188865);
not I_69723 (I1188887,I753217);
nand I_69724 (I1188904,I1188808,I1188887);
DFFARX1 I_69725 (I1188904,I3563,I1188709,I1188930,);
not I_69726 (I1188938,I1188930);
not I_69727 (I1188955,I753226);
nand I_69728 (I1188972,I1188955,I753223);
and I_69729 (I1188989,I1188791,I1188972);
nor I_69730 (I1189006,I1188904,I1188989);
DFFARX1 I_69731 (I1189006,I3563,I1188709,I1188677,);
DFFARX1 I_69732 (I1188989,I3563,I1188709,I1188698,);
nor I_69733 (I1189051,I753226,I753214);
nor I_69734 (I1188689,I1188904,I1189051);
or I_69735 (I1189082,I753226,I753214);
nor I_69736 (I1189099,I753205,I753208);
DFFARX1 I_69737 (I1189099,I3563,I1188709,I1189125,);
not I_69738 (I1189133,I1189125);
nor I_69739 (I1188695,I1189133,I1188938);
nand I_69740 (I1189164,I1189133,I1188783);
not I_69741 (I1189181,I753205);
nand I_69742 (I1189198,I1189181,I1188887);
nand I_69743 (I1189215,I1189133,I1189198);
nand I_69744 (I1188686,I1189215,I1189164);
nand I_69745 (I1188683,I1189198,I1189082);
not I_69746 (I1189287,I3570);
DFFARX1 I_69747 (I769982,I3563,I1189287,I1189313,);
and I_69748 (I1189321,I1189313,I769970);
DFFARX1 I_69749 (I1189321,I3563,I1189287,I1189270,);
DFFARX1 I_69750 (I769973,I3563,I1189287,I1189361,);
not I_69751 (I1189369,I769967);
not I_69752 (I1189386,I769991);
nand I_69753 (I1189403,I1189386,I1189369);
nor I_69754 (I1189258,I1189361,I1189403);
DFFARX1 I_69755 (I1189403,I3563,I1189287,I1189443,);
not I_69756 (I1189279,I1189443);
not I_69757 (I1189465,I769979);
nand I_69758 (I1189482,I1189386,I1189465);
DFFARX1 I_69759 (I1189482,I3563,I1189287,I1189508,);
not I_69760 (I1189516,I1189508);
not I_69761 (I1189533,I769988);
nand I_69762 (I1189550,I1189533,I769985);
and I_69763 (I1189567,I1189369,I1189550);
nor I_69764 (I1189584,I1189482,I1189567);
DFFARX1 I_69765 (I1189584,I3563,I1189287,I1189255,);
DFFARX1 I_69766 (I1189567,I3563,I1189287,I1189276,);
nor I_69767 (I1189629,I769988,I769976);
nor I_69768 (I1189267,I1189482,I1189629);
or I_69769 (I1189660,I769988,I769976);
nor I_69770 (I1189677,I769967,I769970);
DFFARX1 I_69771 (I1189677,I3563,I1189287,I1189703,);
not I_69772 (I1189711,I1189703);
nor I_69773 (I1189273,I1189711,I1189516);
nand I_69774 (I1189742,I1189711,I1189361);
not I_69775 (I1189759,I769967);
nand I_69776 (I1189776,I1189759,I1189465);
nand I_69777 (I1189793,I1189711,I1189776);
nand I_69778 (I1189264,I1189793,I1189742);
nand I_69779 (I1189261,I1189776,I1189660);
not I_69780 (I1189865,I3570);
DFFARX1 I_69781 (I1367850,I3563,I1189865,I1189891,);
and I_69782 (I1189899,I1189891,I1367832);
DFFARX1 I_69783 (I1189899,I3563,I1189865,I1189848,);
DFFARX1 I_69784 (I1367823,I3563,I1189865,I1189939,);
not I_69785 (I1189947,I1367838);
not I_69786 (I1189964,I1367826);
nand I_69787 (I1189981,I1189964,I1189947);
nor I_69788 (I1189836,I1189939,I1189981);
DFFARX1 I_69789 (I1189981,I3563,I1189865,I1190021,);
not I_69790 (I1189857,I1190021);
not I_69791 (I1190043,I1367835);
nand I_69792 (I1190060,I1189964,I1190043);
DFFARX1 I_69793 (I1190060,I3563,I1189865,I1190086,);
not I_69794 (I1190094,I1190086);
not I_69795 (I1190111,I1367844);
nand I_69796 (I1190128,I1190111,I1367823);
and I_69797 (I1190145,I1189947,I1190128);
nor I_69798 (I1190162,I1190060,I1190145);
DFFARX1 I_69799 (I1190162,I3563,I1189865,I1189833,);
DFFARX1 I_69800 (I1190145,I3563,I1189865,I1189854,);
nor I_69801 (I1190207,I1367844,I1367847);
nor I_69802 (I1189845,I1190060,I1190207);
or I_69803 (I1190238,I1367844,I1367847);
nor I_69804 (I1190255,I1367841,I1367829);
DFFARX1 I_69805 (I1190255,I3563,I1189865,I1190281,);
not I_69806 (I1190289,I1190281);
nor I_69807 (I1189851,I1190289,I1190094);
nand I_69808 (I1190320,I1190289,I1189939);
not I_69809 (I1190337,I1367841);
nand I_69810 (I1190354,I1190337,I1190043);
nand I_69811 (I1190371,I1190289,I1190354);
nand I_69812 (I1189842,I1190371,I1190320);
nand I_69813 (I1189839,I1190354,I1190238);
not I_69814 (I1190443,I3570);
DFFARX1 I_69815 (I694842,I3563,I1190443,I1190469,);
and I_69816 (I1190477,I1190469,I694830);
DFFARX1 I_69817 (I1190477,I3563,I1190443,I1190426,);
DFFARX1 I_69818 (I694833,I3563,I1190443,I1190517,);
not I_69819 (I1190525,I694827);
not I_69820 (I1190542,I694851);
nand I_69821 (I1190559,I1190542,I1190525);
nor I_69822 (I1190414,I1190517,I1190559);
DFFARX1 I_69823 (I1190559,I3563,I1190443,I1190599,);
not I_69824 (I1190435,I1190599);
not I_69825 (I1190621,I694839);
nand I_69826 (I1190638,I1190542,I1190621);
DFFARX1 I_69827 (I1190638,I3563,I1190443,I1190664,);
not I_69828 (I1190672,I1190664);
not I_69829 (I1190689,I694848);
nand I_69830 (I1190706,I1190689,I694845);
and I_69831 (I1190723,I1190525,I1190706);
nor I_69832 (I1190740,I1190638,I1190723);
DFFARX1 I_69833 (I1190740,I3563,I1190443,I1190411,);
DFFARX1 I_69834 (I1190723,I3563,I1190443,I1190432,);
nor I_69835 (I1190785,I694848,I694836);
nor I_69836 (I1190423,I1190638,I1190785);
or I_69837 (I1190816,I694848,I694836);
nor I_69838 (I1190833,I694827,I694830);
DFFARX1 I_69839 (I1190833,I3563,I1190443,I1190859,);
not I_69840 (I1190867,I1190859);
nor I_69841 (I1190429,I1190867,I1190672);
nand I_69842 (I1190898,I1190867,I1190517);
not I_69843 (I1190915,I694827);
nand I_69844 (I1190932,I1190915,I1190621);
nand I_69845 (I1190949,I1190867,I1190932);
nand I_69846 (I1190420,I1190949,I1190898);
nand I_69847 (I1190417,I1190932,I1190816);
not I_69848 (I1191021,I3570);
DFFARX1 I_69849 (I405021,I3563,I1191021,I1191047,);
and I_69850 (I1191055,I1191047,I405006);
DFFARX1 I_69851 (I1191055,I3563,I1191021,I1191004,);
DFFARX1 I_69852 (I405012,I3563,I1191021,I1191095,);
not I_69853 (I1191103,I404994);
not I_69854 (I1191120,I405015);
nand I_69855 (I1191137,I1191120,I1191103);
nor I_69856 (I1190992,I1191095,I1191137);
DFFARX1 I_69857 (I1191137,I3563,I1191021,I1191177,);
not I_69858 (I1191013,I1191177);
not I_69859 (I1191199,I405018);
nand I_69860 (I1191216,I1191120,I1191199);
DFFARX1 I_69861 (I1191216,I3563,I1191021,I1191242,);
not I_69862 (I1191250,I1191242);
not I_69863 (I1191267,I405009);
nand I_69864 (I1191284,I1191267,I404997);
and I_69865 (I1191301,I1191103,I1191284);
nor I_69866 (I1191318,I1191216,I1191301);
DFFARX1 I_69867 (I1191318,I3563,I1191021,I1190989,);
DFFARX1 I_69868 (I1191301,I3563,I1191021,I1191010,);
nor I_69869 (I1191363,I405009,I405003);
nor I_69870 (I1191001,I1191216,I1191363);
or I_69871 (I1191394,I405009,I405003);
nor I_69872 (I1191411,I405000,I404994);
DFFARX1 I_69873 (I1191411,I3563,I1191021,I1191437,);
not I_69874 (I1191445,I1191437);
nor I_69875 (I1191007,I1191445,I1191250);
nand I_69876 (I1191476,I1191445,I1191095);
not I_69877 (I1191493,I405000);
nand I_69878 (I1191510,I1191493,I1191199);
nand I_69879 (I1191527,I1191445,I1191510);
nand I_69880 (I1190998,I1191527,I1191476);
nand I_69881 (I1190995,I1191510,I1191394);
not I_69882 (I1191599,I3570);
DFFARX1 I_69883 (I188703,I3563,I1191599,I1191625,);
and I_69884 (I1191633,I1191625,I188706);
DFFARX1 I_69885 (I1191633,I3563,I1191599,I1191582,);
DFFARX1 I_69886 (I188706,I3563,I1191599,I1191673,);
not I_69887 (I1191681,I188721);
not I_69888 (I1191698,I188727);
nand I_69889 (I1191715,I1191698,I1191681);
nor I_69890 (I1191570,I1191673,I1191715);
DFFARX1 I_69891 (I1191715,I3563,I1191599,I1191755,);
not I_69892 (I1191591,I1191755);
not I_69893 (I1191777,I188715);
nand I_69894 (I1191794,I1191698,I1191777);
DFFARX1 I_69895 (I1191794,I3563,I1191599,I1191820,);
not I_69896 (I1191828,I1191820);
not I_69897 (I1191845,I188712);
nand I_69898 (I1191862,I1191845,I188709);
and I_69899 (I1191879,I1191681,I1191862);
nor I_69900 (I1191896,I1191794,I1191879);
DFFARX1 I_69901 (I1191896,I3563,I1191599,I1191567,);
DFFARX1 I_69902 (I1191879,I3563,I1191599,I1191588,);
nor I_69903 (I1191941,I188712,I188703);
nor I_69904 (I1191579,I1191794,I1191941);
or I_69905 (I1191972,I188712,I188703);
nor I_69906 (I1191989,I188718,I188724);
DFFARX1 I_69907 (I1191989,I3563,I1191599,I1192015,);
not I_69908 (I1192023,I1192015);
nor I_69909 (I1191585,I1192023,I1191828);
nand I_69910 (I1192054,I1192023,I1191673);
not I_69911 (I1192071,I188718);
nand I_69912 (I1192088,I1192071,I1191777);
nand I_69913 (I1192105,I1192023,I1192088);
nand I_69914 (I1191576,I1192105,I1192054);
nand I_69915 (I1191573,I1192088,I1191972);
not I_69916 (I1192177,I3570);
DFFARX1 I_69917 (I324917,I3563,I1192177,I1192203,);
and I_69918 (I1192211,I1192203,I324902);
DFFARX1 I_69919 (I1192211,I3563,I1192177,I1192160,);
DFFARX1 I_69920 (I324908,I3563,I1192177,I1192251,);
not I_69921 (I1192259,I324890);
not I_69922 (I1192276,I324911);
nand I_69923 (I1192293,I1192276,I1192259);
nor I_69924 (I1192148,I1192251,I1192293);
DFFARX1 I_69925 (I1192293,I3563,I1192177,I1192333,);
not I_69926 (I1192169,I1192333);
not I_69927 (I1192355,I324914);
nand I_69928 (I1192372,I1192276,I1192355);
DFFARX1 I_69929 (I1192372,I3563,I1192177,I1192398,);
not I_69930 (I1192406,I1192398);
not I_69931 (I1192423,I324905);
nand I_69932 (I1192440,I1192423,I324893);
and I_69933 (I1192457,I1192259,I1192440);
nor I_69934 (I1192474,I1192372,I1192457);
DFFARX1 I_69935 (I1192474,I3563,I1192177,I1192145,);
DFFARX1 I_69936 (I1192457,I3563,I1192177,I1192166,);
nor I_69937 (I1192519,I324905,I324899);
nor I_69938 (I1192157,I1192372,I1192519);
or I_69939 (I1192550,I324905,I324899);
nor I_69940 (I1192567,I324896,I324890);
DFFARX1 I_69941 (I1192567,I3563,I1192177,I1192593,);
not I_69942 (I1192601,I1192593);
nor I_69943 (I1192163,I1192601,I1192406);
nand I_69944 (I1192632,I1192601,I1192251);
not I_69945 (I1192649,I324896);
nand I_69946 (I1192666,I1192649,I1192355);
nand I_69947 (I1192683,I1192601,I1192666);
nand I_69948 (I1192154,I1192683,I1192632);
nand I_69949 (I1192151,I1192666,I1192550);
not I_69950 (I1192755,I3570);
DFFARX1 I_69951 (I1073029,I3563,I1192755,I1192781,);
and I_69952 (I1192789,I1192781,I1073026);
DFFARX1 I_69953 (I1192789,I3563,I1192755,I1192738,);
DFFARX1 I_69954 (I1073032,I3563,I1192755,I1192829,);
not I_69955 (I1192837,I1073035);
not I_69956 (I1192854,I1073029);
nand I_69957 (I1192871,I1192854,I1192837);
nor I_69958 (I1192726,I1192829,I1192871);
DFFARX1 I_69959 (I1192871,I3563,I1192755,I1192911,);
not I_69960 (I1192747,I1192911);
not I_69961 (I1192933,I1073044);
nand I_69962 (I1192950,I1192854,I1192933);
DFFARX1 I_69963 (I1192950,I3563,I1192755,I1192976,);
not I_69964 (I1192984,I1192976);
not I_69965 (I1193001,I1073041);
nand I_69966 (I1193018,I1193001,I1073047);
and I_69967 (I1193035,I1192837,I1193018);
nor I_69968 (I1193052,I1192950,I1193035);
DFFARX1 I_69969 (I1193052,I3563,I1192755,I1192723,);
DFFARX1 I_69970 (I1193035,I3563,I1192755,I1192744,);
nor I_69971 (I1193097,I1073041,I1073026);
nor I_69972 (I1192735,I1192950,I1193097);
or I_69973 (I1193128,I1073041,I1073026);
nor I_69974 (I1193145,I1073038,I1073032);
DFFARX1 I_69975 (I1193145,I3563,I1192755,I1193171,);
not I_69976 (I1193179,I1193171);
nor I_69977 (I1192741,I1193179,I1192984);
nand I_69978 (I1193210,I1193179,I1192829);
not I_69979 (I1193227,I1073038);
nand I_69980 (I1193244,I1193227,I1192933);
nand I_69981 (I1193261,I1193179,I1193244);
nand I_69982 (I1192732,I1193261,I1193210);
nand I_69983 (I1192729,I1193244,I1193128);
not I_69984 (I1193333,I3570);
DFFARX1 I_69985 (I870083,I3563,I1193333,I1193359,);
and I_69986 (I1193367,I1193359,I870089);
DFFARX1 I_69987 (I1193367,I3563,I1193333,I1193316,);
DFFARX1 I_69988 (I870095,I3563,I1193333,I1193407,);
not I_69989 (I1193415,I870080);
not I_69990 (I1193432,I870080);
nand I_69991 (I1193449,I1193432,I1193415);
nor I_69992 (I1193304,I1193407,I1193449);
DFFARX1 I_69993 (I1193449,I3563,I1193333,I1193489,);
not I_69994 (I1193325,I1193489);
not I_69995 (I1193511,I870098);
nand I_69996 (I1193528,I1193432,I1193511);
DFFARX1 I_69997 (I1193528,I3563,I1193333,I1193554,);
not I_69998 (I1193562,I1193554);
not I_69999 (I1193579,I870092);
nand I_70000 (I1193596,I1193579,I870083);
and I_70001 (I1193613,I1193415,I1193596);
nor I_70002 (I1193630,I1193528,I1193613);
DFFARX1 I_70003 (I1193630,I3563,I1193333,I1193301,);
DFFARX1 I_70004 (I1193613,I3563,I1193333,I1193322,);
nor I_70005 (I1193675,I870092,I870101);
nor I_70006 (I1193313,I1193528,I1193675);
or I_70007 (I1193706,I870092,I870101);
nor I_70008 (I1193723,I870086,I870086);
DFFARX1 I_70009 (I1193723,I3563,I1193333,I1193749,);
not I_70010 (I1193757,I1193749);
nor I_70011 (I1193319,I1193757,I1193562);
nand I_70012 (I1193788,I1193757,I1193407);
not I_70013 (I1193805,I870086);
nand I_70014 (I1193822,I1193805,I1193511);
nand I_70015 (I1193839,I1193757,I1193822);
nand I_70016 (I1193310,I1193839,I1193788);
nand I_70017 (I1193307,I1193822,I1193706);
not I_70018 (I1193911,I3570);
DFFARX1 I_70019 (I1383320,I3563,I1193911,I1193937,);
and I_70020 (I1193945,I1193937,I1383302);
DFFARX1 I_70021 (I1193945,I3563,I1193911,I1193894,);
DFFARX1 I_70022 (I1383293,I3563,I1193911,I1193985,);
not I_70023 (I1193993,I1383308);
not I_70024 (I1194010,I1383296);
nand I_70025 (I1194027,I1194010,I1193993);
nor I_70026 (I1193882,I1193985,I1194027);
DFFARX1 I_70027 (I1194027,I3563,I1193911,I1194067,);
not I_70028 (I1193903,I1194067);
not I_70029 (I1194089,I1383305);
nand I_70030 (I1194106,I1194010,I1194089);
DFFARX1 I_70031 (I1194106,I3563,I1193911,I1194132,);
not I_70032 (I1194140,I1194132);
not I_70033 (I1194157,I1383314);
nand I_70034 (I1194174,I1194157,I1383293);
and I_70035 (I1194191,I1193993,I1194174);
nor I_70036 (I1194208,I1194106,I1194191);
DFFARX1 I_70037 (I1194208,I3563,I1193911,I1193879,);
DFFARX1 I_70038 (I1194191,I3563,I1193911,I1193900,);
nor I_70039 (I1194253,I1383314,I1383317);
nor I_70040 (I1193891,I1194106,I1194253);
or I_70041 (I1194284,I1383314,I1383317);
nor I_70042 (I1194301,I1383311,I1383299);
DFFARX1 I_70043 (I1194301,I3563,I1193911,I1194327,);
not I_70044 (I1194335,I1194327);
nor I_70045 (I1193897,I1194335,I1194140);
nand I_70046 (I1194366,I1194335,I1193985);
not I_70047 (I1194383,I1383311);
nand I_70048 (I1194400,I1194383,I1194089);
nand I_70049 (I1194417,I1194335,I1194400);
nand I_70050 (I1193888,I1194417,I1194366);
nand I_70051 (I1193885,I1194400,I1194284);
not I_70052 (I1194489,I3570);
DFFARX1 I_70053 (I929093,I3563,I1194489,I1194515,);
and I_70054 (I1194523,I1194515,I929087);
DFFARX1 I_70055 (I1194523,I3563,I1194489,I1194472,);
DFFARX1 I_70056 (I929105,I3563,I1194489,I1194563,);
not I_70057 (I1194571,I929096);
not I_70058 (I1194588,I929108);
nand I_70059 (I1194605,I1194588,I1194571);
nor I_70060 (I1194460,I1194563,I1194605);
DFFARX1 I_70061 (I1194605,I3563,I1194489,I1194645,);
not I_70062 (I1194481,I1194645);
not I_70063 (I1194667,I929114);
nand I_70064 (I1194684,I1194588,I1194667);
DFFARX1 I_70065 (I1194684,I3563,I1194489,I1194710,);
not I_70066 (I1194718,I1194710);
not I_70067 (I1194735,I929090);
nand I_70068 (I1194752,I1194735,I929111);
and I_70069 (I1194769,I1194571,I1194752);
nor I_70070 (I1194786,I1194684,I1194769);
DFFARX1 I_70071 (I1194786,I3563,I1194489,I1194457,);
DFFARX1 I_70072 (I1194769,I3563,I1194489,I1194478,);
nor I_70073 (I1194831,I929090,I929102);
nor I_70074 (I1194469,I1194684,I1194831);
or I_70075 (I1194862,I929090,I929102);
nor I_70076 (I1194879,I929087,I929099);
DFFARX1 I_70077 (I1194879,I3563,I1194489,I1194905,);
not I_70078 (I1194913,I1194905);
nor I_70079 (I1194475,I1194913,I1194718);
nand I_70080 (I1194944,I1194913,I1194563);
not I_70081 (I1194961,I929087);
nand I_70082 (I1194978,I1194961,I1194667);
nand I_70083 (I1194995,I1194913,I1194978);
nand I_70084 (I1194466,I1194995,I1194944);
nand I_70085 (I1194463,I1194978,I1194862);
not I_70086 (I1195067,I3570);
DFFARX1 I_70087 (I576884,I3563,I1195067,I1195093,);
and I_70088 (I1195101,I1195093,I576899);
DFFARX1 I_70089 (I1195101,I3563,I1195067,I1195050,);
DFFARX1 I_70090 (I576890,I3563,I1195067,I1195141,);
not I_70091 (I1195149,I576884);
not I_70092 (I1195166,I576902);
nand I_70093 (I1195183,I1195166,I1195149);
nor I_70094 (I1195038,I1195141,I1195183);
DFFARX1 I_70095 (I1195183,I3563,I1195067,I1195223,);
not I_70096 (I1195059,I1195223);
not I_70097 (I1195245,I576893);
nand I_70098 (I1195262,I1195166,I1195245);
DFFARX1 I_70099 (I1195262,I3563,I1195067,I1195288,);
not I_70100 (I1195296,I1195288);
not I_70101 (I1195313,I576905);
nand I_70102 (I1195330,I1195313,I576881);
and I_70103 (I1195347,I1195149,I1195330);
nor I_70104 (I1195364,I1195262,I1195347);
DFFARX1 I_70105 (I1195364,I3563,I1195067,I1195035,);
DFFARX1 I_70106 (I1195347,I3563,I1195067,I1195056,);
nor I_70107 (I1195409,I576905,I576881);
nor I_70108 (I1195047,I1195262,I1195409);
or I_70109 (I1195440,I576905,I576881);
nor I_70110 (I1195457,I576887,I576896);
DFFARX1 I_70111 (I1195457,I3563,I1195067,I1195483,);
not I_70112 (I1195491,I1195483);
nor I_70113 (I1195053,I1195491,I1195296);
nand I_70114 (I1195522,I1195491,I1195141);
not I_70115 (I1195539,I576887);
nand I_70116 (I1195556,I1195539,I1195245);
nand I_70117 (I1195573,I1195491,I1195556);
nand I_70118 (I1195044,I1195573,I1195522);
nand I_70119 (I1195041,I1195556,I1195440);
not I_70120 (I1195645,I3570);
DFFARX1 I_70121 (I924571,I3563,I1195645,I1195671,);
and I_70122 (I1195679,I1195671,I924565);
DFFARX1 I_70123 (I1195679,I3563,I1195645,I1195628,);
DFFARX1 I_70124 (I924583,I3563,I1195645,I1195719,);
not I_70125 (I1195727,I924574);
not I_70126 (I1195744,I924586);
nand I_70127 (I1195761,I1195744,I1195727);
nor I_70128 (I1195616,I1195719,I1195761);
DFFARX1 I_70129 (I1195761,I3563,I1195645,I1195801,);
not I_70130 (I1195637,I1195801);
not I_70131 (I1195823,I924592);
nand I_70132 (I1195840,I1195744,I1195823);
DFFARX1 I_70133 (I1195840,I3563,I1195645,I1195866,);
not I_70134 (I1195874,I1195866);
not I_70135 (I1195891,I924568);
nand I_70136 (I1195908,I1195891,I924589);
and I_70137 (I1195925,I1195727,I1195908);
nor I_70138 (I1195942,I1195840,I1195925);
DFFARX1 I_70139 (I1195942,I3563,I1195645,I1195613,);
DFFARX1 I_70140 (I1195925,I3563,I1195645,I1195634,);
nor I_70141 (I1195987,I924568,I924580);
nor I_70142 (I1195625,I1195840,I1195987);
or I_70143 (I1196018,I924568,I924580);
nor I_70144 (I1196035,I924565,I924577);
DFFARX1 I_70145 (I1196035,I3563,I1195645,I1196061,);
not I_70146 (I1196069,I1196061);
nor I_70147 (I1195631,I1196069,I1195874);
nand I_70148 (I1196100,I1196069,I1195719);
not I_70149 (I1196117,I924565);
nand I_70150 (I1196134,I1196117,I1195823);
nand I_70151 (I1196151,I1196069,I1196134);
nand I_70152 (I1195622,I1196151,I1196100);
nand I_70153 (I1195619,I1196134,I1196018);
not I_70154 (I1196223,I3570);
DFFARX1 I_70155 (I87237,I3563,I1196223,I1196249,);
and I_70156 (I1196257,I1196249,I87213);
DFFARX1 I_70157 (I1196257,I3563,I1196223,I1196206,);
DFFARX1 I_70158 (I87231,I3563,I1196223,I1196297,);
not I_70159 (I1196305,I87219);
not I_70160 (I1196322,I87216);
nand I_70161 (I1196339,I1196322,I1196305);
nor I_70162 (I1196194,I1196297,I1196339);
DFFARX1 I_70163 (I1196339,I3563,I1196223,I1196379,);
not I_70164 (I1196215,I1196379);
not I_70165 (I1196401,I87225);
nand I_70166 (I1196418,I1196322,I1196401);
DFFARX1 I_70167 (I1196418,I3563,I1196223,I1196444,);
not I_70168 (I1196452,I1196444);
not I_70169 (I1196469,I87216);
nand I_70170 (I1196486,I1196469,I87234);
and I_70171 (I1196503,I1196305,I1196486);
nor I_70172 (I1196520,I1196418,I1196503);
DFFARX1 I_70173 (I1196520,I3563,I1196223,I1196191,);
DFFARX1 I_70174 (I1196503,I3563,I1196223,I1196212,);
nor I_70175 (I1196565,I87216,I87228);
nor I_70176 (I1196203,I1196418,I1196565);
or I_70177 (I1196596,I87216,I87228);
nor I_70178 (I1196613,I87222,I87213);
DFFARX1 I_70179 (I1196613,I3563,I1196223,I1196639,);
not I_70180 (I1196647,I1196639);
nor I_70181 (I1196209,I1196647,I1196452);
nand I_70182 (I1196678,I1196647,I1196297);
not I_70183 (I1196695,I87222);
nand I_70184 (I1196712,I1196695,I1196401);
nand I_70185 (I1196729,I1196647,I1196712);
nand I_70186 (I1196200,I1196729,I1196678);
nand I_70187 (I1196197,I1196712,I1196596);
not I_70188 (I1196801,I3570);
DFFARX1 I_70189 (I276168,I3563,I1196801,I1196827,);
and I_70190 (I1196835,I1196827,I276171);
DFFARX1 I_70191 (I1196835,I3563,I1196801,I1196784,);
DFFARX1 I_70192 (I276171,I3563,I1196801,I1196875,);
not I_70193 (I1196883,I276186);
not I_70194 (I1196900,I276192);
nand I_70195 (I1196917,I1196900,I1196883);
nor I_70196 (I1196772,I1196875,I1196917);
DFFARX1 I_70197 (I1196917,I3563,I1196801,I1196957,);
not I_70198 (I1196793,I1196957);
not I_70199 (I1196979,I276180);
nand I_70200 (I1196996,I1196900,I1196979);
DFFARX1 I_70201 (I1196996,I3563,I1196801,I1197022,);
not I_70202 (I1197030,I1197022);
not I_70203 (I1197047,I276177);
nand I_70204 (I1197064,I1197047,I276174);
and I_70205 (I1197081,I1196883,I1197064);
nor I_70206 (I1197098,I1196996,I1197081);
DFFARX1 I_70207 (I1197098,I3563,I1196801,I1196769,);
DFFARX1 I_70208 (I1197081,I3563,I1196801,I1196790,);
nor I_70209 (I1197143,I276177,I276168);
nor I_70210 (I1196781,I1196996,I1197143);
or I_70211 (I1197174,I276177,I276168);
nor I_70212 (I1197191,I276183,I276189);
DFFARX1 I_70213 (I1197191,I3563,I1196801,I1197217,);
not I_70214 (I1197225,I1197217);
nor I_70215 (I1196787,I1197225,I1197030);
nand I_70216 (I1197256,I1197225,I1196875);
not I_70217 (I1197273,I276183);
nand I_70218 (I1197290,I1197273,I1196979);
nand I_70219 (I1197307,I1197225,I1197290);
nand I_70220 (I1196778,I1197307,I1197256);
nand I_70221 (I1196775,I1197290,I1197174);
not I_70222 (I1197379,I3570);
DFFARX1 I_70223 (I839517,I3563,I1197379,I1197405,);
and I_70224 (I1197413,I1197405,I839523);
DFFARX1 I_70225 (I1197413,I3563,I1197379,I1197362,);
DFFARX1 I_70226 (I839529,I3563,I1197379,I1197453,);
not I_70227 (I1197461,I839514);
not I_70228 (I1197478,I839514);
nand I_70229 (I1197495,I1197478,I1197461);
nor I_70230 (I1197350,I1197453,I1197495);
DFFARX1 I_70231 (I1197495,I3563,I1197379,I1197535,);
not I_70232 (I1197371,I1197535);
not I_70233 (I1197557,I839532);
nand I_70234 (I1197574,I1197478,I1197557);
DFFARX1 I_70235 (I1197574,I3563,I1197379,I1197600,);
not I_70236 (I1197608,I1197600);
not I_70237 (I1197625,I839526);
nand I_70238 (I1197642,I1197625,I839517);
and I_70239 (I1197659,I1197461,I1197642);
nor I_70240 (I1197676,I1197574,I1197659);
DFFARX1 I_70241 (I1197676,I3563,I1197379,I1197347,);
DFFARX1 I_70242 (I1197659,I3563,I1197379,I1197368,);
nor I_70243 (I1197721,I839526,I839535);
nor I_70244 (I1197359,I1197574,I1197721);
or I_70245 (I1197752,I839526,I839535);
nor I_70246 (I1197769,I839520,I839520);
DFFARX1 I_70247 (I1197769,I3563,I1197379,I1197795,);
not I_70248 (I1197803,I1197795);
nor I_70249 (I1197365,I1197803,I1197608);
nand I_70250 (I1197834,I1197803,I1197453);
not I_70251 (I1197851,I839520);
nand I_70252 (I1197868,I1197851,I1197557);
nand I_70253 (I1197885,I1197803,I1197868);
nand I_70254 (I1197356,I1197885,I1197834);
nand I_70255 (I1197353,I1197868,I1197752);
not I_70256 (I1197957,I3570);
DFFARX1 I_70257 (I739926,I3563,I1197957,I1197983,);
and I_70258 (I1197991,I1197983,I739914);
DFFARX1 I_70259 (I1197991,I3563,I1197957,I1197940,);
DFFARX1 I_70260 (I739917,I3563,I1197957,I1198031,);
not I_70261 (I1198039,I739911);
not I_70262 (I1198056,I739935);
nand I_70263 (I1198073,I1198056,I1198039);
nor I_70264 (I1197928,I1198031,I1198073);
DFFARX1 I_70265 (I1198073,I3563,I1197957,I1198113,);
not I_70266 (I1197949,I1198113);
not I_70267 (I1198135,I739923);
nand I_70268 (I1198152,I1198056,I1198135);
DFFARX1 I_70269 (I1198152,I3563,I1197957,I1198178,);
not I_70270 (I1198186,I1198178);
not I_70271 (I1198203,I739932);
nand I_70272 (I1198220,I1198203,I739929);
and I_70273 (I1198237,I1198039,I1198220);
nor I_70274 (I1198254,I1198152,I1198237);
DFFARX1 I_70275 (I1198254,I3563,I1197957,I1197925,);
DFFARX1 I_70276 (I1198237,I3563,I1197957,I1197946,);
nor I_70277 (I1198299,I739932,I739920);
nor I_70278 (I1197937,I1198152,I1198299);
or I_70279 (I1198330,I739932,I739920);
nor I_70280 (I1198347,I739911,I739914);
DFFARX1 I_70281 (I1198347,I3563,I1197957,I1198373,);
not I_70282 (I1198381,I1198373);
nor I_70283 (I1197943,I1198381,I1198186);
nand I_70284 (I1198412,I1198381,I1198031);
not I_70285 (I1198429,I739911);
nand I_70286 (I1198446,I1198429,I1198135);
nand I_70287 (I1198463,I1198381,I1198446);
nand I_70288 (I1197934,I1198463,I1198412);
nand I_70289 (I1197931,I1198446,I1198330);
not I_70290 (I1198535,I3570);
DFFARX1 I_70291 (I119384,I3563,I1198535,I1198561,);
and I_70292 (I1198569,I1198561,I119360);
DFFARX1 I_70293 (I1198569,I3563,I1198535,I1198518,);
DFFARX1 I_70294 (I119378,I3563,I1198535,I1198609,);
not I_70295 (I1198617,I119366);
not I_70296 (I1198634,I119363);
nand I_70297 (I1198651,I1198634,I1198617);
nor I_70298 (I1198506,I1198609,I1198651);
DFFARX1 I_70299 (I1198651,I3563,I1198535,I1198691,);
not I_70300 (I1198527,I1198691);
not I_70301 (I1198713,I119372);
nand I_70302 (I1198730,I1198634,I1198713);
DFFARX1 I_70303 (I1198730,I3563,I1198535,I1198756,);
not I_70304 (I1198764,I1198756);
not I_70305 (I1198781,I119363);
nand I_70306 (I1198798,I1198781,I119381);
and I_70307 (I1198815,I1198617,I1198798);
nor I_70308 (I1198832,I1198730,I1198815);
DFFARX1 I_70309 (I1198832,I3563,I1198535,I1198503,);
DFFARX1 I_70310 (I1198815,I3563,I1198535,I1198524,);
nor I_70311 (I1198877,I119363,I119375);
nor I_70312 (I1198515,I1198730,I1198877);
or I_70313 (I1198908,I119363,I119375);
nor I_70314 (I1198925,I119369,I119360);
DFFARX1 I_70315 (I1198925,I3563,I1198535,I1198951,);
not I_70316 (I1198959,I1198951);
nor I_70317 (I1198521,I1198959,I1198764);
nand I_70318 (I1198990,I1198959,I1198609);
not I_70319 (I1199007,I119369);
nand I_70320 (I1199024,I1199007,I1198713);
nand I_70321 (I1199041,I1198959,I1199024);
nand I_70322 (I1198512,I1199041,I1198990);
nand I_70323 (I1198509,I1199024,I1198908);
not I_70324 (I1199113,I3570);
DFFARX1 I_70325 (I821072,I3563,I1199113,I1199139,);
and I_70326 (I1199147,I1199139,I821078);
DFFARX1 I_70327 (I1199147,I3563,I1199113,I1199096,);
DFFARX1 I_70328 (I821084,I3563,I1199113,I1199187,);
not I_70329 (I1199195,I821069);
not I_70330 (I1199212,I821069);
nand I_70331 (I1199229,I1199212,I1199195);
nor I_70332 (I1199084,I1199187,I1199229);
DFFARX1 I_70333 (I1199229,I3563,I1199113,I1199269,);
not I_70334 (I1199105,I1199269);
not I_70335 (I1199291,I821087);
nand I_70336 (I1199308,I1199212,I1199291);
DFFARX1 I_70337 (I1199308,I3563,I1199113,I1199334,);
not I_70338 (I1199342,I1199334);
not I_70339 (I1199359,I821081);
nand I_70340 (I1199376,I1199359,I821072);
and I_70341 (I1199393,I1199195,I1199376);
nor I_70342 (I1199410,I1199308,I1199393);
DFFARX1 I_70343 (I1199410,I3563,I1199113,I1199081,);
DFFARX1 I_70344 (I1199393,I3563,I1199113,I1199102,);
nor I_70345 (I1199455,I821081,I821090);
nor I_70346 (I1199093,I1199308,I1199455);
or I_70347 (I1199486,I821081,I821090);
nor I_70348 (I1199503,I821075,I821075);
DFFARX1 I_70349 (I1199503,I3563,I1199113,I1199529,);
not I_70350 (I1199537,I1199529);
nor I_70351 (I1199099,I1199537,I1199342);
nand I_70352 (I1199568,I1199537,I1199187);
not I_70353 (I1199585,I821075);
nand I_70354 (I1199602,I1199585,I1199291);
nand I_70355 (I1199619,I1199537,I1199602);
nand I_70356 (I1199090,I1199619,I1199568);
nand I_70357 (I1199087,I1199602,I1199486);
not I_70358 (I1199691,I3570);
DFFARX1 I_70359 (I60887,I3563,I1199691,I1199717,);
and I_70360 (I1199725,I1199717,I60863);
DFFARX1 I_70361 (I1199725,I3563,I1199691,I1199674,);
DFFARX1 I_70362 (I60881,I3563,I1199691,I1199765,);
not I_70363 (I1199773,I60869);
not I_70364 (I1199790,I60866);
nand I_70365 (I1199807,I1199790,I1199773);
nor I_70366 (I1199662,I1199765,I1199807);
DFFARX1 I_70367 (I1199807,I3563,I1199691,I1199847,);
not I_70368 (I1199683,I1199847);
not I_70369 (I1199869,I60875);
nand I_70370 (I1199886,I1199790,I1199869);
DFFARX1 I_70371 (I1199886,I3563,I1199691,I1199912,);
not I_70372 (I1199920,I1199912);
not I_70373 (I1199937,I60866);
nand I_70374 (I1199954,I1199937,I60884);
and I_70375 (I1199971,I1199773,I1199954);
nor I_70376 (I1199988,I1199886,I1199971);
DFFARX1 I_70377 (I1199988,I3563,I1199691,I1199659,);
DFFARX1 I_70378 (I1199971,I3563,I1199691,I1199680,);
nor I_70379 (I1200033,I60866,I60878);
nor I_70380 (I1199671,I1199886,I1200033);
or I_70381 (I1200064,I60866,I60878);
nor I_70382 (I1200081,I60872,I60863);
DFFARX1 I_70383 (I1200081,I3563,I1199691,I1200107,);
not I_70384 (I1200115,I1200107);
nor I_70385 (I1199677,I1200115,I1199920);
nand I_70386 (I1200146,I1200115,I1199765);
not I_70387 (I1200163,I60872);
nand I_70388 (I1200180,I1200163,I1199869);
nand I_70389 (I1200197,I1200115,I1200180);
nand I_70390 (I1199668,I1200197,I1200146);
nand I_70391 (I1199665,I1200180,I1200064);
not I_70392 (I1200269,I3570);
DFFARX1 I_70393 (I815802,I3563,I1200269,I1200295,);
and I_70394 (I1200303,I1200295,I815808);
DFFARX1 I_70395 (I1200303,I3563,I1200269,I1200252,);
DFFARX1 I_70396 (I815814,I3563,I1200269,I1200343,);
not I_70397 (I1200351,I815799);
not I_70398 (I1200368,I815799);
nand I_70399 (I1200385,I1200368,I1200351);
nor I_70400 (I1200240,I1200343,I1200385);
DFFARX1 I_70401 (I1200385,I3563,I1200269,I1200425,);
not I_70402 (I1200261,I1200425);
not I_70403 (I1200447,I815817);
nand I_70404 (I1200464,I1200368,I1200447);
DFFARX1 I_70405 (I1200464,I3563,I1200269,I1200490,);
not I_70406 (I1200498,I1200490);
not I_70407 (I1200515,I815811);
nand I_70408 (I1200532,I1200515,I815802);
and I_70409 (I1200549,I1200351,I1200532);
nor I_70410 (I1200566,I1200464,I1200549);
DFFARX1 I_70411 (I1200566,I3563,I1200269,I1200237,);
DFFARX1 I_70412 (I1200549,I3563,I1200269,I1200258,);
nor I_70413 (I1200611,I815811,I815820);
nor I_70414 (I1200249,I1200464,I1200611);
or I_70415 (I1200642,I815811,I815820);
nor I_70416 (I1200659,I815805,I815805);
DFFARX1 I_70417 (I1200659,I3563,I1200269,I1200685,);
not I_70418 (I1200693,I1200685);
nor I_70419 (I1200255,I1200693,I1200498);
nand I_70420 (I1200724,I1200693,I1200343);
not I_70421 (I1200741,I815805);
nand I_70422 (I1200758,I1200741,I1200447);
nand I_70423 (I1200775,I1200693,I1200758);
nand I_70424 (I1200246,I1200775,I1200724);
nand I_70425 (I1200243,I1200758,I1200642);
not I_70426 (I1200847,I3570);
DFFARX1 I_70427 (I1336910,I3563,I1200847,I1200873,);
and I_70428 (I1200881,I1200873,I1336892);
DFFARX1 I_70429 (I1200881,I3563,I1200847,I1200830,);
DFFARX1 I_70430 (I1336883,I3563,I1200847,I1200921,);
not I_70431 (I1200929,I1336898);
not I_70432 (I1200946,I1336886);
nand I_70433 (I1200963,I1200946,I1200929);
nor I_70434 (I1200818,I1200921,I1200963);
DFFARX1 I_70435 (I1200963,I3563,I1200847,I1201003,);
not I_70436 (I1200839,I1201003);
not I_70437 (I1201025,I1336895);
nand I_70438 (I1201042,I1200946,I1201025);
DFFARX1 I_70439 (I1201042,I3563,I1200847,I1201068,);
not I_70440 (I1201076,I1201068);
not I_70441 (I1201093,I1336904);
nand I_70442 (I1201110,I1201093,I1336883);
and I_70443 (I1201127,I1200929,I1201110);
nor I_70444 (I1201144,I1201042,I1201127);
DFFARX1 I_70445 (I1201144,I3563,I1200847,I1200815,);
DFFARX1 I_70446 (I1201127,I3563,I1200847,I1200836,);
nor I_70447 (I1201189,I1336904,I1336907);
nor I_70448 (I1200827,I1201042,I1201189);
or I_70449 (I1201220,I1336904,I1336907);
nor I_70450 (I1201237,I1336901,I1336889);
DFFARX1 I_70451 (I1201237,I3563,I1200847,I1201263,);
not I_70452 (I1201271,I1201263);
nor I_70453 (I1200833,I1201271,I1201076);
nand I_70454 (I1201302,I1201271,I1200921);
not I_70455 (I1201319,I1336901);
nand I_70456 (I1201336,I1201319,I1201025);
nand I_70457 (I1201353,I1201271,I1201336);
nand I_70458 (I1200824,I1201353,I1201302);
nand I_70459 (I1200821,I1201336,I1201220);
not I_70460 (I1201425,I3570);
DFFARX1 I_70461 (I1033099,I3563,I1201425,I1201451,);
and I_70462 (I1201459,I1201451,I1033093);
DFFARX1 I_70463 (I1201459,I3563,I1201425,I1201408,);
DFFARX1 I_70464 (I1033111,I3563,I1201425,I1201499,);
not I_70465 (I1201507,I1033102);
not I_70466 (I1201524,I1033114);
nand I_70467 (I1201541,I1201524,I1201507);
nor I_70468 (I1201396,I1201499,I1201541);
DFFARX1 I_70469 (I1201541,I3563,I1201425,I1201581,);
not I_70470 (I1201417,I1201581);
not I_70471 (I1201603,I1033120);
nand I_70472 (I1201620,I1201524,I1201603);
DFFARX1 I_70473 (I1201620,I3563,I1201425,I1201646,);
not I_70474 (I1201654,I1201646);
not I_70475 (I1201671,I1033096);
nand I_70476 (I1201688,I1201671,I1033117);
and I_70477 (I1201705,I1201507,I1201688);
nor I_70478 (I1201722,I1201620,I1201705);
DFFARX1 I_70479 (I1201722,I3563,I1201425,I1201393,);
DFFARX1 I_70480 (I1201705,I3563,I1201425,I1201414,);
nor I_70481 (I1201767,I1033096,I1033108);
nor I_70482 (I1201405,I1201620,I1201767);
or I_70483 (I1201798,I1033096,I1033108);
nor I_70484 (I1201815,I1033093,I1033105);
DFFARX1 I_70485 (I1201815,I3563,I1201425,I1201841,);
not I_70486 (I1201849,I1201841);
nor I_70487 (I1201411,I1201849,I1201654);
nand I_70488 (I1201880,I1201849,I1201499);
not I_70489 (I1201897,I1033093);
nand I_70490 (I1201914,I1201897,I1201603);
nand I_70491 (I1201931,I1201849,I1201914);
nand I_70492 (I1201402,I1201931,I1201880);
nand I_70493 (I1201399,I1201914,I1201798);
not I_70494 (I1202003,I3570);
DFFARX1 I_70495 (I845841,I3563,I1202003,I1202029,);
and I_70496 (I1202037,I1202029,I845847);
DFFARX1 I_70497 (I1202037,I3563,I1202003,I1201986,);
DFFARX1 I_70498 (I845853,I3563,I1202003,I1202077,);
not I_70499 (I1202085,I845838);
not I_70500 (I1202102,I845838);
nand I_70501 (I1202119,I1202102,I1202085);
nor I_70502 (I1201974,I1202077,I1202119);
DFFARX1 I_70503 (I1202119,I3563,I1202003,I1202159,);
not I_70504 (I1201995,I1202159);
not I_70505 (I1202181,I845856);
nand I_70506 (I1202198,I1202102,I1202181);
DFFARX1 I_70507 (I1202198,I3563,I1202003,I1202224,);
not I_70508 (I1202232,I1202224);
not I_70509 (I1202249,I845850);
nand I_70510 (I1202266,I1202249,I845841);
and I_70511 (I1202283,I1202085,I1202266);
nor I_70512 (I1202300,I1202198,I1202283);
DFFARX1 I_70513 (I1202300,I3563,I1202003,I1201971,);
DFFARX1 I_70514 (I1202283,I3563,I1202003,I1201992,);
nor I_70515 (I1202345,I845850,I845859);
nor I_70516 (I1201983,I1202198,I1202345);
or I_70517 (I1202376,I845850,I845859);
nor I_70518 (I1202393,I845844,I845844);
DFFARX1 I_70519 (I1202393,I3563,I1202003,I1202419,);
not I_70520 (I1202427,I1202419);
nor I_70521 (I1201989,I1202427,I1202232);
nand I_70522 (I1202458,I1202427,I1202077);
not I_70523 (I1202475,I845844);
nand I_70524 (I1202492,I1202475,I1202181);
nand I_70525 (I1202509,I1202427,I1202492);
nand I_70526 (I1201980,I1202509,I1202458);
nand I_70527 (I1201977,I1202492,I1202376);
not I_70528 (I1202581,I3570);
DFFARX1 I_70529 (I850057,I3563,I1202581,I1202607,);
and I_70530 (I1202615,I1202607,I850063);
DFFARX1 I_70531 (I1202615,I3563,I1202581,I1202564,);
DFFARX1 I_70532 (I850069,I3563,I1202581,I1202655,);
not I_70533 (I1202663,I850054);
not I_70534 (I1202680,I850054);
nand I_70535 (I1202697,I1202680,I1202663);
nor I_70536 (I1202552,I1202655,I1202697);
DFFARX1 I_70537 (I1202697,I3563,I1202581,I1202737,);
not I_70538 (I1202573,I1202737);
not I_70539 (I1202759,I850072);
nand I_70540 (I1202776,I1202680,I1202759);
DFFARX1 I_70541 (I1202776,I3563,I1202581,I1202802,);
not I_70542 (I1202810,I1202802);
not I_70543 (I1202827,I850066);
nand I_70544 (I1202844,I1202827,I850057);
and I_70545 (I1202861,I1202663,I1202844);
nor I_70546 (I1202878,I1202776,I1202861);
DFFARX1 I_70547 (I1202878,I3563,I1202581,I1202549,);
DFFARX1 I_70548 (I1202861,I3563,I1202581,I1202570,);
nor I_70549 (I1202923,I850066,I850075);
nor I_70550 (I1202561,I1202776,I1202923);
or I_70551 (I1202954,I850066,I850075);
nor I_70552 (I1202971,I850060,I850060);
DFFARX1 I_70553 (I1202971,I3563,I1202581,I1202997,);
not I_70554 (I1203005,I1202997);
nor I_70555 (I1202567,I1203005,I1202810);
nand I_70556 (I1203036,I1203005,I1202655);
not I_70557 (I1203053,I850060);
nand I_70558 (I1203070,I1203053,I1202759);
nand I_70559 (I1203087,I1203005,I1203070);
nand I_70560 (I1202558,I1203087,I1203036);
nand I_70561 (I1202555,I1203070,I1202954);
not I_70562 (I1203159,I3570);
DFFARX1 I_70563 (I796570,I3563,I1203159,I1203185,);
and I_70564 (I1203193,I1203185,I796558);
DFFARX1 I_70565 (I1203193,I3563,I1203159,I1203142,);
DFFARX1 I_70566 (I796561,I3563,I1203159,I1203233,);
not I_70567 (I1203241,I796555);
not I_70568 (I1203258,I796579);
nand I_70569 (I1203275,I1203258,I1203241);
nor I_70570 (I1203130,I1203233,I1203275);
DFFARX1 I_70571 (I1203275,I3563,I1203159,I1203315,);
not I_70572 (I1203151,I1203315);
not I_70573 (I1203337,I796567);
nand I_70574 (I1203354,I1203258,I1203337);
DFFARX1 I_70575 (I1203354,I3563,I1203159,I1203380,);
not I_70576 (I1203388,I1203380);
not I_70577 (I1203405,I796576);
nand I_70578 (I1203422,I1203405,I796573);
and I_70579 (I1203439,I1203241,I1203422);
nor I_70580 (I1203456,I1203354,I1203439);
DFFARX1 I_70581 (I1203456,I3563,I1203159,I1203127,);
DFFARX1 I_70582 (I1203439,I3563,I1203159,I1203148,);
nor I_70583 (I1203501,I796576,I796564);
nor I_70584 (I1203139,I1203354,I1203501);
or I_70585 (I1203532,I796576,I796564);
nor I_70586 (I1203549,I796555,I796558);
DFFARX1 I_70587 (I1203549,I3563,I1203159,I1203575,);
not I_70588 (I1203583,I1203575);
nor I_70589 (I1203145,I1203583,I1203388);
nand I_70590 (I1203614,I1203583,I1203233);
not I_70591 (I1203631,I796555);
nand I_70592 (I1203648,I1203631,I1203337);
nand I_70593 (I1203665,I1203583,I1203648);
nand I_70594 (I1203136,I1203665,I1203614);
nand I_70595 (I1203133,I1203648,I1203532);
not I_70596 (I1203737,I3570);
DFFARX1 I_70597 (I743972,I3563,I1203737,I1203763,);
and I_70598 (I1203771,I1203763,I743960);
DFFARX1 I_70599 (I1203771,I3563,I1203737,I1203720,);
DFFARX1 I_70600 (I743963,I3563,I1203737,I1203811,);
not I_70601 (I1203819,I743957);
not I_70602 (I1203836,I743981);
nand I_70603 (I1203853,I1203836,I1203819);
nor I_70604 (I1203708,I1203811,I1203853);
DFFARX1 I_70605 (I1203853,I3563,I1203737,I1203893,);
not I_70606 (I1203729,I1203893);
not I_70607 (I1203915,I743969);
nand I_70608 (I1203932,I1203836,I1203915);
DFFARX1 I_70609 (I1203932,I3563,I1203737,I1203958,);
not I_70610 (I1203966,I1203958);
not I_70611 (I1203983,I743978);
nand I_70612 (I1204000,I1203983,I743975);
and I_70613 (I1204017,I1203819,I1204000);
nor I_70614 (I1204034,I1203932,I1204017);
DFFARX1 I_70615 (I1204034,I3563,I1203737,I1203705,);
DFFARX1 I_70616 (I1204017,I3563,I1203737,I1203726,);
nor I_70617 (I1204079,I743978,I743966);
nor I_70618 (I1203717,I1203932,I1204079);
or I_70619 (I1204110,I743978,I743966);
nor I_70620 (I1204127,I743957,I743960);
DFFARX1 I_70621 (I1204127,I3563,I1203737,I1204153,);
not I_70622 (I1204161,I1204153);
nor I_70623 (I1203723,I1204161,I1203966);
nand I_70624 (I1204192,I1204161,I1203811);
not I_70625 (I1204209,I743957);
nand I_70626 (I1204226,I1204209,I1203915);
nand I_70627 (I1204243,I1204161,I1204226);
nand I_70628 (I1203714,I1204243,I1204192);
nand I_70629 (I1203711,I1204226,I1204110);
not I_70630 (I1204315,I3570);
DFFARX1 I_70631 (I669410,I3563,I1204315,I1204341,);
and I_70632 (I1204349,I1204341,I669398);
DFFARX1 I_70633 (I1204349,I3563,I1204315,I1204298,);
DFFARX1 I_70634 (I669401,I3563,I1204315,I1204389,);
not I_70635 (I1204397,I669395);
not I_70636 (I1204414,I669419);
nand I_70637 (I1204431,I1204414,I1204397);
nor I_70638 (I1204286,I1204389,I1204431);
DFFARX1 I_70639 (I1204431,I3563,I1204315,I1204471,);
not I_70640 (I1204307,I1204471);
not I_70641 (I1204493,I669407);
nand I_70642 (I1204510,I1204414,I1204493);
DFFARX1 I_70643 (I1204510,I3563,I1204315,I1204536,);
not I_70644 (I1204544,I1204536);
not I_70645 (I1204561,I669416);
nand I_70646 (I1204578,I1204561,I669413);
and I_70647 (I1204595,I1204397,I1204578);
nor I_70648 (I1204612,I1204510,I1204595);
DFFARX1 I_70649 (I1204612,I3563,I1204315,I1204283,);
DFFARX1 I_70650 (I1204595,I3563,I1204315,I1204304,);
nor I_70651 (I1204657,I669416,I669404);
nor I_70652 (I1204295,I1204510,I1204657);
or I_70653 (I1204688,I669416,I669404);
nor I_70654 (I1204705,I669395,I669398);
DFFARX1 I_70655 (I1204705,I3563,I1204315,I1204731,);
not I_70656 (I1204739,I1204731);
nor I_70657 (I1204301,I1204739,I1204544);
nand I_70658 (I1204770,I1204739,I1204389);
not I_70659 (I1204787,I669395);
nand I_70660 (I1204804,I1204787,I1204493);
nand I_70661 (I1204821,I1204739,I1204804);
nand I_70662 (I1204292,I1204821,I1204770);
nand I_70663 (I1204289,I1204804,I1204688);
not I_70664 (I1204893,I3570);
DFFARX1 I_70665 (I216073,I3563,I1204893,I1204919,);
and I_70666 (I1204927,I1204919,I216076);
DFFARX1 I_70667 (I1204927,I3563,I1204893,I1204876,);
DFFARX1 I_70668 (I216076,I3563,I1204893,I1204967,);
not I_70669 (I1204975,I216091);
not I_70670 (I1204992,I216097);
nand I_70671 (I1205009,I1204992,I1204975);
nor I_70672 (I1204864,I1204967,I1205009);
DFFARX1 I_70673 (I1205009,I3563,I1204893,I1205049,);
not I_70674 (I1204885,I1205049);
not I_70675 (I1205071,I216085);
nand I_70676 (I1205088,I1204992,I1205071);
DFFARX1 I_70677 (I1205088,I3563,I1204893,I1205114,);
not I_70678 (I1205122,I1205114);
not I_70679 (I1205139,I216082);
nand I_70680 (I1205156,I1205139,I216079);
and I_70681 (I1205173,I1204975,I1205156);
nor I_70682 (I1205190,I1205088,I1205173);
DFFARX1 I_70683 (I1205190,I3563,I1204893,I1204861,);
DFFARX1 I_70684 (I1205173,I3563,I1204893,I1204882,);
nor I_70685 (I1205235,I216082,I216073);
nor I_70686 (I1204873,I1205088,I1205235);
or I_70687 (I1205266,I216082,I216073);
nor I_70688 (I1205283,I216088,I216094);
DFFARX1 I_70689 (I1205283,I3563,I1204893,I1205309,);
not I_70690 (I1205317,I1205309);
nor I_70691 (I1204879,I1205317,I1205122);
nand I_70692 (I1205348,I1205317,I1204967);
not I_70693 (I1205365,I216088);
nand I_70694 (I1205382,I1205365,I1205071);
nand I_70695 (I1205399,I1205317,I1205382);
nand I_70696 (I1204870,I1205399,I1205348);
nand I_70697 (I1204867,I1205382,I1205266);
not I_70698 (I1205471,I3570);
DFFARX1 I_70699 (I1361900,I3563,I1205471,I1205497,);
and I_70700 (I1205505,I1205497,I1361882);
DFFARX1 I_70701 (I1205505,I3563,I1205471,I1205454,);
DFFARX1 I_70702 (I1361873,I3563,I1205471,I1205545,);
not I_70703 (I1205553,I1361888);
not I_70704 (I1205570,I1361876);
nand I_70705 (I1205587,I1205570,I1205553);
nor I_70706 (I1205442,I1205545,I1205587);
DFFARX1 I_70707 (I1205587,I3563,I1205471,I1205627,);
not I_70708 (I1205463,I1205627);
not I_70709 (I1205649,I1361885);
nand I_70710 (I1205666,I1205570,I1205649);
DFFARX1 I_70711 (I1205666,I3563,I1205471,I1205692,);
not I_70712 (I1205700,I1205692);
not I_70713 (I1205717,I1361894);
nand I_70714 (I1205734,I1205717,I1361873);
and I_70715 (I1205751,I1205553,I1205734);
nor I_70716 (I1205768,I1205666,I1205751);
DFFARX1 I_70717 (I1205768,I3563,I1205471,I1205439,);
DFFARX1 I_70718 (I1205751,I3563,I1205471,I1205460,);
nor I_70719 (I1205813,I1361894,I1361897);
nor I_70720 (I1205451,I1205666,I1205813);
or I_70721 (I1205844,I1361894,I1361897);
nor I_70722 (I1205861,I1361891,I1361879);
DFFARX1 I_70723 (I1205861,I3563,I1205471,I1205887,);
not I_70724 (I1205895,I1205887);
nor I_70725 (I1205457,I1205895,I1205700);
nand I_70726 (I1205926,I1205895,I1205545);
not I_70727 (I1205943,I1361891);
nand I_70728 (I1205960,I1205943,I1205649);
nand I_70729 (I1205977,I1205895,I1205960);
nand I_70730 (I1205448,I1205977,I1205926);
nand I_70731 (I1205445,I1205960,I1205844);
not I_70732 (I1206049,I3570);
DFFARX1 I_70733 (I413453,I3563,I1206049,I1206075,);
and I_70734 (I1206083,I1206075,I413438);
DFFARX1 I_70735 (I1206083,I3563,I1206049,I1206032,);
DFFARX1 I_70736 (I413444,I3563,I1206049,I1206123,);
not I_70737 (I1206131,I413426);
not I_70738 (I1206148,I413447);
nand I_70739 (I1206165,I1206148,I1206131);
nor I_70740 (I1206020,I1206123,I1206165);
DFFARX1 I_70741 (I1206165,I3563,I1206049,I1206205,);
not I_70742 (I1206041,I1206205);
not I_70743 (I1206227,I413450);
nand I_70744 (I1206244,I1206148,I1206227);
DFFARX1 I_70745 (I1206244,I3563,I1206049,I1206270,);
not I_70746 (I1206278,I1206270);
not I_70747 (I1206295,I413441);
nand I_70748 (I1206312,I1206295,I413429);
and I_70749 (I1206329,I1206131,I1206312);
nor I_70750 (I1206346,I1206244,I1206329);
DFFARX1 I_70751 (I1206346,I3563,I1206049,I1206017,);
DFFARX1 I_70752 (I1206329,I3563,I1206049,I1206038,);
nor I_70753 (I1206391,I413441,I413435);
nor I_70754 (I1206029,I1206244,I1206391);
or I_70755 (I1206422,I413441,I413435);
nor I_70756 (I1206439,I413432,I413426);
DFFARX1 I_70757 (I1206439,I3563,I1206049,I1206465,);
not I_70758 (I1206473,I1206465);
nor I_70759 (I1206035,I1206473,I1206278);
nand I_70760 (I1206504,I1206473,I1206123);
not I_70761 (I1206521,I413432);
nand I_70762 (I1206538,I1206521,I1206227);
nand I_70763 (I1206555,I1206473,I1206538);
nand I_70764 (I1206026,I1206555,I1206504);
nand I_70765 (I1206023,I1206538,I1206422);
not I_70766 (I1206627,I3570);
DFFARX1 I_70767 (I521410,I3563,I1206627,I1206653,);
and I_70768 (I1206661,I1206653,I521425);
DFFARX1 I_70769 (I1206661,I3563,I1206627,I1206610,);
DFFARX1 I_70770 (I521428,I3563,I1206627,I1206701,);
not I_70771 (I1206709,I521422);
not I_70772 (I1206726,I521437);
nand I_70773 (I1206743,I1206726,I1206709);
nor I_70774 (I1206598,I1206701,I1206743);
DFFARX1 I_70775 (I1206743,I3563,I1206627,I1206783,);
not I_70776 (I1206619,I1206783);
not I_70777 (I1206805,I521413);
nand I_70778 (I1206822,I1206726,I1206805);
DFFARX1 I_70779 (I1206822,I3563,I1206627,I1206848,);
not I_70780 (I1206856,I1206848);
not I_70781 (I1206873,I521416);
nand I_70782 (I1206890,I1206873,I521410);
and I_70783 (I1206907,I1206709,I1206890);
nor I_70784 (I1206924,I1206822,I1206907);
DFFARX1 I_70785 (I1206924,I3563,I1206627,I1206595,);
DFFARX1 I_70786 (I1206907,I3563,I1206627,I1206616,);
nor I_70787 (I1206969,I521416,I521419);
nor I_70788 (I1206607,I1206822,I1206969);
or I_70789 (I1207000,I521416,I521419);
nor I_70790 (I1207017,I521434,I521431);
DFFARX1 I_70791 (I1207017,I3563,I1206627,I1207043,);
not I_70792 (I1207051,I1207043);
nor I_70793 (I1206613,I1207051,I1206856);
nand I_70794 (I1207082,I1207051,I1206701);
not I_70795 (I1207099,I521434);
nand I_70796 (I1207116,I1207099,I1206805);
nand I_70797 (I1207133,I1207051,I1207116);
nand I_70798 (I1206604,I1207133,I1207082);
nand I_70799 (I1206601,I1207116,I1207000);
not I_70800 (I1207205,I3570);
DFFARX1 I_70801 (I191678,I3563,I1207205,I1207231,);
and I_70802 (I1207239,I1207231,I191681);
DFFARX1 I_70803 (I1207239,I3563,I1207205,I1207188,);
DFFARX1 I_70804 (I191681,I3563,I1207205,I1207279,);
not I_70805 (I1207287,I191696);
not I_70806 (I1207304,I191702);
nand I_70807 (I1207321,I1207304,I1207287);
nor I_70808 (I1207176,I1207279,I1207321);
DFFARX1 I_70809 (I1207321,I3563,I1207205,I1207361,);
not I_70810 (I1207197,I1207361);
not I_70811 (I1207383,I191690);
nand I_70812 (I1207400,I1207304,I1207383);
DFFARX1 I_70813 (I1207400,I3563,I1207205,I1207426,);
not I_70814 (I1207434,I1207426);
not I_70815 (I1207451,I191687);
nand I_70816 (I1207468,I1207451,I191684);
and I_70817 (I1207485,I1207287,I1207468);
nor I_70818 (I1207502,I1207400,I1207485);
DFFARX1 I_70819 (I1207502,I3563,I1207205,I1207173,);
DFFARX1 I_70820 (I1207485,I3563,I1207205,I1207194,);
nor I_70821 (I1207547,I191687,I191678);
nor I_70822 (I1207185,I1207400,I1207547);
or I_70823 (I1207578,I191687,I191678);
nor I_70824 (I1207595,I191693,I191699);
DFFARX1 I_70825 (I1207595,I3563,I1207205,I1207621,);
not I_70826 (I1207629,I1207621);
nor I_70827 (I1207191,I1207629,I1207434);
nand I_70828 (I1207660,I1207629,I1207279);
not I_70829 (I1207677,I191693);
nand I_70830 (I1207694,I1207677,I1207383);
nand I_70831 (I1207711,I1207629,I1207694);
nand I_70832 (I1207182,I1207711,I1207660);
nand I_70833 (I1207179,I1207694,I1207578);
not I_70834 (I1207783,I3570);
DFFARX1 I_70835 (I546539,I3563,I1207783,I1207809,);
and I_70836 (I1207817,I1207809,I546554);
DFFARX1 I_70837 (I1207817,I3563,I1207783,I1207766,);
DFFARX1 I_70838 (I546545,I3563,I1207783,I1207857,);
not I_70839 (I1207865,I546539);
not I_70840 (I1207882,I546557);
nand I_70841 (I1207899,I1207882,I1207865);
nor I_70842 (I1207754,I1207857,I1207899);
DFFARX1 I_70843 (I1207899,I3563,I1207783,I1207939,);
not I_70844 (I1207775,I1207939);
not I_70845 (I1207961,I546548);
nand I_70846 (I1207978,I1207882,I1207961);
DFFARX1 I_70847 (I1207978,I3563,I1207783,I1208004,);
not I_70848 (I1208012,I1208004);
not I_70849 (I1208029,I546560);
nand I_70850 (I1208046,I1208029,I546536);
and I_70851 (I1208063,I1207865,I1208046);
nor I_70852 (I1208080,I1207978,I1208063);
DFFARX1 I_70853 (I1208080,I3563,I1207783,I1207751,);
DFFARX1 I_70854 (I1208063,I3563,I1207783,I1207772,);
nor I_70855 (I1208125,I546560,I546536);
nor I_70856 (I1207763,I1207978,I1208125);
or I_70857 (I1208156,I546560,I546536);
nor I_70858 (I1208173,I546542,I546551);
DFFARX1 I_70859 (I1208173,I3563,I1207783,I1208199,);
not I_70860 (I1208207,I1208199);
nor I_70861 (I1207769,I1208207,I1208012);
nand I_70862 (I1208238,I1208207,I1207857);
not I_70863 (I1208255,I546542);
nand I_70864 (I1208272,I1208255,I1207961);
nand I_70865 (I1208289,I1208207,I1208272);
nand I_70866 (I1207760,I1208289,I1208238);
nand I_70867 (I1207757,I1208272,I1208156);
not I_70868 (I1208361,I3570);
DFFARX1 I_70869 (I478978,I3563,I1208361,I1208387,);
and I_70870 (I1208395,I1208387,I478993);
DFFARX1 I_70871 (I1208395,I3563,I1208361,I1208344,);
DFFARX1 I_70872 (I478996,I3563,I1208361,I1208435,);
not I_70873 (I1208443,I478990);
not I_70874 (I1208460,I479005);
nand I_70875 (I1208477,I1208460,I1208443);
nor I_70876 (I1208332,I1208435,I1208477);
DFFARX1 I_70877 (I1208477,I3563,I1208361,I1208517,);
not I_70878 (I1208353,I1208517);
not I_70879 (I1208539,I478981);
nand I_70880 (I1208556,I1208460,I1208539);
DFFARX1 I_70881 (I1208556,I3563,I1208361,I1208582,);
not I_70882 (I1208590,I1208582);
not I_70883 (I1208607,I478984);
nand I_70884 (I1208624,I1208607,I478978);
and I_70885 (I1208641,I1208443,I1208624);
nor I_70886 (I1208658,I1208556,I1208641);
DFFARX1 I_70887 (I1208658,I3563,I1208361,I1208329,);
DFFARX1 I_70888 (I1208641,I3563,I1208361,I1208350,);
nor I_70889 (I1208703,I478984,I478987);
nor I_70890 (I1208341,I1208556,I1208703);
or I_70891 (I1208734,I478984,I478987);
nor I_70892 (I1208751,I479002,I478999);
DFFARX1 I_70893 (I1208751,I3563,I1208361,I1208777,);
not I_70894 (I1208785,I1208777);
nor I_70895 (I1208347,I1208785,I1208590);
nand I_70896 (I1208816,I1208785,I1208435);
not I_70897 (I1208833,I479002);
nand I_70898 (I1208850,I1208833,I1208539);
nand I_70899 (I1208867,I1208785,I1208850);
nand I_70900 (I1208338,I1208867,I1208816);
nand I_70901 (I1208335,I1208850,I1208734);
not I_70902 (I1208939,I3570);
DFFARX1 I_70903 (I188108,I3563,I1208939,I1208965,);
and I_70904 (I1208973,I1208965,I188111);
DFFARX1 I_70905 (I1208973,I3563,I1208939,I1208922,);
DFFARX1 I_70906 (I188111,I3563,I1208939,I1209013,);
not I_70907 (I1209021,I188126);
not I_70908 (I1209038,I188132);
nand I_70909 (I1209055,I1209038,I1209021);
nor I_70910 (I1208910,I1209013,I1209055);
DFFARX1 I_70911 (I1209055,I3563,I1208939,I1209095,);
not I_70912 (I1208931,I1209095);
not I_70913 (I1209117,I188120);
nand I_70914 (I1209134,I1209038,I1209117);
DFFARX1 I_70915 (I1209134,I3563,I1208939,I1209160,);
not I_70916 (I1209168,I1209160);
not I_70917 (I1209185,I188117);
nand I_70918 (I1209202,I1209185,I188114);
and I_70919 (I1209219,I1209021,I1209202);
nor I_70920 (I1209236,I1209134,I1209219);
DFFARX1 I_70921 (I1209236,I3563,I1208939,I1208907,);
DFFARX1 I_70922 (I1209219,I3563,I1208939,I1208928,);
nor I_70923 (I1209281,I188117,I188108);
nor I_70924 (I1208919,I1209134,I1209281);
or I_70925 (I1209312,I188117,I188108);
nor I_70926 (I1209329,I188123,I188129);
DFFARX1 I_70927 (I1209329,I3563,I1208939,I1209355,);
not I_70928 (I1209363,I1209355);
nor I_70929 (I1208925,I1209363,I1209168);
nand I_70930 (I1209394,I1209363,I1209013);
not I_70931 (I1209411,I188123);
nand I_70932 (I1209428,I1209411,I1209117);
nand I_70933 (I1209445,I1209363,I1209428);
nand I_70934 (I1208916,I1209445,I1209394);
nand I_70935 (I1208913,I1209428,I1209312);
not I_70936 (I1209517,I3570);
DFFARX1 I_70937 (I105155,I3563,I1209517,I1209543,);
and I_70938 (I1209551,I1209543,I105131);
DFFARX1 I_70939 (I1209551,I3563,I1209517,I1209500,);
DFFARX1 I_70940 (I105149,I3563,I1209517,I1209591,);
not I_70941 (I1209599,I105137);
not I_70942 (I1209616,I105134);
nand I_70943 (I1209633,I1209616,I1209599);
nor I_70944 (I1209488,I1209591,I1209633);
DFFARX1 I_70945 (I1209633,I3563,I1209517,I1209673,);
not I_70946 (I1209509,I1209673);
not I_70947 (I1209695,I105143);
nand I_70948 (I1209712,I1209616,I1209695);
DFFARX1 I_70949 (I1209712,I3563,I1209517,I1209738,);
not I_70950 (I1209746,I1209738);
not I_70951 (I1209763,I105134);
nand I_70952 (I1209780,I1209763,I105152);
and I_70953 (I1209797,I1209599,I1209780);
nor I_70954 (I1209814,I1209712,I1209797);
DFFARX1 I_70955 (I1209814,I3563,I1209517,I1209485,);
DFFARX1 I_70956 (I1209797,I3563,I1209517,I1209506,);
nor I_70957 (I1209859,I105134,I105146);
nor I_70958 (I1209497,I1209712,I1209859);
or I_70959 (I1209890,I105134,I105146);
nor I_70960 (I1209907,I105140,I105131);
DFFARX1 I_70961 (I1209907,I3563,I1209517,I1209933,);
not I_70962 (I1209941,I1209933);
nor I_70963 (I1209503,I1209941,I1209746);
nand I_70964 (I1209972,I1209941,I1209591);
not I_70965 (I1209989,I105140);
nand I_70966 (I1210006,I1209989,I1209695);
nand I_70967 (I1210023,I1209941,I1210006);
nand I_70968 (I1209494,I1210023,I1209972);
nand I_70969 (I1209491,I1210006,I1209890);
not I_70970 (I1210095,I3570);
DFFARX1 I_70971 (I1340480,I3563,I1210095,I1210121,);
and I_70972 (I1210129,I1210121,I1340462);
DFFARX1 I_70973 (I1210129,I3563,I1210095,I1210078,);
DFFARX1 I_70974 (I1340453,I3563,I1210095,I1210169,);
not I_70975 (I1210177,I1340468);
not I_70976 (I1210194,I1340456);
nand I_70977 (I1210211,I1210194,I1210177);
nor I_70978 (I1210066,I1210169,I1210211);
DFFARX1 I_70979 (I1210211,I3563,I1210095,I1210251,);
not I_70980 (I1210087,I1210251);
not I_70981 (I1210273,I1340465);
nand I_70982 (I1210290,I1210194,I1210273);
DFFARX1 I_70983 (I1210290,I3563,I1210095,I1210316,);
not I_70984 (I1210324,I1210316);
not I_70985 (I1210341,I1340474);
nand I_70986 (I1210358,I1210341,I1340453);
and I_70987 (I1210375,I1210177,I1210358);
nor I_70988 (I1210392,I1210290,I1210375);
DFFARX1 I_70989 (I1210392,I3563,I1210095,I1210063,);
DFFARX1 I_70990 (I1210375,I3563,I1210095,I1210084,);
nor I_70991 (I1210437,I1340474,I1340477);
nor I_70992 (I1210075,I1210290,I1210437);
or I_70993 (I1210468,I1340474,I1340477);
nor I_70994 (I1210485,I1340471,I1340459);
DFFARX1 I_70995 (I1210485,I3563,I1210095,I1210511,);
not I_70996 (I1210519,I1210511);
nor I_70997 (I1210081,I1210519,I1210324);
nand I_70998 (I1210550,I1210519,I1210169);
not I_70999 (I1210567,I1340471);
nand I_71000 (I1210584,I1210567,I1210273);
nand I_71001 (I1210601,I1210519,I1210584);
nand I_71002 (I1210072,I1210601,I1210550);
nand I_71003 (I1210069,I1210584,I1210468);
not I_71004 (I1210673,I3570);
DFFARX1 I_71005 (I29770,I3563,I1210673,I1210699,);
and I_71006 (I1210707,I1210699,I29773);
DFFARX1 I_71007 (I1210707,I3563,I1210673,I1210656,);
DFFARX1 I_71008 (I29773,I3563,I1210673,I1210747,);
not I_71009 (I1210755,I29776);
not I_71010 (I1210772,I29791);
nand I_71011 (I1210789,I1210772,I1210755);
nor I_71012 (I1210644,I1210747,I1210789);
DFFARX1 I_71013 (I1210789,I3563,I1210673,I1210829,);
not I_71014 (I1210665,I1210829);
not I_71015 (I1210851,I29785);
nand I_71016 (I1210868,I1210772,I1210851);
DFFARX1 I_71017 (I1210868,I3563,I1210673,I1210894,);
not I_71018 (I1210902,I1210894);
not I_71019 (I1210919,I29788);
nand I_71020 (I1210936,I1210919,I29770);
and I_71021 (I1210953,I1210755,I1210936);
nor I_71022 (I1210970,I1210868,I1210953);
DFFARX1 I_71023 (I1210970,I3563,I1210673,I1210641,);
DFFARX1 I_71024 (I1210953,I3563,I1210673,I1210662,);
nor I_71025 (I1211015,I29788,I29782);
nor I_71026 (I1210653,I1210868,I1211015);
or I_71027 (I1211046,I29788,I29782);
nor I_71028 (I1211063,I29779,I29794);
DFFARX1 I_71029 (I1211063,I3563,I1210673,I1211089,);
not I_71030 (I1211097,I1211089);
nor I_71031 (I1210659,I1211097,I1210902);
nand I_71032 (I1211128,I1211097,I1210747);
not I_71033 (I1211145,I29779);
nand I_71034 (I1211162,I1211145,I1210851);
nand I_71035 (I1211179,I1211097,I1211162);
nand I_71036 (I1210650,I1211179,I1211128);
nand I_71037 (I1210647,I1211162,I1211046);
not I_71038 (I1211251,I3570);
DFFARX1 I_71039 (I444162,I3563,I1211251,I1211277,);
and I_71040 (I1211285,I1211277,I444177);
DFFARX1 I_71041 (I1211285,I3563,I1211251,I1211234,);
DFFARX1 I_71042 (I444180,I3563,I1211251,I1211325,);
not I_71043 (I1211333,I444174);
not I_71044 (I1211350,I444189);
nand I_71045 (I1211367,I1211350,I1211333);
nor I_71046 (I1211222,I1211325,I1211367);
DFFARX1 I_71047 (I1211367,I3563,I1211251,I1211407,);
not I_71048 (I1211243,I1211407);
not I_71049 (I1211429,I444165);
nand I_71050 (I1211446,I1211350,I1211429);
DFFARX1 I_71051 (I1211446,I3563,I1211251,I1211472,);
not I_71052 (I1211480,I1211472);
not I_71053 (I1211497,I444168);
nand I_71054 (I1211514,I1211497,I444162);
and I_71055 (I1211531,I1211333,I1211514);
nor I_71056 (I1211548,I1211446,I1211531);
DFFARX1 I_71057 (I1211548,I3563,I1211251,I1211219,);
DFFARX1 I_71058 (I1211531,I3563,I1211251,I1211240,);
nor I_71059 (I1211593,I444168,I444171);
nor I_71060 (I1211231,I1211446,I1211593);
or I_71061 (I1211624,I444168,I444171);
nor I_71062 (I1211641,I444186,I444183);
DFFARX1 I_71063 (I1211641,I3563,I1211251,I1211667,);
not I_71064 (I1211675,I1211667);
nor I_71065 (I1211237,I1211675,I1211480);
nand I_71066 (I1211706,I1211675,I1211325);
not I_71067 (I1211723,I444186);
nand I_71068 (I1211740,I1211723,I1211429);
nand I_71069 (I1211757,I1211675,I1211740);
nand I_71070 (I1211228,I1211757,I1211706);
nand I_71071 (I1211225,I1211740,I1211624);
not I_71072 (I1211829,I3570);
DFFARX1 I_71073 (I1359520,I3563,I1211829,I1211855,);
and I_71074 (I1211863,I1211855,I1359502);
DFFARX1 I_71075 (I1211863,I3563,I1211829,I1211812,);
DFFARX1 I_71076 (I1359493,I3563,I1211829,I1211903,);
not I_71077 (I1211911,I1359508);
not I_71078 (I1211928,I1359496);
nand I_71079 (I1211945,I1211928,I1211911);
nor I_71080 (I1211800,I1211903,I1211945);
DFFARX1 I_71081 (I1211945,I3563,I1211829,I1211985,);
not I_71082 (I1211821,I1211985);
not I_71083 (I1212007,I1359505);
nand I_71084 (I1212024,I1211928,I1212007);
DFFARX1 I_71085 (I1212024,I3563,I1211829,I1212050,);
not I_71086 (I1212058,I1212050);
not I_71087 (I1212075,I1359514);
nand I_71088 (I1212092,I1212075,I1359493);
and I_71089 (I1212109,I1211911,I1212092);
nor I_71090 (I1212126,I1212024,I1212109);
DFFARX1 I_71091 (I1212126,I3563,I1211829,I1211797,);
DFFARX1 I_71092 (I1212109,I3563,I1211829,I1211818,);
nor I_71093 (I1212171,I1359514,I1359517);
nor I_71094 (I1211809,I1212024,I1212171);
or I_71095 (I1212202,I1359514,I1359517);
nor I_71096 (I1212219,I1359511,I1359499);
DFFARX1 I_71097 (I1212219,I3563,I1211829,I1212245,);
not I_71098 (I1212253,I1212245);
nor I_71099 (I1211815,I1212253,I1212058);
nand I_71100 (I1212284,I1212253,I1211903);
not I_71101 (I1212301,I1359511);
nand I_71102 (I1212318,I1212301,I1212007);
nand I_71103 (I1212335,I1212253,I1212318);
nand I_71104 (I1211806,I1212335,I1212284);
nand I_71105 (I1211803,I1212318,I1212202);
not I_71106 (I1212407,I3570);
DFFARX1 I_71107 (I246418,I3563,I1212407,I1212433,);
and I_71108 (I1212441,I1212433,I246421);
DFFARX1 I_71109 (I1212441,I3563,I1212407,I1212390,);
DFFARX1 I_71110 (I246421,I3563,I1212407,I1212481,);
not I_71111 (I1212489,I246436);
not I_71112 (I1212506,I246442);
nand I_71113 (I1212523,I1212506,I1212489);
nor I_71114 (I1212378,I1212481,I1212523);
DFFARX1 I_71115 (I1212523,I3563,I1212407,I1212563,);
not I_71116 (I1212399,I1212563);
not I_71117 (I1212585,I246430);
nand I_71118 (I1212602,I1212506,I1212585);
DFFARX1 I_71119 (I1212602,I3563,I1212407,I1212628,);
not I_71120 (I1212636,I1212628);
not I_71121 (I1212653,I246427);
nand I_71122 (I1212670,I1212653,I246424);
and I_71123 (I1212687,I1212489,I1212670);
nor I_71124 (I1212704,I1212602,I1212687);
DFFARX1 I_71125 (I1212704,I3563,I1212407,I1212375,);
DFFARX1 I_71126 (I1212687,I3563,I1212407,I1212396,);
nor I_71127 (I1212749,I246427,I246418);
nor I_71128 (I1212387,I1212602,I1212749);
or I_71129 (I1212780,I246427,I246418);
nor I_71130 (I1212797,I246433,I246439);
DFFARX1 I_71131 (I1212797,I3563,I1212407,I1212823,);
not I_71132 (I1212831,I1212823);
nor I_71133 (I1212393,I1212831,I1212636);
nand I_71134 (I1212862,I1212831,I1212481);
not I_71135 (I1212879,I246433);
nand I_71136 (I1212896,I1212879,I1212585);
nand I_71137 (I1212913,I1212831,I1212896);
nand I_71138 (I1212384,I1212913,I1212862);
nand I_71139 (I1212381,I1212896,I1212780);
not I_71140 (I1212985,I3570);
DFFARX1 I_71141 (I828977,I3563,I1212985,I1213011,);
and I_71142 (I1213019,I1213011,I828983);
DFFARX1 I_71143 (I1213019,I3563,I1212985,I1212968,);
DFFARX1 I_71144 (I828989,I3563,I1212985,I1213059,);
not I_71145 (I1213067,I828974);
not I_71146 (I1213084,I828974);
nand I_71147 (I1213101,I1213084,I1213067);
nor I_71148 (I1212956,I1213059,I1213101);
DFFARX1 I_71149 (I1213101,I3563,I1212985,I1213141,);
not I_71150 (I1212977,I1213141);
not I_71151 (I1213163,I828992);
nand I_71152 (I1213180,I1213084,I1213163);
DFFARX1 I_71153 (I1213180,I3563,I1212985,I1213206,);
not I_71154 (I1213214,I1213206);
not I_71155 (I1213231,I828986);
nand I_71156 (I1213248,I1213231,I828977);
and I_71157 (I1213265,I1213067,I1213248);
nor I_71158 (I1213282,I1213180,I1213265);
DFFARX1 I_71159 (I1213282,I3563,I1212985,I1212953,);
DFFARX1 I_71160 (I1213265,I3563,I1212985,I1212974,);
nor I_71161 (I1213327,I828986,I828995);
nor I_71162 (I1212965,I1213180,I1213327);
or I_71163 (I1213358,I828986,I828995);
nor I_71164 (I1213375,I828980,I828980);
DFFARX1 I_71165 (I1213375,I3563,I1212985,I1213401,);
not I_71166 (I1213409,I1213401);
nor I_71167 (I1212971,I1213409,I1213214);
nand I_71168 (I1213440,I1213409,I1213059);
not I_71169 (I1213457,I828980);
nand I_71170 (I1213474,I1213457,I1213163);
nand I_71171 (I1213491,I1213409,I1213474);
nand I_71172 (I1212962,I1213491,I1213440);
nand I_71173 (I1212959,I1213474,I1213358);
not I_71174 (I1213563,I3570);
DFFARX1 I_71175 (I1039559,I3563,I1213563,I1213589,);
and I_71176 (I1213597,I1213589,I1039553);
DFFARX1 I_71177 (I1213597,I3563,I1213563,I1213546,);
DFFARX1 I_71178 (I1039571,I3563,I1213563,I1213637,);
not I_71179 (I1213645,I1039562);
not I_71180 (I1213662,I1039574);
nand I_71181 (I1213679,I1213662,I1213645);
nor I_71182 (I1213534,I1213637,I1213679);
DFFARX1 I_71183 (I1213679,I3563,I1213563,I1213719,);
not I_71184 (I1213555,I1213719);
not I_71185 (I1213741,I1039580);
nand I_71186 (I1213758,I1213662,I1213741);
DFFARX1 I_71187 (I1213758,I3563,I1213563,I1213784,);
not I_71188 (I1213792,I1213784);
not I_71189 (I1213809,I1039556);
nand I_71190 (I1213826,I1213809,I1039577);
and I_71191 (I1213843,I1213645,I1213826);
nor I_71192 (I1213860,I1213758,I1213843);
DFFARX1 I_71193 (I1213860,I3563,I1213563,I1213531,);
DFFARX1 I_71194 (I1213843,I3563,I1213563,I1213552,);
nor I_71195 (I1213905,I1039556,I1039568);
nor I_71196 (I1213543,I1213758,I1213905);
or I_71197 (I1213936,I1039556,I1039568);
nor I_71198 (I1213953,I1039553,I1039565);
DFFARX1 I_71199 (I1213953,I3563,I1213563,I1213979,);
not I_71200 (I1213987,I1213979);
nor I_71201 (I1213549,I1213987,I1213792);
nand I_71202 (I1214018,I1213987,I1213637);
not I_71203 (I1214035,I1039553);
nand I_71204 (I1214052,I1214035,I1213741);
nand I_71205 (I1214069,I1213987,I1214052);
nand I_71206 (I1213540,I1214069,I1214018);
nand I_71207 (I1213537,I1214052,I1213936);
not I_71208 (I1214141,I3570);
DFFARX1 I_71209 (I916173,I3563,I1214141,I1214167,);
and I_71210 (I1214175,I1214167,I916167);
DFFARX1 I_71211 (I1214175,I3563,I1214141,I1214124,);
DFFARX1 I_71212 (I916185,I3563,I1214141,I1214215,);
not I_71213 (I1214223,I916176);
not I_71214 (I1214240,I916188);
nand I_71215 (I1214257,I1214240,I1214223);
nor I_71216 (I1214112,I1214215,I1214257);
DFFARX1 I_71217 (I1214257,I3563,I1214141,I1214297,);
not I_71218 (I1214133,I1214297);
not I_71219 (I1214319,I916194);
nand I_71220 (I1214336,I1214240,I1214319);
DFFARX1 I_71221 (I1214336,I3563,I1214141,I1214362,);
not I_71222 (I1214370,I1214362);
not I_71223 (I1214387,I916170);
nand I_71224 (I1214404,I1214387,I916191);
and I_71225 (I1214421,I1214223,I1214404);
nor I_71226 (I1214438,I1214336,I1214421);
DFFARX1 I_71227 (I1214438,I3563,I1214141,I1214109,);
DFFARX1 I_71228 (I1214421,I3563,I1214141,I1214130,);
nor I_71229 (I1214483,I916170,I916182);
nor I_71230 (I1214121,I1214336,I1214483);
or I_71231 (I1214514,I916170,I916182);
nor I_71232 (I1214531,I916167,I916179);
DFFARX1 I_71233 (I1214531,I3563,I1214141,I1214557,);
not I_71234 (I1214565,I1214557);
nor I_71235 (I1214127,I1214565,I1214370);
nand I_71236 (I1214596,I1214565,I1214215);
not I_71237 (I1214613,I916167);
nand I_71238 (I1214630,I1214613,I1214319);
nand I_71239 (I1214647,I1214565,I1214630);
nand I_71240 (I1214118,I1214647,I1214596);
nand I_71241 (I1214115,I1214630,I1214514);
not I_71242 (I1214719,I3570);
DFFARX1 I_71243 (I1033745,I3563,I1214719,I1214745,);
and I_71244 (I1214753,I1214745,I1033739);
DFFARX1 I_71245 (I1214753,I3563,I1214719,I1214702,);
DFFARX1 I_71246 (I1033757,I3563,I1214719,I1214793,);
not I_71247 (I1214801,I1033748);
not I_71248 (I1214818,I1033760);
nand I_71249 (I1214835,I1214818,I1214801);
nor I_71250 (I1214690,I1214793,I1214835);
DFFARX1 I_71251 (I1214835,I3563,I1214719,I1214875,);
not I_71252 (I1214711,I1214875);
not I_71253 (I1214897,I1033766);
nand I_71254 (I1214914,I1214818,I1214897);
DFFARX1 I_71255 (I1214914,I3563,I1214719,I1214940,);
not I_71256 (I1214948,I1214940);
not I_71257 (I1214965,I1033742);
nand I_71258 (I1214982,I1214965,I1033763);
and I_71259 (I1214999,I1214801,I1214982);
nor I_71260 (I1215016,I1214914,I1214999);
DFFARX1 I_71261 (I1215016,I3563,I1214719,I1214687,);
DFFARX1 I_71262 (I1214999,I3563,I1214719,I1214708,);
nor I_71263 (I1215061,I1033742,I1033754);
nor I_71264 (I1214699,I1214914,I1215061);
or I_71265 (I1215092,I1033742,I1033754);
nor I_71266 (I1215109,I1033739,I1033751);
DFFARX1 I_71267 (I1215109,I3563,I1214719,I1215135,);
not I_71268 (I1215143,I1215135);
nor I_71269 (I1214705,I1215143,I1214948);
nand I_71270 (I1215174,I1215143,I1214793);
not I_71271 (I1215191,I1033739);
nand I_71272 (I1215208,I1215191,I1214897);
nand I_71273 (I1215225,I1215143,I1215208);
nand I_71274 (I1214696,I1215225,I1215174);
nand I_71275 (I1214693,I1215208,I1215092);
not I_71276 (I1215297,I3570);
DFFARX1 I_71277 (I1246430,I3563,I1215297,I1215323,);
and I_71278 (I1215331,I1215323,I1246424);
DFFARX1 I_71279 (I1215331,I3563,I1215297,I1215280,);
DFFARX1 I_71280 (I1246409,I3563,I1215297,I1215371,);
not I_71281 (I1215379,I1246415);
not I_71282 (I1215396,I1246427);
nand I_71283 (I1215413,I1215396,I1215379);
nor I_71284 (I1215268,I1215371,I1215413);
DFFARX1 I_71285 (I1215413,I3563,I1215297,I1215453,);
not I_71286 (I1215289,I1215453);
not I_71287 (I1215475,I1246409);
nand I_71288 (I1215492,I1215396,I1215475);
DFFARX1 I_71289 (I1215492,I3563,I1215297,I1215518,);
not I_71290 (I1215526,I1215518);
not I_71291 (I1215543,I1246433);
nand I_71292 (I1215560,I1215543,I1246421);
and I_71293 (I1215577,I1215379,I1215560);
nor I_71294 (I1215594,I1215492,I1215577);
DFFARX1 I_71295 (I1215594,I3563,I1215297,I1215265,);
DFFARX1 I_71296 (I1215577,I3563,I1215297,I1215286,);
nor I_71297 (I1215639,I1246433,I1246412);
nor I_71298 (I1215277,I1215492,I1215639);
or I_71299 (I1215670,I1246433,I1246412);
nor I_71300 (I1215687,I1246418,I1246412);
DFFARX1 I_71301 (I1215687,I3563,I1215297,I1215713,);
not I_71302 (I1215721,I1215713);
nor I_71303 (I1215283,I1215721,I1215526);
nand I_71304 (I1215752,I1215721,I1215371);
not I_71305 (I1215769,I1246418);
nand I_71306 (I1215786,I1215769,I1215475);
nand I_71307 (I1215803,I1215721,I1215786);
nand I_71308 (I1215274,I1215803,I1215752);
nand I_71309 (I1215271,I1215786,I1215670);
not I_71310 (I1215875,I3570);
DFFARX1 I_71311 (I1337505,I3563,I1215875,I1215901,);
and I_71312 (I1215909,I1215901,I1337487);
DFFARX1 I_71313 (I1215909,I3563,I1215875,I1215858,);
DFFARX1 I_71314 (I1337478,I3563,I1215875,I1215949,);
not I_71315 (I1215957,I1337493);
not I_71316 (I1215974,I1337481);
nand I_71317 (I1215991,I1215974,I1215957);
nor I_71318 (I1215846,I1215949,I1215991);
DFFARX1 I_71319 (I1215991,I3563,I1215875,I1216031,);
not I_71320 (I1215867,I1216031);
not I_71321 (I1216053,I1337490);
nand I_71322 (I1216070,I1215974,I1216053);
DFFARX1 I_71323 (I1216070,I3563,I1215875,I1216096,);
not I_71324 (I1216104,I1216096);
not I_71325 (I1216121,I1337499);
nand I_71326 (I1216138,I1216121,I1337478);
and I_71327 (I1216155,I1215957,I1216138);
nor I_71328 (I1216172,I1216070,I1216155);
DFFARX1 I_71329 (I1216172,I3563,I1215875,I1215843,);
DFFARX1 I_71330 (I1216155,I3563,I1215875,I1215864,);
nor I_71331 (I1216217,I1337499,I1337502);
nor I_71332 (I1215855,I1216070,I1216217);
or I_71333 (I1216248,I1337499,I1337502);
nor I_71334 (I1216265,I1337496,I1337484);
DFFARX1 I_71335 (I1216265,I3563,I1215875,I1216291,);
not I_71336 (I1216299,I1216291);
nor I_71337 (I1215861,I1216299,I1216104);
nand I_71338 (I1216330,I1216299,I1215949);
not I_71339 (I1216347,I1337496);
nand I_71340 (I1216364,I1216347,I1216053);
nand I_71341 (I1216381,I1216299,I1216364);
nand I_71342 (I1215852,I1216381,I1216330);
nand I_71343 (I1215849,I1216364,I1216248);
not I_71344 (I1216453,I3570);
DFFARX1 I_71345 (I1356545,I3563,I1216453,I1216479,);
and I_71346 (I1216487,I1216479,I1356527);
DFFARX1 I_71347 (I1216487,I3563,I1216453,I1216436,);
DFFARX1 I_71348 (I1356518,I3563,I1216453,I1216527,);
not I_71349 (I1216535,I1356533);
not I_71350 (I1216552,I1356521);
nand I_71351 (I1216569,I1216552,I1216535);
nor I_71352 (I1216424,I1216527,I1216569);
DFFARX1 I_71353 (I1216569,I3563,I1216453,I1216609,);
not I_71354 (I1216445,I1216609);
not I_71355 (I1216631,I1356530);
nand I_71356 (I1216648,I1216552,I1216631);
DFFARX1 I_71357 (I1216648,I3563,I1216453,I1216674,);
not I_71358 (I1216682,I1216674);
not I_71359 (I1216699,I1356539);
nand I_71360 (I1216716,I1216699,I1356518);
and I_71361 (I1216733,I1216535,I1216716);
nor I_71362 (I1216750,I1216648,I1216733);
DFFARX1 I_71363 (I1216750,I3563,I1216453,I1216421,);
DFFARX1 I_71364 (I1216733,I3563,I1216453,I1216442,);
nor I_71365 (I1216795,I1356539,I1356542);
nor I_71366 (I1216433,I1216648,I1216795);
or I_71367 (I1216826,I1356539,I1356542);
nor I_71368 (I1216843,I1356536,I1356524);
DFFARX1 I_71369 (I1216843,I3563,I1216453,I1216869,);
not I_71370 (I1216877,I1216869);
nor I_71371 (I1216439,I1216877,I1216682);
nand I_71372 (I1216908,I1216877,I1216527);
not I_71373 (I1216925,I1356536);
nand I_71374 (I1216942,I1216925,I1216631);
nand I_71375 (I1216959,I1216877,I1216942);
nand I_71376 (I1216430,I1216959,I1216908);
nand I_71377 (I1216427,I1216942,I1216826);
not I_71378 (I1217031,I3570);
DFFARX1 I_71379 (I1036329,I3563,I1217031,I1217057,);
and I_71380 (I1217065,I1217057,I1036323);
DFFARX1 I_71381 (I1217065,I3563,I1217031,I1217014,);
DFFARX1 I_71382 (I1036341,I3563,I1217031,I1217105,);
not I_71383 (I1217113,I1036332);
not I_71384 (I1217130,I1036344);
nand I_71385 (I1217147,I1217130,I1217113);
nor I_71386 (I1217002,I1217105,I1217147);
DFFARX1 I_71387 (I1217147,I3563,I1217031,I1217187,);
not I_71388 (I1217023,I1217187);
not I_71389 (I1217209,I1036350);
nand I_71390 (I1217226,I1217130,I1217209);
DFFARX1 I_71391 (I1217226,I3563,I1217031,I1217252,);
not I_71392 (I1217260,I1217252);
not I_71393 (I1217277,I1036326);
nand I_71394 (I1217294,I1217277,I1036347);
and I_71395 (I1217311,I1217113,I1217294);
nor I_71396 (I1217328,I1217226,I1217311);
DFFARX1 I_71397 (I1217328,I3563,I1217031,I1216999,);
DFFARX1 I_71398 (I1217311,I3563,I1217031,I1217020,);
nor I_71399 (I1217373,I1036326,I1036338);
nor I_71400 (I1217011,I1217226,I1217373);
or I_71401 (I1217404,I1036326,I1036338);
nor I_71402 (I1217421,I1036323,I1036335);
DFFARX1 I_71403 (I1217421,I3563,I1217031,I1217447,);
not I_71404 (I1217455,I1217447);
nor I_71405 (I1217017,I1217455,I1217260);
nand I_71406 (I1217486,I1217455,I1217105);
not I_71407 (I1217503,I1036323);
nand I_71408 (I1217520,I1217503,I1217209);
nand I_71409 (I1217537,I1217455,I1217520);
nand I_71410 (I1217008,I1217537,I1217486);
nand I_71411 (I1217005,I1217520,I1217404);
not I_71412 (I1217609,I3570);
DFFARX1 I_71413 (I348632,I3563,I1217609,I1217635,);
and I_71414 (I1217643,I1217635,I348617);
DFFARX1 I_71415 (I1217643,I3563,I1217609,I1217592,);
DFFARX1 I_71416 (I348623,I3563,I1217609,I1217683,);
not I_71417 (I1217691,I348605);
not I_71418 (I1217708,I348626);
nand I_71419 (I1217725,I1217708,I1217691);
nor I_71420 (I1217580,I1217683,I1217725);
DFFARX1 I_71421 (I1217725,I3563,I1217609,I1217765,);
not I_71422 (I1217601,I1217765);
not I_71423 (I1217787,I348629);
nand I_71424 (I1217804,I1217708,I1217787);
DFFARX1 I_71425 (I1217804,I3563,I1217609,I1217830,);
not I_71426 (I1217838,I1217830);
not I_71427 (I1217855,I348620);
nand I_71428 (I1217872,I1217855,I348608);
and I_71429 (I1217889,I1217691,I1217872);
nor I_71430 (I1217906,I1217804,I1217889);
DFFARX1 I_71431 (I1217906,I3563,I1217609,I1217577,);
DFFARX1 I_71432 (I1217889,I3563,I1217609,I1217598,);
nor I_71433 (I1217951,I348620,I348614);
nor I_71434 (I1217589,I1217804,I1217951);
or I_71435 (I1217982,I348620,I348614);
nor I_71436 (I1217999,I348611,I348605);
DFFARX1 I_71437 (I1217999,I3563,I1217609,I1218025,);
not I_71438 (I1218033,I1218025);
nor I_71439 (I1217595,I1218033,I1217838);
nand I_71440 (I1218064,I1218033,I1217683);
not I_71441 (I1218081,I348611);
nand I_71442 (I1218098,I1218081,I1217787);
nand I_71443 (I1218115,I1218033,I1218098);
nand I_71444 (I1217586,I1218115,I1218064);
nand I_71445 (I1217583,I1218098,I1217982);
not I_71446 (I1218187,I3570);
DFFARX1 I_71447 (I230353,I3563,I1218187,I1218213,);
and I_71448 (I1218221,I1218213,I230356);
DFFARX1 I_71449 (I1218221,I3563,I1218187,I1218170,);
DFFARX1 I_71450 (I230356,I3563,I1218187,I1218261,);
not I_71451 (I1218269,I230371);
not I_71452 (I1218286,I230377);
nand I_71453 (I1218303,I1218286,I1218269);
nor I_71454 (I1218158,I1218261,I1218303);
DFFARX1 I_71455 (I1218303,I3563,I1218187,I1218343,);
not I_71456 (I1218179,I1218343);
not I_71457 (I1218365,I230365);
nand I_71458 (I1218382,I1218286,I1218365);
DFFARX1 I_71459 (I1218382,I3563,I1218187,I1218408,);
not I_71460 (I1218416,I1218408);
not I_71461 (I1218433,I230362);
nand I_71462 (I1218450,I1218433,I230359);
and I_71463 (I1218467,I1218269,I1218450);
nor I_71464 (I1218484,I1218382,I1218467);
DFFARX1 I_71465 (I1218484,I3563,I1218187,I1218155,);
DFFARX1 I_71466 (I1218467,I3563,I1218187,I1218176,);
nor I_71467 (I1218529,I230362,I230353);
nor I_71468 (I1218167,I1218382,I1218529);
or I_71469 (I1218560,I230362,I230353);
nor I_71470 (I1218577,I230368,I230374);
DFFARX1 I_71471 (I1218577,I3563,I1218187,I1218603,);
not I_71472 (I1218611,I1218603);
nor I_71473 (I1218173,I1218611,I1218416);
nand I_71474 (I1218642,I1218611,I1218261);
not I_71475 (I1218659,I230368);
nand I_71476 (I1218676,I1218659,I1218365);
nand I_71477 (I1218693,I1218611,I1218676);
nand I_71478 (I1218164,I1218693,I1218642);
nand I_71479 (I1218161,I1218676,I1218560);
not I_71480 (I1218765,I3570);
DFFARX1 I_71481 (I387103,I3563,I1218765,I1218791,);
and I_71482 (I1218799,I1218791,I387088);
DFFARX1 I_71483 (I1218799,I3563,I1218765,I1218748,);
DFFARX1 I_71484 (I387094,I3563,I1218765,I1218839,);
not I_71485 (I1218847,I387076);
not I_71486 (I1218864,I387097);
nand I_71487 (I1218881,I1218864,I1218847);
nor I_71488 (I1218736,I1218839,I1218881);
DFFARX1 I_71489 (I1218881,I3563,I1218765,I1218921,);
not I_71490 (I1218757,I1218921);
not I_71491 (I1218943,I387100);
nand I_71492 (I1218960,I1218864,I1218943);
DFFARX1 I_71493 (I1218960,I3563,I1218765,I1218986,);
not I_71494 (I1218994,I1218986);
not I_71495 (I1219011,I387091);
nand I_71496 (I1219028,I1219011,I387079);
and I_71497 (I1219045,I1218847,I1219028);
nor I_71498 (I1219062,I1218960,I1219045);
DFFARX1 I_71499 (I1219062,I3563,I1218765,I1218733,);
DFFARX1 I_71500 (I1219045,I3563,I1218765,I1218754,);
nor I_71501 (I1219107,I387091,I387085);
nor I_71502 (I1218745,I1218960,I1219107);
or I_71503 (I1219138,I387091,I387085);
nor I_71504 (I1219155,I387082,I387076);
DFFARX1 I_71505 (I1219155,I3563,I1218765,I1219181,);
not I_71506 (I1219189,I1219181);
nor I_71507 (I1218751,I1219189,I1218994);
nand I_71508 (I1219220,I1219189,I1218839);
not I_71509 (I1219237,I387082);
nand I_71510 (I1219254,I1219237,I1218943);
nand I_71511 (I1219271,I1219189,I1219254);
nand I_71512 (I1218742,I1219271,I1219220);
nand I_71513 (I1218739,I1219254,I1219138);
not I_71514 (I1219343,I3570);
DFFARX1 I_71515 (I213098,I3563,I1219343,I1219369,);
and I_71516 (I1219377,I1219369,I213101);
DFFARX1 I_71517 (I1219377,I3563,I1219343,I1219326,);
DFFARX1 I_71518 (I213101,I3563,I1219343,I1219417,);
not I_71519 (I1219425,I213116);
not I_71520 (I1219442,I213122);
nand I_71521 (I1219459,I1219442,I1219425);
nor I_71522 (I1219314,I1219417,I1219459);
DFFARX1 I_71523 (I1219459,I3563,I1219343,I1219499,);
not I_71524 (I1219335,I1219499);
not I_71525 (I1219521,I213110);
nand I_71526 (I1219538,I1219442,I1219521);
DFFARX1 I_71527 (I1219538,I3563,I1219343,I1219564,);
not I_71528 (I1219572,I1219564);
not I_71529 (I1219589,I213107);
nand I_71530 (I1219606,I1219589,I213104);
and I_71531 (I1219623,I1219425,I1219606);
nor I_71532 (I1219640,I1219538,I1219623);
DFFARX1 I_71533 (I1219640,I3563,I1219343,I1219311,);
DFFARX1 I_71534 (I1219623,I3563,I1219343,I1219332,);
nor I_71535 (I1219685,I213107,I213098);
nor I_71536 (I1219323,I1219538,I1219685);
or I_71537 (I1219716,I213107,I213098);
nor I_71538 (I1219733,I213113,I213119);
DFFARX1 I_71539 (I1219733,I3563,I1219343,I1219759,);
not I_71540 (I1219767,I1219759);
nor I_71541 (I1219329,I1219767,I1219572);
nand I_71542 (I1219798,I1219767,I1219417);
not I_71543 (I1219815,I213113);
nand I_71544 (I1219832,I1219815,I1219521);
nand I_71545 (I1219849,I1219767,I1219832);
nand I_71546 (I1219320,I1219849,I1219798);
nand I_71547 (I1219317,I1219832,I1219716);
not I_71548 (I1219921,I3570);
DFFARX1 I_71549 (I585022,I3563,I1219921,I1219947,);
and I_71550 (I1219955,I1219947,I585010);
DFFARX1 I_71551 (I1219955,I3563,I1219921,I1219904,);
DFFARX1 I_71552 (I585025,I3563,I1219921,I1219995,);
not I_71553 (I1220003,I585016);
not I_71554 (I1220020,I585007);
nand I_71555 (I1220037,I1220020,I1220003);
nor I_71556 (I1219892,I1219995,I1220037);
DFFARX1 I_71557 (I1220037,I3563,I1219921,I1220077,);
not I_71558 (I1219913,I1220077);
not I_71559 (I1220099,I585013);
nand I_71560 (I1220116,I1220020,I1220099);
DFFARX1 I_71561 (I1220116,I3563,I1219921,I1220142,);
not I_71562 (I1220150,I1220142);
not I_71563 (I1220167,I585028);
nand I_71564 (I1220184,I1220167,I585031);
and I_71565 (I1220201,I1220003,I1220184);
nor I_71566 (I1220218,I1220116,I1220201);
DFFARX1 I_71567 (I1220218,I3563,I1219921,I1219889,);
DFFARX1 I_71568 (I1220201,I3563,I1219921,I1219910,);
nor I_71569 (I1220263,I585028,I585007);
nor I_71570 (I1219901,I1220116,I1220263);
or I_71571 (I1220294,I585028,I585007);
nor I_71572 (I1220311,I585019,I585010);
DFFARX1 I_71573 (I1220311,I3563,I1219921,I1220337,);
not I_71574 (I1220345,I1220337);
nor I_71575 (I1219907,I1220345,I1220150);
nand I_71576 (I1220376,I1220345,I1219995);
not I_71577 (I1220393,I585019);
nand I_71578 (I1220410,I1220393,I1220099);
nand I_71579 (I1220427,I1220345,I1220410);
nand I_71580 (I1219898,I1220427,I1220376);
nand I_71581 (I1219895,I1220410,I1220294);
not I_71582 (I1220499,I3570);
DFFARX1 I_71583 (I1366065,I3563,I1220499,I1220525,);
and I_71584 (I1220533,I1220525,I1366047);
DFFARX1 I_71585 (I1220533,I3563,I1220499,I1220482,);
DFFARX1 I_71586 (I1366038,I3563,I1220499,I1220573,);
not I_71587 (I1220581,I1366053);
not I_71588 (I1220598,I1366041);
nand I_71589 (I1220615,I1220598,I1220581);
nor I_71590 (I1220470,I1220573,I1220615);
DFFARX1 I_71591 (I1220615,I3563,I1220499,I1220655,);
not I_71592 (I1220491,I1220655);
not I_71593 (I1220677,I1366050);
nand I_71594 (I1220694,I1220598,I1220677);
DFFARX1 I_71595 (I1220694,I3563,I1220499,I1220720,);
not I_71596 (I1220728,I1220720);
not I_71597 (I1220745,I1366059);
nand I_71598 (I1220762,I1220745,I1366038);
and I_71599 (I1220779,I1220581,I1220762);
nor I_71600 (I1220796,I1220694,I1220779);
DFFARX1 I_71601 (I1220796,I3563,I1220499,I1220467,);
DFFARX1 I_71602 (I1220779,I3563,I1220499,I1220488,);
nor I_71603 (I1220841,I1366059,I1366062);
nor I_71604 (I1220479,I1220694,I1220841);
or I_71605 (I1220872,I1366059,I1366062);
nor I_71606 (I1220889,I1366056,I1366044);
DFFARX1 I_71607 (I1220889,I3563,I1220499,I1220915,);
not I_71608 (I1220923,I1220915);
nor I_71609 (I1220485,I1220923,I1220728);
nand I_71610 (I1220954,I1220923,I1220573);
not I_71611 (I1220971,I1366056);
nand I_71612 (I1220988,I1220971,I1220677);
nand I_71613 (I1221005,I1220923,I1220988);
nand I_71614 (I1220476,I1221005,I1220954);
nand I_71615 (I1220473,I1220988,I1220872);
not I_71616 (I1221077,I3570);
DFFARX1 I_71617 (I572124,I3563,I1221077,I1221103,);
and I_71618 (I1221111,I1221103,I572139);
DFFARX1 I_71619 (I1221111,I3563,I1221077,I1221060,);
DFFARX1 I_71620 (I572130,I3563,I1221077,I1221151,);
not I_71621 (I1221159,I572124);
not I_71622 (I1221176,I572142);
nand I_71623 (I1221193,I1221176,I1221159);
nor I_71624 (I1221048,I1221151,I1221193);
DFFARX1 I_71625 (I1221193,I3563,I1221077,I1221233,);
not I_71626 (I1221069,I1221233);
not I_71627 (I1221255,I572133);
nand I_71628 (I1221272,I1221176,I1221255);
DFFARX1 I_71629 (I1221272,I3563,I1221077,I1221298,);
not I_71630 (I1221306,I1221298);
not I_71631 (I1221323,I572145);
nand I_71632 (I1221340,I1221323,I572121);
and I_71633 (I1221357,I1221159,I1221340);
nor I_71634 (I1221374,I1221272,I1221357);
DFFARX1 I_71635 (I1221374,I3563,I1221077,I1221045,);
DFFARX1 I_71636 (I1221357,I3563,I1221077,I1221066,);
nor I_71637 (I1221419,I572145,I572121);
nor I_71638 (I1221057,I1221272,I1221419);
or I_71639 (I1221450,I572145,I572121);
nor I_71640 (I1221467,I572127,I572136);
DFFARX1 I_71641 (I1221467,I3563,I1221077,I1221493,);
not I_71642 (I1221501,I1221493);
nor I_71643 (I1221063,I1221501,I1221306);
nand I_71644 (I1221532,I1221501,I1221151);
not I_71645 (I1221549,I572127);
nand I_71646 (I1221566,I1221549,I1221255);
nand I_71647 (I1221583,I1221501,I1221566);
nand I_71648 (I1221054,I1221583,I1221532);
nand I_71649 (I1221051,I1221566,I1221450);
not I_71650 (I1221655,I3570);
DFFARX1 I_71651 (I1303961,I3563,I1221655,I1221681,);
and I_71652 (I1221689,I1221681,I1303943);
DFFARX1 I_71653 (I1221689,I3563,I1221655,I1221638,);
DFFARX1 I_71654 (I1303952,I3563,I1221655,I1221729,);
not I_71655 (I1221737,I1303937);
not I_71656 (I1221754,I1303949);
nand I_71657 (I1221771,I1221754,I1221737);
nor I_71658 (I1221626,I1221729,I1221771);
DFFARX1 I_71659 (I1221771,I3563,I1221655,I1221811,);
not I_71660 (I1221647,I1221811);
not I_71661 (I1221833,I1303940);
nand I_71662 (I1221850,I1221754,I1221833);
DFFARX1 I_71663 (I1221850,I3563,I1221655,I1221876,);
not I_71664 (I1221884,I1221876);
not I_71665 (I1221901,I1303937);
nand I_71666 (I1221918,I1221901,I1303940);
and I_71667 (I1221935,I1221737,I1221918);
nor I_71668 (I1221952,I1221850,I1221935);
DFFARX1 I_71669 (I1221952,I3563,I1221655,I1221623,);
DFFARX1 I_71670 (I1221935,I3563,I1221655,I1221644,);
nor I_71671 (I1221997,I1303937,I1303958);
nor I_71672 (I1221635,I1221850,I1221997);
or I_71673 (I1222028,I1303937,I1303958);
nor I_71674 (I1222045,I1303946,I1303955);
DFFARX1 I_71675 (I1222045,I3563,I1221655,I1222071,);
not I_71676 (I1222079,I1222071);
nor I_71677 (I1221641,I1222079,I1221884);
nand I_71678 (I1222110,I1222079,I1221729);
not I_71679 (I1222127,I1303946);
nand I_71680 (I1222144,I1222127,I1221833);
nand I_71681 (I1222161,I1222079,I1222144);
nand I_71682 (I1221632,I1222161,I1222110);
nand I_71683 (I1221629,I1222144,I1222028);
not I_71684 (I1222233,I3570);
DFFARX1 I_71685 (I648602,I3563,I1222233,I1222259,);
and I_71686 (I1222267,I1222259,I648590);
DFFARX1 I_71687 (I1222267,I3563,I1222233,I1222216,);
DFFARX1 I_71688 (I648605,I3563,I1222233,I1222307,);
not I_71689 (I1222315,I648596);
not I_71690 (I1222332,I648587);
nand I_71691 (I1222349,I1222332,I1222315);
nor I_71692 (I1222204,I1222307,I1222349);
DFFARX1 I_71693 (I1222349,I3563,I1222233,I1222389,);
not I_71694 (I1222225,I1222389);
not I_71695 (I1222411,I648593);
nand I_71696 (I1222428,I1222332,I1222411);
DFFARX1 I_71697 (I1222428,I3563,I1222233,I1222454,);
not I_71698 (I1222462,I1222454);
not I_71699 (I1222479,I648608);
nand I_71700 (I1222496,I1222479,I648611);
and I_71701 (I1222513,I1222315,I1222496);
nor I_71702 (I1222530,I1222428,I1222513);
DFFARX1 I_71703 (I1222530,I3563,I1222233,I1222201,);
DFFARX1 I_71704 (I1222513,I3563,I1222233,I1222222,);
nor I_71705 (I1222575,I648608,I648587);
nor I_71706 (I1222213,I1222428,I1222575);
or I_71707 (I1222606,I648608,I648587);
nor I_71708 (I1222623,I648599,I648590);
DFFARX1 I_71709 (I1222623,I3563,I1222233,I1222649,);
not I_71710 (I1222657,I1222649);
nor I_71711 (I1222219,I1222657,I1222462);
nand I_71712 (I1222688,I1222657,I1222307);
not I_71713 (I1222705,I648599);
nand I_71714 (I1222722,I1222705,I1222411);
nand I_71715 (I1222739,I1222657,I1222722);
nand I_71716 (I1222210,I1222739,I1222688);
nand I_71717 (I1222207,I1222722,I1222606);
not I_71718 (I1222811,I3570);
DFFARX1 I_71719 (I923925,I3563,I1222811,I1222837,);
and I_71720 (I1222845,I1222837,I923919);
DFFARX1 I_71721 (I1222845,I3563,I1222811,I1222794,);
DFFARX1 I_71722 (I923937,I3563,I1222811,I1222885,);
not I_71723 (I1222893,I923928);
not I_71724 (I1222910,I923940);
nand I_71725 (I1222927,I1222910,I1222893);
nor I_71726 (I1222782,I1222885,I1222927);
DFFARX1 I_71727 (I1222927,I3563,I1222811,I1222967,);
not I_71728 (I1222803,I1222967);
not I_71729 (I1222989,I923946);
nand I_71730 (I1223006,I1222910,I1222989);
DFFARX1 I_71731 (I1223006,I3563,I1222811,I1223032,);
not I_71732 (I1223040,I1223032);
not I_71733 (I1223057,I923922);
nand I_71734 (I1223074,I1223057,I923943);
and I_71735 (I1223091,I1222893,I1223074);
nor I_71736 (I1223108,I1223006,I1223091);
DFFARX1 I_71737 (I1223108,I3563,I1222811,I1222779,);
DFFARX1 I_71738 (I1223091,I3563,I1222811,I1222800,);
nor I_71739 (I1223153,I923922,I923934);
nor I_71740 (I1222791,I1223006,I1223153);
or I_71741 (I1223184,I923922,I923934);
nor I_71742 (I1223201,I923919,I923931);
DFFARX1 I_71743 (I1223201,I3563,I1222811,I1223227,);
not I_71744 (I1223235,I1223227);
nor I_71745 (I1222797,I1223235,I1223040);
nand I_71746 (I1223266,I1223235,I1222885);
not I_71747 (I1223283,I923919);
nand I_71748 (I1223300,I1223283,I1222989);
nand I_71749 (I1223317,I1223235,I1223300);
nand I_71750 (I1222788,I1223317,I1223266);
nand I_71751 (I1222785,I1223300,I1223184);
not I_71752 (I1223389,I3570);
DFFARX1 I_71753 (I789056,I3563,I1223389,I1223415,);
and I_71754 (I1223423,I1223415,I789044);
DFFARX1 I_71755 (I1223423,I3563,I1223389,I1223372,);
DFFARX1 I_71756 (I789047,I3563,I1223389,I1223463,);
not I_71757 (I1223471,I789041);
not I_71758 (I1223488,I789065);
nand I_71759 (I1223505,I1223488,I1223471);
nor I_71760 (I1223360,I1223463,I1223505);
DFFARX1 I_71761 (I1223505,I3563,I1223389,I1223545,);
not I_71762 (I1223381,I1223545);
not I_71763 (I1223567,I789053);
nand I_71764 (I1223584,I1223488,I1223567);
DFFARX1 I_71765 (I1223584,I3563,I1223389,I1223610,);
not I_71766 (I1223618,I1223610);
not I_71767 (I1223635,I789062);
nand I_71768 (I1223652,I1223635,I789059);
and I_71769 (I1223669,I1223471,I1223652);
nor I_71770 (I1223686,I1223584,I1223669);
DFFARX1 I_71771 (I1223686,I3563,I1223389,I1223357,);
DFFARX1 I_71772 (I1223669,I3563,I1223389,I1223378,);
nor I_71773 (I1223731,I789062,I789050);
nor I_71774 (I1223369,I1223584,I1223731);
or I_71775 (I1223762,I789062,I789050);
nor I_71776 (I1223779,I789041,I789044);
DFFARX1 I_71777 (I1223779,I3563,I1223389,I1223805,);
not I_71778 (I1223813,I1223805);
nor I_71779 (I1223375,I1223813,I1223618);
nand I_71780 (I1223844,I1223813,I1223463);
not I_71781 (I1223861,I789041);
nand I_71782 (I1223878,I1223861,I1223567);
nand I_71783 (I1223895,I1223813,I1223878);
nand I_71784 (I1223366,I1223895,I1223844);
nand I_71785 (I1223363,I1223878,I1223762);
not I_71786 (I1223967,I3570);
DFFARX1 I_71787 (I704090,I3563,I1223967,I1223993,);
and I_71788 (I1224001,I1223993,I704078);
DFFARX1 I_71789 (I1224001,I3563,I1223967,I1223950,);
DFFARX1 I_71790 (I704081,I3563,I1223967,I1224041,);
not I_71791 (I1224049,I704075);
not I_71792 (I1224066,I704099);
nand I_71793 (I1224083,I1224066,I1224049);
nor I_71794 (I1223938,I1224041,I1224083);
DFFARX1 I_71795 (I1224083,I3563,I1223967,I1224123,);
not I_71796 (I1223959,I1224123);
not I_71797 (I1224145,I704087);
nand I_71798 (I1224162,I1224066,I1224145);
DFFARX1 I_71799 (I1224162,I3563,I1223967,I1224188,);
not I_71800 (I1224196,I1224188);
not I_71801 (I1224213,I704096);
nand I_71802 (I1224230,I1224213,I704093);
and I_71803 (I1224247,I1224049,I1224230);
nor I_71804 (I1224264,I1224162,I1224247);
DFFARX1 I_71805 (I1224264,I3563,I1223967,I1223935,);
DFFARX1 I_71806 (I1224247,I3563,I1223967,I1223956,);
nor I_71807 (I1224309,I704096,I704084);
nor I_71808 (I1223947,I1224162,I1224309);
or I_71809 (I1224340,I704096,I704084);
nor I_71810 (I1224357,I704075,I704078);
DFFARX1 I_71811 (I1224357,I3563,I1223967,I1224383,);
not I_71812 (I1224391,I1224383);
nor I_71813 (I1223953,I1224391,I1224196);
nand I_71814 (I1224422,I1224391,I1224041);
not I_71815 (I1224439,I704075);
nand I_71816 (I1224456,I1224439,I1224145);
nand I_71817 (I1224473,I1224391,I1224456);
nand I_71818 (I1223944,I1224473,I1224422);
nand I_71819 (I1223941,I1224456,I1224340);
not I_71820 (I1224545,I3570);
DFFARX1 I_71821 (I224403,I3563,I1224545,I1224571,);
and I_71822 (I1224579,I1224571,I224406);
DFFARX1 I_71823 (I1224579,I3563,I1224545,I1224528,);
DFFARX1 I_71824 (I224406,I3563,I1224545,I1224619,);
not I_71825 (I1224627,I224421);
not I_71826 (I1224644,I224427);
nand I_71827 (I1224661,I1224644,I1224627);
nor I_71828 (I1224516,I1224619,I1224661);
DFFARX1 I_71829 (I1224661,I3563,I1224545,I1224701,);
not I_71830 (I1224537,I1224701);
not I_71831 (I1224723,I224415);
nand I_71832 (I1224740,I1224644,I1224723);
DFFARX1 I_71833 (I1224740,I3563,I1224545,I1224766,);
not I_71834 (I1224774,I1224766);
not I_71835 (I1224791,I224412);
nand I_71836 (I1224808,I1224791,I224409);
and I_71837 (I1224825,I1224627,I1224808);
nor I_71838 (I1224842,I1224740,I1224825);
DFFARX1 I_71839 (I1224842,I3563,I1224545,I1224513,);
DFFARX1 I_71840 (I1224825,I3563,I1224545,I1224534,);
nor I_71841 (I1224887,I224412,I224403);
nor I_71842 (I1224525,I1224740,I1224887);
or I_71843 (I1224918,I224412,I224403);
nor I_71844 (I1224935,I224418,I224424);
DFFARX1 I_71845 (I1224935,I3563,I1224545,I1224961,);
not I_71846 (I1224969,I1224961);
nor I_71847 (I1224531,I1224969,I1224774);
nand I_71848 (I1225000,I1224969,I1224619);
not I_71849 (I1225017,I224418);
nand I_71850 (I1225034,I1225017,I1224723);
nand I_71851 (I1225051,I1224969,I1225034);
nand I_71852 (I1224522,I1225051,I1225000);
nand I_71853 (I1224519,I1225034,I1224918);
not I_71854 (I1225123,I3570);
DFFARX1 I_71855 (I1367255,I3563,I1225123,I1225149,);
and I_71856 (I1225157,I1225149,I1367237);
DFFARX1 I_71857 (I1225157,I3563,I1225123,I1225106,);
DFFARX1 I_71858 (I1367228,I3563,I1225123,I1225197,);
not I_71859 (I1225205,I1367243);
not I_71860 (I1225222,I1367231);
nand I_71861 (I1225239,I1225222,I1225205);
nor I_71862 (I1225094,I1225197,I1225239);
DFFARX1 I_71863 (I1225239,I3563,I1225123,I1225279,);
not I_71864 (I1225115,I1225279);
not I_71865 (I1225301,I1367240);
nand I_71866 (I1225318,I1225222,I1225301);
DFFARX1 I_71867 (I1225318,I3563,I1225123,I1225344,);
not I_71868 (I1225352,I1225344);
not I_71869 (I1225369,I1367249);
nand I_71870 (I1225386,I1225369,I1367228);
and I_71871 (I1225403,I1225205,I1225386);
nor I_71872 (I1225420,I1225318,I1225403);
DFFARX1 I_71873 (I1225420,I3563,I1225123,I1225091,);
DFFARX1 I_71874 (I1225403,I3563,I1225123,I1225112,);
nor I_71875 (I1225465,I1367249,I1367252);
nor I_71876 (I1225103,I1225318,I1225465);
or I_71877 (I1225496,I1367249,I1367252);
nor I_71878 (I1225513,I1367246,I1367234);
DFFARX1 I_71879 (I1225513,I3563,I1225123,I1225539,);
not I_71880 (I1225547,I1225539);
nor I_71881 (I1225109,I1225547,I1225352);
nand I_71882 (I1225578,I1225547,I1225197);
not I_71883 (I1225595,I1367246);
nand I_71884 (I1225612,I1225595,I1225301);
nand I_71885 (I1225629,I1225547,I1225612);
nand I_71886 (I1225100,I1225629,I1225578);
nand I_71887 (I1225097,I1225612,I1225496);
not I_71888 (I1225701,I3570);
DFFARX1 I_71889 (I657850,I3563,I1225701,I1225727,);
and I_71890 (I1225735,I1225727,I657838);
DFFARX1 I_71891 (I1225735,I3563,I1225701,I1225684,);
DFFARX1 I_71892 (I657853,I3563,I1225701,I1225775,);
not I_71893 (I1225783,I657844);
not I_71894 (I1225800,I657835);
nand I_71895 (I1225817,I1225800,I1225783);
nor I_71896 (I1225672,I1225775,I1225817);
DFFARX1 I_71897 (I1225817,I3563,I1225701,I1225857,);
not I_71898 (I1225693,I1225857);
not I_71899 (I1225879,I657841);
nand I_71900 (I1225896,I1225800,I1225879);
DFFARX1 I_71901 (I1225896,I3563,I1225701,I1225922,);
not I_71902 (I1225930,I1225922);
not I_71903 (I1225947,I657856);
nand I_71904 (I1225964,I1225947,I657859);
and I_71905 (I1225981,I1225783,I1225964);
nor I_71906 (I1225998,I1225896,I1225981);
DFFARX1 I_71907 (I1225998,I3563,I1225701,I1225669,);
DFFARX1 I_71908 (I1225981,I3563,I1225701,I1225690,);
nor I_71909 (I1226043,I657856,I657835);
nor I_71910 (I1225681,I1225896,I1226043);
or I_71911 (I1226074,I657856,I657835);
nor I_71912 (I1226091,I657847,I657838);
DFFARX1 I_71913 (I1226091,I3563,I1225701,I1226117,);
not I_71914 (I1226125,I1226117);
nor I_71915 (I1225687,I1226125,I1225930);
nand I_71916 (I1226156,I1226125,I1225775);
not I_71917 (I1226173,I657847);
nand I_71918 (I1226190,I1226173,I1225879);
nand I_71919 (I1226207,I1226125,I1226190);
nand I_71920 (I1225678,I1226207,I1226156);
nand I_71921 (I1225675,I1226190,I1226074);
not I_71922 (I1226279,I3570);
DFFARX1 I_71923 (I1246974,I3563,I1226279,I1226305,);
and I_71924 (I1226313,I1226305,I1246968);
DFFARX1 I_71925 (I1226313,I3563,I1226279,I1226262,);
DFFARX1 I_71926 (I1246953,I3563,I1226279,I1226353,);
not I_71927 (I1226361,I1246959);
not I_71928 (I1226378,I1246971);
nand I_71929 (I1226395,I1226378,I1226361);
nor I_71930 (I1226250,I1226353,I1226395);
DFFARX1 I_71931 (I1226395,I3563,I1226279,I1226435,);
not I_71932 (I1226271,I1226435);
not I_71933 (I1226457,I1246953);
nand I_71934 (I1226474,I1226378,I1226457);
DFFARX1 I_71935 (I1226474,I3563,I1226279,I1226500,);
not I_71936 (I1226508,I1226500);
not I_71937 (I1226525,I1246977);
nand I_71938 (I1226542,I1226525,I1246965);
and I_71939 (I1226559,I1226361,I1226542);
nor I_71940 (I1226576,I1226474,I1226559);
DFFARX1 I_71941 (I1226576,I3563,I1226279,I1226247,);
DFFARX1 I_71942 (I1226559,I3563,I1226279,I1226268,);
nor I_71943 (I1226621,I1246977,I1246956);
nor I_71944 (I1226259,I1226474,I1226621);
or I_71945 (I1226652,I1246977,I1246956);
nor I_71946 (I1226669,I1246962,I1246956);
DFFARX1 I_71947 (I1226669,I3563,I1226279,I1226695,);
not I_71948 (I1226703,I1226695);
nor I_71949 (I1226265,I1226703,I1226508);
nand I_71950 (I1226734,I1226703,I1226353);
not I_71951 (I1226751,I1246962);
nand I_71952 (I1226768,I1226751,I1226457);
nand I_71953 (I1226785,I1226703,I1226768);
nand I_71954 (I1226256,I1226785,I1226734);
nand I_71955 (I1226253,I1226768,I1226652);
not I_71956 (I1226857,I3570);
DFFARX1 I_71957 (I23973,I3563,I1226857,I1226883,);
and I_71958 (I1226891,I1226883,I23976);
DFFARX1 I_71959 (I1226891,I3563,I1226857,I1226840,);
DFFARX1 I_71960 (I23976,I3563,I1226857,I1226931,);
not I_71961 (I1226939,I23979);
not I_71962 (I1226956,I23994);
nand I_71963 (I1226973,I1226956,I1226939);
nor I_71964 (I1226828,I1226931,I1226973);
DFFARX1 I_71965 (I1226973,I3563,I1226857,I1227013,);
not I_71966 (I1226849,I1227013);
not I_71967 (I1227035,I23988);
nand I_71968 (I1227052,I1226956,I1227035);
DFFARX1 I_71969 (I1227052,I3563,I1226857,I1227078,);
not I_71970 (I1227086,I1227078);
not I_71971 (I1227103,I23991);
nand I_71972 (I1227120,I1227103,I23973);
and I_71973 (I1227137,I1226939,I1227120);
nor I_71974 (I1227154,I1227052,I1227137);
DFFARX1 I_71975 (I1227154,I3563,I1226857,I1226825,);
DFFARX1 I_71976 (I1227137,I3563,I1226857,I1226846,);
nor I_71977 (I1227199,I23991,I23985);
nor I_71978 (I1226837,I1227052,I1227199);
or I_71979 (I1227230,I23991,I23985);
nor I_71980 (I1227247,I23982,I23997);
DFFARX1 I_71981 (I1227247,I3563,I1226857,I1227273,);
not I_71982 (I1227281,I1227273);
nor I_71983 (I1226843,I1227281,I1227086);
nand I_71984 (I1227312,I1227281,I1226931);
not I_71985 (I1227329,I23982);
nand I_71986 (I1227346,I1227329,I1227035);
nand I_71987 (I1227363,I1227281,I1227346);
nand I_71988 (I1226834,I1227363,I1227312);
nand I_71989 (I1226831,I1227346,I1227230);
not I_71990 (I1227435,I3570);
DFFARX1 I_71991 (I512706,I3563,I1227435,I1227461,);
and I_71992 (I1227469,I1227461,I512721);
DFFARX1 I_71993 (I1227469,I3563,I1227435,I1227418,);
DFFARX1 I_71994 (I512724,I3563,I1227435,I1227509,);
not I_71995 (I1227517,I512718);
not I_71996 (I1227534,I512733);
nand I_71997 (I1227551,I1227534,I1227517);
nor I_71998 (I1227406,I1227509,I1227551);
DFFARX1 I_71999 (I1227551,I3563,I1227435,I1227591,);
not I_72000 (I1227427,I1227591);
not I_72001 (I1227613,I512709);
nand I_72002 (I1227630,I1227534,I1227613);
DFFARX1 I_72003 (I1227630,I3563,I1227435,I1227656,);
not I_72004 (I1227664,I1227656);
not I_72005 (I1227681,I512712);
nand I_72006 (I1227698,I1227681,I512706);
and I_72007 (I1227715,I1227517,I1227698);
nor I_72008 (I1227732,I1227630,I1227715);
DFFARX1 I_72009 (I1227732,I3563,I1227435,I1227403,);
DFFARX1 I_72010 (I1227715,I3563,I1227435,I1227424,);
nor I_72011 (I1227777,I512712,I512715);
nor I_72012 (I1227415,I1227630,I1227777);
or I_72013 (I1227808,I512712,I512715);
nor I_72014 (I1227825,I512730,I512727);
DFFARX1 I_72015 (I1227825,I3563,I1227435,I1227851,);
not I_72016 (I1227859,I1227851);
nor I_72017 (I1227421,I1227859,I1227664);
nand I_72018 (I1227890,I1227859,I1227509);
not I_72019 (I1227907,I512730);
nand I_72020 (I1227924,I1227907,I1227613);
nand I_72021 (I1227941,I1227859,I1227924);
nand I_72022 (I1227412,I1227941,I1227890);
nand I_72023 (I1227409,I1227924,I1227808);
not I_72024 (I1228013,I3570);
DFFARX1 I_72025 (I202388,I3563,I1228013,I1228039,);
and I_72026 (I1228047,I1228039,I202391);
DFFARX1 I_72027 (I1228047,I3563,I1228013,I1227996,);
DFFARX1 I_72028 (I202391,I3563,I1228013,I1228087,);
not I_72029 (I1228095,I202406);
not I_72030 (I1228112,I202412);
nand I_72031 (I1228129,I1228112,I1228095);
nor I_72032 (I1227984,I1228087,I1228129);
DFFARX1 I_72033 (I1228129,I3563,I1228013,I1228169,);
not I_72034 (I1228005,I1228169);
not I_72035 (I1228191,I202400);
nand I_72036 (I1228208,I1228112,I1228191);
DFFARX1 I_72037 (I1228208,I3563,I1228013,I1228234,);
not I_72038 (I1228242,I1228234);
not I_72039 (I1228259,I202397);
nand I_72040 (I1228276,I1228259,I202394);
and I_72041 (I1228293,I1228095,I1228276);
nor I_72042 (I1228310,I1228208,I1228293);
DFFARX1 I_72043 (I1228310,I3563,I1228013,I1227981,);
DFFARX1 I_72044 (I1228293,I3563,I1228013,I1228002,);
nor I_72045 (I1228355,I202397,I202388);
nor I_72046 (I1227993,I1228208,I1228355);
or I_72047 (I1228386,I202397,I202388);
nor I_72048 (I1228403,I202403,I202409);
DFFARX1 I_72049 (I1228403,I3563,I1228013,I1228429,);
not I_72050 (I1228437,I1228429);
nor I_72051 (I1227999,I1228437,I1228242);
nand I_72052 (I1228468,I1228437,I1228087);
not I_72053 (I1228485,I202403);
nand I_72054 (I1228502,I1228485,I1228191);
nand I_72055 (I1228519,I1228437,I1228502);
nand I_72056 (I1227990,I1228519,I1228468);
nand I_72057 (I1227987,I1228502,I1228386);
not I_72058 (I1228591,I3570);
DFFARX1 I_72059 (I1256222,I3563,I1228591,I1228617,);
and I_72060 (I1228625,I1228617,I1256216);
DFFARX1 I_72061 (I1228625,I3563,I1228591,I1228574,);
DFFARX1 I_72062 (I1256201,I3563,I1228591,I1228665,);
not I_72063 (I1228673,I1256207);
not I_72064 (I1228690,I1256219);
nand I_72065 (I1228707,I1228690,I1228673);
nor I_72066 (I1228562,I1228665,I1228707);
DFFARX1 I_72067 (I1228707,I3563,I1228591,I1228747,);
not I_72068 (I1228583,I1228747);
not I_72069 (I1228769,I1256201);
nand I_72070 (I1228786,I1228690,I1228769);
DFFARX1 I_72071 (I1228786,I3563,I1228591,I1228812,);
not I_72072 (I1228820,I1228812);
not I_72073 (I1228837,I1256225);
nand I_72074 (I1228854,I1228837,I1256213);
and I_72075 (I1228871,I1228673,I1228854);
nor I_72076 (I1228888,I1228786,I1228871);
DFFARX1 I_72077 (I1228888,I3563,I1228591,I1228559,);
DFFARX1 I_72078 (I1228871,I3563,I1228591,I1228580,);
nor I_72079 (I1228933,I1256225,I1256204);
nor I_72080 (I1228571,I1228786,I1228933);
or I_72081 (I1228964,I1256225,I1256204);
nor I_72082 (I1228981,I1256210,I1256204);
DFFARX1 I_72083 (I1228981,I3563,I1228591,I1229007,);
not I_72084 (I1229015,I1229007);
nor I_72085 (I1228577,I1229015,I1228820);
nand I_72086 (I1229046,I1229015,I1228665);
not I_72087 (I1229063,I1256210);
nand I_72088 (I1229080,I1229063,I1228769);
nand I_72089 (I1229097,I1229015,I1229080);
nand I_72090 (I1228568,I1229097,I1229046);
nand I_72091 (I1228565,I1229080,I1228964);
not I_72092 (I1229169,I3570);
DFFARX1 I_72093 (I874826,I3563,I1229169,I1229195,);
and I_72094 (I1229203,I1229195,I874832);
DFFARX1 I_72095 (I1229203,I3563,I1229169,I1229152,);
DFFARX1 I_72096 (I874838,I3563,I1229169,I1229243,);
not I_72097 (I1229251,I874823);
not I_72098 (I1229268,I874823);
nand I_72099 (I1229285,I1229268,I1229251);
nor I_72100 (I1229140,I1229243,I1229285);
DFFARX1 I_72101 (I1229285,I3563,I1229169,I1229325,);
not I_72102 (I1229161,I1229325);
not I_72103 (I1229347,I874841);
nand I_72104 (I1229364,I1229268,I1229347);
DFFARX1 I_72105 (I1229364,I3563,I1229169,I1229390,);
not I_72106 (I1229398,I1229390);
not I_72107 (I1229415,I874835);
nand I_72108 (I1229432,I1229415,I874826);
and I_72109 (I1229449,I1229251,I1229432);
nor I_72110 (I1229466,I1229364,I1229449);
DFFARX1 I_72111 (I1229466,I3563,I1229169,I1229137,);
DFFARX1 I_72112 (I1229449,I3563,I1229169,I1229158,);
nor I_72113 (I1229511,I874835,I874844);
nor I_72114 (I1229149,I1229364,I1229511);
or I_72115 (I1229542,I874835,I874844);
nor I_72116 (I1229559,I874829,I874829);
DFFARX1 I_72117 (I1229559,I3563,I1229169,I1229585,);
not I_72118 (I1229593,I1229585);
nor I_72119 (I1229155,I1229593,I1229398);
nand I_72120 (I1229624,I1229593,I1229243);
not I_72121 (I1229641,I874829);
nand I_72122 (I1229658,I1229641,I1229347);
nand I_72123 (I1229675,I1229593,I1229658);
nand I_72124 (I1229146,I1229675,I1229624);
nand I_72125 (I1229143,I1229658,I1229542);
not I_72126 (I1229747,I3570);
DFFARX1 I_72127 (I261888,I3563,I1229747,I1229773,);
and I_72128 (I1229781,I1229773,I261891);
DFFARX1 I_72129 (I1229781,I3563,I1229747,I1229730,);
DFFARX1 I_72130 (I261891,I3563,I1229747,I1229821,);
not I_72131 (I1229829,I261906);
not I_72132 (I1229846,I261912);
nand I_72133 (I1229863,I1229846,I1229829);
nor I_72134 (I1229718,I1229821,I1229863);
DFFARX1 I_72135 (I1229863,I3563,I1229747,I1229903,);
not I_72136 (I1229739,I1229903);
not I_72137 (I1229925,I261900);
nand I_72138 (I1229942,I1229846,I1229925);
DFFARX1 I_72139 (I1229942,I3563,I1229747,I1229968,);
not I_72140 (I1229976,I1229968);
not I_72141 (I1229993,I261897);
nand I_72142 (I1230010,I1229993,I261894);
and I_72143 (I1230027,I1229829,I1230010);
nor I_72144 (I1230044,I1229942,I1230027);
DFFARX1 I_72145 (I1230044,I3563,I1229747,I1229715,);
DFFARX1 I_72146 (I1230027,I3563,I1229747,I1229736,);
nor I_72147 (I1230089,I261897,I261888);
nor I_72148 (I1229727,I1229942,I1230089);
or I_72149 (I1230120,I261897,I261888);
nor I_72150 (I1230137,I261903,I261909);
DFFARX1 I_72151 (I1230137,I3563,I1229747,I1230163,);
not I_72152 (I1230171,I1230163);
nor I_72153 (I1229733,I1230171,I1229976);
nand I_72154 (I1230202,I1230171,I1229821);
not I_72155 (I1230219,I261903);
nand I_72156 (I1230236,I1230219,I1229925);
nand I_72157 (I1230253,I1230171,I1230236);
nand I_72158 (I1229724,I1230253,I1230202);
nand I_72159 (I1229721,I1230236,I1230120);
not I_72160 (I1230325,I3570);
DFFARX1 I_72161 (I1287230,I3563,I1230325,I1230351,);
and I_72162 (I1230359,I1230351,I1287224);
DFFARX1 I_72163 (I1230359,I3563,I1230325,I1230308,);
DFFARX1 I_72164 (I1287209,I3563,I1230325,I1230399,);
not I_72165 (I1230407,I1287215);
not I_72166 (I1230424,I1287227);
nand I_72167 (I1230441,I1230424,I1230407);
nor I_72168 (I1230296,I1230399,I1230441);
DFFARX1 I_72169 (I1230441,I3563,I1230325,I1230481,);
not I_72170 (I1230317,I1230481);
not I_72171 (I1230503,I1287209);
nand I_72172 (I1230520,I1230424,I1230503);
DFFARX1 I_72173 (I1230520,I3563,I1230325,I1230546,);
not I_72174 (I1230554,I1230546);
not I_72175 (I1230571,I1287233);
nand I_72176 (I1230588,I1230571,I1287221);
and I_72177 (I1230605,I1230407,I1230588);
nor I_72178 (I1230622,I1230520,I1230605);
DFFARX1 I_72179 (I1230622,I3563,I1230325,I1230293,);
DFFARX1 I_72180 (I1230605,I3563,I1230325,I1230314,);
nor I_72181 (I1230667,I1287233,I1287212);
nor I_72182 (I1230305,I1230520,I1230667);
or I_72183 (I1230698,I1287233,I1287212);
nor I_72184 (I1230715,I1287218,I1287212);
DFFARX1 I_72185 (I1230715,I3563,I1230325,I1230741,);
not I_72186 (I1230749,I1230741);
nor I_72187 (I1230311,I1230749,I1230554);
nand I_72188 (I1230780,I1230749,I1230399);
not I_72189 (I1230797,I1287218);
nand I_72190 (I1230814,I1230797,I1230503);
nand I_72191 (I1230831,I1230749,I1230814);
nand I_72192 (I1230302,I1230831,I1230780);
nand I_72193 (I1230299,I1230814,I1230698);
not I_72194 (I1230903,I3570);
DFFARX1 I_72195 (I90926,I3563,I1230903,I1230929,);
and I_72196 (I1230937,I1230929,I90902);
DFFARX1 I_72197 (I1230937,I3563,I1230903,I1230886,);
DFFARX1 I_72198 (I90920,I3563,I1230903,I1230977,);
not I_72199 (I1230985,I90908);
not I_72200 (I1231002,I90905);
nand I_72201 (I1231019,I1231002,I1230985);
nor I_72202 (I1230874,I1230977,I1231019);
DFFARX1 I_72203 (I1231019,I3563,I1230903,I1231059,);
not I_72204 (I1230895,I1231059);
not I_72205 (I1231081,I90914);
nand I_72206 (I1231098,I1231002,I1231081);
DFFARX1 I_72207 (I1231098,I3563,I1230903,I1231124,);
not I_72208 (I1231132,I1231124);
not I_72209 (I1231149,I90905);
nand I_72210 (I1231166,I1231149,I90923);
and I_72211 (I1231183,I1230985,I1231166);
nor I_72212 (I1231200,I1231098,I1231183);
DFFARX1 I_72213 (I1231200,I3563,I1230903,I1230871,);
DFFARX1 I_72214 (I1231183,I3563,I1230903,I1230892,);
nor I_72215 (I1231245,I90905,I90917);
nor I_72216 (I1230883,I1231098,I1231245);
or I_72217 (I1231276,I90905,I90917);
nor I_72218 (I1231293,I90911,I90902);
DFFARX1 I_72219 (I1231293,I3563,I1230903,I1231319,);
not I_72220 (I1231327,I1231319);
nor I_72221 (I1230889,I1231327,I1231132);
nand I_72222 (I1231358,I1231327,I1230977);
not I_72223 (I1231375,I90911);
nand I_72224 (I1231392,I1231375,I1231081);
nand I_72225 (I1231409,I1231327,I1231392);
nand I_72226 (I1230880,I1231409,I1231358);
nand I_72227 (I1230877,I1231392,I1231276);
not I_72228 (I1231481,I3570);
DFFARX1 I_72229 (I1062931,I3563,I1231481,I1231507,);
and I_72230 (I1231515,I1231507,I1062928);
DFFARX1 I_72231 (I1231515,I3563,I1231481,I1231464,);
DFFARX1 I_72232 (I1062934,I3563,I1231481,I1231555,);
not I_72233 (I1231563,I1062937);
not I_72234 (I1231580,I1062931);
nand I_72235 (I1231597,I1231580,I1231563);
nor I_72236 (I1231452,I1231555,I1231597);
DFFARX1 I_72237 (I1231597,I3563,I1231481,I1231637,);
not I_72238 (I1231473,I1231637);
not I_72239 (I1231659,I1062946);
nand I_72240 (I1231676,I1231580,I1231659);
DFFARX1 I_72241 (I1231676,I3563,I1231481,I1231702,);
not I_72242 (I1231710,I1231702);
not I_72243 (I1231727,I1062943);
nand I_72244 (I1231744,I1231727,I1062949);
and I_72245 (I1231761,I1231563,I1231744);
nor I_72246 (I1231778,I1231676,I1231761);
DFFARX1 I_72247 (I1231778,I3563,I1231481,I1231449,);
DFFARX1 I_72248 (I1231761,I3563,I1231481,I1231470,);
nor I_72249 (I1231823,I1062943,I1062928);
nor I_72250 (I1231461,I1231676,I1231823);
or I_72251 (I1231854,I1062943,I1062928);
nor I_72252 (I1231871,I1062940,I1062934);
DFFARX1 I_72253 (I1231871,I3563,I1231481,I1231897,);
not I_72254 (I1231905,I1231897);
nor I_72255 (I1231467,I1231905,I1231710);
nand I_72256 (I1231936,I1231905,I1231555);
not I_72257 (I1231953,I1062940);
nand I_72258 (I1231970,I1231953,I1231659);
nand I_72259 (I1231987,I1231905,I1231970);
nand I_72260 (I1231458,I1231987,I1231936);
nand I_72261 (I1231455,I1231970,I1231854);
not I_72262 (I1232059,I3570);
DFFARX1 I_72263 (I628372,I3563,I1232059,I1232085,);
and I_72264 (I1232093,I1232085,I628360);
DFFARX1 I_72265 (I1232093,I3563,I1232059,I1232042,);
DFFARX1 I_72266 (I628375,I3563,I1232059,I1232133,);
not I_72267 (I1232141,I628366);
not I_72268 (I1232158,I628357);
nand I_72269 (I1232175,I1232158,I1232141);
nor I_72270 (I1232030,I1232133,I1232175);
DFFARX1 I_72271 (I1232175,I3563,I1232059,I1232215,);
not I_72272 (I1232051,I1232215);
not I_72273 (I1232237,I628363);
nand I_72274 (I1232254,I1232158,I1232237);
DFFARX1 I_72275 (I1232254,I3563,I1232059,I1232280,);
not I_72276 (I1232288,I1232280);
not I_72277 (I1232305,I628378);
nand I_72278 (I1232322,I1232305,I628381);
and I_72279 (I1232339,I1232141,I1232322);
nor I_72280 (I1232356,I1232254,I1232339);
DFFARX1 I_72281 (I1232356,I3563,I1232059,I1232027,);
DFFARX1 I_72282 (I1232339,I3563,I1232059,I1232048,);
nor I_72283 (I1232401,I628378,I628357);
nor I_72284 (I1232039,I1232254,I1232401);
or I_72285 (I1232432,I628378,I628357);
nor I_72286 (I1232449,I628369,I628360);
DFFARX1 I_72287 (I1232449,I3563,I1232059,I1232475,);
not I_72288 (I1232483,I1232475);
nor I_72289 (I1232045,I1232483,I1232288);
nand I_72290 (I1232514,I1232483,I1232133);
not I_72291 (I1232531,I628369);
nand I_72292 (I1232548,I1232531,I1232237);
nand I_72293 (I1232565,I1232483,I1232548);
nand I_72294 (I1232036,I1232565,I1232514);
nand I_72295 (I1232033,I1232548,I1232432);
not I_72296 (I1232637,I3570);
DFFARX1 I_72297 (I117803,I3563,I1232637,I1232663,);
and I_72298 (I1232671,I1232663,I117779);
DFFARX1 I_72299 (I1232671,I3563,I1232637,I1232620,);
DFFARX1 I_72300 (I117797,I3563,I1232637,I1232711,);
not I_72301 (I1232719,I117785);
not I_72302 (I1232736,I117782);
nand I_72303 (I1232753,I1232736,I1232719);
nor I_72304 (I1232608,I1232711,I1232753);
DFFARX1 I_72305 (I1232753,I3563,I1232637,I1232793,);
not I_72306 (I1232629,I1232793);
not I_72307 (I1232815,I117791);
nand I_72308 (I1232832,I1232736,I1232815);
DFFARX1 I_72309 (I1232832,I3563,I1232637,I1232858,);
not I_72310 (I1232866,I1232858);
not I_72311 (I1232883,I117782);
nand I_72312 (I1232900,I1232883,I117800);
and I_72313 (I1232917,I1232719,I1232900);
nor I_72314 (I1232934,I1232832,I1232917);
DFFARX1 I_72315 (I1232934,I3563,I1232637,I1232605,);
DFFARX1 I_72316 (I1232917,I3563,I1232637,I1232626,);
nor I_72317 (I1232979,I117782,I117794);
nor I_72318 (I1232617,I1232832,I1232979);
or I_72319 (I1233010,I117782,I117794);
nor I_72320 (I1233027,I117788,I117779);
DFFARX1 I_72321 (I1233027,I3563,I1232637,I1233053,);
not I_72322 (I1233061,I1233053);
nor I_72323 (I1232623,I1233061,I1232866);
nand I_72324 (I1233092,I1233061,I1232711);
not I_72325 (I1233109,I117788);
nand I_72326 (I1233126,I1233109,I1232815);
nand I_72327 (I1233143,I1233061,I1233126);
nand I_72328 (I1232614,I1233143,I1233092);
nand I_72329 (I1232611,I1233126,I1233010);
not I_72330 (I1233215,I3570);
DFFARX1 I_72331 (I728366,I3563,I1233215,I1233241,);
and I_72332 (I1233249,I1233241,I728354);
DFFARX1 I_72333 (I1233249,I3563,I1233215,I1233198,);
DFFARX1 I_72334 (I728357,I3563,I1233215,I1233289,);
not I_72335 (I1233297,I728351);
not I_72336 (I1233314,I728375);
nand I_72337 (I1233331,I1233314,I1233297);
nor I_72338 (I1233186,I1233289,I1233331);
DFFARX1 I_72339 (I1233331,I3563,I1233215,I1233371,);
not I_72340 (I1233207,I1233371);
not I_72341 (I1233393,I728363);
nand I_72342 (I1233410,I1233314,I1233393);
DFFARX1 I_72343 (I1233410,I3563,I1233215,I1233436,);
not I_72344 (I1233444,I1233436);
not I_72345 (I1233461,I728372);
nand I_72346 (I1233478,I1233461,I728369);
and I_72347 (I1233495,I1233297,I1233478);
nor I_72348 (I1233512,I1233410,I1233495);
DFFARX1 I_72349 (I1233512,I3563,I1233215,I1233183,);
DFFARX1 I_72350 (I1233495,I3563,I1233215,I1233204,);
nor I_72351 (I1233557,I728372,I728360);
nor I_72352 (I1233195,I1233410,I1233557);
or I_72353 (I1233588,I728372,I728360);
nor I_72354 (I1233605,I728351,I728354);
DFFARX1 I_72355 (I1233605,I3563,I1233215,I1233631,);
not I_72356 (I1233639,I1233631);
nor I_72357 (I1233201,I1233639,I1233444);
nand I_72358 (I1233670,I1233639,I1233289);
not I_72359 (I1233687,I728351);
nand I_72360 (I1233704,I1233687,I1233393);
nand I_72361 (I1233721,I1233639,I1233704);
nand I_72362 (I1233192,I1233721,I1233670);
nand I_72363 (I1233189,I1233704,I1233588);
not I_72364 (I1233793,I3570);
DFFARX1 I_72365 (I368131,I3563,I1233793,I1233819,);
and I_72366 (I1233827,I1233819,I368116);
DFFARX1 I_72367 (I1233827,I3563,I1233793,I1233776,);
DFFARX1 I_72368 (I368122,I3563,I1233793,I1233867,);
not I_72369 (I1233875,I368104);
not I_72370 (I1233892,I368125);
nand I_72371 (I1233909,I1233892,I1233875);
nor I_72372 (I1233764,I1233867,I1233909);
DFFARX1 I_72373 (I1233909,I3563,I1233793,I1233949,);
not I_72374 (I1233785,I1233949);
not I_72375 (I1233971,I368128);
nand I_72376 (I1233988,I1233892,I1233971);
DFFARX1 I_72377 (I1233988,I3563,I1233793,I1234014,);
not I_72378 (I1234022,I1234014);
not I_72379 (I1234039,I368119);
nand I_72380 (I1234056,I1234039,I368107);
and I_72381 (I1234073,I1233875,I1234056);
nor I_72382 (I1234090,I1233988,I1234073);
DFFARX1 I_72383 (I1234090,I3563,I1233793,I1233761,);
DFFARX1 I_72384 (I1234073,I3563,I1233793,I1233782,);
nor I_72385 (I1234135,I368119,I368113);
nor I_72386 (I1233773,I1233988,I1234135);
or I_72387 (I1234166,I368119,I368113);
nor I_72388 (I1234183,I368110,I368104);
DFFARX1 I_72389 (I1234183,I3563,I1233793,I1234209,);
not I_72390 (I1234217,I1234209);
nor I_72391 (I1233779,I1234217,I1234022);
nand I_72392 (I1234248,I1234217,I1233867);
not I_72393 (I1234265,I368110);
nand I_72394 (I1234282,I1234265,I1233971);
nand I_72395 (I1234299,I1234217,I1234282);
nand I_72396 (I1233770,I1234299,I1234248);
nand I_72397 (I1233767,I1234282,I1234166);
not I_72398 (I1234371,I3570);
DFFARX1 I_72399 (I567959,I3563,I1234371,I1234397,);
and I_72400 (I1234405,I1234397,I567974);
DFFARX1 I_72401 (I1234405,I3563,I1234371,I1234354,);
DFFARX1 I_72402 (I567965,I3563,I1234371,I1234445,);
not I_72403 (I1234453,I567959);
not I_72404 (I1234470,I567977);
nand I_72405 (I1234487,I1234470,I1234453);
nor I_72406 (I1234342,I1234445,I1234487);
DFFARX1 I_72407 (I1234487,I3563,I1234371,I1234527,);
not I_72408 (I1234363,I1234527);
not I_72409 (I1234549,I567968);
nand I_72410 (I1234566,I1234470,I1234549);
DFFARX1 I_72411 (I1234566,I3563,I1234371,I1234592,);
not I_72412 (I1234600,I1234592);
not I_72413 (I1234617,I567980);
nand I_72414 (I1234634,I1234617,I567956);
and I_72415 (I1234651,I1234453,I1234634);
nor I_72416 (I1234668,I1234566,I1234651);
DFFARX1 I_72417 (I1234668,I3563,I1234371,I1234339,);
DFFARX1 I_72418 (I1234651,I3563,I1234371,I1234360,);
nor I_72419 (I1234713,I567980,I567956);
nor I_72420 (I1234351,I1234566,I1234713);
or I_72421 (I1234744,I567980,I567956);
nor I_72422 (I1234761,I567962,I567971);
DFFARX1 I_72423 (I1234761,I3563,I1234371,I1234787,);
not I_72424 (I1234795,I1234787);
nor I_72425 (I1234357,I1234795,I1234600);
nand I_72426 (I1234826,I1234795,I1234445);
not I_72427 (I1234843,I567962);
nand I_72428 (I1234860,I1234843,I1234549);
nand I_72429 (I1234877,I1234795,I1234860);
nand I_72430 (I1234348,I1234877,I1234826);
nand I_72431 (I1234345,I1234860,I1234744);
not I_72432 (I1234949,I3570);
DFFARX1 I_72433 (I19230,I3563,I1234949,I1234975,);
and I_72434 (I1234983,I1234975,I19233);
DFFARX1 I_72435 (I1234983,I3563,I1234949,I1234932,);
DFFARX1 I_72436 (I19233,I3563,I1234949,I1235023,);
not I_72437 (I1235031,I19236);
not I_72438 (I1235048,I19251);
nand I_72439 (I1235065,I1235048,I1235031);
nor I_72440 (I1234920,I1235023,I1235065);
DFFARX1 I_72441 (I1235065,I3563,I1234949,I1235105,);
not I_72442 (I1234941,I1235105);
not I_72443 (I1235127,I19245);
nand I_72444 (I1235144,I1235048,I1235127);
DFFARX1 I_72445 (I1235144,I3563,I1234949,I1235170,);
not I_72446 (I1235178,I1235170);
not I_72447 (I1235195,I19248);
nand I_72448 (I1235212,I1235195,I19230);
and I_72449 (I1235229,I1235031,I1235212);
nor I_72450 (I1235246,I1235144,I1235229);
DFFARX1 I_72451 (I1235246,I3563,I1234949,I1234917,);
DFFARX1 I_72452 (I1235229,I3563,I1234949,I1234938,);
nor I_72453 (I1235291,I19248,I19242);
nor I_72454 (I1234929,I1235144,I1235291);
or I_72455 (I1235322,I19248,I19242);
nor I_72456 (I1235339,I19239,I19254);
DFFARX1 I_72457 (I1235339,I3563,I1234949,I1235365,);
not I_72458 (I1235373,I1235365);
nor I_72459 (I1234935,I1235373,I1235178);
nand I_72460 (I1235404,I1235373,I1235023);
not I_72461 (I1235421,I19239);
nand I_72462 (I1235438,I1235421,I1235127);
nand I_72463 (I1235455,I1235373,I1235438);
nand I_72464 (I1234926,I1235455,I1235404);
nand I_72465 (I1234923,I1235438,I1235322);
not I_72466 (I1235527,I3570);
DFFARX1 I_72467 (I700044,I3563,I1235527,I1235553,);
and I_72468 (I1235561,I1235553,I700032);
DFFARX1 I_72469 (I1235561,I3563,I1235527,I1235510,);
DFFARX1 I_72470 (I700035,I3563,I1235527,I1235601,);
not I_72471 (I1235609,I700029);
not I_72472 (I1235626,I700053);
nand I_72473 (I1235643,I1235626,I1235609);
nor I_72474 (I1235498,I1235601,I1235643);
DFFARX1 I_72475 (I1235643,I3563,I1235527,I1235683,);
not I_72476 (I1235519,I1235683);
not I_72477 (I1235705,I700041);
nand I_72478 (I1235722,I1235626,I1235705);
DFFARX1 I_72479 (I1235722,I3563,I1235527,I1235748,);
not I_72480 (I1235756,I1235748);
not I_72481 (I1235773,I700050);
nand I_72482 (I1235790,I1235773,I700047);
and I_72483 (I1235807,I1235609,I1235790);
nor I_72484 (I1235824,I1235722,I1235807);
DFFARX1 I_72485 (I1235824,I3563,I1235527,I1235495,);
DFFARX1 I_72486 (I1235807,I3563,I1235527,I1235516,);
nor I_72487 (I1235869,I700050,I700038);
nor I_72488 (I1235507,I1235722,I1235869);
or I_72489 (I1235900,I700050,I700038);
nor I_72490 (I1235917,I700029,I700032);
DFFARX1 I_72491 (I1235917,I3563,I1235527,I1235943,);
not I_72492 (I1235951,I1235943);
nor I_72493 (I1235513,I1235951,I1235756);
nand I_72494 (I1235982,I1235951,I1235601);
not I_72495 (I1235999,I700029);
nand I_72496 (I1236016,I1235999,I1235705);
nand I_72497 (I1236033,I1235951,I1236016);
nand I_72498 (I1235504,I1236033,I1235982);
nand I_72499 (I1235501,I1236016,I1235900);
not I_72500 (I1236105,I3570);
DFFARX1 I_72501 (I179778,I3563,I1236105,I1236131,);
and I_72502 (I1236139,I1236131,I179781);
DFFARX1 I_72503 (I1236139,I3563,I1236105,I1236088,);
DFFARX1 I_72504 (I179781,I3563,I1236105,I1236179,);
not I_72505 (I1236187,I179796);
not I_72506 (I1236204,I179802);
nand I_72507 (I1236221,I1236204,I1236187);
nor I_72508 (I1236076,I1236179,I1236221);
DFFARX1 I_72509 (I1236221,I3563,I1236105,I1236261,);
not I_72510 (I1236097,I1236261);
not I_72511 (I1236283,I179790);
nand I_72512 (I1236300,I1236204,I1236283);
DFFARX1 I_72513 (I1236300,I3563,I1236105,I1236326,);
not I_72514 (I1236334,I1236326);
not I_72515 (I1236351,I179787);
nand I_72516 (I1236368,I1236351,I179784);
and I_72517 (I1236385,I1236187,I1236368);
nor I_72518 (I1236402,I1236300,I1236385);
DFFARX1 I_72519 (I1236402,I3563,I1236105,I1236073,);
DFFARX1 I_72520 (I1236385,I3563,I1236105,I1236094,);
nor I_72521 (I1236447,I179787,I179778);
nor I_72522 (I1236085,I1236300,I1236447);
or I_72523 (I1236478,I179787,I179778);
nor I_72524 (I1236495,I179793,I179799);
DFFARX1 I_72525 (I1236495,I3563,I1236105,I1236521,);
not I_72526 (I1236529,I1236521);
nor I_72527 (I1236091,I1236529,I1236334);
nand I_72528 (I1236560,I1236529,I1236179);
not I_72529 (I1236577,I179793);
nand I_72530 (I1236594,I1236577,I1236283);
nand I_72531 (I1236611,I1236529,I1236594);
nand I_72532 (I1236082,I1236611,I1236560);
nand I_72533 (I1236079,I1236594,I1236478);
not I_72534 (I1236683,I3570);
DFFARX1 I_72535 (I1327533,I3563,I1236683,I1236709,);
and I_72536 (I1236717,I1236709,I1327560);
DFFARX1 I_72537 (I1236717,I3563,I1236683,I1236666,);
DFFARX1 I_72538 (I1327542,I3563,I1236683,I1236757,);
not I_72539 (I1236765,I1327551);
not I_72540 (I1236782,I1327554);
nand I_72541 (I1236799,I1236782,I1236765);
nor I_72542 (I1236654,I1236757,I1236799);
DFFARX1 I_72543 (I1236799,I3563,I1236683,I1236839,);
not I_72544 (I1236675,I1236839);
not I_72545 (I1236861,I1327548);
nand I_72546 (I1236878,I1236782,I1236861);
DFFARX1 I_72547 (I1236878,I3563,I1236683,I1236904,);
not I_72548 (I1236912,I1236904);
not I_72549 (I1236929,I1327536);
nand I_72550 (I1236946,I1236929,I1327539);
and I_72551 (I1236963,I1236765,I1236946);
nor I_72552 (I1236980,I1236878,I1236963);
DFFARX1 I_72553 (I1236980,I3563,I1236683,I1236651,);
DFFARX1 I_72554 (I1236963,I3563,I1236683,I1236672,);
nor I_72555 (I1237025,I1327536,I1327557);
nor I_72556 (I1236663,I1236878,I1237025);
or I_72557 (I1237056,I1327536,I1327557);
nor I_72558 (I1237073,I1327545,I1327533);
DFFARX1 I_72559 (I1237073,I3563,I1236683,I1237099,);
not I_72560 (I1237107,I1237099);
nor I_72561 (I1236669,I1237107,I1236912);
nand I_72562 (I1237138,I1237107,I1236757);
not I_72563 (I1237155,I1327545);
nand I_72564 (I1237172,I1237155,I1236861);
nand I_72565 (I1237189,I1237107,I1237172);
nand I_72566 (I1236660,I1237189,I1237138);
nand I_72567 (I1236657,I1237172,I1237056);
not I_72568 (I1237261,I3570);
DFFARX1 I_72569 (I709292,I3563,I1237261,I1237287,);
and I_72570 (I1237295,I1237287,I709280);
DFFARX1 I_72571 (I1237295,I3563,I1237261,I1237244,);
DFFARX1 I_72572 (I709283,I3563,I1237261,I1237335,);
not I_72573 (I1237343,I709277);
not I_72574 (I1237360,I709301);
nand I_72575 (I1237377,I1237360,I1237343);
nor I_72576 (I1237232,I1237335,I1237377);
DFFARX1 I_72577 (I1237377,I3563,I1237261,I1237417,);
not I_72578 (I1237253,I1237417);
not I_72579 (I1237439,I709289);
nand I_72580 (I1237456,I1237360,I1237439);
DFFARX1 I_72581 (I1237456,I3563,I1237261,I1237482,);
not I_72582 (I1237490,I1237482);
not I_72583 (I1237507,I709298);
nand I_72584 (I1237524,I1237507,I709295);
and I_72585 (I1237541,I1237343,I1237524);
nor I_72586 (I1237558,I1237456,I1237541);
DFFARX1 I_72587 (I1237558,I3563,I1237261,I1237229,);
DFFARX1 I_72588 (I1237541,I3563,I1237261,I1237250,);
nor I_72589 (I1237603,I709298,I709286);
nor I_72590 (I1237241,I1237456,I1237603);
or I_72591 (I1237634,I709298,I709286);
nor I_72592 (I1237651,I709277,I709280);
DFFARX1 I_72593 (I1237651,I3563,I1237261,I1237677,);
not I_72594 (I1237685,I1237677);
nor I_72595 (I1237247,I1237685,I1237490);
nand I_72596 (I1237716,I1237685,I1237335);
not I_72597 (I1237733,I709277);
nand I_72598 (I1237750,I1237733,I1237439);
nand I_72599 (I1237767,I1237685,I1237750);
nand I_72600 (I1237238,I1237767,I1237716);
nand I_72601 (I1237235,I1237750,I1237634);
not I_72602 (I1237839,I3570);
DFFARX1 I_72603 (I487138,I3563,I1237839,I1237865,);
and I_72604 (I1237873,I1237865,I487153);
DFFARX1 I_72605 (I1237873,I3563,I1237839,I1237822,);
DFFARX1 I_72606 (I487156,I3563,I1237839,I1237913,);
not I_72607 (I1237921,I487150);
not I_72608 (I1237938,I487165);
nand I_72609 (I1237955,I1237938,I1237921);
nor I_72610 (I1237810,I1237913,I1237955);
DFFARX1 I_72611 (I1237955,I3563,I1237839,I1237995,);
not I_72612 (I1237831,I1237995);
not I_72613 (I1238017,I487141);
nand I_72614 (I1238034,I1237938,I1238017);
DFFARX1 I_72615 (I1238034,I3563,I1237839,I1238060,);
not I_72616 (I1238068,I1238060);
not I_72617 (I1238085,I487144);
nand I_72618 (I1238102,I1238085,I487138);
and I_72619 (I1238119,I1237921,I1238102);
nor I_72620 (I1238136,I1238034,I1238119);
DFFARX1 I_72621 (I1238136,I3563,I1237839,I1237807,);
DFFARX1 I_72622 (I1238119,I3563,I1237839,I1237828,);
nor I_72623 (I1238181,I487144,I487147);
nor I_72624 (I1237819,I1238034,I1238181);
or I_72625 (I1238212,I487144,I487147);
nor I_72626 (I1238229,I487162,I487159);
DFFARX1 I_72627 (I1238229,I3563,I1237839,I1238255,);
not I_72628 (I1238263,I1238255);
nor I_72629 (I1237825,I1238263,I1238068);
nand I_72630 (I1238294,I1238263,I1237913);
not I_72631 (I1238311,I487162);
nand I_72632 (I1238328,I1238311,I1238017);
nand I_72633 (I1238345,I1238263,I1238328);
nand I_72634 (I1237816,I1238345,I1238294);
nand I_72635 (I1237813,I1238328,I1238212);
not I_72636 (I1238417,I3570);
DFFARX1 I_72637 (I378144,I3563,I1238417,I1238443,);
and I_72638 (I1238451,I1238443,I378129);
DFFARX1 I_72639 (I1238451,I3563,I1238417,I1238400,);
DFFARX1 I_72640 (I378135,I3563,I1238417,I1238491,);
not I_72641 (I1238499,I378117);
not I_72642 (I1238516,I378138);
nand I_72643 (I1238533,I1238516,I1238499);
nor I_72644 (I1238388,I1238491,I1238533);
DFFARX1 I_72645 (I1238533,I3563,I1238417,I1238573,);
not I_72646 (I1238409,I1238573);
not I_72647 (I1238595,I378141);
nand I_72648 (I1238612,I1238516,I1238595);
DFFARX1 I_72649 (I1238612,I3563,I1238417,I1238638,);
not I_72650 (I1238646,I1238638);
not I_72651 (I1238663,I378132);
nand I_72652 (I1238680,I1238663,I378120);
and I_72653 (I1238697,I1238499,I1238680);
nor I_72654 (I1238714,I1238612,I1238697);
DFFARX1 I_72655 (I1238714,I3563,I1238417,I1238385,);
DFFARX1 I_72656 (I1238697,I3563,I1238417,I1238406,);
nor I_72657 (I1238759,I378132,I378126);
nor I_72658 (I1238397,I1238612,I1238759);
or I_72659 (I1238790,I378132,I378126);
nor I_72660 (I1238807,I378123,I378117);
DFFARX1 I_72661 (I1238807,I3563,I1238417,I1238833,);
not I_72662 (I1238841,I1238833);
nor I_72663 (I1238403,I1238841,I1238646);
nand I_72664 (I1238872,I1238841,I1238491);
not I_72665 (I1238889,I378123);
nand I_72666 (I1238906,I1238889,I1238595);
nand I_72667 (I1238923,I1238841,I1238906);
nand I_72668 (I1238394,I1238923,I1238872);
nand I_72669 (I1238391,I1238906,I1238790);
not I_72670 (I1238995,I3570);
DFFARX1 I_72671 (I384995,I3563,I1238995,I1239021,);
and I_72672 (I1239029,I1239021,I384980);
DFFARX1 I_72673 (I1239029,I3563,I1238995,I1238978,);
DFFARX1 I_72674 (I384986,I3563,I1238995,I1239069,);
not I_72675 (I1239077,I384968);
not I_72676 (I1239094,I384989);
nand I_72677 (I1239111,I1239094,I1239077);
nor I_72678 (I1238966,I1239069,I1239111);
DFFARX1 I_72679 (I1239111,I3563,I1238995,I1239151,);
not I_72680 (I1238987,I1239151);
not I_72681 (I1239173,I384992);
nand I_72682 (I1239190,I1239094,I1239173);
DFFARX1 I_72683 (I1239190,I3563,I1238995,I1239216,);
not I_72684 (I1239224,I1239216);
not I_72685 (I1239241,I384983);
nand I_72686 (I1239258,I1239241,I384971);
and I_72687 (I1239275,I1239077,I1239258);
nor I_72688 (I1239292,I1239190,I1239275);
DFFARX1 I_72689 (I1239292,I3563,I1238995,I1238963,);
DFFARX1 I_72690 (I1239275,I3563,I1238995,I1238984,);
nor I_72691 (I1239337,I384983,I384977);
nor I_72692 (I1238975,I1239190,I1239337);
or I_72693 (I1239368,I384983,I384977);
nor I_72694 (I1239385,I384974,I384968);
DFFARX1 I_72695 (I1239385,I3563,I1238995,I1239411,);
not I_72696 (I1239419,I1239411);
nor I_72697 (I1238981,I1239419,I1239224);
nand I_72698 (I1239450,I1239419,I1239069);
not I_72699 (I1239467,I384974);
nand I_72700 (I1239484,I1239467,I1239173);
nand I_72701 (I1239501,I1239419,I1239484);
nand I_72702 (I1238972,I1239501,I1239450);
nand I_72703 (I1238969,I1239484,I1239368);
not I_72704 (I1239573,I3570);
DFFARX1 I_72705 (I719118,I3563,I1239573,I1239599,);
and I_72706 (I1239607,I1239599,I719106);
DFFARX1 I_72707 (I1239607,I3563,I1239573,I1239556,);
DFFARX1 I_72708 (I719109,I3563,I1239573,I1239647,);
not I_72709 (I1239655,I719103);
not I_72710 (I1239672,I719127);
nand I_72711 (I1239689,I1239672,I1239655);
nor I_72712 (I1239544,I1239647,I1239689);
DFFARX1 I_72713 (I1239689,I3563,I1239573,I1239729,);
not I_72714 (I1239565,I1239729);
not I_72715 (I1239751,I719115);
nand I_72716 (I1239768,I1239672,I1239751);
DFFARX1 I_72717 (I1239768,I3563,I1239573,I1239794,);
not I_72718 (I1239802,I1239794);
not I_72719 (I1239819,I719124);
nand I_72720 (I1239836,I1239819,I719121);
and I_72721 (I1239853,I1239655,I1239836);
nor I_72722 (I1239870,I1239768,I1239853);
DFFARX1 I_72723 (I1239870,I3563,I1239573,I1239541,);
DFFARX1 I_72724 (I1239853,I3563,I1239573,I1239562,);
nor I_72725 (I1239915,I719124,I719112);
nor I_72726 (I1239553,I1239768,I1239915);
or I_72727 (I1239946,I719124,I719112);
nor I_72728 (I1239963,I719103,I719106);
DFFARX1 I_72729 (I1239963,I3563,I1239573,I1239989,);
not I_72730 (I1239997,I1239989);
nor I_72731 (I1239559,I1239997,I1239802);
nand I_72732 (I1240028,I1239997,I1239647);
not I_72733 (I1240045,I719103);
nand I_72734 (I1240062,I1240045,I1239751);
nand I_72735 (I1240079,I1239997,I1240062);
nand I_72736 (I1239550,I1240079,I1240028);
nand I_72737 (I1239547,I1240062,I1239946);
not I_72738 (I1240151,I3570);
DFFARX1 I_72739 (I800038,I3563,I1240151,I1240177,);
and I_72740 (I1240185,I1240177,I800026);
DFFARX1 I_72741 (I1240185,I3563,I1240151,I1240134,);
DFFARX1 I_72742 (I800029,I3563,I1240151,I1240225,);
not I_72743 (I1240233,I800023);
not I_72744 (I1240250,I800047);
nand I_72745 (I1240267,I1240250,I1240233);
nor I_72746 (I1240122,I1240225,I1240267);
DFFARX1 I_72747 (I1240267,I3563,I1240151,I1240307,);
not I_72748 (I1240143,I1240307);
not I_72749 (I1240329,I800035);
nand I_72750 (I1240346,I1240250,I1240329);
DFFARX1 I_72751 (I1240346,I3563,I1240151,I1240372,);
not I_72752 (I1240380,I1240372);
not I_72753 (I1240397,I800044);
nand I_72754 (I1240414,I1240397,I800041);
and I_72755 (I1240431,I1240233,I1240414);
nor I_72756 (I1240448,I1240346,I1240431);
DFFARX1 I_72757 (I1240448,I3563,I1240151,I1240119,);
DFFARX1 I_72758 (I1240431,I3563,I1240151,I1240140,);
nor I_72759 (I1240493,I800044,I800032);
nor I_72760 (I1240131,I1240346,I1240493);
or I_72761 (I1240524,I800044,I800032);
nor I_72762 (I1240541,I800023,I800026);
DFFARX1 I_72763 (I1240541,I3563,I1240151,I1240567,);
not I_72764 (I1240575,I1240567);
nor I_72765 (I1240137,I1240575,I1240380);
nand I_72766 (I1240606,I1240575,I1240225);
not I_72767 (I1240623,I800023);
nand I_72768 (I1240640,I1240623,I1240329);
nand I_72769 (I1240657,I1240575,I1240640);
nand I_72770 (I1240128,I1240657,I1240606);
nand I_72771 (I1240125,I1240640,I1240524);
not I_72772 (I1240729,I3570);
DFFARX1 I_72773 (I158358,I3563,I1240729,I1240755,);
and I_72774 (I1240763,I1240755,I158382);
DFFARX1 I_72775 (I1240763,I3563,I1240729,I1240712,);
DFFARX1 I_72776 (I158358,I3563,I1240729,I1240803,);
not I_72777 (I1240811,I158376);
not I_72778 (I1240828,I158361);
nand I_72779 (I1240845,I1240828,I1240811);
nor I_72780 (I1240700,I1240803,I1240845);
DFFARX1 I_72781 (I1240845,I3563,I1240729,I1240885,);
not I_72782 (I1240721,I1240885);
not I_72783 (I1240907,I158370);
nand I_72784 (I1240924,I1240828,I1240907);
DFFARX1 I_72785 (I1240924,I3563,I1240729,I1240950,);
not I_72786 (I1240958,I1240950);
not I_72787 (I1240975,I158367);
nand I_72788 (I1240992,I1240975,I158364);
and I_72789 (I1241009,I1240811,I1240992);
nor I_72790 (I1241026,I1240924,I1241009);
DFFARX1 I_72791 (I1241026,I3563,I1240729,I1240697,);
DFFARX1 I_72792 (I1241009,I3563,I1240729,I1240718,);
nor I_72793 (I1241071,I158367,I158373);
nor I_72794 (I1240709,I1240924,I1241071);
or I_72795 (I1241102,I158367,I158373);
nor I_72796 (I1241119,I158379,I158385);
DFFARX1 I_72797 (I1241119,I3563,I1240729,I1241145,);
not I_72798 (I1241153,I1241145);
nor I_72799 (I1240715,I1241153,I1240958);
nand I_72800 (I1241184,I1241153,I1240803);
not I_72801 (I1241201,I158379);
nand I_72802 (I1241218,I1241201,I1240907);
nand I_72803 (I1241235,I1241153,I1241218);
nand I_72804 (I1240706,I1241235,I1241184);
nand I_72805 (I1240703,I1241218,I1241102);
not I_72806 (I1241307,I3570);
DFFARX1 I_72807 (I253558,I3563,I1241307,I1241333,);
and I_72808 (I1241341,I1241333,I253561);
DFFARX1 I_72809 (I1241341,I3563,I1241307,I1241290,);
DFFARX1 I_72810 (I253561,I3563,I1241307,I1241381,);
not I_72811 (I1241389,I253576);
not I_72812 (I1241406,I253582);
nand I_72813 (I1241423,I1241406,I1241389);
nor I_72814 (I1241278,I1241381,I1241423);
DFFARX1 I_72815 (I1241423,I3563,I1241307,I1241463,);
not I_72816 (I1241299,I1241463);
not I_72817 (I1241485,I253570);
nand I_72818 (I1241502,I1241406,I1241485);
DFFARX1 I_72819 (I1241502,I3563,I1241307,I1241528,);
not I_72820 (I1241536,I1241528);
not I_72821 (I1241553,I253567);
nand I_72822 (I1241570,I1241553,I253564);
and I_72823 (I1241587,I1241389,I1241570);
nor I_72824 (I1241604,I1241502,I1241587);
DFFARX1 I_72825 (I1241604,I3563,I1241307,I1241275,);
DFFARX1 I_72826 (I1241587,I3563,I1241307,I1241296,);
nor I_72827 (I1241649,I253567,I253558);
nor I_72828 (I1241287,I1241502,I1241649);
or I_72829 (I1241680,I253567,I253558);
nor I_72830 (I1241697,I253573,I253579);
DFFARX1 I_72831 (I1241697,I3563,I1241307,I1241723,);
not I_72832 (I1241731,I1241723);
nor I_72833 (I1241293,I1241731,I1241536);
nand I_72834 (I1241762,I1241731,I1241381);
not I_72835 (I1241779,I253573);
nand I_72836 (I1241796,I1241779,I1241485);
nand I_72837 (I1241813,I1241731,I1241796);
nand I_72838 (I1241284,I1241813,I1241762);
nand I_72839 (I1241281,I1241796,I1241680);
not I_72840 (I1241885,I3570);
DFFARX1 I_72841 (I487682,I3563,I1241885,I1241911,);
and I_72842 (I1241919,I1241911,I487697);
DFFARX1 I_72843 (I1241919,I3563,I1241885,I1241868,);
DFFARX1 I_72844 (I487700,I3563,I1241885,I1241959,);
not I_72845 (I1241967,I487694);
not I_72846 (I1241984,I487709);
nand I_72847 (I1242001,I1241984,I1241967);
nor I_72848 (I1241856,I1241959,I1242001);
DFFARX1 I_72849 (I1242001,I3563,I1241885,I1242041,);
not I_72850 (I1241877,I1242041);
not I_72851 (I1242063,I487685);
nand I_72852 (I1242080,I1241984,I1242063);
DFFARX1 I_72853 (I1242080,I3563,I1241885,I1242106,);
not I_72854 (I1242114,I1242106);
not I_72855 (I1242131,I487688);
nand I_72856 (I1242148,I1242131,I487682);
and I_72857 (I1242165,I1241967,I1242148);
nor I_72858 (I1242182,I1242080,I1242165);
DFFARX1 I_72859 (I1242182,I3563,I1241885,I1241853,);
DFFARX1 I_72860 (I1242165,I3563,I1241885,I1241874,);
nor I_72861 (I1242227,I487688,I487691);
nor I_72862 (I1241865,I1242080,I1242227);
or I_72863 (I1242258,I487688,I487691);
nor I_72864 (I1242275,I487706,I487703);
DFFARX1 I_72865 (I1242275,I3563,I1241885,I1242301,);
not I_72866 (I1242309,I1242301);
nor I_72867 (I1241871,I1242309,I1242114);
nand I_72868 (I1242340,I1242309,I1241959);
not I_72869 (I1242357,I487706);
nand I_72870 (I1242374,I1242357,I1242063);
nand I_72871 (I1242391,I1242309,I1242374);
nand I_72872 (I1241862,I1242391,I1242340);
nand I_72873 (I1241859,I1242374,I1242258);
not I_72874 (I1242463,I3570);
DFFARX1 I_72875 (I225593,I3563,I1242463,I1242489,);
and I_72876 (I1242497,I1242489,I225596);
DFFARX1 I_72877 (I1242497,I3563,I1242463,I1242446,);
DFFARX1 I_72878 (I225596,I3563,I1242463,I1242537,);
not I_72879 (I1242545,I225611);
not I_72880 (I1242562,I225617);
nand I_72881 (I1242579,I1242562,I1242545);
nor I_72882 (I1242434,I1242537,I1242579);
DFFARX1 I_72883 (I1242579,I3563,I1242463,I1242619,);
not I_72884 (I1242455,I1242619);
not I_72885 (I1242641,I225605);
nand I_72886 (I1242658,I1242562,I1242641);
DFFARX1 I_72887 (I1242658,I3563,I1242463,I1242684,);
not I_72888 (I1242692,I1242684);
not I_72889 (I1242709,I225602);
nand I_72890 (I1242726,I1242709,I225599);
and I_72891 (I1242743,I1242545,I1242726);
nor I_72892 (I1242760,I1242658,I1242743);
DFFARX1 I_72893 (I1242760,I3563,I1242463,I1242431,);
DFFARX1 I_72894 (I1242743,I3563,I1242463,I1242452,);
nor I_72895 (I1242805,I225602,I225593);
nor I_72896 (I1242443,I1242658,I1242805);
or I_72897 (I1242836,I225602,I225593);
nor I_72898 (I1242853,I225608,I225614);
DFFARX1 I_72899 (I1242853,I3563,I1242463,I1242879,);
not I_72900 (I1242887,I1242879);
nor I_72901 (I1242449,I1242887,I1242692);
nand I_72902 (I1242918,I1242887,I1242537);
not I_72903 (I1242935,I225608);
nand I_72904 (I1242952,I1242935,I1242641);
nand I_72905 (I1242969,I1242887,I1242952);
nand I_72906 (I1242440,I1242969,I1242918);
nand I_72907 (I1242437,I1242952,I1242836);
not I_72908 (I1243041,I3570);
DFFARX1 I_72909 (I330714,I3563,I1243041,I1243067,);
and I_72910 (I1243075,I1243067,I330699);
DFFARX1 I_72911 (I1243075,I3563,I1243041,I1243024,);
DFFARX1 I_72912 (I330705,I3563,I1243041,I1243115,);
not I_72913 (I1243123,I330687);
not I_72914 (I1243140,I330708);
nand I_72915 (I1243157,I1243140,I1243123);
nor I_72916 (I1243012,I1243115,I1243157);
DFFARX1 I_72917 (I1243157,I3563,I1243041,I1243197,);
not I_72918 (I1243033,I1243197);
not I_72919 (I1243219,I330711);
nand I_72920 (I1243236,I1243140,I1243219);
DFFARX1 I_72921 (I1243236,I3563,I1243041,I1243262,);
not I_72922 (I1243270,I1243262);
not I_72923 (I1243287,I330702);
nand I_72924 (I1243304,I1243287,I330690);
and I_72925 (I1243321,I1243123,I1243304);
nor I_72926 (I1243338,I1243236,I1243321);
DFFARX1 I_72927 (I1243338,I3563,I1243041,I1243009,);
DFFARX1 I_72928 (I1243321,I3563,I1243041,I1243030,);
nor I_72929 (I1243383,I330702,I330696);
nor I_72930 (I1243021,I1243236,I1243383);
or I_72931 (I1243414,I330702,I330696);
nor I_72932 (I1243431,I330693,I330687);
DFFARX1 I_72933 (I1243431,I3563,I1243041,I1243457,);
not I_72934 (I1243465,I1243457);
nor I_72935 (I1243027,I1243465,I1243270);
nand I_72936 (I1243496,I1243465,I1243115);
not I_72937 (I1243513,I330693);
nand I_72938 (I1243530,I1243513,I1243219);
nand I_72939 (I1243547,I1243465,I1243530);
nand I_72940 (I1243018,I1243547,I1243496);
nand I_72941 (I1243015,I1243530,I1243414);
not I_72942 (I1243619,I3570);
DFFARX1 I_72943 (I427298,I3563,I1243619,I1243645,);
and I_72944 (I1243653,I1243645,I427313);
DFFARX1 I_72945 (I1243653,I3563,I1243619,I1243602,);
DFFARX1 I_72946 (I427316,I3563,I1243619,I1243693,);
not I_72947 (I1243701,I427310);
not I_72948 (I1243718,I427325);
nand I_72949 (I1243735,I1243718,I1243701);
nor I_72950 (I1243590,I1243693,I1243735);
DFFARX1 I_72951 (I1243735,I3563,I1243619,I1243775,);
not I_72952 (I1243611,I1243775);
not I_72953 (I1243797,I427301);
nand I_72954 (I1243814,I1243718,I1243797);
DFFARX1 I_72955 (I1243814,I3563,I1243619,I1243840,);
not I_72956 (I1243848,I1243840);
not I_72957 (I1243865,I427304);
nand I_72958 (I1243882,I1243865,I427298);
and I_72959 (I1243899,I1243701,I1243882);
nor I_72960 (I1243916,I1243814,I1243899);
DFFARX1 I_72961 (I1243916,I3563,I1243619,I1243587,);
DFFARX1 I_72962 (I1243899,I3563,I1243619,I1243608,);
nor I_72963 (I1243961,I427304,I427307);
nor I_72964 (I1243599,I1243814,I1243961);
or I_72965 (I1243992,I427304,I427307);
nor I_72966 (I1244009,I427322,I427319);
DFFARX1 I_72967 (I1244009,I3563,I1243619,I1244035,);
not I_72968 (I1244043,I1244035);
nor I_72969 (I1243605,I1244043,I1243848);
nand I_72970 (I1244074,I1244043,I1243693);
not I_72971 (I1244091,I427322);
nand I_72972 (I1244108,I1244091,I1243797);
nand I_72973 (I1244125,I1244043,I1244108);
nand I_72974 (I1243596,I1244125,I1244074);
nand I_72975 (I1243593,I1244108,I1243992);
not I_72976 (I1244197,I3570);
DFFARX1 I_72977 (I1317255,I3563,I1244197,I1244223,);
and I_72978 (I1244231,I1244223,I1317237);
DFFARX1 I_72979 (I1244231,I3563,I1244197,I1244180,);
DFFARX1 I_72980 (I1317246,I3563,I1244197,I1244271,);
not I_72981 (I1244279,I1317231);
not I_72982 (I1244296,I1317243);
nand I_72983 (I1244313,I1244296,I1244279);
nor I_72984 (I1244168,I1244271,I1244313);
DFFARX1 I_72985 (I1244313,I3563,I1244197,I1244353,);
not I_72986 (I1244189,I1244353);
not I_72987 (I1244375,I1317234);
nand I_72988 (I1244392,I1244296,I1244375);
DFFARX1 I_72989 (I1244392,I3563,I1244197,I1244418,);
not I_72990 (I1244426,I1244418);
not I_72991 (I1244443,I1317231);
nand I_72992 (I1244460,I1244443,I1317234);
and I_72993 (I1244477,I1244279,I1244460);
nor I_72994 (I1244494,I1244392,I1244477);
DFFARX1 I_72995 (I1244494,I3563,I1244197,I1244165,);
DFFARX1 I_72996 (I1244477,I3563,I1244197,I1244186,);
nor I_72997 (I1244539,I1317231,I1317252);
nor I_72998 (I1244177,I1244392,I1244539);
or I_72999 (I1244570,I1317231,I1317252);
nor I_73000 (I1244587,I1317240,I1317249);
DFFARX1 I_73001 (I1244587,I3563,I1244197,I1244613,);
not I_73002 (I1244621,I1244613);
nor I_73003 (I1244183,I1244621,I1244426);
nand I_73004 (I1244652,I1244621,I1244271);
not I_73005 (I1244669,I1317240);
nand I_73006 (I1244686,I1244669,I1244375);
nand I_73007 (I1244703,I1244621,I1244686);
nand I_73008 (I1244174,I1244703,I1244652);
nand I_73009 (I1244171,I1244686,I1244570);
not I_73010 (I1244775,I3570);
DFFARX1 I_73011 (I801194,I3563,I1244775,I1244801,);
and I_73012 (I1244809,I1244801,I801182);
DFFARX1 I_73013 (I1244809,I3563,I1244775,I1244758,);
DFFARX1 I_73014 (I801185,I3563,I1244775,I1244849,);
not I_73015 (I1244857,I801179);
not I_73016 (I1244874,I801203);
nand I_73017 (I1244891,I1244874,I1244857);
nor I_73018 (I1244746,I1244849,I1244891);
DFFARX1 I_73019 (I1244891,I3563,I1244775,I1244931,);
not I_73020 (I1244767,I1244931);
not I_73021 (I1244953,I801191);
nand I_73022 (I1244970,I1244874,I1244953);
DFFARX1 I_73023 (I1244970,I3563,I1244775,I1244996,);
not I_73024 (I1245004,I1244996);
not I_73025 (I1245021,I801200);
nand I_73026 (I1245038,I1245021,I801197);
and I_73027 (I1245055,I1244857,I1245038);
nor I_73028 (I1245072,I1244970,I1245055);
DFFARX1 I_73029 (I1245072,I3563,I1244775,I1244743,);
DFFARX1 I_73030 (I1245055,I3563,I1244775,I1244764,);
nor I_73031 (I1245117,I801200,I801188);
nor I_73032 (I1244755,I1244970,I1245117);
or I_73033 (I1245148,I801200,I801188);
nor I_73034 (I1245165,I801179,I801182);
DFFARX1 I_73035 (I1245165,I3563,I1244775,I1245191,);
not I_73036 (I1245199,I1245191);
nor I_73037 (I1244761,I1245199,I1245004);
nand I_73038 (I1245230,I1245199,I1244849);
not I_73039 (I1245247,I801179);
nand I_73040 (I1245264,I1245247,I1244953);
nand I_73041 (I1245281,I1245199,I1245264);
nand I_73042 (I1244752,I1245281,I1245230);
nand I_73043 (I1244749,I1245264,I1245148);
not I_73044 (I1245353,I3570);
DFFARX1 I_73045 (I1324755,I3563,I1245353,I1245379,);
nand I_73046 (I1245387,I1245379,I1324740);
DFFARX1 I_73047 (I1324752,I3563,I1245353,I1245413,);
DFFARX1 I_73048 (I1245413,I3563,I1245353,I1245430,);
not I_73049 (I1245345,I1245430);
not I_73050 (I1245452,I1324746);
nor I_73051 (I1245469,I1324746,I1324737);
not I_73052 (I1245486,I1324731);
nand I_73053 (I1245503,I1245452,I1245486);
nor I_73054 (I1245520,I1324731,I1324746);
and I_73055 (I1245324,I1245520,I1245387);
not I_73056 (I1245551,I1324743);
nand I_73057 (I1245568,I1245551,I1324728);
nor I_73058 (I1245585,I1324743,I1324749);
not I_73059 (I1245602,I1245585);
nand I_73060 (I1245327,I1245469,I1245602);
DFFARX1 I_73061 (I1245585,I3563,I1245353,I1245342,);
nor I_73062 (I1245647,I1324734,I1324731);
nor I_73063 (I1245664,I1245647,I1324737);
and I_73064 (I1245681,I1245664,I1245568);
DFFARX1 I_73065 (I1245681,I3563,I1245353,I1245339,);
nor I_73066 (I1245336,I1245647,I1245503);
or I_73067 (I1245333,I1245585,I1245647);
nor I_73068 (I1245740,I1324734,I1324728);
DFFARX1 I_73069 (I1245740,I3563,I1245353,I1245766,);
not I_73070 (I1245774,I1245766);
nand I_73071 (I1245791,I1245774,I1245452);
nor I_73072 (I1245808,I1245791,I1324737);
DFFARX1 I_73073 (I1245808,I3563,I1245353,I1245321,);
nor I_73074 (I1245839,I1245774,I1245503);
nor I_73075 (I1245330,I1245647,I1245839);
not I_73076 (I1245897,I3570);
DFFARX1 I_73077 (I838993,I3563,I1245897,I1245923,);
nand I_73078 (I1245931,I1245923,I838987);
DFFARX1 I_73079 (I838990,I3563,I1245897,I1245957,);
DFFARX1 I_73080 (I1245957,I3563,I1245897,I1245974,);
not I_73081 (I1245889,I1245974);
not I_73082 (I1245996,I838996);
nor I_73083 (I1246013,I838996,I838990);
not I_73084 (I1246030,I838999);
nand I_73085 (I1246047,I1245996,I1246030);
nor I_73086 (I1246064,I838999,I838996);
and I_73087 (I1245868,I1246064,I1245931);
not I_73088 (I1246095,I839008);
nand I_73089 (I1246112,I1246095,I839002);
nor I_73090 (I1246129,I839008,I839005);
not I_73091 (I1246146,I1246129);
nand I_73092 (I1245871,I1246013,I1246146);
DFFARX1 I_73093 (I1246129,I3563,I1245897,I1245886,);
nor I_73094 (I1246191,I838987,I838999);
nor I_73095 (I1246208,I1246191,I838990);
and I_73096 (I1246225,I1246208,I1246112);
DFFARX1 I_73097 (I1246225,I3563,I1245897,I1245883,);
nor I_73098 (I1245880,I1246191,I1246047);
or I_73099 (I1245877,I1246129,I1246191);
nor I_73100 (I1246284,I838987,I838993);
DFFARX1 I_73101 (I1246284,I3563,I1245897,I1246310,);
not I_73102 (I1246318,I1246310);
nand I_73103 (I1246335,I1246318,I1245996);
nor I_73104 (I1246352,I1246335,I838990);
DFFARX1 I_73105 (I1246352,I3563,I1245897,I1245865,);
nor I_73106 (I1246383,I1246318,I1246047);
nor I_73107 (I1245874,I1246191,I1246383);
not I_73108 (I1246441,I3570);
DFFARX1 I_73109 (I597744,I3563,I1246441,I1246467,);
nand I_73110 (I1246475,I1246467,I597732);
DFFARX1 I_73111 (I597738,I3563,I1246441,I1246501,);
DFFARX1 I_73112 (I1246501,I3563,I1246441,I1246518,);
not I_73113 (I1246433,I1246518);
not I_73114 (I1246540,I597723);
nor I_73115 (I1246557,I597723,I597735);
not I_73116 (I1246574,I597726);
nand I_73117 (I1246591,I1246540,I1246574);
nor I_73118 (I1246608,I597726,I597723);
and I_73119 (I1246412,I1246608,I1246475);
not I_73120 (I1246639,I597741);
nand I_73121 (I1246656,I1246639,I597723);
nor I_73122 (I1246673,I597741,I597747);
not I_73123 (I1246690,I1246673);
nand I_73124 (I1246415,I1246557,I1246690);
DFFARX1 I_73125 (I1246673,I3563,I1246441,I1246430,);
nor I_73126 (I1246735,I597729,I597726);
nor I_73127 (I1246752,I1246735,I597735);
and I_73128 (I1246769,I1246752,I1246656);
DFFARX1 I_73129 (I1246769,I3563,I1246441,I1246427,);
nor I_73130 (I1246424,I1246735,I1246591);
or I_73131 (I1246421,I1246673,I1246735);
nor I_73132 (I1246828,I597729,I597726);
DFFARX1 I_73133 (I1246828,I3563,I1246441,I1246854,);
not I_73134 (I1246862,I1246854);
nand I_73135 (I1246879,I1246862,I1246540);
nor I_73136 (I1246896,I1246879,I597735);
DFFARX1 I_73137 (I1246896,I3563,I1246441,I1246409,);
nor I_73138 (I1246927,I1246862,I1246591);
nor I_73139 (I1246418,I1246735,I1246927);
not I_73140 (I1246985,I3570);
DFFARX1 I_73141 (I665930,I3563,I1246985,I1247011,);
nand I_73142 (I1247019,I1247011,I665945);
DFFARX1 I_73143 (I665939,I3563,I1246985,I1247045,);
DFFARX1 I_73144 (I1247045,I3563,I1246985,I1247062,);
not I_73145 (I1246977,I1247062);
not I_73146 (I1247084,I665942);
nor I_73147 (I1247101,I665942,I665948);
not I_73148 (I1247118,I665930);
nand I_73149 (I1247135,I1247084,I1247118);
nor I_73150 (I1247152,I665930,I665942);
and I_73151 (I1246956,I1247152,I1247019);
not I_73152 (I1247183,I665927);
nand I_73153 (I1247200,I1247183,I665933);
nor I_73154 (I1247217,I665927,I665927);
not I_73155 (I1247234,I1247217);
nand I_73156 (I1246959,I1247101,I1247234);
DFFARX1 I_73157 (I1247217,I3563,I1246985,I1246974,);
nor I_73158 (I1247279,I665936,I665930);
nor I_73159 (I1247296,I1247279,I665948);
and I_73160 (I1247313,I1247296,I1247200);
DFFARX1 I_73161 (I1247313,I3563,I1246985,I1246971,);
nor I_73162 (I1246968,I1247279,I1247135);
or I_73163 (I1246965,I1247217,I1247279);
nor I_73164 (I1247372,I665936,I665951);
DFFARX1 I_73165 (I1247372,I3563,I1246985,I1247398,);
not I_73166 (I1247406,I1247398);
nand I_73167 (I1247423,I1247406,I1247084);
nor I_73168 (I1247440,I1247423,I665948);
DFFARX1 I_73169 (I1247440,I3563,I1246985,I1246953,);
nor I_73170 (I1247471,I1247406,I1247135);
nor I_73171 (I1246962,I1247279,I1247471);
not I_73172 (I1247529,I3570);
DFFARX1 I_73173 (I235122,I3563,I1247529,I1247555,);
nand I_73174 (I1247563,I1247555,I235137);
DFFARX1 I_73175 (I235134,I3563,I1247529,I1247589,);
DFFARX1 I_73176 (I1247589,I3563,I1247529,I1247606,);
not I_73177 (I1247521,I1247606);
not I_73178 (I1247628,I235113);
nor I_73179 (I1247645,I235113,I235119);
not I_73180 (I1247662,I235125);
nand I_73181 (I1247679,I1247628,I1247662);
nor I_73182 (I1247696,I235125,I235113);
and I_73183 (I1247500,I1247696,I1247563);
not I_73184 (I1247727,I235131);
nand I_73185 (I1247744,I1247727,I235113);
nor I_73186 (I1247761,I235131,I235116);
not I_73187 (I1247778,I1247761);
nand I_73188 (I1247503,I1247645,I1247778);
DFFARX1 I_73189 (I1247761,I3563,I1247529,I1247518,);
nor I_73190 (I1247823,I235116,I235125);
nor I_73191 (I1247840,I1247823,I235119);
and I_73192 (I1247857,I1247840,I1247744);
DFFARX1 I_73193 (I1247857,I3563,I1247529,I1247515,);
nor I_73194 (I1247512,I1247823,I1247679);
or I_73195 (I1247509,I1247761,I1247823);
nor I_73196 (I1247916,I235116,I235128);
DFFARX1 I_73197 (I1247916,I3563,I1247529,I1247942,);
not I_73198 (I1247950,I1247942);
nand I_73199 (I1247967,I1247950,I1247628);
nor I_73200 (I1247984,I1247967,I235119);
DFFARX1 I_73201 (I1247984,I3563,I1247529,I1247497,);
nor I_73202 (I1248015,I1247950,I1247679);
nor I_73203 (I1247506,I1247823,I1248015);
not I_73204 (I1248073,I3570);
DFFARX1 I_73205 (I974953,I3563,I1248073,I1248099,);
nand I_73206 (I1248107,I1248099,I974953);
DFFARX1 I_73207 (I974965,I3563,I1248073,I1248133,);
DFFARX1 I_73208 (I1248133,I3563,I1248073,I1248150,);
not I_73209 (I1248065,I1248150);
not I_73210 (I1248172,I974959);
nor I_73211 (I1248189,I974959,I974980);
not I_73212 (I1248206,I974968);
nand I_73213 (I1248223,I1248172,I1248206);
nor I_73214 (I1248240,I974968,I974959);
and I_73215 (I1248044,I1248240,I1248107);
not I_73216 (I1248271,I974962);
nand I_73217 (I1248288,I1248271,I974977);
nor I_73218 (I1248305,I974962,I974971);
not I_73219 (I1248322,I1248305);
nand I_73220 (I1248047,I1248189,I1248322);
DFFARX1 I_73221 (I1248305,I3563,I1248073,I1248062,);
nor I_73222 (I1248367,I974974,I974968);
nor I_73223 (I1248384,I1248367,I974980);
and I_73224 (I1248401,I1248384,I1248288);
DFFARX1 I_73225 (I1248401,I3563,I1248073,I1248059,);
nor I_73226 (I1248056,I1248367,I1248223);
or I_73227 (I1248053,I1248305,I1248367);
nor I_73228 (I1248460,I974974,I974956);
DFFARX1 I_73229 (I1248460,I3563,I1248073,I1248486,);
not I_73230 (I1248494,I1248486);
nand I_73231 (I1248511,I1248494,I1248172);
nor I_73232 (I1248528,I1248511,I974980);
DFFARX1 I_73233 (I1248528,I3563,I1248073,I1248041,);
nor I_73234 (I1248559,I1248494,I1248223);
nor I_73235 (I1248050,I1248367,I1248559);
not I_73236 (I1248617,I3570);
DFFARX1 I_73237 (I630112,I3563,I1248617,I1248643,);
nand I_73238 (I1248651,I1248643,I630100);
DFFARX1 I_73239 (I630106,I3563,I1248617,I1248677,);
DFFARX1 I_73240 (I1248677,I3563,I1248617,I1248694,);
not I_73241 (I1248609,I1248694);
not I_73242 (I1248716,I630091);
nor I_73243 (I1248733,I630091,I630103);
not I_73244 (I1248750,I630094);
nand I_73245 (I1248767,I1248716,I1248750);
nor I_73246 (I1248784,I630094,I630091);
and I_73247 (I1248588,I1248784,I1248651);
not I_73248 (I1248815,I630109);
nand I_73249 (I1248832,I1248815,I630091);
nor I_73250 (I1248849,I630109,I630115);
not I_73251 (I1248866,I1248849);
nand I_73252 (I1248591,I1248733,I1248866);
DFFARX1 I_73253 (I1248849,I3563,I1248617,I1248606,);
nor I_73254 (I1248911,I630097,I630094);
nor I_73255 (I1248928,I1248911,I630103);
and I_73256 (I1248945,I1248928,I1248832);
DFFARX1 I_73257 (I1248945,I3563,I1248617,I1248603,);
nor I_73258 (I1248600,I1248911,I1248767);
or I_73259 (I1248597,I1248849,I1248911);
nor I_73260 (I1249004,I630097,I630094);
DFFARX1 I_73261 (I1249004,I3563,I1248617,I1249030,);
not I_73262 (I1249038,I1249030);
nand I_73263 (I1249055,I1249038,I1248716);
nor I_73264 (I1249072,I1249055,I630103);
DFFARX1 I_73265 (I1249072,I3563,I1248617,I1248585,);
nor I_73266 (I1249103,I1249038,I1248767);
nor I_73267 (I1248594,I1248911,I1249103);
not I_73268 (I1249161,I3570);
DFFARX1 I_73269 (I476826,I3563,I1249161,I1249187,);
nand I_73270 (I1249195,I1249187,I476823);
DFFARX1 I_73271 (I476802,I3563,I1249161,I1249221,);
DFFARX1 I_73272 (I1249221,I3563,I1249161,I1249238,);
not I_73273 (I1249153,I1249238);
not I_73274 (I1249260,I476817);
nor I_73275 (I1249277,I476817,I476820);
not I_73276 (I1249294,I476811);
nand I_73277 (I1249311,I1249260,I1249294);
nor I_73278 (I1249328,I476811,I476817);
and I_73279 (I1249132,I1249328,I1249195);
not I_73280 (I1249359,I476808);
nand I_73281 (I1249376,I1249359,I476829);
nor I_73282 (I1249393,I476808,I476805);
not I_73283 (I1249410,I1249393);
nand I_73284 (I1249135,I1249277,I1249410);
DFFARX1 I_73285 (I1249393,I3563,I1249161,I1249150,);
nor I_73286 (I1249455,I476814,I476811);
nor I_73287 (I1249472,I1249455,I476820);
and I_73288 (I1249489,I1249472,I1249376);
DFFARX1 I_73289 (I1249489,I3563,I1249161,I1249147,);
nor I_73290 (I1249144,I1249455,I1249311);
or I_73291 (I1249141,I1249393,I1249455);
nor I_73292 (I1249548,I476814,I476802);
DFFARX1 I_73293 (I1249548,I3563,I1249161,I1249574,);
not I_73294 (I1249582,I1249574);
nand I_73295 (I1249599,I1249582,I1249260);
nor I_73296 (I1249616,I1249599,I476820);
DFFARX1 I_73297 (I1249616,I3563,I1249161,I1249129,);
nor I_73298 (I1249647,I1249582,I1249311);
nor I_73299 (I1249138,I1249455,I1249647);
not I_73300 (I1249705,I3570);
DFFARX1 I_73301 (I746272,I3563,I1249705,I1249731,);
nand I_73302 (I1249739,I1249731,I746287);
DFFARX1 I_73303 (I746281,I3563,I1249705,I1249765,);
DFFARX1 I_73304 (I1249765,I3563,I1249705,I1249782,);
not I_73305 (I1249697,I1249782);
not I_73306 (I1249804,I746284);
nor I_73307 (I1249821,I746284,I746290);
not I_73308 (I1249838,I746272);
nand I_73309 (I1249855,I1249804,I1249838);
nor I_73310 (I1249872,I746272,I746284);
and I_73311 (I1249676,I1249872,I1249739);
not I_73312 (I1249903,I746269);
nand I_73313 (I1249920,I1249903,I746275);
nor I_73314 (I1249937,I746269,I746269);
not I_73315 (I1249954,I1249937);
nand I_73316 (I1249679,I1249821,I1249954);
DFFARX1 I_73317 (I1249937,I3563,I1249705,I1249694,);
nor I_73318 (I1249999,I746278,I746272);
nor I_73319 (I1250016,I1249999,I746290);
and I_73320 (I1250033,I1250016,I1249920);
DFFARX1 I_73321 (I1250033,I3563,I1249705,I1249691,);
nor I_73322 (I1249688,I1249999,I1249855);
or I_73323 (I1249685,I1249937,I1249999);
nor I_73324 (I1250092,I746278,I746293);
DFFARX1 I_73325 (I1250092,I3563,I1249705,I1250118,);
not I_73326 (I1250126,I1250118);
nand I_73327 (I1250143,I1250126,I1249804);
nor I_73328 (I1250160,I1250143,I746290);
DFFARX1 I_73329 (I1250160,I3563,I1249705,I1249673,);
nor I_73330 (I1250191,I1250126,I1249855);
nor I_73331 (I1249682,I1249999,I1250191);
not I_73332 (I1250249,I3570);
DFFARX1 I_73333 (I369697,I3563,I1250249,I1250275,);
nand I_73334 (I1250283,I1250275,I369700);
DFFARX1 I_73335 (I369694,I3563,I1250249,I1250309,);
DFFARX1 I_73336 (I1250309,I3563,I1250249,I1250326,);
not I_73337 (I1250241,I1250326);
not I_73338 (I1250348,I369703);
nor I_73339 (I1250365,I369703,I369688);
not I_73340 (I1250382,I369712);
nand I_73341 (I1250399,I1250348,I1250382);
nor I_73342 (I1250416,I369712,I369703);
and I_73343 (I1250220,I1250416,I1250283);
not I_73344 (I1250447,I369691);
nand I_73345 (I1250464,I1250447,I369709);
nor I_73346 (I1250481,I369691,I369685);
not I_73347 (I1250498,I1250481);
nand I_73348 (I1250223,I1250365,I1250498);
DFFARX1 I_73349 (I1250481,I3563,I1250249,I1250238,);
nor I_73350 (I1250543,I369706,I369712);
nor I_73351 (I1250560,I1250543,I369688);
and I_73352 (I1250577,I1250560,I1250464);
DFFARX1 I_73353 (I1250577,I3563,I1250249,I1250235,);
nor I_73354 (I1250232,I1250543,I1250399);
or I_73355 (I1250229,I1250481,I1250543);
nor I_73356 (I1250636,I369706,I369685);
DFFARX1 I_73357 (I1250636,I3563,I1250249,I1250662,);
not I_73358 (I1250670,I1250662);
nand I_73359 (I1250687,I1250670,I1250348);
nor I_73360 (I1250704,I1250687,I369688);
DFFARX1 I_73361 (I1250704,I3563,I1250249,I1250217,);
nor I_73362 (I1250735,I1250670,I1250399);
nor I_73363 (I1250226,I1250543,I1250735);
not I_73364 (I1250793,I3570);
DFFARX1 I_73365 (I277962,I3563,I1250793,I1250819,);
nand I_73366 (I1250827,I1250819,I277977);
DFFARX1 I_73367 (I277974,I3563,I1250793,I1250853,);
DFFARX1 I_73368 (I1250853,I3563,I1250793,I1250870,);
not I_73369 (I1250785,I1250870);
not I_73370 (I1250892,I277953);
nor I_73371 (I1250909,I277953,I277959);
not I_73372 (I1250926,I277965);
nand I_73373 (I1250943,I1250892,I1250926);
nor I_73374 (I1250960,I277965,I277953);
and I_73375 (I1250764,I1250960,I1250827);
not I_73376 (I1250991,I277971);
nand I_73377 (I1251008,I1250991,I277953);
nor I_73378 (I1251025,I277971,I277956);
not I_73379 (I1251042,I1251025);
nand I_73380 (I1250767,I1250909,I1251042);
DFFARX1 I_73381 (I1251025,I3563,I1250793,I1250782,);
nor I_73382 (I1251087,I277956,I277965);
nor I_73383 (I1251104,I1251087,I277959);
and I_73384 (I1251121,I1251104,I1251008);
DFFARX1 I_73385 (I1251121,I3563,I1250793,I1250779,);
nor I_73386 (I1250776,I1251087,I1250943);
or I_73387 (I1250773,I1251025,I1251087);
nor I_73388 (I1251180,I277956,I277968);
DFFARX1 I_73389 (I1251180,I3563,I1250793,I1251206,);
not I_73390 (I1251214,I1251206);
nand I_73391 (I1251231,I1251214,I1250892);
nor I_73392 (I1251248,I1251231,I277959);
DFFARX1 I_73393 (I1251248,I3563,I1250793,I1250761,);
nor I_73394 (I1251279,I1251214,I1250943);
nor I_73395 (I1250770,I1251087,I1251279);
not I_73396 (I1251337,I3570);
DFFARX1 I_73397 (I689628,I3563,I1251337,I1251363,);
nand I_73398 (I1251371,I1251363,I689643);
DFFARX1 I_73399 (I689637,I3563,I1251337,I1251397,);
DFFARX1 I_73400 (I1251397,I3563,I1251337,I1251414,);
not I_73401 (I1251329,I1251414);
not I_73402 (I1251436,I689640);
nor I_73403 (I1251453,I689640,I689646);
not I_73404 (I1251470,I689628);
nand I_73405 (I1251487,I1251436,I1251470);
nor I_73406 (I1251504,I689628,I689640);
and I_73407 (I1251308,I1251504,I1251371);
not I_73408 (I1251535,I689625);
nand I_73409 (I1251552,I1251535,I689631);
nor I_73410 (I1251569,I689625,I689625);
not I_73411 (I1251586,I1251569);
nand I_73412 (I1251311,I1251453,I1251586);
DFFARX1 I_73413 (I1251569,I3563,I1251337,I1251326,);
nor I_73414 (I1251631,I689634,I689628);
nor I_73415 (I1251648,I1251631,I689646);
and I_73416 (I1251665,I1251648,I1251552);
DFFARX1 I_73417 (I1251665,I3563,I1251337,I1251323,);
nor I_73418 (I1251320,I1251631,I1251487);
or I_73419 (I1251317,I1251569,I1251631);
nor I_73420 (I1251724,I689634,I689649);
DFFARX1 I_73421 (I1251724,I3563,I1251337,I1251750,);
not I_73422 (I1251758,I1251750);
nand I_73423 (I1251775,I1251758,I1251436);
nor I_73424 (I1251792,I1251775,I689646);
DFFARX1 I_73425 (I1251792,I3563,I1251337,I1251305,);
nor I_73426 (I1251823,I1251758,I1251487);
nor I_73427 (I1251314,I1251631,I1251823);
not I_73428 (I1251881,I3570);
DFFARX1 I_73429 (I344928,I3563,I1251881,I1251907,);
nand I_73430 (I1251915,I1251907,I344931);
DFFARX1 I_73431 (I344925,I3563,I1251881,I1251941,);
DFFARX1 I_73432 (I1251941,I3563,I1251881,I1251958,);
not I_73433 (I1251873,I1251958);
not I_73434 (I1251980,I344934);
nor I_73435 (I1251997,I344934,I344919);
not I_73436 (I1252014,I344943);
nand I_73437 (I1252031,I1251980,I1252014);
nor I_73438 (I1252048,I344943,I344934);
and I_73439 (I1251852,I1252048,I1251915);
not I_73440 (I1252079,I344922);
nand I_73441 (I1252096,I1252079,I344940);
nor I_73442 (I1252113,I344922,I344916);
not I_73443 (I1252130,I1252113);
nand I_73444 (I1251855,I1251997,I1252130);
DFFARX1 I_73445 (I1252113,I3563,I1251881,I1251870,);
nor I_73446 (I1252175,I344937,I344943);
nor I_73447 (I1252192,I1252175,I344919);
and I_73448 (I1252209,I1252192,I1252096);
DFFARX1 I_73449 (I1252209,I3563,I1251881,I1251867,);
nor I_73450 (I1251864,I1252175,I1252031);
or I_73451 (I1251861,I1252113,I1252175);
nor I_73452 (I1252268,I344937,I344916);
DFFARX1 I_73453 (I1252268,I3563,I1251881,I1252294,);
not I_73454 (I1252302,I1252294);
nand I_73455 (I1252319,I1252302,I1251980);
nor I_73456 (I1252336,I1252319,I344919);
DFFARX1 I_73457 (I1252336,I3563,I1251881,I1251849,);
nor I_73458 (I1252367,I1252302,I1252031);
nor I_73459 (I1251858,I1252175,I1252367);
not I_73460 (I1252425,I3570);
DFFARX1 I_73461 (I1225693,I3563,I1252425,I1252451,);
nand I_73462 (I1252459,I1252451,I1225672);
DFFARX1 I_73463 (I1225669,I3563,I1252425,I1252485,);
DFFARX1 I_73464 (I1252485,I3563,I1252425,I1252502,);
not I_73465 (I1252417,I1252502);
not I_73466 (I1252524,I1225681);
nor I_73467 (I1252541,I1225681,I1225690);
not I_73468 (I1252558,I1225678);
nand I_73469 (I1252575,I1252524,I1252558);
nor I_73470 (I1252592,I1225678,I1225681);
and I_73471 (I1252396,I1252592,I1252459);
not I_73472 (I1252623,I1225687);
nand I_73473 (I1252640,I1252623,I1225684);
nor I_73474 (I1252657,I1225687,I1225669);
not I_73475 (I1252674,I1252657);
nand I_73476 (I1252399,I1252541,I1252674);
DFFARX1 I_73477 (I1252657,I3563,I1252425,I1252414,);
nor I_73478 (I1252719,I1225672,I1225678);
nor I_73479 (I1252736,I1252719,I1225690);
and I_73480 (I1252753,I1252736,I1252640);
DFFARX1 I_73481 (I1252753,I3563,I1252425,I1252411,);
nor I_73482 (I1252408,I1252719,I1252575);
or I_73483 (I1252405,I1252657,I1252719);
nor I_73484 (I1252812,I1225672,I1225675);
DFFARX1 I_73485 (I1252812,I3563,I1252425,I1252838,);
not I_73486 (I1252846,I1252838);
nand I_73487 (I1252863,I1252846,I1252524);
nor I_73488 (I1252880,I1252863,I1225690);
DFFARX1 I_73489 (I1252880,I3563,I1252425,I1252393,);
nor I_73490 (I1252911,I1252846,I1252575);
nor I_73491 (I1252402,I1252719,I1252911);
not I_73492 (I1252969,I3570);
DFFARX1 I_73493 (I604102,I3563,I1252969,I1252995,);
nand I_73494 (I1253003,I1252995,I604090);
DFFARX1 I_73495 (I604096,I3563,I1252969,I1253029,);
DFFARX1 I_73496 (I1253029,I3563,I1252969,I1253046,);
not I_73497 (I1252961,I1253046);
not I_73498 (I1253068,I604081);
nor I_73499 (I1253085,I604081,I604093);
not I_73500 (I1253102,I604084);
nand I_73501 (I1253119,I1253068,I1253102);
nor I_73502 (I1253136,I604084,I604081);
and I_73503 (I1252940,I1253136,I1253003);
not I_73504 (I1253167,I604099);
nand I_73505 (I1253184,I1253167,I604081);
nor I_73506 (I1253201,I604099,I604105);
not I_73507 (I1253218,I1253201);
nand I_73508 (I1252943,I1253085,I1253218);
DFFARX1 I_73509 (I1253201,I3563,I1252969,I1252958,);
nor I_73510 (I1253263,I604087,I604084);
nor I_73511 (I1253280,I1253263,I604093);
and I_73512 (I1253297,I1253280,I1253184);
DFFARX1 I_73513 (I1253297,I3563,I1252969,I1252955,);
nor I_73514 (I1252952,I1253263,I1253119);
or I_73515 (I1252949,I1253201,I1253263);
nor I_73516 (I1253356,I604087,I604084);
DFFARX1 I_73517 (I1253356,I3563,I1252969,I1253382,);
not I_73518 (I1253390,I1253382);
nand I_73519 (I1253407,I1253390,I1253068);
nor I_73520 (I1253424,I1253407,I604093);
DFFARX1 I_73521 (I1253424,I3563,I1252969,I1252937,);
nor I_73522 (I1253455,I1253390,I1253119);
nor I_73523 (I1252946,I1253263,I1253455);
not I_73524 (I1253513,I3570);
DFFARX1 I_73525 (I730088,I3563,I1253513,I1253539,);
nand I_73526 (I1253547,I1253539,I730103);
DFFARX1 I_73527 (I730097,I3563,I1253513,I1253573,);
DFFARX1 I_73528 (I1253573,I3563,I1253513,I1253590,);
not I_73529 (I1253505,I1253590);
not I_73530 (I1253612,I730100);
nor I_73531 (I1253629,I730100,I730106);
not I_73532 (I1253646,I730088);
nand I_73533 (I1253663,I1253612,I1253646);
nor I_73534 (I1253680,I730088,I730100);
and I_73535 (I1253484,I1253680,I1253547);
not I_73536 (I1253711,I730085);
nand I_73537 (I1253728,I1253711,I730091);
nor I_73538 (I1253745,I730085,I730085);
not I_73539 (I1253762,I1253745);
nand I_73540 (I1253487,I1253629,I1253762);
DFFARX1 I_73541 (I1253745,I3563,I1253513,I1253502,);
nor I_73542 (I1253807,I730094,I730088);
nor I_73543 (I1253824,I1253807,I730106);
and I_73544 (I1253841,I1253824,I1253728);
DFFARX1 I_73545 (I1253841,I3563,I1253513,I1253499,);
nor I_73546 (I1253496,I1253807,I1253663);
or I_73547 (I1253493,I1253745,I1253807);
nor I_73548 (I1253900,I730094,I730109);
DFFARX1 I_73549 (I1253900,I3563,I1253513,I1253926,);
not I_73550 (I1253934,I1253926);
nand I_73551 (I1253951,I1253934,I1253612);
nor I_73552 (I1253968,I1253951,I730106);
DFFARX1 I_73553 (I1253968,I3563,I1253513,I1253481,);
nor I_73554 (I1253999,I1253934,I1253663);
nor I_73555 (I1253490,I1253807,I1253999);
not I_73556 (I1254057,I3570);
DFFARX1 I_73557 (I1021465,I3563,I1254057,I1254083,);
nand I_73558 (I1254091,I1254083,I1021465);
DFFARX1 I_73559 (I1021477,I3563,I1254057,I1254117,);
DFFARX1 I_73560 (I1254117,I3563,I1254057,I1254134,);
not I_73561 (I1254049,I1254134);
not I_73562 (I1254156,I1021471);
nor I_73563 (I1254173,I1021471,I1021492);
not I_73564 (I1254190,I1021480);
nand I_73565 (I1254207,I1254156,I1254190);
nor I_73566 (I1254224,I1021480,I1021471);
and I_73567 (I1254028,I1254224,I1254091);
not I_73568 (I1254255,I1021474);
nand I_73569 (I1254272,I1254255,I1021489);
nor I_73570 (I1254289,I1021474,I1021483);
not I_73571 (I1254306,I1254289);
nand I_73572 (I1254031,I1254173,I1254306);
DFFARX1 I_73573 (I1254289,I3563,I1254057,I1254046,);
nor I_73574 (I1254351,I1021486,I1021480);
nor I_73575 (I1254368,I1254351,I1021492);
and I_73576 (I1254385,I1254368,I1254272);
DFFARX1 I_73577 (I1254385,I3563,I1254057,I1254043,);
nor I_73578 (I1254040,I1254351,I1254207);
or I_73579 (I1254037,I1254289,I1254351);
nor I_73580 (I1254444,I1021486,I1021468);
DFFARX1 I_73581 (I1254444,I3563,I1254057,I1254470,);
not I_73582 (I1254478,I1254470);
nand I_73583 (I1254495,I1254478,I1254156);
nor I_73584 (I1254512,I1254495,I1021492);
DFFARX1 I_73585 (I1254512,I3563,I1254057,I1254025,);
nor I_73586 (I1254543,I1254478,I1254207);
nor I_73587 (I1254034,I1254351,I1254543);
not I_73588 (I1254601,I3570);
DFFARX1 I_73589 (I1082581,I3563,I1254601,I1254627,);
nand I_73590 (I1254635,I1254627,I1082569);
DFFARX1 I_73591 (I1082563,I3563,I1254601,I1254661,);
DFFARX1 I_73592 (I1254661,I3563,I1254601,I1254678,);
not I_73593 (I1254593,I1254678);
not I_73594 (I1254700,I1082563);
nor I_73595 (I1254717,I1082563,I1082575);
not I_73596 (I1254734,I1082572);
nand I_73597 (I1254751,I1254700,I1254734);
nor I_73598 (I1254768,I1082572,I1082563);
and I_73599 (I1254572,I1254768,I1254635);
not I_73600 (I1254799,I1082566);
nand I_73601 (I1254816,I1254799,I1082578);
nor I_73602 (I1254833,I1082566,I1082584);
not I_73603 (I1254850,I1254833);
nand I_73604 (I1254575,I1254717,I1254850);
DFFARX1 I_73605 (I1254833,I3563,I1254601,I1254590,);
nor I_73606 (I1254895,I1082569,I1082572);
nor I_73607 (I1254912,I1254895,I1082575);
and I_73608 (I1254929,I1254912,I1254816);
DFFARX1 I_73609 (I1254929,I3563,I1254601,I1254587,);
nor I_73610 (I1254584,I1254895,I1254751);
or I_73611 (I1254581,I1254833,I1254895);
nor I_73612 (I1254988,I1082569,I1082566);
DFFARX1 I_73613 (I1254988,I3563,I1254601,I1255014,);
not I_73614 (I1255022,I1255014);
nand I_73615 (I1255039,I1255022,I1254700);
nor I_73616 (I1255056,I1255039,I1082575);
DFFARX1 I_73617 (I1255056,I3563,I1254601,I1254569,);
nor I_73618 (I1255087,I1255022,I1254751);
nor I_73619 (I1254578,I1254895,I1255087);
not I_73620 (I1255145,I3570);
DFFARX1 I_73621 (I518170,I3563,I1255145,I1255171,);
nand I_73622 (I1255179,I1255171,I518167);
DFFARX1 I_73623 (I518146,I3563,I1255145,I1255205,);
DFFARX1 I_73624 (I1255205,I3563,I1255145,I1255222,);
not I_73625 (I1255137,I1255222);
not I_73626 (I1255244,I518161);
nor I_73627 (I1255261,I518161,I518164);
not I_73628 (I1255278,I518155);
nand I_73629 (I1255295,I1255244,I1255278);
nor I_73630 (I1255312,I518155,I518161);
and I_73631 (I1255116,I1255312,I1255179);
not I_73632 (I1255343,I518152);
nand I_73633 (I1255360,I1255343,I518173);
nor I_73634 (I1255377,I518152,I518149);
not I_73635 (I1255394,I1255377);
nand I_73636 (I1255119,I1255261,I1255394);
DFFARX1 I_73637 (I1255377,I3563,I1255145,I1255134,);
nor I_73638 (I1255439,I518158,I518155);
nor I_73639 (I1255456,I1255439,I518164);
and I_73640 (I1255473,I1255456,I1255360);
DFFARX1 I_73641 (I1255473,I3563,I1255145,I1255131,);
nor I_73642 (I1255128,I1255439,I1255295);
or I_73643 (I1255125,I1255377,I1255439);
nor I_73644 (I1255532,I518158,I518146);
DFFARX1 I_73645 (I1255532,I3563,I1255145,I1255558,);
not I_73646 (I1255566,I1255558);
nand I_73647 (I1255583,I1255566,I1255244);
nor I_73648 (I1255600,I1255583,I518164);
DFFARX1 I_73649 (I1255600,I3563,I1255145,I1255113,);
nor I_73650 (I1255631,I1255566,I1255295);
nor I_73651 (I1255122,I1255439,I1255631);
not I_73652 (I1255689,I3570);
DFFARX1 I_73653 (I316997,I3563,I1255689,I1255715,);
nand I_73654 (I1255723,I1255715,I317000);
DFFARX1 I_73655 (I316994,I3563,I1255689,I1255749,);
DFFARX1 I_73656 (I1255749,I3563,I1255689,I1255766,);
not I_73657 (I1255681,I1255766);
not I_73658 (I1255788,I317003);
nor I_73659 (I1255805,I317003,I316988);
not I_73660 (I1255822,I317012);
nand I_73661 (I1255839,I1255788,I1255822);
nor I_73662 (I1255856,I317012,I317003);
and I_73663 (I1255660,I1255856,I1255723);
not I_73664 (I1255887,I316991);
nand I_73665 (I1255904,I1255887,I317009);
nor I_73666 (I1255921,I316991,I316985);
not I_73667 (I1255938,I1255921);
nand I_73668 (I1255663,I1255805,I1255938);
DFFARX1 I_73669 (I1255921,I3563,I1255689,I1255678,);
nor I_73670 (I1255983,I317006,I317012);
nor I_73671 (I1256000,I1255983,I316988);
and I_73672 (I1256017,I1256000,I1255904);
DFFARX1 I_73673 (I1256017,I3563,I1255689,I1255675,);
nor I_73674 (I1255672,I1255983,I1255839);
or I_73675 (I1255669,I1255921,I1255983);
nor I_73676 (I1256076,I317006,I316985);
DFFARX1 I_73677 (I1256076,I3563,I1255689,I1256102,);
not I_73678 (I1256110,I1256102);
nand I_73679 (I1256127,I1256110,I1255788);
nor I_73680 (I1256144,I1256127,I316988);
DFFARX1 I_73681 (I1256144,I3563,I1255689,I1255657,);
nor I_73682 (I1256175,I1256110,I1255839);
nor I_73683 (I1255666,I1255983,I1256175);
not I_73684 (I1256233,I3570);
DFFARX1 I_73685 (I182167,I3563,I1256233,I1256259,);
nand I_73686 (I1256267,I1256259,I182182);
DFFARX1 I_73687 (I182179,I3563,I1256233,I1256293,);
DFFARX1 I_73688 (I1256293,I3563,I1256233,I1256310,);
not I_73689 (I1256225,I1256310);
not I_73690 (I1256332,I182158);
nor I_73691 (I1256349,I182158,I182164);
not I_73692 (I1256366,I182170);
nand I_73693 (I1256383,I1256332,I1256366);
nor I_73694 (I1256400,I182170,I182158);
and I_73695 (I1256204,I1256400,I1256267);
not I_73696 (I1256431,I182176);
nand I_73697 (I1256448,I1256431,I182158);
nor I_73698 (I1256465,I182176,I182161);
not I_73699 (I1256482,I1256465);
nand I_73700 (I1256207,I1256349,I1256482);
DFFARX1 I_73701 (I1256465,I3563,I1256233,I1256222,);
nor I_73702 (I1256527,I182161,I182170);
nor I_73703 (I1256544,I1256527,I182164);
and I_73704 (I1256561,I1256544,I1256448);
DFFARX1 I_73705 (I1256561,I3563,I1256233,I1256219,);
nor I_73706 (I1256216,I1256527,I1256383);
or I_73707 (I1256213,I1256465,I1256527);
nor I_73708 (I1256620,I182161,I182173);
DFFARX1 I_73709 (I1256620,I3563,I1256233,I1256646,);
not I_73710 (I1256654,I1256646);
nand I_73711 (I1256671,I1256654,I1256332);
nor I_73712 (I1256688,I1256671,I182164);
DFFARX1 I_73713 (I1256688,I3563,I1256233,I1256201,);
nor I_73714 (I1256719,I1256654,I1256383);
nor I_73715 (I1256210,I1256527,I1256719);
not I_73716 (I1256777,I3570);
DFFARX1 I_73717 (I22928,I3563,I1256777,I1256803,);
nand I_73718 (I1256811,I1256803,I22922);
DFFARX1 I_73719 (I22943,I3563,I1256777,I1256837,);
DFFARX1 I_73720 (I1256837,I3563,I1256777,I1256854,);
not I_73721 (I1256769,I1256854);
not I_73722 (I1256876,I22931);
nor I_73723 (I1256893,I22931,I22940);
not I_73724 (I1256910,I22919);
nand I_73725 (I1256927,I1256876,I1256910);
nor I_73726 (I1256944,I22919,I22931);
and I_73727 (I1256748,I1256944,I1256811);
not I_73728 (I1256975,I22937);
nand I_73729 (I1256992,I1256975,I22925);
nor I_73730 (I1257009,I22937,I22919);
not I_73731 (I1257026,I1257009);
nand I_73732 (I1256751,I1256893,I1257026);
DFFARX1 I_73733 (I1257009,I3563,I1256777,I1256766,);
nor I_73734 (I1257071,I22922,I22919);
nor I_73735 (I1257088,I1257071,I22940);
and I_73736 (I1257105,I1257088,I1256992);
DFFARX1 I_73737 (I1257105,I3563,I1256777,I1256763,);
nor I_73738 (I1256760,I1257071,I1256927);
or I_73739 (I1256757,I1257009,I1257071);
nor I_73740 (I1257164,I22922,I22934);
DFFARX1 I_73741 (I1257164,I3563,I1256777,I1257190,);
not I_73742 (I1257198,I1257190);
nand I_73743 (I1257215,I1257198,I1256876);
nor I_73744 (I1257232,I1257215,I22940);
DFFARX1 I_73745 (I1257232,I3563,I1256777,I1256745,);
nor I_73746 (I1257263,I1257198,I1256927);
nor I_73747 (I1256754,I1257071,I1257263);
not I_73748 (I1257321,I3570);
DFFARX1 I_73749 (I1373800,I3563,I1257321,I1257347,);
nand I_73750 (I1257355,I1257347,I1373785);
DFFARX1 I_73751 (I1373779,I3563,I1257321,I1257381,);
DFFARX1 I_73752 (I1257381,I3563,I1257321,I1257398,);
not I_73753 (I1257313,I1257398);
not I_73754 (I1257420,I1373773);
nor I_73755 (I1257437,I1373773,I1373794);
not I_73756 (I1257454,I1373782);
nand I_73757 (I1257471,I1257420,I1257454);
nor I_73758 (I1257488,I1373782,I1373773);
and I_73759 (I1257292,I1257488,I1257355);
not I_73760 (I1257519,I1373791);
nand I_73761 (I1257536,I1257519,I1373797);
nor I_73762 (I1257553,I1373791,I1373788);
not I_73763 (I1257570,I1257553);
nand I_73764 (I1257295,I1257437,I1257570);
DFFARX1 I_73765 (I1257553,I3563,I1257321,I1257310,);
nor I_73766 (I1257615,I1373776,I1373782);
nor I_73767 (I1257632,I1257615,I1373794);
and I_73768 (I1257649,I1257632,I1257536);
DFFARX1 I_73769 (I1257649,I3563,I1257321,I1257307,);
nor I_73770 (I1257304,I1257615,I1257471);
or I_73771 (I1257301,I1257553,I1257615);
nor I_73772 (I1257708,I1373776,I1373773);
DFFARX1 I_73773 (I1257708,I3563,I1257321,I1257734,);
not I_73774 (I1257742,I1257734);
nand I_73775 (I1257759,I1257742,I1257420);
nor I_73776 (I1257776,I1257759,I1373794);
DFFARX1 I_73777 (I1257776,I3563,I1257321,I1257289,);
nor I_73778 (I1257807,I1257742,I1257471);
nor I_73779 (I1257298,I1257615,I1257807);
not I_73780 (I1257865,I3570);
DFFARX1 I_73781 (I1060141,I3563,I1257865,I1257891,);
nand I_73782 (I1257899,I1257891,I1060129);
DFFARX1 I_73783 (I1060123,I3563,I1257865,I1257925,);
DFFARX1 I_73784 (I1257925,I3563,I1257865,I1257942,);
not I_73785 (I1257857,I1257942);
not I_73786 (I1257964,I1060123);
nor I_73787 (I1257981,I1060123,I1060135);
not I_73788 (I1257998,I1060132);
nand I_73789 (I1258015,I1257964,I1257998);
nor I_73790 (I1258032,I1060132,I1060123);
and I_73791 (I1257836,I1258032,I1257899);
not I_73792 (I1258063,I1060126);
nand I_73793 (I1258080,I1258063,I1060138);
nor I_73794 (I1258097,I1060126,I1060144);
not I_73795 (I1258114,I1258097);
nand I_73796 (I1257839,I1257981,I1258114);
DFFARX1 I_73797 (I1258097,I3563,I1257865,I1257854,);
nor I_73798 (I1258159,I1060129,I1060132);
nor I_73799 (I1258176,I1258159,I1060135);
and I_73800 (I1258193,I1258176,I1258080);
DFFARX1 I_73801 (I1258193,I3563,I1257865,I1257851,);
nor I_73802 (I1257848,I1258159,I1258015);
or I_73803 (I1257845,I1258097,I1258159);
nor I_73804 (I1258252,I1060129,I1060126);
DFFARX1 I_73805 (I1258252,I3563,I1257865,I1258278,);
not I_73806 (I1258286,I1258278);
nand I_73807 (I1258303,I1258286,I1257964);
nor I_73808 (I1258320,I1258303,I1060135);
DFFARX1 I_73809 (I1258320,I3563,I1257865,I1257833,);
nor I_73810 (I1258351,I1258286,I1258015);
nor I_73811 (I1257842,I1258159,I1258351);
not I_73812 (I1258409,I3570);
DFFARX1 I_73813 (I131502,I3563,I1258409,I1258435,);
nand I_73814 (I1258443,I1258435,I131484);
DFFARX1 I_73815 (I131481,I3563,I1258409,I1258469,);
DFFARX1 I_73816 (I1258469,I3563,I1258409,I1258486,);
not I_73817 (I1258401,I1258486);
not I_73818 (I1258508,I131499);
nor I_73819 (I1258525,I131499,I131493);
not I_73820 (I1258542,I131481);
nand I_73821 (I1258559,I1258508,I1258542);
nor I_73822 (I1258576,I131481,I131499);
and I_73823 (I1258380,I1258576,I1258443);
not I_73824 (I1258607,I131490);
nand I_73825 (I1258624,I1258607,I131496);
nor I_73826 (I1258641,I131490,I131484);
not I_73827 (I1258658,I1258641);
nand I_73828 (I1258383,I1258525,I1258658);
DFFARX1 I_73829 (I1258641,I3563,I1258409,I1258398,);
nor I_73830 (I1258703,I131487,I131481);
nor I_73831 (I1258720,I1258703,I131493);
and I_73832 (I1258737,I1258720,I1258624);
DFFARX1 I_73833 (I1258737,I3563,I1258409,I1258395,);
nor I_73834 (I1258392,I1258703,I1258559);
or I_73835 (I1258389,I1258641,I1258703);
nor I_73836 (I1258796,I131487,I131505);
DFFARX1 I_73837 (I1258796,I3563,I1258409,I1258822,);
not I_73838 (I1258830,I1258822);
nand I_73839 (I1258847,I1258830,I1258508);
nor I_73840 (I1258864,I1258847,I131493);
DFFARX1 I_73841 (I1258864,I3563,I1258409,I1258377,);
nor I_73842 (I1258895,I1258830,I1258559);
nor I_73843 (I1258386,I1258703,I1258895);
not I_73844 (I1258953,I3570);
DFFARX1 I_73845 (I560221,I3563,I1258953,I1258979,);
nand I_73846 (I1258987,I1258979,I560245);
DFFARX1 I_73847 (I560224,I3563,I1258953,I1259013,);
DFFARX1 I_73848 (I1259013,I3563,I1258953,I1259030,);
not I_73849 (I1258945,I1259030);
not I_73850 (I1259052,I560227);
nor I_73851 (I1259069,I560227,I560242);
not I_73852 (I1259086,I560233);
nand I_73853 (I1259103,I1259052,I1259086);
nor I_73854 (I1259120,I560233,I560227);
and I_73855 (I1258924,I1259120,I1258987);
not I_73856 (I1259151,I560230);
nand I_73857 (I1259168,I1259151,I560224);
nor I_73858 (I1259185,I560230,I560239);
not I_73859 (I1259202,I1259185);
nand I_73860 (I1258927,I1259069,I1259202);
DFFARX1 I_73861 (I1259185,I3563,I1258953,I1258942,);
nor I_73862 (I1259247,I560236,I560233);
nor I_73863 (I1259264,I1259247,I560242);
and I_73864 (I1259281,I1259264,I1259168);
DFFARX1 I_73865 (I1259281,I3563,I1258953,I1258939,);
nor I_73866 (I1258936,I1259247,I1259103);
or I_73867 (I1258933,I1259185,I1259247);
nor I_73868 (I1259340,I560236,I560221);
DFFARX1 I_73869 (I1259340,I3563,I1258953,I1259366,);
not I_73870 (I1259374,I1259366);
nand I_73871 (I1259391,I1259374,I1259052);
nor I_73872 (I1259408,I1259391,I560242);
DFFARX1 I_73873 (I1259408,I3563,I1258953,I1258921,);
nor I_73874 (I1259439,I1259374,I1259103);
nor I_73875 (I1258930,I1259247,I1259439);
not I_73876 (I1259497,I3570);
DFFARX1 I_73877 (I1186967,I3563,I1259497,I1259523,);
nand I_73878 (I1259531,I1259523,I1186946);
DFFARX1 I_73879 (I1186943,I3563,I1259497,I1259557,);
DFFARX1 I_73880 (I1259557,I3563,I1259497,I1259574,);
not I_73881 (I1259489,I1259574);
not I_73882 (I1259596,I1186955);
nor I_73883 (I1259613,I1186955,I1186964);
not I_73884 (I1259630,I1186952);
nand I_73885 (I1259647,I1259596,I1259630);
nor I_73886 (I1259664,I1186952,I1186955);
and I_73887 (I1259468,I1259664,I1259531);
not I_73888 (I1259695,I1186961);
nand I_73889 (I1259712,I1259695,I1186958);
nor I_73890 (I1259729,I1186961,I1186943);
not I_73891 (I1259746,I1259729);
nand I_73892 (I1259471,I1259613,I1259746);
DFFARX1 I_73893 (I1259729,I3563,I1259497,I1259486,);
nor I_73894 (I1259791,I1186946,I1186952);
nor I_73895 (I1259808,I1259791,I1186964);
and I_73896 (I1259825,I1259808,I1259712);
DFFARX1 I_73897 (I1259825,I3563,I1259497,I1259483,);
nor I_73898 (I1259480,I1259791,I1259647);
or I_73899 (I1259477,I1259729,I1259791);
nor I_73900 (I1259884,I1186946,I1186949);
DFFARX1 I_73901 (I1259884,I3563,I1259497,I1259910,);
not I_73902 (I1259918,I1259910);
nand I_73903 (I1259935,I1259918,I1259596);
nor I_73904 (I1259952,I1259935,I1186964);
DFFARX1 I_73905 (I1259952,I3563,I1259497,I1259465,);
nor I_73906 (I1259983,I1259918,I1259647);
nor I_73907 (I1259474,I1259791,I1259983);
not I_73908 (I1260041,I3570);
DFFARX1 I_73909 (I823710,I3563,I1260041,I1260067,);
nand I_73910 (I1260075,I1260067,I823704);
DFFARX1 I_73911 (I823707,I3563,I1260041,I1260101,);
DFFARX1 I_73912 (I1260101,I3563,I1260041,I1260118,);
not I_73913 (I1260033,I1260118);
not I_73914 (I1260140,I823713);
nor I_73915 (I1260157,I823713,I823707);
not I_73916 (I1260174,I823716);
nand I_73917 (I1260191,I1260140,I1260174);
nor I_73918 (I1260208,I823716,I823713);
and I_73919 (I1260012,I1260208,I1260075);
not I_73920 (I1260239,I823725);
nand I_73921 (I1260256,I1260239,I823719);
nor I_73922 (I1260273,I823725,I823722);
not I_73923 (I1260290,I1260273);
nand I_73924 (I1260015,I1260157,I1260290);
DFFARX1 I_73925 (I1260273,I3563,I1260041,I1260030,);
nor I_73926 (I1260335,I823704,I823716);
nor I_73927 (I1260352,I1260335,I823707);
and I_73928 (I1260369,I1260352,I1260256);
DFFARX1 I_73929 (I1260369,I3563,I1260041,I1260027,);
nor I_73930 (I1260024,I1260335,I1260191);
or I_73931 (I1260021,I1260273,I1260335);
nor I_73932 (I1260428,I823704,I823710);
DFFARX1 I_73933 (I1260428,I3563,I1260041,I1260454,);
not I_73934 (I1260462,I1260454);
nand I_73935 (I1260479,I1260462,I1260140);
nor I_73936 (I1260496,I1260479,I823707);
DFFARX1 I_73937 (I1260496,I3563,I1260041,I1260009,);
nor I_73938 (I1260527,I1260462,I1260191);
nor I_73939 (I1260018,I1260335,I1260527);
not I_73940 (I1260585,I3570);
DFFARX1 I_73941 (I1208931,I3563,I1260585,I1260611,);
nand I_73942 (I1260619,I1260611,I1208910);
DFFARX1 I_73943 (I1208907,I3563,I1260585,I1260645,);
DFFARX1 I_73944 (I1260645,I3563,I1260585,I1260662,);
not I_73945 (I1260577,I1260662);
not I_73946 (I1260684,I1208919);
nor I_73947 (I1260701,I1208919,I1208928);
not I_73948 (I1260718,I1208916);
nand I_73949 (I1260735,I1260684,I1260718);
nor I_73950 (I1260752,I1208916,I1208919);
and I_73951 (I1260556,I1260752,I1260619);
not I_73952 (I1260783,I1208925);
nand I_73953 (I1260800,I1260783,I1208922);
nor I_73954 (I1260817,I1208925,I1208907);
not I_73955 (I1260834,I1260817);
nand I_73956 (I1260559,I1260701,I1260834);
DFFARX1 I_73957 (I1260817,I3563,I1260585,I1260574,);
nor I_73958 (I1260879,I1208910,I1208916);
nor I_73959 (I1260896,I1260879,I1208928);
and I_73960 (I1260913,I1260896,I1260800);
DFFARX1 I_73961 (I1260913,I3563,I1260585,I1260571,);
nor I_73962 (I1260568,I1260879,I1260735);
or I_73963 (I1260565,I1260817,I1260879);
nor I_73964 (I1260972,I1208910,I1208913);
DFFARX1 I_73965 (I1260972,I3563,I1260585,I1260998,);
not I_73966 (I1261006,I1260998);
nand I_73967 (I1261023,I1261006,I1260684);
nor I_73968 (I1261040,I1261023,I1208928);
DFFARX1 I_73969 (I1261040,I3563,I1260585,I1260553,);
nor I_73970 (I1261071,I1261006,I1260735);
nor I_73971 (I1260562,I1260879,I1261071);
not I_73972 (I1261129,I3570);
DFFARX1 I_73973 (I311200,I3563,I1261129,I1261155,);
nand I_73974 (I1261163,I1261155,I311203);
DFFARX1 I_73975 (I311197,I3563,I1261129,I1261189,);
DFFARX1 I_73976 (I1261189,I3563,I1261129,I1261206,);
not I_73977 (I1261121,I1261206);
not I_73978 (I1261228,I311206);
nor I_73979 (I1261245,I311206,I311191);
not I_73980 (I1261262,I311215);
nand I_73981 (I1261279,I1261228,I1261262);
nor I_73982 (I1261296,I311215,I311206);
and I_73983 (I1261100,I1261296,I1261163);
not I_73984 (I1261327,I311194);
nand I_73985 (I1261344,I1261327,I311212);
nor I_73986 (I1261361,I311194,I311188);
not I_73987 (I1261378,I1261361);
nand I_73988 (I1261103,I1261245,I1261378);
DFFARX1 I_73989 (I1261361,I3563,I1261129,I1261118,);
nor I_73990 (I1261423,I311209,I311215);
nor I_73991 (I1261440,I1261423,I311191);
and I_73992 (I1261457,I1261440,I1261344);
DFFARX1 I_73993 (I1261457,I3563,I1261129,I1261115,);
nor I_73994 (I1261112,I1261423,I1261279);
or I_73995 (I1261109,I1261361,I1261423);
nor I_73996 (I1261516,I311209,I311188);
DFFARX1 I_73997 (I1261516,I3563,I1261129,I1261542,);
not I_73998 (I1261550,I1261542);
nand I_73999 (I1261567,I1261550,I1261228);
nor I_74000 (I1261584,I1261567,I311191);
DFFARX1 I_74001 (I1261584,I3563,I1261129,I1261097,);
nor I_74002 (I1261615,I1261550,I1261279);
nor I_74003 (I1261106,I1261423,I1261615);
not I_74004 (I1261673,I3570);
DFFARX1 I_74005 (I74059,I3563,I1261673,I1261699,);
nand I_74006 (I1261707,I1261699,I74041);
DFFARX1 I_74007 (I74038,I3563,I1261673,I1261733,);
DFFARX1 I_74008 (I1261733,I3563,I1261673,I1261750,);
not I_74009 (I1261665,I1261750);
not I_74010 (I1261772,I74056);
nor I_74011 (I1261789,I74056,I74050);
not I_74012 (I1261806,I74038);
nand I_74013 (I1261823,I1261772,I1261806);
nor I_74014 (I1261840,I74038,I74056);
and I_74015 (I1261644,I1261840,I1261707);
not I_74016 (I1261871,I74047);
nand I_74017 (I1261888,I1261871,I74053);
nor I_74018 (I1261905,I74047,I74041);
not I_74019 (I1261922,I1261905);
nand I_74020 (I1261647,I1261789,I1261922);
DFFARX1 I_74021 (I1261905,I3563,I1261673,I1261662,);
nor I_74022 (I1261967,I74044,I74038);
nor I_74023 (I1261984,I1261967,I74050);
and I_74024 (I1262001,I1261984,I1261888);
DFFARX1 I_74025 (I1262001,I3563,I1261673,I1261659,);
nor I_74026 (I1261656,I1261967,I1261823);
or I_74027 (I1261653,I1261905,I1261967);
nor I_74028 (I1262060,I74044,I74062);
DFFARX1 I_74029 (I1262060,I3563,I1261673,I1262086,);
not I_74030 (I1262094,I1262086);
nand I_74031 (I1262111,I1262094,I1261772);
nor I_74032 (I1262128,I1262111,I74050);
DFFARX1 I_74033 (I1262128,I3563,I1261673,I1261641,);
nor I_74034 (I1262159,I1262094,I1261823);
nor I_74035 (I1261650,I1261967,I1262159);
not I_74036 (I1262217,I3570);
DFFARX1 I_74037 (I575691,I3563,I1262217,I1262243,);
nand I_74038 (I1262251,I1262243,I575715);
DFFARX1 I_74039 (I575694,I3563,I1262217,I1262277,);
DFFARX1 I_74040 (I1262277,I3563,I1262217,I1262294,);
not I_74041 (I1262209,I1262294);
not I_74042 (I1262316,I575697);
nor I_74043 (I1262333,I575697,I575712);
not I_74044 (I1262350,I575703);
nand I_74045 (I1262367,I1262316,I1262350);
nor I_74046 (I1262384,I575703,I575697);
and I_74047 (I1262188,I1262384,I1262251);
not I_74048 (I1262415,I575700);
nand I_74049 (I1262432,I1262415,I575694);
nor I_74050 (I1262449,I575700,I575709);
not I_74051 (I1262466,I1262449);
nand I_74052 (I1262191,I1262333,I1262466);
DFFARX1 I_74053 (I1262449,I3563,I1262217,I1262206,);
nor I_74054 (I1262511,I575706,I575703);
nor I_74055 (I1262528,I1262511,I575712);
and I_74056 (I1262545,I1262528,I1262432);
DFFARX1 I_74057 (I1262545,I3563,I1262217,I1262203,);
nor I_74058 (I1262200,I1262511,I1262367);
or I_74059 (I1262197,I1262449,I1262511);
nor I_74060 (I1262604,I575706,I575691);
DFFARX1 I_74061 (I1262604,I3563,I1262217,I1262630,);
not I_74062 (I1262638,I1262630);
nand I_74063 (I1262655,I1262638,I1262316);
nor I_74064 (I1262672,I1262655,I575712);
DFFARX1 I_74065 (I1262672,I3563,I1262217,I1262185,);
nor I_74066 (I1262703,I1262638,I1262367);
nor I_74067 (I1262194,I1262511,I1262703);
not I_74068 (I1262761,I3570);
DFFARX1 I_74069 (I1108359,I3563,I1262761,I1262787,);
nand I_74070 (I1262795,I1262787,I1108338);
DFFARX1 I_74071 (I1108335,I3563,I1262761,I1262821,);
DFFARX1 I_74072 (I1262821,I3563,I1262761,I1262838,);
not I_74073 (I1262753,I1262838);
not I_74074 (I1262860,I1108347);
nor I_74075 (I1262877,I1108347,I1108356);
not I_74076 (I1262894,I1108344);
nand I_74077 (I1262911,I1262860,I1262894);
nor I_74078 (I1262928,I1108344,I1108347);
and I_74079 (I1262732,I1262928,I1262795);
not I_74080 (I1262959,I1108353);
nand I_74081 (I1262976,I1262959,I1108350);
nor I_74082 (I1262993,I1108353,I1108335);
not I_74083 (I1263010,I1262993);
nand I_74084 (I1262735,I1262877,I1263010);
DFFARX1 I_74085 (I1262993,I3563,I1262761,I1262750,);
nor I_74086 (I1263055,I1108338,I1108344);
nor I_74087 (I1263072,I1263055,I1108356);
and I_74088 (I1263089,I1263072,I1262976);
DFFARX1 I_74089 (I1263089,I3563,I1262761,I1262747,);
nor I_74090 (I1262744,I1263055,I1262911);
or I_74091 (I1262741,I1262993,I1263055);
nor I_74092 (I1263148,I1108338,I1108341);
DFFARX1 I_74093 (I1263148,I3563,I1262761,I1263174,);
not I_74094 (I1263182,I1263174);
nand I_74095 (I1263199,I1263182,I1262860);
nor I_74096 (I1263216,I1263199,I1108356);
DFFARX1 I_74097 (I1263216,I3563,I1262761,I1262729,);
nor I_74098 (I1263247,I1263182,I1262911);
nor I_74099 (I1262738,I1263055,I1263247);
not I_74100 (I1263305,I3570);
DFFARX1 I_74101 (I1113561,I3563,I1263305,I1263331,);
nand I_74102 (I1263339,I1263331,I1113540);
DFFARX1 I_74103 (I1113537,I3563,I1263305,I1263365,);
DFFARX1 I_74104 (I1263365,I3563,I1263305,I1263382,);
not I_74105 (I1263297,I1263382);
not I_74106 (I1263404,I1113549);
nor I_74107 (I1263421,I1113549,I1113558);
not I_74108 (I1263438,I1113546);
nand I_74109 (I1263455,I1263404,I1263438);
nor I_74110 (I1263472,I1113546,I1113549);
and I_74111 (I1263276,I1263472,I1263339);
not I_74112 (I1263503,I1113555);
nand I_74113 (I1263520,I1263503,I1113552);
nor I_74114 (I1263537,I1113555,I1113537);
not I_74115 (I1263554,I1263537);
nand I_74116 (I1263279,I1263421,I1263554);
DFFARX1 I_74117 (I1263537,I3563,I1263305,I1263294,);
nor I_74118 (I1263599,I1113540,I1113546);
nor I_74119 (I1263616,I1263599,I1113558);
and I_74120 (I1263633,I1263616,I1263520);
DFFARX1 I_74121 (I1263633,I3563,I1263305,I1263291,);
nor I_74122 (I1263288,I1263599,I1263455);
or I_74123 (I1263285,I1263537,I1263599);
nor I_74124 (I1263692,I1113540,I1113543);
DFFARX1 I_74125 (I1263692,I3563,I1263305,I1263718,);
not I_74126 (I1263726,I1263718);
nand I_74127 (I1263743,I1263726,I1263404);
nor I_74128 (I1263760,I1263743,I1113558);
DFFARX1 I_74129 (I1263760,I3563,I1263305,I1263273,);
nor I_74130 (I1263791,I1263726,I1263455);
nor I_74131 (I1263282,I1263599,I1263791);
not I_74132 (I1263849,I3570);
DFFARX1 I_74133 (I524698,I3563,I1263849,I1263875,);
nand I_74134 (I1263883,I1263875,I524695);
DFFARX1 I_74135 (I524674,I3563,I1263849,I1263909,);
DFFARX1 I_74136 (I1263909,I3563,I1263849,I1263926,);
not I_74137 (I1263841,I1263926);
not I_74138 (I1263948,I524689);
nor I_74139 (I1263965,I524689,I524692);
not I_74140 (I1263982,I524683);
nand I_74141 (I1263999,I1263948,I1263982);
nor I_74142 (I1264016,I524683,I524689);
and I_74143 (I1263820,I1264016,I1263883);
not I_74144 (I1264047,I524680);
nand I_74145 (I1264064,I1264047,I524701);
nor I_74146 (I1264081,I524680,I524677);
not I_74147 (I1264098,I1264081);
nand I_74148 (I1263823,I1263965,I1264098);
DFFARX1 I_74149 (I1264081,I3563,I1263849,I1263838,);
nor I_74150 (I1264143,I524686,I524683);
nor I_74151 (I1264160,I1264143,I524692);
and I_74152 (I1264177,I1264160,I1264064);
DFFARX1 I_74153 (I1264177,I3563,I1263849,I1263835,);
nor I_74154 (I1263832,I1264143,I1263999);
or I_74155 (I1263829,I1264081,I1264143);
nor I_74156 (I1264236,I524686,I524674);
DFFARX1 I_74157 (I1264236,I3563,I1263849,I1264262,);
not I_74158 (I1264270,I1264262);
nand I_74159 (I1264287,I1264270,I1263948);
nor I_74160 (I1264304,I1264287,I524692);
DFFARX1 I_74161 (I1264304,I3563,I1263849,I1263817,);
nor I_74162 (I1264335,I1264270,I1263999);
nor I_74163 (I1263826,I1264143,I1264335);
not I_74164 (I1264393,I3570);
DFFARX1 I_74165 (I804072,I3563,I1264393,I1264419,);
nand I_74166 (I1264427,I1264419,I804087);
DFFARX1 I_74167 (I804081,I3563,I1264393,I1264453,);
DFFARX1 I_74168 (I1264453,I3563,I1264393,I1264470,);
not I_74169 (I1264385,I1264470);
not I_74170 (I1264492,I804084);
nor I_74171 (I1264509,I804084,I804090);
not I_74172 (I1264526,I804072);
nand I_74173 (I1264543,I1264492,I1264526);
nor I_74174 (I1264560,I804072,I804084);
and I_74175 (I1264364,I1264560,I1264427);
not I_74176 (I1264591,I804069);
nand I_74177 (I1264608,I1264591,I804075);
nor I_74178 (I1264625,I804069,I804069);
not I_74179 (I1264642,I1264625);
nand I_74180 (I1264367,I1264509,I1264642);
DFFARX1 I_74181 (I1264625,I3563,I1264393,I1264382,);
nor I_74182 (I1264687,I804078,I804072);
nor I_74183 (I1264704,I1264687,I804090);
and I_74184 (I1264721,I1264704,I1264608);
DFFARX1 I_74185 (I1264721,I3563,I1264393,I1264379,);
nor I_74186 (I1264376,I1264687,I1264543);
or I_74187 (I1264373,I1264625,I1264687);
nor I_74188 (I1264780,I804078,I804093);
DFFARX1 I_74189 (I1264780,I3563,I1264393,I1264806,);
not I_74190 (I1264814,I1264806);
nand I_74191 (I1264831,I1264814,I1264492);
nor I_74192 (I1264848,I1264831,I804090);
DFFARX1 I_74193 (I1264848,I3563,I1264393,I1264361,);
nor I_74194 (I1264879,I1264814,I1264543);
nor I_74195 (I1264370,I1264687,I1264879);
not I_74196 (I1264937,I3570);
DFFARX1 I_74197 (I983997,I3563,I1264937,I1264963,);
nand I_74198 (I1264971,I1264963,I983997);
DFFARX1 I_74199 (I984009,I3563,I1264937,I1264997,);
DFFARX1 I_74200 (I1264997,I3563,I1264937,I1265014,);
not I_74201 (I1264929,I1265014);
not I_74202 (I1265036,I984003);
nor I_74203 (I1265053,I984003,I984024);
not I_74204 (I1265070,I984012);
nand I_74205 (I1265087,I1265036,I1265070);
nor I_74206 (I1265104,I984012,I984003);
and I_74207 (I1264908,I1265104,I1264971);
not I_74208 (I1265135,I984006);
nand I_74209 (I1265152,I1265135,I984021);
nor I_74210 (I1265169,I984006,I984015);
not I_74211 (I1265186,I1265169);
nand I_74212 (I1264911,I1265053,I1265186);
DFFARX1 I_74213 (I1265169,I3563,I1264937,I1264926,);
nor I_74214 (I1265231,I984018,I984012);
nor I_74215 (I1265248,I1265231,I984024);
and I_74216 (I1265265,I1265248,I1265152);
DFFARX1 I_74217 (I1265265,I3563,I1264937,I1264923,);
nor I_74218 (I1264920,I1265231,I1265087);
or I_74219 (I1264917,I1265169,I1265231);
nor I_74220 (I1265324,I984018,I984000);
DFFARX1 I_74221 (I1265324,I3563,I1264937,I1265350,);
not I_74222 (I1265358,I1265350);
nand I_74223 (I1265375,I1265358,I1265036);
nor I_74224 (I1265392,I1265375,I984024);
DFFARX1 I_74225 (I1265392,I3563,I1264937,I1264905,);
nor I_74226 (I1265423,I1265358,I1265087);
nor I_74227 (I1264914,I1265231,I1265423);
not I_74228 (I1265481,I3570);
DFFARX1 I_74229 (I1142461,I3563,I1265481,I1265507,);
nand I_74230 (I1265515,I1265507,I1142440);
DFFARX1 I_74231 (I1142437,I3563,I1265481,I1265541,);
DFFARX1 I_74232 (I1265541,I3563,I1265481,I1265558,);
not I_74233 (I1265473,I1265558);
not I_74234 (I1265580,I1142449);
nor I_74235 (I1265597,I1142449,I1142458);
not I_74236 (I1265614,I1142446);
nand I_74237 (I1265631,I1265580,I1265614);
nor I_74238 (I1265648,I1142446,I1142449);
and I_74239 (I1265452,I1265648,I1265515);
not I_74240 (I1265679,I1142455);
nand I_74241 (I1265696,I1265679,I1142452);
nor I_74242 (I1265713,I1142455,I1142437);
not I_74243 (I1265730,I1265713);
nand I_74244 (I1265455,I1265597,I1265730);
DFFARX1 I_74245 (I1265713,I3563,I1265481,I1265470,);
nor I_74246 (I1265775,I1142440,I1142446);
nor I_74247 (I1265792,I1265775,I1142458);
and I_74248 (I1265809,I1265792,I1265696);
DFFARX1 I_74249 (I1265809,I3563,I1265481,I1265467,);
nor I_74250 (I1265464,I1265775,I1265631);
or I_74251 (I1265461,I1265713,I1265775);
nor I_74252 (I1265868,I1142440,I1142443);
DFFARX1 I_74253 (I1265868,I3563,I1265481,I1265894,);
not I_74254 (I1265902,I1265894);
nand I_74255 (I1265919,I1265902,I1265580);
nor I_74256 (I1265936,I1265919,I1142458);
DFFARX1 I_74257 (I1265936,I3563,I1265481,I1265449,);
nor I_74258 (I1265967,I1265902,I1265631);
nor I_74259 (I1265458,I1265775,I1265967);
not I_74260 (I1266025,I3570);
DFFARX1 I_74261 (I55075,I3563,I1266025,I1266051,);
nand I_74262 (I1266059,I1266051,I55069);
DFFARX1 I_74263 (I55090,I3563,I1266025,I1266085,);
DFFARX1 I_74264 (I1266085,I3563,I1266025,I1266102,);
not I_74265 (I1266017,I1266102);
not I_74266 (I1266124,I55078);
nor I_74267 (I1266141,I55078,I55087);
not I_74268 (I1266158,I55066);
nand I_74269 (I1266175,I1266124,I1266158);
nor I_74270 (I1266192,I55066,I55078);
and I_74271 (I1265996,I1266192,I1266059);
not I_74272 (I1266223,I55084);
nand I_74273 (I1266240,I1266223,I55072);
nor I_74274 (I1266257,I55084,I55066);
not I_74275 (I1266274,I1266257);
nand I_74276 (I1265999,I1266141,I1266274);
DFFARX1 I_74277 (I1266257,I3563,I1266025,I1266014,);
nor I_74278 (I1266319,I55069,I55066);
nor I_74279 (I1266336,I1266319,I55087);
and I_74280 (I1266353,I1266336,I1266240);
DFFARX1 I_74281 (I1266353,I3563,I1266025,I1266011,);
nor I_74282 (I1266008,I1266319,I1266175);
or I_74283 (I1266005,I1266257,I1266319);
nor I_74284 (I1266412,I55069,I55081);
DFFARX1 I_74285 (I1266412,I3563,I1266025,I1266438,);
not I_74286 (I1266446,I1266438);
nand I_74287 (I1266463,I1266446,I1266124);
nor I_74288 (I1266480,I1266463,I55087);
DFFARX1 I_74289 (I1266480,I3563,I1266025,I1265993,);
nor I_74290 (I1266511,I1266446,I1266175);
nor I_74291 (I1266002,I1266319,I1266511);
not I_74292 (I1266569,I3570);
DFFARX1 I_74293 (I1027279,I3563,I1266569,I1266595,);
nand I_74294 (I1266603,I1266595,I1027279);
DFFARX1 I_74295 (I1027291,I3563,I1266569,I1266629,);
DFFARX1 I_74296 (I1266629,I3563,I1266569,I1266646,);
not I_74297 (I1266561,I1266646);
not I_74298 (I1266668,I1027285);
nor I_74299 (I1266685,I1027285,I1027306);
not I_74300 (I1266702,I1027294);
nand I_74301 (I1266719,I1266668,I1266702);
nor I_74302 (I1266736,I1027294,I1027285);
and I_74303 (I1266540,I1266736,I1266603);
not I_74304 (I1266767,I1027288);
nand I_74305 (I1266784,I1266767,I1027303);
nor I_74306 (I1266801,I1027288,I1027297);
not I_74307 (I1266818,I1266801);
nand I_74308 (I1266543,I1266685,I1266818);
DFFARX1 I_74309 (I1266801,I3563,I1266569,I1266558,);
nor I_74310 (I1266863,I1027300,I1027294);
nor I_74311 (I1266880,I1266863,I1027306);
and I_74312 (I1266897,I1266880,I1266784);
DFFARX1 I_74313 (I1266897,I3563,I1266569,I1266555,);
nor I_74314 (I1266552,I1266863,I1266719);
or I_74315 (I1266549,I1266801,I1266863);
nor I_74316 (I1266956,I1027300,I1027282);
DFFARX1 I_74317 (I1266956,I3563,I1266569,I1266982,);
not I_74318 (I1266990,I1266982);
nand I_74319 (I1267007,I1266990,I1266668);
nor I_74320 (I1267024,I1267007,I1027306);
DFFARX1 I_74321 (I1267024,I3563,I1266569,I1266537,);
nor I_74322 (I1267055,I1266990,I1266719);
nor I_74323 (I1266546,I1266863,I1267055);
not I_74324 (I1267113,I3570);
DFFARX1 I_74325 (I371805,I3563,I1267113,I1267139,);
nand I_74326 (I1267147,I1267139,I371808);
DFFARX1 I_74327 (I371802,I3563,I1267113,I1267173,);
DFFARX1 I_74328 (I1267173,I3563,I1267113,I1267190,);
not I_74329 (I1267105,I1267190);
not I_74330 (I1267212,I371811);
nor I_74331 (I1267229,I371811,I371796);
not I_74332 (I1267246,I371820);
nand I_74333 (I1267263,I1267212,I1267246);
nor I_74334 (I1267280,I371820,I371811);
and I_74335 (I1267084,I1267280,I1267147);
not I_74336 (I1267311,I371799);
nand I_74337 (I1267328,I1267311,I371817);
nor I_74338 (I1267345,I371799,I371793);
not I_74339 (I1267362,I1267345);
nand I_74340 (I1267087,I1267229,I1267362);
DFFARX1 I_74341 (I1267345,I3563,I1267113,I1267102,);
nor I_74342 (I1267407,I371814,I371820);
nor I_74343 (I1267424,I1267407,I371796);
and I_74344 (I1267441,I1267424,I1267328);
DFFARX1 I_74345 (I1267441,I3563,I1267113,I1267099,);
nor I_74346 (I1267096,I1267407,I1267263);
or I_74347 (I1267093,I1267345,I1267407);
nor I_74348 (I1267500,I371814,I371793);
DFFARX1 I_74349 (I1267500,I3563,I1267113,I1267526,);
not I_74350 (I1267534,I1267526);
nand I_74351 (I1267551,I1267534,I1267212);
nor I_74352 (I1267568,I1267551,I371796);
DFFARX1 I_74353 (I1267568,I3563,I1267113,I1267081,);
nor I_74354 (I1267599,I1267534,I1267263);
nor I_74355 (I1267090,I1267407,I1267599);
not I_74356 (I1267657,I3570);
DFFARX1 I_74357 (I577476,I3563,I1267657,I1267683,);
nand I_74358 (I1267691,I1267683,I577500);
DFFARX1 I_74359 (I577479,I3563,I1267657,I1267717,);
DFFARX1 I_74360 (I1267717,I3563,I1267657,I1267734,);
not I_74361 (I1267649,I1267734);
not I_74362 (I1267756,I577482);
nor I_74363 (I1267773,I577482,I577497);
not I_74364 (I1267790,I577488);
nand I_74365 (I1267807,I1267756,I1267790);
nor I_74366 (I1267824,I577488,I577482);
and I_74367 (I1267628,I1267824,I1267691);
not I_74368 (I1267855,I577485);
nand I_74369 (I1267872,I1267855,I577479);
nor I_74370 (I1267889,I577485,I577494);
not I_74371 (I1267906,I1267889);
nand I_74372 (I1267631,I1267773,I1267906);
DFFARX1 I_74373 (I1267889,I3563,I1267657,I1267646,);
nor I_74374 (I1267951,I577491,I577488);
nor I_74375 (I1267968,I1267951,I577497);
and I_74376 (I1267985,I1267968,I1267872);
DFFARX1 I_74377 (I1267985,I3563,I1267657,I1267643,);
nor I_74378 (I1267640,I1267951,I1267807);
or I_74379 (I1267637,I1267889,I1267951);
nor I_74380 (I1268044,I577491,I577476);
DFFARX1 I_74381 (I1268044,I3563,I1267657,I1268070,);
not I_74382 (I1268078,I1268070);
nand I_74383 (I1268095,I1268078,I1267756);
nor I_74384 (I1268112,I1268095,I577497);
DFFARX1 I_74385 (I1268112,I3563,I1267657,I1267625,);
nor I_74386 (I1268143,I1268078,I1267807);
nor I_74387 (I1267634,I1267951,I1268143);
not I_74388 (I1268201,I3570);
DFFARX1 I_74389 (I239287,I3563,I1268201,I1268227,);
nand I_74390 (I1268235,I1268227,I239302);
DFFARX1 I_74391 (I239299,I3563,I1268201,I1268261,);
DFFARX1 I_74392 (I1268261,I3563,I1268201,I1268278,);
not I_74393 (I1268193,I1268278);
not I_74394 (I1268300,I239278);
nor I_74395 (I1268317,I239278,I239284);
not I_74396 (I1268334,I239290);
nand I_74397 (I1268351,I1268300,I1268334);
nor I_74398 (I1268368,I239290,I239278);
and I_74399 (I1268172,I1268368,I1268235);
not I_74400 (I1268399,I239296);
nand I_74401 (I1268416,I1268399,I239278);
nor I_74402 (I1268433,I239296,I239281);
not I_74403 (I1268450,I1268433);
nand I_74404 (I1268175,I1268317,I1268450);
DFFARX1 I_74405 (I1268433,I3563,I1268201,I1268190,);
nor I_74406 (I1268495,I239281,I239290);
nor I_74407 (I1268512,I1268495,I239284);
and I_74408 (I1268529,I1268512,I1268416);
DFFARX1 I_74409 (I1268529,I3563,I1268201,I1268187,);
nor I_74410 (I1268184,I1268495,I1268351);
or I_74411 (I1268181,I1268433,I1268495);
nor I_74412 (I1268588,I239281,I239293);
DFFARX1 I_74413 (I1268588,I3563,I1268201,I1268614,);
not I_74414 (I1268622,I1268614);
nand I_74415 (I1268639,I1268622,I1268300);
nor I_74416 (I1268656,I1268639,I239284);
DFFARX1 I_74417 (I1268656,I3563,I1268201,I1268169,);
nor I_74418 (I1268687,I1268622,I1268351);
nor I_74419 (I1268178,I1268495,I1268687);
not I_74420 (I1268745,I3570);
DFFARX1 I_74421 (I132029,I3563,I1268745,I1268771,);
nand I_74422 (I1268779,I1268771,I132011);
DFFARX1 I_74423 (I132008,I3563,I1268745,I1268805,);
DFFARX1 I_74424 (I1268805,I3563,I1268745,I1268822,);
not I_74425 (I1268737,I1268822);
not I_74426 (I1268844,I132026);
nor I_74427 (I1268861,I132026,I132020);
not I_74428 (I1268878,I132008);
nand I_74429 (I1268895,I1268844,I1268878);
nor I_74430 (I1268912,I132008,I132026);
and I_74431 (I1268716,I1268912,I1268779);
not I_74432 (I1268943,I132017);
nand I_74433 (I1268960,I1268943,I132023);
nor I_74434 (I1268977,I132017,I132011);
not I_74435 (I1268994,I1268977);
nand I_74436 (I1268719,I1268861,I1268994);
DFFARX1 I_74437 (I1268977,I3563,I1268745,I1268734,);
nor I_74438 (I1269039,I132014,I132008);
nor I_74439 (I1269056,I1269039,I132020);
and I_74440 (I1269073,I1269056,I1268960);
DFFARX1 I_74441 (I1269073,I3563,I1268745,I1268731,);
nor I_74442 (I1268728,I1269039,I1268895);
or I_74443 (I1268725,I1268977,I1269039);
nor I_74444 (I1269132,I132014,I132032);
DFFARX1 I_74445 (I1269132,I3563,I1268745,I1269158,);
not I_74446 (I1269166,I1269158);
nand I_74447 (I1269183,I1269166,I1268844);
nor I_74448 (I1269200,I1269183,I132020);
DFFARX1 I_74449 (I1269200,I3563,I1268745,I1268713,);
nor I_74450 (I1269231,I1269166,I1268895);
nor I_74451 (I1268722,I1269039,I1269231);
not I_74452 (I1269289,I3570);
DFFARX1 I_74453 (I843209,I3563,I1269289,I1269315,);
nand I_74454 (I1269323,I1269315,I843203);
DFFARX1 I_74455 (I843206,I3563,I1269289,I1269349,);
DFFARX1 I_74456 (I1269349,I3563,I1269289,I1269366,);
not I_74457 (I1269281,I1269366);
not I_74458 (I1269388,I843212);
nor I_74459 (I1269405,I843212,I843206);
not I_74460 (I1269422,I843215);
nand I_74461 (I1269439,I1269388,I1269422);
nor I_74462 (I1269456,I843215,I843212);
and I_74463 (I1269260,I1269456,I1269323);
not I_74464 (I1269487,I843224);
nand I_74465 (I1269504,I1269487,I843218);
nor I_74466 (I1269521,I843224,I843221);
not I_74467 (I1269538,I1269521);
nand I_74468 (I1269263,I1269405,I1269538);
DFFARX1 I_74469 (I1269521,I3563,I1269289,I1269278,);
nor I_74470 (I1269583,I843203,I843215);
nor I_74471 (I1269600,I1269583,I843206);
and I_74472 (I1269617,I1269600,I1269504);
DFFARX1 I_74473 (I1269617,I3563,I1269289,I1269275,);
nor I_74474 (I1269272,I1269583,I1269439);
or I_74475 (I1269269,I1269521,I1269583);
nor I_74476 (I1269676,I843203,I843209);
DFFARX1 I_74477 (I1269676,I3563,I1269289,I1269702,);
not I_74478 (I1269710,I1269702);
nand I_74479 (I1269727,I1269710,I1269388);
nor I_74480 (I1269744,I1269727,I843206);
DFFARX1 I_74481 (I1269744,I3563,I1269289,I1269257,);
nor I_74482 (I1269775,I1269710,I1269439);
nor I_74483 (I1269266,I1269583,I1269775);
not I_74484 (I1269833,I3570);
DFFARX1 I_74485 (I600634,I3563,I1269833,I1269859,);
nand I_74486 (I1269867,I1269859,I600622);
DFFARX1 I_74487 (I600628,I3563,I1269833,I1269893,);
DFFARX1 I_74488 (I1269893,I3563,I1269833,I1269910,);
not I_74489 (I1269825,I1269910);
not I_74490 (I1269932,I600613);
nor I_74491 (I1269949,I600613,I600625);
not I_74492 (I1269966,I600616);
nand I_74493 (I1269983,I1269932,I1269966);
nor I_74494 (I1270000,I600616,I600613);
and I_74495 (I1269804,I1270000,I1269867);
not I_74496 (I1270031,I600631);
nand I_74497 (I1270048,I1270031,I600613);
nor I_74498 (I1270065,I600631,I600637);
not I_74499 (I1270082,I1270065);
nand I_74500 (I1269807,I1269949,I1270082);
DFFARX1 I_74501 (I1270065,I3563,I1269833,I1269822,);
nor I_74502 (I1270127,I600619,I600616);
nor I_74503 (I1270144,I1270127,I600625);
and I_74504 (I1270161,I1270144,I1270048);
DFFARX1 I_74505 (I1270161,I3563,I1269833,I1269819,);
nor I_74506 (I1269816,I1270127,I1269983);
or I_74507 (I1269813,I1270065,I1270127);
nor I_74508 (I1270220,I600619,I600616);
DFFARX1 I_74509 (I1270220,I3563,I1269833,I1270246,);
not I_74510 (I1270254,I1270246);
nand I_74511 (I1270271,I1270254,I1269932);
nor I_74512 (I1270288,I1270271,I600625);
DFFARX1 I_74513 (I1270288,I3563,I1269833,I1269801,);
nor I_74514 (I1270319,I1270254,I1269983);
nor I_74515 (I1269810,I1270127,I1270319);
not I_74516 (I1270377,I3570);
DFFARX1 I_74517 (I598900,I3563,I1270377,I1270403,);
nand I_74518 (I1270411,I1270403,I598888);
DFFARX1 I_74519 (I598894,I3563,I1270377,I1270437,);
DFFARX1 I_74520 (I1270437,I3563,I1270377,I1270454,);
not I_74521 (I1270369,I1270454);
not I_74522 (I1270476,I598879);
nor I_74523 (I1270493,I598879,I598891);
not I_74524 (I1270510,I598882);
nand I_74525 (I1270527,I1270476,I1270510);
nor I_74526 (I1270544,I598882,I598879);
and I_74527 (I1270348,I1270544,I1270411);
not I_74528 (I1270575,I598897);
nand I_74529 (I1270592,I1270575,I598879);
nor I_74530 (I1270609,I598897,I598903);
not I_74531 (I1270626,I1270609);
nand I_74532 (I1270351,I1270493,I1270626);
DFFARX1 I_74533 (I1270609,I3563,I1270377,I1270366,);
nor I_74534 (I1270671,I598885,I598882);
nor I_74535 (I1270688,I1270671,I598891);
and I_74536 (I1270705,I1270688,I1270592);
DFFARX1 I_74537 (I1270705,I3563,I1270377,I1270363,);
nor I_74538 (I1270360,I1270671,I1270527);
or I_74539 (I1270357,I1270609,I1270671);
nor I_74540 (I1270764,I598885,I598882);
DFFARX1 I_74541 (I1270764,I3563,I1270377,I1270790,);
not I_74542 (I1270798,I1270790);
nand I_74543 (I1270815,I1270798,I1270476);
nor I_74544 (I1270832,I1270815,I598891);
DFFARX1 I_74545 (I1270832,I3563,I1270377,I1270345,);
nor I_74546 (I1270863,I1270798,I1270527);
nor I_74547 (I1270354,I1270671,I1270863);
not I_74548 (I1270921,I3570);
DFFARX1 I_74549 (I901179,I3563,I1270921,I1270947,);
nand I_74550 (I1270955,I1270947,I901173);
DFFARX1 I_74551 (I901176,I3563,I1270921,I1270981,);
DFFARX1 I_74552 (I1270981,I3563,I1270921,I1270998,);
not I_74553 (I1270913,I1270998);
not I_74554 (I1271020,I901182);
nor I_74555 (I1271037,I901182,I901176);
not I_74556 (I1271054,I901185);
nand I_74557 (I1271071,I1271020,I1271054);
nor I_74558 (I1271088,I901185,I901182);
and I_74559 (I1270892,I1271088,I1270955);
not I_74560 (I1271119,I901194);
nand I_74561 (I1271136,I1271119,I901188);
nor I_74562 (I1271153,I901194,I901191);
not I_74563 (I1271170,I1271153);
nand I_74564 (I1270895,I1271037,I1271170);
DFFARX1 I_74565 (I1271153,I3563,I1270921,I1270910,);
nor I_74566 (I1271215,I901173,I901185);
nor I_74567 (I1271232,I1271215,I901176);
and I_74568 (I1271249,I1271232,I1271136);
DFFARX1 I_74569 (I1271249,I3563,I1270921,I1270907,);
nor I_74570 (I1270904,I1271215,I1271071);
or I_74571 (I1270901,I1271153,I1271215);
nor I_74572 (I1271308,I901173,I901179);
DFFARX1 I_74573 (I1271308,I3563,I1270921,I1271334,);
not I_74574 (I1271342,I1271334);
nand I_74575 (I1271359,I1271342,I1271020);
nor I_74576 (I1271376,I1271359,I901176);
DFFARX1 I_74577 (I1271376,I3563,I1270921,I1270889,);
nor I_74578 (I1271407,I1271342,I1271071);
nor I_74579 (I1270898,I1271215,I1271407);
not I_74580 (I1271465,I3570);
DFFARX1 I_74581 (I1133791,I3563,I1271465,I1271491,);
nand I_74582 (I1271499,I1271491,I1133770);
DFFARX1 I_74583 (I1133767,I3563,I1271465,I1271525,);
DFFARX1 I_74584 (I1271525,I3563,I1271465,I1271542,);
not I_74585 (I1271457,I1271542);
not I_74586 (I1271564,I1133779);
nor I_74587 (I1271581,I1133779,I1133788);
not I_74588 (I1271598,I1133776);
nand I_74589 (I1271615,I1271564,I1271598);
nor I_74590 (I1271632,I1133776,I1133779);
and I_74591 (I1271436,I1271632,I1271499);
not I_74592 (I1271663,I1133785);
nand I_74593 (I1271680,I1271663,I1133782);
nor I_74594 (I1271697,I1133785,I1133767);
not I_74595 (I1271714,I1271697);
nand I_74596 (I1271439,I1271581,I1271714);
DFFARX1 I_74597 (I1271697,I3563,I1271465,I1271454,);
nor I_74598 (I1271759,I1133770,I1133776);
nor I_74599 (I1271776,I1271759,I1133788);
and I_74600 (I1271793,I1271776,I1271680);
DFFARX1 I_74601 (I1271793,I3563,I1271465,I1271451,);
nor I_74602 (I1271448,I1271759,I1271615);
or I_74603 (I1271445,I1271697,I1271759);
nor I_74604 (I1271852,I1133770,I1133773);
DFFARX1 I_74605 (I1271852,I3563,I1271465,I1271878,);
not I_74606 (I1271886,I1271878);
nand I_74607 (I1271903,I1271886,I1271564);
nor I_74608 (I1271920,I1271903,I1133788);
DFFARX1 I_74609 (I1271920,I3563,I1271465,I1271433,);
nor I_74610 (I1271951,I1271886,I1271615);
nor I_74611 (I1271442,I1271759,I1271951);
not I_74612 (I1272009,I3570);
DFFARX1 I_74613 (I1160957,I3563,I1272009,I1272035,);
nand I_74614 (I1272043,I1272035,I1160936);
DFFARX1 I_74615 (I1160933,I3563,I1272009,I1272069,);
DFFARX1 I_74616 (I1272069,I3563,I1272009,I1272086,);
not I_74617 (I1272001,I1272086);
not I_74618 (I1272108,I1160945);
nor I_74619 (I1272125,I1160945,I1160954);
not I_74620 (I1272142,I1160942);
nand I_74621 (I1272159,I1272108,I1272142);
nor I_74622 (I1272176,I1160942,I1160945);
and I_74623 (I1271980,I1272176,I1272043);
not I_74624 (I1272207,I1160951);
nand I_74625 (I1272224,I1272207,I1160948);
nor I_74626 (I1272241,I1160951,I1160933);
not I_74627 (I1272258,I1272241);
nand I_74628 (I1271983,I1272125,I1272258);
DFFARX1 I_74629 (I1272241,I3563,I1272009,I1271998,);
nor I_74630 (I1272303,I1160936,I1160942);
nor I_74631 (I1272320,I1272303,I1160954);
and I_74632 (I1272337,I1272320,I1272224);
DFFARX1 I_74633 (I1272337,I3563,I1272009,I1271995,);
nor I_74634 (I1271992,I1272303,I1272159);
or I_74635 (I1271989,I1272241,I1272303);
nor I_74636 (I1272396,I1160936,I1160939);
DFFARX1 I_74637 (I1272396,I3563,I1272009,I1272422,);
not I_74638 (I1272430,I1272422);
nand I_74639 (I1272447,I1272430,I1272108);
nor I_74640 (I1272464,I1272447,I1160954);
DFFARX1 I_74641 (I1272464,I3563,I1272009,I1271977,);
nor I_74642 (I1272495,I1272430,I1272159);
nor I_74643 (I1271986,I1272303,I1272495);
not I_74644 (I1272553,I3570);
DFFARX1 I_74645 (I1406525,I3563,I1272553,I1272579,);
nand I_74646 (I1272587,I1272579,I1406510);
DFFARX1 I_74647 (I1406504,I3563,I1272553,I1272613,);
DFFARX1 I_74648 (I1272613,I3563,I1272553,I1272630,);
not I_74649 (I1272545,I1272630);
not I_74650 (I1272652,I1406498);
nor I_74651 (I1272669,I1406498,I1406519);
not I_74652 (I1272686,I1406507);
nand I_74653 (I1272703,I1272652,I1272686);
nor I_74654 (I1272720,I1406507,I1406498);
and I_74655 (I1272524,I1272720,I1272587);
not I_74656 (I1272751,I1406516);
nand I_74657 (I1272768,I1272751,I1406522);
nor I_74658 (I1272785,I1406516,I1406513);
not I_74659 (I1272802,I1272785);
nand I_74660 (I1272527,I1272669,I1272802);
DFFARX1 I_74661 (I1272785,I3563,I1272553,I1272542,);
nor I_74662 (I1272847,I1406501,I1406507);
nor I_74663 (I1272864,I1272847,I1406519);
and I_74664 (I1272881,I1272864,I1272768);
DFFARX1 I_74665 (I1272881,I3563,I1272553,I1272539,);
nor I_74666 (I1272536,I1272847,I1272703);
or I_74667 (I1272533,I1272785,I1272847);
nor I_74668 (I1272940,I1406501,I1406498);
DFFARX1 I_74669 (I1272940,I3563,I1272553,I1272966,);
not I_74670 (I1272974,I1272966);
nand I_74671 (I1272991,I1272974,I1272652);
nor I_74672 (I1273008,I1272991,I1406519);
DFFARX1 I_74673 (I1273008,I3563,I1272553,I1272521,);
nor I_74674 (I1273039,I1272974,I1272703);
nor I_74675 (I1272530,I1272847,I1273039);
not I_74676 (I1273097,I3570);
DFFARX1 I_74677 (I111476,I3563,I1273097,I1273123,);
nand I_74678 (I1273131,I1273123,I111458);
DFFARX1 I_74679 (I111455,I3563,I1273097,I1273157,);
DFFARX1 I_74680 (I1273157,I3563,I1273097,I1273174,);
not I_74681 (I1273089,I1273174);
not I_74682 (I1273196,I111473);
nor I_74683 (I1273213,I111473,I111467);
not I_74684 (I1273230,I111455);
nand I_74685 (I1273247,I1273196,I1273230);
nor I_74686 (I1273264,I111455,I111473);
and I_74687 (I1273068,I1273264,I1273131);
not I_74688 (I1273295,I111464);
nand I_74689 (I1273312,I1273295,I111470);
nor I_74690 (I1273329,I111464,I111458);
not I_74691 (I1273346,I1273329);
nand I_74692 (I1273071,I1273213,I1273346);
DFFARX1 I_74693 (I1273329,I3563,I1273097,I1273086,);
nor I_74694 (I1273391,I111461,I111455);
nor I_74695 (I1273408,I1273391,I111467);
and I_74696 (I1273425,I1273408,I1273312);
DFFARX1 I_74697 (I1273425,I3563,I1273097,I1273083,);
nor I_74698 (I1273080,I1273391,I1273247);
or I_74699 (I1273077,I1273329,I1273391);
nor I_74700 (I1273484,I111461,I111479);
DFFARX1 I_74701 (I1273484,I3563,I1273097,I1273510,);
not I_74702 (I1273518,I1273510);
nand I_74703 (I1273535,I1273518,I1273196);
nor I_74704 (I1273552,I1273535,I111467);
DFFARX1 I_74705 (I1273552,I3563,I1273097,I1273065,);
nor I_74706 (I1273583,I1273518,I1273247);
nor I_74707 (I1273074,I1273391,I1273583);
not I_74708 (I1273641,I3570);
DFFARX1 I_74709 (I988519,I3563,I1273641,I1273667,);
nand I_74710 (I1273675,I1273667,I988519);
DFFARX1 I_74711 (I988531,I3563,I1273641,I1273701,);
DFFARX1 I_74712 (I1273701,I3563,I1273641,I1273718,);
not I_74713 (I1273633,I1273718);
not I_74714 (I1273740,I988525);
nor I_74715 (I1273757,I988525,I988546);
not I_74716 (I1273774,I988534);
nand I_74717 (I1273791,I1273740,I1273774);
nor I_74718 (I1273808,I988534,I988525);
and I_74719 (I1273612,I1273808,I1273675);
not I_74720 (I1273839,I988528);
nand I_74721 (I1273856,I1273839,I988543);
nor I_74722 (I1273873,I988528,I988537);
not I_74723 (I1273890,I1273873);
nand I_74724 (I1273615,I1273757,I1273890);
DFFARX1 I_74725 (I1273873,I3563,I1273641,I1273630,);
nor I_74726 (I1273935,I988540,I988534);
nor I_74727 (I1273952,I1273935,I988546);
and I_74728 (I1273969,I1273952,I1273856);
DFFARX1 I_74729 (I1273969,I3563,I1273641,I1273627,);
nor I_74730 (I1273624,I1273935,I1273791);
or I_74731 (I1273621,I1273873,I1273935);
nor I_74732 (I1274028,I988540,I988522);
DFFARX1 I_74733 (I1274028,I3563,I1273641,I1274054,);
not I_74734 (I1274062,I1274054);
nand I_74735 (I1274079,I1274062,I1273740);
nor I_74736 (I1274096,I1274079,I988546);
DFFARX1 I_74737 (I1274096,I3563,I1273641,I1273609,);
nor I_74738 (I1274127,I1274062,I1273791);
nor I_74739 (I1273618,I1273935,I1274127);
not I_74740 (I1274185,I3570);
DFFARX1 I_74741 (I447450,I3563,I1274185,I1274211,);
nand I_74742 (I1274219,I1274211,I447447);
DFFARX1 I_74743 (I447426,I3563,I1274185,I1274245,);
DFFARX1 I_74744 (I1274245,I3563,I1274185,I1274262,);
not I_74745 (I1274177,I1274262);
not I_74746 (I1274284,I447441);
nor I_74747 (I1274301,I447441,I447444);
not I_74748 (I1274318,I447435);
nand I_74749 (I1274335,I1274284,I1274318);
nor I_74750 (I1274352,I447435,I447441);
and I_74751 (I1274156,I1274352,I1274219);
not I_74752 (I1274383,I447432);
nand I_74753 (I1274400,I1274383,I447453);
nor I_74754 (I1274417,I447432,I447429);
not I_74755 (I1274434,I1274417);
nand I_74756 (I1274159,I1274301,I1274434);
DFFARX1 I_74757 (I1274417,I3563,I1274185,I1274174,);
nor I_74758 (I1274479,I447438,I447435);
nor I_74759 (I1274496,I1274479,I447444);
and I_74760 (I1274513,I1274496,I1274400);
DFFARX1 I_74761 (I1274513,I3563,I1274185,I1274171,);
nor I_74762 (I1274168,I1274479,I1274335);
or I_74763 (I1274165,I1274417,I1274479);
nor I_74764 (I1274572,I447438,I447426);
DFFARX1 I_74765 (I1274572,I3563,I1274185,I1274598,);
not I_74766 (I1274606,I1274598);
nand I_74767 (I1274623,I1274606,I1274284);
nor I_74768 (I1274640,I1274623,I447444);
DFFARX1 I_74769 (I1274640,I3563,I1274185,I1274153,);
nor I_74770 (I1274671,I1274606,I1274335);
nor I_74771 (I1274162,I1274479,I1274671);
not I_74772 (I1274729,I3570);
DFFARX1 I_74773 (I455610,I3563,I1274729,I1274755,);
nand I_74774 (I1274763,I1274755,I455607);
DFFARX1 I_74775 (I455586,I3563,I1274729,I1274789,);
DFFARX1 I_74776 (I1274789,I3563,I1274729,I1274806,);
not I_74777 (I1274721,I1274806);
not I_74778 (I1274828,I455601);
nor I_74779 (I1274845,I455601,I455604);
not I_74780 (I1274862,I455595);
nand I_74781 (I1274879,I1274828,I1274862);
nor I_74782 (I1274896,I455595,I455601);
and I_74783 (I1274700,I1274896,I1274763);
not I_74784 (I1274927,I455592);
nand I_74785 (I1274944,I1274927,I455613);
nor I_74786 (I1274961,I455592,I455589);
not I_74787 (I1274978,I1274961);
nand I_74788 (I1274703,I1274845,I1274978);
DFFARX1 I_74789 (I1274961,I3563,I1274729,I1274718,);
nor I_74790 (I1275023,I455598,I455595);
nor I_74791 (I1275040,I1275023,I455604);
and I_74792 (I1275057,I1275040,I1274944);
DFFARX1 I_74793 (I1275057,I3563,I1274729,I1274715,);
nor I_74794 (I1274712,I1275023,I1274879);
or I_74795 (I1274709,I1274961,I1275023);
nor I_74796 (I1275116,I455598,I455586);
DFFARX1 I_74797 (I1275116,I3563,I1274729,I1275142,);
not I_74798 (I1275150,I1275142);
nand I_74799 (I1275167,I1275150,I1274828);
nor I_74800 (I1275184,I1275167,I455604);
DFFARX1 I_74801 (I1275184,I3563,I1274729,I1274697,);
nor I_74802 (I1275215,I1275150,I1274879);
nor I_74803 (I1274706,I1275023,I1275215);
not I_74804 (I1275273,I3570);
DFFARX1 I_74805 (I4177,I3563,I1275273,I1275299,);
nand I_74806 (I1275307,I1275299,I4189);
DFFARX1 I_74807 (I4186,I3563,I1275273,I1275333,);
DFFARX1 I_74808 (I1275333,I3563,I1275273,I1275350,);
not I_74809 (I1275265,I1275350);
not I_74810 (I1275372,I4174);
nor I_74811 (I1275389,I4174,I4174);
not I_74812 (I1275406,I4168);
nand I_74813 (I1275423,I1275372,I1275406);
nor I_74814 (I1275440,I4168,I4174);
and I_74815 (I1275244,I1275440,I1275307);
not I_74816 (I1275471,I4171);
nand I_74817 (I1275488,I1275471,I4171);
nor I_74818 (I1275505,I4171,I4180);
not I_74819 (I1275522,I1275505);
nand I_74820 (I1275247,I1275389,I1275522);
DFFARX1 I_74821 (I1275505,I3563,I1275273,I1275262,);
nor I_74822 (I1275567,I4168,I4168);
nor I_74823 (I1275584,I1275567,I4174);
and I_74824 (I1275601,I1275584,I1275488);
DFFARX1 I_74825 (I1275601,I3563,I1275273,I1275259,);
nor I_74826 (I1275256,I1275567,I1275423);
or I_74827 (I1275253,I1275505,I1275567);
nor I_74828 (I1275660,I4168,I4183);
DFFARX1 I_74829 (I1275660,I3563,I1275273,I1275686,);
not I_74830 (I1275694,I1275686);
nand I_74831 (I1275711,I1275694,I1275372);
nor I_74832 (I1275728,I1275711,I4174);
DFFARX1 I_74833 (I1275728,I3563,I1275273,I1275241,);
nor I_74834 (I1275759,I1275694,I1275423);
nor I_74835 (I1275250,I1275567,I1275759);
not I_74836 (I1275817,I3570);
DFFARX1 I_74837 (I400790,I3563,I1275817,I1275843,);
nand I_74838 (I1275851,I1275843,I400793);
DFFARX1 I_74839 (I400787,I3563,I1275817,I1275877,);
DFFARX1 I_74840 (I1275877,I3563,I1275817,I1275894,);
not I_74841 (I1275809,I1275894);
not I_74842 (I1275916,I400796);
nor I_74843 (I1275933,I400796,I400781);
not I_74844 (I1275950,I400805);
nand I_74845 (I1275967,I1275916,I1275950);
nor I_74846 (I1275984,I400805,I400796);
and I_74847 (I1275788,I1275984,I1275851);
not I_74848 (I1276015,I400784);
nand I_74849 (I1276032,I1276015,I400802);
nor I_74850 (I1276049,I400784,I400778);
not I_74851 (I1276066,I1276049);
nand I_74852 (I1275791,I1275933,I1276066);
DFFARX1 I_74853 (I1276049,I3563,I1275817,I1275806,);
nor I_74854 (I1276111,I400799,I400805);
nor I_74855 (I1276128,I1276111,I400781);
and I_74856 (I1276145,I1276128,I1276032);
DFFARX1 I_74857 (I1276145,I3563,I1275817,I1275803,);
nor I_74858 (I1275800,I1276111,I1275967);
or I_74859 (I1275797,I1276049,I1276111);
nor I_74860 (I1276204,I400799,I400778);
DFFARX1 I_74861 (I1276204,I3563,I1275817,I1276230,);
not I_74862 (I1276238,I1276230);
nand I_74863 (I1276255,I1276238,I1275916);
nor I_74864 (I1276272,I1276255,I400781);
DFFARX1 I_74865 (I1276272,I3563,I1275817,I1275785,);
nor I_74866 (I1276303,I1276238,I1275967);
nor I_74867 (I1275794,I1276111,I1276303);
not I_74868 (I1276361,I3570);
DFFARX1 I_74869 (I1184655,I3563,I1276361,I1276387,);
nand I_74870 (I1276395,I1276387,I1184634);
DFFARX1 I_74871 (I1184631,I3563,I1276361,I1276421,);
DFFARX1 I_74872 (I1276421,I3563,I1276361,I1276438,);
not I_74873 (I1276353,I1276438);
not I_74874 (I1276460,I1184643);
nor I_74875 (I1276477,I1184643,I1184652);
not I_74876 (I1276494,I1184640);
nand I_74877 (I1276511,I1276460,I1276494);
nor I_74878 (I1276528,I1184640,I1184643);
and I_74879 (I1276332,I1276528,I1276395);
not I_74880 (I1276559,I1184649);
nand I_74881 (I1276576,I1276559,I1184646);
nor I_74882 (I1276593,I1184649,I1184631);
not I_74883 (I1276610,I1276593);
nand I_74884 (I1276335,I1276477,I1276610);
DFFARX1 I_74885 (I1276593,I3563,I1276361,I1276350,);
nor I_74886 (I1276655,I1184634,I1184640);
nor I_74887 (I1276672,I1276655,I1184652);
and I_74888 (I1276689,I1276672,I1276576);
DFFARX1 I_74889 (I1276689,I3563,I1276361,I1276347,);
nor I_74890 (I1276344,I1276655,I1276511);
or I_74891 (I1276341,I1276593,I1276655);
nor I_74892 (I1276748,I1184634,I1184637);
DFFARX1 I_74893 (I1276748,I3563,I1276361,I1276774,);
not I_74894 (I1276782,I1276774);
nand I_74895 (I1276799,I1276782,I1276460);
nor I_74896 (I1276816,I1276799,I1184652);
DFFARX1 I_74897 (I1276816,I3563,I1276361,I1276329,);
nor I_74898 (I1276847,I1276782,I1276511);
nor I_74899 (I1276338,I1276655,I1276847);
not I_74900 (I1276905,I3570);
DFFARX1 I_74901 (I696564,I3563,I1276905,I1276931,);
nand I_74902 (I1276939,I1276931,I696579);
DFFARX1 I_74903 (I696573,I3563,I1276905,I1276965,);
DFFARX1 I_74904 (I1276965,I3563,I1276905,I1276982,);
not I_74905 (I1276897,I1276982);
not I_74906 (I1277004,I696576);
nor I_74907 (I1277021,I696576,I696582);
not I_74908 (I1277038,I696564);
nand I_74909 (I1277055,I1277004,I1277038);
nor I_74910 (I1277072,I696564,I696576);
and I_74911 (I1276876,I1277072,I1276939);
not I_74912 (I1277103,I696561);
nand I_74913 (I1277120,I1277103,I696567);
nor I_74914 (I1277137,I696561,I696561);
not I_74915 (I1277154,I1277137);
nand I_74916 (I1276879,I1277021,I1277154);
DFFARX1 I_74917 (I1277137,I3563,I1276905,I1276894,);
nor I_74918 (I1277199,I696570,I696564);
nor I_74919 (I1277216,I1277199,I696582);
and I_74920 (I1277233,I1277216,I1277120);
DFFARX1 I_74921 (I1277233,I3563,I1276905,I1276891,);
nor I_74922 (I1276888,I1277199,I1277055);
or I_74923 (I1276885,I1277137,I1277199);
nor I_74924 (I1277292,I696570,I696585);
DFFARX1 I_74925 (I1277292,I3563,I1276905,I1277318,);
not I_74926 (I1277326,I1277318);
nand I_74927 (I1277343,I1277326,I1277004);
nor I_74928 (I1277360,I1277343,I696582);
DFFARX1 I_74929 (I1277360,I3563,I1276905,I1276873,);
nor I_74930 (I1277391,I1277326,I1277055);
nor I_74931 (I1276882,I1277199,I1277391);
not I_74932 (I1277449,I3570);
DFFARX1 I_74933 (I730666,I3563,I1277449,I1277475,);
nand I_74934 (I1277483,I1277475,I730681);
DFFARX1 I_74935 (I730675,I3563,I1277449,I1277509,);
DFFARX1 I_74936 (I1277509,I3563,I1277449,I1277526,);
not I_74937 (I1277441,I1277526);
not I_74938 (I1277548,I730678);
nor I_74939 (I1277565,I730678,I730684);
not I_74940 (I1277582,I730666);
nand I_74941 (I1277599,I1277548,I1277582);
nor I_74942 (I1277616,I730666,I730678);
and I_74943 (I1277420,I1277616,I1277483);
not I_74944 (I1277647,I730663);
nand I_74945 (I1277664,I1277647,I730669);
nor I_74946 (I1277681,I730663,I730663);
not I_74947 (I1277698,I1277681);
nand I_74948 (I1277423,I1277565,I1277698);
DFFARX1 I_74949 (I1277681,I3563,I1277449,I1277438,);
nor I_74950 (I1277743,I730672,I730666);
nor I_74951 (I1277760,I1277743,I730684);
and I_74952 (I1277777,I1277760,I1277664);
DFFARX1 I_74953 (I1277777,I3563,I1277449,I1277435,);
nor I_74954 (I1277432,I1277743,I1277599);
or I_74955 (I1277429,I1277681,I1277743);
nor I_74956 (I1277836,I730672,I730687);
DFFARX1 I_74957 (I1277836,I3563,I1277449,I1277862,);
not I_74958 (I1277870,I1277862);
nand I_74959 (I1277887,I1277870,I1277548);
nor I_74960 (I1277904,I1277887,I730684);
DFFARX1 I_74961 (I1277904,I3563,I1277449,I1277417,);
nor I_74962 (I1277935,I1277870,I1277599);
nor I_74963 (I1277426,I1277743,I1277935);
not I_74964 (I1277993,I3570);
DFFARX1 I_74965 (I934901,I3563,I1277993,I1278019,);
nand I_74966 (I1278027,I1278019,I934901);
DFFARX1 I_74967 (I934913,I3563,I1277993,I1278053,);
DFFARX1 I_74968 (I1278053,I3563,I1277993,I1278070,);
not I_74969 (I1277985,I1278070);
not I_74970 (I1278092,I934907);
nor I_74971 (I1278109,I934907,I934928);
not I_74972 (I1278126,I934916);
nand I_74973 (I1278143,I1278092,I1278126);
nor I_74974 (I1278160,I934916,I934907);
and I_74975 (I1277964,I1278160,I1278027);
not I_74976 (I1278191,I934910);
nand I_74977 (I1278208,I1278191,I934925);
nor I_74978 (I1278225,I934910,I934919);
not I_74979 (I1278242,I1278225);
nand I_74980 (I1277967,I1278109,I1278242);
DFFARX1 I_74981 (I1278225,I3563,I1277993,I1277982,);
nor I_74982 (I1278287,I934922,I934916);
nor I_74983 (I1278304,I1278287,I934928);
and I_74984 (I1278321,I1278304,I1278208);
DFFARX1 I_74985 (I1278321,I3563,I1277993,I1277979,);
nor I_74986 (I1277976,I1278287,I1278143);
or I_74987 (I1277973,I1278225,I1278287);
nor I_74988 (I1278380,I934922,I934904);
DFFARX1 I_74989 (I1278380,I3563,I1277993,I1278406,);
not I_74990 (I1278414,I1278406);
nand I_74991 (I1278431,I1278414,I1278092);
nor I_74992 (I1278448,I1278431,I934928);
DFFARX1 I_74993 (I1278448,I3563,I1277993,I1277961,);
nor I_74994 (I1278479,I1278414,I1278143);
nor I_74995 (I1277970,I1278287,I1278479);
not I_74996 (I1278537,I3570);
DFFARX1 I_74997 (I1121075,I3563,I1278537,I1278563,);
nand I_74998 (I1278571,I1278563,I1121054);
DFFARX1 I_74999 (I1121051,I3563,I1278537,I1278597,);
DFFARX1 I_75000 (I1278597,I3563,I1278537,I1278614,);
not I_75001 (I1278529,I1278614);
not I_75002 (I1278636,I1121063);
nor I_75003 (I1278653,I1121063,I1121072);
not I_75004 (I1278670,I1121060);
nand I_75005 (I1278687,I1278636,I1278670);
nor I_75006 (I1278704,I1121060,I1121063);
and I_75007 (I1278508,I1278704,I1278571);
not I_75008 (I1278735,I1121069);
nand I_75009 (I1278752,I1278735,I1121066);
nor I_75010 (I1278769,I1121069,I1121051);
not I_75011 (I1278786,I1278769);
nand I_75012 (I1278511,I1278653,I1278786);
DFFARX1 I_75013 (I1278769,I3563,I1278537,I1278526,);
nor I_75014 (I1278831,I1121054,I1121060);
nor I_75015 (I1278848,I1278831,I1121072);
and I_75016 (I1278865,I1278848,I1278752);
DFFARX1 I_75017 (I1278865,I3563,I1278537,I1278523,);
nor I_75018 (I1278520,I1278831,I1278687);
or I_75019 (I1278517,I1278769,I1278831);
nor I_75020 (I1278924,I1121054,I1121057);
DFFARX1 I_75021 (I1278924,I3563,I1278537,I1278950,);
not I_75022 (I1278958,I1278950);
nand I_75023 (I1278975,I1278958,I1278636);
nor I_75024 (I1278992,I1278975,I1121072);
DFFARX1 I_75025 (I1278992,I3563,I1278537,I1278505,);
nor I_75026 (I1279023,I1278958,I1278687);
nor I_75027 (I1278514,I1278831,I1279023);
not I_75028 (I1279081,I3570);
DFFARX1 I_75029 (I338604,I3563,I1279081,I1279107,);
nand I_75030 (I1279115,I1279107,I338607);
DFFARX1 I_75031 (I338601,I3563,I1279081,I1279141,);
DFFARX1 I_75032 (I1279141,I3563,I1279081,I1279158,);
not I_75033 (I1279073,I1279158);
not I_75034 (I1279180,I338610);
nor I_75035 (I1279197,I338610,I338595);
not I_75036 (I1279214,I338619);
nand I_75037 (I1279231,I1279180,I1279214);
nor I_75038 (I1279248,I338619,I338610);
and I_75039 (I1279052,I1279248,I1279115);
not I_75040 (I1279279,I338598);
nand I_75041 (I1279296,I1279279,I338616);
nor I_75042 (I1279313,I338598,I338592);
not I_75043 (I1279330,I1279313);
nand I_75044 (I1279055,I1279197,I1279330);
DFFARX1 I_75045 (I1279313,I3563,I1279081,I1279070,);
nor I_75046 (I1279375,I338613,I338619);
nor I_75047 (I1279392,I1279375,I338595);
and I_75048 (I1279409,I1279392,I1279296);
DFFARX1 I_75049 (I1279409,I3563,I1279081,I1279067,);
nor I_75050 (I1279064,I1279375,I1279231);
or I_75051 (I1279061,I1279313,I1279375);
nor I_75052 (I1279468,I338613,I338592);
DFFARX1 I_75053 (I1279468,I3563,I1279081,I1279494,);
not I_75054 (I1279502,I1279494);
nand I_75055 (I1279519,I1279502,I1279180);
nor I_75056 (I1279536,I1279519,I338595);
DFFARX1 I_75057 (I1279536,I3563,I1279081,I1279049,);
nor I_75058 (I1279567,I1279502,I1279231);
nor I_75059 (I1279058,I1279375,I1279567);
not I_75060 (I1279625,I3570);
DFFARX1 I_75061 (I762456,I3563,I1279625,I1279651,);
nand I_75062 (I1279659,I1279651,I762471);
DFFARX1 I_75063 (I762465,I3563,I1279625,I1279685,);
DFFARX1 I_75064 (I1279685,I3563,I1279625,I1279702,);
not I_75065 (I1279617,I1279702);
not I_75066 (I1279724,I762468);
nor I_75067 (I1279741,I762468,I762474);
not I_75068 (I1279758,I762456);
nand I_75069 (I1279775,I1279724,I1279758);
nor I_75070 (I1279792,I762456,I762468);
and I_75071 (I1279596,I1279792,I1279659);
not I_75072 (I1279823,I762453);
nand I_75073 (I1279840,I1279823,I762459);
nor I_75074 (I1279857,I762453,I762453);
not I_75075 (I1279874,I1279857);
nand I_75076 (I1279599,I1279741,I1279874);
DFFARX1 I_75077 (I1279857,I3563,I1279625,I1279614,);
nor I_75078 (I1279919,I762462,I762456);
nor I_75079 (I1279936,I1279919,I762474);
and I_75080 (I1279953,I1279936,I1279840);
DFFARX1 I_75081 (I1279953,I3563,I1279625,I1279611,);
nor I_75082 (I1279608,I1279919,I1279775);
or I_75083 (I1279605,I1279857,I1279919);
nor I_75084 (I1280012,I762462,I762477);
DFFARX1 I_75085 (I1280012,I3563,I1279625,I1280038,);
not I_75086 (I1280046,I1280038);
nand I_75087 (I1280063,I1280046,I1279724);
nor I_75088 (I1280080,I1280063,I762474);
DFFARX1 I_75089 (I1280080,I3563,I1279625,I1279593,);
nor I_75090 (I1280111,I1280046,I1279775);
nor I_75091 (I1279602,I1279919,I1280111);
not I_75092 (I1280169,I3570);
DFFARX1 I_75093 (I1326438,I3563,I1280169,I1280195,);
nand I_75094 (I1280203,I1280195,I1326423);
DFFARX1 I_75095 (I1326435,I3563,I1280169,I1280229,);
DFFARX1 I_75096 (I1280229,I3563,I1280169,I1280246,);
not I_75097 (I1280161,I1280246);
not I_75098 (I1280268,I1326429);
nor I_75099 (I1280285,I1326429,I1326420);
not I_75100 (I1280302,I1326414);
nand I_75101 (I1280319,I1280268,I1280302);
nor I_75102 (I1280336,I1326414,I1326429);
and I_75103 (I1280140,I1280336,I1280203);
not I_75104 (I1280367,I1326426);
nand I_75105 (I1280384,I1280367,I1326411);
nor I_75106 (I1280401,I1326426,I1326432);
not I_75107 (I1280418,I1280401);
nand I_75108 (I1280143,I1280285,I1280418);
DFFARX1 I_75109 (I1280401,I3563,I1280169,I1280158,);
nor I_75110 (I1280463,I1326417,I1326414);
nor I_75111 (I1280480,I1280463,I1326420);
and I_75112 (I1280497,I1280480,I1280384);
DFFARX1 I_75113 (I1280497,I3563,I1280169,I1280155,);
nor I_75114 (I1280152,I1280463,I1280319);
or I_75115 (I1280149,I1280401,I1280463);
nor I_75116 (I1280556,I1326417,I1326411);
DFFARX1 I_75117 (I1280556,I3563,I1280169,I1280582,);
not I_75118 (I1280590,I1280582);
nand I_75119 (I1280607,I1280590,I1280268);
nor I_75120 (I1280624,I1280607,I1326420);
DFFARX1 I_75121 (I1280624,I3563,I1280169,I1280137,);
nor I_75122 (I1280655,I1280590,I1280319);
nor I_75123 (I1280146,I1280463,I1280655);
not I_75124 (I1280713,I3570);
DFFARX1 I_75125 (I1214711,I3563,I1280713,I1280739,);
nand I_75126 (I1280747,I1280739,I1214690);
DFFARX1 I_75127 (I1214687,I3563,I1280713,I1280773,);
DFFARX1 I_75128 (I1280773,I3563,I1280713,I1280790,);
not I_75129 (I1280705,I1280790);
not I_75130 (I1280812,I1214699);
nor I_75131 (I1280829,I1214699,I1214708);
not I_75132 (I1280846,I1214696);
nand I_75133 (I1280863,I1280812,I1280846);
nor I_75134 (I1280880,I1214696,I1214699);
and I_75135 (I1280684,I1280880,I1280747);
not I_75136 (I1280911,I1214705);
nand I_75137 (I1280928,I1280911,I1214702);
nor I_75138 (I1280945,I1214705,I1214687);
not I_75139 (I1280962,I1280945);
nand I_75140 (I1280687,I1280829,I1280962);
DFFARX1 I_75141 (I1280945,I3563,I1280713,I1280702,);
nor I_75142 (I1281007,I1214690,I1214696);
nor I_75143 (I1281024,I1281007,I1214708);
and I_75144 (I1281041,I1281024,I1280928);
DFFARX1 I_75145 (I1281041,I3563,I1280713,I1280699,);
nor I_75146 (I1280696,I1281007,I1280863);
or I_75147 (I1280693,I1280945,I1281007);
nor I_75148 (I1281100,I1214690,I1214693);
DFFARX1 I_75149 (I1281100,I3563,I1280713,I1281126,);
not I_75150 (I1281134,I1281126);
nand I_75151 (I1281151,I1281134,I1280812);
nor I_75152 (I1281168,I1281151,I1214708);
DFFARX1 I_75153 (I1281168,I3563,I1280713,I1280681,);
nor I_75154 (I1281199,I1281134,I1280863);
nor I_75155 (I1280690,I1281007,I1281199);
not I_75156 (I1281257,I3570);
DFFARX1 I_75157 (I438746,I3563,I1281257,I1281283,);
nand I_75158 (I1281291,I1281283,I438743);
DFFARX1 I_75159 (I438722,I3563,I1281257,I1281317,);
DFFARX1 I_75160 (I1281317,I3563,I1281257,I1281334,);
not I_75161 (I1281249,I1281334);
not I_75162 (I1281356,I438737);
nor I_75163 (I1281373,I438737,I438740);
not I_75164 (I1281390,I438731);
nand I_75165 (I1281407,I1281356,I1281390);
nor I_75166 (I1281424,I438731,I438737);
and I_75167 (I1281228,I1281424,I1281291);
not I_75168 (I1281455,I438728);
nand I_75169 (I1281472,I1281455,I438749);
nor I_75170 (I1281489,I438728,I438725);
not I_75171 (I1281506,I1281489);
nand I_75172 (I1281231,I1281373,I1281506);
DFFARX1 I_75173 (I1281489,I3563,I1281257,I1281246,);
nor I_75174 (I1281551,I438734,I438731);
nor I_75175 (I1281568,I1281551,I438740);
and I_75176 (I1281585,I1281568,I1281472);
DFFARX1 I_75177 (I1281585,I3563,I1281257,I1281243,);
nor I_75178 (I1281240,I1281551,I1281407);
or I_75179 (I1281237,I1281489,I1281551);
nor I_75180 (I1281644,I438734,I438722);
DFFARX1 I_75181 (I1281644,I3563,I1281257,I1281670,);
not I_75182 (I1281678,I1281670);
nand I_75183 (I1281695,I1281678,I1281356);
nor I_75184 (I1281712,I1281695,I438740);
DFFARX1 I_75185 (I1281712,I3563,I1281257,I1281225,);
nor I_75186 (I1281743,I1281678,I1281407);
nor I_75187 (I1281234,I1281551,I1281743);
not I_75188 (I1281801,I3570);
DFFARX1 I_75189 (I754942,I3563,I1281801,I1281827,);
nand I_75190 (I1281835,I1281827,I754957);
DFFARX1 I_75191 (I754951,I3563,I1281801,I1281861,);
DFFARX1 I_75192 (I1281861,I3563,I1281801,I1281878,);
not I_75193 (I1281793,I1281878);
not I_75194 (I1281900,I754954);
nor I_75195 (I1281917,I754954,I754960);
not I_75196 (I1281934,I754942);
nand I_75197 (I1281951,I1281900,I1281934);
nor I_75198 (I1281968,I754942,I754954);
and I_75199 (I1281772,I1281968,I1281835);
not I_75200 (I1281999,I754939);
nand I_75201 (I1282016,I1281999,I754945);
nor I_75202 (I1282033,I754939,I754939);
not I_75203 (I1282050,I1282033);
nand I_75204 (I1281775,I1281917,I1282050);
DFFARX1 I_75205 (I1282033,I3563,I1281801,I1281790,);
nor I_75206 (I1282095,I754948,I754942);
nor I_75207 (I1282112,I1282095,I754960);
and I_75208 (I1282129,I1282112,I1282016);
DFFARX1 I_75209 (I1282129,I3563,I1281801,I1281787,);
nor I_75210 (I1281784,I1282095,I1281951);
or I_75211 (I1281781,I1282033,I1282095);
nor I_75212 (I1282188,I754948,I754963);
DFFARX1 I_75213 (I1282188,I3563,I1281801,I1282214,);
not I_75214 (I1282222,I1282214);
nand I_75215 (I1282239,I1282222,I1281900);
nor I_75216 (I1282256,I1282239,I754960);
DFFARX1 I_75217 (I1282256,I3563,I1281801,I1281769,);
nor I_75218 (I1282287,I1282222,I1281951);
nor I_75219 (I1281778,I1282095,I1282287);
not I_75220 (I1282345,I3570);
DFFARX1 I_75221 (I476282,I3563,I1282345,I1282371,);
nand I_75222 (I1282379,I1282371,I476279);
DFFARX1 I_75223 (I476258,I3563,I1282345,I1282405,);
DFFARX1 I_75224 (I1282405,I3563,I1282345,I1282422,);
not I_75225 (I1282337,I1282422);
not I_75226 (I1282444,I476273);
nor I_75227 (I1282461,I476273,I476276);
not I_75228 (I1282478,I476267);
nand I_75229 (I1282495,I1282444,I1282478);
nor I_75230 (I1282512,I476267,I476273);
and I_75231 (I1282316,I1282512,I1282379);
not I_75232 (I1282543,I476264);
nand I_75233 (I1282560,I1282543,I476285);
nor I_75234 (I1282577,I476264,I476261);
not I_75235 (I1282594,I1282577);
nand I_75236 (I1282319,I1282461,I1282594);
DFFARX1 I_75237 (I1282577,I3563,I1282345,I1282334,);
nor I_75238 (I1282639,I476270,I476267);
nor I_75239 (I1282656,I1282639,I476276);
and I_75240 (I1282673,I1282656,I1282560);
DFFARX1 I_75241 (I1282673,I3563,I1282345,I1282331,);
nor I_75242 (I1282328,I1282639,I1282495);
or I_75243 (I1282325,I1282577,I1282639);
nor I_75244 (I1282732,I476270,I476258);
DFFARX1 I_75245 (I1282732,I3563,I1282345,I1282758,);
not I_75246 (I1282766,I1282758);
nand I_75247 (I1282783,I1282766,I1282444);
nor I_75248 (I1282800,I1282783,I476276);
DFFARX1 I_75249 (I1282800,I3563,I1282345,I1282313,);
nor I_75250 (I1282831,I1282766,I1282495);
nor I_75251 (I1282322,I1282639,I1282831);
not I_75252 (I1282889,I3570);
DFFARX1 I_75253 (I813697,I3563,I1282889,I1282915,);
nand I_75254 (I1282923,I1282915,I813691);
DFFARX1 I_75255 (I813694,I3563,I1282889,I1282949,);
DFFARX1 I_75256 (I1282949,I3563,I1282889,I1282966,);
not I_75257 (I1282881,I1282966);
not I_75258 (I1282988,I813700);
nor I_75259 (I1283005,I813700,I813694);
not I_75260 (I1283022,I813703);
nand I_75261 (I1283039,I1282988,I1283022);
nor I_75262 (I1283056,I813703,I813700);
and I_75263 (I1282860,I1283056,I1282923);
not I_75264 (I1283087,I813712);
nand I_75265 (I1283104,I1283087,I813706);
nor I_75266 (I1283121,I813712,I813709);
not I_75267 (I1283138,I1283121);
nand I_75268 (I1282863,I1283005,I1283138);
DFFARX1 I_75269 (I1283121,I3563,I1282889,I1282878,);
nor I_75270 (I1283183,I813691,I813703);
nor I_75271 (I1283200,I1283183,I813694);
and I_75272 (I1283217,I1283200,I1283104);
DFFARX1 I_75273 (I1283217,I3563,I1282889,I1282875,);
nor I_75274 (I1282872,I1283183,I1283039);
or I_75275 (I1282869,I1283121,I1283183);
nor I_75276 (I1283276,I813691,I813697);
DFFARX1 I_75277 (I1283276,I3563,I1282889,I1283302,);
not I_75278 (I1283310,I1283302);
nand I_75279 (I1283327,I1283310,I1282988);
nor I_75280 (I1283344,I1283327,I813694);
DFFARX1 I_75281 (I1283344,I3563,I1282889,I1282857,);
nor I_75282 (I1283375,I1283310,I1283039);
nor I_75283 (I1282866,I1283183,I1283375);
not I_75284 (I1283433,I3570);
DFFARX1 I_75285 (I1398195,I3563,I1283433,I1283459,);
nand I_75286 (I1283467,I1283459,I1398180);
DFFARX1 I_75287 (I1398174,I3563,I1283433,I1283493,);
DFFARX1 I_75288 (I1283493,I3563,I1283433,I1283510,);
not I_75289 (I1283425,I1283510);
not I_75290 (I1283532,I1398168);
nor I_75291 (I1283549,I1398168,I1398189);
not I_75292 (I1283566,I1398177);
nand I_75293 (I1283583,I1283532,I1283566);
nor I_75294 (I1283600,I1398177,I1398168);
and I_75295 (I1283404,I1283600,I1283467);
not I_75296 (I1283631,I1398186);
nand I_75297 (I1283648,I1283631,I1398192);
nor I_75298 (I1283665,I1398186,I1398183);
not I_75299 (I1283682,I1283665);
nand I_75300 (I1283407,I1283549,I1283682);
DFFARX1 I_75301 (I1283665,I3563,I1283433,I1283422,);
nor I_75302 (I1283727,I1398171,I1398177);
nor I_75303 (I1283744,I1283727,I1398189);
and I_75304 (I1283761,I1283744,I1283648);
DFFARX1 I_75305 (I1283761,I3563,I1283433,I1283419,);
nor I_75306 (I1283416,I1283727,I1283583);
or I_75307 (I1283413,I1283665,I1283727);
nor I_75308 (I1283820,I1398171,I1398168);
DFFARX1 I_75309 (I1283820,I3563,I1283433,I1283846,);
not I_75310 (I1283854,I1283846);
nand I_75311 (I1283871,I1283854,I1283532);
nor I_75312 (I1283888,I1283871,I1398189);
DFFARX1 I_75313 (I1283888,I3563,I1283433,I1283401,);
nor I_75314 (I1283919,I1283854,I1283583);
nor I_75315 (I1283410,I1283727,I1283919);
not I_75316 (I1283977,I3570);
DFFARX1 I_75317 (I678068,I3563,I1283977,I1284003,);
nand I_75318 (I1284011,I1284003,I678083);
DFFARX1 I_75319 (I678077,I3563,I1283977,I1284037,);
DFFARX1 I_75320 (I1284037,I3563,I1283977,I1284054,);
not I_75321 (I1283969,I1284054);
not I_75322 (I1284076,I678080);
nor I_75323 (I1284093,I678080,I678086);
not I_75324 (I1284110,I678068);
nand I_75325 (I1284127,I1284076,I1284110);
nor I_75326 (I1284144,I678068,I678080);
and I_75327 (I1283948,I1284144,I1284011);
not I_75328 (I1284175,I678065);
nand I_75329 (I1284192,I1284175,I678071);
nor I_75330 (I1284209,I678065,I678065);
not I_75331 (I1284226,I1284209);
nand I_75332 (I1283951,I1284093,I1284226);
DFFARX1 I_75333 (I1284209,I3563,I1283977,I1283966,);
nor I_75334 (I1284271,I678074,I678068);
nor I_75335 (I1284288,I1284271,I678086);
and I_75336 (I1284305,I1284288,I1284192);
DFFARX1 I_75337 (I1284305,I3563,I1283977,I1283963,);
nor I_75338 (I1283960,I1284271,I1284127);
or I_75339 (I1283957,I1284209,I1284271);
nor I_75340 (I1284364,I678074,I678089);
DFFARX1 I_75341 (I1284364,I3563,I1283977,I1284390,);
not I_75342 (I1284398,I1284390);
nand I_75343 (I1284415,I1284398,I1284076);
nor I_75344 (I1284432,I1284415,I678086);
DFFARX1 I_75345 (I1284432,I3563,I1283977,I1283945,);
nor I_75346 (I1284463,I1284398,I1284127);
nor I_75347 (I1283954,I1284271,I1284463);
not I_75348 (I1284521,I3570);
DFFARX1 I_75349 (I34522,I3563,I1284521,I1284547,);
nand I_75350 (I1284555,I1284547,I34516);
DFFARX1 I_75351 (I34537,I3563,I1284521,I1284581,);
DFFARX1 I_75352 (I1284581,I3563,I1284521,I1284598,);
not I_75353 (I1284513,I1284598);
not I_75354 (I1284620,I34525);
nor I_75355 (I1284637,I34525,I34534);
not I_75356 (I1284654,I34513);
nand I_75357 (I1284671,I1284620,I1284654);
nor I_75358 (I1284688,I34513,I34525);
and I_75359 (I1284492,I1284688,I1284555);
not I_75360 (I1284719,I34531);
nand I_75361 (I1284736,I1284719,I34519);
nor I_75362 (I1284753,I34531,I34513);
not I_75363 (I1284770,I1284753);
nand I_75364 (I1284495,I1284637,I1284770);
DFFARX1 I_75365 (I1284753,I3563,I1284521,I1284510,);
nor I_75366 (I1284815,I34516,I34513);
nor I_75367 (I1284832,I1284815,I34534);
and I_75368 (I1284849,I1284832,I1284736);
DFFARX1 I_75369 (I1284849,I3563,I1284521,I1284507,);
nor I_75370 (I1284504,I1284815,I1284671);
or I_75371 (I1284501,I1284753,I1284815);
nor I_75372 (I1284908,I34516,I34528);
DFFARX1 I_75373 (I1284908,I3563,I1284521,I1284934,);
not I_75374 (I1284942,I1284934);
nand I_75375 (I1284959,I1284942,I1284620);
nor I_75376 (I1284976,I1284959,I34534);
DFFARX1 I_75377 (I1284976,I3563,I1284521,I1284489,);
nor I_75378 (I1285007,I1284942,I1284671);
nor I_75379 (I1284498,I1284815,I1285007);
not I_75380 (I1285065,I3570);
DFFARX1 I_75381 (I584450,I3563,I1285065,I1285091,);
nand I_75382 (I1285099,I1285091,I584438);
DFFARX1 I_75383 (I584444,I3563,I1285065,I1285125,);
DFFARX1 I_75384 (I1285125,I3563,I1285065,I1285142,);
not I_75385 (I1285057,I1285142);
not I_75386 (I1285164,I584429);
nor I_75387 (I1285181,I584429,I584441);
not I_75388 (I1285198,I584432);
nand I_75389 (I1285215,I1285164,I1285198);
nor I_75390 (I1285232,I584432,I584429);
and I_75391 (I1285036,I1285232,I1285099);
not I_75392 (I1285263,I584447);
nand I_75393 (I1285280,I1285263,I584429);
nor I_75394 (I1285297,I584447,I584453);
not I_75395 (I1285314,I1285297);
nand I_75396 (I1285039,I1285181,I1285314);
DFFARX1 I_75397 (I1285297,I3563,I1285065,I1285054,);
nor I_75398 (I1285359,I584435,I584432);
nor I_75399 (I1285376,I1285359,I584441);
and I_75400 (I1285393,I1285376,I1285280);
DFFARX1 I_75401 (I1285393,I3563,I1285065,I1285051,);
nor I_75402 (I1285048,I1285359,I1285215);
or I_75403 (I1285045,I1285297,I1285359);
nor I_75404 (I1285452,I584435,I584432);
DFFARX1 I_75405 (I1285452,I3563,I1285065,I1285478,);
not I_75406 (I1285486,I1285478);
nand I_75407 (I1285503,I1285486,I1285164);
nor I_75408 (I1285520,I1285503,I584441);
DFFARX1 I_75409 (I1285520,I3563,I1285065,I1285033,);
nor I_75410 (I1285551,I1285486,I1285215);
nor I_75411 (I1285042,I1285359,I1285551);
not I_75412 (I1285609,I3570);
DFFARX1 I_75413 (I663040,I3563,I1285609,I1285635,);
nand I_75414 (I1285643,I1285635,I663055);
DFFARX1 I_75415 (I663049,I3563,I1285609,I1285669,);
DFFARX1 I_75416 (I1285669,I3563,I1285609,I1285686,);
not I_75417 (I1285601,I1285686);
not I_75418 (I1285708,I663052);
nor I_75419 (I1285725,I663052,I663058);
not I_75420 (I1285742,I663040);
nand I_75421 (I1285759,I1285708,I1285742);
nor I_75422 (I1285776,I663040,I663052);
and I_75423 (I1285580,I1285776,I1285643);
not I_75424 (I1285807,I663037);
nand I_75425 (I1285824,I1285807,I663043);
nor I_75426 (I1285841,I663037,I663037);
not I_75427 (I1285858,I1285841);
nand I_75428 (I1285583,I1285725,I1285858);
DFFARX1 I_75429 (I1285841,I3563,I1285609,I1285598,);
nor I_75430 (I1285903,I663046,I663040);
nor I_75431 (I1285920,I1285903,I663058);
and I_75432 (I1285937,I1285920,I1285824);
DFFARX1 I_75433 (I1285937,I3563,I1285609,I1285595,);
nor I_75434 (I1285592,I1285903,I1285759);
or I_75435 (I1285589,I1285841,I1285903);
nor I_75436 (I1285996,I663046,I663061);
DFFARX1 I_75437 (I1285996,I3563,I1285609,I1286022,);
not I_75438 (I1286030,I1286022);
nand I_75439 (I1286047,I1286030,I1285708);
nor I_75440 (I1286064,I1286047,I663058);
DFFARX1 I_75441 (I1286064,I3563,I1285609,I1285577,);
nor I_75442 (I1286095,I1286030,I1285759);
nor I_75443 (I1285586,I1285903,I1286095);
not I_75444 (I1286153,I3570);
DFFARX1 I_75445 (I1154599,I3563,I1286153,I1286179,);
nand I_75446 (I1286187,I1286179,I1154578);
DFFARX1 I_75447 (I1154575,I3563,I1286153,I1286213,);
DFFARX1 I_75448 (I1286213,I3563,I1286153,I1286230,);
not I_75449 (I1286145,I1286230);
not I_75450 (I1286252,I1154587);
nor I_75451 (I1286269,I1154587,I1154596);
not I_75452 (I1286286,I1154584);
nand I_75453 (I1286303,I1286252,I1286286);
nor I_75454 (I1286320,I1154584,I1154587);
and I_75455 (I1286124,I1286320,I1286187);
not I_75456 (I1286351,I1154593);
nand I_75457 (I1286368,I1286351,I1154590);
nor I_75458 (I1286385,I1154593,I1154575);
not I_75459 (I1286402,I1286385);
nand I_75460 (I1286127,I1286269,I1286402);
DFFARX1 I_75461 (I1286385,I3563,I1286153,I1286142,);
nor I_75462 (I1286447,I1154578,I1154584);
nor I_75463 (I1286464,I1286447,I1154596);
and I_75464 (I1286481,I1286464,I1286368);
DFFARX1 I_75465 (I1286481,I3563,I1286153,I1286139,);
nor I_75466 (I1286136,I1286447,I1286303);
or I_75467 (I1286133,I1286385,I1286447);
nor I_75468 (I1286540,I1154578,I1154581);
DFFARX1 I_75469 (I1286540,I3563,I1286153,I1286566,);
not I_75470 (I1286574,I1286566);
nand I_75471 (I1286591,I1286574,I1286252);
nor I_75472 (I1286608,I1286591,I1154596);
DFFARX1 I_75473 (I1286608,I3563,I1286153,I1286121,);
nor I_75474 (I1286639,I1286574,I1286303);
nor I_75475 (I1286130,I1286447,I1286639);
not I_75476 (I1286697,I3570);
DFFARX1 I_75477 (I1193325,I3563,I1286697,I1286723,);
nand I_75478 (I1286731,I1286723,I1193304);
DFFARX1 I_75479 (I1193301,I3563,I1286697,I1286757,);
DFFARX1 I_75480 (I1286757,I3563,I1286697,I1286774,);
not I_75481 (I1286689,I1286774);
not I_75482 (I1286796,I1193313);
nor I_75483 (I1286813,I1193313,I1193322);
not I_75484 (I1286830,I1193310);
nand I_75485 (I1286847,I1286796,I1286830);
nor I_75486 (I1286864,I1193310,I1193313);
and I_75487 (I1286668,I1286864,I1286731);
not I_75488 (I1286895,I1193319);
nand I_75489 (I1286912,I1286895,I1193316);
nor I_75490 (I1286929,I1193319,I1193301);
not I_75491 (I1286946,I1286929);
nand I_75492 (I1286671,I1286813,I1286946);
DFFARX1 I_75493 (I1286929,I3563,I1286697,I1286686,);
nor I_75494 (I1286991,I1193304,I1193310);
nor I_75495 (I1287008,I1286991,I1193322);
and I_75496 (I1287025,I1287008,I1286912);
DFFARX1 I_75497 (I1287025,I3563,I1286697,I1286683,);
nor I_75498 (I1286680,I1286991,I1286847);
or I_75499 (I1286677,I1286929,I1286991);
nor I_75500 (I1287084,I1193304,I1193307);
DFFARX1 I_75501 (I1287084,I3563,I1286697,I1287110,);
not I_75502 (I1287118,I1287110);
nand I_75503 (I1287135,I1287118,I1286796);
nor I_75504 (I1287152,I1287135,I1193322);
DFFARX1 I_75505 (I1287152,I3563,I1286697,I1286665,);
nor I_75506 (I1287183,I1287118,I1286847);
nor I_75507 (I1286674,I1286991,I1287183);
not I_75508 (I1287241,I3570);
DFFARX1 I_75509 (I638204,I3563,I1287241,I1287267,);
nand I_75510 (I1287275,I1287267,I638192);
DFFARX1 I_75511 (I638198,I3563,I1287241,I1287301,);
DFFARX1 I_75512 (I1287301,I3563,I1287241,I1287318,);
not I_75513 (I1287233,I1287318);
not I_75514 (I1287340,I638183);
nor I_75515 (I1287357,I638183,I638195);
not I_75516 (I1287374,I638186);
nand I_75517 (I1287391,I1287340,I1287374);
nor I_75518 (I1287408,I638186,I638183);
and I_75519 (I1287212,I1287408,I1287275);
not I_75520 (I1287439,I638201);
nand I_75521 (I1287456,I1287439,I638183);
nor I_75522 (I1287473,I638201,I638207);
not I_75523 (I1287490,I1287473);
nand I_75524 (I1287215,I1287357,I1287490);
DFFARX1 I_75525 (I1287473,I3563,I1287241,I1287230,);
nor I_75526 (I1287535,I638189,I638186);
nor I_75527 (I1287552,I1287535,I638195);
and I_75528 (I1287569,I1287552,I1287456);
DFFARX1 I_75529 (I1287569,I3563,I1287241,I1287227,);
nor I_75530 (I1287224,I1287535,I1287391);
or I_75531 (I1287221,I1287473,I1287535);
nor I_75532 (I1287628,I638189,I638186);
DFFARX1 I_75533 (I1287628,I3563,I1287241,I1287654,);
not I_75534 (I1287662,I1287654);
nand I_75535 (I1287679,I1287662,I1287340);
nor I_75536 (I1287696,I1287679,I638195);
DFFARX1 I_75537 (I1287696,I3563,I1287241,I1287209,);
nor I_75538 (I1287727,I1287662,I1287391);
nor I_75539 (I1287218,I1287535,I1287727);
not I_75540 (I1287785,I3570);
DFFARX1 I_75541 (I33465,I3563,I1287785,I1287811,);
nand I_75542 (I1287819,I1287811,I33459);
not I_75543 (I1287836,I1287819);
DFFARX1 I_75544 (I33477,I3563,I1287785,I1287862,);
not I_75545 (I1287870,I1287862);
not I_75546 (I1287887,I33480);
or I_75547 (I1287904,I33483,I33480);
nor I_75548 (I1287921,I33483,I33480);
or I_75549 (I1287938,I33468,I33483);
DFFARX1 I_75550 (I1287938,I3563,I1287785,I1287777,);
not I_75551 (I1287969,I33471);
nand I_75552 (I1287986,I1287969,I33474);
nand I_75553 (I1288003,I1287887,I1287986);
and I_75554 (I1287756,I1287870,I1288003);
nor I_75555 (I1288034,I33471,I33462);
and I_75556 (I1288051,I1287870,I1288034);
nor I_75557 (I1287762,I1287836,I1288051);
DFFARX1 I_75558 (I1288034,I3563,I1287785,I1288091,);
not I_75559 (I1288099,I1288091);
nor I_75560 (I1287771,I1287870,I1288099);
or I_75561 (I1288130,I1287938,I33462);
nor I_75562 (I1288147,I33462,I33468);
nand I_75563 (I1288164,I1288003,I1288147);
nand I_75564 (I1288181,I1288130,I1288164);
DFFARX1 I_75565 (I1288181,I3563,I1287785,I1287774,);
nor I_75566 (I1288212,I1288147,I1287904);
DFFARX1 I_75567 (I1288212,I3563,I1287785,I1287753,);
nor I_75568 (I1288243,I33462,I33459);
DFFARX1 I_75569 (I1288243,I3563,I1287785,I1288269,);
DFFARX1 I_75570 (I1288269,I3563,I1287785,I1287768,);
not I_75571 (I1288291,I1288269);
nand I_75572 (I1287765,I1288291,I1287819);
nand I_75573 (I1287759,I1288291,I1287921);
not I_75574 (I1288363,I3570);
DFFARX1 I_75575 (I72996,I3563,I1288363,I1288389,);
nand I_75576 (I1288397,I1288389,I72987);
not I_75577 (I1288414,I1288397);
DFFARX1 I_75578 (I72984,I3563,I1288363,I1288440,);
not I_75579 (I1288448,I1288440);
not I_75580 (I1288465,I72993);
or I_75581 (I1288482,I72984,I72993);
nor I_75582 (I1288499,I72984,I72993);
or I_75583 (I1288516,I72990,I72984);
DFFARX1 I_75584 (I1288516,I3563,I1288363,I1288355,);
not I_75585 (I1288547,I72999);
nand I_75586 (I1288564,I1288547,I73008);
nand I_75587 (I1288581,I1288465,I1288564);
and I_75588 (I1288334,I1288448,I1288581);
nor I_75589 (I1288612,I72999,I73002);
and I_75590 (I1288629,I1288448,I1288612);
nor I_75591 (I1288340,I1288414,I1288629);
DFFARX1 I_75592 (I1288612,I3563,I1288363,I1288669,);
not I_75593 (I1288677,I1288669);
nor I_75594 (I1288349,I1288448,I1288677);
or I_75595 (I1288708,I1288516,I72987);
nor I_75596 (I1288725,I72987,I72990);
nand I_75597 (I1288742,I1288581,I1288725);
nand I_75598 (I1288759,I1288708,I1288742);
DFFARX1 I_75599 (I1288759,I3563,I1288363,I1288352,);
nor I_75600 (I1288790,I1288725,I1288482);
DFFARX1 I_75601 (I1288790,I3563,I1288363,I1288331,);
nor I_75602 (I1288821,I72987,I73005);
DFFARX1 I_75603 (I1288821,I3563,I1288363,I1288847,);
DFFARX1 I_75604 (I1288847,I3563,I1288363,I1288346,);
not I_75605 (I1288869,I1288847);
nand I_75606 (I1288343,I1288869,I1288397);
nand I_75607 (I1288337,I1288869,I1288499);
not I_75608 (I1288941,I3570);
DFFARX1 I_75609 (I587900,I3563,I1288941,I1288967,);
nand I_75610 (I1288975,I1288967,I587915);
not I_75611 (I1288992,I1288975);
DFFARX1 I_75612 (I587897,I3563,I1288941,I1289018,);
not I_75613 (I1289026,I1289018);
not I_75614 (I1289043,I587906);
or I_75615 (I1289060,I587900,I587906);
nor I_75616 (I1289077,I587900,I587906);
or I_75617 (I1289094,I587897,I587900);
DFFARX1 I_75618 (I1289094,I3563,I1288941,I1288933,);
not I_75619 (I1289125,I587918);
nand I_75620 (I1289142,I1289125,I587921);
nand I_75621 (I1289159,I1289043,I1289142);
and I_75622 (I1288912,I1289026,I1289159);
nor I_75623 (I1289190,I587918,I587903);
and I_75624 (I1289207,I1289026,I1289190);
nor I_75625 (I1288918,I1288992,I1289207);
DFFARX1 I_75626 (I1289190,I3563,I1288941,I1289247,);
not I_75627 (I1289255,I1289247);
nor I_75628 (I1288927,I1289026,I1289255);
or I_75629 (I1289286,I1289094,I587909);
nor I_75630 (I1289303,I587909,I587897);
nand I_75631 (I1289320,I1289159,I1289303);
nand I_75632 (I1289337,I1289286,I1289320);
DFFARX1 I_75633 (I1289337,I3563,I1288941,I1288930,);
nor I_75634 (I1289368,I1289303,I1289060);
DFFARX1 I_75635 (I1289368,I3563,I1288941,I1288909,);
nor I_75636 (I1289399,I587909,I587912);
DFFARX1 I_75637 (I1289399,I3563,I1288941,I1289425,);
DFFARX1 I_75638 (I1289425,I3563,I1288941,I1288924,);
not I_75639 (I1289447,I1289425);
nand I_75640 (I1288921,I1289447,I1288975);
nand I_75641 (I1288915,I1289447,I1289077);
not I_75642 (I1289519,I3570);
DFFARX1 I_75643 (I232733,I3563,I1289519,I1289545,);
nand I_75644 (I1289553,I1289545,I232736);
not I_75645 (I1289570,I1289553);
DFFARX1 I_75646 (I232745,I3563,I1289519,I1289596,);
not I_75647 (I1289604,I1289596);
not I_75648 (I1289621,I232748);
or I_75649 (I1289638,I232739,I232748);
nor I_75650 (I1289655,I232739,I232748);
or I_75651 (I1289672,I232751,I232739);
DFFARX1 I_75652 (I1289672,I3563,I1289519,I1289511,);
not I_75653 (I1289703,I232736);
nand I_75654 (I1289720,I1289703,I232742);
nand I_75655 (I1289737,I1289621,I1289720);
and I_75656 (I1289490,I1289604,I1289737);
nor I_75657 (I1289768,I232736,I232754);
and I_75658 (I1289785,I1289604,I1289768);
nor I_75659 (I1289496,I1289570,I1289785);
DFFARX1 I_75660 (I1289768,I3563,I1289519,I1289825,);
not I_75661 (I1289833,I1289825);
nor I_75662 (I1289505,I1289604,I1289833);
or I_75663 (I1289864,I1289672,I232733);
nor I_75664 (I1289881,I232733,I232751);
nand I_75665 (I1289898,I1289737,I1289881);
nand I_75666 (I1289915,I1289864,I1289898);
DFFARX1 I_75667 (I1289915,I3563,I1289519,I1289508,);
nor I_75668 (I1289946,I1289881,I1289638);
DFFARX1 I_75669 (I1289946,I3563,I1289519,I1289487,);
nor I_75670 (I1289977,I232733,I232757);
DFFARX1 I_75671 (I1289977,I3563,I1289519,I1290003,);
DFFARX1 I_75672 (I1290003,I3563,I1289519,I1289502,);
not I_75673 (I1290025,I1290003);
nand I_75674 (I1289499,I1290025,I1289553);
nand I_75675 (I1289493,I1290025,I1289655);
not I_75676 (I1290097,I3570);
DFFARX1 I_75677 (I881150,I3563,I1290097,I1290123,);
nand I_75678 (I1290131,I1290123,I881150);
not I_75679 (I1290148,I1290131);
DFFARX1 I_75680 (I881156,I3563,I1290097,I1290174,);
not I_75681 (I1290182,I1290174);
not I_75682 (I1290199,I881168);
or I_75683 (I1290216,I881153,I881168);
nor I_75684 (I1290233,I881153,I881168);
or I_75685 (I1290250,I881147,I881153);
DFFARX1 I_75686 (I1290250,I3563,I1290097,I1290089,);
not I_75687 (I1290281,I881165);
nand I_75688 (I1290298,I1290281,I881159);
nand I_75689 (I1290315,I1290199,I1290298);
and I_75690 (I1290068,I1290182,I1290315);
nor I_75691 (I1290346,I881165,I881147);
and I_75692 (I1290363,I1290182,I1290346);
nor I_75693 (I1290074,I1290148,I1290363);
DFFARX1 I_75694 (I1290346,I3563,I1290097,I1290403,);
not I_75695 (I1290411,I1290403);
nor I_75696 (I1290083,I1290182,I1290411);
or I_75697 (I1290442,I1290250,I881162);
nor I_75698 (I1290459,I881162,I881147);
nand I_75699 (I1290476,I1290315,I1290459);
nand I_75700 (I1290493,I1290442,I1290476);
DFFARX1 I_75701 (I1290493,I3563,I1290097,I1290086,);
nor I_75702 (I1290524,I1290459,I1290216);
DFFARX1 I_75703 (I1290524,I3563,I1290097,I1290065,);
nor I_75704 (I1290555,I881162,I881153);
DFFARX1 I_75705 (I1290555,I3563,I1290097,I1290581,);
DFFARX1 I_75706 (I1290581,I3563,I1290097,I1290080,);
not I_75707 (I1290603,I1290581);
nand I_75708 (I1290077,I1290603,I1290131);
nand I_75709 (I1290071,I1290603,I1290233);
not I_75710 (I1290675,I3570);
DFFARX1 I_75711 (I76158,I3563,I1290675,I1290701,);
nand I_75712 (I1290709,I1290701,I76149);
not I_75713 (I1290726,I1290709);
DFFARX1 I_75714 (I76146,I3563,I1290675,I1290752,);
not I_75715 (I1290760,I1290752);
not I_75716 (I1290777,I76155);
or I_75717 (I1290794,I76146,I76155);
nor I_75718 (I1290811,I76146,I76155);
or I_75719 (I1290828,I76152,I76146);
DFFARX1 I_75720 (I1290828,I3563,I1290675,I1290667,);
not I_75721 (I1290859,I76161);
nand I_75722 (I1290876,I1290859,I76170);
nand I_75723 (I1290893,I1290777,I1290876);
and I_75724 (I1290646,I1290760,I1290893);
nor I_75725 (I1290924,I76161,I76164);
and I_75726 (I1290941,I1290760,I1290924);
nor I_75727 (I1290652,I1290726,I1290941);
DFFARX1 I_75728 (I1290924,I3563,I1290675,I1290981,);
not I_75729 (I1290989,I1290981);
nor I_75730 (I1290661,I1290760,I1290989);
or I_75731 (I1291020,I1290828,I76149);
nor I_75732 (I1291037,I76149,I76152);
nand I_75733 (I1291054,I1290893,I1291037);
nand I_75734 (I1291071,I1291020,I1291054);
DFFARX1 I_75735 (I1291071,I3563,I1290675,I1290664,);
nor I_75736 (I1291102,I1291037,I1290794);
DFFARX1 I_75737 (I1291102,I3563,I1290675,I1290643,);
nor I_75738 (I1291133,I76149,I76167);
DFFARX1 I_75739 (I1291133,I3563,I1290675,I1291159,);
DFFARX1 I_75740 (I1291159,I3563,I1290675,I1290658,);
not I_75741 (I1291181,I1291159);
nand I_75742 (I1290655,I1291181,I1290709);
nand I_75743 (I1290649,I1291181,I1290811);
not I_75744 (I1291253,I3570);
DFFARX1 I_75745 (I855854,I3563,I1291253,I1291279,);
nand I_75746 (I1291287,I1291279,I855854);
not I_75747 (I1291304,I1291287);
DFFARX1 I_75748 (I855860,I3563,I1291253,I1291330,);
not I_75749 (I1291338,I1291330);
not I_75750 (I1291355,I855872);
or I_75751 (I1291372,I855857,I855872);
nor I_75752 (I1291389,I855857,I855872);
or I_75753 (I1291406,I855851,I855857);
DFFARX1 I_75754 (I1291406,I3563,I1291253,I1291245,);
not I_75755 (I1291437,I855869);
nand I_75756 (I1291454,I1291437,I855863);
nand I_75757 (I1291471,I1291355,I1291454);
and I_75758 (I1291224,I1291338,I1291471);
nor I_75759 (I1291502,I855869,I855851);
and I_75760 (I1291519,I1291338,I1291502);
nor I_75761 (I1291230,I1291304,I1291519);
DFFARX1 I_75762 (I1291502,I3563,I1291253,I1291559,);
not I_75763 (I1291567,I1291559);
nor I_75764 (I1291239,I1291338,I1291567);
or I_75765 (I1291598,I1291406,I855866);
nor I_75766 (I1291615,I855866,I855851);
nand I_75767 (I1291632,I1291471,I1291615);
nand I_75768 (I1291649,I1291598,I1291632);
DFFARX1 I_75769 (I1291649,I3563,I1291253,I1291242,);
nor I_75770 (I1291680,I1291615,I1291372);
DFFARX1 I_75771 (I1291680,I3563,I1291253,I1291221,);
nor I_75772 (I1291711,I855866,I855857);
DFFARX1 I_75773 (I1291711,I3563,I1291253,I1291737,);
DFFARX1 I_75774 (I1291737,I3563,I1291253,I1291236,);
not I_75775 (I1291759,I1291737);
nand I_75776 (I1291233,I1291759,I1291287);
nand I_75777 (I1291227,I1291759,I1291389);
not I_75778 (I1291831,I3570);
DFFARX1 I_75779 (I1384507,I3563,I1291831,I1291857,);
nand I_75780 (I1291865,I1291857,I1384498);
not I_75781 (I1291882,I1291865);
DFFARX1 I_75782 (I1384483,I3563,I1291831,I1291908,);
not I_75783 (I1291916,I1291908);
not I_75784 (I1291933,I1384486);
or I_75785 (I1291950,I1384495,I1384486);
nor I_75786 (I1291967,I1384495,I1384486);
or I_75787 (I1291984,I1384492,I1384495);
DFFARX1 I_75788 (I1291984,I3563,I1291831,I1291823,);
not I_75789 (I1292015,I1384504);
nand I_75790 (I1292032,I1292015,I1384483);
nand I_75791 (I1292049,I1291933,I1292032);
and I_75792 (I1291802,I1291916,I1292049);
nor I_75793 (I1292080,I1384504,I1384489);
and I_75794 (I1292097,I1291916,I1292080);
nor I_75795 (I1291808,I1291882,I1292097);
DFFARX1 I_75796 (I1292080,I3563,I1291831,I1292137,);
not I_75797 (I1292145,I1292137);
nor I_75798 (I1291817,I1291916,I1292145);
or I_75799 (I1292176,I1291984,I1384510);
nor I_75800 (I1292193,I1384510,I1384492);
nand I_75801 (I1292210,I1292049,I1292193);
nand I_75802 (I1292227,I1292176,I1292210);
DFFARX1 I_75803 (I1292227,I3563,I1291831,I1291820,);
nor I_75804 (I1292258,I1292193,I1291950);
DFFARX1 I_75805 (I1292258,I3563,I1291831,I1291799,);
nor I_75806 (I1292289,I1384510,I1384501);
DFFARX1 I_75807 (I1292289,I3563,I1291831,I1292315,);
DFFARX1 I_75808 (I1292315,I3563,I1291831,I1291814,);
not I_75809 (I1292337,I1292315);
nand I_75810 (I1291811,I1292337,I1291865);
nand I_75811 (I1291805,I1292337,I1291967);
not I_75812 (I1292409,I3570);
DFFARX1 I_75813 (I1206035,I3563,I1292409,I1292435,);
nand I_75814 (I1292443,I1292435,I1206020);
not I_75815 (I1292460,I1292443);
DFFARX1 I_75816 (I1206023,I3563,I1292409,I1292486,);
not I_75817 (I1292494,I1292486);
not I_75818 (I1292511,I1206038);
or I_75819 (I1292528,I1206041,I1206038);
nor I_75820 (I1292545,I1206041,I1206038);
or I_75821 (I1292562,I1206017,I1206041);
DFFARX1 I_75822 (I1292562,I3563,I1292409,I1292401,);
not I_75823 (I1292593,I1206029);
nand I_75824 (I1292610,I1292593,I1206032);
nand I_75825 (I1292627,I1292511,I1292610);
and I_75826 (I1292380,I1292494,I1292627);
nor I_75827 (I1292658,I1206029,I1206026);
and I_75828 (I1292675,I1292494,I1292658);
nor I_75829 (I1292386,I1292460,I1292675);
DFFARX1 I_75830 (I1292658,I3563,I1292409,I1292715,);
not I_75831 (I1292723,I1292715);
nor I_75832 (I1292395,I1292494,I1292723);
or I_75833 (I1292754,I1292562,I1206017);
nor I_75834 (I1292771,I1206017,I1206017);
nand I_75835 (I1292788,I1292627,I1292771);
nand I_75836 (I1292805,I1292754,I1292788);
DFFARX1 I_75837 (I1292805,I3563,I1292409,I1292398,);
nor I_75838 (I1292836,I1292771,I1292528);
DFFARX1 I_75839 (I1292836,I3563,I1292409,I1292377,);
nor I_75840 (I1292867,I1206017,I1206020);
DFFARX1 I_75841 (I1292867,I3563,I1292409,I1292893,);
DFFARX1 I_75842 (I1292893,I3563,I1292409,I1292392,);
not I_75843 (I1292915,I1292893);
nand I_75844 (I1292389,I1292915,I1292443);
nand I_75845 (I1292383,I1292915,I1292545);
not I_75846 (I1292987,I3570);
DFFARX1 I_75847 (I822653,I3563,I1292987,I1293013,);
nand I_75848 (I1293021,I1293013,I822653);
not I_75849 (I1293038,I1293021);
DFFARX1 I_75850 (I822659,I3563,I1292987,I1293064,);
not I_75851 (I1293072,I1293064);
not I_75852 (I1293089,I822671);
or I_75853 (I1293106,I822656,I822671);
nor I_75854 (I1293123,I822656,I822671);
or I_75855 (I1293140,I822650,I822656);
DFFARX1 I_75856 (I1293140,I3563,I1292987,I1292979,);
not I_75857 (I1293171,I822668);
nand I_75858 (I1293188,I1293171,I822662);
nand I_75859 (I1293205,I1293089,I1293188);
and I_75860 (I1292958,I1293072,I1293205);
nor I_75861 (I1293236,I822668,I822650);
and I_75862 (I1293253,I1293072,I1293236);
nor I_75863 (I1292964,I1293038,I1293253);
DFFARX1 I_75864 (I1293236,I3563,I1292987,I1293293,);
not I_75865 (I1293301,I1293293);
nor I_75866 (I1292973,I1293072,I1293301);
or I_75867 (I1293332,I1293140,I822665);
nor I_75868 (I1293349,I822665,I822650);
nand I_75869 (I1293366,I1293205,I1293349);
nand I_75870 (I1293383,I1293332,I1293366);
DFFARX1 I_75871 (I1293383,I3563,I1292987,I1292976,);
nor I_75872 (I1293414,I1293349,I1293106);
DFFARX1 I_75873 (I1293414,I3563,I1292987,I1292955,);
nor I_75874 (I1293445,I822665,I822656);
DFFARX1 I_75875 (I1293445,I3563,I1292987,I1293471,);
DFFARX1 I_75876 (I1293471,I3563,I1292987,I1292970,);
not I_75877 (I1293493,I1293471);
nand I_75878 (I1292967,I1293493,I1293021);
nand I_75879 (I1292961,I1293493,I1293123);
not I_75880 (I1293565,I3570);
DFFARX1 I_75881 (I1268728,I3563,I1293565,I1293591,);
nand I_75882 (I1293599,I1293591,I1268737);
not I_75883 (I1293616,I1293599);
DFFARX1 I_75884 (I1268713,I3563,I1293565,I1293642,);
not I_75885 (I1293650,I1293642);
not I_75886 (I1293667,I1268716);
or I_75887 (I1293684,I1268713,I1268716);
nor I_75888 (I1293701,I1268713,I1268716);
or I_75889 (I1293718,I1268731,I1268713);
DFFARX1 I_75890 (I1293718,I3563,I1293565,I1293557,);
not I_75891 (I1293749,I1268719);
nand I_75892 (I1293766,I1293749,I1268734);
nand I_75893 (I1293783,I1293667,I1293766);
and I_75894 (I1293536,I1293650,I1293783);
nor I_75895 (I1293814,I1268719,I1268722);
and I_75896 (I1293831,I1293650,I1293814);
nor I_75897 (I1293542,I1293616,I1293831);
DFFARX1 I_75898 (I1293814,I3563,I1293565,I1293871,);
not I_75899 (I1293879,I1293871);
nor I_75900 (I1293551,I1293650,I1293879);
or I_75901 (I1293910,I1293718,I1268725);
nor I_75902 (I1293927,I1268725,I1268731);
nand I_75903 (I1293944,I1293783,I1293927);
nand I_75904 (I1293961,I1293910,I1293944);
DFFARX1 I_75905 (I1293961,I3563,I1293565,I1293554,);
nor I_75906 (I1293992,I1293927,I1293684);
DFFARX1 I_75907 (I1293992,I3563,I1293565,I1293533,);
nor I_75908 (I1294023,I1268725,I1268716);
DFFARX1 I_75909 (I1294023,I3563,I1293565,I1294049,);
DFFARX1 I_75910 (I1294049,I3563,I1293565,I1293548,);
not I_75911 (I1294071,I1294049);
nand I_75912 (I1293545,I1294071,I1293599);
nand I_75913 (I1293539,I1294071,I1293701);
not I_75914 (I1294143,I3570);
DFFARX1 I_75915 (I101454,I3563,I1294143,I1294169,);
nand I_75916 (I1294177,I1294169,I101445);
not I_75917 (I1294194,I1294177);
DFFARX1 I_75918 (I101442,I3563,I1294143,I1294220,);
not I_75919 (I1294228,I1294220);
not I_75920 (I1294245,I101451);
or I_75921 (I1294262,I101442,I101451);
nor I_75922 (I1294279,I101442,I101451);
or I_75923 (I1294296,I101448,I101442);
DFFARX1 I_75924 (I1294296,I3563,I1294143,I1294135,);
not I_75925 (I1294327,I101457);
nand I_75926 (I1294344,I1294327,I101466);
nand I_75927 (I1294361,I1294245,I1294344);
and I_75928 (I1294114,I1294228,I1294361);
nor I_75929 (I1294392,I101457,I101460);
and I_75930 (I1294409,I1294228,I1294392);
nor I_75931 (I1294120,I1294194,I1294409);
DFFARX1 I_75932 (I1294392,I3563,I1294143,I1294449,);
not I_75933 (I1294457,I1294449);
nor I_75934 (I1294129,I1294228,I1294457);
or I_75935 (I1294488,I1294296,I101445);
nor I_75936 (I1294505,I101445,I101448);
nand I_75937 (I1294522,I1294361,I1294505);
nand I_75938 (I1294539,I1294488,I1294522);
DFFARX1 I_75939 (I1294539,I3563,I1294143,I1294132,);
nor I_75940 (I1294570,I1294505,I1294262);
DFFARX1 I_75941 (I1294570,I3563,I1294143,I1294111,);
nor I_75942 (I1294601,I101445,I101463);
DFFARX1 I_75943 (I1294601,I3563,I1294143,I1294627,);
DFFARX1 I_75944 (I1294627,I3563,I1294143,I1294126,);
not I_75945 (I1294649,I1294627);
nand I_75946 (I1294123,I1294649,I1294177);
nand I_75947 (I1294117,I1294649,I1294279);
not I_75948 (I1294721,I3570);
DFFARX1 I_75949 (I575096,I3563,I1294721,I1294747,);
nand I_75950 (I1294755,I1294747,I575105);
not I_75951 (I1294772,I1294755);
DFFARX1 I_75952 (I575117,I3563,I1294721,I1294798,);
not I_75953 (I1294806,I1294798);
not I_75954 (I1294823,I575108);
or I_75955 (I1294840,I575102,I575108);
nor I_75956 (I1294857,I575102,I575108);
or I_75957 (I1294874,I575096,I575102);
DFFARX1 I_75958 (I1294874,I3563,I1294721,I1294713,);
not I_75959 (I1294905,I575099);
nand I_75960 (I1294922,I1294905,I575111);
nand I_75961 (I1294939,I1294823,I1294922);
and I_75962 (I1294692,I1294806,I1294939);
nor I_75963 (I1294970,I575099,I575120);
and I_75964 (I1294987,I1294806,I1294970);
nor I_75965 (I1294698,I1294772,I1294987);
DFFARX1 I_75966 (I1294970,I3563,I1294721,I1295027,);
not I_75967 (I1295035,I1295027);
nor I_75968 (I1294707,I1294806,I1295035);
or I_75969 (I1295066,I1294874,I575114);
nor I_75970 (I1295083,I575114,I575096);
nand I_75971 (I1295100,I1294939,I1295083);
nand I_75972 (I1295117,I1295066,I1295100);
DFFARX1 I_75973 (I1295117,I3563,I1294721,I1294710,);
nor I_75974 (I1295148,I1295083,I1294840);
DFFARX1 I_75975 (I1295148,I3563,I1294721,I1294689,);
nor I_75976 (I1295179,I575114,I575099);
DFFARX1 I_75977 (I1295179,I3563,I1294721,I1295205,);
DFFARX1 I_75978 (I1295205,I3563,I1294721,I1294704,);
not I_75979 (I1295227,I1295205);
nand I_75980 (I1294701,I1295227,I1294755);
nand I_75981 (I1294695,I1295227,I1294857);
not I_75982 (I1295299,I3570);
DFFARX1 I_75983 (I1222219,I3563,I1295299,I1295325,);
nand I_75984 (I1295333,I1295325,I1222204);
not I_75985 (I1295350,I1295333);
DFFARX1 I_75986 (I1222207,I3563,I1295299,I1295376,);
not I_75987 (I1295384,I1295376);
not I_75988 (I1295401,I1222222);
or I_75989 (I1295418,I1222225,I1222222);
nor I_75990 (I1295435,I1222225,I1222222);
or I_75991 (I1295452,I1222201,I1222225);
DFFARX1 I_75992 (I1295452,I3563,I1295299,I1295291,);
not I_75993 (I1295483,I1222213);
nand I_75994 (I1295500,I1295483,I1222216);
nand I_75995 (I1295517,I1295401,I1295500);
and I_75996 (I1295270,I1295384,I1295517);
nor I_75997 (I1295548,I1222213,I1222210);
and I_75998 (I1295565,I1295384,I1295548);
nor I_75999 (I1295276,I1295350,I1295565);
DFFARX1 I_76000 (I1295548,I3563,I1295299,I1295605,);
not I_76001 (I1295613,I1295605);
nor I_76002 (I1295285,I1295384,I1295613);
or I_76003 (I1295644,I1295452,I1222201);
nor I_76004 (I1295661,I1222201,I1222201);
nand I_76005 (I1295678,I1295517,I1295661);
nand I_76006 (I1295695,I1295644,I1295678);
DFFARX1 I_76007 (I1295695,I3563,I1295299,I1295288,);
nor I_76008 (I1295726,I1295661,I1295418);
DFFARX1 I_76009 (I1295726,I3563,I1295299,I1295267,);
nor I_76010 (I1295757,I1222201,I1222204);
DFFARX1 I_76011 (I1295757,I3563,I1295299,I1295783,);
DFFARX1 I_76012 (I1295783,I3563,I1295299,I1295282,);
not I_76013 (I1295805,I1295783);
nand I_76014 (I1295279,I1295805,I1295333);
nand I_76015 (I1295273,I1295805,I1295435);
not I_76016 (I1295877,I3570);
DFFARX1 I_76017 (I251773,I3563,I1295877,I1295903,);
nand I_76018 (I1295911,I1295903,I251776);
not I_76019 (I1295928,I1295911);
DFFARX1 I_76020 (I251785,I3563,I1295877,I1295954,);
not I_76021 (I1295962,I1295954);
not I_76022 (I1295979,I251788);
or I_76023 (I1295996,I251779,I251788);
nor I_76024 (I1296013,I251779,I251788);
or I_76025 (I1296030,I251791,I251779);
DFFARX1 I_76026 (I1296030,I3563,I1295877,I1295869,);
not I_76027 (I1296061,I251776);
nand I_76028 (I1296078,I1296061,I251782);
nand I_76029 (I1296095,I1295979,I1296078);
and I_76030 (I1295848,I1295962,I1296095);
nor I_76031 (I1296126,I251776,I251794);
and I_76032 (I1296143,I1295962,I1296126);
nor I_76033 (I1295854,I1295928,I1296143);
DFFARX1 I_76034 (I1296126,I3563,I1295877,I1296183,);
not I_76035 (I1296191,I1296183);
nor I_76036 (I1295863,I1295962,I1296191);
or I_76037 (I1296222,I1296030,I251773);
nor I_76038 (I1296239,I251773,I251791);
nand I_76039 (I1296256,I1296095,I1296239);
nand I_76040 (I1296273,I1296222,I1296256);
DFFARX1 I_76041 (I1296273,I3563,I1295877,I1295866,);
nor I_76042 (I1296304,I1296239,I1295996);
DFFARX1 I_76043 (I1296304,I3563,I1295877,I1295845,);
nor I_76044 (I1296335,I251773,I251797);
DFFARX1 I_76045 (I1296335,I3563,I1295877,I1296361,);
DFFARX1 I_76046 (I1296361,I3563,I1295877,I1295860,);
not I_76047 (I1296383,I1296361);
nand I_76048 (I1295857,I1296383,I1295911);
nand I_76049 (I1295851,I1296383,I1296013);
not I_76050 (I1296455,I3570);
DFFARX1 I_76051 (I244633,I3563,I1296455,I1296481,);
nand I_76052 (I1296489,I1296481,I244636);
not I_76053 (I1296506,I1296489);
DFFARX1 I_76054 (I244645,I3563,I1296455,I1296532,);
not I_76055 (I1296540,I1296532);
not I_76056 (I1296557,I244648);
or I_76057 (I1296574,I244639,I244648);
nor I_76058 (I1296591,I244639,I244648);
or I_76059 (I1296608,I244651,I244639);
DFFARX1 I_76060 (I1296608,I3563,I1296455,I1296447,);
not I_76061 (I1296639,I244636);
nand I_76062 (I1296656,I1296639,I244642);
nand I_76063 (I1296673,I1296557,I1296656);
and I_76064 (I1296426,I1296540,I1296673);
nor I_76065 (I1296704,I244636,I244654);
and I_76066 (I1296721,I1296540,I1296704);
nor I_76067 (I1296432,I1296506,I1296721);
DFFARX1 I_76068 (I1296704,I3563,I1296455,I1296761,);
not I_76069 (I1296769,I1296761);
nor I_76070 (I1296441,I1296540,I1296769);
or I_76071 (I1296800,I1296608,I244633);
nor I_76072 (I1296817,I244633,I244651);
nand I_76073 (I1296834,I1296673,I1296817);
nand I_76074 (I1296851,I1296800,I1296834);
DFFARX1 I_76075 (I1296851,I3563,I1296455,I1296444,);
nor I_76076 (I1296882,I1296817,I1296574);
DFFARX1 I_76077 (I1296882,I3563,I1296455,I1296423,);
nor I_76078 (I1296913,I244633,I244657);
DFFARX1 I_76079 (I1296913,I3563,I1296455,I1296939,);
DFFARX1 I_76080 (I1296939,I3563,I1296455,I1296438,);
not I_76081 (I1296961,I1296939);
nand I_76082 (I1296435,I1296961,I1296489);
nand I_76083 (I1296429,I1296961,I1296591);
not I_76084 (I1297033,I3570);
DFFARX1 I_76085 (I155208,I3563,I1297033,I1297059,);
nand I_76086 (I1297067,I1297059,I155199);
not I_76087 (I1297084,I1297067);
DFFARX1 I_76088 (I155196,I3563,I1297033,I1297110,);
not I_76089 (I1297118,I1297110);
not I_76090 (I1297135,I155205);
or I_76091 (I1297152,I155196,I155205);
nor I_76092 (I1297169,I155196,I155205);
or I_76093 (I1297186,I155202,I155196);
DFFARX1 I_76094 (I1297186,I3563,I1297033,I1297025,);
not I_76095 (I1297217,I155211);
nand I_76096 (I1297234,I1297217,I155220);
nand I_76097 (I1297251,I1297135,I1297234);
and I_76098 (I1297004,I1297118,I1297251);
nor I_76099 (I1297282,I155211,I155214);
and I_76100 (I1297299,I1297118,I1297282);
nor I_76101 (I1297010,I1297084,I1297299);
DFFARX1 I_76102 (I1297282,I3563,I1297033,I1297339,);
not I_76103 (I1297347,I1297339);
nor I_76104 (I1297019,I1297118,I1297347);
or I_76105 (I1297378,I1297186,I155199);
nor I_76106 (I1297395,I155199,I155202);
nand I_76107 (I1297412,I1297251,I1297395);
nand I_76108 (I1297429,I1297378,I1297412);
DFFARX1 I_76109 (I1297429,I3563,I1297033,I1297022,);
nor I_76110 (I1297460,I1297395,I1297152);
DFFARX1 I_76111 (I1297460,I3563,I1297033,I1297001,);
nor I_76112 (I1297491,I155199,I155217);
DFFARX1 I_76113 (I1297491,I3563,I1297033,I1297517,);
DFFARX1 I_76114 (I1297517,I3563,I1297033,I1297016,);
not I_76115 (I1297539,I1297517);
nand I_76116 (I1297013,I1297539,I1297067);
nand I_76117 (I1297007,I1297539,I1297169);
not I_76118 (I1297611,I3570);
DFFARX1 I_76119 (I904865,I3563,I1297611,I1297637,);
nand I_76120 (I1297645,I1297637,I904865);
not I_76121 (I1297662,I1297645);
DFFARX1 I_76122 (I904871,I3563,I1297611,I1297688,);
not I_76123 (I1297696,I1297688);
not I_76124 (I1297713,I904883);
or I_76125 (I1297730,I904868,I904883);
nor I_76126 (I1297747,I904868,I904883);
or I_76127 (I1297764,I904862,I904868);
DFFARX1 I_76128 (I1297764,I3563,I1297611,I1297603,);
not I_76129 (I1297795,I904880);
nand I_76130 (I1297812,I1297795,I904874);
nand I_76131 (I1297829,I1297713,I1297812);
and I_76132 (I1297582,I1297696,I1297829);
nor I_76133 (I1297860,I904880,I904862);
and I_76134 (I1297877,I1297696,I1297860);
nor I_76135 (I1297588,I1297662,I1297877);
DFFARX1 I_76136 (I1297860,I3563,I1297611,I1297917,);
not I_76137 (I1297925,I1297917);
nor I_76138 (I1297597,I1297696,I1297925);
or I_76139 (I1297956,I1297764,I904877);
nor I_76140 (I1297973,I904877,I904862);
nand I_76141 (I1297990,I1297829,I1297973);
nand I_76142 (I1298007,I1297956,I1297990);
DFFARX1 I_76143 (I1298007,I3563,I1297611,I1297600,);
nor I_76144 (I1298038,I1297973,I1297730);
DFFARX1 I_76145 (I1298038,I3563,I1297611,I1297579,);
nor I_76146 (I1298069,I904877,I904868);
DFFARX1 I_76147 (I1298069,I3563,I1297611,I1298095,);
DFFARX1 I_76148 (I1298095,I3563,I1297611,I1297594,);
not I_76149 (I1298117,I1298095);
nand I_76150 (I1297591,I1298117,I1297645);
nand I_76151 (I1297585,I1298117,I1297747);
not I_76152 (I1298189,I3570);
DFFARX1 I_76153 (I859016,I3563,I1298189,I1298215,);
nand I_76154 (I1298223,I1298215,I859016);
not I_76155 (I1298240,I1298223);
DFFARX1 I_76156 (I859022,I3563,I1298189,I1298266,);
not I_76157 (I1298274,I1298266);
not I_76158 (I1298291,I859034);
or I_76159 (I1298308,I859019,I859034);
nor I_76160 (I1298325,I859019,I859034);
or I_76161 (I1298342,I859013,I859019);
DFFARX1 I_76162 (I1298342,I3563,I1298189,I1298181,);
not I_76163 (I1298373,I859031);
nand I_76164 (I1298390,I1298373,I859025);
nand I_76165 (I1298407,I1298291,I1298390);
and I_76166 (I1298160,I1298274,I1298407);
nor I_76167 (I1298438,I859031,I859013);
and I_76168 (I1298455,I1298274,I1298438);
nor I_76169 (I1298166,I1298240,I1298455);
DFFARX1 I_76170 (I1298438,I3563,I1298189,I1298495,);
not I_76171 (I1298503,I1298495);
nor I_76172 (I1298175,I1298274,I1298503);
or I_76173 (I1298534,I1298342,I859028);
nor I_76174 (I1298551,I859028,I859013);
nand I_76175 (I1298568,I1298407,I1298551);
nand I_76176 (I1298585,I1298534,I1298568);
DFFARX1 I_76177 (I1298585,I3563,I1298189,I1298178,);
nor I_76178 (I1298616,I1298551,I1298308);
DFFARX1 I_76179 (I1298616,I3563,I1298189,I1298157,);
nor I_76180 (I1298647,I859028,I859019);
DFFARX1 I_76181 (I1298647,I3563,I1298189,I1298673,);
DFFARX1 I_76182 (I1298673,I3563,I1298189,I1298172,);
not I_76183 (I1298695,I1298673);
nand I_76184 (I1298169,I1298695,I1298223);
nand I_76185 (I1298163,I1298695,I1298325);
not I_76186 (I1298767,I3570);
DFFARX1 I_76187 (I927801,I3563,I1298767,I1298793,);
nand I_76188 (I1298801,I1298793,I927822);
not I_76189 (I1298818,I1298801);
DFFARX1 I_76190 (I927795,I3563,I1298767,I1298844,);
not I_76191 (I1298852,I1298844);
not I_76192 (I1298869,I927816);
or I_76193 (I1298886,I927807,I927816);
nor I_76194 (I1298903,I927807,I927816);
or I_76195 (I1298920,I927810,I927807);
DFFARX1 I_76196 (I1298920,I3563,I1298767,I1298759,);
not I_76197 (I1298951,I927798);
nand I_76198 (I1298968,I1298951,I927813);
nand I_76199 (I1298985,I1298869,I1298968);
and I_76200 (I1298738,I1298852,I1298985);
nor I_76201 (I1299016,I927798,I927795);
and I_76202 (I1299033,I1298852,I1299016);
nor I_76203 (I1298744,I1298818,I1299033);
DFFARX1 I_76204 (I1299016,I3563,I1298767,I1299073,);
not I_76205 (I1299081,I1299073);
nor I_76206 (I1298753,I1298852,I1299081);
or I_76207 (I1299112,I1298920,I927819);
nor I_76208 (I1299129,I927819,I927810);
nand I_76209 (I1299146,I1298985,I1299129);
nand I_76210 (I1299163,I1299112,I1299146);
DFFARX1 I_76211 (I1299163,I3563,I1298767,I1298756,);
nor I_76212 (I1299194,I1299129,I1298886);
DFFARX1 I_76213 (I1299194,I3563,I1298767,I1298735,);
nor I_76214 (I1299225,I927819,I927804);
DFFARX1 I_76215 (I1299225,I3563,I1298767,I1299251,);
DFFARX1 I_76216 (I1299251,I3563,I1298767,I1298750,);
not I_76217 (I1299273,I1299251);
nand I_76218 (I1298747,I1299273,I1298801);
nand I_76219 (I1298741,I1299273,I1298903);
not I_76220 (I1299345,I3570);
DFFARX1 I_76221 (I1227421,I3563,I1299345,I1299371,);
nand I_76222 (I1299379,I1299371,I1227406);
not I_76223 (I1299396,I1299379);
DFFARX1 I_76224 (I1227409,I3563,I1299345,I1299422,);
not I_76225 (I1299430,I1299422);
not I_76226 (I1299447,I1227424);
or I_76227 (I1299464,I1227427,I1227424);
nor I_76228 (I1299481,I1227427,I1227424);
or I_76229 (I1299498,I1227403,I1227427);
DFFARX1 I_76230 (I1299498,I3563,I1299345,I1299337,);
not I_76231 (I1299529,I1227415);
nand I_76232 (I1299546,I1299529,I1227418);
nand I_76233 (I1299563,I1299447,I1299546);
and I_76234 (I1299316,I1299430,I1299563);
nor I_76235 (I1299594,I1227415,I1227412);
and I_76236 (I1299611,I1299430,I1299594);
nor I_76237 (I1299322,I1299396,I1299611);
DFFARX1 I_76238 (I1299594,I3563,I1299345,I1299651,);
not I_76239 (I1299659,I1299651);
nor I_76240 (I1299331,I1299430,I1299659);
or I_76241 (I1299690,I1299498,I1227403);
nor I_76242 (I1299707,I1227403,I1227403);
nand I_76243 (I1299724,I1299563,I1299707);
nand I_76244 (I1299741,I1299690,I1299724);
DFFARX1 I_76245 (I1299741,I3563,I1299345,I1299334,);
nor I_76246 (I1299772,I1299707,I1299464);
DFFARX1 I_76247 (I1299772,I3563,I1299345,I1299313,);
nor I_76248 (I1299803,I1227403,I1227406);
DFFARX1 I_76249 (I1299803,I3563,I1299345,I1299829,);
DFFARX1 I_76250 (I1299829,I3563,I1299345,I1299328,);
not I_76251 (I1299851,I1299829);
nand I_76252 (I1299325,I1299851,I1299379);
nand I_76253 (I1299319,I1299851,I1299481);
not I_76254 (I1299923,I3570);
DFFARX1 I_76255 (I842679,I3563,I1299923,I1299949,);
nand I_76256 (I1299957,I1299949,I842679);
not I_76257 (I1299974,I1299957);
DFFARX1 I_76258 (I842685,I3563,I1299923,I1300000,);
not I_76259 (I1300008,I1300000);
not I_76260 (I1300025,I842697);
or I_76261 (I1300042,I842682,I842697);
nor I_76262 (I1300059,I842682,I842697);
or I_76263 (I1300076,I842676,I842682);
DFFARX1 I_76264 (I1300076,I3563,I1299923,I1299915,);
not I_76265 (I1300107,I842694);
nand I_76266 (I1300124,I1300107,I842688);
nand I_76267 (I1300141,I1300025,I1300124);
and I_76268 (I1299894,I1300008,I1300141);
nor I_76269 (I1300172,I842694,I842676);
and I_76270 (I1300189,I1300008,I1300172);
nor I_76271 (I1299900,I1299974,I1300189);
DFFARX1 I_76272 (I1300172,I3563,I1299923,I1300229,);
not I_76273 (I1300237,I1300229);
nor I_76274 (I1299909,I1300008,I1300237);
or I_76275 (I1300268,I1300076,I842691);
nor I_76276 (I1300285,I842691,I842676);
nand I_76277 (I1300302,I1300141,I1300285);
nand I_76278 (I1300319,I1300268,I1300302);
DFFARX1 I_76279 (I1300319,I3563,I1299923,I1299912,);
nor I_76280 (I1300350,I1300285,I1300042);
DFFARX1 I_76281 (I1300350,I3563,I1299923,I1299891,);
nor I_76282 (I1300381,I842691,I842682);
DFFARX1 I_76283 (I1300381,I3563,I1299923,I1300407,);
DFFARX1 I_76284 (I1300407,I3563,I1299923,I1299906,);
not I_76285 (I1300429,I1300407);
nand I_76286 (I1299903,I1300429,I1299957);
nand I_76287 (I1299897,I1300429,I1300059);
not I_76288 (I1300501,I3570);
DFFARX1 I_76289 (I914351,I3563,I1300501,I1300527,);
nand I_76290 (I1300535,I1300527,I914351);
not I_76291 (I1300552,I1300535);
DFFARX1 I_76292 (I914357,I3563,I1300501,I1300578,);
not I_76293 (I1300586,I1300578);
not I_76294 (I1300603,I914369);
or I_76295 (I1300620,I914354,I914369);
nor I_76296 (I1300637,I914354,I914369);
or I_76297 (I1300654,I914348,I914354);
DFFARX1 I_76298 (I1300654,I3563,I1300501,I1300493,);
not I_76299 (I1300685,I914366);
nand I_76300 (I1300702,I1300685,I914360);
nand I_76301 (I1300719,I1300603,I1300702);
and I_76302 (I1300472,I1300586,I1300719);
nor I_76303 (I1300750,I914366,I914348);
and I_76304 (I1300767,I1300586,I1300750);
nor I_76305 (I1300478,I1300552,I1300767);
DFFARX1 I_76306 (I1300750,I3563,I1300501,I1300807,);
not I_76307 (I1300815,I1300807);
nor I_76308 (I1300487,I1300586,I1300815);
or I_76309 (I1300846,I1300654,I914363);
nor I_76310 (I1300863,I914363,I914348);
nand I_76311 (I1300880,I1300719,I1300863);
nand I_76312 (I1300897,I1300846,I1300880);
DFFARX1 I_76313 (I1300897,I3563,I1300501,I1300490,);
nor I_76314 (I1300928,I1300863,I1300620);
DFFARX1 I_76315 (I1300928,I3563,I1300501,I1300469,);
nor I_76316 (I1300959,I914363,I914354);
DFFARX1 I_76317 (I1300959,I3563,I1300501,I1300985,);
DFFARX1 I_76318 (I1300985,I3563,I1300501,I1300484,);
not I_76319 (I1301007,I1300985);
nand I_76320 (I1300481,I1301007,I1300535);
nand I_76321 (I1300475,I1301007,I1300637);
not I_76322 (I1301079,I3570);
DFFARX1 I_76323 (I1079767,I3563,I1301079,I1301105,);
nand I_76324 (I1301113,I1301105,I1079764);
not I_76325 (I1301130,I1301113);
DFFARX1 I_76326 (I1079764,I3563,I1301079,I1301156,);
not I_76327 (I1301164,I1301156);
not I_76328 (I1301181,I1079761);
or I_76329 (I1301198,I1079770,I1079761);
nor I_76330 (I1301215,I1079770,I1079761);
or I_76331 (I1301232,I1079773,I1079770);
DFFARX1 I_76332 (I1301232,I3563,I1301079,I1301071,);
not I_76333 (I1301263,I1079761);
nand I_76334 (I1301280,I1301263,I1079758);
nand I_76335 (I1301297,I1301181,I1301280);
and I_76336 (I1301050,I1301164,I1301297);
nor I_76337 (I1301328,I1079761,I1079776);
and I_76338 (I1301345,I1301164,I1301328);
nor I_76339 (I1301056,I1301130,I1301345);
DFFARX1 I_76340 (I1301328,I3563,I1301079,I1301385,);
not I_76341 (I1301393,I1301385);
nor I_76342 (I1301065,I1301164,I1301393);
or I_76343 (I1301424,I1301232,I1079779);
nor I_76344 (I1301441,I1079779,I1079773);
nand I_76345 (I1301458,I1301297,I1301441);
nand I_76346 (I1301475,I1301424,I1301458);
DFFARX1 I_76347 (I1301475,I3563,I1301079,I1301068,);
nor I_76348 (I1301506,I1301441,I1301198);
DFFARX1 I_76349 (I1301506,I3563,I1301079,I1301047,);
nor I_76350 (I1301537,I1079779,I1079758);
DFFARX1 I_76351 (I1301537,I3563,I1301079,I1301563,);
DFFARX1 I_76352 (I1301563,I3563,I1301079,I1301062,);
not I_76353 (I1301585,I1301563);
nand I_76354 (I1301059,I1301585,I1301113);
nand I_76355 (I1301053,I1301585,I1301215);
not I_76356 (I1301657,I3570);
DFFARX1 I_76357 (I95657,I3563,I1301657,I1301683,);
nand I_76358 (I1301691,I1301683,I95648);
not I_76359 (I1301708,I1301691);
DFFARX1 I_76360 (I95645,I3563,I1301657,I1301734,);
not I_76361 (I1301742,I1301734);
not I_76362 (I1301759,I95654);
or I_76363 (I1301776,I95645,I95654);
nor I_76364 (I1301793,I95645,I95654);
or I_76365 (I1301810,I95651,I95645);
DFFARX1 I_76366 (I1301810,I3563,I1301657,I1301649,);
not I_76367 (I1301841,I95660);
nand I_76368 (I1301858,I1301841,I95669);
nand I_76369 (I1301875,I1301759,I1301858);
and I_76370 (I1301628,I1301742,I1301875);
nor I_76371 (I1301906,I95660,I95663);
and I_76372 (I1301923,I1301742,I1301906);
nor I_76373 (I1301634,I1301708,I1301923);
DFFARX1 I_76374 (I1301906,I3563,I1301657,I1301963,);
not I_76375 (I1301971,I1301963);
nor I_76376 (I1301643,I1301742,I1301971);
or I_76377 (I1302002,I1301810,I95648);
nor I_76378 (I1302019,I95648,I95651);
nand I_76379 (I1302036,I1301875,I1302019);
nand I_76380 (I1302053,I1302002,I1302036);
DFFARX1 I_76381 (I1302053,I3563,I1301657,I1301646,);
nor I_76382 (I1302084,I1302019,I1301776);
DFFARX1 I_76383 (I1302084,I3563,I1301657,I1301625,);
nor I_76384 (I1302115,I95648,I95666);
DFFARX1 I_76385 (I1302115,I3563,I1301657,I1302141,);
DFFARX1 I_76386 (I1302141,I3563,I1301657,I1301640,);
not I_76387 (I1302163,I1302141);
nand I_76388 (I1301637,I1302163,I1301691);
nand I_76389 (I1301631,I1302163,I1301793);
not I_76390 (I1302235,I3570);
DFFARX1 I_76391 (I738755,I3563,I1302235,I1302261,);
nand I_76392 (I1302269,I1302261,I738758);
not I_76393 (I1302286,I1302269);
DFFARX1 I_76394 (I738770,I3563,I1302235,I1302312,);
not I_76395 (I1302320,I1302312);
not I_76396 (I1302337,I738755);
or I_76397 (I1302354,I738764,I738755);
nor I_76398 (I1302371,I738764,I738755);
or I_76399 (I1302388,I738773,I738764);
DFFARX1 I_76400 (I1302388,I3563,I1302235,I1302227,);
not I_76401 (I1302419,I738776);
nand I_76402 (I1302436,I1302419,I738758);
nand I_76403 (I1302453,I1302337,I1302436);
and I_76404 (I1302206,I1302320,I1302453);
nor I_76405 (I1302484,I738776,I738761);
and I_76406 (I1302501,I1302320,I1302484);
nor I_76407 (I1302212,I1302286,I1302501);
DFFARX1 I_76408 (I1302484,I3563,I1302235,I1302541,);
not I_76409 (I1302549,I1302541);
nor I_76410 (I1302221,I1302320,I1302549);
or I_76411 (I1302580,I1302388,I738767);
nor I_76412 (I1302597,I738767,I738773);
nand I_76413 (I1302614,I1302453,I1302597);
nand I_76414 (I1302631,I1302580,I1302614);
DFFARX1 I_76415 (I1302631,I3563,I1302235,I1302224,);
nor I_76416 (I1302662,I1302597,I1302354);
DFFARX1 I_76417 (I1302662,I3563,I1302235,I1302203,);
nor I_76418 (I1302693,I738767,I738779);
DFFARX1 I_76419 (I1302693,I3563,I1302235,I1302719,);
DFFARX1 I_76420 (I1302719,I3563,I1302235,I1302218,);
not I_76421 (I1302741,I1302719);
nand I_76422 (I1302215,I1302741,I1302269);
nand I_76423 (I1302209,I1302741,I1302371);
not I_76424 (I1302813,I3570);
DFFARX1 I_76425 (I1069108,I3563,I1302813,I1302839,);
nand I_76426 (I1302847,I1302839,I1069105);
not I_76427 (I1302864,I1302847);
DFFARX1 I_76428 (I1069105,I3563,I1302813,I1302890,);
not I_76429 (I1302898,I1302890);
not I_76430 (I1302915,I1069102);
or I_76431 (I1302932,I1069111,I1069102);
nor I_76432 (I1302949,I1069111,I1069102);
or I_76433 (I1302966,I1069114,I1069111);
DFFARX1 I_76434 (I1302966,I3563,I1302813,I1302805,);
not I_76435 (I1302997,I1069102);
nand I_76436 (I1303014,I1302997,I1069099);
nand I_76437 (I1303031,I1302915,I1303014);
and I_76438 (I1302784,I1302898,I1303031);
nor I_76439 (I1303062,I1069102,I1069117);
and I_76440 (I1303079,I1302898,I1303062);
nor I_76441 (I1302790,I1302864,I1303079);
DFFARX1 I_76442 (I1303062,I3563,I1302813,I1303119,);
not I_76443 (I1303127,I1303119);
nor I_76444 (I1302799,I1302898,I1303127);
or I_76445 (I1303158,I1302966,I1069120);
nor I_76446 (I1303175,I1069120,I1069114);
nand I_76447 (I1303192,I1303031,I1303175);
nand I_76448 (I1303209,I1303158,I1303192);
DFFARX1 I_76449 (I1303209,I3563,I1302813,I1302802,);
nor I_76450 (I1303240,I1303175,I1302932);
DFFARX1 I_76451 (I1303240,I3563,I1302813,I1302781,);
nor I_76452 (I1303271,I1069120,I1069099);
DFFARX1 I_76453 (I1303271,I3563,I1302813,I1303297,);
DFFARX1 I_76454 (I1303297,I3563,I1302813,I1302796,);
not I_76455 (I1303319,I1303297);
nand I_76456 (I1302793,I1303319,I1302847);
nand I_76457 (I1302787,I1303319,I1302949);
not I_76458 (I1303391,I3570);
DFFARX1 I_76459 (I553081,I3563,I1303391,I1303417,);
nand I_76460 (I1303425,I1303417,I553090);
not I_76461 (I1303442,I1303425);
DFFARX1 I_76462 (I553102,I3563,I1303391,I1303468,);
not I_76463 (I1303476,I1303468);
not I_76464 (I1303493,I553093);
or I_76465 (I1303510,I553087,I553093);
nor I_76466 (I1303527,I553087,I553093);
or I_76467 (I1303544,I553081,I553087);
DFFARX1 I_76468 (I1303544,I3563,I1303391,I1303383,);
not I_76469 (I1303575,I553084);
nand I_76470 (I1303592,I1303575,I553096);
nand I_76471 (I1303609,I1303493,I1303592);
and I_76472 (I1303362,I1303476,I1303609);
nor I_76473 (I1303640,I553084,I553105);
and I_76474 (I1303657,I1303476,I1303640);
nor I_76475 (I1303368,I1303442,I1303657);
DFFARX1 I_76476 (I1303640,I3563,I1303391,I1303697,);
not I_76477 (I1303705,I1303697);
nor I_76478 (I1303377,I1303476,I1303705);
or I_76479 (I1303736,I1303544,I553099);
nor I_76480 (I1303753,I553099,I553081);
nand I_76481 (I1303770,I1303609,I1303753);
nand I_76482 (I1303787,I1303736,I1303770);
DFFARX1 I_76483 (I1303787,I3563,I1303391,I1303380,);
nor I_76484 (I1303818,I1303753,I1303510);
DFFARX1 I_76485 (I1303818,I3563,I1303391,I1303359,);
nor I_76486 (I1303849,I553099,I553084);
DFFARX1 I_76487 (I1303849,I3563,I1303391,I1303875,);
DFFARX1 I_76488 (I1303875,I3563,I1303391,I1303374,);
not I_76489 (I1303897,I1303875);
nand I_76490 (I1303371,I1303897,I1303425);
nand I_76491 (I1303365,I1303897,I1303527);
not I_76492 (I1303969,I3570);
DFFARX1 I_76493 (I79320,I3563,I1303969,I1303995,);
nand I_76494 (I1304003,I1303995,I79311);
not I_76495 (I1304020,I1304003);
DFFARX1 I_76496 (I79308,I3563,I1303969,I1304046,);
not I_76497 (I1304054,I1304046);
not I_76498 (I1304071,I79317);
or I_76499 (I1304088,I79308,I79317);
nor I_76500 (I1304105,I79308,I79317);
or I_76501 (I1304122,I79314,I79308);
DFFARX1 I_76502 (I1304122,I3563,I1303969,I1303961,);
not I_76503 (I1304153,I79323);
nand I_76504 (I1304170,I1304153,I79332);
nand I_76505 (I1304187,I1304071,I1304170);
and I_76506 (I1303940,I1304054,I1304187);
nor I_76507 (I1304218,I79323,I79326);
and I_76508 (I1304235,I1304054,I1304218);
nor I_76509 (I1303946,I1304020,I1304235);
DFFARX1 I_76510 (I1304218,I3563,I1303969,I1304275,);
not I_76511 (I1304283,I1304275);
nor I_76512 (I1303955,I1304054,I1304283);
or I_76513 (I1304314,I1304122,I79311);
nor I_76514 (I1304331,I79311,I79314);
nand I_76515 (I1304348,I1304187,I1304331);
nand I_76516 (I1304365,I1304314,I1304348);
DFFARX1 I_76517 (I1304365,I3563,I1303969,I1303958,);
nor I_76518 (I1304396,I1304331,I1304088);
DFFARX1 I_76519 (I1304396,I3563,I1303969,I1303937,);
nor I_76520 (I1304427,I79311,I79329);
DFFARX1 I_76521 (I1304427,I3563,I1303969,I1304453,);
DFFARX1 I_76522 (I1304453,I3563,I1303969,I1303952,);
not I_76523 (I1304475,I1304453);
nand I_76524 (I1303949,I1304475,I1304003);
nand I_76525 (I1303943,I1304475,I1304105);
not I_76526 (I1304547,I3570);
DFFARX1 I_76527 (I340706,I3563,I1304547,I1304573,);
nand I_76528 (I1304581,I1304573,I340727);
not I_76529 (I1304598,I1304581);
DFFARX1 I_76530 (I340721,I3563,I1304547,I1304624,);
not I_76531 (I1304632,I1304624);
not I_76532 (I1304649,I340709);
or I_76533 (I1304666,I340724,I340709);
nor I_76534 (I1304683,I340724,I340709);
or I_76535 (I1304700,I340715,I340724);
DFFARX1 I_76536 (I1304700,I3563,I1304547,I1304539,);
not I_76537 (I1304731,I340703);
nand I_76538 (I1304748,I1304731,I340700);
nand I_76539 (I1304765,I1304649,I1304748);
and I_76540 (I1304518,I1304632,I1304765);
nor I_76541 (I1304796,I340703,I340712);
and I_76542 (I1304813,I1304632,I1304796);
nor I_76543 (I1304524,I1304598,I1304813);
DFFARX1 I_76544 (I1304796,I3563,I1304547,I1304853,);
not I_76545 (I1304861,I1304853);
nor I_76546 (I1304533,I1304632,I1304861);
or I_76547 (I1304892,I1304700,I340718);
nor I_76548 (I1304909,I340718,I340715);
nand I_76549 (I1304926,I1304765,I1304909);
nand I_76550 (I1304943,I1304892,I1304926);
DFFARX1 I_76551 (I1304943,I3563,I1304547,I1304536,);
nor I_76552 (I1304974,I1304909,I1304666);
DFFARX1 I_76553 (I1304974,I3563,I1304547,I1304515,);
nor I_76554 (I1305005,I340718,I340700);
DFFARX1 I_76555 (I1305005,I3563,I1304547,I1305031,);
DFFARX1 I_76556 (I1305031,I3563,I1304547,I1304530,);
not I_76557 (I1305053,I1305031);
nand I_76558 (I1304527,I1305053,I1304581);
nand I_76559 (I1304521,I1305053,I1304683);
not I_76560 (I1305125,I3570);
DFFARX1 I_76561 (I849530,I3563,I1305125,I1305151,);
nand I_76562 (I1305159,I1305151,I849530);
not I_76563 (I1305176,I1305159);
DFFARX1 I_76564 (I849536,I3563,I1305125,I1305202,);
not I_76565 (I1305210,I1305202);
not I_76566 (I1305227,I849548);
or I_76567 (I1305244,I849533,I849548);
nor I_76568 (I1305261,I849533,I849548);
or I_76569 (I1305278,I849527,I849533);
DFFARX1 I_76570 (I1305278,I3563,I1305125,I1305117,);
not I_76571 (I1305309,I849545);
nand I_76572 (I1305326,I1305309,I849539);
nand I_76573 (I1305343,I1305227,I1305326);
and I_76574 (I1305096,I1305210,I1305343);
nor I_76575 (I1305374,I849545,I849527);
and I_76576 (I1305391,I1305210,I1305374);
nor I_76577 (I1305102,I1305176,I1305391);
DFFARX1 I_76578 (I1305374,I3563,I1305125,I1305431,);
not I_76579 (I1305439,I1305431);
nor I_76580 (I1305111,I1305210,I1305439);
or I_76581 (I1305470,I1305278,I849542);
nor I_76582 (I1305487,I849542,I849527);
nand I_76583 (I1305504,I1305343,I1305487);
nand I_76584 (I1305521,I1305470,I1305504);
DFFARX1 I_76585 (I1305521,I3563,I1305125,I1305114,);
nor I_76586 (I1305552,I1305487,I1305244);
DFFARX1 I_76587 (I1305552,I3563,I1305125,I1305093,);
nor I_76588 (I1305583,I849542,I849533);
DFFARX1 I_76589 (I1305583,I3563,I1305125,I1305609,);
DFFARX1 I_76590 (I1305609,I3563,I1305125,I1305108,);
not I_76591 (I1305631,I1305609);
nand I_76592 (I1305105,I1305631,I1305159);
nand I_76593 (I1305099,I1305631,I1305261);
not I_76594 (I1305703,I3570);
DFFARX1 I_76595 (I1077523,I3563,I1305703,I1305729,);
nand I_76596 (I1305737,I1305729,I1077520);
not I_76597 (I1305754,I1305737);
DFFARX1 I_76598 (I1077520,I3563,I1305703,I1305780,);
not I_76599 (I1305788,I1305780);
not I_76600 (I1305805,I1077517);
or I_76601 (I1305822,I1077526,I1077517);
nor I_76602 (I1305839,I1077526,I1077517);
or I_76603 (I1305856,I1077529,I1077526);
DFFARX1 I_76604 (I1305856,I3563,I1305703,I1305695,);
not I_76605 (I1305887,I1077517);
nand I_76606 (I1305904,I1305887,I1077514);
nand I_76607 (I1305921,I1305805,I1305904);
and I_76608 (I1305674,I1305788,I1305921);
nor I_76609 (I1305952,I1077517,I1077532);
and I_76610 (I1305969,I1305788,I1305952);
nor I_76611 (I1305680,I1305754,I1305969);
DFFARX1 I_76612 (I1305952,I3563,I1305703,I1306009,);
not I_76613 (I1306017,I1306009);
nor I_76614 (I1305689,I1305788,I1306017);
or I_76615 (I1306048,I1305856,I1077535);
nor I_76616 (I1306065,I1077535,I1077529);
nand I_76617 (I1306082,I1305921,I1306065);
nand I_76618 (I1306099,I1306048,I1306082);
DFFARX1 I_76619 (I1306099,I3563,I1305703,I1305692,);
nor I_76620 (I1306130,I1306065,I1305822);
DFFARX1 I_76621 (I1306130,I3563,I1305703,I1305671,);
nor I_76622 (I1306161,I1077535,I1077514);
DFFARX1 I_76623 (I1306161,I3563,I1305703,I1306187,);
DFFARX1 I_76624 (I1306187,I3563,I1305703,I1305686,);
not I_76625 (I1306209,I1306187);
nand I_76626 (I1305683,I1306209,I1305737);
nand I_76627 (I1305677,I1306209,I1305839);
not I_76628 (I1306281,I3570);
DFFARX1 I_76629 (I909608,I3563,I1306281,I1306307,);
nand I_76630 (I1306315,I1306307,I909608);
not I_76631 (I1306332,I1306315);
DFFARX1 I_76632 (I909614,I3563,I1306281,I1306358,);
not I_76633 (I1306366,I1306358);
not I_76634 (I1306383,I909626);
or I_76635 (I1306400,I909611,I909626);
nor I_76636 (I1306417,I909611,I909626);
or I_76637 (I1306434,I909605,I909611);
DFFARX1 I_76638 (I1306434,I3563,I1306281,I1306273,);
not I_76639 (I1306465,I909623);
nand I_76640 (I1306482,I1306465,I909617);
nand I_76641 (I1306499,I1306383,I1306482);
and I_76642 (I1306252,I1306366,I1306499);
nor I_76643 (I1306530,I909623,I909605);
and I_76644 (I1306547,I1306366,I1306530);
nor I_76645 (I1306258,I1306332,I1306547);
DFFARX1 I_76646 (I1306530,I3563,I1306281,I1306587,);
not I_76647 (I1306595,I1306587);
nor I_76648 (I1306267,I1306366,I1306595);
or I_76649 (I1306626,I1306434,I909620);
nor I_76650 (I1306643,I909620,I909605);
nand I_76651 (I1306660,I1306499,I1306643);
nand I_76652 (I1306677,I1306626,I1306660);
DFFARX1 I_76653 (I1306677,I3563,I1306281,I1306270,);
nor I_76654 (I1306708,I1306643,I1306400);
DFFARX1 I_76655 (I1306708,I3563,I1306281,I1306249,);
nor I_76656 (I1306739,I909620,I909611);
DFFARX1 I_76657 (I1306739,I3563,I1306281,I1306765,);
DFFARX1 I_76658 (I1306765,I3563,I1306281,I1306264,);
not I_76659 (I1306787,I1306765);
nand I_76660 (I1306261,I1306787,I1306315);
nand I_76661 (I1306255,I1306787,I1306417);
not I_76662 (I1306859,I3570);
DFFARX1 I_76663 (I1026639,I3563,I1306859,I1306885,);
nand I_76664 (I1306893,I1306885,I1026660);
not I_76665 (I1306910,I1306893);
DFFARX1 I_76666 (I1026633,I3563,I1306859,I1306936,);
not I_76667 (I1306944,I1306936);
not I_76668 (I1306961,I1026654);
or I_76669 (I1306978,I1026645,I1026654);
nor I_76670 (I1306995,I1026645,I1026654);
or I_76671 (I1307012,I1026648,I1026645);
DFFARX1 I_76672 (I1307012,I3563,I1306859,I1306851,);
not I_76673 (I1307043,I1026636);
nand I_76674 (I1307060,I1307043,I1026651);
nand I_76675 (I1307077,I1306961,I1307060);
and I_76676 (I1306830,I1306944,I1307077);
nor I_76677 (I1307108,I1026636,I1026633);
and I_76678 (I1307125,I1306944,I1307108);
nor I_76679 (I1306836,I1306910,I1307125);
DFFARX1 I_76680 (I1307108,I3563,I1306859,I1307165,);
not I_76681 (I1307173,I1307165);
nor I_76682 (I1306845,I1306944,I1307173);
or I_76683 (I1307204,I1307012,I1026657);
nor I_76684 (I1307221,I1026657,I1026648);
nand I_76685 (I1307238,I1307077,I1307221);
nand I_76686 (I1307255,I1307204,I1307238);
DFFARX1 I_76687 (I1307255,I3563,I1306859,I1306848,);
nor I_76688 (I1307286,I1307221,I1306978);
DFFARX1 I_76689 (I1307286,I3563,I1306859,I1306827,);
nor I_76690 (I1307317,I1026657,I1026642);
DFFARX1 I_76691 (I1307317,I3563,I1306859,I1307343,);
DFFARX1 I_76692 (I1307343,I3563,I1306859,I1306842,);
not I_76693 (I1307365,I1307343);
nand I_76694 (I1306839,I1307365,I1306893);
nand I_76695 (I1306833,I1307365,I1306995);
not I_76696 (I1307437,I3570);
DFFARX1 I_76697 (I875353,I3563,I1307437,I1307463,);
nand I_76698 (I1307471,I1307463,I875353);
not I_76699 (I1307488,I1307471);
DFFARX1 I_76700 (I875359,I3563,I1307437,I1307514,);
not I_76701 (I1307522,I1307514);
not I_76702 (I1307539,I875371);
or I_76703 (I1307556,I875356,I875371);
nor I_76704 (I1307573,I875356,I875371);
or I_76705 (I1307590,I875350,I875356);
DFFARX1 I_76706 (I1307590,I3563,I1307437,I1307429,);
not I_76707 (I1307621,I875368);
nand I_76708 (I1307638,I1307621,I875362);
nand I_76709 (I1307655,I1307539,I1307638);
and I_76710 (I1307408,I1307522,I1307655);
nor I_76711 (I1307686,I875368,I875350);
and I_76712 (I1307703,I1307522,I1307686);
nor I_76713 (I1307414,I1307488,I1307703);
DFFARX1 I_76714 (I1307686,I3563,I1307437,I1307743,);
not I_76715 (I1307751,I1307743);
nor I_76716 (I1307423,I1307522,I1307751);
or I_76717 (I1307782,I1307590,I875365);
nor I_76718 (I1307799,I875365,I875350);
nand I_76719 (I1307816,I1307655,I1307799);
nand I_76720 (I1307833,I1307782,I1307816);
DFFARX1 I_76721 (I1307833,I3563,I1307437,I1307426,);
nor I_76722 (I1307864,I1307799,I1307556);
DFFARX1 I_76723 (I1307864,I3563,I1307437,I1307405,);
nor I_76724 (I1307895,I875365,I875356);
DFFARX1 I_76725 (I1307895,I3563,I1307437,I1307921,);
DFFARX1 I_76726 (I1307921,I3563,I1307437,I1307420,);
not I_76727 (I1307943,I1307921);
nand I_76728 (I1307417,I1307943,I1307471);
nand I_76729 (I1307411,I1307943,I1307573);
not I_76730 (I1308015,I3570);
DFFARX1 I_76731 (I1110665,I3563,I1308015,I1308041,);
nand I_76732 (I1308049,I1308041,I1110650);
not I_76733 (I1308066,I1308049);
DFFARX1 I_76734 (I1110653,I3563,I1308015,I1308092,);
not I_76735 (I1308100,I1308092);
not I_76736 (I1308117,I1110668);
or I_76737 (I1308134,I1110671,I1110668);
nor I_76738 (I1308151,I1110671,I1110668);
or I_76739 (I1308168,I1110647,I1110671);
DFFARX1 I_76740 (I1308168,I3563,I1308015,I1308007,);
not I_76741 (I1308199,I1110659);
nand I_76742 (I1308216,I1308199,I1110662);
nand I_76743 (I1308233,I1308117,I1308216);
and I_76744 (I1307986,I1308100,I1308233);
nor I_76745 (I1308264,I1110659,I1110656);
and I_76746 (I1308281,I1308100,I1308264);
nor I_76747 (I1307992,I1308066,I1308281);
DFFARX1 I_76748 (I1308264,I3563,I1308015,I1308321,);
not I_76749 (I1308329,I1308321);
nor I_76750 (I1308001,I1308100,I1308329);
or I_76751 (I1308360,I1308168,I1110647);
nor I_76752 (I1308377,I1110647,I1110647);
nand I_76753 (I1308394,I1308233,I1308377);
nand I_76754 (I1308411,I1308360,I1308394);
DFFARX1 I_76755 (I1308411,I3563,I1308015,I1308004,);
nor I_76756 (I1308442,I1308377,I1308134);
DFFARX1 I_76757 (I1308442,I3563,I1308015,I1307983,);
nor I_76758 (I1308473,I1110647,I1110650);
DFFARX1 I_76759 (I1308473,I3563,I1308015,I1308499,);
DFFARX1 I_76760 (I1308499,I3563,I1308015,I1307998,);
not I_76761 (I1308521,I1308499);
nand I_76762 (I1307995,I1308521,I1308049);
nand I_76763 (I1307989,I1308521,I1308151);
not I_76764 (I1308593,I3570);
DFFARX1 I_76765 (I1215861,I3563,I1308593,I1308619,);
nand I_76766 (I1308627,I1308619,I1215846);
not I_76767 (I1308644,I1308627);
DFFARX1 I_76768 (I1215849,I3563,I1308593,I1308670,);
not I_76769 (I1308678,I1308670);
not I_76770 (I1308695,I1215864);
or I_76771 (I1308712,I1215867,I1215864);
nor I_76772 (I1308729,I1215867,I1215864);
or I_76773 (I1308746,I1215843,I1215867);
DFFARX1 I_76774 (I1308746,I3563,I1308593,I1308585,);
not I_76775 (I1308777,I1215855);
nand I_76776 (I1308794,I1308777,I1215858);
nand I_76777 (I1308811,I1308695,I1308794);
and I_76778 (I1308564,I1308678,I1308811);
nor I_76779 (I1308842,I1215855,I1215852);
and I_76780 (I1308859,I1308678,I1308842);
nor I_76781 (I1308570,I1308644,I1308859);
DFFARX1 I_76782 (I1308842,I3563,I1308593,I1308899,);
not I_76783 (I1308907,I1308899);
nor I_76784 (I1308579,I1308678,I1308907);
or I_76785 (I1308938,I1308746,I1215843);
nor I_76786 (I1308955,I1215843,I1215843);
nand I_76787 (I1308972,I1308811,I1308955);
nand I_76788 (I1308989,I1308938,I1308972);
DFFARX1 I_76789 (I1308989,I3563,I1308593,I1308582,);
nor I_76790 (I1309020,I1308955,I1308712);
DFFARX1 I_76791 (I1309020,I3563,I1308593,I1308561,);
nor I_76792 (I1309051,I1215843,I1215846);
DFFARX1 I_76793 (I1309051,I3563,I1308593,I1309077,);
DFFARX1 I_76794 (I1309077,I3563,I1308593,I1308576,);
not I_76795 (I1309099,I1309077);
nand I_76796 (I1308573,I1309099,I1308627);
nand I_76797 (I1308567,I1309099,I1308729);
not I_76798 (I1309171,I3570);
DFFARX1 I_76799 (I1386887,I3563,I1309171,I1309197,);
nand I_76800 (I1309205,I1309197,I1386878);
not I_76801 (I1309222,I1309205);
DFFARX1 I_76802 (I1386863,I3563,I1309171,I1309248,);
not I_76803 (I1309256,I1309248);
not I_76804 (I1309273,I1386866);
or I_76805 (I1309290,I1386875,I1386866);
nor I_76806 (I1309307,I1386875,I1386866);
or I_76807 (I1309324,I1386872,I1386875);
DFFARX1 I_76808 (I1309324,I3563,I1309171,I1309163,);
not I_76809 (I1309355,I1386884);
nand I_76810 (I1309372,I1309355,I1386863);
nand I_76811 (I1309389,I1309273,I1309372);
and I_76812 (I1309142,I1309256,I1309389);
nor I_76813 (I1309420,I1386884,I1386869);
and I_76814 (I1309437,I1309256,I1309420);
nor I_76815 (I1309148,I1309222,I1309437);
DFFARX1 I_76816 (I1309420,I3563,I1309171,I1309477,);
not I_76817 (I1309485,I1309477);
nor I_76818 (I1309157,I1309256,I1309485);
or I_76819 (I1309516,I1309324,I1386890);
nor I_76820 (I1309533,I1386890,I1386872);
nand I_76821 (I1309550,I1309389,I1309533);
nand I_76822 (I1309567,I1309516,I1309550);
DFFARX1 I_76823 (I1309567,I3563,I1309171,I1309160,);
nor I_76824 (I1309598,I1309533,I1309290);
DFFARX1 I_76825 (I1309598,I3563,I1309171,I1309139,);
nor I_76826 (I1309629,I1386890,I1386881);
DFFARX1 I_76827 (I1309629,I3563,I1309171,I1309655,);
DFFARX1 I_76828 (I1309655,I3563,I1309171,I1309154,);
not I_76829 (I1309677,I1309655);
nand I_76830 (I1309151,I1309677,I1309205);
nand I_76831 (I1309145,I1309677,I1309307);
not I_76832 (I1309749,I3570);
DFFARX1 I_76833 (I742801,I3563,I1309749,I1309775,);
nand I_76834 (I1309783,I1309775,I742804);
not I_76835 (I1309800,I1309783);
DFFARX1 I_76836 (I742816,I3563,I1309749,I1309826,);
not I_76837 (I1309834,I1309826);
not I_76838 (I1309851,I742801);
or I_76839 (I1309868,I742810,I742801);
nor I_76840 (I1309885,I742810,I742801);
or I_76841 (I1309902,I742819,I742810);
DFFARX1 I_76842 (I1309902,I3563,I1309749,I1309741,);
not I_76843 (I1309933,I742822);
nand I_76844 (I1309950,I1309933,I742804);
nand I_76845 (I1309967,I1309851,I1309950);
and I_76846 (I1309720,I1309834,I1309967);
nor I_76847 (I1309998,I742822,I742807);
and I_76848 (I1310015,I1309834,I1309998);
nor I_76849 (I1309726,I1309800,I1310015);
DFFARX1 I_76850 (I1309998,I3563,I1309749,I1310055,);
not I_76851 (I1310063,I1310055);
nor I_76852 (I1309735,I1309834,I1310063);
or I_76853 (I1310094,I1309902,I742813);
nor I_76854 (I1310111,I742813,I742819);
nand I_76855 (I1310128,I1309967,I1310111);
nand I_76856 (I1310145,I1310094,I1310128);
DFFARX1 I_76857 (I1310145,I3563,I1309749,I1309738,);
nor I_76858 (I1310176,I1310111,I1309868);
DFFARX1 I_76859 (I1310176,I3563,I1309749,I1309717,);
nor I_76860 (I1310207,I742813,I742825);
DFFARX1 I_76861 (I1310207,I3563,I1309749,I1310233,);
DFFARX1 I_76862 (I1310233,I3563,I1309749,I1309732,);
not I_76863 (I1310255,I1310233);
nand I_76864 (I1309729,I1310255,I1309783);
nand I_76865 (I1309723,I1310255,I1309885);
not I_76866 (I1310327,I3570);
DFFARX1 I_76867 (I310667,I3563,I1310327,I1310353,);
nand I_76868 (I1310361,I1310353,I310688);
not I_76869 (I1310378,I1310361);
DFFARX1 I_76870 (I310682,I3563,I1310327,I1310404,);
not I_76871 (I1310412,I1310404);
not I_76872 (I1310429,I310670);
or I_76873 (I1310446,I310685,I310670);
nor I_76874 (I1310463,I310685,I310670);
or I_76875 (I1310480,I310676,I310685);
DFFARX1 I_76876 (I1310480,I3563,I1310327,I1310319,);
not I_76877 (I1310511,I310664);
nand I_76878 (I1310528,I1310511,I310661);
nand I_76879 (I1310545,I1310429,I1310528);
and I_76880 (I1310298,I1310412,I1310545);
nor I_76881 (I1310576,I310664,I310673);
and I_76882 (I1310593,I1310412,I1310576);
nor I_76883 (I1310304,I1310378,I1310593);
DFFARX1 I_76884 (I1310576,I3563,I1310327,I1310633,);
not I_76885 (I1310641,I1310633);
nor I_76886 (I1310313,I1310412,I1310641);
or I_76887 (I1310672,I1310480,I310679);
nor I_76888 (I1310689,I310679,I310676);
nand I_76889 (I1310706,I1310545,I1310689);
nand I_76890 (I1310723,I1310672,I1310706);
DFFARX1 I_76891 (I1310723,I3563,I1310327,I1310316,);
nor I_76892 (I1310754,I1310689,I1310446);
DFFARX1 I_76893 (I1310754,I3563,I1310327,I1310295,);
nor I_76894 (I1310785,I310679,I310661);
DFFARX1 I_76895 (I1310785,I3563,I1310327,I1310811,);
DFFARX1 I_76896 (I1310811,I3563,I1310327,I1310310,);
not I_76897 (I1310833,I1310811);
nand I_76898 (I1310307,I1310833,I1310361);
nand I_76899 (I1310301,I1310833,I1310463);
not I_76900 (I1310905,I3570);
DFFARX1 I_76901 (I1105463,I3563,I1310905,I1310931,);
nand I_76902 (I1310939,I1310931,I1105448);
not I_76903 (I1310956,I1310939);
DFFARX1 I_76904 (I1105451,I3563,I1310905,I1310982,);
not I_76905 (I1310990,I1310982);
not I_76906 (I1311007,I1105466);
or I_76907 (I1311024,I1105469,I1105466);
nor I_76908 (I1311041,I1105469,I1105466);
or I_76909 (I1311058,I1105445,I1105469);
DFFARX1 I_76910 (I1311058,I3563,I1310905,I1310897,);
not I_76911 (I1311089,I1105457);
nand I_76912 (I1311106,I1311089,I1105460);
nand I_76913 (I1311123,I1311007,I1311106);
and I_76914 (I1310876,I1310990,I1311123);
nor I_76915 (I1311154,I1105457,I1105454);
and I_76916 (I1311171,I1310990,I1311154);
nor I_76917 (I1310882,I1310956,I1311171);
DFFARX1 I_76918 (I1311154,I3563,I1310905,I1311211,);
not I_76919 (I1311219,I1311211);
nor I_76920 (I1310891,I1310990,I1311219);
or I_76921 (I1311250,I1311058,I1105445);
nor I_76922 (I1311267,I1105445,I1105445);
nand I_76923 (I1311284,I1311123,I1311267);
nand I_76924 (I1311301,I1311250,I1311284);
DFFARX1 I_76925 (I1311301,I3563,I1310905,I1310894,);
nor I_76926 (I1311332,I1311267,I1311024);
DFFARX1 I_76927 (I1311332,I3563,I1310905,I1310873,);
nor I_76928 (I1311363,I1105445,I1105448);
DFFARX1 I_76929 (I1311363,I3563,I1310905,I1311389,);
DFFARX1 I_76930 (I1311389,I3563,I1310905,I1310888,);
not I_76931 (I1311411,I1311389);
nand I_76932 (I1310885,I1311411,I1310939);
nand I_76933 (I1310879,I1311411,I1311041);
not I_76934 (I1311483,I3570);
DFFARX1 I_76935 (I784995,I3563,I1311483,I1311509,);
nand I_76936 (I1311517,I1311509,I784998);
not I_76937 (I1311534,I1311517);
DFFARX1 I_76938 (I785010,I3563,I1311483,I1311560,);
not I_76939 (I1311568,I1311560);
not I_76940 (I1311585,I784995);
or I_76941 (I1311602,I785004,I784995);
nor I_76942 (I1311619,I785004,I784995);
or I_76943 (I1311636,I785013,I785004);
DFFARX1 I_76944 (I1311636,I3563,I1311483,I1311475,);
not I_76945 (I1311667,I785016);
nand I_76946 (I1311684,I1311667,I784998);
nand I_76947 (I1311701,I1311585,I1311684);
and I_76948 (I1311454,I1311568,I1311701);
nor I_76949 (I1311732,I785016,I785001);
and I_76950 (I1311749,I1311568,I1311732);
nor I_76951 (I1311460,I1311534,I1311749);
DFFARX1 I_76952 (I1311732,I3563,I1311483,I1311789,);
not I_76953 (I1311797,I1311789);
nor I_76954 (I1311469,I1311568,I1311797);
or I_76955 (I1311828,I1311636,I785007);
nor I_76956 (I1311845,I785007,I785013);
nand I_76957 (I1311862,I1311701,I1311845);
nand I_76958 (I1311879,I1311828,I1311862);
DFFARX1 I_76959 (I1311879,I3563,I1311483,I1311472,);
nor I_76960 (I1311910,I1311845,I1311602);
DFFARX1 I_76961 (I1311910,I3563,I1311483,I1311451,);
nor I_76962 (I1311941,I785007,I785019);
DFFARX1 I_76963 (I1311941,I3563,I1311483,I1311967,);
DFFARX1 I_76964 (I1311967,I3563,I1311483,I1311466,);
not I_76965 (I1311989,I1311967);
nand I_76966 (I1311463,I1311989,I1311517);
nand I_76967 (I1311457,I1311989,I1311619);
not I_76968 (I1312061,I3570);
DFFARX1 I_76969 (I280333,I3563,I1312061,I1312087,);
nand I_76970 (I1312095,I1312087,I280336);
not I_76971 (I1312112,I1312095);
DFFARX1 I_76972 (I280345,I3563,I1312061,I1312138,);
not I_76973 (I1312146,I1312138);
not I_76974 (I1312163,I280348);
or I_76975 (I1312180,I280339,I280348);
nor I_76976 (I1312197,I280339,I280348);
or I_76977 (I1312214,I280351,I280339);
DFFARX1 I_76978 (I1312214,I3563,I1312061,I1312053,);
not I_76979 (I1312245,I280336);
nand I_76980 (I1312262,I1312245,I280342);
nand I_76981 (I1312279,I1312163,I1312262);
and I_76982 (I1312032,I1312146,I1312279);
nor I_76983 (I1312310,I280336,I280354);
and I_76984 (I1312327,I1312146,I1312310);
nor I_76985 (I1312038,I1312112,I1312327);
DFFARX1 I_76986 (I1312310,I3563,I1312061,I1312367,);
not I_76987 (I1312375,I1312367);
nor I_76988 (I1312047,I1312146,I1312375);
or I_76989 (I1312406,I1312214,I280333);
nor I_76990 (I1312423,I280333,I280351);
nand I_76991 (I1312440,I1312279,I1312423);
nand I_76992 (I1312457,I1312406,I1312440);
DFFARX1 I_76993 (I1312457,I3563,I1312061,I1312050,);
nor I_76994 (I1312488,I1312423,I1312180);
DFFARX1 I_76995 (I1312488,I3563,I1312061,I1312029,);
nor I_76996 (I1312519,I280333,I280357);
DFFARX1 I_76997 (I1312519,I3563,I1312061,I1312545,);
DFFARX1 I_76998 (I1312545,I3563,I1312061,I1312044,);
not I_76999 (I1312567,I1312545);
nand I_77000 (I1312041,I1312567,I1312095);
nand I_77001 (I1312035,I1312567,I1312197);
not I_77002 (I1312639,I3570);
DFFARX1 I_77003 (I702341,I3563,I1312639,I1312665,);
nand I_77004 (I1312673,I1312665,I702344);
not I_77005 (I1312690,I1312673);
DFFARX1 I_77006 (I702356,I3563,I1312639,I1312716,);
not I_77007 (I1312724,I1312716);
not I_77008 (I1312741,I702341);
or I_77009 (I1312758,I702350,I702341);
nor I_77010 (I1312775,I702350,I702341);
or I_77011 (I1312792,I702359,I702350);
DFFARX1 I_77012 (I1312792,I3563,I1312639,I1312631,);
not I_77013 (I1312823,I702362);
nand I_77014 (I1312840,I1312823,I702344);
nand I_77015 (I1312857,I1312741,I1312840);
and I_77016 (I1312610,I1312724,I1312857);
nor I_77017 (I1312888,I702362,I702347);
and I_77018 (I1312905,I1312724,I1312888);
nor I_77019 (I1312616,I1312690,I1312905);
DFFARX1 I_77020 (I1312888,I3563,I1312639,I1312945,);
not I_77021 (I1312953,I1312945);
nor I_77022 (I1312625,I1312724,I1312953);
or I_77023 (I1312984,I1312792,I702353);
nor I_77024 (I1313001,I702353,I702359);
nand I_77025 (I1313018,I1312857,I1313001);
nand I_77026 (I1313035,I1312984,I1313018);
DFFARX1 I_77027 (I1313035,I3563,I1312639,I1312628,);
nor I_77028 (I1313066,I1313001,I1312758);
DFFARX1 I_77029 (I1313066,I3563,I1312639,I1312607,);
nor I_77030 (I1313097,I702353,I702365);
DFFARX1 I_77031 (I1313097,I3563,I1312639,I1313123,);
DFFARX1 I_77032 (I1313123,I3563,I1312639,I1312622,);
not I_77033 (I1313145,I1313123);
nand I_77034 (I1312619,I1313145,I1312673);
nand I_77035 (I1312613,I1313145,I1312775);
not I_77036 (I1313217,I3570);
DFFARX1 I_77037 (I1254040,I3563,I1313217,I1313243,);
nand I_77038 (I1313251,I1313243,I1254049);
not I_77039 (I1313268,I1313251);
DFFARX1 I_77040 (I1254025,I3563,I1313217,I1313294,);
not I_77041 (I1313302,I1313294);
not I_77042 (I1313319,I1254028);
or I_77043 (I1313336,I1254025,I1254028);
nor I_77044 (I1313353,I1254025,I1254028);
or I_77045 (I1313370,I1254043,I1254025);
DFFARX1 I_77046 (I1313370,I3563,I1313217,I1313209,);
not I_77047 (I1313401,I1254031);
nand I_77048 (I1313418,I1313401,I1254046);
nand I_77049 (I1313435,I1313319,I1313418);
and I_77050 (I1313188,I1313302,I1313435);
nor I_77051 (I1313466,I1254031,I1254034);
and I_77052 (I1313483,I1313302,I1313466);
nor I_77053 (I1313194,I1313268,I1313483);
DFFARX1 I_77054 (I1313466,I3563,I1313217,I1313523,);
not I_77055 (I1313531,I1313523);
nor I_77056 (I1313203,I1313302,I1313531);
or I_77057 (I1313562,I1313370,I1254037);
nor I_77058 (I1313579,I1254037,I1254043);
nand I_77059 (I1313596,I1313435,I1313579);
nand I_77060 (I1313613,I1313562,I1313596);
DFFARX1 I_77061 (I1313613,I3563,I1313217,I1313206,);
nor I_77062 (I1313644,I1313579,I1313336);
DFFARX1 I_77063 (I1313644,I3563,I1313217,I1313185,);
nor I_77064 (I1313675,I1254037,I1254028);
DFFARX1 I_77065 (I1313675,I3563,I1313217,I1313701,);
DFFARX1 I_77066 (I1313701,I3563,I1313217,I1313200,);
not I_77067 (I1313723,I1313701);
nand I_77068 (I1313197,I1313723,I1313251);
nand I_77069 (I1313191,I1313723,I1313353);
not I_77070 (I1313795,I3570);
DFFARX1 I_77071 (I134128,I3563,I1313795,I1313821,);
nand I_77072 (I1313829,I1313821,I134119);
not I_77073 (I1313846,I1313829);
DFFARX1 I_77074 (I134116,I3563,I1313795,I1313872,);
not I_77075 (I1313880,I1313872);
not I_77076 (I1313897,I134125);
or I_77077 (I1313914,I134116,I134125);
nor I_77078 (I1313931,I134116,I134125);
or I_77079 (I1313948,I134122,I134116);
DFFARX1 I_77080 (I1313948,I3563,I1313795,I1313787,);
not I_77081 (I1313979,I134131);
nand I_77082 (I1313996,I1313979,I134140);
nand I_77083 (I1314013,I1313897,I1313996);
and I_77084 (I1313766,I1313880,I1314013);
nor I_77085 (I1314044,I134131,I134134);
and I_77086 (I1314061,I1313880,I1314044);
nor I_77087 (I1313772,I1313846,I1314061);
DFFARX1 I_77088 (I1314044,I3563,I1313795,I1314101,);
not I_77089 (I1314109,I1314101);
nor I_77090 (I1313781,I1313880,I1314109);
or I_77091 (I1314140,I1313948,I134119);
nor I_77092 (I1314157,I134119,I134122);
nand I_77093 (I1314174,I1314013,I1314157);
nand I_77094 (I1314191,I1314140,I1314174);
DFFARX1 I_77095 (I1314191,I3563,I1313795,I1313784,);
nor I_77096 (I1314222,I1314157,I1313914);
DFFARX1 I_77097 (I1314222,I3563,I1313795,I1313763,);
nor I_77098 (I1314253,I134119,I134137);
DFFARX1 I_77099 (I1314253,I3563,I1313795,I1314279,);
DFFARX1 I_77100 (I1314279,I3563,I1313795,I1313778,);
not I_77101 (I1314301,I1314279);
nand I_77102 (I1313775,I1314301,I1313829);
nand I_77103 (I1313769,I1314301,I1313931);
not I_77104 (I1314373,I3570);
DFFARX1 I_77105 (I1354162,I3563,I1314373,I1314399,);
nand I_77106 (I1314407,I1314399,I1354153);
not I_77107 (I1314424,I1314407);
DFFARX1 I_77108 (I1354138,I3563,I1314373,I1314450,);
not I_77109 (I1314458,I1314450);
not I_77110 (I1314475,I1354141);
or I_77111 (I1314492,I1354150,I1354141);
nor I_77112 (I1314509,I1354150,I1354141);
or I_77113 (I1314526,I1354147,I1354150);
DFFARX1 I_77114 (I1314526,I3563,I1314373,I1314365,);
not I_77115 (I1314557,I1354159);
nand I_77116 (I1314574,I1314557,I1354138);
nand I_77117 (I1314591,I1314475,I1314574);
and I_77118 (I1314344,I1314458,I1314591);
nor I_77119 (I1314622,I1354159,I1354144);
and I_77120 (I1314639,I1314458,I1314622);
nor I_77121 (I1314350,I1314424,I1314639);
DFFARX1 I_77122 (I1314622,I3563,I1314373,I1314679,);
not I_77123 (I1314687,I1314679);
nor I_77124 (I1314359,I1314458,I1314687);
or I_77125 (I1314718,I1314526,I1354165);
nor I_77126 (I1314735,I1354165,I1354147);
nand I_77127 (I1314752,I1314591,I1314735);
nand I_77128 (I1314769,I1314718,I1314752);
DFFARX1 I_77129 (I1314769,I3563,I1314373,I1314362,);
nor I_77130 (I1314800,I1314735,I1314492);
DFFARX1 I_77131 (I1314800,I3563,I1314373,I1314341,);
nor I_77132 (I1314831,I1354165,I1354156);
DFFARX1 I_77133 (I1314831,I3563,I1314373,I1314857,);
DFFARX1 I_77134 (I1314857,I3563,I1314373,I1314356,);
not I_77135 (I1314879,I1314857);
nand I_77136 (I1314353,I1314879,I1314407);
nand I_77137 (I1314347,I1314879,I1314509);
not I_77138 (I1314951,I3570);
DFFARX1 I_77139 (I568551,I3563,I1314951,I1314977,);
nand I_77140 (I1314985,I1314977,I568560);
not I_77141 (I1315002,I1314985);
DFFARX1 I_77142 (I568572,I3563,I1314951,I1315028,);
not I_77143 (I1315036,I1315028);
not I_77144 (I1315053,I568563);
or I_77145 (I1315070,I568557,I568563);
nor I_77146 (I1315087,I568557,I568563);
or I_77147 (I1315104,I568551,I568557);
DFFARX1 I_77148 (I1315104,I3563,I1314951,I1314943,);
not I_77149 (I1315135,I568554);
nand I_77150 (I1315152,I1315135,I568566);
nand I_77151 (I1315169,I1315053,I1315152);
and I_77152 (I1314922,I1315036,I1315169);
nor I_77153 (I1315200,I568554,I568575);
and I_77154 (I1315217,I1315036,I1315200);
nor I_77155 (I1314928,I1315002,I1315217);
DFFARX1 I_77156 (I1315200,I3563,I1314951,I1315257,);
not I_77157 (I1315265,I1315257);
nor I_77158 (I1314937,I1315036,I1315265);
or I_77159 (I1315296,I1315104,I568569);
nor I_77160 (I1315313,I568569,I568551);
nand I_77161 (I1315330,I1315169,I1315313);
nand I_77162 (I1315347,I1315296,I1315330);
DFFARX1 I_77163 (I1315347,I3563,I1314951,I1314940,);
nor I_77164 (I1315378,I1315313,I1315070);
DFFARX1 I_77165 (I1315378,I3563,I1314951,I1314919,);
nor I_77166 (I1315409,I568569,I568554);
DFFARX1 I_77167 (I1315409,I3563,I1314951,I1315435,);
DFFARX1 I_77168 (I1315435,I3563,I1314951,I1314934,);
not I_77169 (I1315457,I1315435);
nand I_77170 (I1314931,I1315457,I1314985);
nand I_77171 (I1314925,I1315457,I1315087);
not I_77172 (I1315529,I3570);
DFFARX1 I_77173 (I1163263,I3563,I1315529,I1315555,);
nand I_77174 (I1315563,I1315555,I1163248);
not I_77175 (I1315580,I1315563);
DFFARX1 I_77176 (I1163251,I3563,I1315529,I1315606,);
not I_77177 (I1315614,I1315606);
not I_77178 (I1315631,I1163266);
or I_77179 (I1315648,I1163269,I1163266);
nor I_77180 (I1315665,I1163269,I1163266);
or I_77181 (I1315682,I1163245,I1163269);
DFFARX1 I_77182 (I1315682,I3563,I1315529,I1315521,);
not I_77183 (I1315713,I1163257);
nand I_77184 (I1315730,I1315713,I1163260);
nand I_77185 (I1315747,I1315631,I1315730);
and I_77186 (I1315500,I1315614,I1315747);
nor I_77187 (I1315778,I1163257,I1163254);
and I_77188 (I1315795,I1315614,I1315778);
nor I_77189 (I1315506,I1315580,I1315795);
DFFARX1 I_77190 (I1315778,I3563,I1315529,I1315835,);
not I_77191 (I1315843,I1315835);
nor I_77192 (I1315515,I1315614,I1315843);
or I_77193 (I1315874,I1315682,I1163245);
nor I_77194 (I1315891,I1163245,I1163245);
nand I_77195 (I1315908,I1315747,I1315891);
nand I_77196 (I1315925,I1315874,I1315908);
DFFARX1 I_77197 (I1315925,I3563,I1315529,I1315518,);
nor I_77198 (I1315956,I1315891,I1315648);
DFFARX1 I_77199 (I1315956,I3563,I1315529,I1315497,);
nor I_77200 (I1315987,I1163245,I1163248);
DFFARX1 I_77201 (I1315987,I3563,I1315529,I1316013,);
DFFARX1 I_77202 (I1316013,I3563,I1315529,I1315512,);
not I_77203 (I1316035,I1316013);
nand I_77204 (I1315509,I1316035,I1315563);
nand I_77205 (I1315503,I1316035,I1315665);
not I_77206 (I1316107,I3570);
DFFARX1 I_77207 (I1050034,I3563,I1316107,I1316133,);
nand I_77208 (I1316141,I1316133,I1050031);
not I_77209 (I1316158,I1316141);
DFFARX1 I_77210 (I1050031,I3563,I1316107,I1316184,);
not I_77211 (I1316192,I1316184);
not I_77212 (I1316209,I1050028);
or I_77213 (I1316226,I1050037,I1050028);
nor I_77214 (I1316243,I1050037,I1050028);
or I_77215 (I1316260,I1050040,I1050037);
DFFARX1 I_77216 (I1316260,I3563,I1316107,I1316099,);
not I_77217 (I1316291,I1050028);
nand I_77218 (I1316308,I1316291,I1050025);
nand I_77219 (I1316325,I1316209,I1316308);
and I_77220 (I1316078,I1316192,I1316325);
nor I_77221 (I1316356,I1050028,I1050043);
and I_77222 (I1316373,I1316192,I1316356);
nor I_77223 (I1316084,I1316158,I1316373);
DFFARX1 I_77224 (I1316356,I3563,I1316107,I1316413,);
not I_77225 (I1316421,I1316413);
nor I_77226 (I1316093,I1316192,I1316421);
or I_77227 (I1316452,I1316260,I1050046);
nor I_77228 (I1316469,I1050046,I1050040);
nand I_77229 (I1316486,I1316325,I1316469);
nand I_77230 (I1316503,I1316452,I1316486);
DFFARX1 I_77231 (I1316503,I3563,I1316107,I1316096,);
nor I_77232 (I1316534,I1316469,I1316226);
DFFARX1 I_77233 (I1316534,I3563,I1316107,I1316075,);
nor I_77234 (I1316565,I1050046,I1050025);
DFFARX1 I_77235 (I1316565,I3563,I1316107,I1316591,);
DFFARX1 I_77236 (I1316591,I3563,I1316107,I1316090,);
not I_77237 (I1316613,I1316591);
nand I_77238 (I1316087,I1316613,I1316141);
nand I_77239 (I1316081,I1316613,I1316243);
not I_77240 (I1316685,I3570);
DFFARX1 I_77241 (I58767,I3563,I1316685,I1316711,);
nand I_77242 (I1316719,I1316711,I58758);
not I_77243 (I1316736,I1316719);
DFFARX1 I_77244 (I58755,I3563,I1316685,I1316762,);
not I_77245 (I1316770,I1316762);
not I_77246 (I1316787,I58764);
or I_77247 (I1316804,I58755,I58764);
nor I_77248 (I1316821,I58755,I58764);
or I_77249 (I1316838,I58761,I58755);
DFFARX1 I_77250 (I1316838,I3563,I1316685,I1316677,);
not I_77251 (I1316869,I58770);
nand I_77252 (I1316886,I1316869,I58779);
nand I_77253 (I1316903,I1316787,I1316886);
and I_77254 (I1316656,I1316770,I1316903);
nor I_77255 (I1316934,I58770,I58773);
and I_77256 (I1316951,I1316770,I1316934);
nor I_77257 (I1316662,I1316736,I1316951);
DFFARX1 I_77258 (I1316934,I3563,I1316685,I1316991,);
not I_77259 (I1316999,I1316991);
nor I_77260 (I1316671,I1316770,I1316999);
or I_77261 (I1317030,I1316838,I58758);
nor I_77262 (I1317047,I58758,I58761);
nand I_77263 (I1317064,I1316903,I1317047);
nand I_77264 (I1317081,I1317030,I1317064);
DFFARX1 I_77265 (I1317081,I3563,I1316685,I1316674,);
nor I_77266 (I1317112,I1317047,I1316804);
DFFARX1 I_77267 (I1317112,I3563,I1316685,I1316653,);
nor I_77268 (I1317143,I58758,I58776);
DFFARX1 I_77269 (I1317143,I3563,I1316685,I1317169,);
DFFARX1 I_77270 (I1317169,I3563,I1316685,I1316668,);
not I_77271 (I1317191,I1317169);
nand I_77272 (I1316665,I1317191,I1316719);
nand I_77273 (I1316659,I1317191,I1316821);
not I_77274 (I1317263,I3570);
DFFARX1 I_77275 (I966561,I3563,I1317263,I1317289,);
nand I_77276 (I1317297,I1317289,I966582);
not I_77277 (I1317314,I1317297);
DFFARX1 I_77278 (I966555,I3563,I1317263,I1317340,);
not I_77279 (I1317348,I1317340);
not I_77280 (I1317365,I966576);
or I_77281 (I1317382,I966567,I966576);
nor I_77282 (I1317399,I966567,I966576);
or I_77283 (I1317416,I966570,I966567);
DFFARX1 I_77284 (I1317416,I3563,I1317263,I1317255,);
not I_77285 (I1317447,I966558);
nand I_77286 (I1317464,I1317447,I966573);
nand I_77287 (I1317481,I1317365,I1317464);
and I_77288 (I1317234,I1317348,I1317481);
nor I_77289 (I1317512,I966558,I966555);
and I_77290 (I1317529,I1317348,I1317512);
nor I_77291 (I1317240,I1317314,I1317529);
DFFARX1 I_77292 (I1317512,I3563,I1317263,I1317569,);
not I_77293 (I1317577,I1317569);
nor I_77294 (I1317249,I1317348,I1317577);
or I_77295 (I1317608,I1317416,I966579);
nor I_77296 (I1317625,I966579,I966570);
nand I_77297 (I1317642,I1317481,I1317625);
nand I_77298 (I1317659,I1317608,I1317642);
DFFARX1 I_77299 (I1317659,I3563,I1317263,I1317252,);
nor I_77300 (I1317690,I1317625,I1317382);
DFFARX1 I_77301 (I1317690,I3563,I1317263,I1317231,);
nor I_77302 (I1317721,I966579,I966564);
DFFARX1 I_77303 (I1317721,I3563,I1317263,I1317747,);
DFFARX1 I_77304 (I1317747,I3563,I1317263,I1317246,);
not I_77305 (I1317769,I1317747);
nand I_77306 (I1317243,I1317769,I1317297);
nand I_77307 (I1317237,I1317769,I1317399);
not I_77308 (I1317841,I3570);
DFFARX1 I_77309 (I687891,I3563,I1317841,I1317867,);
nand I_77310 (I1317875,I1317867,I687894);
not I_77311 (I1317892,I1317875);
DFFARX1 I_77312 (I687906,I3563,I1317841,I1317918,);
not I_77313 (I1317926,I1317918);
not I_77314 (I1317943,I687891);
or I_77315 (I1317960,I687900,I687891);
nor I_77316 (I1317977,I687900,I687891);
or I_77317 (I1317994,I687909,I687900);
DFFARX1 I_77318 (I1317994,I3563,I1317841,I1317833,);
not I_77319 (I1318025,I687912);
nand I_77320 (I1318042,I1318025,I687894);
nand I_77321 (I1318059,I1317943,I1318042);
and I_77322 (I1317812,I1317926,I1318059);
nor I_77323 (I1318090,I687912,I687897);
and I_77324 (I1318107,I1317926,I1318090);
nor I_77325 (I1317818,I1317892,I1318107);
DFFARX1 I_77326 (I1318090,I3563,I1317841,I1318147,);
not I_77327 (I1318155,I1318147);
nor I_77328 (I1317827,I1317926,I1318155);
or I_77329 (I1318186,I1317994,I687903);
nor I_77330 (I1318203,I687903,I687909);
nand I_77331 (I1318220,I1318059,I1318203);
nand I_77332 (I1318237,I1318186,I1318220);
DFFARX1 I_77333 (I1318237,I3563,I1317841,I1317830,);
nor I_77334 (I1318268,I1318203,I1317960);
DFFARX1 I_77335 (I1318268,I3563,I1317841,I1317809,);
nor I_77336 (I1318299,I687903,I687915);
DFFARX1 I_77337 (I1318299,I3563,I1317841,I1318325,);
DFFARX1 I_77338 (I1318325,I3563,I1317841,I1317824,);
not I_77339 (I1318347,I1318325);
nand I_77340 (I1317821,I1318347,I1317875);
nand I_77341 (I1317815,I1318347,I1317977);
not I_77342 (I1318419,I3570);
DFFARX1 I_77343 (I545346,I3563,I1318419,I1318445,);
nand I_77344 (I1318453,I1318445,I545355);
not I_77345 (I1318470,I1318453);
DFFARX1 I_77346 (I545367,I3563,I1318419,I1318496,);
not I_77347 (I1318504,I1318496);
not I_77348 (I1318521,I545358);
or I_77349 (I1318538,I545352,I545358);
nor I_77350 (I1318555,I545352,I545358);
or I_77351 (I1318572,I545346,I545352);
DFFARX1 I_77352 (I1318572,I3563,I1318419,I1318411,);
not I_77353 (I1318603,I545349);
nand I_77354 (I1318620,I1318603,I545361);
nand I_77355 (I1318637,I1318521,I1318620);
and I_77356 (I1318390,I1318504,I1318637);
nor I_77357 (I1318668,I545349,I545370);
and I_77358 (I1318685,I1318504,I1318668);
nor I_77359 (I1318396,I1318470,I1318685);
DFFARX1 I_77360 (I1318668,I3563,I1318419,I1318725,);
not I_77361 (I1318733,I1318725);
nor I_77362 (I1318405,I1318504,I1318733);
or I_77363 (I1318764,I1318572,I545364);
nor I_77364 (I1318781,I545364,I545346);
nand I_77365 (I1318798,I1318637,I1318781);
nand I_77366 (I1318815,I1318764,I1318798);
DFFARX1 I_77367 (I1318815,I3563,I1318419,I1318408,);
nor I_77368 (I1318846,I1318781,I1318538);
DFFARX1 I_77369 (I1318846,I3563,I1318419,I1318387,);
nor I_77370 (I1318877,I545364,I545349);
DFFARX1 I_77371 (I1318877,I3563,I1318419,I1318903,);
DFFARX1 I_77372 (I1318903,I3563,I1318419,I1318402,);
not I_77373 (I1318925,I1318903);
nand I_77374 (I1318399,I1318925,I1318453);
nand I_77375 (I1318393,I1318925,I1318555);
not I_77376 (I1318997,I3570);
DFFARX1 I_77377 (I1338692,I3563,I1318997,I1319023,);
nand I_77378 (I1319031,I1319023,I1338683);
not I_77379 (I1319048,I1319031);
DFFARX1 I_77380 (I1338668,I3563,I1318997,I1319074,);
not I_77381 (I1319082,I1319074);
not I_77382 (I1319099,I1338671);
or I_77383 (I1319116,I1338680,I1338671);
nor I_77384 (I1319133,I1338680,I1338671);
or I_77385 (I1319150,I1338677,I1338680);
DFFARX1 I_77386 (I1319150,I3563,I1318997,I1318989,);
not I_77387 (I1319181,I1338689);
nand I_77388 (I1319198,I1319181,I1338668);
nand I_77389 (I1319215,I1319099,I1319198);
and I_77390 (I1318968,I1319082,I1319215);
nor I_77391 (I1319246,I1338689,I1338674);
and I_77392 (I1319263,I1319082,I1319246);
nor I_77393 (I1318974,I1319048,I1319263);
DFFARX1 I_77394 (I1319246,I3563,I1318997,I1319303,);
not I_77395 (I1319311,I1319303);
nor I_77396 (I1318983,I1319082,I1319311);
or I_77397 (I1319342,I1319150,I1338695);
nor I_77398 (I1319359,I1338695,I1338677);
nand I_77399 (I1319376,I1319215,I1319359);
nand I_77400 (I1319393,I1319342,I1319376);
DFFARX1 I_77401 (I1319393,I3563,I1318997,I1318986,);
nor I_77402 (I1319424,I1319359,I1319116);
DFFARX1 I_77403 (I1319424,I3563,I1318997,I1318965,);
nor I_77404 (I1319455,I1338695,I1338686);
DFFARX1 I_77405 (I1319455,I3563,I1318997,I1319481,);
DFFARX1 I_77406 (I1319481,I3563,I1318997,I1318980,);
not I_77407 (I1319503,I1319481);
nand I_77408 (I1318977,I1319503,I1319031);
nand I_77409 (I1318971,I1319503,I1319133);
not I_77410 (I1319575,I3570);
DFFARX1 I_77411 (I376542,I3563,I1319575,I1319601,);
nand I_77412 (I1319609,I1319601,I376563);
not I_77413 (I1319626,I1319609);
DFFARX1 I_77414 (I376557,I3563,I1319575,I1319652,);
not I_77415 (I1319660,I1319652);
not I_77416 (I1319677,I376545);
or I_77417 (I1319694,I376560,I376545);
nor I_77418 (I1319711,I376560,I376545);
or I_77419 (I1319728,I376551,I376560);
DFFARX1 I_77420 (I1319728,I3563,I1319575,I1319567,);
not I_77421 (I1319759,I376539);
nand I_77422 (I1319776,I1319759,I376536);
nand I_77423 (I1319793,I1319677,I1319776);
and I_77424 (I1319546,I1319660,I1319793);
nor I_77425 (I1319824,I376539,I376548);
and I_77426 (I1319841,I1319660,I1319824);
nor I_77427 (I1319552,I1319626,I1319841);
DFFARX1 I_77428 (I1319824,I3563,I1319575,I1319881,);
not I_77429 (I1319889,I1319881);
nor I_77430 (I1319561,I1319660,I1319889);
or I_77431 (I1319920,I1319728,I376554);
nor I_77432 (I1319937,I376554,I376551);
nand I_77433 (I1319954,I1319793,I1319937);
nand I_77434 (I1319971,I1319920,I1319954);
DFFARX1 I_77435 (I1319971,I3563,I1319575,I1319564,);
nor I_77436 (I1320002,I1319937,I1319694);
DFFARX1 I_77437 (I1320002,I3563,I1319575,I1319543,);
nor I_77438 (I1320033,I376554,I376536);
DFFARX1 I_77439 (I1320033,I3563,I1319575,I1320059,);
DFFARX1 I_77440 (I1320059,I3563,I1319575,I1319558,);
not I_77441 (I1320081,I1320059);
nand I_77442 (I1319555,I1320081,I1319609);
nand I_77443 (I1319549,I1320081,I1319711);
not I_77444 (I1320153,I3570);
DFFARX1 I_77445 (I1188695,I3563,I1320153,I1320179,);
nand I_77446 (I1320187,I1320179,I1188680);
not I_77447 (I1320204,I1320187);
DFFARX1 I_77448 (I1188683,I3563,I1320153,I1320230,);
not I_77449 (I1320238,I1320230);
not I_77450 (I1320255,I1188698);
or I_77451 (I1320272,I1188701,I1188698);
nor I_77452 (I1320289,I1188701,I1188698);
or I_77453 (I1320306,I1188677,I1188701);
DFFARX1 I_77454 (I1320306,I3563,I1320153,I1320145,);
not I_77455 (I1320337,I1188689);
nand I_77456 (I1320354,I1320337,I1188692);
nand I_77457 (I1320371,I1320255,I1320354);
and I_77458 (I1320124,I1320238,I1320371);
nor I_77459 (I1320402,I1188689,I1188686);
and I_77460 (I1320419,I1320238,I1320402);
nor I_77461 (I1320130,I1320204,I1320419);
DFFARX1 I_77462 (I1320402,I3563,I1320153,I1320459,);
not I_77463 (I1320467,I1320459);
nor I_77464 (I1320139,I1320238,I1320467);
or I_77465 (I1320498,I1320306,I1188677);
nor I_77466 (I1320515,I1188677,I1188677);
nand I_77467 (I1320532,I1320371,I1320515);
nand I_77468 (I1320549,I1320498,I1320532);
DFFARX1 I_77469 (I1320549,I3563,I1320153,I1320142,);
nor I_77470 (I1320580,I1320515,I1320272);
DFFARX1 I_77471 (I1320580,I3563,I1320153,I1320121,);
nor I_77472 (I1320611,I1188677,I1188680);
DFFARX1 I_77473 (I1320611,I3563,I1320153,I1320637,);
DFFARX1 I_77474 (I1320637,I3563,I1320153,I1320136,);
not I_77475 (I1320659,I1320637);
nand I_77476 (I1320133,I1320659,I1320187);
nand I_77477 (I1320127,I1320659,I1320289);
not I_77478 (I1320731,I3570);
DFFARX1 I_77479 (I1047790,I3563,I1320731,I1320757,);
nand I_77480 (I1320765,I1320757,I1047787);
not I_77481 (I1320782,I1320765);
DFFARX1 I_77482 (I1047787,I3563,I1320731,I1320808,);
not I_77483 (I1320816,I1320808);
not I_77484 (I1320833,I1047784);
or I_77485 (I1320850,I1047793,I1047784);
nor I_77486 (I1320867,I1047793,I1047784);
or I_77487 (I1320884,I1047796,I1047793);
DFFARX1 I_77488 (I1320884,I3563,I1320731,I1320723,);
not I_77489 (I1320915,I1047784);
nand I_77490 (I1320932,I1320915,I1047781);
nand I_77491 (I1320949,I1320833,I1320932);
and I_77492 (I1320702,I1320816,I1320949);
nor I_77493 (I1320980,I1047784,I1047799);
and I_77494 (I1320997,I1320816,I1320980);
nor I_77495 (I1320708,I1320782,I1320997);
DFFARX1 I_77496 (I1320980,I3563,I1320731,I1321037,);
not I_77497 (I1321045,I1321037);
nor I_77498 (I1320717,I1320816,I1321045);
or I_77499 (I1321076,I1320884,I1047802);
nor I_77500 (I1321093,I1047802,I1047796);
nand I_77501 (I1321110,I1320949,I1321093);
nand I_77502 (I1321127,I1321076,I1321110);
DFFARX1 I_77503 (I1321127,I3563,I1320731,I1320720,);
nor I_77504 (I1321158,I1321093,I1320850);
DFFARX1 I_77505 (I1321158,I3563,I1320731,I1320699,);
nor I_77506 (I1321189,I1047802,I1047781);
DFFARX1 I_77507 (I1321189,I3563,I1320731,I1321215,);
DFFARX1 I_77508 (I1321215,I3563,I1320731,I1320714,);
not I_77509 (I1321237,I1321215);
nand I_77510 (I1320711,I1321237,I1320765);
nand I_77511 (I1320705,I1321237,I1320867);
not I_77512 (I1321309,I3570);
DFFARX1 I_77513 (I363894,I3563,I1321309,I1321335,);
nand I_77514 (I1321343,I1321335,I363915);
not I_77515 (I1321360,I1321343);
DFFARX1 I_77516 (I363909,I3563,I1321309,I1321386,);
not I_77517 (I1321394,I1321386);
not I_77518 (I1321411,I363897);
or I_77519 (I1321428,I363912,I363897);
nor I_77520 (I1321445,I363912,I363897);
or I_77521 (I1321462,I363903,I363912);
DFFARX1 I_77522 (I1321462,I3563,I1321309,I1321301,);
not I_77523 (I1321493,I363891);
nand I_77524 (I1321510,I1321493,I363888);
nand I_77525 (I1321527,I1321411,I1321510);
and I_77526 (I1321280,I1321394,I1321527);
nor I_77527 (I1321558,I363891,I363900);
and I_77528 (I1321575,I1321394,I1321558);
nor I_77529 (I1321286,I1321360,I1321575);
DFFARX1 I_77530 (I1321558,I3563,I1321309,I1321615,);
not I_77531 (I1321623,I1321615);
nor I_77532 (I1321295,I1321394,I1321623);
or I_77533 (I1321654,I1321462,I363906);
nor I_77534 (I1321671,I363906,I363903);
nand I_77535 (I1321688,I1321527,I1321671);
nand I_77536 (I1321705,I1321654,I1321688);
DFFARX1 I_77537 (I1321705,I3563,I1321309,I1321298,);
nor I_77538 (I1321736,I1321671,I1321428);
DFFARX1 I_77539 (I1321736,I3563,I1321309,I1321277,);
nor I_77540 (I1321767,I363906,I363888);
DFFARX1 I_77541 (I1321767,I3563,I1321309,I1321793,);
DFFARX1 I_77542 (I1321793,I3563,I1321309,I1321292,);
not I_77543 (I1321815,I1321793);
nand I_77544 (I1321289,I1321815,I1321343);
nand I_77545 (I1321283,I1321815,I1321445);
not I_77546 (I1321887,I3570);
DFFARX1 I_77547 (I474629,I3563,I1321887,I1321913,);
nand I_77548 (I1321921,I1321913,I474638);
not I_77549 (I1321938,I1321921);
DFFARX1 I_77550 (I474626,I3563,I1321887,I1321964,);
not I_77551 (I1321972,I1321964);
not I_77552 (I1321989,I474632);
or I_77553 (I1322006,I474626,I474632);
nor I_77554 (I1322023,I474626,I474632);
or I_77555 (I1322040,I474641,I474626);
DFFARX1 I_77556 (I1322040,I3563,I1321887,I1321879,);
not I_77557 (I1322071,I474635);
nand I_77558 (I1322088,I1322071,I474650);
nand I_77559 (I1322105,I1321989,I1322088);
and I_77560 (I1321858,I1321972,I1322105);
nor I_77561 (I1322136,I474635,I474653);
and I_77562 (I1322153,I1321972,I1322136);
nor I_77563 (I1321864,I1321938,I1322153);
DFFARX1 I_77564 (I1322136,I3563,I1321887,I1322193,);
not I_77565 (I1322201,I1322193);
nor I_77566 (I1321873,I1321972,I1322201);
or I_77567 (I1322232,I1322040,I474644);
nor I_77568 (I1322249,I474644,I474641);
nand I_77569 (I1322266,I1322105,I1322249);
nand I_77570 (I1322283,I1322232,I1322266);
DFFARX1 I_77571 (I1322283,I3563,I1321887,I1321876,);
nor I_77572 (I1322314,I1322249,I1322006);
DFFARX1 I_77573 (I1322314,I3563,I1321887,I1321855,);
nor I_77574 (I1322345,I474644,I474647);
DFFARX1 I_77575 (I1322345,I3563,I1321887,I1322371,);
DFFARX1 I_77576 (I1322371,I3563,I1321887,I1321870,);
not I_77577 (I1322393,I1322371);
nand I_77578 (I1321867,I1322393,I1321921);
nand I_77579 (I1321861,I1322393,I1322023);
not I_77580 (I1322465,I3570);
DFFARX1 I_77581 (I254153,I3563,I1322465,I1322491,);
nand I_77582 (I1322499,I1322491,I254156);
not I_77583 (I1322516,I1322499);
DFFARX1 I_77584 (I254165,I3563,I1322465,I1322542,);
not I_77585 (I1322550,I1322542);
not I_77586 (I1322567,I254168);
or I_77587 (I1322584,I254159,I254168);
nor I_77588 (I1322601,I254159,I254168);
or I_77589 (I1322618,I254171,I254159);
DFFARX1 I_77590 (I1322618,I3563,I1322465,I1322457,);
not I_77591 (I1322649,I254156);
nand I_77592 (I1322666,I1322649,I254162);
nand I_77593 (I1322683,I1322567,I1322666);
and I_77594 (I1322436,I1322550,I1322683);
nor I_77595 (I1322714,I254156,I254174);
and I_77596 (I1322731,I1322550,I1322714);
nor I_77597 (I1322442,I1322516,I1322731);
DFFARX1 I_77598 (I1322714,I3563,I1322465,I1322771,);
not I_77599 (I1322779,I1322771);
nor I_77600 (I1322451,I1322550,I1322779);
or I_77601 (I1322810,I1322618,I254153);
nor I_77602 (I1322827,I254153,I254171);
nand I_77603 (I1322844,I1322683,I1322827);
nand I_77604 (I1322861,I1322810,I1322844);
DFFARX1 I_77605 (I1322861,I3563,I1322465,I1322454,);
nor I_77606 (I1322892,I1322827,I1322584);
DFFARX1 I_77607 (I1322892,I3563,I1322465,I1322433,);
nor I_77608 (I1322923,I254153,I254177);
DFFARX1 I_77609 (I1322923,I3563,I1322465,I1322949,);
DFFARX1 I_77610 (I1322949,I3563,I1322465,I1322448,);
not I_77611 (I1322971,I1322949);
nand I_77612 (I1322445,I1322971,I1322499);
nand I_77613 (I1322439,I1322971,I1322601);
not I_77614 (I1323043,I3570);
DFFARX1 I_77615 (I999507,I3563,I1323043,I1323069,);
nand I_77616 (I1323077,I1323069,I999528);
not I_77617 (I1323094,I1323077);
DFFARX1 I_77618 (I999501,I3563,I1323043,I1323120,);
not I_77619 (I1323128,I1323120);
not I_77620 (I1323145,I999522);
or I_77621 (I1323162,I999513,I999522);
nor I_77622 (I1323179,I999513,I999522);
or I_77623 (I1323196,I999516,I999513);
DFFARX1 I_77624 (I1323196,I3563,I1323043,I1323035,);
not I_77625 (I1323227,I999504);
nand I_77626 (I1323244,I1323227,I999519);
nand I_77627 (I1323261,I1323145,I1323244);
and I_77628 (I1323014,I1323128,I1323261);
nor I_77629 (I1323292,I999504,I999501);
and I_77630 (I1323309,I1323128,I1323292);
nor I_77631 (I1323020,I1323094,I1323309);
DFFARX1 I_77632 (I1323292,I3563,I1323043,I1323349,);
not I_77633 (I1323357,I1323349);
nor I_77634 (I1323029,I1323128,I1323357);
or I_77635 (I1323388,I1323196,I999525);
nor I_77636 (I1323405,I999525,I999516);
nand I_77637 (I1323422,I1323261,I1323405);
nand I_77638 (I1323439,I1323388,I1323422);
DFFARX1 I_77639 (I1323439,I3563,I1323043,I1323032,);
nor I_77640 (I1323470,I1323405,I1323162);
DFFARX1 I_77641 (I1323470,I3563,I1323043,I1323011,);
nor I_77642 (I1323501,I999525,I999510);
DFFARX1 I_77643 (I1323501,I3563,I1323043,I1323527,);
DFFARX1 I_77644 (I1323527,I3563,I1323043,I1323026,);
not I_77645 (I1323549,I1323527);
nand I_77646 (I1323023,I1323549,I1323077);
nand I_77647 (I1323017,I1323549,I1323179);
not I_77648 (I1323621,I3570);
DFFARX1 I_77649 (I384447,I3563,I1323621,I1323647,);
nand I_77650 (I1323655,I1323647,I384468);
not I_77651 (I1323672,I1323655);
DFFARX1 I_77652 (I384462,I3563,I1323621,I1323698,);
not I_77653 (I1323706,I1323698);
not I_77654 (I1323723,I384450);
or I_77655 (I1323740,I384465,I384450);
nor I_77656 (I1323757,I384465,I384450);
or I_77657 (I1323774,I384456,I384465);
DFFARX1 I_77658 (I1323774,I3563,I1323621,I1323613,);
not I_77659 (I1323805,I384444);
nand I_77660 (I1323822,I1323805,I384441);
nand I_77661 (I1323839,I1323723,I1323822);
and I_77662 (I1323592,I1323706,I1323839);
nor I_77663 (I1323870,I384444,I384453);
and I_77664 (I1323887,I1323706,I1323870);
nor I_77665 (I1323598,I1323672,I1323887);
DFFARX1 I_77666 (I1323870,I3563,I1323621,I1323927,);
not I_77667 (I1323935,I1323927);
nor I_77668 (I1323607,I1323706,I1323935);
or I_77669 (I1323966,I1323774,I384459);
nor I_77670 (I1323983,I384459,I384456);
nand I_77671 (I1324000,I1323839,I1323983);
nand I_77672 (I1324017,I1323966,I1324000);
DFFARX1 I_77673 (I1324017,I3563,I1323621,I1323610,);
nor I_77674 (I1324048,I1323983,I1323740);
DFFARX1 I_77675 (I1324048,I3563,I1323621,I1323589,);
nor I_77676 (I1324079,I384459,I384441);
DFFARX1 I_77677 (I1324079,I3563,I1323621,I1324105,);
DFFARX1 I_77678 (I1324105,I3563,I1323621,I1323604,);
not I_77679 (I1324127,I1324105);
nand I_77680 (I1323601,I1324127,I1323655);
nand I_77681 (I1323595,I1324127,I1323757);
not I_77682 (I1324202,I3570);
DFFARX1 I_77683 (I130978,I3563,I1324202,I1324228,);
nand I_77684 (I1324236,I1324228,I130969);
not I_77685 (I1324253,I1324236);
DFFARX1 I_77686 (I130957,I3563,I1324202,I1324279,);
not I_77687 (I1324287,I1324279);
nor I_77688 (I1324304,I130960,I130957);
not I_77689 (I1324321,I1324304);
DFFARX1 I_77690 (I1324321,I3563,I1324202,I1324188,);
or I_77691 (I1324352,I130954,I130960);
DFFARX1 I_77692 (I1324352,I3563,I1324202,I1324191,);
not I_77693 (I1324383,I130963);
nor I_77694 (I1324400,I1324383,I130954);
nor I_77695 (I1324417,I1324400,I130957);
nor I_77696 (I1324434,I130954,I130966);
nor I_77697 (I1324451,I1324287,I1324434);
nor I_77698 (I1324176,I1324253,I1324451);
not I_77699 (I1324482,I1324434);
nand I_77700 (I1324179,I1324482,I1324236);
nand I_77701 (I1324173,I1324482,I1324304);
nor I_77702 (I1324170,I1324434,I1324417);
nor I_77703 (I1324541,I130972,I130954);
not I_77704 (I1324558,I1324541);
DFFARX1 I_77705 (I1324541,I3563,I1324202,I1324584,);
not I_77706 (I1324194,I1324584);
nor I_77707 (I1324606,I130972,I130975);
DFFARX1 I_77708 (I1324606,I3563,I1324202,I1324632,);
and I_77709 (I1324640,I1324632,I130960);
nor I_77710 (I1324657,I1324640,I1324558);
DFFARX1 I_77711 (I1324657,I3563,I1324202,I1324185,);
nor I_77712 (I1324688,I1324632,I1324417);
DFFARX1 I_77713 (I1324688,I3563,I1324202,I1324167,);
nor I_77714 (I1324182,I1324632,I1324321);
not I_77715 (I1324763,I3570);
DFFARX1 I_77716 (I145207,I3563,I1324763,I1324789,);
nand I_77717 (I1324797,I1324789,I145198);
not I_77718 (I1324814,I1324797);
DFFARX1 I_77719 (I145186,I3563,I1324763,I1324840,);
not I_77720 (I1324848,I1324840);
nor I_77721 (I1324865,I145189,I145186);
not I_77722 (I1324882,I1324865);
DFFARX1 I_77723 (I1324882,I3563,I1324763,I1324749,);
or I_77724 (I1324913,I145183,I145189);
DFFARX1 I_77725 (I1324913,I3563,I1324763,I1324752,);
not I_77726 (I1324944,I145192);
nor I_77727 (I1324961,I1324944,I145183);
nor I_77728 (I1324978,I1324961,I145186);
nor I_77729 (I1324995,I145183,I145195);
nor I_77730 (I1325012,I1324848,I1324995);
nor I_77731 (I1324737,I1324814,I1325012);
not I_77732 (I1325043,I1324995);
nand I_77733 (I1324740,I1325043,I1324797);
nand I_77734 (I1324734,I1325043,I1324865);
nor I_77735 (I1324731,I1324995,I1324978);
nor I_77736 (I1325102,I145201,I145183);
not I_77737 (I1325119,I1325102);
DFFARX1 I_77738 (I1325102,I3563,I1324763,I1325145,);
not I_77739 (I1324755,I1325145);
nor I_77740 (I1325167,I145201,I145204);
DFFARX1 I_77741 (I1325167,I3563,I1324763,I1325193,);
and I_77742 (I1325201,I1325193,I145189);
nor I_77743 (I1325218,I1325201,I1325119);
DFFARX1 I_77744 (I1325218,I3563,I1324763,I1324746,);
nor I_77745 (I1325249,I1325193,I1324978);
DFFARX1 I_77746 (I1325249,I3563,I1324763,I1324728,);
nor I_77747 (I1324743,I1325193,I1324882);
not I_77748 (I1325324,I3570);
DFFARX1 I_77749 (I1139550,I3563,I1325324,I1325350,);
nand I_77750 (I1325358,I1325350,I1139547);
not I_77751 (I1325375,I1325358);
DFFARX1 I_77752 (I1139550,I3563,I1325324,I1325401,);
not I_77753 (I1325409,I1325401);
nor I_77754 (I1325426,I1139568,I1139562);
not I_77755 (I1325443,I1325426);
DFFARX1 I_77756 (I1325443,I3563,I1325324,I1325310,);
or I_77757 (I1325474,I1139571,I1139568);
DFFARX1 I_77758 (I1325474,I3563,I1325324,I1325313,);
not I_77759 (I1325505,I1139559);
nor I_77760 (I1325522,I1325505,I1139556);
nor I_77761 (I1325539,I1325522,I1139562);
nor I_77762 (I1325556,I1139556,I1139547);
nor I_77763 (I1325573,I1325409,I1325556);
nor I_77764 (I1325298,I1325375,I1325573);
not I_77765 (I1325604,I1325556);
nand I_77766 (I1325301,I1325604,I1325358);
nand I_77767 (I1325295,I1325604,I1325426);
nor I_77768 (I1325292,I1325556,I1325539);
nor I_77769 (I1325663,I1139553,I1139571);
not I_77770 (I1325680,I1325663);
DFFARX1 I_77771 (I1325663,I3563,I1325324,I1325706,);
not I_77772 (I1325316,I1325706);
nor I_77773 (I1325728,I1139553,I1139565);
DFFARX1 I_77774 (I1325728,I3563,I1325324,I1325754,);
and I_77775 (I1325762,I1325754,I1139568);
nor I_77776 (I1325779,I1325762,I1325680);
DFFARX1 I_77777 (I1325779,I3563,I1325324,I1325307,);
nor I_77778 (I1325810,I1325754,I1325539);
DFFARX1 I_77779 (I1325810,I3563,I1325324,I1325289,);
nor I_77780 (I1325304,I1325754,I1325443);
not I_77781 (I1325885,I3570);
DFFARX1 I_77782 (I827923,I3563,I1325885,I1325911,);
nand I_77783 (I1325919,I1325911,I827941);
not I_77784 (I1325936,I1325919);
DFFARX1 I_77785 (I827920,I3563,I1325885,I1325962,);
not I_77786 (I1325970,I1325962);
nor I_77787 (I1325987,I827935,I827929);
not I_77788 (I1326004,I1325987);
DFFARX1 I_77789 (I1326004,I3563,I1325885,I1325871,);
or I_77790 (I1326035,I827926,I827935);
DFFARX1 I_77791 (I1326035,I3563,I1325885,I1325874,);
not I_77792 (I1326066,I827926);
nor I_77793 (I1326083,I1326066,I827932);
nor I_77794 (I1326100,I1326083,I827929);
nor I_77795 (I1326117,I827932,I827920);
nor I_77796 (I1326134,I1325970,I1326117);
nor I_77797 (I1325859,I1325936,I1326134);
not I_77798 (I1326165,I1326117);
nand I_77799 (I1325862,I1326165,I1325919);
nand I_77800 (I1325856,I1326165,I1325987);
nor I_77801 (I1325853,I1326117,I1326100);
nor I_77802 (I1326224,I827923,I827926);
not I_77803 (I1326241,I1326224);
DFFARX1 I_77804 (I1326224,I3563,I1325885,I1326267,);
not I_77805 (I1325877,I1326267);
nor I_77806 (I1326289,I827923,I827938);
DFFARX1 I_77807 (I1326289,I3563,I1325885,I1326315,);
and I_77808 (I1326323,I1326315,I827935);
nor I_77809 (I1326340,I1326323,I1326241);
DFFARX1 I_77810 (I1326340,I3563,I1325885,I1325868,);
nor I_77811 (I1326371,I1326315,I1326100);
DFFARX1 I_77812 (I1326371,I3563,I1325885,I1325850,);
nor I_77813 (I1325865,I1326315,I1326004);
not I_77814 (I1326446,I3570);
DFFARX1 I_77815 (I103574,I3563,I1326446,I1326472,);
nand I_77816 (I1326480,I1326472,I103565);
not I_77817 (I1326497,I1326480);
DFFARX1 I_77818 (I103553,I3563,I1326446,I1326523,);
not I_77819 (I1326531,I1326523);
nor I_77820 (I1326548,I103556,I103553);
not I_77821 (I1326565,I1326548);
DFFARX1 I_77822 (I1326565,I3563,I1326446,I1326432,);
or I_77823 (I1326596,I103550,I103556);
DFFARX1 I_77824 (I1326596,I3563,I1326446,I1326435,);
not I_77825 (I1326627,I103559);
nor I_77826 (I1326644,I1326627,I103550);
nor I_77827 (I1326661,I1326644,I103553);
nor I_77828 (I1326678,I103550,I103562);
nor I_77829 (I1326695,I1326531,I1326678);
nor I_77830 (I1326420,I1326497,I1326695);
not I_77831 (I1326726,I1326678);
nand I_77832 (I1326423,I1326726,I1326480);
nand I_77833 (I1326417,I1326726,I1326548);
nor I_77834 (I1326414,I1326678,I1326661);
nor I_77835 (I1326785,I103568,I103550);
not I_77836 (I1326802,I1326785);
DFFARX1 I_77837 (I1326785,I3563,I1326446,I1326828,);
not I_77838 (I1326438,I1326828);
nor I_77839 (I1326850,I103568,I103571);
DFFARX1 I_77840 (I1326850,I3563,I1326446,I1326876,);
and I_77841 (I1326884,I1326876,I103556);
nor I_77842 (I1326901,I1326884,I1326802);
DFFARX1 I_77843 (I1326901,I3563,I1326446,I1326429,);
nor I_77844 (I1326932,I1326876,I1326661);
DFFARX1 I_77845 (I1326932,I3563,I1326446,I1326411,);
nor I_77846 (I1326426,I1326876,I1326565);
not I_77847 (I1327007,I3570);
DFFARX1 I_77848 (I106736,I3563,I1327007,I1327033,);
nand I_77849 (I1327041,I1327033,I106727);
not I_77850 (I1327058,I1327041);
DFFARX1 I_77851 (I106715,I3563,I1327007,I1327084,);
not I_77852 (I1327092,I1327084);
nor I_77853 (I1327109,I106718,I106715);
not I_77854 (I1327126,I1327109);
DFFARX1 I_77855 (I1327126,I3563,I1327007,I1326993,);
or I_77856 (I1327157,I106712,I106718);
DFFARX1 I_77857 (I1327157,I3563,I1327007,I1326996,);
not I_77858 (I1327188,I106721);
nor I_77859 (I1327205,I1327188,I106712);
nor I_77860 (I1327222,I1327205,I106715);
nor I_77861 (I1327239,I106712,I106724);
nor I_77862 (I1327256,I1327092,I1327239);
nor I_77863 (I1326981,I1327058,I1327256);
not I_77864 (I1327287,I1327239);
nand I_77865 (I1326984,I1327287,I1327041);
nand I_77866 (I1326978,I1327287,I1327109);
nor I_77867 (I1326975,I1327239,I1327222);
nor I_77868 (I1327346,I106730,I106712);
not I_77869 (I1327363,I1327346);
DFFARX1 I_77870 (I1327346,I3563,I1327007,I1327389,);
not I_77871 (I1326999,I1327389);
nor I_77872 (I1327411,I106730,I106733);
DFFARX1 I_77873 (I1327411,I3563,I1327007,I1327437,);
and I_77874 (I1327445,I1327437,I106718);
nor I_77875 (I1327462,I1327445,I1327363);
DFFARX1 I_77876 (I1327462,I3563,I1327007,I1326990,);
nor I_77877 (I1327493,I1327437,I1327222);
DFFARX1 I_77878 (I1327493,I3563,I1327007,I1326972,);
nor I_77879 (I1326987,I1327437,I1327126);
not I_77880 (I1327568,I3570);
DFFARX1 I_77881 (I591967,I3563,I1327568,I1327594,);
nand I_77882 (I1327602,I1327594,I591946);
not I_77883 (I1327619,I1327602);
DFFARX1 I_77884 (I591958,I3563,I1327568,I1327645,);
not I_77885 (I1327653,I1327645);
nor I_77886 (I1327670,I591946,I591955);
not I_77887 (I1327687,I1327670);
DFFARX1 I_77888 (I1327687,I3563,I1327568,I1327554,);
or I_77889 (I1327718,I591949,I591946);
DFFARX1 I_77890 (I1327718,I3563,I1327568,I1327557,);
not I_77891 (I1327749,I591952);
nor I_77892 (I1327766,I1327749,I591943);
nor I_77893 (I1327783,I1327766,I591955);
nor I_77894 (I1327800,I591943,I591961);
nor I_77895 (I1327817,I1327653,I1327800);
nor I_77896 (I1327542,I1327619,I1327817);
not I_77897 (I1327848,I1327800);
nand I_77898 (I1327545,I1327848,I1327602);
nand I_77899 (I1327539,I1327848,I1327670);
nor I_77900 (I1327536,I1327800,I1327783);
nor I_77901 (I1327907,I591964,I591949);
not I_77902 (I1327924,I1327907);
DFFARX1 I_77903 (I1327907,I3563,I1327568,I1327950,);
not I_77904 (I1327560,I1327950);
nor I_77905 (I1327972,I591964,I591943);
DFFARX1 I_77906 (I1327972,I3563,I1327568,I1327998,);
and I_77907 (I1328006,I1327998,I591946);
nor I_77908 (I1328023,I1328006,I1327924);
DFFARX1 I_77909 (I1328023,I3563,I1327568,I1327551,);
nor I_77910 (I1328054,I1327998,I1327783);
DFFARX1 I_77911 (I1328054,I3563,I1327568,I1327533,);
nor I_77912 (I1327548,I1327998,I1327687);
not I_77913 (I1328129,I3570);
DFFARX1 I_77914 (I465399,I3563,I1328129,I1328155,);
nand I_77915 (I1328163,I1328155,I465381);
not I_77916 (I1328180,I1328163);
DFFARX1 I_77917 (I465378,I3563,I1328129,I1328206,);
not I_77918 (I1328214,I1328206);
nor I_77919 (I1328231,I465384,I465378);
not I_77920 (I1328248,I1328231);
DFFARX1 I_77921 (I1328248,I3563,I1328129,I1328115,);
or I_77922 (I1328279,I465387,I465384);
DFFARX1 I_77923 (I1328279,I3563,I1328129,I1328118,);
not I_77924 (I1328310,I465393);
nor I_77925 (I1328327,I1328310,I465405);
nor I_77926 (I1328344,I1328327,I465378);
nor I_77927 (I1328361,I465405,I465390);
nor I_77928 (I1328378,I1328214,I1328361);
nor I_77929 (I1328103,I1328180,I1328378);
not I_77930 (I1328409,I1328361);
nand I_77931 (I1328106,I1328409,I1328163);
nand I_77932 (I1328100,I1328409,I1328231);
nor I_77933 (I1328097,I1328361,I1328344);
nor I_77934 (I1328468,I465396,I465387);
not I_77935 (I1328485,I1328468);
DFFARX1 I_77936 (I1328468,I3563,I1328129,I1328511,);
not I_77937 (I1328121,I1328511);
nor I_77938 (I1328533,I465396,I465402);
DFFARX1 I_77939 (I1328533,I3563,I1328129,I1328559,);
and I_77940 (I1328567,I1328559,I465384);
nor I_77941 (I1328584,I1328567,I1328485);
DFFARX1 I_77942 (I1328584,I3563,I1328129,I1328112,);
nor I_77943 (I1328615,I1328559,I1328344);
DFFARX1 I_77944 (I1328615,I3563,I1328129,I1328094,);
nor I_77945 (I1328109,I1328559,I1328248);
not I_77946 (I1328690,I3570);
DFFARX1 I_77947 (I891690,I3563,I1328690,I1328716,);
nand I_77948 (I1328724,I1328716,I891708);
not I_77949 (I1328741,I1328724);
DFFARX1 I_77950 (I891687,I3563,I1328690,I1328767,);
not I_77951 (I1328775,I1328767);
nor I_77952 (I1328792,I891702,I891696);
not I_77953 (I1328809,I1328792);
DFFARX1 I_77954 (I1328809,I3563,I1328690,I1328676,);
or I_77955 (I1328840,I891693,I891702);
DFFARX1 I_77956 (I1328840,I3563,I1328690,I1328679,);
not I_77957 (I1328871,I891693);
nor I_77958 (I1328888,I1328871,I891699);
nor I_77959 (I1328905,I1328888,I891696);
nor I_77960 (I1328922,I891699,I891687);
nor I_77961 (I1328939,I1328775,I1328922);
nor I_77962 (I1328664,I1328741,I1328939);
not I_77963 (I1328970,I1328922);
nand I_77964 (I1328667,I1328970,I1328724);
nand I_77965 (I1328661,I1328970,I1328792);
nor I_77966 (I1328658,I1328922,I1328905);
nor I_77967 (I1329029,I891690,I891693);
not I_77968 (I1329046,I1329029);
DFFARX1 I_77969 (I1329029,I3563,I1328690,I1329072,);
not I_77970 (I1328682,I1329072);
nor I_77971 (I1329094,I891690,I891705);
DFFARX1 I_77972 (I1329094,I3563,I1328690,I1329120,);
and I_77973 (I1329128,I1329120,I891702);
nor I_77974 (I1329145,I1329128,I1329046);
DFFARX1 I_77975 (I1329145,I3563,I1328690,I1328673,);
nor I_77976 (I1329176,I1329120,I1328905);
DFFARX1 I_77977 (I1329176,I3563,I1328690,I1328655,);
nor I_77978 (I1328670,I1329120,I1328809);
not I_77979 (I1329251,I3570);
DFFARX1 I_77980 (I1155156,I3563,I1329251,I1329277,);
nand I_77981 (I1329285,I1329277,I1155153);
not I_77982 (I1329302,I1329285);
DFFARX1 I_77983 (I1155156,I3563,I1329251,I1329328,);
not I_77984 (I1329336,I1329328);
nor I_77985 (I1329353,I1155174,I1155168);
not I_77986 (I1329370,I1329353);
DFFARX1 I_77987 (I1329370,I3563,I1329251,I1329237,);
or I_77988 (I1329401,I1155177,I1155174);
DFFARX1 I_77989 (I1329401,I3563,I1329251,I1329240,);
not I_77990 (I1329432,I1155165);
nor I_77991 (I1329449,I1329432,I1155162);
nor I_77992 (I1329466,I1329449,I1155168);
nor I_77993 (I1329483,I1155162,I1155153);
nor I_77994 (I1329500,I1329336,I1329483);
nor I_77995 (I1329225,I1329302,I1329500);
not I_77996 (I1329531,I1329483);
nand I_77997 (I1329228,I1329531,I1329285);
nand I_77998 (I1329222,I1329531,I1329353);
nor I_77999 (I1329219,I1329483,I1329466);
nor I_78000 (I1329590,I1155159,I1155177);
not I_78001 (I1329607,I1329590);
DFFARX1 I_78002 (I1329590,I3563,I1329251,I1329633,);
not I_78003 (I1329243,I1329633);
nor I_78004 (I1329655,I1155159,I1155171);
DFFARX1 I_78005 (I1329655,I3563,I1329251,I1329681,);
and I_78006 (I1329689,I1329681,I1155174);
nor I_78007 (I1329706,I1329689,I1329607);
DFFARX1 I_78008 (I1329706,I3563,I1329251,I1329234,);
nor I_78009 (I1329737,I1329681,I1329466);
DFFARX1 I_78010 (I1329737,I3563,I1329251,I1329216,);
nor I_78011 (I1329231,I1329681,I1329370);
not I_78012 (I1329812,I3570);
DFFARX1 I_78013 (I534053,I3563,I1329812,I1329838,);
nand I_78014 (I1329846,I1329838,I534044);
not I_78015 (I1329863,I1329846);
DFFARX1 I_78016 (I534044,I3563,I1329812,I1329889,);
not I_78017 (I1329897,I1329889);
nor I_78018 (I1329914,I534041,I534062);
not I_78019 (I1329931,I1329914);
DFFARX1 I_78020 (I1329931,I3563,I1329812,I1329798,);
or I_78021 (I1329962,I534056,I534041);
DFFARX1 I_78022 (I1329962,I3563,I1329812,I1329801,);
not I_78023 (I1329993,I534047);
nor I_78024 (I1330010,I1329993,I534041);
nor I_78025 (I1330027,I1330010,I534062);
nor I_78026 (I1330044,I534041,I534050);
nor I_78027 (I1330061,I1329897,I1330044);
nor I_78028 (I1329786,I1329863,I1330061);
not I_78029 (I1330092,I1330044);
nand I_78030 (I1329789,I1330092,I1329846);
nand I_78031 (I1329783,I1330092,I1329914);
nor I_78032 (I1329780,I1330044,I1330027);
nor I_78033 (I1330151,I534065,I534056);
not I_78034 (I1330168,I1330151);
DFFARX1 I_78035 (I1330151,I3563,I1329812,I1330194,);
not I_78036 (I1329804,I1330194);
nor I_78037 (I1330216,I534065,I534059);
DFFARX1 I_78038 (I1330216,I3563,I1329812,I1330242,);
and I_78039 (I1330250,I1330242,I534041);
nor I_78040 (I1330267,I1330250,I1330168);
DFFARX1 I_78041 (I1330267,I3563,I1329812,I1329795,);
nor I_78042 (I1330298,I1330242,I1330027);
DFFARX1 I_78043 (I1330298,I3563,I1329812,I1329777,);
nor I_78044 (I1329792,I1330242,I1329931);
not I_78045 (I1330373,I3570);
DFFARX1 I_78046 (I1029223,I3563,I1330373,I1330399,);
DFFARX1 I_78047 (I1029241,I3563,I1330373,I1330416,);
not I_78048 (I1330424,I1330416);
nor I_78049 (I1330341,I1330399,I1330424);
DFFARX1 I_78050 (I1330424,I3563,I1330373,I1330356,);
nor I_78051 (I1330469,I1029220,I1029232);
and I_78052 (I1330486,I1330469,I1029217);
nor I_78053 (I1330503,I1330486,I1029220);
not I_78054 (I1330520,I1029220);
and I_78055 (I1330537,I1330520,I1029226);
nand I_78056 (I1330554,I1330537,I1029238);
nor I_78057 (I1330571,I1330520,I1330554);
DFFARX1 I_78058 (I1330571,I3563,I1330373,I1330338,);
not I_78059 (I1330602,I1330554);
nand I_78060 (I1330619,I1330424,I1330602);
nand I_78061 (I1330350,I1330486,I1330602);
DFFARX1 I_78062 (I1330520,I3563,I1330373,I1330365,);
not I_78063 (I1330664,I1029229);
nor I_78064 (I1330681,I1330664,I1029226);
nor I_78065 (I1330698,I1330681,I1330503);
DFFARX1 I_78066 (I1330698,I3563,I1330373,I1330362,);
not I_78067 (I1330729,I1330681);
DFFARX1 I_78068 (I1330729,I3563,I1330373,I1330755,);
not I_78069 (I1330763,I1330755);
nor I_78070 (I1330359,I1330763,I1330681);
nor I_78071 (I1330794,I1330664,I1029217);
and I_78072 (I1330811,I1330794,I1029244);
or I_78073 (I1330828,I1330811,I1029235);
DFFARX1 I_78074 (I1330828,I3563,I1330373,I1330854,);
not I_78075 (I1330862,I1330854);
nand I_78076 (I1330879,I1330862,I1330602);
not I_78077 (I1330353,I1330879);
nand I_78078 (I1330347,I1330879,I1330619);
nand I_78079 (I1330344,I1330862,I1330486);
not I_78080 (I1330968,I3570);
DFFARX1 I_78081 (I289075,I3563,I1330968,I1330994,);
DFFARX1 I_78082 (I289069,I3563,I1330968,I1331011,);
not I_78083 (I1331019,I1331011);
nor I_78084 (I1330936,I1330994,I1331019);
DFFARX1 I_78085 (I1331019,I3563,I1330968,I1330951,);
nor I_78086 (I1331064,I289057,I289078);
and I_78087 (I1331081,I1331064,I289072);
nor I_78088 (I1331098,I1331081,I289057);
not I_78089 (I1331115,I289057);
and I_78090 (I1331132,I1331115,I289054);
nand I_78091 (I1331149,I1331132,I289066);
nor I_78092 (I1331166,I1331115,I1331149);
DFFARX1 I_78093 (I1331166,I3563,I1330968,I1330933,);
not I_78094 (I1331197,I1331149);
nand I_78095 (I1331214,I1331019,I1331197);
nand I_78096 (I1330945,I1331081,I1331197);
DFFARX1 I_78097 (I1331115,I3563,I1330968,I1330960,);
not I_78098 (I1331259,I289081);
nor I_78099 (I1331276,I1331259,I289054);
nor I_78100 (I1331293,I1331276,I1331098);
DFFARX1 I_78101 (I1331293,I3563,I1330968,I1330957,);
not I_78102 (I1331324,I1331276);
DFFARX1 I_78103 (I1331324,I3563,I1330968,I1331350,);
not I_78104 (I1331358,I1331350);
nor I_78105 (I1330954,I1331358,I1331276);
nor I_78106 (I1331389,I1331259,I289063);
and I_78107 (I1331406,I1331389,I289060);
or I_78108 (I1331423,I1331406,I289054);
DFFARX1 I_78109 (I1331423,I3563,I1330968,I1331449,);
not I_78110 (I1331457,I1331449);
nand I_78111 (I1331474,I1331457,I1331197);
not I_78112 (I1330948,I1331474);
nand I_78113 (I1330942,I1331474,I1331214);
nand I_78114 (I1330939,I1331457,I1331081);
not I_78115 (I1331563,I3570);
DFFARX1 I_78116 (I726060,I3563,I1331563,I1331589,);
DFFARX1 I_78117 (I726042,I3563,I1331563,I1331606,);
not I_78118 (I1331614,I1331606);
nor I_78119 (I1331531,I1331589,I1331614);
DFFARX1 I_78120 (I1331614,I3563,I1331563,I1331546,);
nor I_78121 (I1331659,I726048,I726051);
and I_78122 (I1331676,I1331659,I726039);
nor I_78123 (I1331693,I1331676,I726048);
not I_78124 (I1331710,I726048);
and I_78125 (I1331727,I1331710,I726057);
nand I_78126 (I1331744,I1331727,I726045);
nor I_78127 (I1331761,I1331710,I1331744);
DFFARX1 I_78128 (I1331761,I3563,I1331563,I1331528,);
not I_78129 (I1331792,I1331744);
nand I_78130 (I1331809,I1331614,I1331792);
nand I_78131 (I1331540,I1331676,I1331792);
DFFARX1 I_78132 (I1331710,I3563,I1331563,I1331555,);
not I_78133 (I1331854,I726042);
nor I_78134 (I1331871,I1331854,I726057);
nor I_78135 (I1331888,I1331871,I1331693);
DFFARX1 I_78136 (I1331888,I3563,I1331563,I1331552,);
not I_78137 (I1331919,I1331871);
DFFARX1 I_78138 (I1331919,I3563,I1331563,I1331945,);
not I_78139 (I1331953,I1331945);
nor I_78140 (I1331549,I1331953,I1331871);
nor I_78141 (I1331984,I1331854,I726054);
and I_78142 (I1332001,I1331984,I726063);
or I_78143 (I1332018,I1332001,I726039);
DFFARX1 I_78144 (I1332018,I3563,I1331563,I1332044,);
not I_78145 (I1332052,I1332044);
nand I_78146 (I1332069,I1332052,I1331792);
not I_78147 (I1331543,I1332069);
nand I_78148 (I1331537,I1332069,I1331809);
nand I_78149 (I1331534,I1332052,I1331676);
not I_78150 (I1332158,I3570);
DFFARX1 I_78151 (I347045,I3563,I1332158,I1332184,);
DFFARX1 I_78152 (I347039,I3563,I1332158,I1332201,);
not I_78153 (I1332209,I1332201);
nor I_78154 (I1332126,I1332184,I1332209);
DFFARX1 I_78155 (I1332209,I3563,I1332158,I1332141,);
nor I_78156 (I1332254,I347027,I347048);
and I_78157 (I1332271,I1332254,I347042);
nor I_78158 (I1332288,I1332271,I347027);
not I_78159 (I1332305,I347027);
and I_78160 (I1332322,I1332305,I347024);
nand I_78161 (I1332339,I1332322,I347036);
nor I_78162 (I1332356,I1332305,I1332339);
DFFARX1 I_78163 (I1332356,I3563,I1332158,I1332123,);
not I_78164 (I1332387,I1332339);
nand I_78165 (I1332404,I1332209,I1332387);
nand I_78166 (I1332135,I1332271,I1332387);
DFFARX1 I_78167 (I1332305,I3563,I1332158,I1332150,);
not I_78168 (I1332449,I347051);
nor I_78169 (I1332466,I1332449,I347024);
nor I_78170 (I1332483,I1332466,I1332288);
DFFARX1 I_78171 (I1332483,I3563,I1332158,I1332147,);
not I_78172 (I1332514,I1332466);
DFFARX1 I_78173 (I1332514,I3563,I1332158,I1332540,);
not I_78174 (I1332548,I1332540);
nor I_78175 (I1332144,I1332548,I1332466);
nor I_78176 (I1332579,I1332449,I347033);
and I_78177 (I1332596,I1332579,I347030);
or I_78178 (I1332613,I1332596,I347024);
DFFARX1 I_78179 (I1332613,I3563,I1332158,I1332639,);
not I_78180 (I1332647,I1332639);
nand I_78181 (I1332664,I1332647,I1332387);
not I_78182 (I1332138,I1332664);
nand I_78183 (I1332132,I1332664,I1332404);
nand I_78184 (I1332129,I1332647,I1332271);
not I_78185 (I1332753,I3570);
DFFARX1 I_78186 (I1020825,I3563,I1332753,I1332779,);
DFFARX1 I_78187 (I1020843,I3563,I1332753,I1332796,);
not I_78188 (I1332804,I1332796);
nor I_78189 (I1332721,I1332779,I1332804);
DFFARX1 I_78190 (I1332804,I3563,I1332753,I1332736,);
nor I_78191 (I1332849,I1020822,I1020834);
and I_78192 (I1332866,I1332849,I1020819);
nor I_78193 (I1332883,I1332866,I1020822);
not I_78194 (I1332900,I1020822);
and I_78195 (I1332917,I1332900,I1020828);
nand I_78196 (I1332934,I1332917,I1020840);
nor I_78197 (I1332951,I1332900,I1332934);
DFFARX1 I_78198 (I1332951,I3563,I1332753,I1332718,);
not I_78199 (I1332982,I1332934);
nand I_78200 (I1332999,I1332804,I1332982);
nand I_78201 (I1332730,I1332866,I1332982);
DFFARX1 I_78202 (I1332900,I3563,I1332753,I1332745,);
not I_78203 (I1333044,I1020831);
nor I_78204 (I1333061,I1333044,I1020828);
nor I_78205 (I1333078,I1333061,I1332883);
DFFARX1 I_78206 (I1333078,I3563,I1332753,I1332742,);
not I_78207 (I1333109,I1333061);
DFFARX1 I_78208 (I1333109,I3563,I1332753,I1333135,);
not I_78209 (I1333143,I1333135);
nor I_78210 (I1332739,I1333143,I1333061);
nor I_78211 (I1333174,I1333044,I1020819);
and I_78212 (I1333191,I1333174,I1020846);
or I_78213 (I1333208,I1333191,I1020837);
DFFARX1 I_78214 (I1333208,I3563,I1332753,I1333234,);
not I_78215 (I1333242,I1333234);
nand I_78216 (I1333259,I1333242,I1332982);
not I_78217 (I1332733,I1333259);
nand I_78218 (I1332727,I1333259,I1332999);
nand I_78219 (I1332724,I1333242,I1332866);
not I_78220 (I1333348,I3570);
DFFARX1 I_78221 (I978189,I3563,I1333348,I1333374,);
DFFARX1 I_78222 (I978207,I3563,I1333348,I1333391,);
not I_78223 (I1333399,I1333391);
nor I_78224 (I1333316,I1333374,I1333399);
DFFARX1 I_78225 (I1333399,I3563,I1333348,I1333331,);
nor I_78226 (I1333444,I978186,I978198);
and I_78227 (I1333461,I1333444,I978183);
nor I_78228 (I1333478,I1333461,I978186);
not I_78229 (I1333495,I978186);
and I_78230 (I1333512,I1333495,I978192);
nand I_78231 (I1333529,I1333512,I978204);
nor I_78232 (I1333546,I1333495,I1333529);
DFFARX1 I_78233 (I1333546,I3563,I1333348,I1333313,);
not I_78234 (I1333577,I1333529);
nand I_78235 (I1333594,I1333399,I1333577);
nand I_78236 (I1333325,I1333461,I1333577);
DFFARX1 I_78237 (I1333495,I3563,I1333348,I1333340,);
not I_78238 (I1333639,I978195);
nor I_78239 (I1333656,I1333639,I978192);
nor I_78240 (I1333673,I1333656,I1333478);
DFFARX1 I_78241 (I1333673,I3563,I1333348,I1333337,);
not I_78242 (I1333704,I1333656);
DFFARX1 I_78243 (I1333704,I3563,I1333348,I1333730,);
not I_78244 (I1333738,I1333730);
nor I_78245 (I1333334,I1333738,I1333656);
nor I_78246 (I1333769,I1333639,I978183);
and I_78247 (I1333786,I1333769,I978210);
or I_78248 (I1333803,I1333786,I978201);
DFFARX1 I_78249 (I1333803,I3563,I1333348,I1333829,);
not I_78250 (I1333837,I1333829);
nand I_78251 (I1333854,I1333837,I1333577);
not I_78252 (I1333328,I1333854);
nand I_78253 (I1333322,I1333854,I1333594);
nand I_78254 (I1333319,I1333837,I1333461);
not I_78255 (I1333943,I3570);
DFFARX1 I_78256 (I398691,I3563,I1333943,I1333969,);
DFFARX1 I_78257 (I398685,I3563,I1333943,I1333986,);
not I_78258 (I1333994,I1333986);
nor I_78259 (I1333911,I1333969,I1333994);
DFFARX1 I_78260 (I1333994,I3563,I1333943,I1333926,);
nor I_78261 (I1334039,I398673,I398694);
and I_78262 (I1334056,I1334039,I398688);
nor I_78263 (I1334073,I1334056,I398673);
not I_78264 (I1334090,I398673);
and I_78265 (I1334107,I1334090,I398670);
nand I_78266 (I1334124,I1334107,I398682);
nor I_78267 (I1334141,I1334090,I1334124);
DFFARX1 I_78268 (I1334141,I3563,I1333943,I1333908,);
not I_78269 (I1334172,I1334124);
nand I_78270 (I1334189,I1333994,I1334172);
nand I_78271 (I1333920,I1334056,I1334172);
DFFARX1 I_78272 (I1334090,I3563,I1333943,I1333935,);
not I_78273 (I1334234,I398697);
nor I_78274 (I1334251,I1334234,I398670);
nor I_78275 (I1334268,I1334251,I1334073);
DFFARX1 I_78276 (I1334268,I3563,I1333943,I1333932,);
not I_78277 (I1334299,I1334251);
DFFARX1 I_78278 (I1334299,I3563,I1333943,I1334325,);
not I_78279 (I1334333,I1334325);
nor I_78280 (I1333929,I1334333,I1334251);
nor I_78281 (I1334364,I1334234,I398679);
and I_78282 (I1334381,I1334364,I398676);
or I_78283 (I1334398,I1334381,I398670);
DFFARX1 I_78284 (I1334398,I3563,I1333943,I1334424,);
not I_78285 (I1334432,I1334424);
nand I_78286 (I1334449,I1334432,I1334172);
not I_78287 (I1333923,I1334449);
nand I_78288 (I1333917,I1334449,I1334189);
nand I_78289 (I1333914,I1334432,I1334056);
not I_78290 (I1334538,I3570);
DFFARX1 I_78291 (I687334,I3563,I1334538,I1334564,);
DFFARX1 I_78292 (I687316,I3563,I1334538,I1334581,);
not I_78293 (I1334589,I1334581);
nor I_78294 (I1334506,I1334564,I1334589);
DFFARX1 I_78295 (I1334589,I3563,I1334538,I1334521,);
nor I_78296 (I1334634,I687322,I687325);
and I_78297 (I1334651,I1334634,I687313);
nor I_78298 (I1334668,I1334651,I687322);
not I_78299 (I1334685,I687322);
and I_78300 (I1334702,I1334685,I687331);
nand I_78301 (I1334719,I1334702,I687319);
nor I_78302 (I1334736,I1334685,I1334719);
DFFARX1 I_78303 (I1334736,I3563,I1334538,I1334503,);
not I_78304 (I1334767,I1334719);
nand I_78305 (I1334784,I1334589,I1334767);
nand I_78306 (I1334515,I1334651,I1334767);
DFFARX1 I_78307 (I1334685,I3563,I1334538,I1334530,);
not I_78308 (I1334829,I687316);
nor I_78309 (I1334846,I1334829,I687331);
nor I_78310 (I1334863,I1334846,I1334668);
DFFARX1 I_78311 (I1334863,I3563,I1334538,I1334527,);
not I_78312 (I1334894,I1334846);
DFFARX1 I_78313 (I1334894,I3563,I1334538,I1334920,);
not I_78314 (I1334928,I1334920);
nor I_78315 (I1334524,I1334928,I1334846);
nor I_78316 (I1334959,I1334829,I687328);
and I_78317 (I1334976,I1334959,I687337);
or I_78318 (I1334993,I1334976,I687313);
DFFARX1 I_78319 (I1334993,I3563,I1334538,I1335019,);
not I_78320 (I1335027,I1335019);
nand I_78321 (I1335044,I1335027,I1334767);
not I_78322 (I1334518,I1335044);
nand I_78323 (I1334512,I1335044,I1334784);
nand I_78324 (I1334509,I1335027,I1334651);
not I_78325 (I1335133,I3570);
DFFARX1 I_78326 (I1121632,I3563,I1335133,I1335159,);
DFFARX1 I_78327 (I1121644,I3563,I1335133,I1335176,);
not I_78328 (I1335184,I1335176);
nor I_78329 (I1335101,I1335159,I1335184);
DFFARX1 I_78330 (I1335184,I3563,I1335133,I1335116,);
nor I_78331 (I1335229,I1121641,I1121635);
and I_78332 (I1335246,I1335229,I1121629);
nor I_78333 (I1335263,I1335246,I1121641);
not I_78334 (I1335280,I1121641);
and I_78335 (I1335297,I1335280,I1121638);
nand I_78336 (I1335314,I1335297,I1121629);
nor I_78337 (I1335331,I1335280,I1335314);
DFFARX1 I_78338 (I1335331,I3563,I1335133,I1335098,);
not I_78339 (I1335362,I1335314);
nand I_78340 (I1335379,I1335184,I1335362);
nand I_78341 (I1335110,I1335246,I1335362);
DFFARX1 I_78342 (I1335280,I3563,I1335133,I1335125,);
not I_78343 (I1335424,I1121653);
nor I_78344 (I1335441,I1335424,I1121638);
nor I_78345 (I1335458,I1335441,I1335263);
DFFARX1 I_78346 (I1335458,I3563,I1335133,I1335122,);
not I_78347 (I1335489,I1335441);
DFFARX1 I_78348 (I1335489,I3563,I1335133,I1335515,);
not I_78349 (I1335523,I1335515);
nor I_78350 (I1335119,I1335523,I1335441);
nor I_78351 (I1335554,I1335424,I1121647);
and I_78352 (I1335571,I1335554,I1121650);
or I_78353 (I1335588,I1335571,I1121632);
DFFARX1 I_78354 (I1335588,I3563,I1335133,I1335614,);
not I_78355 (I1335622,I1335614);
nand I_78356 (I1335639,I1335622,I1335362);
not I_78357 (I1335113,I1335639);
nand I_78358 (I1335107,I1335639,I1335379);
nand I_78359 (I1335104,I1335622,I1335246);
not I_78360 (I1335728,I3570);
DFFARX1 I_78361 (I1196194,I3563,I1335728,I1335754,);
DFFARX1 I_78362 (I1196206,I3563,I1335728,I1335771,);
not I_78363 (I1335779,I1335771);
nor I_78364 (I1335696,I1335754,I1335779);
DFFARX1 I_78365 (I1335779,I3563,I1335728,I1335711,);
nor I_78366 (I1335824,I1196203,I1196197);
and I_78367 (I1335841,I1335824,I1196191);
nor I_78368 (I1335858,I1335841,I1196203);
not I_78369 (I1335875,I1196203);
and I_78370 (I1335892,I1335875,I1196200);
nand I_78371 (I1335909,I1335892,I1196191);
nor I_78372 (I1335926,I1335875,I1335909);
DFFARX1 I_78373 (I1335926,I3563,I1335728,I1335693,);
not I_78374 (I1335957,I1335909);
nand I_78375 (I1335974,I1335779,I1335957);
nand I_78376 (I1335705,I1335841,I1335957);
DFFARX1 I_78377 (I1335875,I3563,I1335728,I1335720,);
not I_78378 (I1336019,I1196215);
nor I_78379 (I1336036,I1336019,I1196200);
nor I_78380 (I1336053,I1336036,I1335858);
DFFARX1 I_78381 (I1336053,I3563,I1335728,I1335717,);
not I_78382 (I1336084,I1336036);
DFFARX1 I_78383 (I1336084,I3563,I1335728,I1336110,);
not I_78384 (I1336118,I1336110);
nor I_78385 (I1335714,I1336118,I1336036);
nor I_78386 (I1336149,I1336019,I1196209);
and I_78387 (I1336166,I1336149,I1196212);
or I_78388 (I1336183,I1336166,I1196194);
DFFARX1 I_78389 (I1336183,I3563,I1335728,I1336209,);
not I_78390 (I1336217,I1336209);
nand I_78391 (I1336234,I1336217,I1335957);
not I_78392 (I1335708,I1336234);
nand I_78393 (I1335702,I1336234,I1335974);
nand I_78394 (I1335699,I1336217,I1335841);
not I_78395 (I1336323,I3570);
DFFARX1 I_78396 (I1099668,I3563,I1336323,I1336349,);
DFFARX1 I_78397 (I1099680,I3563,I1336323,I1336366,);
not I_78398 (I1336374,I1336366);
nor I_78399 (I1336291,I1336349,I1336374);
DFFARX1 I_78400 (I1336374,I3563,I1336323,I1336306,);
nor I_78401 (I1336419,I1099677,I1099671);
and I_78402 (I1336436,I1336419,I1099665);
nor I_78403 (I1336453,I1336436,I1099677);
not I_78404 (I1336470,I1099677);
and I_78405 (I1336487,I1336470,I1099674);
nand I_78406 (I1336504,I1336487,I1099665);
nor I_78407 (I1336521,I1336470,I1336504);
DFFARX1 I_78408 (I1336521,I3563,I1336323,I1336288,);
not I_78409 (I1336552,I1336504);
nand I_78410 (I1336569,I1336374,I1336552);
nand I_78411 (I1336300,I1336436,I1336552);
DFFARX1 I_78412 (I1336470,I3563,I1336323,I1336315,);
not I_78413 (I1336614,I1099689);
nor I_78414 (I1336631,I1336614,I1099674);
nor I_78415 (I1336648,I1336631,I1336453);
DFFARX1 I_78416 (I1336648,I3563,I1336323,I1336312,);
not I_78417 (I1336679,I1336631);
DFFARX1 I_78418 (I1336679,I3563,I1336323,I1336705,);
not I_78419 (I1336713,I1336705);
nor I_78420 (I1336309,I1336713,I1336631);
nor I_78421 (I1336744,I1336614,I1099683);
and I_78422 (I1336761,I1336744,I1099686);
or I_78423 (I1336778,I1336761,I1099668);
DFFARX1 I_78424 (I1336778,I3563,I1336323,I1336804,);
not I_78425 (I1336812,I1336804);
nand I_78426 (I1336829,I1336812,I1336552);
not I_78427 (I1336303,I1336829);
nand I_78428 (I1336297,I1336829,I1336569);
nand I_78429 (I1336294,I1336812,I1336436);
not I_78430 (I1336918,I3570);
DFFARX1 I_78431 (I701784,I3563,I1336918,I1336944,);
DFFARX1 I_78432 (I701766,I3563,I1336918,I1336961,);
not I_78433 (I1336969,I1336961);
nor I_78434 (I1336886,I1336944,I1336969);
DFFARX1 I_78435 (I1336969,I3563,I1336918,I1336901,);
nor I_78436 (I1337014,I701772,I701775);
and I_78437 (I1337031,I1337014,I701763);
nor I_78438 (I1337048,I1337031,I701772);
not I_78439 (I1337065,I701772);
and I_78440 (I1337082,I1337065,I701781);
nand I_78441 (I1337099,I1337082,I701769);
nor I_78442 (I1337116,I1337065,I1337099);
DFFARX1 I_78443 (I1337116,I3563,I1336918,I1336883,);
not I_78444 (I1337147,I1337099);
nand I_78445 (I1337164,I1336969,I1337147);
nand I_78446 (I1336895,I1337031,I1337147);
DFFARX1 I_78447 (I1337065,I3563,I1336918,I1336910,);
not I_78448 (I1337209,I701766);
nor I_78449 (I1337226,I1337209,I701781);
nor I_78450 (I1337243,I1337226,I1337048);
DFFARX1 I_78451 (I1337243,I3563,I1336918,I1336907,);
not I_78452 (I1337274,I1337226);
DFFARX1 I_78453 (I1337274,I3563,I1336918,I1337300,);
not I_78454 (I1337308,I1337300);
nor I_78455 (I1336904,I1337308,I1337226);
nor I_78456 (I1337339,I1337209,I701778);
and I_78457 (I1337356,I1337339,I701787);
or I_78458 (I1337373,I1337356,I701763);
DFFARX1 I_78459 (I1337373,I3563,I1336918,I1337399,);
not I_78460 (I1337407,I1337399);
nand I_78461 (I1337424,I1337407,I1337147);
not I_78462 (I1336898,I1337424);
nand I_78463 (I1336892,I1337424,I1337164);
nand I_78464 (I1336889,I1337407,I1337031);
not I_78465 (I1337513,I3570);
DFFARX1 I_78466 (I172638,I3563,I1337513,I1337539,);
DFFARX1 I_78467 (I172641,I3563,I1337513,I1337556,);
not I_78468 (I1337564,I1337556);
nor I_78469 (I1337481,I1337539,I1337564);
DFFARX1 I_78470 (I1337564,I3563,I1337513,I1337496,);
nor I_78471 (I1337609,I172647,I172641);
and I_78472 (I1337626,I1337609,I172644);
nor I_78473 (I1337643,I1337626,I172647);
not I_78474 (I1337660,I172647);
and I_78475 (I1337677,I1337660,I172638);
nand I_78476 (I1337694,I1337677,I172656);
nor I_78477 (I1337711,I1337660,I1337694);
DFFARX1 I_78478 (I1337711,I3563,I1337513,I1337478,);
not I_78479 (I1337742,I1337694);
nand I_78480 (I1337759,I1337564,I1337742);
nand I_78481 (I1337490,I1337626,I1337742);
DFFARX1 I_78482 (I1337660,I3563,I1337513,I1337505,);
not I_78483 (I1337804,I172650);
nor I_78484 (I1337821,I1337804,I172638);
nor I_78485 (I1337838,I1337821,I1337643);
DFFARX1 I_78486 (I1337838,I3563,I1337513,I1337502,);
not I_78487 (I1337869,I1337821);
DFFARX1 I_78488 (I1337869,I3563,I1337513,I1337895,);
not I_78489 (I1337903,I1337895);
nor I_78490 (I1337499,I1337903,I1337821);
nor I_78491 (I1337934,I1337804,I172653);
and I_78492 (I1337951,I1337934,I172659);
or I_78493 (I1337968,I1337951,I172662);
DFFARX1 I_78494 (I1337968,I3563,I1337513,I1337994,);
not I_78495 (I1338002,I1337994);
nand I_78496 (I1338019,I1338002,I1337742);
not I_78497 (I1337493,I1338019);
nand I_78498 (I1337487,I1338019,I1337759);
nand I_78499 (I1337484,I1338002,I1337626);
not I_78500 (I1338108,I3570);
DFFARX1 I_78501 (I1156890,I3563,I1338108,I1338134,);
DFFARX1 I_78502 (I1156902,I3563,I1338108,I1338151,);
not I_78503 (I1338159,I1338151);
nor I_78504 (I1338076,I1338134,I1338159);
DFFARX1 I_78505 (I1338159,I3563,I1338108,I1338091,);
nor I_78506 (I1338204,I1156899,I1156893);
and I_78507 (I1338221,I1338204,I1156887);
nor I_78508 (I1338238,I1338221,I1156899);
not I_78509 (I1338255,I1156899);
and I_78510 (I1338272,I1338255,I1156896);
nand I_78511 (I1338289,I1338272,I1156887);
nor I_78512 (I1338306,I1338255,I1338289);
DFFARX1 I_78513 (I1338306,I3563,I1338108,I1338073,);
not I_78514 (I1338337,I1338289);
nand I_78515 (I1338354,I1338159,I1338337);
nand I_78516 (I1338085,I1338221,I1338337);
DFFARX1 I_78517 (I1338255,I3563,I1338108,I1338100,);
not I_78518 (I1338399,I1156911);
nor I_78519 (I1338416,I1338399,I1156896);
nor I_78520 (I1338433,I1338416,I1338238);
DFFARX1 I_78521 (I1338433,I3563,I1338108,I1338097,);
not I_78522 (I1338464,I1338416);
DFFARX1 I_78523 (I1338464,I3563,I1338108,I1338490,);
not I_78524 (I1338498,I1338490);
nor I_78525 (I1338094,I1338498,I1338416);
nor I_78526 (I1338529,I1338399,I1156905);
and I_78527 (I1338546,I1338529,I1156908);
or I_78528 (I1338563,I1338546,I1156890);
DFFARX1 I_78529 (I1338563,I3563,I1338108,I1338589,);
not I_78530 (I1338597,I1338589);
nand I_78531 (I1338614,I1338597,I1338337);
not I_78532 (I1338088,I1338614);
nand I_78533 (I1338082,I1338614,I1338354);
nand I_78534 (I1338079,I1338597,I1338221);
not I_78535 (I1338703,I3570);
DFFARX1 I_78536 (I528091,I3563,I1338703,I1338729,);
DFFARX1 I_78537 (I528094,I3563,I1338703,I1338746,);
not I_78538 (I1338754,I1338746);
nor I_78539 (I1338671,I1338729,I1338754);
DFFARX1 I_78540 (I1338754,I3563,I1338703,I1338686,);
nor I_78541 (I1338799,I528097,I528115);
and I_78542 (I1338816,I1338799,I528100);
nor I_78543 (I1338833,I1338816,I528097);
not I_78544 (I1338850,I528097);
and I_78545 (I1338867,I1338850,I528109);
nand I_78546 (I1338884,I1338867,I528112);
nor I_78547 (I1338901,I1338850,I1338884);
DFFARX1 I_78548 (I1338901,I3563,I1338703,I1338668,);
not I_78549 (I1338932,I1338884);
nand I_78550 (I1338949,I1338754,I1338932);
nand I_78551 (I1338680,I1338816,I1338932);
DFFARX1 I_78552 (I1338850,I3563,I1338703,I1338695,);
not I_78553 (I1338994,I528103);
nor I_78554 (I1339011,I1338994,I528109);
nor I_78555 (I1339028,I1339011,I1338833);
DFFARX1 I_78556 (I1339028,I3563,I1338703,I1338692,);
not I_78557 (I1339059,I1339011);
DFFARX1 I_78558 (I1339059,I3563,I1338703,I1339085,);
not I_78559 (I1339093,I1339085);
nor I_78560 (I1338689,I1339093,I1339011);
nor I_78561 (I1339124,I1338994,I528091);
and I_78562 (I1339141,I1339124,I528106);
or I_78563 (I1339158,I1339141,I528094);
DFFARX1 I_78564 (I1339158,I3563,I1338703,I1339184,);
not I_78565 (I1339192,I1339184);
nand I_78566 (I1339209,I1339192,I1338932);
not I_78567 (I1338683,I1339209);
nand I_78568 (I1338677,I1339209,I1338949);
nand I_78569 (I1338674,I1339192,I1338816);
not I_78570 (I1339298,I3570);
DFFARX1 I_78571 (I187513,I3563,I1339298,I1339324,);
DFFARX1 I_78572 (I187516,I3563,I1339298,I1339341,);
not I_78573 (I1339349,I1339341);
nor I_78574 (I1339266,I1339324,I1339349);
DFFARX1 I_78575 (I1339349,I3563,I1339298,I1339281,);
nor I_78576 (I1339394,I187522,I187516);
and I_78577 (I1339411,I1339394,I187519);
nor I_78578 (I1339428,I1339411,I187522);
not I_78579 (I1339445,I187522);
and I_78580 (I1339462,I1339445,I187513);
nand I_78581 (I1339479,I1339462,I187531);
nor I_78582 (I1339496,I1339445,I1339479);
DFFARX1 I_78583 (I1339496,I3563,I1339298,I1339263,);
not I_78584 (I1339527,I1339479);
nand I_78585 (I1339544,I1339349,I1339527);
nand I_78586 (I1339275,I1339411,I1339527);
DFFARX1 I_78587 (I1339445,I3563,I1339298,I1339290,);
not I_78588 (I1339589,I187525);
nor I_78589 (I1339606,I1339589,I187513);
nor I_78590 (I1339623,I1339606,I1339428);
DFFARX1 I_78591 (I1339623,I3563,I1339298,I1339287,);
not I_78592 (I1339654,I1339606);
DFFARX1 I_78593 (I1339654,I3563,I1339298,I1339680,);
not I_78594 (I1339688,I1339680);
nor I_78595 (I1339284,I1339688,I1339606);
nor I_78596 (I1339719,I1339589,I187528);
and I_78597 (I1339736,I1339719,I187534);
or I_78598 (I1339753,I1339736,I187537);
DFFARX1 I_78599 (I1339753,I3563,I1339298,I1339779,);
not I_78600 (I1339787,I1339779);
nand I_78601 (I1339804,I1339787,I1339527);
not I_78602 (I1339278,I1339804);
nand I_78603 (I1339272,I1339804,I1339544);
nand I_78604 (I1339269,I1339787,I1339411);
not I_78605 (I1339893,I3570);
DFFARX1 I_78606 (I275573,I3563,I1339893,I1339919,);
DFFARX1 I_78607 (I275576,I3563,I1339893,I1339936,);
not I_78608 (I1339944,I1339936);
nor I_78609 (I1339861,I1339919,I1339944);
DFFARX1 I_78610 (I1339944,I3563,I1339893,I1339876,);
nor I_78611 (I1339989,I275582,I275576);
and I_78612 (I1340006,I1339989,I275579);
nor I_78613 (I1340023,I1340006,I275582);
not I_78614 (I1340040,I275582);
and I_78615 (I1340057,I1340040,I275573);
nand I_78616 (I1340074,I1340057,I275591);
nor I_78617 (I1340091,I1340040,I1340074);
DFFARX1 I_78618 (I1340091,I3563,I1339893,I1339858,);
not I_78619 (I1340122,I1340074);
nand I_78620 (I1340139,I1339944,I1340122);
nand I_78621 (I1339870,I1340006,I1340122);
DFFARX1 I_78622 (I1340040,I3563,I1339893,I1339885,);
not I_78623 (I1340184,I275585);
nor I_78624 (I1340201,I1340184,I275573);
nor I_78625 (I1340218,I1340201,I1340023);
DFFARX1 I_78626 (I1340218,I3563,I1339893,I1339882,);
not I_78627 (I1340249,I1340201);
DFFARX1 I_78628 (I1340249,I3563,I1339893,I1340275,);
not I_78629 (I1340283,I1340275);
nor I_78630 (I1339879,I1340283,I1340201);
nor I_78631 (I1340314,I1340184,I275588);
and I_78632 (I1340331,I1340314,I275594);
or I_78633 (I1340348,I1340331,I275597);
DFFARX1 I_78634 (I1340348,I3563,I1339893,I1340374,);
not I_78635 (I1340382,I1340374);
nand I_78636 (I1340399,I1340382,I1340122);
not I_78637 (I1339873,I1340399);
nand I_78638 (I1339867,I1340399,I1340139);
nand I_78639 (I1339864,I1340382,I1340006);
not I_78640 (I1340488,I3570);
DFFARX1 I_78641 (I1257289,I3563,I1340488,I1340514,);
DFFARX1 I_78642 (I1257292,I3563,I1340488,I1340531,);
not I_78643 (I1340539,I1340531);
nor I_78644 (I1340456,I1340514,I1340539);
DFFARX1 I_78645 (I1340539,I3563,I1340488,I1340471,);
nor I_78646 (I1340584,I1257292,I1257307);
and I_78647 (I1340601,I1340584,I1257301);
nor I_78648 (I1340618,I1340601,I1257292);
not I_78649 (I1340635,I1257292);
and I_78650 (I1340652,I1340635,I1257310);
nand I_78651 (I1340669,I1340652,I1257298);
nor I_78652 (I1340686,I1340635,I1340669);
DFFARX1 I_78653 (I1340686,I3563,I1340488,I1340453,);
not I_78654 (I1340717,I1340669);
nand I_78655 (I1340734,I1340539,I1340717);
nand I_78656 (I1340465,I1340601,I1340717);
DFFARX1 I_78657 (I1340635,I3563,I1340488,I1340480,);
not I_78658 (I1340779,I1257304);
nor I_78659 (I1340796,I1340779,I1257310);
nor I_78660 (I1340813,I1340796,I1340618);
DFFARX1 I_78661 (I1340813,I3563,I1340488,I1340477,);
not I_78662 (I1340844,I1340796);
DFFARX1 I_78663 (I1340844,I3563,I1340488,I1340870,);
not I_78664 (I1340878,I1340870);
nor I_78665 (I1340474,I1340878,I1340796);
nor I_78666 (I1340909,I1340779,I1257289);
and I_78667 (I1340926,I1340909,I1257313);
or I_78668 (I1340943,I1340926,I1257295);
DFFARX1 I_78669 (I1340943,I3563,I1340488,I1340969,);
not I_78670 (I1340977,I1340969);
nand I_78671 (I1340994,I1340977,I1340717);
not I_78672 (I1340468,I1340994);
nand I_78673 (I1340462,I1340994,I1340734);
nand I_78674 (I1340459,I1340977,I1340601);
not I_78675 (I1341083,I3570);
DFFARX1 I_78676 (I517058,I3563,I1341083,I1341109,);
DFFARX1 I_78677 (I517064,I3563,I1341083,I1341126,);
not I_78678 (I1341134,I1341126);
nor I_78679 (I1341051,I1341109,I1341134);
DFFARX1 I_78680 (I1341134,I3563,I1341083,I1341066,);
nor I_78681 (I1341179,I517073,I517058);
and I_78682 (I1341196,I1341179,I517085);
nor I_78683 (I1341213,I1341196,I517073);
not I_78684 (I1341230,I517073);
and I_78685 (I1341247,I1341230,I517061);
nand I_78686 (I1341264,I1341247,I517082);
nor I_78687 (I1341281,I1341230,I1341264);
DFFARX1 I_78688 (I1341281,I3563,I1341083,I1341048,);
not I_78689 (I1341312,I1341264);
nand I_78690 (I1341329,I1341134,I1341312);
nand I_78691 (I1341060,I1341196,I1341312);
DFFARX1 I_78692 (I1341230,I3563,I1341083,I1341075,);
not I_78693 (I1341374,I517070);
nor I_78694 (I1341391,I1341374,I517061);
nor I_78695 (I1341408,I1341391,I1341213);
DFFARX1 I_78696 (I1341408,I3563,I1341083,I1341072,);
not I_78697 (I1341439,I1341391);
DFFARX1 I_78698 (I1341439,I3563,I1341083,I1341465,);
not I_78699 (I1341473,I1341465);
nor I_78700 (I1341069,I1341473,I1341391);
nor I_78701 (I1341504,I1341374,I517067);
and I_78702 (I1341521,I1341504,I517079);
or I_78703 (I1341538,I1341521,I517076);
DFFARX1 I_78704 (I1341538,I3563,I1341083,I1341564,);
not I_78705 (I1341572,I1341564);
nand I_78706 (I1341589,I1341572,I1341312);
not I_78707 (I1341063,I1341589);
nand I_78708 (I1341057,I1341589,I1341329);
nand I_78709 (I1341054,I1341572,I1341196);
not I_78710 (I1341678,I3570);
DFFARX1 I_78711 (I1283401,I3563,I1341678,I1341704,);
DFFARX1 I_78712 (I1283404,I3563,I1341678,I1341721,);
not I_78713 (I1341729,I1341721);
nor I_78714 (I1341646,I1341704,I1341729);
DFFARX1 I_78715 (I1341729,I3563,I1341678,I1341661,);
nor I_78716 (I1341774,I1283404,I1283419);
and I_78717 (I1341791,I1341774,I1283413);
nor I_78718 (I1341808,I1341791,I1283404);
not I_78719 (I1341825,I1283404);
and I_78720 (I1341842,I1341825,I1283422);
nand I_78721 (I1341859,I1341842,I1283410);
nor I_78722 (I1341876,I1341825,I1341859);
DFFARX1 I_78723 (I1341876,I3563,I1341678,I1341643,);
not I_78724 (I1341907,I1341859);
nand I_78725 (I1341924,I1341729,I1341907);
nand I_78726 (I1341655,I1341791,I1341907);
DFFARX1 I_78727 (I1341825,I3563,I1341678,I1341670,);
not I_78728 (I1341969,I1283416);
nor I_78729 (I1341986,I1341969,I1283422);
nor I_78730 (I1342003,I1341986,I1341808);
DFFARX1 I_78731 (I1342003,I3563,I1341678,I1341667,);
not I_78732 (I1342034,I1341986);
DFFARX1 I_78733 (I1342034,I3563,I1341678,I1342060,);
not I_78734 (I1342068,I1342060);
nor I_78735 (I1341664,I1342068,I1341986);
nor I_78736 (I1342099,I1341969,I1283401);
and I_78737 (I1342116,I1342099,I1283425);
or I_78738 (I1342133,I1342116,I1283407);
DFFARX1 I_78739 (I1342133,I3563,I1341678,I1342159,);
not I_78740 (I1342167,I1342159);
nand I_78741 (I1342184,I1342167,I1341907);
not I_78742 (I1341658,I1342184);
nand I_78743 (I1341652,I1342184,I1341924);
nand I_78744 (I1341649,I1342167,I1341791);
not I_78745 (I1342273,I3570);
DFFARX1 I_78746 (I1210066,I3563,I1342273,I1342299,);
DFFARX1 I_78747 (I1210078,I3563,I1342273,I1342316,);
not I_78748 (I1342324,I1342316);
nor I_78749 (I1342241,I1342299,I1342324);
DFFARX1 I_78750 (I1342324,I3563,I1342273,I1342256,);
nor I_78751 (I1342369,I1210075,I1210069);
and I_78752 (I1342386,I1342369,I1210063);
nor I_78753 (I1342403,I1342386,I1210075);
not I_78754 (I1342420,I1210075);
and I_78755 (I1342437,I1342420,I1210072);
nand I_78756 (I1342454,I1342437,I1210063);
nor I_78757 (I1342471,I1342420,I1342454);
DFFARX1 I_78758 (I1342471,I3563,I1342273,I1342238,);
not I_78759 (I1342502,I1342454);
nand I_78760 (I1342519,I1342324,I1342502);
nand I_78761 (I1342250,I1342386,I1342502);
DFFARX1 I_78762 (I1342420,I3563,I1342273,I1342265,);
not I_78763 (I1342564,I1210087);
nor I_78764 (I1342581,I1342564,I1210072);
nor I_78765 (I1342598,I1342581,I1342403);
DFFARX1 I_78766 (I1342598,I3563,I1342273,I1342262,);
not I_78767 (I1342629,I1342581);
DFFARX1 I_78768 (I1342629,I3563,I1342273,I1342655,);
not I_78769 (I1342663,I1342655);
nor I_78770 (I1342259,I1342663,I1342581);
nor I_78771 (I1342694,I1342564,I1210081);
and I_78772 (I1342711,I1342694,I1210084);
or I_78773 (I1342728,I1342711,I1210066);
DFFARX1 I_78774 (I1342728,I3563,I1342273,I1342754,);
not I_78775 (I1342762,I1342754);
nand I_78776 (I1342779,I1342762,I1342502);
not I_78777 (I1342253,I1342779);
nand I_78778 (I1342247,I1342779,I1342519);
nand I_78779 (I1342244,I1342762,I1342386);
not I_78780 (I1342868,I3570);
DFFARX1 I_78781 (I1040851,I3563,I1342868,I1342894,);
DFFARX1 I_78782 (I1040869,I3563,I1342868,I1342911,);
not I_78783 (I1342919,I1342911);
nor I_78784 (I1342836,I1342894,I1342919);
DFFARX1 I_78785 (I1342919,I3563,I1342868,I1342851,);
nor I_78786 (I1342964,I1040848,I1040860);
and I_78787 (I1342981,I1342964,I1040845);
nor I_78788 (I1342998,I1342981,I1040848);
not I_78789 (I1343015,I1040848);
and I_78790 (I1343032,I1343015,I1040854);
nand I_78791 (I1343049,I1343032,I1040866);
nor I_78792 (I1343066,I1343015,I1343049);
DFFARX1 I_78793 (I1343066,I3563,I1342868,I1342833,);
not I_78794 (I1343097,I1343049);
nand I_78795 (I1343114,I1342919,I1343097);
nand I_78796 (I1342845,I1342981,I1343097);
DFFARX1 I_78797 (I1343015,I3563,I1342868,I1342860,);
not I_78798 (I1343159,I1040857);
nor I_78799 (I1343176,I1343159,I1040854);
nor I_78800 (I1343193,I1343176,I1342998);
DFFARX1 I_78801 (I1343193,I3563,I1342868,I1342857,);
not I_78802 (I1343224,I1343176);
DFFARX1 I_78803 (I1343224,I3563,I1342868,I1343250,);
not I_78804 (I1343258,I1343250);
nor I_78805 (I1342854,I1343258,I1343176);
nor I_78806 (I1343289,I1343159,I1040845);
and I_78807 (I1343306,I1343289,I1040872);
or I_78808 (I1343323,I1343306,I1040863);
DFFARX1 I_78809 (I1343323,I3563,I1342868,I1343349,);
not I_78810 (I1343357,I1343349);
nand I_78811 (I1343374,I1343357,I1343097);
not I_78812 (I1342848,I1343374);
nand I_78813 (I1342842,I1343374,I1343114);
nand I_78814 (I1342839,I1343357,I1342981);
not I_78815 (I1343463,I3570);
DFFARX1 I_78816 (I1052842,I3563,I1343463,I1343489,);
DFFARX1 I_78817 (I1052833,I3563,I1343463,I1343506,);
not I_78818 (I1343514,I1343506);
nor I_78819 (I1343431,I1343489,I1343514);
DFFARX1 I_78820 (I1343514,I3563,I1343463,I1343446,);
nor I_78821 (I1343559,I1052839,I1052848);
and I_78822 (I1343576,I1343559,I1052851);
nor I_78823 (I1343593,I1343576,I1052839);
not I_78824 (I1343610,I1052839);
and I_78825 (I1343627,I1343610,I1052830);
nand I_78826 (I1343644,I1343627,I1052836);
nor I_78827 (I1343661,I1343610,I1343644);
DFFARX1 I_78828 (I1343661,I3563,I1343463,I1343428,);
not I_78829 (I1343692,I1343644);
nand I_78830 (I1343709,I1343514,I1343692);
nand I_78831 (I1343440,I1343576,I1343692);
DFFARX1 I_78832 (I1343610,I3563,I1343463,I1343455,);
not I_78833 (I1343754,I1052845);
nor I_78834 (I1343771,I1343754,I1052830);
nor I_78835 (I1343788,I1343771,I1343593);
DFFARX1 I_78836 (I1343788,I3563,I1343463,I1343452,);
not I_78837 (I1343819,I1343771);
DFFARX1 I_78838 (I1343819,I3563,I1343463,I1343845,);
not I_78839 (I1343853,I1343845);
nor I_78840 (I1343449,I1343853,I1343771);
nor I_78841 (I1343884,I1343754,I1052830);
and I_78842 (I1343901,I1343884,I1052833);
or I_78843 (I1343918,I1343901,I1052836);
DFFARX1 I_78844 (I1343918,I3563,I1343463,I1343944,);
not I_78845 (I1343952,I1343944);
nand I_78846 (I1343969,I1343952,I1343692);
not I_78847 (I1343443,I1343969);
nand I_78848 (I1343437,I1343969,I1343709);
nand I_78849 (I1343434,I1343952,I1343576);
not I_78850 (I1344058,I3570);
DFFARX1 I_78851 (I997569,I3563,I1344058,I1344084,);
DFFARX1 I_78852 (I997587,I3563,I1344058,I1344101,);
not I_78853 (I1344109,I1344101);
nor I_78854 (I1344026,I1344084,I1344109);
DFFARX1 I_78855 (I1344109,I3563,I1344058,I1344041,);
nor I_78856 (I1344154,I997566,I997578);
and I_78857 (I1344171,I1344154,I997563);
nor I_78858 (I1344188,I1344171,I997566);
not I_78859 (I1344205,I997566);
and I_78860 (I1344222,I1344205,I997572);
nand I_78861 (I1344239,I1344222,I997584);
nor I_78862 (I1344256,I1344205,I1344239);
DFFARX1 I_78863 (I1344256,I3563,I1344058,I1344023,);
not I_78864 (I1344287,I1344239);
nand I_78865 (I1344304,I1344109,I1344287);
nand I_78866 (I1344035,I1344171,I1344287);
DFFARX1 I_78867 (I1344205,I3563,I1344058,I1344050,);
not I_78868 (I1344349,I997575);
nor I_78869 (I1344366,I1344349,I997572);
nor I_78870 (I1344383,I1344366,I1344188);
DFFARX1 I_78871 (I1344383,I3563,I1344058,I1344047,);
not I_78872 (I1344414,I1344366);
DFFARX1 I_78873 (I1344414,I3563,I1344058,I1344440,);
not I_78874 (I1344448,I1344440);
nor I_78875 (I1344044,I1344448,I1344366);
nor I_78876 (I1344479,I1344349,I997563);
and I_78877 (I1344496,I1344479,I997590);
or I_78878 (I1344513,I1344496,I997581);
DFFARX1 I_78879 (I1344513,I3563,I1344058,I1344539,);
not I_78880 (I1344547,I1344539);
nand I_78881 (I1344564,I1344547,I1344287);
not I_78882 (I1344038,I1344564);
nand I_78883 (I1344032,I1344564,I1344304);
nand I_78884 (I1344029,I1344547,I1344171);
not I_78885 (I1344653,I3570);
DFFARX1 I_78886 (I1197350,I3563,I1344653,I1344679,);
DFFARX1 I_78887 (I1197362,I3563,I1344653,I1344696,);
not I_78888 (I1344704,I1344696);
nor I_78889 (I1344621,I1344679,I1344704);
DFFARX1 I_78890 (I1344704,I3563,I1344653,I1344636,);
nor I_78891 (I1344749,I1197359,I1197353);
and I_78892 (I1344766,I1344749,I1197347);
nor I_78893 (I1344783,I1344766,I1197359);
not I_78894 (I1344800,I1197359);
and I_78895 (I1344817,I1344800,I1197356);
nand I_78896 (I1344834,I1344817,I1197347);
nor I_78897 (I1344851,I1344800,I1344834);
DFFARX1 I_78898 (I1344851,I3563,I1344653,I1344618,);
not I_78899 (I1344882,I1344834);
nand I_78900 (I1344899,I1344704,I1344882);
nand I_78901 (I1344630,I1344766,I1344882);
DFFARX1 I_78902 (I1344800,I3563,I1344653,I1344645,);
not I_78903 (I1344944,I1197371);
nor I_78904 (I1344961,I1344944,I1197356);
nor I_78905 (I1344978,I1344961,I1344783);
DFFARX1 I_78906 (I1344978,I3563,I1344653,I1344642,);
not I_78907 (I1345009,I1344961);
DFFARX1 I_78908 (I1345009,I3563,I1344653,I1345035,);
not I_78909 (I1345043,I1345035);
nor I_78910 (I1344639,I1345043,I1344961);
nor I_78911 (I1345074,I1344944,I1197365);
and I_78912 (I1345091,I1345074,I1197368);
or I_78913 (I1345108,I1345091,I1197350);
DFFARX1 I_78914 (I1345108,I3563,I1344653,I1345134,);
not I_78915 (I1345142,I1345134);
nand I_78916 (I1345159,I1345142,I1344882);
not I_78917 (I1344633,I1345159);
nand I_78918 (I1344627,I1345159,I1344899);
nand I_78919 (I1344624,I1345142,I1344766);
not I_78920 (I1345248,I3570);
DFFARX1 I_78921 (I292764,I3563,I1345248,I1345274,);
DFFARX1 I_78922 (I292758,I3563,I1345248,I1345291,);
not I_78923 (I1345299,I1345291);
nor I_78924 (I1345216,I1345274,I1345299);
DFFARX1 I_78925 (I1345299,I3563,I1345248,I1345231,);
nor I_78926 (I1345344,I292746,I292767);
and I_78927 (I1345361,I1345344,I292761);
nor I_78928 (I1345378,I1345361,I292746);
not I_78929 (I1345395,I292746);
and I_78930 (I1345412,I1345395,I292743);
nand I_78931 (I1345429,I1345412,I292755);
nor I_78932 (I1345446,I1345395,I1345429);
DFFARX1 I_78933 (I1345446,I3563,I1345248,I1345213,);
not I_78934 (I1345477,I1345429);
nand I_78935 (I1345494,I1345299,I1345477);
nand I_78936 (I1345225,I1345361,I1345477);
DFFARX1 I_78937 (I1345395,I3563,I1345248,I1345240,);
not I_78938 (I1345539,I292770);
nor I_78939 (I1345556,I1345539,I292743);
nor I_78940 (I1345573,I1345556,I1345378);
DFFARX1 I_78941 (I1345573,I3563,I1345248,I1345237,);
not I_78942 (I1345604,I1345556);
DFFARX1 I_78943 (I1345604,I3563,I1345248,I1345630,);
not I_78944 (I1345638,I1345630);
nor I_78945 (I1345234,I1345638,I1345556);
nor I_78946 (I1345669,I1345539,I292752);
and I_78947 (I1345686,I1345669,I292749);
or I_78948 (I1345703,I1345686,I292743);
DFFARX1 I_78949 (I1345703,I3563,I1345248,I1345729,);
not I_78950 (I1345737,I1345729);
nand I_78951 (I1345754,I1345737,I1345477);
not I_78952 (I1345228,I1345754);
nand I_78953 (I1345222,I1345754,I1345494);
nand I_78954 (I1345219,I1345737,I1345361);
not I_78955 (I1345843,I3570);
DFFARX1 I_78956 (I319114,I3563,I1345843,I1345869,);
DFFARX1 I_78957 (I319108,I3563,I1345843,I1345886,);
not I_78958 (I1345894,I1345886);
nor I_78959 (I1345811,I1345869,I1345894);
DFFARX1 I_78960 (I1345894,I3563,I1345843,I1345826,);
nor I_78961 (I1345939,I319096,I319117);
and I_78962 (I1345956,I1345939,I319111);
nor I_78963 (I1345973,I1345956,I319096);
not I_78964 (I1345990,I319096);
and I_78965 (I1346007,I1345990,I319093);
nand I_78966 (I1346024,I1346007,I319105);
nor I_78967 (I1346041,I1345990,I1346024);
DFFARX1 I_78968 (I1346041,I3563,I1345843,I1345808,);
not I_78969 (I1346072,I1346024);
nand I_78970 (I1346089,I1345894,I1346072);
nand I_78971 (I1345820,I1345956,I1346072);
DFFARX1 I_78972 (I1345990,I3563,I1345843,I1345835,);
not I_78973 (I1346134,I319120);
nor I_78974 (I1346151,I1346134,I319093);
nor I_78975 (I1346168,I1346151,I1345973);
DFFARX1 I_78976 (I1346168,I3563,I1345843,I1345832,);
not I_78977 (I1346199,I1346151);
DFFARX1 I_78978 (I1346199,I3563,I1345843,I1346225,);
not I_78979 (I1346233,I1346225);
nor I_78980 (I1345829,I1346233,I1346151);
nor I_78981 (I1346264,I1346134,I319102);
and I_78982 (I1346281,I1346264,I319099);
or I_78983 (I1346298,I1346281,I319093);
DFFARX1 I_78984 (I1346298,I3563,I1345843,I1346324,);
not I_78985 (I1346332,I1346324);
nand I_78986 (I1346349,I1346332,I1346072);
not I_78987 (I1345823,I1346349);
nand I_78988 (I1345817,I1346349,I1346089);
nand I_78989 (I1345814,I1346332,I1345956);
not I_78990 (I1346438,I3570);
DFFARX1 I_78991 (I1231452,I3563,I1346438,I1346464,);
DFFARX1 I_78992 (I1231464,I3563,I1346438,I1346481,);
not I_78993 (I1346489,I1346481);
nor I_78994 (I1346406,I1346464,I1346489);
DFFARX1 I_78995 (I1346489,I3563,I1346438,I1346421,);
nor I_78996 (I1346534,I1231461,I1231455);
and I_78997 (I1346551,I1346534,I1231449);
nor I_78998 (I1346568,I1346551,I1231461);
not I_78999 (I1346585,I1231461);
and I_79000 (I1346602,I1346585,I1231458);
nand I_79001 (I1346619,I1346602,I1231449);
nor I_79002 (I1346636,I1346585,I1346619);
DFFARX1 I_79003 (I1346636,I3563,I1346438,I1346403,);
not I_79004 (I1346667,I1346619);
nand I_79005 (I1346684,I1346489,I1346667);
nand I_79006 (I1346415,I1346551,I1346667);
DFFARX1 I_79007 (I1346585,I3563,I1346438,I1346430,);
not I_79008 (I1346729,I1231473);
nor I_79009 (I1346746,I1346729,I1231458);
nor I_79010 (I1346763,I1346746,I1346568);
DFFARX1 I_79011 (I1346763,I3563,I1346438,I1346427,);
not I_79012 (I1346794,I1346746);
DFFARX1 I_79013 (I1346794,I3563,I1346438,I1346820,);
not I_79014 (I1346828,I1346820);
nor I_79015 (I1346424,I1346828,I1346746);
nor I_79016 (I1346859,I1346729,I1231467);
and I_79017 (I1346876,I1346859,I1231470);
or I_79018 (I1346893,I1346876,I1231452);
DFFARX1 I_79019 (I1346893,I3563,I1346438,I1346919,);
not I_79020 (I1346927,I1346919);
nand I_79021 (I1346944,I1346927,I1346667);
not I_79022 (I1346418,I1346944);
nand I_79023 (I1346412,I1346944,I1346684);
nand I_79024 (I1346409,I1346927,I1346551);
not I_79025 (I1347033,I3570);
DFFARX1 I_79026 (I209528,I3563,I1347033,I1347059,);
DFFARX1 I_79027 (I209531,I3563,I1347033,I1347076,);
not I_79028 (I1347084,I1347076);
nor I_79029 (I1347001,I1347059,I1347084);
DFFARX1 I_79030 (I1347084,I3563,I1347033,I1347016,);
nor I_79031 (I1347129,I209537,I209531);
and I_79032 (I1347146,I1347129,I209534);
nor I_79033 (I1347163,I1347146,I209537);
not I_79034 (I1347180,I209537);
and I_79035 (I1347197,I1347180,I209528);
nand I_79036 (I1347214,I1347197,I209546);
nor I_79037 (I1347231,I1347180,I1347214);
DFFARX1 I_79038 (I1347231,I3563,I1347033,I1346998,);
not I_79039 (I1347262,I1347214);
nand I_79040 (I1347279,I1347084,I1347262);
nand I_79041 (I1347010,I1347146,I1347262);
DFFARX1 I_79042 (I1347180,I3563,I1347033,I1347025,);
not I_79043 (I1347324,I209540);
nor I_79044 (I1347341,I1347324,I209528);
nor I_79045 (I1347358,I1347341,I1347163);
DFFARX1 I_79046 (I1347358,I3563,I1347033,I1347022,);
not I_79047 (I1347389,I1347341);
DFFARX1 I_79048 (I1347389,I3563,I1347033,I1347415,);
not I_79049 (I1347423,I1347415);
nor I_79050 (I1347019,I1347423,I1347341);
nor I_79051 (I1347454,I1347324,I209543);
and I_79052 (I1347471,I1347454,I209549);
or I_79053 (I1347488,I1347471,I209552);
DFFARX1 I_79054 (I1347488,I3563,I1347033,I1347514,);
not I_79055 (I1347522,I1347514);
nand I_79056 (I1347539,I1347522,I1347262);
not I_79057 (I1347013,I1347539);
nand I_79058 (I1347007,I1347539,I1347279);
nand I_79059 (I1347004,I1347522,I1347146);
not I_79060 (I1347628,I3570);
DFFARX1 I_79061 (I598322,I3563,I1347628,I1347654,);
DFFARX1 I_79062 (I598316,I3563,I1347628,I1347671,);
not I_79063 (I1347679,I1347671);
nor I_79064 (I1347596,I1347654,I1347679);
DFFARX1 I_79065 (I1347679,I3563,I1347628,I1347611,);
nor I_79066 (I1347724,I598313,I598304);
and I_79067 (I1347741,I1347724,I598301);
nor I_79068 (I1347758,I1347741,I598313);
not I_79069 (I1347775,I598313);
and I_79070 (I1347792,I1347775,I598307);
nand I_79071 (I1347809,I1347792,I598319);
nor I_79072 (I1347826,I1347775,I1347809);
DFFARX1 I_79073 (I1347826,I3563,I1347628,I1347593,);
not I_79074 (I1347857,I1347809);
nand I_79075 (I1347874,I1347679,I1347857);
nand I_79076 (I1347605,I1347741,I1347857);
DFFARX1 I_79077 (I1347775,I3563,I1347628,I1347620,);
not I_79078 (I1347919,I598325);
nor I_79079 (I1347936,I1347919,I598307);
nor I_79080 (I1347953,I1347936,I1347758);
DFFARX1 I_79081 (I1347953,I3563,I1347628,I1347617,);
not I_79082 (I1347984,I1347936);
DFFARX1 I_79083 (I1347984,I3563,I1347628,I1348010,);
not I_79084 (I1348018,I1348010);
nor I_79085 (I1347614,I1348018,I1347936);
nor I_79086 (I1348049,I1347919,I598304);
and I_79087 (I1348066,I1348049,I598310);
or I_79088 (I1348083,I1348066,I598301);
DFFARX1 I_79089 (I1348083,I3563,I1347628,I1348109,);
not I_79090 (I1348117,I1348109);
nand I_79091 (I1348134,I1348117,I1347857);
not I_79092 (I1347608,I1348134);
nand I_79093 (I1347602,I1348134,I1347874);
nand I_79094 (I1347599,I1348117,I1347741);
not I_79095 (I1348223,I3570);
DFFARX1 I_79096 (I973021,I3563,I1348223,I1348249,);
DFFARX1 I_79097 (I973039,I3563,I1348223,I1348266,);
not I_79098 (I1348274,I1348266);
nor I_79099 (I1348191,I1348249,I1348274);
DFFARX1 I_79100 (I1348274,I3563,I1348223,I1348206,);
nor I_79101 (I1348319,I973018,I973030);
and I_79102 (I1348336,I1348319,I973015);
nor I_79103 (I1348353,I1348336,I973018);
not I_79104 (I1348370,I973018);
and I_79105 (I1348387,I1348370,I973024);
nand I_79106 (I1348404,I1348387,I973036);
nor I_79107 (I1348421,I1348370,I1348404);
DFFARX1 I_79108 (I1348421,I3563,I1348223,I1348188,);
not I_79109 (I1348452,I1348404);
nand I_79110 (I1348469,I1348274,I1348452);
nand I_79111 (I1348200,I1348336,I1348452);
DFFARX1 I_79112 (I1348370,I3563,I1348223,I1348215,);
not I_79113 (I1348514,I973027);
nor I_79114 (I1348531,I1348514,I973024);
nor I_79115 (I1348548,I1348531,I1348353);
DFFARX1 I_79116 (I1348548,I3563,I1348223,I1348212,);
not I_79117 (I1348579,I1348531);
DFFARX1 I_79118 (I1348579,I3563,I1348223,I1348605,);
not I_79119 (I1348613,I1348605);
nor I_79120 (I1348209,I1348613,I1348531);
nor I_79121 (I1348644,I1348514,I973015);
and I_79122 (I1348661,I1348644,I973042);
or I_79123 (I1348678,I1348661,I973033);
DFFARX1 I_79124 (I1348678,I3563,I1348223,I1348704,);
not I_79125 (I1348712,I1348704);
nand I_79126 (I1348729,I1348712,I1348452);
not I_79127 (I1348203,I1348729);
nand I_79128 (I1348197,I1348729,I1348469);
nand I_79129 (I1348194,I1348712,I1348336);
not I_79130 (I1348818,I3570);
DFFARX1 I_79131 (I972375,I3563,I1348818,I1348844,);
DFFARX1 I_79132 (I972393,I3563,I1348818,I1348861,);
not I_79133 (I1348869,I1348861);
nor I_79134 (I1348786,I1348844,I1348869);
DFFARX1 I_79135 (I1348869,I3563,I1348818,I1348801,);
nor I_79136 (I1348914,I972372,I972384);
and I_79137 (I1348931,I1348914,I972369);
nor I_79138 (I1348948,I1348931,I972372);
not I_79139 (I1348965,I972372);
and I_79140 (I1348982,I1348965,I972378);
nand I_79141 (I1348999,I1348982,I972390);
nor I_79142 (I1349016,I1348965,I1348999);
DFFARX1 I_79143 (I1349016,I3563,I1348818,I1348783,);
not I_79144 (I1349047,I1348999);
nand I_79145 (I1349064,I1348869,I1349047);
nand I_79146 (I1348795,I1348931,I1349047);
DFFARX1 I_79147 (I1348965,I3563,I1348818,I1348810,);
not I_79148 (I1349109,I972381);
nor I_79149 (I1349126,I1349109,I972378);
nor I_79150 (I1349143,I1349126,I1348948);
DFFARX1 I_79151 (I1349143,I3563,I1348818,I1348807,);
not I_79152 (I1349174,I1349126);
DFFARX1 I_79153 (I1349174,I3563,I1348818,I1349200,);
not I_79154 (I1349208,I1349200);
nor I_79155 (I1348804,I1349208,I1349126);
nor I_79156 (I1349239,I1349109,I972369);
and I_79157 (I1349256,I1349239,I972396);
or I_79158 (I1349273,I1349256,I972387);
DFFARX1 I_79159 (I1349273,I3563,I1348818,I1349299,);
not I_79160 (I1349307,I1349299);
nand I_79161 (I1349324,I1349307,I1349047);
not I_79162 (I1348798,I1349324);
nand I_79163 (I1348792,I1349324,I1349064);
nand I_79164 (I1348789,I1349307,I1348931);
not I_79165 (I1349413,I3570);
DFFARX1 I_79166 (I1281225,I3563,I1349413,I1349439,);
DFFARX1 I_79167 (I1281228,I3563,I1349413,I1349456,);
not I_79168 (I1349464,I1349456);
nor I_79169 (I1349381,I1349439,I1349464);
DFFARX1 I_79170 (I1349464,I3563,I1349413,I1349396,);
nor I_79171 (I1349509,I1281228,I1281243);
and I_79172 (I1349526,I1349509,I1281237);
nor I_79173 (I1349543,I1349526,I1281228);
not I_79174 (I1349560,I1281228);
and I_79175 (I1349577,I1349560,I1281246);
nand I_79176 (I1349594,I1349577,I1281234);
nor I_79177 (I1349611,I1349560,I1349594);
DFFARX1 I_79178 (I1349611,I3563,I1349413,I1349378,);
not I_79179 (I1349642,I1349594);
nand I_79180 (I1349659,I1349464,I1349642);
nand I_79181 (I1349390,I1349526,I1349642);
DFFARX1 I_79182 (I1349560,I3563,I1349413,I1349405,);
not I_79183 (I1349704,I1281240);
nor I_79184 (I1349721,I1349704,I1281246);
nor I_79185 (I1349738,I1349721,I1349543);
DFFARX1 I_79186 (I1349738,I3563,I1349413,I1349402,);
not I_79187 (I1349769,I1349721);
DFFARX1 I_79188 (I1349769,I3563,I1349413,I1349795,);
not I_79189 (I1349803,I1349795);
nor I_79190 (I1349399,I1349803,I1349721);
nor I_79191 (I1349834,I1349704,I1281225);
and I_79192 (I1349851,I1349834,I1281249);
or I_79193 (I1349868,I1349851,I1281231);
DFFARX1 I_79194 (I1349868,I3563,I1349413,I1349894,);
not I_79195 (I1349902,I1349894);
nand I_79196 (I1349919,I1349902,I1349642);
not I_79197 (I1349393,I1349919);
nand I_79198 (I1349387,I1349919,I1349659);
nand I_79199 (I1349384,I1349902,I1349526);
not I_79200 (I1350008,I3570);
DFFARX1 I_79201 (I293291,I3563,I1350008,I1350034,);
DFFARX1 I_79202 (I293285,I3563,I1350008,I1350051,);
not I_79203 (I1350059,I1350051);
nor I_79204 (I1349976,I1350034,I1350059);
DFFARX1 I_79205 (I1350059,I3563,I1350008,I1349991,);
nor I_79206 (I1350104,I293273,I293294);
and I_79207 (I1350121,I1350104,I293288);
nor I_79208 (I1350138,I1350121,I293273);
not I_79209 (I1350155,I293273);
and I_79210 (I1350172,I1350155,I293270);
nand I_79211 (I1350189,I1350172,I293282);
nor I_79212 (I1350206,I1350155,I1350189);
DFFARX1 I_79213 (I1350206,I3563,I1350008,I1349973,);
not I_79214 (I1350237,I1350189);
nand I_79215 (I1350254,I1350059,I1350237);
nand I_79216 (I1349985,I1350121,I1350237);
DFFARX1 I_79217 (I1350155,I3563,I1350008,I1350000,);
not I_79218 (I1350299,I293297);
nor I_79219 (I1350316,I1350299,I293270);
nor I_79220 (I1350333,I1350316,I1350138);
DFFARX1 I_79221 (I1350333,I3563,I1350008,I1349997,);
not I_79222 (I1350364,I1350316);
DFFARX1 I_79223 (I1350364,I3563,I1350008,I1350390,);
not I_79224 (I1350398,I1350390);
nor I_79225 (I1349994,I1350398,I1350316);
nor I_79226 (I1350429,I1350299,I293279);
and I_79227 (I1350446,I1350429,I293276);
or I_79228 (I1350463,I1350446,I293270);
DFFARX1 I_79229 (I1350463,I3563,I1350008,I1350489,);
not I_79230 (I1350497,I1350489);
nand I_79231 (I1350514,I1350497,I1350237);
not I_79232 (I1349988,I1350514);
nand I_79233 (I1349982,I1350514,I1350254);
nand I_79234 (I1349979,I1350497,I1350121);
not I_79235 (I1350603,I3570);
DFFARX1 I_79236 (I177398,I3563,I1350603,I1350629,);
DFFARX1 I_79237 (I177401,I3563,I1350603,I1350646,);
not I_79238 (I1350654,I1350646);
nor I_79239 (I1350571,I1350629,I1350654);
DFFARX1 I_79240 (I1350654,I3563,I1350603,I1350586,);
nor I_79241 (I1350699,I177407,I177401);
and I_79242 (I1350716,I1350699,I177404);
nor I_79243 (I1350733,I1350716,I177407);
not I_79244 (I1350750,I177407);
and I_79245 (I1350767,I1350750,I177398);
nand I_79246 (I1350784,I1350767,I177416);
nor I_79247 (I1350801,I1350750,I1350784);
DFFARX1 I_79248 (I1350801,I3563,I1350603,I1350568,);
not I_79249 (I1350832,I1350784);
nand I_79250 (I1350849,I1350654,I1350832);
nand I_79251 (I1350580,I1350716,I1350832);
DFFARX1 I_79252 (I1350750,I3563,I1350603,I1350595,);
not I_79253 (I1350894,I177410);
nor I_79254 (I1350911,I1350894,I177398);
nor I_79255 (I1350928,I1350911,I1350733);
DFFARX1 I_79256 (I1350928,I3563,I1350603,I1350592,);
not I_79257 (I1350959,I1350911);
DFFARX1 I_79258 (I1350959,I3563,I1350603,I1350985,);
not I_79259 (I1350993,I1350985);
nor I_79260 (I1350589,I1350993,I1350911);
nor I_79261 (I1351024,I1350894,I177413);
and I_79262 (I1351041,I1351024,I177419);
or I_79263 (I1351058,I1351041,I177422);
DFFARX1 I_79264 (I1351058,I3563,I1350603,I1351084,);
not I_79265 (I1351092,I1351084);
nand I_79266 (I1351109,I1351092,I1350832);
not I_79267 (I1350583,I1351109);
nand I_79268 (I1350577,I1351109,I1350849);
nand I_79269 (I1350574,I1351092,I1350716);
not I_79270 (I1351198,I3570);
DFFARX1 I_79271 (I507810,I3563,I1351198,I1351224,);
DFFARX1 I_79272 (I507816,I3563,I1351198,I1351241,);
not I_79273 (I1351249,I1351241);
nor I_79274 (I1351166,I1351224,I1351249);
DFFARX1 I_79275 (I1351249,I3563,I1351198,I1351181,);
nor I_79276 (I1351294,I507825,I507810);
and I_79277 (I1351311,I1351294,I507837);
nor I_79278 (I1351328,I1351311,I507825);
not I_79279 (I1351345,I507825);
and I_79280 (I1351362,I1351345,I507813);
nand I_79281 (I1351379,I1351362,I507834);
nor I_79282 (I1351396,I1351345,I1351379);
DFFARX1 I_79283 (I1351396,I3563,I1351198,I1351163,);
not I_79284 (I1351427,I1351379);
nand I_79285 (I1351444,I1351249,I1351427);
nand I_79286 (I1351175,I1351311,I1351427);
DFFARX1 I_79287 (I1351345,I3563,I1351198,I1351190,);
not I_79288 (I1351489,I507822);
nor I_79289 (I1351506,I1351489,I507813);
nor I_79290 (I1351523,I1351506,I1351328);
DFFARX1 I_79291 (I1351523,I3563,I1351198,I1351187,);
not I_79292 (I1351554,I1351506);
DFFARX1 I_79293 (I1351554,I3563,I1351198,I1351580,);
not I_79294 (I1351588,I1351580);
nor I_79295 (I1351184,I1351588,I1351506);
nor I_79296 (I1351619,I1351489,I507819);
and I_79297 (I1351636,I1351619,I507831);
or I_79298 (I1351653,I1351636,I507828);
DFFARX1 I_79299 (I1351653,I3563,I1351198,I1351679,);
not I_79300 (I1351687,I1351679);
nand I_79301 (I1351704,I1351687,I1351427);
not I_79302 (I1351178,I1351704);
nand I_79303 (I1351172,I1351704,I1351444);
nand I_79304 (I1351169,I1351687,I1351311);
not I_79305 (I1351793,I3570);
DFFARX1 I_79306 (I426754,I3563,I1351793,I1351819,);
DFFARX1 I_79307 (I426760,I3563,I1351793,I1351836,);
not I_79308 (I1351844,I1351836);
nor I_79309 (I1351761,I1351819,I1351844);
DFFARX1 I_79310 (I1351844,I3563,I1351793,I1351776,);
nor I_79311 (I1351889,I426769,I426754);
and I_79312 (I1351906,I1351889,I426781);
nor I_79313 (I1351923,I1351906,I426769);
not I_79314 (I1351940,I426769);
and I_79315 (I1351957,I1351940,I426757);
nand I_79316 (I1351974,I1351957,I426778);
nor I_79317 (I1351991,I1351940,I1351974);
DFFARX1 I_79318 (I1351991,I3563,I1351793,I1351758,);
not I_79319 (I1352022,I1351974);
nand I_79320 (I1352039,I1351844,I1352022);
nand I_79321 (I1351770,I1351906,I1352022);
DFFARX1 I_79322 (I1351940,I3563,I1351793,I1351785,);
not I_79323 (I1352084,I426766);
nor I_79324 (I1352101,I1352084,I426757);
nor I_79325 (I1352118,I1352101,I1351923);
DFFARX1 I_79326 (I1352118,I3563,I1351793,I1351782,);
not I_79327 (I1352149,I1352101);
DFFARX1 I_79328 (I1352149,I3563,I1351793,I1352175,);
not I_79329 (I1352183,I1352175);
nor I_79330 (I1351779,I1352183,I1352101);
nor I_79331 (I1352214,I1352084,I426763);
and I_79332 (I1352231,I1352214,I426775);
or I_79333 (I1352248,I1352231,I426772);
DFFARX1 I_79334 (I1352248,I3563,I1351793,I1352274,);
not I_79335 (I1352282,I1352274);
nand I_79336 (I1352299,I1352282,I1352022);
not I_79337 (I1351773,I1352299);
nand I_79338 (I1351767,I1352299,I1352039);
nand I_79339 (I1351764,I1352282,I1351906);
not I_79340 (I1352388,I3570);
DFFARX1 I_79341 (I1252393,I3563,I1352388,I1352414,);
DFFARX1 I_79342 (I1252396,I3563,I1352388,I1352431,);
not I_79343 (I1352439,I1352431);
nor I_79344 (I1352356,I1352414,I1352439);
DFFARX1 I_79345 (I1352439,I3563,I1352388,I1352371,);
nor I_79346 (I1352484,I1252396,I1252411);
and I_79347 (I1352501,I1352484,I1252405);
nor I_79348 (I1352518,I1352501,I1252396);
not I_79349 (I1352535,I1252396);
and I_79350 (I1352552,I1352535,I1252414);
nand I_79351 (I1352569,I1352552,I1252402);
nor I_79352 (I1352586,I1352535,I1352569);
DFFARX1 I_79353 (I1352586,I3563,I1352388,I1352353,);
not I_79354 (I1352617,I1352569);
nand I_79355 (I1352634,I1352439,I1352617);
nand I_79356 (I1352365,I1352501,I1352617);
DFFARX1 I_79357 (I1352535,I3563,I1352388,I1352380,);
not I_79358 (I1352679,I1252408);
nor I_79359 (I1352696,I1352679,I1252414);
nor I_79360 (I1352713,I1352696,I1352518);
DFFARX1 I_79361 (I1352713,I3563,I1352388,I1352377,);
not I_79362 (I1352744,I1352696);
DFFARX1 I_79363 (I1352744,I3563,I1352388,I1352770,);
not I_79364 (I1352778,I1352770);
nor I_79365 (I1352374,I1352778,I1352696);
nor I_79366 (I1352809,I1352679,I1252393);
and I_79367 (I1352826,I1352809,I1252417);
or I_79368 (I1352843,I1352826,I1252399);
DFFARX1 I_79369 (I1352843,I3563,I1352388,I1352869,);
not I_79370 (I1352877,I1352869);
nand I_79371 (I1352894,I1352877,I1352617);
not I_79372 (I1352368,I1352894);
nand I_79373 (I1352362,I1352894,I1352634);
nand I_79374 (I1352359,I1352877,I1352501);
not I_79375 (I1352983,I3570);
DFFARX1 I_79376 (I1312047,I3563,I1352983,I1353009,);
DFFARX1 I_79377 (I1312038,I3563,I1352983,I1353026,);
not I_79378 (I1353034,I1353026);
nor I_79379 (I1352951,I1353009,I1353034);
DFFARX1 I_79380 (I1353034,I3563,I1352983,I1352966,);
nor I_79381 (I1353079,I1312029,I1312044);
and I_79382 (I1353096,I1353079,I1312032);
nor I_79383 (I1353113,I1353096,I1312029);
not I_79384 (I1353130,I1312029);
and I_79385 (I1353147,I1353130,I1312035);
nand I_79386 (I1353164,I1353147,I1312053);
nor I_79387 (I1353181,I1353130,I1353164);
DFFARX1 I_79388 (I1353181,I3563,I1352983,I1352948,);
not I_79389 (I1353212,I1353164);
nand I_79390 (I1353229,I1353034,I1353212);
nand I_79391 (I1352960,I1353096,I1353212);
DFFARX1 I_79392 (I1353130,I3563,I1352983,I1352975,);
not I_79393 (I1353274,I1312029);
nor I_79394 (I1353291,I1353274,I1312035);
nor I_79395 (I1353308,I1353291,I1353113);
DFFARX1 I_79396 (I1353308,I3563,I1352983,I1352972,);
not I_79397 (I1353339,I1353291);
DFFARX1 I_79398 (I1353339,I3563,I1352983,I1353365,);
not I_79399 (I1353373,I1353365);
nor I_79400 (I1352969,I1353373,I1353291);
nor I_79401 (I1353404,I1353274,I1312032);
and I_79402 (I1353421,I1353404,I1312041);
or I_79403 (I1353438,I1353421,I1312050);
DFFARX1 I_79404 (I1353438,I3563,I1352983,I1353464,);
not I_79405 (I1353472,I1353464);
nand I_79406 (I1353489,I1353472,I1353212);
not I_79407 (I1352963,I1353489);
nand I_79408 (I1352957,I1353489,I1353229);
nand I_79409 (I1352954,I1353472,I1353096);
not I_79410 (I1353578,I3570);
DFFARX1 I_79411 (I255938,I3563,I1353578,I1353604,);
DFFARX1 I_79412 (I255941,I3563,I1353578,I1353621,);
not I_79413 (I1353629,I1353621);
nor I_79414 (I1353546,I1353604,I1353629);
DFFARX1 I_79415 (I1353629,I3563,I1353578,I1353561,);
nor I_79416 (I1353674,I255947,I255941);
and I_79417 (I1353691,I1353674,I255944);
nor I_79418 (I1353708,I1353691,I255947);
not I_79419 (I1353725,I255947);
and I_79420 (I1353742,I1353725,I255938);
nand I_79421 (I1353759,I1353742,I255956);
nor I_79422 (I1353776,I1353725,I1353759);
DFFARX1 I_79423 (I1353776,I3563,I1353578,I1353543,);
not I_79424 (I1353807,I1353759);
nand I_79425 (I1353824,I1353629,I1353807);
nand I_79426 (I1353555,I1353691,I1353807);
DFFARX1 I_79427 (I1353725,I3563,I1353578,I1353570,);
not I_79428 (I1353869,I255950);
nor I_79429 (I1353886,I1353869,I255938);
nor I_79430 (I1353903,I1353886,I1353708);
DFFARX1 I_79431 (I1353903,I3563,I1353578,I1353567,);
not I_79432 (I1353934,I1353886);
DFFARX1 I_79433 (I1353934,I3563,I1353578,I1353960,);
not I_79434 (I1353968,I1353960);
nor I_79435 (I1353564,I1353968,I1353886);
nor I_79436 (I1353999,I1353869,I255953);
and I_79437 (I1354016,I1353999,I255959);
or I_79438 (I1354033,I1354016,I255962);
DFFARX1 I_79439 (I1354033,I3563,I1353578,I1354059,);
not I_79440 (I1354067,I1354059);
nand I_79441 (I1354084,I1354067,I1353807);
not I_79442 (I1353558,I1354084);
nand I_79443 (I1353552,I1354084,I1353824);
nand I_79444 (I1353549,I1354067,I1353691);
not I_79445 (I1354173,I3570);
DFFARX1 I_79446 (I895385,I3563,I1354173,I1354199,);
DFFARX1 I_79447 (I895382,I3563,I1354173,I1354216,);
not I_79448 (I1354224,I1354216);
nor I_79449 (I1354141,I1354199,I1354224);
DFFARX1 I_79450 (I1354224,I3563,I1354173,I1354156,);
nor I_79451 (I1354269,I895397,I895379);
and I_79452 (I1354286,I1354269,I895376);
nor I_79453 (I1354303,I1354286,I895397);
not I_79454 (I1354320,I895397);
and I_79455 (I1354337,I1354320,I895382);
nand I_79456 (I1354354,I1354337,I895394);
nor I_79457 (I1354371,I1354320,I1354354);
DFFARX1 I_79458 (I1354371,I3563,I1354173,I1354138,);
not I_79459 (I1354402,I1354354);
nand I_79460 (I1354419,I1354224,I1354402);
nand I_79461 (I1354150,I1354286,I1354402);
DFFARX1 I_79462 (I1354320,I3563,I1354173,I1354165,);
not I_79463 (I1354464,I895388);
nor I_79464 (I1354481,I1354464,I895382);
nor I_79465 (I1354498,I1354481,I1354303);
DFFARX1 I_79466 (I1354498,I3563,I1354173,I1354162,);
not I_79467 (I1354529,I1354481);
DFFARX1 I_79468 (I1354529,I3563,I1354173,I1354555,);
not I_79469 (I1354563,I1354555);
nor I_79470 (I1354159,I1354563,I1354481);
nor I_79471 (I1354594,I1354464,I895376);
and I_79472 (I1354611,I1354594,I895391);
or I_79473 (I1354628,I1354611,I895379);
DFFARX1 I_79474 (I1354628,I3563,I1354173,I1354654,);
not I_79475 (I1354662,I1354654);
nand I_79476 (I1354679,I1354662,I1354402);
not I_79477 (I1354153,I1354679);
nand I_79478 (I1354147,I1354679,I1354419);
nand I_79479 (I1354144,I1354662,I1354286);
not I_79480 (I1354768,I3570);
DFFARX1 I_79481 (I247013,I3563,I1354768,I1354794,);
DFFARX1 I_79482 (I247016,I3563,I1354768,I1354811,);
not I_79483 (I1354819,I1354811);
nor I_79484 (I1354736,I1354794,I1354819);
DFFARX1 I_79485 (I1354819,I3563,I1354768,I1354751,);
nor I_79486 (I1354864,I247022,I247016);
and I_79487 (I1354881,I1354864,I247019);
nor I_79488 (I1354898,I1354881,I247022);
not I_79489 (I1354915,I247022);
and I_79490 (I1354932,I1354915,I247013);
nand I_79491 (I1354949,I1354932,I247031);
nor I_79492 (I1354966,I1354915,I1354949);
DFFARX1 I_79493 (I1354966,I3563,I1354768,I1354733,);
not I_79494 (I1354997,I1354949);
nand I_79495 (I1355014,I1354819,I1354997);
nand I_79496 (I1354745,I1354881,I1354997);
DFFARX1 I_79497 (I1354915,I3563,I1354768,I1354760,);
not I_79498 (I1355059,I247025);
nor I_79499 (I1355076,I1355059,I247013);
nor I_79500 (I1355093,I1355076,I1354898);
DFFARX1 I_79501 (I1355093,I3563,I1354768,I1354757,);
not I_79502 (I1355124,I1355076);
DFFARX1 I_79503 (I1355124,I3563,I1354768,I1355150,);
not I_79504 (I1355158,I1355150);
nor I_79505 (I1354754,I1355158,I1355076);
nor I_79506 (I1355189,I1355059,I247028);
and I_79507 (I1355206,I1355189,I247034);
or I_79508 (I1355223,I1355206,I247037);
DFFARX1 I_79509 (I1355223,I3563,I1354768,I1355249,);
not I_79510 (I1355257,I1355249);
nand I_79511 (I1355274,I1355257,I1354997);
not I_79512 (I1354748,I1355274);
nand I_79513 (I1354742,I1355274,I1355014);
nand I_79514 (I1354739,I1355257,I1354881);
not I_79515 (I1355363,I3570);
DFFARX1 I_79516 (I127286,I3563,I1355363,I1355389,);
DFFARX1 I_79517 (I127274,I3563,I1355363,I1355406,);
not I_79518 (I1355414,I1355406);
nor I_79519 (I1355331,I1355389,I1355414);
DFFARX1 I_79520 (I1355414,I3563,I1355363,I1355346,);
nor I_79521 (I1355459,I127265,I127289);
and I_79522 (I1355476,I1355459,I127268);
nor I_79523 (I1355493,I1355476,I127265);
not I_79524 (I1355510,I127265);
and I_79525 (I1355527,I1355510,I127271);
nand I_79526 (I1355544,I1355527,I127283);
nor I_79527 (I1355561,I1355510,I1355544);
DFFARX1 I_79528 (I1355561,I3563,I1355363,I1355328,);
not I_79529 (I1355592,I1355544);
nand I_79530 (I1355609,I1355414,I1355592);
nand I_79531 (I1355340,I1355476,I1355592);
DFFARX1 I_79532 (I1355510,I3563,I1355363,I1355355,);
not I_79533 (I1355654,I127265);
nor I_79534 (I1355671,I1355654,I127271);
nor I_79535 (I1355688,I1355671,I1355493);
DFFARX1 I_79536 (I1355688,I3563,I1355363,I1355352,);
not I_79537 (I1355719,I1355671);
DFFARX1 I_79538 (I1355719,I3563,I1355363,I1355745,);
not I_79539 (I1355753,I1355745);
nor I_79540 (I1355349,I1355753,I1355671);
nor I_79541 (I1355784,I1355654,I127268);
and I_79542 (I1355801,I1355784,I127277);
or I_79543 (I1355818,I1355801,I127280);
DFFARX1 I_79544 (I1355818,I3563,I1355363,I1355844,);
not I_79545 (I1355852,I1355844);
nand I_79546 (I1355869,I1355852,I1355592);
not I_79547 (I1355343,I1355869);
nand I_79548 (I1355337,I1355869,I1355609);
nand I_79549 (I1355334,I1355852,I1355476);
not I_79550 (I1355958,I3570);
DFFARX1 I_79551 (I877467,I3563,I1355958,I1355984,);
DFFARX1 I_79552 (I877464,I3563,I1355958,I1356001,);
not I_79553 (I1356009,I1356001);
nor I_79554 (I1355926,I1355984,I1356009);
DFFARX1 I_79555 (I1356009,I3563,I1355958,I1355941,);
nor I_79556 (I1356054,I877479,I877461);
and I_79557 (I1356071,I1356054,I877458);
nor I_79558 (I1356088,I1356071,I877479);
not I_79559 (I1356105,I877479);
and I_79560 (I1356122,I1356105,I877464);
nand I_79561 (I1356139,I1356122,I877476);
nor I_79562 (I1356156,I1356105,I1356139);
DFFARX1 I_79563 (I1356156,I3563,I1355958,I1355923,);
not I_79564 (I1356187,I1356139);
nand I_79565 (I1356204,I1356009,I1356187);
nand I_79566 (I1355935,I1356071,I1356187);
DFFARX1 I_79567 (I1356105,I3563,I1355958,I1355950,);
not I_79568 (I1356249,I877470);
nor I_79569 (I1356266,I1356249,I877464);
nor I_79570 (I1356283,I1356266,I1356088);
DFFARX1 I_79571 (I1356283,I3563,I1355958,I1355947,);
not I_79572 (I1356314,I1356266);
DFFARX1 I_79573 (I1356314,I3563,I1355958,I1356340,);
not I_79574 (I1356348,I1356340);
nor I_79575 (I1355944,I1356348,I1356266);
nor I_79576 (I1356379,I1356249,I877458);
and I_79577 (I1356396,I1356379,I877473);
or I_79578 (I1356413,I1356396,I877461);
DFFARX1 I_79579 (I1356413,I3563,I1355958,I1356439,);
not I_79580 (I1356447,I1356439);
nand I_79581 (I1356464,I1356447,I1356187);
not I_79582 (I1355938,I1356464);
nand I_79583 (I1355932,I1356464,I1356204);
nand I_79584 (I1355929,I1356447,I1356071);
not I_79585 (I1356553,I3570);
DFFARX1 I_79586 (I1187524,I3563,I1356553,I1356579,);
DFFARX1 I_79587 (I1187536,I3563,I1356553,I1356596,);
not I_79588 (I1356604,I1356596);
nor I_79589 (I1356521,I1356579,I1356604);
DFFARX1 I_79590 (I1356604,I3563,I1356553,I1356536,);
nor I_79591 (I1356649,I1187533,I1187527);
and I_79592 (I1356666,I1356649,I1187521);
nor I_79593 (I1356683,I1356666,I1187533);
not I_79594 (I1356700,I1187533);
and I_79595 (I1356717,I1356700,I1187530);
nand I_79596 (I1356734,I1356717,I1187521);
nor I_79597 (I1356751,I1356700,I1356734);
DFFARX1 I_79598 (I1356751,I3563,I1356553,I1356518,);
not I_79599 (I1356782,I1356734);
nand I_79600 (I1356799,I1356604,I1356782);
nand I_79601 (I1356530,I1356666,I1356782);
DFFARX1 I_79602 (I1356700,I3563,I1356553,I1356545,);
not I_79603 (I1356844,I1187545);
nor I_79604 (I1356861,I1356844,I1187530);
nor I_79605 (I1356878,I1356861,I1356683);
DFFARX1 I_79606 (I1356878,I3563,I1356553,I1356542,);
not I_79607 (I1356909,I1356861);
DFFARX1 I_79608 (I1356909,I3563,I1356553,I1356935,);
not I_79609 (I1356943,I1356935);
nor I_79610 (I1356539,I1356943,I1356861);
nor I_79611 (I1356974,I1356844,I1187539);
and I_79612 (I1356991,I1356974,I1187542);
or I_79613 (I1357008,I1356991,I1187524);
DFFARX1 I_79614 (I1357008,I3563,I1356553,I1357034,);
not I_79615 (I1357042,I1357034);
nand I_79616 (I1357059,I1357042,I1356782);
not I_79617 (I1356533,I1357059);
nand I_79618 (I1356527,I1357059,I1356799);
nand I_79619 (I1356524,I1357042,I1356666);
not I_79620 (I1357148,I3570);
DFFARX1 I_79621 (I496386,I3563,I1357148,I1357174,);
DFFARX1 I_79622 (I496392,I3563,I1357148,I1357191,);
not I_79623 (I1357199,I1357191);
nor I_79624 (I1357116,I1357174,I1357199);
DFFARX1 I_79625 (I1357199,I3563,I1357148,I1357131,);
nor I_79626 (I1357244,I496401,I496386);
and I_79627 (I1357261,I1357244,I496413);
nor I_79628 (I1357278,I1357261,I496401);
not I_79629 (I1357295,I496401);
and I_79630 (I1357312,I1357295,I496389);
nand I_79631 (I1357329,I1357312,I496410);
nor I_79632 (I1357346,I1357295,I1357329);
DFFARX1 I_79633 (I1357346,I3563,I1357148,I1357113,);
not I_79634 (I1357377,I1357329);
nand I_79635 (I1357394,I1357199,I1357377);
nand I_79636 (I1357125,I1357261,I1357377);
DFFARX1 I_79637 (I1357295,I3563,I1357148,I1357140,);
not I_79638 (I1357439,I496398);
nor I_79639 (I1357456,I1357439,I496389);
nor I_79640 (I1357473,I1357456,I1357278);
DFFARX1 I_79641 (I1357473,I3563,I1357148,I1357137,);
not I_79642 (I1357504,I1357456);
DFFARX1 I_79643 (I1357504,I3563,I1357148,I1357530,);
not I_79644 (I1357538,I1357530);
nor I_79645 (I1357134,I1357538,I1357456);
nor I_79646 (I1357569,I1357439,I496395);
and I_79647 (I1357586,I1357569,I496407);
or I_79648 (I1357603,I1357586,I496404);
DFFARX1 I_79649 (I1357603,I3563,I1357148,I1357629,);
not I_79650 (I1357637,I1357629);
nand I_79651 (I1357654,I1357637,I1357377);
not I_79652 (I1357128,I1357654);
nand I_79653 (I1357122,I1357654,I1357394);
nand I_79654 (I1357119,I1357637,I1357261);
not I_79655 (I1357743,I3570);
DFFARX1 I_79656 (I569741,I3563,I1357743,I1357769,);
DFFARX1 I_79657 (I569744,I3563,I1357743,I1357786,);
not I_79658 (I1357794,I1357786);
nor I_79659 (I1357711,I1357769,I1357794);
DFFARX1 I_79660 (I1357794,I3563,I1357743,I1357726,);
nor I_79661 (I1357839,I569747,I569765);
and I_79662 (I1357856,I1357839,I569750);
nor I_79663 (I1357873,I1357856,I569747);
not I_79664 (I1357890,I569747);
and I_79665 (I1357907,I1357890,I569759);
nand I_79666 (I1357924,I1357907,I569762);
nor I_79667 (I1357941,I1357890,I1357924);
DFFARX1 I_79668 (I1357941,I3563,I1357743,I1357708,);
not I_79669 (I1357972,I1357924);
nand I_79670 (I1357989,I1357794,I1357972);
nand I_79671 (I1357720,I1357856,I1357972);
DFFARX1 I_79672 (I1357890,I3563,I1357743,I1357735,);
not I_79673 (I1358034,I569753);
nor I_79674 (I1358051,I1358034,I569759);
nor I_79675 (I1358068,I1358051,I1357873);
DFFARX1 I_79676 (I1358068,I3563,I1357743,I1357732,);
not I_79677 (I1358099,I1358051);
DFFARX1 I_79678 (I1358099,I3563,I1357743,I1358125,);
not I_79679 (I1358133,I1358125);
nor I_79680 (I1357729,I1358133,I1358051);
nor I_79681 (I1358164,I1358034,I569741);
and I_79682 (I1358181,I1358164,I569756);
or I_79683 (I1358198,I1358181,I569744);
DFFARX1 I_79684 (I1358198,I3563,I1357743,I1358224,);
not I_79685 (I1358232,I1358224);
nand I_79686 (I1358249,I1358232,I1357972);
not I_79687 (I1357723,I1358249);
nand I_79688 (I1357717,I1358249,I1357989);
nand I_79689 (I1357714,I1358232,I1357856);
not I_79690 (I1358338,I3570);
DFFARX1 I_79691 (I1224516,I3563,I1358338,I1358364,);
DFFARX1 I_79692 (I1224528,I3563,I1358338,I1358381,);
not I_79693 (I1358389,I1358381);
nor I_79694 (I1358306,I1358364,I1358389);
DFFARX1 I_79695 (I1358389,I3563,I1358338,I1358321,);
nor I_79696 (I1358434,I1224525,I1224519);
and I_79697 (I1358451,I1358434,I1224513);
nor I_79698 (I1358468,I1358451,I1224525);
not I_79699 (I1358485,I1224525);
and I_79700 (I1358502,I1358485,I1224522);
nand I_79701 (I1358519,I1358502,I1224513);
nor I_79702 (I1358536,I1358485,I1358519);
DFFARX1 I_79703 (I1358536,I3563,I1358338,I1358303,);
not I_79704 (I1358567,I1358519);
nand I_79705 (I1358584,I1358389,I1358567);
nand I_79706 (I1358315,I1358451,I1358567);
DFFARX1 I_79707 (I1358485,I3563,I1358338,I1358330,);
not I_79708 (I1358629,I1224537);
nor I_79709 (I1358646,I1358629,I1224522);
nor I_79710 (I1358663,I1358646,I1358468);
DFFARX1 I_79711 (I1358663,I3563,I1358338,I1358327,);
not I_79712 (I1358694,I1358646);
DFFARX1 I_79713 (I1358694,I3563,I1358338,I1358720,);
not I_79714 (I1358728,I1358720);
nor I_79715 (I1358324,I1358728,I1358646);
nor I_79716 (I1358759,I1358629,I1224531);
and I_79717 (I1358776,I1358759,I1224534);
or I_79718 (I1358793,I1358776,I1224516);
DFFARX1 I_79719 (I1358793,I3563,I1358338,I1358819,);
not I_79720 (I1358827,I1358819);
nand I_79721 (I1358844,I1358827,I1358567);
not I_79722 (I1358318,I1358844);
nand I_79723 (I1358312,I1358844,I1358584);
nand I_79724 (I1358309,I1358827,I1358451);
not I_79725 (I1358933,I3570);
DFFARX1 I_79726 (I434914,I3563,I1358933,I1358959,);
DFFARX1 I_79727 (I434920,I3563,I1358933,I1358976,);
not I_79728 (I1358984,I1358976);
nor I_79729 (I1358901,I1358959,I1358984);
DFFARX1 I_79730 (I1358984,I3563,I1358933,I1358916,);
nor I_79731 (I1359029,I434929,I434914);
and I_79732 (I1359046,I1359029,I434941);
nor I_79733 (I1359063,I1359046,I434929);
not I_79734 (I1359080,I434929);
and I_79735 (I1359097,I1359080,I434917);
nand I_79736 (I1359114,I1359097,I434938);
nor I_79737 (I1359131,I1359080,I1359114);
DFFARX1 I_79738 (I1359131,I3563,I1358933,I1358898,);
not I_79739 (I1359162,I1359114);
nand I_79740 (I1359179,I1358984,I1359162);
nand I_79741 (I1358910,I1359046,I1359162);
DFFARX1 I_79742 (I1359080,I3563,I1358933,I1358925,);
not I_79743 (I1359224,I434926);
nor I_79744 (I1359241,I1359224,I434917);
nor I_79745 (I1359258,I1359241,I1359063);
DFFARX1 I_79746 (I1359258,I3563,I1358933,I1358922,);
not I_79747 (I1359289,I1359241);
DFFARX1 I_79748 (I1359289,I3563,I1358933,I1359315,);
not I_79749 (I1359323,I1359315);
nor I_79750 (I1358919,I1359323,I1359241);
nor I_79751 (I1359354,I1359224,I434923);
and I_79752 (I1359371,I1359354,I434935);
or I_79753 (I1359388,I1359371,I434932);
DFFARX1 I_79754 (I1359388,I3563,I1358933,I1359414,);
not I_79755 (I1359422,I1359414);
nand I_79756 (I1359439,I1359422,I1359162);
not I_79757 (I1358913,I1359439);
nand I_79758 (I1358907,I1359439,I1359179);
nand I_79759 (I1358904,I1359422,I1359046);
not I_79760 (I1359528,I3570);
DFFARX1 I_79761 (I951703,I3563,I1359528,I1359554,);
DFFARX1 I_79762 (I951721,I3563,I1359528,I1359571,);
not I_79763 (I1359579,I1359571);
nor I_79764 (I1359496,I1359554,I1359579);
DFFARX1 I_79765 (I1359579,I3563,I1359528,I1359511,);
nor I_79766 (I1359624,I951700,I951712);
and I_79767 (I1359641,I1359624,I951697);
nor I_79768 (I1359658,I1359641,I951700);
not I_79769 (I1359675,I951700);
and I_79770 (I1359692,I1359675,I951706);
nand I_79771 (I1359709,I1359692,I951718);
nor I_79772 (I1359726,I1359675,I1359709);
DFFARX1 I_79773 (I1359726,I3563,I1359528,I1359493,);
not I_79774 (I1359757,I1359709);
nand I_79775 (I1359774,I1359579,I1359757);
nand I_79776 (I1359505,I1359641,I1359757);
DFFARX1 I_79777 (I1359675,I3563,I1359528,I1359520,);
not I_79778 (I1359819,I951709);
nor I_79779 (I1359836,I1359819,I951706);
nor I_79780 (I1359853,I1359836,I1359658);
DFFARX1 I_79781 (I1359853,I3563,I1359528,I1359517,);
not I_79782 (I1359884,I1359836);
DFFARX1 I_79783 (I1359884,I3563,I1359528,I1359910,);
not I_79784 (I1359918,I1359910);
nor I_79785 (I1359514,I1359918,I1359836);
nor I_79786 (I1359949,I1359819,I951697);
and I_79787 (I1359966,I1359949,I951724);
or I_79788 (I1359983,I1359966,I951715);
DFFARX1 I_79789 (I1359983,I3563,I1359528,I1360009,);
not I_79790 (I1360017,I1360009);
nand I_79791 (I1360034,I1360017,I1359757);
not I_79792 (I1359508,I1360034);
nand I_79793 (I1359502,I1360034,I1359774);
nand I_79794 (I1359499,I1360017,I1359641);
not I_79795 (I1360123,I3570);
DFFARX1 I_79796 (I850590,I3563,I1360123,I1360149,);
DFFARX1 I_79797 (I850587,I3563,I1360123,I1360166,);
not I_79798 (I1360174,I1360166);
nor I_79799 (I1360091,I1360149,I1360174);
DFFARX1 I_79800 (I1360174,I3563,I1360123,I1360106,);
nor I_79801 (I1360219,I850602,I850584);
and I_79802 (I1360236,I1360219,I850581);
nor I_79803 (I1360253,I1360236,I850602);
not I_79804 (I1360270,I850602);
and I_79805 (I1360287,I1360270,I850587);
nand I_79806 (I1360304,I1360287,I850599);
nor I_79807 (I1360321,I1360270,I1360304);
DFFARX1 I_79808 (I1360321,I3563,I1360123,I1360088,);
not I_79809 (I1360352,I1360304);
nand I_79810 (I1360369,I1360174,I1360352);
nand I_79811 (I1360100,I1360236,I1360352);
DFFARX1 I_79812 (I1360270,I3563,I1360123,I1360115,);
not I_79813 (I1360414,I850593);
nor I_79814 (I1360431,I1360414,I850587);
nor I_79815 (I1360448,I1360431,I1360253);
DFFARX1 I_79816 (I1360448,I3563,I1360123,I1360112,);
not I_79817 (I1360479,I1360431);
DFFARX1 I_79818 (I1360479,I3563,I1360123,I1360505,);
not I_79819 (I1360513,I1360505);
nor I_79820 (I1360109,I1360513,I1360431);
nor I_79821 (I1360544,I1360414,I850581);
and I_79822 (I1360561,I1360544,I850596);
or I_79823 (I1360578,I1360561,I850584);
DFFARX1 I_79824 (I1360578,I3563,I1360123,I1360604,);
not I_79825 (I1360612,I1360604);
nand I_79826 (I1360629,I1360612,I1360352);
not I_79827 (I1360103,I1360629);
nand I_79828 (I1360097,I1360629,I1360369);
nand I_79829 (I1360094,I1360612,I1360236);
not I_79830 (I1360718,I3570);
DFFARX1 I_79831 (I482242,I3563,I1360718,I1360744,);
DFFARX1 I_79832 (I482248,I3563,I1360718,I1360761,);
not I_79833 (I1360769,I1360761);
nor I_79834 (I1360686,I1360744,I1360769);
DFFARX1 I_79835 (I1360769,I3563,I1360718,I1360701,);
nor I_79836 (I1360814,I482257,I482242);
and I_79837 (I1360831,I1360814,I482269);
nor I_79838 (I1360848,I1360831,I482257);
not I_79839 (I1360865,I482257);
and I_79840 (I1360882,I1360865,I482245);
nand I_79841 (I1360899,I1360882,I482266);
nor I_79842 (I1360916,I1360865,I1360899);
DFFARX1 I_79843 (I1360916,I3563,I1360718,I1360683,);
not I_79844 (I1360947,I1360899);
nand I_79845 (I1360964,I1360769,I1360947);
nand I_79846 (I1360695,I1360831,I1360947);
DFFARX1 I_79847 (I1360865,I3563,I1360718,I1360710,);
not I_79848 (I1361009,I482254);
nor I_79849 (I1361026,I1361009,I482245);
nor I_79850 (I1361043,I1361026,I1360848);
DFFARX1 I_79851 (I1361043,I3563,I1360718,I1360707,);
not I_79852 (I1361074,I1361026);
DFFARX1 I_79853 (I1361074,I3563,I1360718,I1361100,);
not I_79854 (I1361108,I1361100);
nor I_79855 (I1360704,I1361108,I1361026);
nor I_79856 (I1361139,I1361009,I482251);
and I_79857 (I1361156,I1361139,I482263);
or I_79858 (I1361173,I1361156,I482260);
DFFARX1 I_79859 (I1361173,I3563,I1360718,I1361199,);
not I_79860 (I1361207,I1361199);
nand I_79861 (I1361224,I1361207,I1360947);
not I_79862 (I1360698,I1361224);
nand I_79863 (I1360692,I1361224,I1360964);
nand I_79864 (I1360689,I1361207,I1360831);
not I_79865 (I1361313,I3570);
DFFARX1 I_79866 (I293818,I3563,I1361313,I1361339,);
DFFARX1 I_79867 (I293812,I3563,I1361313,I1361356,);
not I_79868 (I1361364,I1361356);
nor I_79869 (I1361281,I1361339,I1361364);
DFFARX1 I_79870 (I1361364,I3563,I1361313,I1361296,);
nor I_79871 (I1361409,I293800,I293821);
and I_79872 (I1361426,I1361409,I293815);
nor I_79873 (I1361443,I1361426,I293800);
not I_79874 (I1361460,I293800);
and I_79875 (I1361477,I1361460,I293797);
nand I_79876 (I1361494,I1361477,I293809);
nor I_79877 (I1361511,I1361460,I1361494);
DFFARX1 I_79878 (I1361511,I3563,I1361313,I1361278,);
not I_79879 (I1361542,I1361494);
nand I_79880 (I1361559,I1361364,I1361542);
nand I_79881 (I1361290,I1361426,I1361542);
DFFARX1 I_79882 (I1361460,I3563,I1361313,I1361305,);
not I_79883 (I1361604,I293824);
nor I_79884 (I1361621,I1361604,I293797);
nor I_79885 (I1361638,I1361621,I1361443);
DFFARX1 I_79886 (I1361638,I3563,I1361313,I1361302,);
not I_79887 (I1361669,I1361621);
DFFARX1 I_79888 (I1361669,I3563,I1361313,I1361695,);
not I_79889 (I1361703,I1361695);
nor I_79890 (I1361299,I1361703,I1361621);
nor I_79891 (I1361734,I1361604,I293806);
and I_79892 (I1361751,I1361734,I293803);
or I_79893 (I1361768,I1361751,I293797);
DFFARX1 I_79894 (I1361768,I3563,I1361313,I1361794,);
not I_79895 (I1361802,I1361794);
nand I_79896 (I1361819,I1361802,I1361542);
not I_79897 (I1361293,I1361819);
nand I_79898 (I1361287,I1361819,I1361559);
nand I_79899 (I1361284,I1361802,I1361426);
not I_79900 (I1361908,I3570);
DFFARX1 I_79901 (I1059574,I3563,I1361908,I1361934,);
DFFARX1 I_79902 (I1059565,I3563,I1361908,I1361951,);
not I_79903 (I1361959,I1361951);
nor I_79904 (I1361876,I1361934,I1361959);
DFFARX1 I_79905 (I1361959,I3563,I1361908,I1361891,);
nor I_79906 (I1362004,I1059571,I1059580);
and I_79907 (I1362021,I1362004,I1059583);
nor I_79908 (I1362038,I1362021,I1059571);
not I_79909 (I1362055,I1059571);
and I_79910 (I1362072,I1362055,I1059562);
nand I_79911 (I1362089,I1362072,I1059568);
nor I_79912 (I1362106,I1362055,I1362089);
DFFARX1 I_79913 (I1362106,I3563,I1361908,I1361873,);
not I_79914 (I1362137,I1362089);
nand I_79915 (I1362154,I1361959,I1362137);
nand I_79916 (I1361885,I1362021,I1362137);
DFFARX1 I_79917 (I1362055,I3563,I1361908,I1361900,);
not I_79918 (I1362199,I1059577);
nor I_79919 (I1362216,I1362199,I1059562);
nor I_79920 (I1362233,I1362216,I1362038);
DFFARX1 I_79921 (I1362233,I3563,I1361908,I1361897,);
not I_79922 (I1362264,I1362216);
DFFARX1 I_79923 (I1362264,I3563,I1361908,I1362290,);
not I_79924 (I1362298,I1362290);
nor I_79925 (I1361894,I1362298,I1362216);
nor I_79926 (I1362329,I1362199,I1059562);
and I_79927 (I1362346,I1362329,I1059565);
or I_79928 (I1362363,I1362346,I1059568);
DFFARX1 I_79929 (I1362363,I3563,I1361908,I1362389,);
not I_79930 (I1362397,I1362389);
nand I_79931 (I1362414,I1362397,I1362137);
not I_79932 (I1361888,I1362414);
nand I_79933 (I1361882,I1362414,I1362154);
nand I_79934 (I1361879,I1362397,I1362021);
not I_79935 (I1362503,I3570);
DFFARX1 I_79936 (I499650,I3563,I1362503,I1362529,);
DFFARX1 I_79937 (I499656,I3563,I1362503,I1362546,);
not I_79938 (I1362554,I1362546);
nor I_79939 (I1362471,I1362529,I1362554);
DFFARX1 I_79940 (I1362554,I3563,I1362503,I1362486,);
nor I_79941 (I1362599,I499665,I499650);
and I_79942 (I1362616,I1362599,I499677);
nor I_79943 (I1362633,I1362616,I499665);
not I_79944 (I1362650,I499665);
and I_79945 (I1362667,I1362650,I499653);
nand I_79946 (I1362684,I1362667,I499674);
nor I_79947 (I1362701,I1362650,I1362684);
DFFARX1 I_79948 (I1362701,I3563,I1362503,I1362468,);
not I_79949 (I1362732,I1362684);
nand I_79950 (I1362749,I1362554,I1362732);
nand I_79951 (I1362480,I1362616,I1362732);
DFFARX1 I_79952 (I1362650,I3563,I1362503,I1362495,);
not I_79953 (I1362794,I499662);
nor I_79954 (I1362811,I1362794,I499653);
nor I_79955 (I1362828,I1362811,I1362633);
DFFARX1 I_79956 (I1362828,I3563,I1362503,I1362492,);
not I_79957 (I1362859,I1362811);
DFFARX1 I_79958 (I1362859,I3563,I1362503,I1362885,);
not I_79959 (I1362893,I1362885);
nor I_79960 (I1362489,I1362893,I1362811);
nor I_79961 (I1362924,I1362794,I499659);
and I_79962 (I1362941,I1362924,I499671);
or I_79963 (I1362958,I1362941,I499668);
DFFARX1 I_79964 (I1362958,I3563,I1362503,I1362984,);
not I_79965 (I1362992,I1362984);
nand I_79966 (I1363009,I1362992,I1362732);
not I_79967 (I1362483,I1363009);
nand I_79968 (I1362477,I1363009,I1362749);
nand I_79969 (I1362474,I1362992,I1362616);
not I_79970 (I1363098,I3570);
DFFARX1 I_79971 (I505090,I3563,I1363098,I1363124,);
DFFARX1 I_79972 (I505096,I3563,I1363098,I1363141,);
not I_79973 (I1363149,I1363141);
nor I_79974 (I1363066,I1363124,I1363149);
DFFARX1 I_79975 (I1363149,I3563,I1363098,I1363081,);
nor I_79976 (I1363194,I505105,I505090);
and I_79977 (I1363211,I1363194,I505117);
nor I_79978 (I1363228,I1363211,I505105);
not I_79979 (I1363245,I505105);
and I_79980 (I1363262,I1363245,I505093);
nand I_79981 (I1363279,I1363262,I505114);
nor I_79982 (I1363296,I1363245,I1363279);
DFFARX1 I_79983 (I1363296,I3563,I1363098,I1363063,);
not I_79984 (I1363327,I1363279);
nand I_79985 (I1363344,I1363149,I1363327);
nand I_79986 (I1363075,I1363211,I1363327);
DFFARX1 I_79987 (I1363245,I3563,I1363098,I1363090,);
not I_79988 (I1363389,I505102);
nor I_79989 (I1363406,I1363389,I505093);
nor I_79990 (I1363423,I1363406,I1363228);
DFFARX1 I_79991 (I1363423,I3563,I1363098,I1363087,);
not I_79992 (I1363454,I1363406);
DFFARX1 I_79993 (I1363454,I3563,I1363098,I1363480,);
not I_79994 (I1363488,I1363480);
nor I_79995 (I1363084,I1363488,I1363406);
nor I_79996 (I1363519,I1363389,I505099);
and I_79997 (I1363536,I1363519,I505111);
or I_79998 (I1363553,I1363536,I505108);
DFFARX1 I_79999 (I1363553,I3563,I1363098,I1363579,);
not I_80000 (I1363587,I1363579);
nand I_80001 (I1363604,I1363587,I1363327);
not I_80002 (I1363078,I1363604);
nand I_80003 (I1363072,I1363604,I1363344);
nand I_80004 (I1363069,I1363587,I1363211);
not I_80005 (I1363693,I3570);
DFFARX1 I_80006 (I112003,I3563,I1363693,I1363719,);
DFFARX1 I_80007 (I111991,I3563,I1363693,I1363736,);
not I_80008 (I1363744,I1363736);
nor I_80009 (I1363661,I1363719,I1363744);
DFFARX1 I_80010 (I1363744,I3563,I1363693,I1363676,);
nor I_80011 (I1363789,I111982,I112006);
and I_80012 (I1363806,I1363789,I111985);
nor I_80013 (I1363823,I1363806,I111982);
not I_80014 (I1363840,I111982);
and I_80015 (I1363857,I1363840,I111988);
nand I_80016 (I1363874,I1363857,I112000);
nor I_80017 (I1363891,I1363840,I1363874);
DFFARX1 I_80018 (I1363891,I3563,I1363693,I1363658,);
not I_80019 (I1363922,I1363874);
nand I_80020 (I1363939,I1363744,I1363922);
nand I_80021 (I1363670,I1363806,I1363922);
DFFARX1 I_80022 (I1363840,I3563,I1363693,I1363685,);
not I_80023 (I1363984,I111982);
nor I_80024 (I1364001,I1363984,I111988);
nor I_80025 (I1364018,I1364001,I1363823);
DFFARX1 I_80026 (I1364018,I3563,I1363693,I1363682,);
not I_80027 (I1364049,I1364001);
DFFARX1 I_80028 (I1364049,I3563,I1363693,I1364075,);
not I_80029 (I1364083,I1364075);
nor I_80030 (I1363679,I1364083,I1364001);
nor I_80031 (I1364114,I1363984,I111985);
and I_80032 (I1364131,I1364114,I111994);
or I_80033 (I1364148,I1364131,I111997);
DFFARX1 I_80034 (I1364148,I3563,I1363693,I1364174,);
not I_80035 (I1364182,I1364174);
nand I_80036 (I1364199,I1364182,I1363922);
not I_80037 (I1363673,I1364199);
nand I_80038 (I1363667,I1364199,I1363939);
nand I_80039 (I1363664,I1364182,I1363806);
not I_80040 (I1364288,I3570);
DFFARX1 I_80041 (I470274,I3563,I1364288,I1364314,);
DFFARX1 I_80042 (I470280,I3563,I1364288,I1364331,);
not I_80043 (I1364339,I1364331);
nor I_80044 (I1364256,I1364314,I1364339);
DFFARX1 I_80045 (I1364339,I3563,I1364288,I1364271,);
nor I_80046 (I1364384,I470289,I470274);
and I_80047 (I1364401,I1364384,I470301);
nor I_80048 (I1364418,I1364401,I470289);
not I_80049 (I1364435,I470289);
and I_80050 (I1364452,I1364435,I470277);
nand I_80051 (I1364469,I1364452,I470298);
nor I_80052 (I1364486,I1364435,I1364469);
DFFARX1 I_80053 (I1364486,I3563,I1364288,I1364253,);
not I_80054 (I1364517,I1364469);
nand I_80055 (I1364534,I1364339,I1364517);
nand I_80056 (I1364265,I1364401,I1364517);
DFFARX1 I_80057 (I1364435,I3563,I1364288,I1364280,);
not I_80058 (I1364579,I470286);
nor I_80059 (I1364596,I1364579,I470277);
nor I_80060 (I1364613,I1364596,I1364418);
DFFARX1 I_80061 (I1364613,I3563,I1364288,I1364277,);
not I_80062 (I1364644,I1364596);
DFFARX1 I_80063 (I1364644,I3563,I1364288,I1364670,);
not I_80064 (I1364678,I1364670);
nor I_80065 (I1364274,I1364678,I1364596);
nor I_80066 (I1364709,I1364579,I470283);
and I_80067 (I1364726,I1364709,I470295);
or I_80068 (I1364743,I1364726,I470292);
DFFARX1 I_80069 (I1364743,I3563,I1364288,I1364769,);
not I_80070 (I1364777,I1364769);
nand I_80071 (I1364794,I1364777,I1364517);
not I_80072 (I1364268,I1364794);
nand I_80073 (I1364262,I1364794,I1364534);
nand I_80074 (I1364259,I1364777,I1364401);
not I_80075 (I1364883,I3570);
DFFARX1 I_80076 (I869562,I3563,I1364883,I1364909,);
DFFARX1 I_80077 (I869559,I3563,I1364883,I1364926,);
not I_80078 (I1364934,I1364926);
nor I_80079 (I1364851,I1364909,I1364934);
DFFARX1 I_80080 (I1364934,I3563,I1364883,I1364866,);
nor I_80081 (I1364979,I869574,I869556);
and I_80082 (I1364996,I1364979,I869553);
nor I_80083 (I1365013,I1364996,I869574);
not I_80084 (I1365030,I869574);
and I_80085 (I1365047,I1365030,I869559);
nand I_80086 (I1365064,I1365047,I869571);
nor I_80087 (I1365081,I1365030,I1365064);
DFFARX1 I_80088 (I1365081,I3563,I1364883,I1364848,);
not I_80089 (I1365112,I1365064);
nand I_80090 (I1365129,I1364934,I1365112);
nand I_80091 (I1364860,I1364996,I1365112);
DFFARX1 I_80092 (I1365030,I3563,I1364883,I1364875,);
not I_80093 (I1365174,I869565);
nor I_80094 (I1365191,I1365174,I869559);
nor I_80095 (I1365208,I1365191,I1365013);
DFFARX1 I_80096 (I1365208,I3563,I1364883,I1364872,);
not I_80097 (I1365239,I1365191);
DFFARX1 I_80098 (I1365239,I3563,I1364883,I1365265,);
not I_80099 (I1365273,I1365265);
nor I_80100 (I1364869,I1365273,I1365191);
nor I_80101 (I1365304,I1365174,I869553);
and I_80102 (I1365321,I1365304,I869568);
or I_80103 (I1365338,I1365321,I869556);
DFFARX1 I_80104 (I1365338,I3563,I1364883,I1365364,);
not I_80105 (I1365372,I1365364);
nand I_80106 (I1365389,I1365372,I1365112);
not I_80107 (I1364863,I1365389);
nand I_80108 (I1364857,I1365389,I1365129);
nand I_80109 (I1364854,I1365372,I1364996);
not I_80110 (I1365478,I3570);
DFFARX1 I_80111 (I302777,I3563,I1365478,I1365504,);
DFFARX1 I_80112 (I302771,I3563,I1365478,I1365521,);
not I_80113 (I1365529,I1365521);
nor I_80114 (I1365446,I1365504,I1365529);
DFFARX1 I_80115 (I1365529,I3563,I1365478,I1365461,);
nor I_80116 (I1365574,I302759,I302780);
and I_80117 (I1365591,I1365574,I302774);
nor I_80118 (I1365608,I1365591,I302759);
not I_80119 (I1365625,I302759);
and I_80120 (I1365642,I1365625,I302756);
nand I_80121 (I1365659,I1365642,I302768);
nor I_80122 (I1365676,I1365625,I1365659);
DFFARX1 I_80123 (I1365676,I3563,I1365478,I1365443,);
not I_80124 (I1365707,I1365659);
nand I_80125 (I1365724,I1365529,I1365707);
nand I_80126 (I1365455,I1365591,I1365707);
DFFARX1 I_80127 (I1365625,I3563,I1365478,I1365470,);
not I_80128 (I1365769,I302783);
nor I_80129 (I1365786,I1365769,I302756);
nor I_80130 (I1365803,I1365786,I1365608);
DFFARX1 I_80131 (I1365803,I3563,I1365478,I1365467,);
not I_80132 (I1365834,I1365786);
DFFARX1 I_80133 (I1365834,I3563,I1365478,I1365860,);
not I_80134 (I1365868,I1365860);
nor I_80135 (I1365464,I1365868,I1365786);
nor I_80136 (I1365899,I1365769,I302765);
and I_80137 (I1365916,I1365899,I302762);
or I_80138 (I1365933,I1365916,I302756);
DFFARX1 I_80139 (I1365933,I3563,I1365478,I1365959,);
not I_80140 (I1365967,I1365959);
nand I_80141 (I1365984,I1365967,I1365707);
not I_80142 (I1365458,I1365984);
nand I_80143 (I1365452,I1365984,I1365724);
nand I_80144 (I1365449,I1365967,I1365591);
not I_80145 (I1366073,I3570);
DFFARX1 I_80146 (I1296441,I3563,I1366073,I1366099,);
DFFARX1 I_80147 (I1296432,I3563,I1366073,I1366116,);
not I_80148 (I1366124,I1366116);
nor I_80149 (I1366041,I1366099,I1366124);
DFFARX1 I_80150 (I1366124,I3563,I1366073,I1366056,);
nor I_80151 (I1366169,I1296423,I1296438);
and I_80152 (I1366186,I1366169,I1296426);
nor I_80153 (I1366203,I1366186,I1296423);
not I_80154 (I1366220,I1296423);
and I_80155 (I1366237,I1366220,I1296429);
nand I_80156 (I1366254,I1366237,I1296447);
nor I_80157 (I1366271,I1366220,I1366254);
DFFARX1 I_80158 (I1366271,I3563,I1366073,I1366038,);
not I_80159 (I1366302,I1366254);
nand I_80160 (I1366319,I1366124,I1366302);
nand I_80161 (I1366050,I1366186,I1366302);
DFFARX1 I_80162 (I1366220,I3563,I1366073,I1366065,);
not I_80163 (I1366364,I1296423);
nor I_80164 (I1366381,I1366364,I1296429);
nor I_80165 (I1366398,I1366381,I1366203);
DFFARX1 I_80166 (I1366398,I3563,I1366073,I1366062,);
not I_80167 (I1366429,I1366381);
DFFARX1 I_80168 (I1366429,I3563,I1366073,I1366455,);
not I_80169 (I1366463,I1366455);
nor I_80170 (I1366059,I1366463,I1366381);
nor I_80171 (I1366494,I1366364,I1296426);
and I_80172 (I1366511,I1366494,I1296435);
or I_80173 (I1366528,I1366511,I1296444);
DFFARX1 I_80174 (I1366528,I3563,I1366073,I1366554,);
not I_80175 (I1366562,I1366554);
nand I_80176 (I1366579,I1366562,I1366302);
not I_80177 (I1366053,I1366579);
nand I_80178 (I1366047,I1366579,I1366319);
nand I_80179 (I1366044,I1366562,I1366186);
not I_80180 (I1366668,I3570);
DFFARX1 I_80181 (I1037621,I3563,I1366668,I1366694,);
DFFARX1 I_80182 (I1037639,I3563,I1366668,I1366711,);
not I_80183 (I1366719,I1366711);
nor I_80184 (I1366636,I1366694,I1366719);
DFFARX1 I_80185 (I1366719,I3563,I1366668,I1366651,);
nor I_80186 (I1366764,I1037618,I1037630);
and I_80187 (I1366781,I1366764,I1037615);
nor I_80188 (I1366798,I1366781,I1037618);
not I_80189 (I1366815,I1037618);
and I_80190 (I1366832,I1366815,I1037624);
nand I_80191 (I1366849,I1366832,I1037636);
nor I_80192 (I1366866,I1366815,I1366849);
DFFARX1 I_80193 (I1366866,I3563,I1366668,I1366633,);
not I_80194 (I1366897,I1366849);
nand I_80195 (I1366914,I1366719,I1366897);
nand I_80196 (I1366645,I1366781,I1366897);
DFFARX1 I_80197 (I1366815,I3563,I1366668,I1366660,);
not I_80198 (I1366959,I1037627);
nor I_80199 (I1366976,I1366959,I1037624);
nor I_80200 (I1366993,I1366976,I1366798);
DFFARX1 I_80201 (I1366993,I3563,I1366668,I1366657,);
not I_80202 (I1367024,I1366976);
DFFARX1 I_80203 (I1367024,I3563,I1366668,I1367050,);
not I_80204 (I1367058,I1367050);
nor I_80205 (I1366654,I1367058,I1366976);
nor I_80206 (I1367089,I1366959,I1037615);
and I_80207 (I1367106,I1367089,I1037642);
or I_80208 (I1367123,I1367106,I1037633);
DFFARX1 I_80209 (I1367123,I3563,I1366668,I1367149,);
not I_80210 (I1367157,I1367149);
nand I_80211 (I1367174,I1367157,I1366897);
not I_80212 (I1366648,I1367174);
nand I_80213 (I1366642,I1367174,I1366914);
nand I_80214 (I1366639,I1367157,I1366781);
not I_80215 (I1367263,I3570);
DFFARX1 I_80216 (I893277,I3563,I1367263,I1367289,);
DFFARX1 I_80217 (I893274,I3563,I1367263,I1367306,);
not I_80218 (I1367314,I1367306);
nor I_80219 (I1367231,I1367289,I1367314);
DFFARX1 I_80220 (I1367314,I3563,I1367263,I1367246,);
nor I_80221 (I1367359,I893289,I893271);
and I_80222 (I1367376,I1367359,I893268);
nor I_80223 (I1367393,I1367376,I893289);
not I_80224 (I1367410,I893289);
and I_80225 (I1367427,I1367410,I893274);
nand I_80226 (I1367444,I1367427,I893286);
nor I_80227 (I1367461,I1367410,I1367444);
DFFARX1 I_80228 (I1367461,I3563,I1367263,I1367228,);
not I_80229 (I1367492,I1367444);
nand I_80230 (I1367509,I1367314,I1367492);
nand I_80231 (I1367240,I1367376,I1367492);
DFFARX1 I_80232 (I1367410,I3563,I1367263,I1367255,);
not I_80233 (I1367554,I893280);
nor I_80234 (I1367571,I1367554,I893274);
nor I_80235 (I1367588,I1367571,I1367393);
DFFARX1 I_80236 (I1367588,I3563,I1367263,I1367252,);
not I_80237 (I1367619,I1367571);
DFFARX1 I_80238 (I1367619,I3563,I1367263,I1367645,);
not I_80239 (I1367653,I1367645);
nor I_80240 (I1367249,I1367653,I1367571);
nor I_80241 (I1367684,I1367554,I893268);
and I_80242 (I1367701,I1367684,I893283);
or I_80243 (I1367718,I1367701,I893271);
DFFARX1 I_80244 (I1367718,I3563,I1367263,I1367744,);
not I_80245 (I1367752,I1367744);
nand I_80246 (I1367769,I1367752,I1367492);
not I_80247 (I1367243,I1367769);
nand I_80248 (I1367237,I1367769,I1367509);
nand I_80249 (I1367234,I1367752,I1367376);
not I_80250 (I1367858,I3570);
DFFARX1 I_80251 (I1041497,I3563,I1367858,I1367884,);
DFFARX1 I_80252 (I1041515,I3563,I1367858,I1367901,);
not I_80253 (I1367909,I1367901);
nor I_80254 (I1367826,I1367884,I1367909);
DFFARX1 I_80255 (I1367909,I3563,I1367858,I1367841,);
nor I_80256 (I1367954,I1041494,I1041506);
and I_80257 (I1367971,I1367954,I1041491);
nor I_80258 (I1367988,I1367971,I1041494);
not I_80259 (I1368005,I1041494);
and I_80260 (I1368022,I1368005,I1041500);
nand I_80261 (I1368039,I1368022,I1041512);
nor I_80262 (I1368056,I1368005,I1368039);
DFFARX1 I_80263 (I1368056,I3563,I1367858,I1367823,);
not I_80264 (I1368087,I1368039);
nand I_80265 (I1368104,I1367909,I1368087);
nand I_80266 (I1367835,I1367971,I1368087);
DFFARX1 I_80267 (I1368005,I3563,I1367858,I1367850,);
not I_80268 (I1368149,I1041503);
nor I_80269 (I1368166,I1368149,I1041500);
nor I_80270 (I1368183,I1368166,I1367988);
DFFARX1 I_80271 (I1368183,I3563,I1367858,I1367847,);
not I_80272 (I1368214,I1368166);
DFFARX1 I_80273 (I1368214,I3563,I1367858,I1368240,);
not I_80274 (I1368248,I1368240);
nor I_80275 (I1367844,I1368248,I1368166);
nor I_80276 (I1368279,I1368149,I1041491);
and I_80277 (I1368296,I1368279,I1041518);
or I_80278 (I1368313,I1368296,I1041509);
DFFARX1 I_80279 (I1368313,I3563,I1367858,I1368339,);
not I_80280 (I1368347,I1368339);
nand I_80281 (I1368364,I1368347,I1368087);
not I_80282 (I1367838,I1368364);
nand I_80283 (I1367832,I1368364,I1368104);
nand I_80284 (I1367829,I1368347,I1367971);
not I_80285 (I1368453,I3570);
DFFARX1 I_80286 (I559626,I3563,I1368453,I1368479,);
DFFARX1 I_80287 (I559629,I3563,I1368453,I1368496,);
not I_80288 (I1368504,I1368496);
nor I_80289 (I1368421,I1368479,I1368504);
DFFARX1 I_80290 (I1368504,I3563,I1368453,I1368436,);
nor I_80291 (I1368549,I559632,I559650);
and I_80292 (I1368566,I1368549,I559635);
nor I_80293 (I1368583,I1368566,I559632);
not I_80294 (I1368600,I559632);
and I_80295 (I1368617,I1368600,I559644);
nand I_80296 (I1368634,I1368617,I559647);
nor I_80297 (I1368651,I1368600,I1368634);
DFFARX1 I_80298 (I1368651,I3563,I1368453,I1368418,);
not I_80299 (I1368682,I1368634);
nand I_80300 (I1368699,I1368504,I1368682);
nand I_80301 (I1368430,I1368566,I1368682);
DFFARX1 I_80302 (I1368600,I3563,I1368453,I1368445,);
not I_80303 (I1368744,I559638);
nor I_80304 (I1368761,I1368744,I559644);
nor I_80305 (I1368778,I1368761,I1368583);
DFFARX1 I_80306 (I1368778,I3563,I1368453,I1368442,);
not I_80307 (I1368809,I1368761);
DFFARX1 I_80308 (I1368809,I3563,I1368453,I1368835,);
not I_80309 (I1368843,I1368835);
nor I_80310 (I1368439,I1368843,I1368761);
nor I_80311 (I1368874,I1368744,I559626);
and I_80312 (I1368891,I1368874,I559641);
or I_80313 (I1368908,I1368891,I559629);
DFFARX1 I_80314 (I1368908,I3563,I1368453,I1368934,);
not I_80315 (I1368942,I1368934);
nand I_80316 (I1368959,I1368942,I1368682);
not I_80317 (I1368433,I1368959);
nand I_80318 (I1368427,I1368959,I1368699);
nand I_80319 (I1368424,I1368942,I1368566);
not I_80320 (I1369048,I3570);
DFFARX1 I_80321 (I619708,I3563,I1369048,I1369074,);
DFFARX1 I_80322 (I619702,I3563,I1369048,I1369091,);
not I_80323 (I1369099,I1369091);
nor I_80324 (I1369016,I1369074,I1369099);
DFFARX1 I_80325 (I1369099,I3563,I1369048,I1369031,);
nor I_80326 (I1369144,I619699,I619690);
and I_80327 (I1369161,I1369144,I619687);
nor I_80328 (I1369178,I1369161,I619699);
not I_80329 (I1369195,I619699);
and I_80330 (I1369212,I1369195,I619693);
nand I_80331 (I1369229,I1369212,I619705);
nor I_80332 (I1369246,I1369195,I1369229);
DFFARX1 I_80333 (I1369246,I3563,I1369048,I1369013,);
not I_80334 (I1369277,I1369229);
nand I_80335 (I1369294,I1369099,I1369277);
nand I_80336 (I1369025,I1369161,I1369277);
DFFARX1 I_80337 (I1369195,I3563,I1369048,I1369040,);
not I_80338 (I1369339,I619711);
nor I_80339 (I1369356,I1369339,I619693);
nor I_80340 (I1369373,I1369356,I1369178);
DFFARX1 I_80341 (I1369373,I3563,I1369048,I1369037,);
not I_80342 (I1369404,I1369356);
DFFARX1 I_80343 (I1369404,I3563,I1369048,I1369430,);
not I_80344 (I1369438,I1369430);
nor I_80345 (I1369034,I1369438,I1369356);
nor I_80346 (I1369469,I1369339,I619690);
and I_80347 (I1369486,I1369469,I619696);
or I_80348 (I1369503,I1369486,I619687);
DFFARX1 I_80349 (I1369503,I3563,I1369048,I1369529,);
not I_80350 (I1369537,I1369529);
nand I_80351 (I1369554,I1369537,I1369277);
not I_80352 (I1369028,I1369554);
nand I_80353 (I1369022,I1369554,I1369294);
nand I_80354 (I1369019,I1369537,I1369161);
not I_80355 (I1369643,I3570);
DFFARX1 I_80356 (I712188,I3563,I1369643,I1369669,);
DFFARX1 I_80357 (I712170,I3563,I1369643,I1369686,);
not I_80358 (I1369694,I1369686);
nor I_80359 (I1369611,I1369669,I1369694);
DFFARX1 I_80360 (I1369694,I3563,I1369643,I1369626,);
nor I_80361 (I1369739,I712176,I712179);
and I_80362 (I1369756,I1369739,I712167);
nor I_80363 (I1369773,I1369756,I712176);
not I_80364 (I1369790,I712176);
and I_80365 (I1369807,I1369790,I712185);
nand I_80366 (I1369824,I1369807,I712173);
nor I_80367 (I1369841,I1369790,I1369824);
DFFARX1 I_80368 (I1369841,I3563,I1369643,I1369608,);
not I_80369 (I1369872,I1369824);
nand I_80370 (I1369889,I1369694,I1369872);
nand I_80371 (I1369620,I1369756,I1369872);
DFFARX1 I_80372 (I1369790,I3563,I1369643,I1369635,);
not I_80373 (I1369934,I712170);
nor I_80374 (I1369951,I1369934,I712185);
nor I_80375 (I1369968,I1369951,I1369773);
DFFARX1 I_80376 (I1369968,I3563,I1369643,I1369632,);
not I_80377 (I1369999,I1369951);
DFFARX1 I_80378 (I1369999,I3563,I1369643,I1370025,);
not I_80379 (I1370033,I1370025);
nor I_80380 (I1369629,I1370033,I1369951);
nor I_80381 (I1370064,I1369934,I712182);
and I_80382 (I1370081,I1370064,I712191);
or I_80383 (I1370098,I1370081,I712167);
DFFARX1 I_80384 (I1370098,I3563,I1369643,I1370124,);
not I_80385 (I1370132,I1370124);
nand I_80386 (I1370149,I1370132,I1369872);
not I_80387 (I1369623,I1370149);
nand I_80388 (I1369617,I1370149,I1369889);
nand I_80389 (I1369614,I1370132,I1369756);
not I_80390 (I1370238,I3570);
DFFARX1 I_80391 (I941367,I3563,I1370238,I1370264,);
DFFARX1 I_80392 (I941385,I3563,I1370238,I1370281,);
not I_80393 (I1370289,I1370281);
nor I_80394 (I1370206,I1370264,I1370289);
DFFARX1 I_80395 (I1370289,I3563,I1370238,I1370221,);
nor I_80396 (I1370334,I941364,I941376);
and I_80397 (I1370351,I1370334,I941361);
nor I_80398 (I1370368,I1370351,I941364);
not I_80399 (I1370385,I941364);
and I_80400 (I1370402,I1370385,I941370);
nand I_80401 (I1370419,I1370402,I941382);
nor I_80402 (I1370436,I1370385,I1370419);
DFFARX1 I_80403 (I1370436,I3563,I1370238,I1370203,);
not I_80404 (I1370467,I1370419);
nand I_80405 (I1370484,I1370289,I1370467);
nand I_80406 (I1370215,I1370351,I1370467);
DFFARX1 I_80407 (I1370385,I3563,I1370238,I1370230,);
not I_80408 (I1370529,I941373);
nor I_80409 (I1370546,I1370529,I941370);
nor I_80410 (I1370563,I1370546,I1370368);
DFFARX1 I_80411 (I1370563,I3563,I1370238,I1370227,);
not I_80412 (I1370594,I1370546);
DFFARX1 I_80413 (I1370594,I3563,I1370238,I1370620,);
not I_80414 (I1370628,I1370620);
nor I_80415 (I1370224,I1370628,I1370546);
nor I_80416 (I1370659,I1370529,I941361);
and I_80417 (I1370676,I1370659,I941388);
or I_80418 (I1370693,I1370676,I941379);
DFFARX1 I_80419 (I1370693,I3563,I1370238,I1370719,);
not I_80420 (I1370727,I1370719);
nand I_80421 (I1370744,I1370727,I1370467);
not I_80422 (I1370218,I1370744);
nand I_80423 (I1370212,I1370744,I1370484);
nand I_80424 (I1370209,I1370727,I1370351);
not I_80425 (I1370833,I3570);
DFFARX1 I_80426 (I1272521,I3563,I1370833,I1370859,);
DFFARX1 I_80427 (I1272524,I3563,I1370833,I1370876,);
not I_80428 (I1370884,I1370876);
nor I_80429 (I1370801,I1370859,I1370884);
DFFARX1 I_80430 (I1370884,I3563,I1370833,I1370816,);
nor I_80431 (I1370929,I1272524,I1272539);
and I_80432 (I1370946,I1370929,I1272533);
nor I_80433 (I1370963,I1370946,I1272524);
not I_80434 (I1370980,I1272524);
and I_80435 (I1370997,I1370980,I1272542);
nand I_80436 (I1371014,I1370997,I1272530);
nor I_80437 (I1371031,I1370980,I1371014);
DFFARX1 I_80438 (I1371031,I3563,I1370833,I1370798,);
not I_80439 (I1371062,I1371014);
nand I_80440 (I1371079,I1370884,I1371062);
nand I_80441 (I1370810,I1370946,I1371062);
DFFARX1 I_80442 (I1370980,I3563,I1370833,I1370825,);
not I_80443 (I1371124,I1272536);
nor I_80444 (I1371141,I1371124,I1272542);
nor I_80445 (I1371158,I1371141,I1370963);
DFFARX1 I_80446 (I1371158,I3563,I1370833,I1370822,);
not I_80447 (I1371189,I1371141);
DFFARX1 I_80448 (I1371189,I3563,I1370833,I1371215,);
not I_80449 (I1371223,I1371215);
nor I_80450 (I1370819,I1371223,I1371141);
nor I_80451 (I1371254,I1371124,I1272521);
and I_80452 (I1371271,I1371254,I1272545);
or I_80453 (I1371288,I1371271,I1272527);
DFFARX1 I_80454 (I1371288,I3563,I1370833,I1371314,);
not I_80455 (I1371322,I1371314);
nand I_80456 (I1371339,I1371322,I1371062);
not I_80457 (I1370813,I1371339);
nand I_80458 (I1370807,I1371339,I1371079);
nand I_80459 (I1370804,I1371322,I1370946);
not I_80460 (I1371428,I3570);
DFFARX1 I_80461 (I418717,I3563,I1371428,I1371454,);
DFFARX1 I_80462 (I418711,I3563,I1371428,I1371471,);
not I_80463 (I1371479,I1371471);
nor I_80464 (I1371396,I1371454,I1371479);
DFFARX1 I_80465 (I1371479,I3563,I1371428,I1371411,);
nor I_80466 (I1371524,I418699,I418720);
and I_80467 (I1371541,I1371524,I418714);
nor I_80468 (I1371558,I1371541,I418699);
not I_80469 (I1371575,I418699);
and I_80470 (I1371592,I1371575,I418696);
nand I_80471 (I1371609,I1371592,I418708);
nor I_80472 (I1371626,I1371575,I1371609);
DFFARX1 I_80473 (I1371626,I3563,I1371428,I1371393,);
not I_80474 (I1371657,I1371609);
nand I_80475 (I1371674,I1371479,I1371657);
nand I_80476 (I1371405,I1371541,I1371657);
DFFARX1 I_80477 (I1371575,I3563,I1371428,I1371420,);
not I_80478 (I1371719,I418723);
nor I_80479 (I1371736,I1371719,I418696);
nor I_80480 (I1371753,I1371736,I1371558);
DFFARX1 I_80481 (I1371753,I3563,I1371428,I1371417,);
not I_80482 (I1371784,I1371736);
DFFARX1 I_80483 (I1371784,I3563,I1371428,I1371810,);
not I_80484 (I1371818,I1371810);
nor I_80485 (I1371414,I1371818,I1371736);
nor I_80486 (I1371849,I1371719,I418705);
and I_80487 (I1371866,I1371849,I418702);
or I_80488 (I1371883,I1371866,I418696);
DFFARX1 I_80489 (I1371883,I3563,I1371428,I1371909,);
not I_80490 (I1371917,I1371909);
nand I_80491 (I1371934,I1371917,I1371657);
not I_80492 (I1371408,I1371934);
nand I_80493 (I1371402,I1371934,I1371674);
nand I_80494 (I1371399,I1371917,I1371541);
not I_80495 (I1372023,I3570);
DFFARX1 I_80496 (I403434,I3563,I1372023,I1372049,);
DFFARX1 I_80497 (I403428,I3563,I1372023,I1372066,);
not I_80498 (I1372074,I1372066);
nor I_80499 (I1371991,I1372049,I1372074);
DFFARX1 I_80500 (I1372074,I3563,I1372023,I1372006,);
nor I_80501 (I1372119,I403416,I403437);
and I_80502 (I1372136,I1372119,I403431);
nor I_80503 (I1372153,I1372136,I403416);
not I_80504 (I1372170,I403416);
and I_80505 (I1372187,I1372170,I403413);
nand I_80506 (I1372204,I1372187,I403425);
nor I_80507 (I1372221,I1372170,I1372204);
DFFARX1 I_80508 (I1372221,I3563,I1372023,I1371988,);
not I_80509 (I1372252,I1372204);
nand I_80510 (I1372269,I1372074,I1372252);
nand I_80511 (I1372000,I1372136,I1372252);
DFFARX1 I_80512 (I1372170,I3563,I1372023,I1372015,);
not I_80513 (I1372314,I403440);
nor I_80514 (I1372331,I1372314,I403413);
nor I_80515 (I1372348,I1372331,I1372153);
DFFARX1 I_80516 (I1372348,I3563,I1372023,I1372012,);
not I_80517 (I1372379,I1372331);
DFFARX1 I_80518 (I1372379,I3563,I1372023,I1372405,);
not I_80519 (I1372413,I1372405);
nor I_80520 (I1372009,I1372413,I1372331);
nor I_80521 (I1372444,I1372314,I403422);
and I_80522 (I1372461,I1372444,I403419);
or I_80523 (I1372478,I1372461,I403413);
DFFARX1 I_80524 (I1372478,I3563,I1372023,I1372504,);
not I_80525 (I1372512,I1372504);
nand I_80526 (I1372529,I1372512,I1372252);
not I_80527 (I1372003,I1372529);
nand I_80528 (I1371997,I1372529,I1372269);
nand I_80529 (I1371994,I1372512,I1372136);
not I_80530 (I1372618,I3570);
DFFARX1 I_80531 (I68789,I3563,I1372618,I1372644,);
DFFARX1 I_80532 (I68777,I3563,I1372618,I1372661,);
not I_80533 (I1372669,I1372661);
nor I_80534 (I1372586,I1372644,I1372669);
DFFARX1 I_80535 (I1372669,I3563,I1372618,I1372601,);
nor I_80536 (I1372714,I68768,I68792);
and I_80537 (I1372731,I1372714,I68771);
nor I_80538 (I1372748,I1372731,I68768);
not I_80539 (I1372765,I68768);
and I_80540 (I1372782,I1372765,I68774);
nand I_80541 (I1372799,I1372782,I68786);
nor I_80542 (I1372816,I1372765,I1372799);
DFFARX1 I_80543 (I1372816,I3563,I1372618,I1372583,);
not I_80544 (I1372847,I1372799);
nand I_80545 (I1372864,I1372669,I1372847);
nand I_80546 (I1372595,I1372731,I1372847);
DFFARX1 I_80547 (I1372765,I3563,I1372618,I1372610,);
not I_80548 (I1372909,I68768);
nor I_80549 (I1372926,I1372909,I68774);
nor I_80550 (I1372943,I1372926,I1372748);
DFFARX1 I_80551 (I1372943,I3563,I1372618,I1372607,);
not I_80552 (I1372974,I1372926);
DFFARX1 I_80553 (I1372974,I3563,I1372618,I1373000,);
not I_80554 (I1373008,I1373000);
nor I_80555 (I1372604,I1373008,I1372926);
nor I_80556 (I1373039,I1372909,I68771);
and I_80557 (I1373056,I1373039,I68780);
or I_80558 (I1373073,I1373056,I68783);
DFFARX1 I_80559 (I1373073,I3563,I1372618,I1373099,);
not I_80560 (I1373107,I1373099);
nand I_80561 (I1373124,I1373107,I1372847);
not I_80562 (I1372598,I1373124);
nand I_80563 (I1372592,I1373124,I1372864);
nand I_80564 (I1372589,I1373107,I1372731);
not I_80565 (I1373213,I3570);
DFFARX1 I_80566 (I312790,I3563,I1373213,I1373239,);
DFFARX1 I_80567 (I312784,I3563,I1373213,I1373256,);
not I_80568 (I1373264,I1373256);
nor I_80569 (I1373181,I1373239,I1373264);
DFFARX1 I_80570 (I1373264,I3563,I1373213,I1373196,);
nor I_80571 (I1373309,I312772,I312793);
and I_80572 (I1373326,I1373309,I312787);
nor I_80573 (I1373343,I1373326,I312772);
not I_80574 (I1373360,I312772);
and I_80575 (I1373377,I1373360,I312769);
nand I_80576 (I1373394,I1373377,I312781);
nor I_80577 (I1373411,I1373360,I1373394);
DFFARX1 I_80578 (I1373411,I3563,I1373213,I1373178,);
not I_80579 (I1373442,I1373394);
nand I_80580 (I1373459,I1373264,I1373442);
nand I_80581 (I1373190,I1373326,I1373442);
DFFARX1 I_80582 (I1373360,I3563,I1373213,I1373205,);
not I_80583 (I1373504,I312796);
nor I_80584 (I1373521,I1373504,I312769);
nor I_80585 (I1373538,I1373521,I1373343);
DFFARX1 I_80586 (I1373538,I3563,I1373213,I1373202,);
not I_80587 (I1373569,I1373521);
DFFARX1 I_80588 (I1373569,I3563,I1373213,I1373595,);
not I_80589 (I1373603,I1373595);
nor I_80590 (I1373199,I1373603,I1373521);
nor I_80591 (I1373634,I1373504,I312778);
and I_80592 (I1373651,I1373634,I312775);
or I_80593 (I1373668,I1373651,I312769);
DFFARX1 I_80594 (I1373668,I3563,I1373213,I1373694,);
not I_80595 (I1373702,I1373694);
nand I_80596 (I1373719,I1373702,I1373442);
not I_80597 (I1373193,I1373719);
nand I_80598 (I1373187,I1373719,I1373459);
nand I_80599 (I1373184,I1373702,I1373326);
not I_80600 (I1373808,I3570);
DFFARX1 I_80601 (I784438,I3563,I1373808,I1373834,);
DFFARX1 I_80602 (I784420,I3563,I1373808,I1373851,);
not I_80603 (I1373859,I1373851);
nor I_80604 (I1373776,I1373834,I1373859);
DFFARX1 I_80605 (I1373859,I3563,I1373808,I1373791,);
nor I_80606 (I1373904,I784426,I784429);
and I_80607 (I1373921,I1373904,I784417);
nor I_80608 (I1373938,I1373921,I784426);
not I_80609 (I1373955,I784426);
and I_80610 (I1373972,I1373955,I784435);
nand I_80611 (I1373989,I1373972,I784423);
nor I_80612 (I1374006,I1373955,I1373989);
DFFARX1 I_80613 (I1374006,I3563,I1373808,I1373773,);
not I_80614 (I1374037,I1373989);
nand I_80615 (I1374054,I1373859,I1374037);
nand I_80616 (I1373785,I1373921,I1374037);
DFFARX1 I_80617 (I1373955,I3563,I1373808,I1373800,);
not I_80618 (I1374099,I784420);
nor I_80619 (I1374116,I1374099,I784435);
nor I_80620 (I1374133,I1374116,I1373938);
DFFARX1 I_80621 (I1374133,I3563,I1373808,I1373797,);
not I_80622 (I1374164,I1374116);
DFFARX1 I_80623 (I1374164,I3563,I1373808,I1374190,);
not I_80624 (I1374198,I1374190);
nor I_80625 (I1373794,I1374198,I1374116);
nor I_80626 (I1374229,I1374099,I784432);
and I_80627 (I1374246,I1374229,I784441);
or I_80628 (I1374263,I1374246,I784417);
DFFARX1 I_80629 (I1374263,I3563,I1373808,I1374289,);
not I_80630 (I1374297,I1374289);
nand I_80631 (I1374314,I1374297,I1374037);
not I_80632 (I1373788,I1374314);
nand I_80633 (I1373782,I1374314,I1374054);
nand I_80634 (I1373779,I1374297,I1373921);
not I_80635 (I1374403,I3570);
DFFARX1 I_80636 (I7146,I3563,I1374403,I1374429,);
DFFARX1 I_80637 (I7143,I3563,I1374403,I1374446,);
not I_80638 (I1374454,I1374446);
nor I_80639 (I1374371,I1374429,I1374454);
DFFARX1 I_80640 (I1374454,I3563,I1374403,I1374386,);
nor I_80641 (I1374499,I7161,I7158);
and I_80642 (I1374516,I1374499,I7149);
nor I_80643 (I1374533,I1374516,I7161);
not I_80644 (I1374550,I7161);
and I_80645 (I1374567,I1374550,I7146);
nand I_80646 (I1374584,I1374567,I7155);
nor I_80647 (I1374601,I1374550,I1374584);
DFFARX1 I_80648 (I1374601,I3563,I1374403,I1374368,);
not I_80649 (I1374632,I1374584);
nand I_80650 (I1374649,I1374454,I1374632);
nand I_80651 (I1374380,I1374516,I1374632);
DFFARX1 I_80652 (I1374550,I3563,I1374403,I1374395,);
not I_80653 (I1374694,I7164);
nor I_80654 (I1374711,I1374694,I7146);
nor I_80655 (I1374728,I1374711,I1374533);
DFFARX1 I_80656 (I1374728,I3563,I1374403,I1374392,);
not I_80657 (I1374759,I1374711);
DFFARX1 I_80658 (I1374759,I3563,I1374403,I1374785,);
not I_80659 (I1374793,I1374785);
nor I_80660 (I1374389,I1374793,I1374711);
nor I_80661 (I1374824,I1374694,I7143);
and I_80662 (I1374841,I1374824,I7149);
or I_80663 (I1374858,I1374841,I7152);
DFFARX1 I_80664 (I1374858,I3563,I1374403,I1374884,);
not I_80665 (I1374892,I1374884);
nand I_80666 (I1374909,I1374892,I1374632);
not I_80667 (I1374383,I1374909);
nand I_80668 (I1374377,I1374909,I1374649);
nand I_80669 (I1374374,I1374892,I1374516);
not I_80670 (I1374998,I3570);
DFFARX1 I_80671 (I1320717,I3563,I1374998,I1375024,);
DFFARX1 I_80672 (I1320708,I3563,I1374998,I1375041,);
not I_80673 (I1375049,I1375041);
nor I_80674 (I1374966,I1375024,I1375049);
DFFARX1 I_80675 (I1375049,I3563,I1374998,I1374981,);
nor I_80676 (I1375094,I1320699,I1320714);
and I_80677 (I1375111,I1375094,I1320702);
nor I_80678 (I1375128,I1375111,I1320699);
not I_80679 (I1375145,I1320699);
and I_80680 (I1375162,I1375145,I1320705);
nand I_80681 (I1375179,I1375162,I1320723);
nor I_80682 (I1375196,I1375145,I1375179);
DFFARX1 I_80683 (I1375196,I3563,I1374998,I1374963,);
not I_80684 (I1375227,I1375179);
nand I_80685 (I1375244,I1375049,I1375227);
nand I_80686 (I1374975,I1375111,I1375227);
DFFARX1 I_80687 (I1375145,I3563,I1374998,I1374990,);
not I_80688 (I1375289,I1320699);
nor I_80689 (I1375306,I1375289,I1320705);
nor I_80690 (I1375323,I1375306,I1375128);
DFFARX1 I_80691 (I1375323,I3563,I1374998,I1374987,);
not I_80692 (I1375354,I1375306);
DFFARX1 I_80693 (I1375354,I3563,I1374998,I1375380,);
not I_80694 (I1375388,I1375380);
nor I_80695 (I1374984,I1375388,I1375306);
nor I_80696 (I1375419,I1375289,I1320702);
and I_80697 (I1375436,I1375419,I1320711);
or I_80698 (I1375453,I1375436,I1320720);
DFFARX1 I_80699 (I1375453,I3563,I1374998,I1375479,);
not I_80700 (I1375487,I1375479);
nand I_80701 (I1375504,I1375487,I1375227);
not I_80702 (I1374978,I1375504);
nand I_80703 (I1374972,I1375504,I1375244);
nand I_80704 (I1374969,I1375487,I1375111);
not I_80705 (I1375593,I3570);
DFFARX1 I_80706 (I720858,I3563,I1375593,I1375619,);
DFFARX1 I_80707 (I720840,I3563,I1375593,I1375636,);
not I_80708 (I1375644,I1375636);
nor I_80709 (I1375561,I1375619,I1375644);
DFFARX1 I_80710 (I1375644,I3563,I1375593,I1375576,);
nor I_80711 (I1375689,I720846,I720849);
and I_80712 (I1375706,I1375689,I720837);
nor I_80713 (I1375723,I1375706,I720846);
not I_80714 (I1375740,I720846);
and I_80715 (I1375757,I1375740,I720855);
nand I_80716 (I1375774,I1375757,I720843);
nor I_80717 (I1375791,I1375740,I1375774);
DFFARX1 I_80718 (I1375791,I3563,I1375593,I1375558,);
not I_80719 (I1375822,I1375774);
nand I_80720 (I1375839,I1375644,I1375822);
nand I_80721 (I1375570,I1375706,I1375822);
DFFARX1 I_80722 (I1375740,I3563,I1375593,I1375585,);
not I_80723 (I1375884,I720840);
nor I_80724 (I1375901,I1375884,I720855);
nor I_80725 (I1375918,I1375901,I1375723);
DFFARX1 I_80726 (I1375918,I3563,I1375593,I1375582,);
not I_80727 (I1375949,I1375901);
DFFARX1 I_80728 (I1375949,I3563,I1375593,I1375975,);
not I_80729 (I1375983,I1375975);
nor I_80730 (I1375579,I1375983,I1375901);
nor I_80731 (I1376014,I1375884,I720852);
and I_80732 (I1376031,I1376014,I720861);
or I_80733 (I1376048,I1376031,I720837);
DFFARX1 I_80734 (I1376048,I3563,I1375593,I1376074,);
not I_80735 (I1376082,I1376074);
nand I_80736 (I1376099,I1376082,I1375822);
not I_80737 (I1375573,I1376099);
nand I_80738 (I1375567,I1376099,I1375839);
nand I_80739 (I1375564,I1376082,I1375706);
not I_80740 (I1376188,I3570);
DFFARX1 I_80741 (I753804,I3563,I1376188,I1376214,);
DFFARX1 I_80742 (I753786,I3563,I1376188,I1376231,);
not I_80743 (I1376239,I1376231);
nor I_80744 (I1376156,I1376214,I1376239);
DFFARX1 I_80745 (I1376239,I3563,I1376188,I1376171,);
nor I_80746 (I1376284,I753792,I753795);
and I_80747 (I1376301,I1376284,I753783);
nor I_80748 (I1376318,I1376301,I753792);
not I_80749 (I1376335,I753792);
and I_80750 (I1376352,I1376335,I753801);
nand I_80751 (I1376369,I1376352,I753789);
nor I_80752 (I1376386,I1376335,I1376369);
DFFARX1 I_80753 (I1376386,I3563,I1376188,I1376153,);
not I_80754 (I1376417,I1376369);
nand I_80755 (I1376434,I1376239,I1376417);
nand I_80756 (I1376165,I1376301,I1376417);
DFFARX1 I_80757 (I1376335,I3563,I1376188,I1376180,);
not I_80758 (I1376479,I753786);
nor I_80759 (I1376496,I1376479,I753801);
nor I_80760 (I1376513,I1376496,I1376318);
DFFARX1 I_80761 (I1376513,I3563,I1376188,I1376177,);
not I_80762 (I1376544,I1376496);
DFFARX1 I_80763 (I1376544,I3563,I1376188,I1376570,);
not I_80764 (I1376578,I1376570);
nor I_80765 (I1376174,I1376578,I1376496);
nor I_80766 (I1376609,I1376479,I753798);
and I_80767 (I1376626,I1376609,I753807);
or I_80768 (I1376643,I1376626,I753783);
DFFARX1 I_80769 (I1376643,I3563,I1376188,I1376669,);
not I_80770 (I1376677,I1376669);
nand I_80771 (I1376694,I1376677,I1376417);
not I_80772 (I1376168,I1376694);
nand I_80773 (I1376162,I1376694,I1376434);
nand I_80774 (I1376159,I1376677,I1376301);
not I_80775 (I1376783,I3570);
DFFARX1 I_80776 (I1322451,I3563,I1376783,I1376809,);
DFFARX1 I_80777 (I1322442,I3563,I1376783,I1376826,);
not I_80778 (I1376834,I1376826);
nor I_80779 (I1376751,I1376809,I1376834);
DFFARX1 I_80780 (I1376834,I3563,I1376783,I1376766,);
nor I_80781 (I1376879,I1322433,I1322448);
and I_80782 (I1376896,I1376879,I1322436);
nor I_80783 (I1376913,I1376896,I1322433);
not I_80784 (I1376930,I1322433);
and I_80785 (I1376947,I1376930,I1322439);
nand I_80786 (I1376964,I1376947,I1322457);
nor I_80787 (I1376981,I1376930,I1376964);
DFFARX1 I_80788 (I1376981,I3563,I1376783,I1376748,);
not I_80789 (I1377012,I1376964);
nand I_80790 (I1377029,I1376834,I1377012);
nand I_80791 (I1376760,I1376896,I1377012);
DFFARX1 I_80792 (I1376930,I3563,I1376783,I1376775,);
not I_80793 (I1377074,I1322433);
nor I_80794 (I1377091,I1377074,I1322439);
nor I_80795 (I1377108,I1377091,I1376913);
DFFARX1 I_80796 (I1377108,I3563,I1376783,I1376772,);
not I_80797 (I1377139,I1377091);
DFFARX1 I_80798 (I1377139,I3563,I1376783,I1377165,);
not I_80799 (I1377173,I1377165);
nor I_80800 (I1376769,I1377173,I1377091);
nor I_80801 (I1377204,I1377074,I1322436);
and I_80802 (I1377221,I1377204,I1322445);
or I_80803 (I1377238,I1377221,I1322454);
DFFARX1 I_80804 (I1377238,I3563,I1376783,I1377264,);
not I_80805 (I1377272,I1377264);
nand I_80806 (I1377289,I1377272,I1377012);
not I_80807 (I1376763,I1377289);
nand I_80808 (I1376757,I1377289,I1377029);
nand I_80809 (I1376754,I1377272,I1376896);
not I_80810 (I1377378,I3570);
DFFARX1 I_80811 (I325965,I3563,I1377378,I1377404,);
DFFARX1 I_80812 (I325959,I3563,I1377378,I1377421,);
not I_80813 (I1377429,I1377421);
nor I_80814 (I1377346,I1377404,I1377429);
DFFARX1 I_80815 (I1377429,I3563,I1377378,I1377361,);
nor I_80816 (I1377474,I325947,I325968);
and I_80817 (I1377491,I1377474,I325962);
nor I_80818 (I1377508,I1377491,I325947);
not I_80819 (I1377525,I325947);
and I_80820 (I1377542,I1377525,I325944);
nand I_80821 (I1377559,I1377542,I325956);
nor I_80822 (I1377576,I1377525,I1377559);
DFFARX1 I_80823 (I1377576,I3563,I1377378,I1377343,);
not I_80824 (I1377607,I1377559);
nand I_80825 (I1377624,I1377429,I1377607);
nand I_80826 (I1377355,I1377491,I1377607);
DFFARX1 I_80827 (I1377525,I3563,I1377378,I1377370,);
not I_80828 (I1377669,I325971);
nor I_80829 (I1377686,I1377669,I325944);
nor I_80830 (I1377703,I1377686,I1377508);
DFFARX1 I_80831 (I1377703,I3563,I1377378,I1377367,);
not I_80832 (I1377734,I1377686);
DFFARX1 I_80833 (I1377734,I3563,I1377378,I1377760,);
not I_80834 (I1377768,I1377760);
nor I_80835 (I1377364,I1377768,I1377686);
nor I_80836 (I1377799,I1377669,I325953);
and I_80837 (I1377816,I1377799,I325950);
or I_80838 (I1377833,I1377816,I325944);
DFFARX1 I_80839 (I1377833,I3563,I1377378,I1377859,);
not I_80840 (I1377867,I1377859);
nand I_80841 (I1377884,I1377867,I1377607);
not I_80842 (I1377358,I1377884);
nand I_80843 (I1377352,I1377884,I1377624);
nand I_80844 (I1377349,I1377867,I1377491);
not I_80845 (I1377973,I3570);
DFFARX1 I_80846 (I1195616,I3563,I1377973,I1377999,);
DFFARX1 I_80847 (I1195628,I3563,I1377973,I1378016,);
not I_80848 (I1378024,I1378016);
nor I_80849 (I1377941,I1377999,I1378024);
DFFARX1 I_80850 (I1378024,I3563,I1377973,I1377956,);
nor I_80851 (I1378069,I1195625,I1195619);
and I_80852 (I1378086,I1378069,I1195613);
nor I_80853 (I1378103,I1378086,I1195625);
not I_80854 (I1378120,I1195625);
and I_80855 (I1378137,I1378120,I1195622);
nand I_80856 (I1378154,I1378137,I1195613);
nor I_80857 (I1378171,I1378120,I1378154);
DFFARX1 I_80858 (I1378171,I3563,I1377973,I1377938,);
not I_80859 (I1378202,I1378154);
nand I_80860 (I1378219,I1378024,I1378202);
nand I_80861 (I1377950,I1378086,I1378202);
DFFARX1 I_80862 (I1378120,I3563,I1377973,I1377965,);
not I_80863 (I1378264,I1195637);
nor I_80864 (I1378281,I1378264,I1195622);
nor I_80865 (I1378298,I1378281,I1378103);
DFFARX1 I_80866 (I1378298,I3563,I1377973,I1377962,);
not I_80867 (I1378329,I1378281);
DFFARX1 I_80868 (I1378329,I3563,I1377973,I1378355,);
not I_80869 (I1378363,I1378355);
nor I_80870 (I1377959,I1378363,I1378281);
nor I_80871 (I1378394,I1378264,I1195631);
and I_80872 (I1378411,I1378394,I1195634);
or I_80873 (I1378428,I1378411,I1195616);
DFFARX1 I_80874 (I1378428,I3563,I1377973,I1378454,);
not I_80875 (I1378462,I1378454);
nand I_80876 (I1378479,I1378462,I1378202);
not I_80877 (I1377953,I1378479);
nand I_80878 (I1377947,I1378479,I1378219);
nand I_80879 (I1377944,I1378462,I1378086);
not I_80880 (I1378568,I3570);
DFFARX1 I_80881 (I5956,I3563,I1378568,I1378594,);
DFFARX1 I_80882 (I5953,I3563,I1378568,I1378611,);
not I_80883 (I1378619,I1378611);
nor I_80884 (I1378536,I1378594,I1378619);
DFFARX1 I_80885 (I1378619,I3563,I1378568,I1378551,);
nor I_80886 (I1378664,I5971,I5968);
and I_80887 (I1378681,I1378664,I5959);
nor I_80888 (I1378698,I1378681,I5971);
not I_80889 (I1378715,I5971);
and I_80890 (I1378732,I1378715,I5956);
nand I_80891 (I1378749,I1378732,I5965);
nor I_80892 (I1378766,I1378715,I1378749);
DFFARX1 I_80893 (I1378766,I3563,I1378568,I1378533,);
not I_80894 (I1378797,I1378749);
nand I_80895 (I1378814,I1378619,I1378797);
nand I_80896 (I1378545,I1378681,I1378797);
DFFARX1 I_80897 (I1378715,I3563,I1378568,I1378560,);
not I_80898 (I1378859,I5974);
nor I_80899 (I1378876,I1378859,I5956);
nor I_80900 (I1378893,I1378876,I1378698);
DFFARX1 I_80901 (I1378893,I3563,I1378568,I1378557,);
not I_80902 (I1378924,I1378876);
DFFARX1 I_80903 (I1378924,I3563,I1378568,I1378950,);
not I_80904 (I1378958,I1378950);
nor I_80905 (I1378554,I1378958,I1378876);
nor I_80906 (I1378989,I1378859,I5953);
and I_80907 (I1379006,I1378989,I5959);
or I_80908 (I1379023,I1379006,I5962);
DFFARX1 I_80909 (I1379023,I3563,I1378568,I1379049,);
not I_80910 (I1379057,I1379049);
nand I_80911 (I1379074,I1379057,I1378797);
not I_80912 (I1378548,I1379074);
nand I_80913 (I1378542,I1379074,I1378814);
nand I_80914 (I1378539,I1379057,I1378681);
not I_80915 (I1379163,I3570);
DFFARX1 I_80916 (I676930,I3563,I1379163,I1379189,);
DFFARX1 I_80917 (I676912,I3563,I1379163,I1379206,);
not I_80918 (I1379214,I1379206);
nor I_80919 (I1379131,I1379189,I1379214);
DFFARX1 I_80920 (I1379214,I3563,I1379163,I1379146,);
nor I_80921 (I1379259,I676918,I676921);
and I_80922 (I1379276,I1379259,I676909);
nor I_80923 (I1379293,I1379276,I676918);
not I_80924 (I1379310,I676918);
and I_80925 (I1379327,I1379310,I676927);
nand I_80926 (I1379344,I1379327,I676915);
nor I_80927 (I1379361,I1379310,I1379344);
DFFARX1 I_80928 (I1379361,I3563,I1379163,I1379128,);
not I_80929 (I1379392,I1379344);
nand I_80930 (I1379409,I1379214,I1379392);
nand I_80931 (I1379140,I1379276,I1379392);
DFFARX1 I_80932 (I1379310,I3563,I1379163,I1379155,);
not I_80933 (I1379454,I676912);
nor I_80934 (I1379471,I1379454,I676927);
nor I_80935 (I1379488,I1379471,I1379293);
DFFARX1 I_80936 (I1379488,I3563,I1379163,I1379152,);
not I_80937 (I1379519,I1379471);
DFFARX1 I_80938 (I1379519,I3563,I1379163,I1379545,);
not I_80939 (I1379553,I1379545);
nor I_80940 (I1379149,I1379553,I1379471);
nor I_80941 (I1379584,I1379454,I676924);
and I_80942 (I1379601,I1379584,I676933);
or I_80943 (I1379618,I1379601,I676909);
DFFARX1 I_80944 (I1379618,I3563,I1379163,I1379644,);
not I_80945 (I1379652,I1379644);
nand I_80946 (I1379669,I1379652,I1379392);
not I_80947 (I1379143,I1379669);
nand I_80948 (I1379137,I1379669,I1379409);
nand I_80949 (I1379134,I1379652,I1379276);
not I_80950 (I1379758,I3570);
DFFARX1 I_80951 (I691380,I3563,I1379758,I1379784,);
DFFARX1 I_80952 (I691362,I3563,I1379758,I1379801,);
not I_80953 (I1379809,I1379801);
nor I_80954 (I1379726,I1379784,I1379809);
DFFARX1 I_80955 (I1379809,I3563,I1379758,I1379741,);
nor I_80956 (I1379854,I691368,I691371);
and I_80957 (I1379871,I1379854,I691359);
nor I_80958 (I1379888,I1379871,I691368);
not I_80959 (I1379905,I691368);
and I_80960 (I1379922,I1379905,I691377);
nand I_80961 (I1379939,I1379922,I691365);
nor I_80962 (I1379956,I1379905,I1379939);
DFFARX1 I_80963 (I1379956,I3563,I1379758,I1379723,);
not I_80964 (I1379987,I1379939);
nand I_80965 (I1380004,I1379809,I1379987);
nand I_80966 (I1379735,I1379871,I1379987);
DFFARX1 I_80967 (I1379905,I3563,I1379758,I1379750,);
not I_80968 (I1380049,I691362);
nor I_80969 (I1380066,I1380049,I691377);
nor I_80970 (I1380083,I1380066,I1379888);
DFFARX1 I_80971 (I1380083,I3563,I1379758,I1379747,);
not I_80972 (I1380114,I1380066);
DFFARX1 I_80973 (I1380114,I3563,I1379758,I1380140,);
not I_80974 (I1380148,I1380140);
nor I_80975 (I1379744,I1380148,I1380066);
nor I_80976 (I1380179,I1380049,I691374);
and I_80977 (I1380196,I1380179,I691383);
or I_80978 (I1380213,I1380196,I691359);
DFFARX1 I_80979 (I1380213,I3563,I1379758,I1380239,);
not I_80980 (I1380247,I1380239);
nand I_80981 (I1380264,I1380247,I1379987);
not I_80982 (I1379738,I1380264);
nand I_80983 (I1379732,I1380264,I1380004);
nand I_80984 (I1379729,I1380247,I1379871);
not I_80985 (I1380353,I3570);
DFFARX1 I_80986 (I483330,I3563,I1380353,I1380379,);
DFFARX1 I_80987 (I483336,I3563,I1380353,I1380396,);
not I_80988 (I1380404,I1380396);
nor I_80989 (I1380321,I1380379,I1380404);
DFFARX1 I_80990 (I1380404,I3563,I1380353,I1380336,);
nor I_80991 (I1380449,I483345,I483330);
and I_80992 (I1380466,I1380449,I483357);
nor I_80993 (I1380483,I1380466,I483345);
not I_80994 (I1380500,I483345);
and I_80995 (I1380517,I1380500,I483333);
nand I_80996 (I1380534,I1380517,I483354);
nor I_80997 (I1380551,I1380500,I1380534);
DFFARX1 I_80998 (I1380551,I3563,I1380353,I1380318,);
not I_80999 (I1380582,I1380534);
nand I_81000 (I1380599,I1380404,I1380582);
nand I_81001 (I1380330,I1380466,I1380582);
DFFARX1 I_81002 (I1380500,I3563,I1380353,I1380345,);
not I_81003 (I1380644,I483342);
nor I_81004 (I1380661,I1380644,I483333);
nor I_81005 (I1380678,I1380661,I1380483);
DFFARX1 I_81006 (I1380678,I3563,I1380353,I1380342,);
not I_81007 (I1380709,I1380661);
DFFARX1 I_81008 (I1380709,I3563,I1380353,I1380735,);
not I_81009 (I1380743,I1380735);
nor I_81010 (I1380339,I1380743,I1380661);
nor I_81011 (I1380774,I1380644,I483339);
and I_81012 (I1380791,I1380774,I483351);
or I_81013 (I1380808,I1380791,I483348);
DFFARX1 I_81014 (I1380808,I3563,I1380353,I1380834,);
not I_81015 (I1380842,I1380834);
nand I_81016 (I1380859,I1380842,I1380582);
not I_81017 (I1380333,I1380859);
nand I_81018 (I1380327,I1380859,I1380599);
nand I_81019 (I1380324,I1380842,I1380466);
not I_81020 (I1380948,I3570);
DFFARX1 I_81021 (I1325316,I3563,I1380948,I1380974,);
DFFARX1 I_81022 (I1325301,I3563,I1380948,I1380991,);
not I_81023 (I1380999,I1380991);
nor I_81024 (I1380916,I1380974,I1380999);
DFFARX1 I_81025 (I1380999,I3563,I1380948,I1380931,);
nor I_81026 (I1381044,I1325298,I1325307);
and I_81027 (I1381061,I1381044,I1325313);
nor I_81028 (I1381078,I1381061,I1325298);
not I_81029 (I1381095,I1325298);
and I_81030 (I1381112,I1381095,I1325295);
nand I_81031 (I1381129,I1381112,I1325289);
nor I_81032 (I1381146,I1381095,I1381129);
DFFARX1 I_81033 (I1381146,I3563,I1380948,I1380913,);
not I_81034 (I1381177,I1381129);
nand I_81035 (I1381194,I1380999,I1381177);
nand I_81036 (I1380925,I1381061,I1381177);
DFFARX1 I_81037 (I1381095,I3563,I1380948,I1380940,);
not I_81038 (I1381239,I1325289);
nor I_81039 (I1381256,I1381239,I1325295);
nor I_81040 (I1381273,I1381256,I1381078);
DFFARX1 I_81041 (I1381273,I3563,I1380948,I1380937,);
not I_81042 (I1381304,I1381256);
DFFARX1 I_81043 (I1381304,I3563,I1380948,I1381330,);
not I_81044 (I1381338,I1381330);
nor I_81045 (I1380934,I1381338,I1381256);
nor I_81046 (I1381369,I1381239,I1325304);
and I_81047 (I1381386,I1381369,I1325310);
or I_81048 (I1381403,I1381386,I1325292);
DFFARX1 I_81049 (I1381403,I3563,I1380948,I1381429,);
not I_81050 (I1381437,I1381429);
nand I_81051 (I1381454,I1381437,I1381177);
not I_81052 (I1380928,I1381454);
nand I_81053 (I1380922,I1381454,I1381194);
nand I_81054 (I1380919,I1381437,I1381061);
not I_81055 (I1381543,I3570);
DFFARX1 I_81056 (I1305689,I3563,I1381543,I1381569,);
DFFARX1 I_81057 (I1305680,I3563,I1381543,I1381586,);
not I_81058 (I1381594,I1381586);
nor I_81059 (I1381511,I1381569,I1381594);
DFFARX1 I_81060 (I1381594,I3563,I1381543,I1381526,);
nor I_81061 (I1381639,I1305671,I1305686);
and I_81062 (I1381656,I1381639,I1305674);
nor I_81063 (I1381673,I1381656,I1305671);
not I_81064 (I1381690,I1305671);
and I_81065 (I1381707,I1381690,I1305677);
nand I_81066 (I1381724,I1381707,I1305695);
nor I_81067 (I1381741,I1381690,I1381724);
DFFARX1 I_81068 (I1381741,I3563,I1381543,I1381508,);
not I_81069 (I1381772,I1381724);
nand I_81070 (I1381789,I1381594,I1381772);
nand I_81071 (I1381520,I1381656,I1381772);
DFFARX1 I_81072 (I1381690,I3563,I1381543,I1381535,);
not I_81073 (I1381834,I1305671);
nor I_81074 (I1381851,I1381834,I1305677);
nor I_81075 (I1381868,I1381851,I1381673);
DFFARX1 I_81076 (I1381868,I3563,I1381543,I1381532,);
not I_81077 (I1381899,I1381851);
DFFARX1 I_81078 (I1381899,I3563,I1381543,I1381925,);
not I_81079 (I1381933,I1381925);
nor I_81080 (I1381529,I1381933,I1381851);
nor I_81081 (I1381964,I1381834,I1305674);
and I_81082 (I1381981,I1381964,I1305683);
or I_81083 (I1381998,I1381981,I1305692);
DFFARX1 I_81084 (I1381998,I3563,I1381543,I1382024,);
not I_81085 (I1382032,I1382024);
nand I_81086 (I1382049,I1382032,I1381772);
not I_81087 (I1381523,I1382049);
nand I_81088 (I1381517,I1382049,I1381789);
nand I_81089 (I1381514,I1382032,I1381656);
not I_81090 (I1382138,I3570);
DFFARX1 I_81091 (I20829,I3563,I1382138,I1382164,);
DFFARX1 I_81092 (I20811,I3563,I1382138,I1382181,);
not I_81093 (I1382189,I1382181);
nor I_81094 (I1382106,I1382164,I1382189);
DFFARX1 I_81095 (I1382189,I3563,I1382138,I1382121,);
nor I_81096 (I1382234,I20811,I20826);
and I_81097 (I1382251,I1382234,I20820);
nor I_81098 (I1382268,I1382251,I20811);
not I_81099 (I1382285,I20811);
and I_81100 (I1382302,I1382285,I20814);
nand I_81101 (I1382319,I1382302,I20817);
nor I_81102 (I1382336,I1382285,I1382319);
DFFARX1 I_81103 (I1382336,I3563,I1382138,I1382103,);
not I_81104 (I1382367,I1382319);
nand I_81105 (I1382384,I1382189,I1382367);
nand I_81106 (I1382115,I1382251,I1382367);
DFFARX1 I_81107 (I1382285,I3563,I1382138,I1382130,);
not I_81108 (I1382429,I20823);
nor I_81109 (I1382446,I1382429,I20814);
nor I_81110 (I1382463,I1382446,I1382268);
DFFARX1 I_81111 (I1382463,I3563,I1382138,I1382127,);
not I_81112 (I1382494,I1382446);
DFFARX1 I_81113 (I1382494,I3563,I1382138,I1382520,);
not I_81114 (I1382528,I1382520);
nor I_81115 (I1382124,I1382528,I1382446);
nor I_81116 (I1382559,I1382429,I20835);
and I_81117 (I1382576,I1382559,I20832);
or I_81118 (I1382593,I1382576,I20814);
DFFARX1 I_81119 (I1382593,I3563,I1382138,I1382619,);
not I_81120 (I1382627,I1382619);
nand I_81121 (I1382644,I1382627,I1382367);
not I_81122 (I1382118,I1382644);
nand I_81123 (I1382112,I1382644,I1382384);
nand I_81124 (I1382109,I1382627,I1382251);
not I_81125 (I1382733,I3570);
DFFARX1 I_81126 (I1055086,I3563,I1382733,I1382759,);
DFFARX1 I_81127 (I1055077,I3563,I1382733,I1382776,);
not I_81128 (I1382784,I1382776);
nor I_81129 (I1382701,I1382759,I1382784);
DFFARX1 I_81130 (I1382784,I3563,I1382733,I1382716,);
nor I_81131 (I1382829,I1055083,I1055092);
and I_81132 (I1382846,I1382829,I1055095);
nor I_81133 (I1382863,I1382846,I1055083);
not I_81134 (I1382880,I1055083);
and I_81135 (I1382897,I1382880,I1055074);
nand I_81136 (I1382914,I1382897,I1055080);
nor I_81137 (I1382931,I1382880,I1382914);
DFFARX1 I_81138 (I1382931,I3563,I1382733,I1382698,);
not I_81139 (I1382962,I1382914);
nand I_81140 (I1382979,I1382784,I1382962);
nand I_81141 (I1382710,I1382846,I1382962);
DFFARX1 I_81142 (I1382880,I3563,I1382733,I1382725,);
not I_81143 (I1383024,I1055089);
nor I_81144 (I1383041,I1383024,I1055074);
nor I_81145 (I1383058,I1383041,I1382863);
DFFARX1 I_81146 (I1383058,I3563,I1382733,I1382722,);
not I_81147 (I1383089,I1383041);
DFFARX1 I_81148 (I1383089,I3563,I1382733,I1383115,);
not I_81149 (I1383123,I1383115);
nor I_81150 (I1382719,I1383123,I1383041);
nor I_81151 (I1383154,I1383024,I1055074);
and I_81152 (I1383171,I1383154,I1055077);
or I_81153 (I1383188,I1383171,I1055080);
DFFARX1 I_81154 (I1383188,I3563,I1382733,I1383214,);
not I_81155 (I1383222,I1383214);
nand I_81156 (I1383239,I1383222,I1382962);
not I_81157 (I1382713,I1383239);
nand I_81158 (I1382707,I1383239,I1382979);
nand I_81159 (I1382704,I1383222,I1382846);
not I_81160 (I1383328,I3570);
DFFARX1 I_81161 (I605258,I3563,I1383328,I1383354,);
DFFARX1 I_81162 (I605252,I3563,I1383328,I1383371,);
not I_81163 (I1383379,I1383371);
nor I_81164 (I1383296,I1383354,I1383379);
DFFARX1 I_81165 (I1383379,I3563,I1383328,I1383311,);
nor I_81166 (I1383424,I605249,I605240);
and I_81167 (I1383441,I1383424,I605237);
nor I_81168 (I1383458,I1383441,I605249);
not I_81169 (I1383475,I605249);
and I_81170 (I1383492,I1383475,I605243);
nand I_81171 (I1383509,I1383492,I605255);
nor I_81172 (I1383526,I1383475,I1383509);
DFFARX1 I_81173 (I1383526,I3563,I1383328,I1383293,);
not I_81174 (I1383557,I1383509);
nand I_81175 (I1383574,I1383379,I1383557);
nand I_81176 (I1383305,I1383441,I1383557);
DFFARX1 I_81177 (I1383475,I3563,I1383328,I1383320,);
not I_81178 (I1383619,I605261);
nor I_81179 (I1383636,I1383619,I605243);
nor I_81180 (I1383653,I1383636,I1383458);
DFFARX1 I_81181 (I1383653,I3563,I1383328,I1383317,);
not I_81182 (I1383684,I1383636);
DFFARX1 I_81183 (I1383684,I3563,I1383328,I1383710,);
not I_81184 (I1383718,I1383710);
nor I_81185 (I1383314,I1383718,I1383636);
nor I_81186 (I1383749,I1383619,I605240);
and I_81187 (I1383766,I1383749,I605246);
or I_81188 (I1383783,I1383766,I605237);
DFFARX1 I_81189 (I1383783,I3563,I1383328,I1383809,);
not I_81190 (I1383817,I1383809);
nand I_81191 (I1383834,I1383817,I1383557);
not I_81192 (I1383308,I1383834);
nand I_81193 (I1383302,I1383834,I1383574);
nand I_81194 (I1383299,I1383817,I1383441);
not I_81195 (I1383923,I3570);
DFFARX1 I_81196 (I54030,I3563,I1383923,I1383949,);
DFFARX1 I_81197 (I54012,I3563,I1383923,I1383966,);
not I_81198 (I1383974,I1383966);
nor I_81199 (I1383891,I1383949,I1383974);
DFFARX1 I_81200 (I1383974,I3563,I1383923,I1383906,);
nor I_81201 (I1384019,I54012,I54027);
and I_81202 (I1384036,I1384019,I54021);
nor I_81203 (I1384053,I1384036,I54012);
not I_81204 (I1384070,I54012);
and I_81205 (I1384087,I1384070,I54015);
nand I_81206 (I1384104,I1384087,I54018);
nor I_81207 (I1384121,I1384070,I1384104);
DFFARX1 I_81208 (I1384121,I3563,I1383923,I1383888,);
not I_81209 (I1384152,I1384104);
nand I_81210 (I1384169,I1383974,I1384152);
nand I_81211 (I1383900,I1384036,I1384152);
DFFARX1 I_81212 (I1384070,I3563,I1383923,I1383915,);
not I_81213 (I1384214,I54024);
nor I_81214 (I1384231,I1384214,I54015);
nor I_81215 (I1384248,I1384231,I1384053);
DFFARX1 I_81216 (I1384248,I3563,I1383923,I1383912,);
not I_81217 (I1384279,I1384231);
DFFARX1 I_81218 (I1384279,I3563,I1383923,I1384305,);
not I_81219 (I1384313,I1384305);
nor I_81220 (I1383909,I1384313,I1384231);
nor I_81221 (I1384344,I1384214,I54036);
and I_81222 (I1384361,I1384344,I54033);
or I_81223 (I1384378,I1384361,I54015);
DFFARX1 I_81224 (I1384378,I3563,I1383923,I1384404,);
not I_81225 (I1384412,I1384404);
nand I_81226 (I1384429,I1384412,I1384152);
not I_81227 (I1383903,I1384429);
nand I_81228 (I1383897,I1384429,I1384169);
nand I_81229 (I1383894,I1384412,I1384036);
not I_81230 (I1384518,I3570);
DFFARX1 I_81231 (I2820,I3563,I1384518,I1384544,);
DFFARX1 I_81232 (I2404,I3563,I1384518,I1384561,);
not I_81233 (I1384569,I1384561);
nor I_81234 (I1384486,I1384544,I1384569);
DFFARX1 I_81235 (I1384569,I3563,I1384518,I1384501,);
nor I_81236 (I1384614,I2676,I1964);
and I_81237 (I1384631,I1384614,I3220);
nor I_81238 (I1384648,I1384631,I2676);
not I_81239 (I1384665,I2676);
and I_81240 (I1384682,I1384665,I3452);
nand I_81241 (I1384699,I1384682,I1596);
nor I_81242 (I1384716,I1384665,I1384699);
DFFARX1 I_81243 (I1384716,I3563,I1384518,I1384483,);
not I_81244 (I1384747,I1384699);
nand I_81245 (I1384764,I1384569,I1384747);
nand I_81246 (I1384495,I1384631,I1384747);
DFFARX1 I_81247 (I1384665,I3563,I1384518,I1384510,);
not I_81248 (I1384809,I2996);
nor I_81249 (I1384826,I1384809,I3452);
nor I_81250 (I1384843,I1384826,I1384648);
DFFARX1 I_81251 (I1384843,I3563,I1384518,I1384507,);
not I_81252 (I1384874,I1384826);
DFFARX1 I_81253 (I1384874,I3563,I1384518,I1384900,);
not I_81254 (I1384908,I1384900);
nor I_81255 (I1384504,I1384908,I1384826);
nor I_81256 (I1384939,I1384809,I1692);
and I_81257 (I1384956,I1384939,I2508);
or I_81258 (I1384973,I1384956,I2068);
DFFARX1 I_81259 (I1384973,I3563,I1384518,I1384999,);
not I_81260 (I1385007,I1384999);
nand I_81261 (I1385024,I1385007,I1384747);
not I_81262 (I1384498,I1385024);
nand I_81263 (I1384492,I1385024,I1384764);
nand I_81264 (I1384489,I1385007,I1384631);
not I_81265 (I1385113,I3570);
DFFARX1 I_81266 (I95139,I3563,I1385113,I1385139,);
DFFARX1 I_81267 (I95127,I3563,I1385113,I1385156,);
not I_81268 (I1385164,I1385156);
nor I_81269 (I1385081,I1385139,I1385164);
DFFARX1 I_81270 (I1385164,I3563,I1385113,I1385096,);
nor I_81271 (I1385209,I95118,I95142);
and I_81272 (I1385226,I1385209,I95121);
nor I_81273 (I1385243,I1385226,I95118);
not I_81274 (I1385260,I95118);
and I_81275 (I1385277,I1385260,I95124);
nand I_81276 (I1385294,I1385277,I95136);
nor I_81277 (I1385311,I1385260,I1385294);
DFFARX1 I_81278 (I1385311,I3563,I1385113,I1385078,);
not I_81279 (I1385342,I1385294);
nand I_81280 (I1385359,I1385164,I1385342);
nand I_81281 (I1385090,I1385226,I1385342);
DFFARX1 I_81282 (I1385260,I3563,I1385113,I1385105,);
not I_81283 (I1385404,I95118);
nor I_81284 (I1385421,I1385404,I95124);
nor I_81285 (I1385438,I1385421,I1385243);
DFFARX1 I_81286 (I1385438,I3563,I1385113,I1385102,);
not I_81287 (I1385469,I1385421);
DFFARX1 I_81288 (I1385469,I3563,I1385113,I1385495,);
not I_81289 (I1385503,I1385495);
nor I_81290 (I1385099,I1385503,I1385421);
nor I_81291 (I1385534,I1385404,I95121);
and I_81292 (I1385551,I1385534,I95130);
or I_81293 (I1385568,I1385551,I95133);
DFFARX1 I_81294 (I1385568,I3563,I1385113,I1385594,);
not I_81295 (I1385602,I1385594);
nand I_81296 (I1385619,I1385602,I1385342);
not I_81297 (I1385093,I1385619);
nand I_81298 (I1385087,I1385619,I1385359);
nand I_81299 (I1385084,I1385602,I1385226);
not I_81300 (I1385708,I3570);
DFFARX1 I_81301 (I1220470,I3563,I1385708,I1385734,);
DFFARX1 I_81302 (I1220482,I3563,I1385708,I1385751,);
not I_81303 (I1385759,I1385751);
nor I_81304 (I1385676,I1385734,I1385759);
DFFARX1 I_81305 (I1385759,I3563,I1385708,I1385691,);
nor I_81306 (I1385804,I1220479,I1220473);
and I_81307 (I1385821,I1385804,I1220467);
nor I_81308 (I1385838,I1385821,I1220479);
not I_81309 (I1385855,I1220479);
and I_81310 (I1385872,I1385855,I1220476);
nand I_81311 (I1385889,I1385872,I1220467);
nor I_81312 (I1385906,I1385855,I1385889);
DFFARX1 I_81313 (I1385906,I3563,I1385708,I1385673,);
not I_81314 (I1385937,I1385889);
nand I_81315 (I1385954,I1385759,I1385937);
nand I_81316 (I1385685,I1385821,I1385937);
DFFARX1 I_81317 (I1385855,I3563,I1385708,I1385700,);
not I_81318 (I1385999,I1220491);
nor I_81319 (I1386016,I1385999,I1220476);
nor I_81320 (I1386033,I1386016,I1385838);
DFFARX1 I_81321 (I1386033,I3563,I1385708,I1385697,);
not I_81322 (I1386064,I1386016);
DFFARX1 I_81323 (I1386064,I3563,I1385708,I1386090,);
not I_81324 (I1386098,I1386090);
nor I_81325 (I1385694,I1386098,I1386016);
nor I_81326 (I1386129,I1385999,I1220485);
and I_81327 (I1386146,I1386129,I1220488);
or I_81328 (I1386163,I1386146,I1220470);
DFFARX1 I_81329 (I1386163,I3563,I1385708,I1386189,);
not I_81330 (I1386197,I1386189);
nand I_81331 (I1386214,I1386197,I1385937);
not I_81332 (I1385688,I1386214);
nand I_81333 (I1385682,I1386214,I1385954);
nand I_81334 (I1385679,I1386197,I1385821);
not I_81335 (I1386303,I3570);
DFFARX1 I_81336 (I26099,I3563,I1386303,I1386329,);
DFFARX1 I_81337 (I26081,I3563,I1386303,I1386346,);
not I_81338 (I1386354,I1386346);
nor I_81339 (I1386271,I1386329,I1386354);
DFFARX1 I_81340 (I1386354,I3563,I1386303,I1386286,);
nor I_81341 (I1386399,I26081,I26096);
and I_81342 (I1386416,I1386399,I26090);
nor I_81343 (I1386433,I1386416,I26081);
not I_81344 (I1386450,I26081);
and I_81345 (I1386467,I1386450,I26084);
nand I_81346 (I1386484,I1386467,I26087);
nor I_81347 (I1386501,I1386450,I1386484);
DFFARX1 I_81348 (I1386501,I3563,I1386303,I1386268,);
not I_81349 (I1386532,I1386484);
nand I_81350 (I1386549,I1386354,I1386532);
nand I_81351 (I1386280,I1386416,I1386532);
DFFARX1 I_81352 (I1386450,I3563,I1386303,I1386295,);
not I_81353 (I1386594,I26093);
nor I_81354 (I1386611,I1386594,I26084);
nor I_81355 (I1386628,I1386611,I1386433);
DFFARX1 I_81356 (I1386628,I3563,I1386303,I1386292,);
not I_81357 (I1386659,I1386611);
DFFARX1 I_81358 (I1386659,I3563,I1386303,I1386685,);
not I_81359 (I1386693,I1386685);
nor I_81360 (I1386289,I1386693,I1386611);
nor I_81361 (I1386724,I1386594,I26105);
and I_81362 (I1386741,I1386724,I26102);
or I_81363 (I1386758,I1386741,I26084);
DFFARX1 I_81364 (I1386758,I3563,I1386303,I1386784,);
not I_81365 (I1386792,I1386784);
nand I_81366 (I1386809,I1386792,I1386532);
not I_81367 (I1386283,I1386809);
nand I_81368 (I1386277,I1386809,I1386549);
nand I_81369 (I1386274,I1386792,I1386416);
not I_81370 (I1386898,I3570);
DFFARX1 I_81371 (I566171,I3563,I1386898,I1386924,);
DFFARX1 I_81372 (I566174,I3563,I1386898,I1386941,);
not I_81373 (I1386949,I1386941);
nor I_81374 (I1386866,I1386924,I1386949);
DFFARX1 I_81375 (I1386949,I3563,I1386898,I1386881,);
nor I_81376 (I1386994,I566177,I566195);
and I_81377 (I1387011,I1386994,I566180);
nor I_81378 (I1387028,I1387011,I566177);
not I_81379 (I1387045,I566177);
and I_81380 (I1387062,I1387045,I566189);
nand I_81381 (I1387079,I1387062,I566192);
nor I_81382 (I1387096,I1387045,I1387079);
DFFARX1 I_81383 (I1387096,I3563,I1386898,I1386863,);
not I_81384 (I1387127,I1387079);
nand I_81385 (I1387144,I1386949,I1387127);
nand I_81386 (I1386875,I1387011,I1387127);
DFFARX1 I_81387 (I1387045,I3563,I1386898,I1386890,);
not I_81388 (I1387189,I566183);
nor I_81389 (I1387206,I1387189,I566189);
nor I_81390 (I1387223,I1387206,I1387028);
DFFARX1 I_81391 (I1387223,I3563,I1386898,I1386887,);
not I_81392 (I1387254,I1387206);
DFFARX1 I_81393 (I1387254,I3563,I1386898,I1387280,);
not I_81394 (I1387288,I1387280);
nor I_81395 (I1386884,I1387288,I1387206);
nor I_81396 (I1387319,I1387189,I566171);
and I_81397 (I1387336,I1387319,I566186);
or I_81398 (I1387353,I1387336,I566174);
DFFARX1 I_81399 (I1387353,I3563,I1386898,I1387379,);
not I_81400 (I1387387,I1387379);
nand I_81401 (I1387404,I1387387,I1387127);
not I_81402 (I1386878,I1387404);
nand I_81403 (I1386872,I1387404,I1387144);
nand I_81404 (I1386869,I1387387,I1387011);
not I_81405 (I1387493,I3570);
DFFARX1 I_81406 (I434370,I3563,I1387493,I1387519,);
DFFARX1 I_81407 (I434376,I3563,I1387493,I1387536,);
not I_81408 (I1387544,I1387536);
nor I_81409 (I1387461,I1387519,I1387544);
DFFARX1 I_81410 (I1387544,I3563,I1387493,I1387476,);
nor I_81411 (I1387589,I434385,I434370);
and I_81412 (I1387606,I1387589,I434397);
nor I_81413 (I1387623,I1387606,I434385);
not I_81414 (I1387640,I434385);
and I_81415 (I1387657,I1387640,I434373);
nand I_81416 (I1387674,I1387657,I434394);
nor I_81417 (I1387691,I1387640,I1387674);
DFFARX1 I_81418 (I1387691,I3563,I1387493,I1387458,);
not I_81419 (I1387722,I1387674);
nand I_81420 (I1387739,I1387544,I1387722);
nand I_81421 (I1387470,I1387606,I1387722);
DFFARX1 I_81422 (I1387640,I3563,I1387493,I1387485,);
not I_81423 (I1387784,I434382);
nor I_81424 (I1387801,I1387784,I434373);
nor I_81425 (I1387818,I1387801,I1387623);
DFFARX1 I_81426 (I1387818,I3563,I1387493,I1387482,);
not I_81427 (I1387849,I1387801);
DFFARX1 I_81428 (I1387849,I3563,I1387493,I1387875,);
not I_81429 (I1387883,I1387875);
nor I_81430 (I1387479,I1387883,I1387801);
nor I_81431 (I1387914,I1387784,I434379);
and I_81432 (I1387931,I1387914,I434391);
or I_81433 (I1387948,I1387931,I434388);
DFFARX1 I_81434 (I1387948,I3563,I1387493,I1387974,);
not I_81435 (I1387982,I1387974);
nand I_81436 (I1387999,I1387982,I1387722);
not I_81437 (I1387473,I1387999);
nand I_81438 (I1387467,I1387999,I1387739);
nand I_81439 (I1387464,I1387982,I1387606);
not I_81440 (I1388088,I3570);
DFFARX1 I_81441 (I301196,I3563,I1388088,I1388114,);
DFFARX1 I_81442 (I301190,I3563,I1388088,I1388131,);
not I_81443 (I1388139,I1388131);
nor I_81444 (I1388056,I1388114,I1388139);
DFFARX1 I_81445 (I1388139,I3563,I1388088,I1388071,);
nor I_81446 (I1388184,I301178,I301199);
and I_81447 (I1388201,I1388184,I301193);
nor I_81448 (I1388218,I1388201,I301178);
not I_81449 (I1388235,I301178);
and I_81450 (I1388252,I1388235,I301175);
nand I_81451 (I1388269,I1388252,I301187);
nor I_81452 (I1388286,I1388235,I1388269);
DFFARX1 I_81453 (I1388286,I3563,I1388088,I1388053,);
not I_81454 (I1388317,I1388269);
nand I_81455 (I1388334,I1388139,I1388317);
nand I_81456 (I1388065,I1388201,I1388317);
DFFARX1 I_81457 (I1388235,I3563,I1388088,I1388080,);
not I_81458 (I1388379,I301202);
nor I_81459 (I1388396,I1388379,I301175);
nor I_81460 (I1388413,I1388396,I1388218);
DFFARX1 I_81461 (I1388413,I3563,I1388088,I1388077,);
not I_81462 (I1388444,I1388396);
DFFARX1 I_81463 (I1388444,I3563,I1388088,I1388470,);
not I_81464 (I1388478,I1388470);
nor I_81465 (I1388074,I1388478,I1388396);
nor I_81466 (I1388509,I1388379,I301184);
and I_81467 (I1388526,I1388509,I301181);
or I_81468 (I1388543,I1388526,I301175);
DFFARX1 I_81469 (I1388543,I3563,I1388088,I1388569,);
not I_81470 (I1388577,I1388569);
nand I_81471 (I1388594,I1388577,I1388317);
not I_81472 (I1388068,I1388594);
nand I_81473 (I1388062,I1388594,I1388334);
nand I_81474 (I1388059,I1388577,I1388201);
not I_81475 (I1388683,I3570);
DFFARX1 I_81476 (I420298,I3563,I1388683,I1388709,);
DFFARX1 I_81477 (I420292,I3563,I1388683,I1388726,);
not I_81478 (I1388734,I1388726);
nor I_81479 (I1388651,I1388709,I1388734);
DFFARX1 I_81480 (I1388734,I3563,I1388683,I1388666,);
nor I_81481 (I1388779,I420280,I420301);
and I_81482 (I1388796,I1388779,I420295);
nor I_81483 (I1388813,I1388796,I420280);
not I_81484 (I1388830,I420280);
and I_81485 (I1388847,I1388830,I420277);
nand I_81486 (I1388864,I1388847,I420289);
nor I_81487 (I1388881,I1388830,I1388864);
DFFARX1 I_81488 (I1388881,I3563,I1388683,I1388648,);
not I_81489 (I1388912,I1388864);
nand I_81490 (I1388929,I1388734,I1388912);
nand I_81491 (I1388660,I1388796,I1388912);
DFFARX1 I_81492 (I1388830,I3563,I1388683,I1388675,);
not I_81493 (I1388974,I420304);
nor I_81494 (I1388991,I1388974,I420277);
nor I_81495 (I1389008,I1388991,I1388813);
DFFARX1 I_81496 (I1389008,I3563,I1388683,I1388672,);
not I_81497 (I1389039,I1388991);
DFFARX1 I_81498 (I1389039,I3563,I1388683,I1389065,);
not I_81499 (I1389073,I1389065);
nor I_81500 (I1388669,I1389073,I1388991);
nor I_81501 (I1389104,I1388974,I420286);
and I_81502 (I1389121,I1389104,I420283);
or I_81503 (I1389138,I1389121,I420277);
DFFARX1 I_81504 (I1389138,I3563,I1388683,I1389164,);
not I_81505 (I1389172,I1389164);
nand I_81506 (I1389189,I1389172,I1388912);
not I_81507 (I1388663,I1389189);
nand I_81508 (I1388657,I1389189,I1388929);
nand I_81509 (I1388654,I1389172,I1388796);
not I_81510 (I1389278,I3570);
DFFARX1 I_81511 (I830037,I3563,I1389278,I1389304,);
DFFARX1 I_81512 (I830034,I3563,I1389278,I1389321,);
not I_81513 (I1389329,I1389321);
nor I_81514 (I1389246,I1389304,I1389329);
DFFARX1 I_81515 (I1389329,I3563,I1389278,I1389261,);
nor I_81516 (I1389374,I830049,I830031);
and I_81517 (I1389391,I1389374,I830028);
nor I_81518 (I1389408,I1389391,I830049);
not I_81519 (I1389425,I830049);
and I_81520 (I1389442,I1389425,I830034);
nand I_81521 (I1389459,I1389442,I830046);
nor I_81522 (I1389476,I1389425,I1389459);
DFFARX1 I_81523 (I1389476,I3563,I1389278,I1389243,);
not I_81524 (I1389507,I1389459);
nand I_81525 (I1389524,I1389329,I1389507);
nand I_81526 (I1389255,I1389391,I1389507);
DFFARX1 I_81527 (I1389425,I3563,I1389278,I1389270,);
not I_81528 (I1389569,I830040);
nor I_81529 (I1389586,I1389569,I830034);
nor I_81530 (I1389603,I1389586,I1389408);
DFFARX1 I_81531 (I1389603,I3563,I1389278,I1389267,);
not I_81532 (I1389634,I1389586);
DFFARX1 I_81533 (I1389634,I3563,I1389278,I1389660,);
not I_81534 (I1389668,I1389660);
nor I_81535 (I1389264,I1389668,I1389586);
nor I_81536 (I1389699,I1389569,I830028);
and I_81537 (I1389716,I1389699,I830043);
or I_81538 (I1389733,I1389716,I830031);
DFFARX1 I_81539 (I1389733,I3563,I1389278,I1389759,);
not I_81540 (I1389767,I1389759);
nand I_81541 (I1389784,I1389767,I1389507);
not I_81542 (I1389258,I1389784);
nand I_81543 (I1389252,I1389784,I1389524);
nand I_81544 (I1389249,I1389767,I1389391);
not I_81545 (I1389873,I3570);
DFFARX1 I_81546 (I910668,I3563,I1389873,I1389899,);
DFFARX1 I_81547 (I910665,I3563,I1389873,I1389916,);
not I_81548 (I1389924,I1389916);
nor I_81549 (I1389841,I1389899,I1389924);
DFFARX1 I_81550 (I1389924,I3563,I1389873,I1389856,);
nor I_81551 (I1389969,I910680,I910662);
and I_81552 (I1389986,I1389969,I910659);
nor I_81553 (I1390003,I1389986,I910680);
not I_81554 (I1390020,I910680);
and I_81555 (I1390037,I1390020,I910665);
nand I_81556 (I1390054,I1390037,I910677);
nor I_81557 (I1390071,I1390020,I1390054);
DFFARX1 I_81558 (I1390071,I3563,I1389873,I1389838,);
not I_81559 (I1390102,I1390054);
nand I_81560 (I1390119,I1389924,I1390102);
nand I_81561 (I1389850,I1389986,I1390102);
DFFARX1 I_81562 (I1390020,I3563,I1389873,I1389865,);
not I_81563 (I1390164,I910671);
nor I_81564 (I1390181,I1390164,I910665);
nor I_81565 (I1390198,I1390181,I1390003);
DFFARX1 I_81566 (I1390198,I3563,I1389873,I1389862,);
not I_81567 (I1390229,I1390181);
DFFARX1 I_81568 (I1390229,I3563,I1389873,I1390255,);
not I_81569 (I1390263,I1390255);
nor I_81570 (I1389859,I1390263,I1390181);
nor I_81571 (I1390294,I1390164,I910659);
and I_81572 (I1390311,I1390294,I910674);
or I_81573 (I1390328,I1390311,I910662);
DFFARX1 I_81574 (I1390328,I3563,I1389873,I1390354,);
not I_81575 (I1390362,I1390354);
nand I_81576 (I1390379,I1390362,I1390102);
not I_81577 (I1389853,I1390379);
nand I_81578 (I1389847,I1390379,I1390119);
nand I_81579 (I1389844,I1390362,I1389986);
not I_81580 (I1390468,I3570);
DFFARX1 I_81581 (I717968,I3563,I1390468,I1390494,);
DFFARX1 I_81582 (I717950,I3563,I1390468,I1390511,);
not I_81583 (I1390519,I1390511);
nor I_81584 (I1390436,I1390494,I1390519);
DFFARX1 I_81585 (I1390519,I3563,I1390468,I1390451,);
nor I_81586 (I1390564,I717956,I717959);
and I_81587 (I1390581,I1390564,I717947);
nor I_81588 (I1390598,I1390581,I717956);
not I_81589 (I1390615,I717956);
and I_81590 (I1390632,I1390615,I717965);
nand I_81591 (I1390649,I1390632,I717953);
nor I_81592 (I1390666,I1390615,I1390649);
DFFARX1 I_81593 (I1390666,I3563,I1390468,I1390433,);
not I_81594 (I1390697,I1390649);
nand I_81595 (I1390714,I1390519,I1390697);
nand I_81596 (I1390445,I1390581,I1390697);
DFFARX1 I_81597 (I1390615,I3563,I1390468,I1390460,);
not I_81598 (I1390759,I717950);
nor I_81599 (I1390776,I1390759,I717965);
nor I_81600 (I1390793,I1390776,I1390598);
DFFARX1 I_81601 (I1390793,I3563,I1390468,I1390457,);
not I_81602 (I1390824,I1390776);
DFFARX1 I_81603 (I1390824,I3563,I1390468,I1390850,);
not I_81604 (I1390858,I1390850);
nor I_81605 (I1390454,I1390858,I1390776);
nor I_81606 (I1390889,I1390759,I717962);
and I_81607 (I1390906,I1390889,I717971);
or I_81608 (I1390923,I1390906,I717947);
DFFARX1 I_81609 (I1390923,I3563,I1390468,I1390949,);
not I_81610 (I1390957,I1390949);
nand I_81611 (I1390974,I1390957,I1390697);
not I_81612 (I1390448,I1390974);
nand I_81613 (I1390442,I1390974,I1390714);
nand I_81614 (I1390439,I1390957,I1390581);
not I_81615 (I1391063,I3570);
DFFARX1 I_81616 (I884845,I3563,I1391063,I1391089,);
DFFARX1 I_81617 (I884842,I3563,I1391063,I1391106,);
not I_81618 (I1391114,I1391106);
nor I_81619 (I1391031,I1391089,I1391114);
DFFARX1 I_81620 (I1391114,I3563,I1391063,I1391046,);
nor I_81621 (I1391159,I884857,I884839);
and I_81622 (I1391176,I1391159,I884836);
nor I_81623 (I1391193,I1391176,I884857);
not I_81624 (I1391210,I884857);
and I_81625 (I1391227,I1391210,I884842);
nand I_81626 (I1391244,I1391227,I884854);
nor I_81627 (I1391261,I1391210,I1391244);
DFFARX1 I_81628 (I1391261,I3563,I1391063,I1391028,);
not I_81629 (I1391292,I1391244);
nand I_81630 (I1391309,I1391114,I1391292);
nand I_81631 (I1391040,I1391176,I1391292);
DFFARX1 I_81632 (I1391210,I3563,I1391063,I1391055,);
not I_81633 (I1391354,I884848);
nor I_81634 (I1391371,I1391354,I884842);
nor I_81635 (I1391388,I1391371,I1391193);
DFFARX1 I_81636 (I1391388,I3563,I1391063,I1391052,);
not I_81637 (I1391419,I1391371);
DFFARX1 I_81638 (I1391419,I3563,I1391063,I1391445,);
not I_81639 (I1391453,I1391445);
nor I_81640 (I1391049,I1391453,I1391371);
nor I_81641 (I1391484,I1391354,I884836);
and I_81642 (I1391501,I1391484,I884851);
or I_81643 (I1391518,I1391501,I884839);
DFFARX1 I_81644 (I1391518,I3563,I1391063,I1391544,);
not I_81645 (I1391552,I1391544);
nand I_81646 (I1391569,I1391552,I1391292);
not I_81647 (I1391043,I1391569);
nand I_81648 (I1391037,I1391569,I1391309);
nand I_81649 (I1391034,I1391552,I1391176);
not I_81650 (I1391658,I3570);
DFFARX1 I_81651 (I504546,I3563,I1391658,I1391684,);
DFFARX1 I_81652 (I504552,I3563,I1391658,I1391701,);
not I_81653 (I1391709,I1391701);
nor I_81654 (I1391626,I1391684,I1391709);
DFFARX1 I_81655 (I1391709,I3563,I1391658,I1391641,);
nor I_81656 (I1391754,I504561,I504546);
and I_81657 (I1391771,I1391754,I504573);
nor I_81658 (I1391788,I1391771,I504561);
not I_81659 (I1391805,I504561);
and I_81660 (I1391822,I1391805,I504549);
nand I_81661 (I1391839,I1391822,I504570);
nor I_81662 (I1391856,I1391805,I1391839);
DFFARX1 I_81663 (I1391856,I3563,I1391658,I1391623,);
not I_81664 (I1391887,I1391839);
nand I_81665 (I1391904,I1391709,I1391887);
nand I_81666 (I1391635,I1391771,I1391887);
DFFARX1 I_81667 (I1391805,I3563,I1391658,I1391650,);
not I_81668 (I1391949,I504558);
nor I_81669 (I1391966,I1391949,I504549);
nor I_81670 (I1391983,I1391966,I1391788);
DFFARX1 I_81671 (I1391983,I3563,I1391658,I1391647,);
not I_81672 (I1392014,I1391966);
DFFARX1 I_81673 (I1392014,I3563,I1391658,I1392040,);
not I_81674 (I1392048,I1392040);
nor I_81675 (I1391644,I1392048,I1391966);
nor I_81676 (I1392079,I1391949,I504555);
and I_81677 (I1392096,I1392079,I504567);
or I_81678 (I1392113,I1392096,I504564);
DFFARX1 I_81679 (I1392113,I3563,I1391658,I1392139,);
not I_81680 (I1392147,I1392139);
nand I_81681 (I1392164,I1392147,I1391887);
not I_81682 (I1391638,I1392164);
nand I_81683 (I1391632,I1392164,I1391904);
nand I_81684 (I1391629,I1392147,I1391771);
not I_81685 (I1392253,I3570);
DFFARX1 I_81686 (I47706,I3563,I1392253,I1392279,);
DFFARX1 I_81687 (I47688,I3563,I1392253,I1392296,);
not I_81688 (I1392304,I1392296);
nor I_81689 (I1392221,I1392279,I1392304);
DFFARX1 I_81690 (I1392304,I3563,I1392253,I1392236,);
nor I_81691 (I1392349,I47688,I47703);
and I_81692 (I1392366,I1392349,I47697);
nor I_81693 (I1392383,I1392366,I47688);
not I_81694 (I1392400,I47688);
and I_81695 (I1392417,I1392400,I47691);
nand I_81696 (I1392434,I1392417,I47694);
nor I_81697 (I1392451,I1392400,I1392434);
DFFARX1 I_81698 (I1392451,I3563,I1392253,I1392218,);
not I_81699 (I1392482,I1392434);
nand I_81700 (I1392499,I1392304,I1392482);
nand I_81701 (I1392230,I1392366,I1392482);
DFFARX1 I_81702 (I1392400,I3563,I1392253,I1392245,);
not I_81703 (I1392544,I47700);
nor I_81704 (I1392561,I1392544,I47691);
nor I_81705 (I1392578,I1392561,I1392383);
DFFARX1 I_81706 (I1392578,I3563,I1392253,I1392242,);
not I_81707 (I1392609,I1392561);
DFFARX1 I_81708 (I1392609,I3563,I1392253,I1392635,);
not I_81709 (I1392643,I1392635);
nor I_81710 (I1392239,I1392643,I1392561);
nor I_81711 (I1392674,I1392544,I47712);
and I_81712 (I1392691,I1392674,I47709);
or I_81713 (I1392708,I1392691,I47691);
DFFARX1 I_81714 (I1392708,I3563,I1392253,I1392734,);
not I_81715 (I1392742,I1392734);
nand I_81716 (I1392759,I1392742,I1392482);
not I_81717 (I1392233,I1392759);
nand I_81718 (I1392227,I1392759,I1392499);
nand I_81719 (I1392224,I1392742,I1392366);
not I_81720 (I1392848,I3570);
DFFARX1 I_81721 (I272003,I3563,I1392848,I1392874,);
DFFARX1 I_81722 (I272006,I3563,I1392848,I1392891,);
not I_81723 (I1392899,I1392891);
nor I_81724 (I1392816,I1392874,I1392899);
DFFARX1 I_81725 (I1392899,I3563,I1392848,I1392831,);
nor I_81726 (I1392944,I272012,I272006);
and I_81727 (I1392961,I1392944,I272009);
nor I_81728 (I1392978,I1392961,I272012);
not I_81729 (I1392995,I272012);
and I_81730 (I1393012,I1392995,I272003);
nand I_81731 (I1393029,I1393012,I272021);
nor I_81732 (I1393046,I1392995,I1393029);
DFFARX1 I_81733 (I1393046,I3563,I1392848,I1392813,);
not I_81734 (I1393077,I1393029);
nand I_81735 (I1393094,I1392899,I1393077);
nand I_81736 (I1392825,I1392961,I1393077);
DFFARX1 I_81737 (I1392995,I3563,I1392848,I1392840,);
not I_81738 (I1393139,I272015);
nor I_81739 (I1393156,I1393139,I272003);
nor I_81740 (I1393173,I1393156,I1392978);
DFFARX1 I_81741 (I1393173,I3563,I1392848,I1392837,);
not I_81742 (I1393204,I1393156);
DFFARX1 I_81743 (I1393204,I3563,I1392848,I1393230,);
not I_81744 (I1393238,I1393230);
nor I_81745 (I1392834,I1393238,I1393156);
nor I_81746 (I1393269,I1393139,I272018);
and I_81747 (I1393286,I1393269,I272024);
or I_81748 (I1393303,I1393286,I272027);
DFFARX1 I_81749 (I1393303,I3563,I1392848,I1393329,);
not I_81750 (I1393337,I1393329);
nand I_81751 (I1393354,I1393337,I1393077);
not I_81752 (I1392828,I1393354);
nand I_81753 (I1392822,I1393354,I1393094);
nand I_81754 (I1392819,I1393337,I1392961);
not I_81755 (I1393443,I3570);
DFFARX1 I_81756 (I371287,I3563,I1393443,I1393469,);
DFFARX1 I_81757 (I371281,I3563,I1393443,I1393486,);
not I_81758 (I1393494,I1393486);
nor I_81759 (I1393411,I1393469,I1393494);
DFFARX1 I_81760 (I1393494,I3563,I1393443,I1393426,);
nor I_81761 (I1393539,I371269,I371290);
and I_81762 (I1393556,I1393539,I371284);
nor I_81763 (I1393573,I1393556,I371269);
not I_81764 (I1393590,I371269);
and I_81765 (I1393607,I1393590,I371266);
nand I_81766 (I1393624,I1393607,I371278);
nor I_81767 (I1393641,I1393590,I1393624);
DFFARX1 I_81768 (I1393641,I3563,I1393443,I1393408,);
not I_81769 (I1393672,I1393624);
nand I_81770 (I1393689,I1393494,I1393672);
nand I_81771 (I1393420,I1393556,I1393672);
DFFARX1 I_81772 (I1393590,I3563,I1393443,I1393435,);
not I_81773 (I1393734,I371293);
nor I_81774 (I1393751,I1393734,I371266);
nor I_81775 (I1393768,I1393751,I1393573);
DFFARX1 I_81776 (I1393768,I3563,I1393443,I1393432,);
not I_81777 (I1393799,I1393751);
DFFARX1 I_81778 (I1393799,I3563,I1393443,I1393825,);
not I_81779 (I1393833,I1393825);
nor I_81780 (I1393429,I1393833,I1393751);
nor I_81781 (I1393864,I1393734,I371275);
and I_81782 (I1393881,I1393864,I371272);
or I_81783 (I1393898,I1393881,I371266);
DFFARX1 I_81784 (I1393898,I3563,I1393443,I1393924,);
not I_81785 (I1393932,I1393924);
nand I_81786 (I1393949,I1393932,I1393672);
not I_81787 (I1393423,I1393949);
nand I_81788 (I1393417,I1393949,I1393689);
nand I_81789 (I1393414,I1393932,I1393556);
not I_81790 (I1394038,I3570);
DFFARX1 I_81791 (I68262,I3563,I1394038,I1394064,);
DFFARX1 I_81792 (I68250,I3563,I1394038,I1394081,);
not I_81793 (I1394089,I1394081);
nor I_81794 (I1394006,I1394064,I1394089);
DFFARX1 I_81795 (I1394089,I3563,I1394038,I1394021,);
nor I_81796 (I1394134,I68241,I68265);
and I_81797 (I1394151,I1394134,I68244);
nor I_81798 (I1394168,I1394151,I68241);
not I_81799 (I1394185,I68241);
and I_81800 (I1394202,I1394185,I68247);
nand I_81801 (I1394219,I1394202,I68259);
nor I_81802 (I1394236,I1394185,I1394219);
DFFARX1 I_81803 (I1394236,I3563,I1394038,I1394003,);
not I_81804 (I1394267,I1394219);
nand I_81805 (I1394284,I1394089,I1394267);
nand I_81806 (I1394015,I1394151,I1394267);
DFFARX1 I_81807 (I1394185,I3563,I1394038,I1394030,);
not I_81808 (I1394329,I68241);
nor I_81809 (I1394346,I1394329,I68247);
nor I_81810 (I1394363,I1394346,I1394168);
DFFARX1 I_81811 (I1394363,I3563,I1394038,I1394027,);
not I_81812 (I1394394,I1394346);
DFFARX1 I_81813 (I1394394,I3563,I1394038,I1394420,);
not I_81814 (I1394428,I1394420);
nor I_81815 (I1394024,I1394428,I1394346);
nor I_81816 (I1394459,I1394329,I68244);
and I_81817 (I1394476,I1394459,I68253);
or I_81818 (I1394493,I1394476,I68256);
DFFARX1 I_81819 (I1394493,I3563,I1394038,I1394519,);
not I_81820 (I1394527,I1394519);
nand I_81821 (I1394544,I1394527,I1394267);
not I_81822 (I1394018,I1394544);
nand I_81823 (I1394012,I1394544,I1394284);
nand I_81824 (I1394009,I1394527,I1394151);
not I_81825 (I1394633,I3570);
DFFARX1 I_81826 (I548321,I3563,I1394633,I1394659,);
DFFARX1 I_81827 (I548324,I3563,I1394633,I1394676,);
not I_81828 (I1394684,I1394676);
nor I_81829 (I1394601,I1394659,I1394684);
DFFARX1 I_81830 (I1394684,I3563,I1394633,I1394616,);
nor I_81831 (I1394729,I548327,I548345);
and I_81832 (I1394746,I1394729,I548330);
nor I_81833 (I1394763,I1394746,I548327);
not I_81834 (I1394780,I548327);
and I_81835 (I1394797,I1394780,I548339);
nand I_81836 (I1394814,I1394797,I548342);
nor I_81837 (I1394831,I1394780,I1394814);
DFFARX1 I_81838 (I1394831,I3563,I1394633,I1394598,);
not I_81839 (I1394862,I1394814);
nand I_81840 (I1394879,I1394684,I1394862);
nand I_81841 (I1394610,I1394746,I1394862);
DFFARX1 I_81842 (I1394780,I3563,I1394633,I1394625,);
not I_81843 (I1394924,I548333);
nor I_81844 (I1394941,I1394924,I548339);
nor I_81845 (I1394958,I1394941,I1394763);
DFFARX1 I_81846 (I1394958,I3563,I1394633,I1394622,);
not I_81847 (I1394989,I1394941);
DFFARX1 I_81848 (I1394989,I3563,I1394633,I1395015,);
not I_81849 (I1395023,I1395015);
nor I_81850 (I1394619,I1395023,I1394941);
nor I_81851 (I1395054,I1394924,I548321);
and I_81852 (I1395071,I1395054,I548336);
or I_81853 (I1395088,I1395071,I548324);
DFFARX1 I_81854 (I1395088,I3563,I1394633,I1395114,);
not I_81855 (I1395122,I1395114);
nand I_81856 (I1395139,I1395122,I1394862);
not I_81857 (I1394613,I1395139);
nand I_81858 (I1394607,I1395139,I1394879);
nand I_81859 (I1394604,I1395122,I1394746);
not I_81860 (I1395228,I3570);
DFFARX1 I_81861 (I463202,I3563,I1395228,I1395254,);
DFFARX1 I_81862 (I463208,I3563,I1395228,I1395271,);
not I_81863 (I1395279,I1395271);
nor I_81864 (I1395196,I1395254,I1395279);
DFFARX1 I_81865 (I1395279,I3563,I1395228,I1395211,);
nor I_81866 (I1395324,I463217,I463202);
and I_81867 (I1395341,I1395324,I463229);
nor I_81868 (I1395358,I1395341,I463217);
not I_81869 (I1395375,I463217);
and I_81870 (I1395392,I1395375,I463205);
nand I_81871 (I1395409,I1395392,I463226);
nor I_81872 (I1395426,I1395375,I1395409);
DFFARX1 I_81873 (I1395426,I3563,I1395228,I1395193,);
not I_81874 (I1395457,I1395409);
nand I_81875 (I1395474,I1395279,I1395457);
nand I_81876 (I1395205,I1395341,I1395457);
DFFARX1 I_81877 (I1395375,I3563,I1395228,I1395220,);
not I_81878 (I1395519,I463214);
nor I_81879 (I1395536,I1395519,I463205);
nor I_81880 (I1395553,I1395536,I1395358);
DFFARX1 I_81881 (I1395553,I3563,I1395228,I1395217,);
not I_81882 (I1395584,I1395536);
DFFARX1 I_81883 (I1395584,I3563,I1395228,I1395610,);
not I_81884 (I1395618,I1395610);
nor I_81885 (I1395214,I1395618,I1395536);
nor I_81886 (I1395649,I1395519,I463211);
and I_81887 (I1395666,I1395649,I463223);
or I_81888 (I1395683,I1395666,I463220);
DFFARX1 I_81889 (I1395683,I3563,I1395228,I1395709,);
not I_81890 (I1395717,I1395709);
nand I_81891 (I1395734,I1395717,I1395457);
not I_81892 (I1395208,I1395734);
nand I_81893 (I1395202,I1395734,I1395474);
nand I_81894 (I1395199,I1395717,I1395341);
not I_81895 (I1395823,I3570);
DFFARX1 I_81896 (I441442,I3563,I1395823,I1395849,);
DFFARX1 I_81897 (I441448,I3563,I1395823,I1395866,);
not I_81898 (I1395874,I1395866);
nor I_81899 (I1395791,I1395849,I1395874);
DFFARX1 I_81900 (I1395874,I3563,I1395823,I1395806,);
nor I_81901 (I1395919,I441457,I441442);
and I_81902 (I1395936,I1395919,I441469);
nor I_81903 (I1395953,I1395936,I441457);
not I_81904 (I1395970,I441457);
and I_81905 (I1395987,I1395970,I441445);
nand I_81906 (I1396004,I1395987,I441466);
nor I_81907 (I1396021,I1395970,I1396004);
DFFARX1 I_81908 (I1396021,I3563,I1395823,I1395788,);
not I_81909 (I1396052,I1396004);
nand I_81910 (I1396069,I1395874,I1396052);
nand I_81911 (I1395800,I1395936,I1396052);
DFFARX1 I_81912 (I1395970,I3563,I1395823,I1395815,);
not I_81913 (I1396114,I441454);
nor I_81914 (I1396131,I1396114,I441445);
nor I_81915 (I1396148,I1396131,I1395953);
DFFARX1 I_81916 (I1396148,I3563,I1395823,I1395812,);
not I_81917 (I1396179,I1396131);
DFFARX1 I_81918 (I1396179,I3563,I1395823,I1396205,);
not I_81919 (I1396213,I1396205);
nor I_81920 (I1395809,I1396213,I1396131);
nor I_81921 (I1396244,I1396114,I441451);
and I_81922 (I1396261,I1396244,I441463);
or I_81923 (I1396278,I1396261,I441460);
DFFARX1 I_81924 (I1396278,I3563,I1395823,I1396304,);
not I_81925 (I1396312,I1396304);
nand I_81926 (I1396329,I1396312,I1396052);
not I_81927 (I1395803,I1396329);
nand I_81928 (I1395797,I1396329,I1396069);
nand I_81929 (I1395794,I1396312,I1395936);
not I_81930 (I1396418,I3570);
DFFARX1 I_81931 (I561411,I3563,I1396418,I1396444,);
DFFARX1 I_81932 (I561414,I3563,I1396418,I1396461,);
not I_81933 (I1396469,I1396461);
nor I_81934 (I1396386,I1396444,I1396469);
DFFARX1 I_81935 (I1396469,I3563,I1396418,I1396401,);
nor I_81936 (I1396514,I561417,I561435);
and I_81937 (I1396531,I1396514,I561420);
nor I_81938 (I1396548,I1396531,I561417);
not I_81939 (I1396565,I561417);
and I_81940 (I1396582,I1396565,I561429);
nand I_81941 (I1396599,I1396582,I561432);
nor I_81942 (I1396616,I1396565,I1396599);
DFFARX1 I_81943 (I1396616,I3563,I1396418,I1396383,);
not I_81944 (I1396647,I1396599);
nand I_81945 (I1396664,I1396469,I1396647);
nand I_81946 (I1396395,I1396531,I1396647);
DFFARX1 I_81947 (I1396565,I3563,I1396418,I1396410,);
not I_81948 (I1396709,I561423);
nor I_81949 (I1396726,I1396709,I561429);
nor I_81950 (I1396743,I1396726,I1396548);
DFFARX1 I_81951 (I1396743,I3563,I1396418,I1396407,);
not I_81952 (I1396774,I1396726);
DFFARX1 I_81953 (I1396774,I3563,I1396418,I1396800,);
not I_81954 (I1396808,I1396800);
nor I_81955 (I1396404,I1396808,I1396726);
nor I_81956 (I1396839,I1396709,I561411);
and I_81957 (I1396856,I1396839,I561426);
or I_81958 (I1396873,I1396856,I561414);
DFFARX1 I_81959 (I1396873,I3563,I1396418,I1396899,);
not I_81960 (I1396907,I1396899);
nand I_81961 (I1396924,I1396907,I1396647);
not I_81962 (I1396398,I1396924);
nand I_81963 (I1396392,I1396924,I1396664);
nand I_81964 (I1396389,I1396907,I1396531);
not I_81965 (I1397013,I3570);
DFFARX1 I_81966 (I1291817,I3563,I1397013,I1397039,);
DFFARX1 I_81967 (I1291808,I3563,I1397013,I1397056,);
not I_81968 (I1397064,I1397056);
nor I_81969 (I1396981,I1397039,I1397064);
DFFARX1 I_81970 (I1397064,I3563,I1397013,I1396996,);
nor I_81971 (I1397109,I1291799,I1291814);
and I_81972 (I1397126,I1397109,I1291802);
nor I_81973 (I1397143,I1397126,I1291799);
not I_81974 (I1397160,I1291799);
and I_81975 (I1397177,I1397160,I1291805);
nand I_81976 (I1397194,I1397177,I1291823);
nor I_81977 (I1397211,I1397160,I1397194);
DFFARX1 I_81978 (I1397211,I3563,I1397013,I1396978,);
not I_81979 (I1397242,I1397194);
nand I_81980 (I1397259,I1397064,I1397242);
nand I_81981 (I1396990,I1397126,I1397242);
DFFARX1 I_81982 (I1397160,I3563,I1397013,I1397005,);
not I_81983 (I1397304,I1291799);
nor I_81984 (I1397321,I1397304,I1291805);
nor I_81985 (I1397338,I1397321,I1397143);
DFFARX1 I_81986 (I1397338,I3563,I1397013,I1397002,);
not I_81987 (I1397369,I1397321);
DFFARX1 I_81988 (I1397369,I3563,I1397013,I1397395,);
not I_81989 (I1397403,I1397395);
nor I_81990 (I1396999,I1397403,I1397321);
nor I_81991 (I1397434,I1397304,I1291802);
and I_81992 (I1397451,I1397434,I1291811);
or I_81993 (I1397468,I1397451,I1291820);
DFFARX1 I_81994 (I1397468,I3563,I1397013,I1397494,);
not I_81995 (I1397502,I1397494);
nand I_81996 (I1397519,I1397502,I1397242);
not I_81997 (I1396993,I1397519);
nand I_81998 (I1396987,I1397519,I1397259);
nand I_81999 (I1396984,I1397502,I1397126);
not I_82000 (I1397608,I3570);
DFFARX1 I_82001 (I240468,I3563,I1397608,I1397634,);
DFFARX1 I_82002 (I240471,I3563,I1397608,I1397651,);
not I_82003 (I1397659,I1397651);
nor I_82004 (I1397576,I1397634,I1397659);
DFFARX1 I_82005 (I1397659,I3563,I1397608,I1397591,);
nor I_82006 (I1397704,I240477,I240471);
and I_82007 (I1397721,I1397704,I240474);
nor I_82008 (I1397738,I1397721,I240477);
not I_82009 (I1397755,I240477);
and I_82010 (I1397772,I1397755,I240468);
nand I_82011 (I1397789,I1397772,I240486);
nor I_82012 (I1397806,I1397755,I1397789);
DFFARX1 I_82013 (I1397806,I3563,I1397608,I1397573,);
not I_82014 (I1397837,I1397789);
nand I_82015 (I1397854,I1397659,I1397837);
nand I_82016 (I1397585,I1397721,I1397837);
DFFARX1 I_82017 (I1397755,I3563,I1397608,I1397600,);
not I_82018 (I1397899,I240480);
nor I_82019 (I1397916,I1397899,I240468);
nor I_82020 (I1397933,I1397916,I1397738);
DFFARX1 I_82021 (I1397933,I3563,I1397608,I1397597,);
not I_82022 (I1397964,I1397916);
DFFARX1 I_82023 (I1397964,I3563,I1397608,I1397990,);
not I_82024 (I1397998,I1397990);
nor I_82025 (I1397594,I1397998,I1397916);
nor I_82026 (I1398029,I1397899,I240483);
and I_82027 (I1398046,I1398029,I240489);
or I_82028 (I1398063,I1398046,I240492);
DFFARX1 I_82029 (I1398063,I3563,I1397608,I1398089,);
not I_82030 (I1398097,I1398089);
nand I_82031 (I1398114,I1398097,I1397837);
not I_82032 (I1397588,I1398114);
nand I_82033 (I1397582,I1398114,I1397854);
nand I_82034 (I1397579,I1398097,I1397721);
not I_82035 (I1398203,I3570);
DFFARX1 I_82036 (I795420,I3563,I1398203,I1398229,);
DFFARX1 I_82037 (I795402,I3563,I1398203,I1398246,);
not I_82038 (I1398254,I1398246);
nor I_82039 (I1398171,I1398229,I1398254);
DFFARX1 I_82040 (I1398254,I3563,I1398203,I1398186,);
nor I_82041 (I1398299,I795408,I795411);
and I_82042 (I1398316,I1398299,I795399);
nor I_82043 (I1398333,I1398316,I795408);
not I_82044 (I1398350,I795408);
and I_82045 (I1398367,I1398350,I795417);
nand I_82046 (I1398384,I1398367,I795405);
nor I_82047 (I1398401,I1398350,I1398384);
DFFARX1 I_82048 (I1398401,I3563,I1398203,I1398168,);
not I_82049 (I1398432,I1398384);
nand I_82050 (I1398449,I1398254,I1398432);
nand I_82051 (I1398180,I1398316,I1398432);
DFFARX1 I_82052 (I1398350,I3563,I1398203,I1398195,);
not I_82053 (I1398494,I795402);
nor I_82054 (I1398511,I1398494,I795417);
nor I_82055 (I1398528,I1398511,I1398333);
DFFARX1 I_82056 (I1398528,I3563,I1398203,I1398192,);
not I_82057 (I1398559,I1398511);
DFFARX1 I_82058 (I1398559,I3563,I1398203,I1398585,);
not I_82059 (I1398593,I1398585);
nor I_82060 (I1398189,I1398593,I1398511);
nor I_82061 (I1398624,I1398494,I795414);
and I_82062 (I1398641,I1398624,I795423);
or I_82063 (I1398658,I1398641,I795399);
DFFARX1 I_82064 (I1398658,I3563,I1398203,I1398684,);
not I_82065 (I1398692,I1398684);
nand I_82066 (I1398709,I1398692,I1398432);
not I_82067 (I1398183,I1398709);
nand I_82068 (I1398177,I1398709,I1398449);
nand I_82069 (I1398174,I1398692,I1398316);
not I_82070 (I1398798,I3570);
DFFARX1 I_82071 (I1151110,I3563,I1398798,I1398824,);
DFFARX1 I_82072 (I1151122,I3563,I1398798,I1398841,);
not I_82073 (I1398849,I1398841);
nor I_82074 (I1398766,I1398824,I1398849);
DFFARX1 I_82075 (I1398849,I3563,I1398798,I1398781,);
nor I_82076 (I1398894,I1151119,I1151113);
and I_82077 (I1398911,I1398894,I1151107);
nor I_82078 (I1398928,I1398911,I1151119);
not I_82079 (I1398945,I1151119);
and I_82080 (I1398962,I1398945,I1151116);
nand I_82081 (I1398979,I1398962,I1151107);
nor I_82082 (I1398996,I1398945,I1398979);
DFFARX1 I_82083 (I1398996,I3563,I1398798,I1398763,);
not I_82084 (I1399027,I1398979);
nand I_82085 (I1399044,I1398849,I1399027);
nand I_82086 (I1398775,I1398911,I1399027);
DFFARX1 I_82087 (I1398945,I3563,I1398798,I1398790,);
not I_82088 (I1399089,I1151131);
nor I_82089 (I1399106,I1399089,I1151116);
nor I_82090 (I1399123,I1399106,I1398928);
DFFARX1 I_82091 (I1399123,I3563,I1398798,I1398787,);
not I_82092 (I1399154,I1399106);
DFFARX1 I_82093 (I1399154,I3563,I1398798,I1399180,);
not I_82094 (I1399188,I1399180);
nor I_82095 (I1398784,I1399188,I1399106);
nor I_82096 (I1399219,I1399089,I1151125);
and I_82097 (I1399236,I1399219,I1151128);
or I_82098 (I1399253,I1399236,I1151110);
DFFARX1 I_82099 (I1399253,I3563,I1398798,I1399279,);
not I_82100 (I1399287,I1399279);
nand I_82101 (I1399304,I1399287,I1399027);
not I_82102 (I1398778,I1399304);
nand I_82103 (I1398772,I1399304,I1399044);
nand I_82104 (I1398769,I1399287,I1398911);
not I_82105 (I1399393,I3570);
DFFARX1 I_82106 (I1302799,I3563,I1399393,I1399419,);
DFFARX1 I_82107 (I1302790,I3563,I1399393,I1399436,);
not I_82108 (I1399444,I1399436);
nor I_82109 (I1399361,I1399419,I1399444);
DFFARX1 I_82110 (I1399444,I3563,I1399393,I1399376,);
nor I_82111 (I1399489,I1302781,I1302796);
and I_82112 (I1399506,I1399489,I1302784);
nor I_82113 (I1399523,I1399506,I1302781);
not I_82114 (I1399540,I1302781);
and I_82115 (I1399557,I1399540,I1302787);
nand I_82116 (I1399574,I1399557,I1302805);
nor I_82117 (I1399591,I1399540,I1399574);
DFFARX1 I_82118 (I1399591,I3563,I1399393,I1399358,);
not I_82119 (I1399622,I1399574);
nand I_82120 (I1399639,I1399444,I1399622);
nand I_82121 (I1399370,I1399506,I1399622);
DFFARX1 I_82122 (I1399540,I3563,I1399393,I1399385,);
not I_82123 (I1399684,I1302781);
nor I_82124 (I1399701,I1399684,I1302787);
nor I_82125 (I1399718,I1399701,I1399523);
DFFARX1 I_82126 (I1399718,I3563,I1399393,I1399382,);
not I_82127 (I1399749,I1399701);
DFFARX1 I_82128 (I1399749,I3563,I1399393,I1399775,);
not I_82129 (I1399783,I1399775);
nor I_82130 (I1399379,I1399783,I1399701);
nor I_82131 (I1399814,I1399684,I1302784);
and I_82132 (I1399831,I1399814,I1302793);
or I_82133 (I1399848,I1399831,I1302802);
DFFARX1 I_82134 (I1399848,I3563,I1399393,I1399874,);
not I_82135 (I1399882,I1399874);
nand I_82136 (I1399899,I1399882,I1399622);
not I_82137 (I1399373,I1399899);
nand I_82138 (I1399367,I1399899,I1399639);
nand I_82139 (I1399364,I1399882,I1399506);
not I_82140 (I1399988,I3570);
DFFARX1 I_82141 (I571526,I3563,I1399988,I1400014,);
DFFARX1 I_82142 (I571529,I3563,I1399988,I1400031,);
not I_82143 (I1400039,I1400031);
nor I_82144 (I1399956,I1400014,I1400039);
DFFARX1 I_82145 (I1400039,I3563,I1399988,I1399971,);
nor I_82146 (I1400084,I571532,I571550);
and I_82147 (I1400101,I1400084,I571535);
nor I_82148 (I1400118,I1400101,I571532);
not I_82149 (I1400135,I571532);
and I_82150 (I1400152,I1400135,I571544);
nand I_82151 (I1400169,I1400152,I571547);
nor I_82152 (I1400186,I1400135,I1400169);
DFFARX1 I_82153 (I1400186,I3563,I1399988,I1399953,);
not I_82154 (I1400217,I1400169);
nand I_82155 (I1400234,I1400039,I1400217);
nand I_82156 (I1399965,I1400101,I1400217);
DFFARX1 I_82157 (I1400135,I3563,I1399988,I1399980,);
not I_82158 (I1400279,I571538);
nor I_82159 (I1400296,I1400279,I571544);
nor I_82160 (I1400313,I1400296,I1400118);
DFFARX1 I_82161 (I1400313,I3563,I1399988,I1399977,);
not I_82162 (I1400344,I1400296);
DFFARX1 I_82163 (I1400344,I3563,I1399988,I1400370,);
not I_82164 (I1400378,I1400370);
nor I_82165 (I1399974,I1400378,I1400296);
nor I_82166 (I1400409,I1400279,I571526);
and I_82167 (I1400426,I1400409,I571541);
or I_82168 (I1400443,I1400426,I571529);
DFFARX1 I_82169 (I1400443,I3563,I1399988,I1400469,);
not I_82170 (I1400477,I1400469);
nand I_82171 (I1400494,I1400477,I1400217);
not I_82172 (I1399968,I1400494);
nand I_82173 (I1399962,I1400494,I1400234);
nand I_82174 (I1399959,I1400477,I1400101);
not I_82175 (I1400583,I3570);
DFFARX1 I_82176 (I709876,I3563,I1400583,I1400609,);
DFFARX1 I_82177 (I709858,I3563,I1400583,I1400626,);
not I_82178 (I1400634,I1400626);
nor I_82179 (I1400551,I1400609,I1400634);
DFFARX1 I_82180 (I1400634,I3563,I1400583,I1400566,);
nor I_82181 (I1400679,I709864,I709867);
and I_82182 (I1400696,I1400679,I709855);
nor I_82183 (I1400713,I1400696,I709864);
not I_82184 (I1400730,I709864);
and I_82185 (I1400747,I1400730,I709873);
nand I_82186 (I1400764,I1400747,I709861);
nor I_82187 (I1400781,I1400730,I1400764);
DFFARX1 I_82188 (I1400781,I3563,I1400583,I1400548,);
not I_82189 (I1400812,I1400764);
nand I_82190 (I1400829,I1400634,I1400812);
nand I_82191 (I1400560,I1400696,I1400812);
DFFARX1 I_82192 (I1400730,I3563,I1400583,I1400575,);
not I_82193 (I1400874,I709858);
nor I_82194 (I1400891,I1400874,I709873);
nor I_82195 (I1400908,I1400891,I1400713);
DFFARX1 I_82196 (I1400908,I3563,I1400583,I1400572,);
not I_82197 (I1400939,I1400891);
DFFARX1 I_82198 (I1400939,I3563,I1400583,I1400965,);
not I_82199 (I1400973,I1400965);
nor I_82200 (I1400569,I1400973,I1400891);
nor I_82201 (I1401004,I1400874,I709870);
and I_82202 (I1401021,I1401004,I709879);
or I_82203 (I1401038,I1401021,I709855);
DFFARX1 I_82204 (I1401038,I3563,I1400583,I1401064,);
not I_82205 (I1401072,I1401064);
nand I_82206 (I1401089,I1401072,I1400812);
not I_82207 (I1400563,I1401089);
nand I_82208 (I1400557,I1401089,I1400829);
nand I_82209 (I1400554,I1401072,I1400696);
not I_82210 (I1401178,I3570);
DFFARX1 I_82211 (I443074,I3563,I1401178,I1401204,);
DFFARX1 I_82212 (I443080,I3563,I1401178,I1401221,);
not I_82213 (I1401229,I1401221);
nor I_82214 (I1401146,I1401204,I1401229);
DFFARX1 I_82215 (I1401229,I3563,I1401178,I1401161,);
nor I_82216 (I1401274,I443089,I443074);
and I_82217 (I1401291,I1401274,I443101);
nor I_82218 (I1401308,I1401291,I443089);
not I_82219 (I1401325,I443089);
and I_82220 (I1401342,I1401325,I443077);
nand I_82221 (I1401359,I1401342,I443098);
nor I_82222 (I1401376,I1401325,I1401359);
DFFARX1 I_82223 (I1401376,I3563,I1401178,I1401143,);
not I_82224 (I1401407,I1401359);
nand I_82225 (I1401424,I1401229,I1401407);
nand I_82226 (I1401155,I1401291,I1401407);
DFFARX1 I_82227 (I1401325,I3563,I1401178,I1401170,);
not I_82228 (I1401469,I443086);
nor I_82229 (I1401486,I1401469,I443077);
nor I_82230 (I1401503,I1401486,I1401308);
DFFARX1 I_82231 (I1401503,I3563,I1401178,I1401167,);
not I_82232 (I1401534,I1401486);
DFFARX1 I_82233 (I1401534,I3563,I1401178,I1401560,);
not I_82234 (I1401568,I1401560);
nor I_82235 (I1401164,I1401568,I1401486);
nor I_82236 (I1401599,I1401469,I443083);
and I_82237 (I1401616,I1401599,I443095);
or I_82238 (I1401633,I1401616,I443092);
DFFARX1 I_82239 (I1401633,I3563,I1401178,I1401659,);
not I_82240 (I1401667,I1401659);
nand I_82241 (I1401684,I1401667,I1401407);
not I_82242 (I1401158,I1401684);
nand I_82243 (I1401152,I1401684,I1401424);
nand I_82244 (I1401149,I1401667,I1401291);
not I_82245 (I1401773,I3570);
DFFARX1 I_82246 (I853752,I3563,I1401773,I1401799,);
DFFARX1 I_82247 (I853749,I3563,I1401773,I1401816,);
not I_82248 (I1401824,I1401816);
nor I_82249 (I1401741,I1401799,I1401824);
DFFARX1 I_82250 (I1401824,I3563,I1401773,I1401756,);
nor I_82251 (I1401869,I853764,I853746);
and I_82252 (I1401886,I1401869,I853743);
nor I_82253 (I1401903,I1401886,I853764);
not I_82254 (I1401920,I853764);
and I_82255 (I1401937,I1401920,I853749);
nand I_82256 (I1401954,I1401937,I853761);
nor I_82257 (I1401971,I1401920,I1401954);
DFFARX1 I_82258 (I1401971,I3563,I1401773,I1401738,);
not I_82259 (I1402002,I1401954);
nand I_82260 (I1402019,I1401824,I1402002);
nand I_82261 (I1401750,I1401886,I1402002);
DFFARX1 I_82262 (I1401920,I3563,I1401773,I1401765,);
not I_82263 (I1402064,I853755);
nor I_82264 (I1402081,I1402064,I853749);
nor I_82265 (I1402098,I1402081,I1401903);
DFFARX1 I_82266 (I1402098,I3563,I1401773,I1401762,);
not I_82267 (I1402129,I1402081);
DFFARX1 I_82268 (I1402129,I3563,I1401773,I1402155,);
not I_82269 (I1402163,I1402155);
nor I_82270 (I1401759,I1402163,I1402081);
nor I_82271 (I1402194,I1402064,I853743);
and I_82272 (I1402211,I1402194,I853758);
or I_82273 (I1402228,I1402211,I853746);
DFFARX1 I_82274 (I1402228,I3563,I1401773,I1402254,);
not I_82275 (I1402262,I1402254);
nand I_82276 (I1402279,I1402262,I1402002);
not I_82277 (I1401753,I1402279);
nand I_82278 (I1401747,I1402279,I1402019);
nand I_82279 (I1401744,I1402262,I1401886);
not I_82280 (I1402368,I3570);
DFFARX1 I_82281 (I936845,I3563,I1402368,I1402394,);
DFFARX1 I_82282 (I936863,I3563,I1402368,I1402411,);
not I_82283 (I1402419,I1402411);
nor I_82284 (I1402336,I1402394,I1402419);
DFFARX1 I_82285 (I1402419,I3563,I1402368,I1402351,);
nor I_82286 (I1402464,I936842,I936854);
and I_82287 (I1402481,I1402464,I936839);
nor I_82288 (I1402498,I1402481,I936842);
not I_82289 (I1402515,I936842);
and I_82290 (I1402532,I1402515,I936848);
nand I_82291 (I1402549,I1402532,I936860);
nor I_82292 (I1402566,I1402515,I1402549);
DFFARX1 I_82293 (I1402566,I3563,I1402368,I1402333,);
not I_82294 (I1402597,I1402549);
nand I_82295 (I1402614,I1402419,I1402597);
nand I_82296 (I1402345,I1402481,I1402597);
DFFARX1 I_82297 (I1402515,I3563,I1402368,I1402360,);
not I_82298 (I1402659,I936851);
nor I_82299 (I1402676,I1402659,I936848);
nor I_82300 (I1402693,I1402676,I1402498);
DFFARX1 I_82301 (I1402693,I3563,I1402368,I1402357,);
not I_82302 (I1402724,I1402676);
DFFARX1 I_82303 (I1402724,I3563,I1402368,I1402750,);
not I_82304 (I1402758,I1402750);
nor I_82305 (I1402354,I1402758,I1402676);
nor I_82306 (I1402789,I1402659,I936839);
and I_82307 (I1402806,I1402789,I936866);
or I_82308 (I1402823,I1402806,I936857);
DFFARX1 I_82309 (I1402823,I3563,I1402368,I1402849,);
not I_82310 (I1402857,I1402849);
nand I_82311 (I1402874,I1402857,I1402597);
not I_82312 (I1402348,I1402874);
nand I_82313 (I1402342,I1402874,I1402614);
nand I_82314 (I1402339,I1402857,I1402481);
not I_82315 (I1402963,I3570);
DFFARX1 I_82316 (I258318,I3563,I1402963,I1402989,);
DFFARX1 I_82317 (I258321,I3563,I1402963,I1403006,);
not I_82318 (I1403014,I1403006);
nor I_82319 (I1402931,I1402989,I1403014);
DFFARX1 I_82320 (I1403014,I3563,I1402963,I1402946,);
nor I_82321 (I1403059,I258327,I258321);
and I_82322 (I1403076,I1403059,I258324);
nor I_82323 (I1403093,I1403076,I258327);
not I_82324 (I1403110,I258327);
and I_82325 (I1403127,I1403110,I258318);
nand I_82326 (I1403144,I1403127,I258336);
nor I_82327 (I1403161,I1403110,I1403144);
DFFARX1 I_82328 (I1403161,I3563,I1402963,I1402928,);
not I_82329 (I1403192,I1403144);
nand I_82330 (I1403209,I1403014,I1403192);
nand I_82331 (I1402940,I1403076,I1403192);
DFFARX1 I_82332 (I1403110,I3563,I1402963,I1402955,);
not I_82333 (I1403254,I258330);
nor I_82334 (I1403271,I1403254,I258318);
nor I_82335 (I1403288,I1403271,I1403093);
DFFARX1 I_82336 (I1403288,I3563,I1402963,I1402952,);
not I_82337 (I1403319,I1403271);
DFFARX1 I_82338 (I1403319,I3563,I1402963,I1403345,);
not I_82339 (I1403353,I1403345);
nor I_82340 (I1402949,I1403353,I1403271);
nor I_82341 (I1403384,I1403254,I258333);
and I_82342 (I1403401,I1403384,I258339);
or I_82343 (I1403418,I1403401,I258342);
DFFARX1 I_82344 (I1403418,I3563,I1402963,I1403444,);
not I_82345 (I1403452,I1403444);
nand I_82346 (I1403469,I1403452,I1403192);
not I_82347 (I1402943,I1403469);
nand I_82348 (I1402937,I1403469,I1403209);
nand I_82349 (I1402934,I1403452,I1403076);
not I_82350 (I1403558,I3570);
DFFARX1 I_82351 (I1063501,I3563,I1403558,I1403584,);
DFFARX1 I_82352 (I1063492,I3563,I1403558,I1403601,);
not I_82353 (I1403609,I1403601);
nor I_82354 (I1403526,I1403584,I1403609);
DFFARX1 I_82355 (I1403609,I3563,I1403558,I1403541,);
nor I_82356 (I1403654,I1063498,I1063507);
and I_82357 (I1403671,I1403654,I1063510);
nor I_82358 (I1403688,I1403671,I1063498);
not I_82359 (I1403705,I1063498);
and I_82360 (I1403722,I1403705,I1063489);
nand I_82361 (I1403739,I1403722,I1063495);
nor I_82362 (I1403756,I1403705,I1403739);
DFFARX1 I_82363 (I1403756,I3563,I1403558,I1403523,);
not I_82364 (I1403787,I1403739);
nand I_82365 (I1403804,I1403609,I1403787);
nand I_82366 (I1403535,I1403671,I1403787);
DFFARX1 I_82367 (I1403705,I3563,I1403558,I1403550,);
not I_82368 (I1403849,I1063504);
nor I_82369 (I1403866,I1403849,I1063489);
nor I_82370 (I1403883,I1403866,I1403688);
DFFARX1 I_82371 (I1403883,I3563,I1403558,I1403547,);
not I_82372 (I1403914,I1403866);
DFFARX1 I_82373 (I1403914,I3563,I1403558,I1403940,);
not I_82374 (I1403948,I1403940);
nor I_82375 (I1403544,I1403948,I1403866);
nor I_82376 (I1403979,I1403849,I1063489);
and I_82377 (I1403996,I1403979,I1063492);
or I_82378 (I1404013,I1403996,I1063495);
DFFARX1 I_82379 (I1404013,I3563,I1403558,I1404039,);
not I_82380 (I1404047,I1404039);
nand I_82381 (I1404064,I1404047,I1403787);
not I_82382 (I1403538,I1404064);
nand I_82383 (I1403532,I1404064,I1403804);
nand I_82384 (I1403529,I1404047,I1403671);
not I_82385 (I1404153,I3570);
DFFARX1 I_82386 (I291183,I3563,I1404153,I1404179,);
DFFARX1 I_82387 (I291177,I3563,I1404153,I1404196,);
not I_82388 (I1404204,I1404196);
nor I_82389 (I1404121,I1404179,I1404204);
DFFARX1 I_82390 (I1404204,I3563,I1404153,I1404136,);
nor I_82391 (I1404249,I291165,I291186);
and I_82392 (I1404266,I1404249,I291180);
nor I_82393 (I1404283,I1404266,I291165);
not I_82394 (I1404300,I291165);
and I_82395 (I1404317,I1404300,I291162);
nand I_82396 (I1404334,I1404317,I291174);
nor I_82397 (I1404351,I1404300,I1404334);
DFFARX1 I_82398 (I1404351,I3563,I1404153,I1404118,);
not I_82399 (I1404382,I1404334);
nand I_82400 (I1404399,I1404204,I1404382);
nand I_82401 (I1404130,I1404266,I1404382);
DFFARX1 I_82402 (I1404300,I3563,I1404153,I1404145,);
not I_82403 (I1404444,I291189);
nor I_82404 (I1404461,I1404444,I291162);
nor I_82405 (I1404478,I1404461,I1404283);
DFFARX1 I_82406 (I1404478,I3563,I1404153,I1404142,);
not I_82407 (I1404509,I1404461);
DFFARX1 I_82408 (I1404509,I3563,I1404153,I1404535,);
not I_82409 (I1404543,I1404535);
nor I_82410 (I1404139,I1404543,I1404461);
nor I_82411 (I1404574,I1404444,I291171);
and I_82412 (I1404591,I1404574,I291168);
or I_82413 (I1404608,I1404591,I291162);
DFFARX1 I_82414 (I1404608,I3563,I1404153,I1404634,);
not I_82415 (I1404642,I1404634);
nand I_82416 (I1404659,I1404642,I1404382);
not I_82417 (I1404133,I1404659);
nand I_82418 (I1404127,I1404659,I1404399);
nand I_82419 (I1404124,I1404642,I1404266);
not I_82420 (I1404748,I3570);
DFFARX1 I_82421 (I439810,I3563,I1404748,I1404774,);
DFFARX1 I_82422 (I439816,I3563,I1404748,I1404791,);
not I_82423 (I1404799,I1404791);
nor I_82424 (I1404716,I1404774,I1404799);
DFFARX1 I_82425 (I1404799,I3563,I1404748,I1404731,);
nor I_82426 (I1404844,I439825,I439810);
and I_82427 (I1404861,I1404844,I439837);
nor I_82428 (I1404878,I1404861,I439825);
not I_82429 (I1404895,I439825);
and I_82430 (I1404912,I1404895,I439813);
nand I_82431 (I1404929,I1404912,I439834);
nor I_82432 (I1404946,I1404895,I1404929);
DFFARX1 I_82433 (I1404946,I3563,I1404748,I1404713,);
not I_82434 (I1404977,I1404929);
nand I_82435 (I1404994,I1404799,I1404977);
nand I_82436 (I1404725,I1404861,I1404977);
DFFARX1 I_82437 (I1404895,I3563,I1404748,I1404740,);
not I_82438 (I1405039,I439822);
nor I_82439 (I1405056,I1405039,I439813);
nor I_82440 (I1405073,I1405056,I1404878);
DFFARX1 I_82441 (I1405073,I3563,I1404748,I1404737,);
not I_82442 (I1405104,I1405056);
DFFARX1 I_82443 (I1405104,I3563,I1404748,I1405130,);
not I_82444 (I1405138,I1405130);
nor I_82445 (I1404734,I1405138,I1405056);
nor I_82446 (I1405169,I1405039,I439819);
and I_82447 (I1405186,I1405169,I439831);
or I_82448 (I1405203,I1405186,I439828);
DFFARX1 I_82449 (I1405203,I3563,I1404748,I1405229,);
not I_82450 (I1405237,I1405229);
nand I_82451 (I1405254,I1405237,I1404977);
not I_82452 (I1404728,I1405254);
nand I_82453 (I1404722,I1405254,I1404994);
nand I_82454 (I1404719,I1405237,I1404861);
not I_82455 (I1405343,I3570);
DFFARX1 I_82456 (I269028,I3563,I1405343,I1405369,);
DFFARX1 I_82457 (I269031,I3563,I1405343,I1405386,);
not I_82458 (I1405394,I1405386);
nor I_82459 (I1405311,I1405369,I1405394);
DFFARX1 I_82460 (I1405394,I3563,I1405343,I1405326,);
nor I_82461 (I1405439,I269037,I269031);
and I_82462 (I1405456,I1405439,I269034);
nor I_82463 (I1405473,I1405456,I269037);
not I_82464 (I1405490,I269037);
and I_82465 (I1405507,I1405490,I269028);
nand I_82466 (I1405524,I1405507,I269046);
nor I_82467 (I1405541,I1405490,I1405524);
DFFARX1 I_82468 (I1405541,I3563,I1405343,I1405308,);
not I_82469 (I1405572,I1405524);
nand I_82470 (I1405589,I1405394,I1405572);
nand I_82471 (I1405320,I1405456,I1405572);
DFFARX1 I_82472 (I1405490,I3563,I1405343,I1405335,);
not I_82473 (I1405634,I269040);
nor I_82474 (I1405651,I1405634,I269028);
nor I_82475 (I1405668,I1405651,I1405473);
DFFARX1 I_82476 (I1405668,I3563,I1405343,I1405332,);
not I_82477 (I1405699,I1405651);
DFFARX1 I_82478 (I1405699,I3563,I1405343,I1405725,);
not I_82479 (I1405733,I1405725);
nor I_82480 (I1405329,I1405733,I1405651);
nor I_82481 (I1405764,I1405634,I269043);
and I_82482 (I1405781,I1405764,I269049);
or I_82483 (I1405798,I1405781,I269052);
DFFARX1 I_82484 (I1405798,I3563,I1405343,I1405824,);
not I_82485 (I1405832,I1405824);
nand I_82486 (I1405849,I1405832,I1405572);
not I_82487 (I1405323,I1405849);
nand I_82488 (I1405317,I1405849,I1405589);
nand I_82489 (I1405314,I1405832,I1405456);
not I_82490 (I1405938,I3570);
DFFARX1 I_82491 (I231543,I3563,I1405938,I1405964,);
DFFARX1 I_82492 (I231546,I3563,I1405938,I1405981,);
not I_82493 (I1405989,I1405981);
nor I_82494 (I1405906,I1405964,I1405989);
DFFARX1 I_82495 (I1405989,I3563,I1405938,I1405921,);
nor I_82496 (I1406034,I231552,I231546);
and I_82497 (I1406051,I1406034,I231549);
nor I_82498 (I1406068,I1406051,I231552);
not I_82499 (I1406085,I231552);
and I_82500 (I1406102,I1406085,I231543);
nand I_82501 (I1406119,I1406102,I231561);
nor I_82502 (I1406136,I1406085,I1406119);
DFFARX1 I_82503 (I1406136,I3563,I1405938,I1405903,);
not I_82504 (I1406167,I1406119);
nand I_82505 (I1406184,I1405989,I1406167);
nand I_82506 (I1405915,I1406051,I1406167);
DFFARX1 I_82507 (I1406085,I3563,I1405938,I1405930,);
not I_82508 (I1406229,I231555);
nor I_82509 (I1406246,I1406229,I231543);
nor I_82510 (I1406263,I1406246,I1406068);
DFFARX1 I_82511 (I1406263,I3563,I1405938,I1405927,);
not I_82512 (I1406294,I1406246);
DFFARX1 I_82513 (I1406294,I3563,I1405938,I1406320,);
not I_82514 (I1406328,I1406320);
nor I_82515 (I1405924,I1406328,I1406246);
nor I_82516 (I1406359,I1406229,I231558);
and I_82517 (I1406376,I1406359,I231564);
or I_82518 (I1406393,I1406376,I231567);
DFFARX1 I_82519 (I1406393,I3563,I1405938,I1406419,);
not I_82520 (I1406427,I1406419);
nand I_82521 (I1406444,I1406427,I1406167);
not I_82522 (I1405918,I1406444);
nand I_82523 (I1405912,I1406444,I1406184);
nand I_82524 (I1405909,I1406427,I1406051);
not I_82525 (I1406533,I3570);
DFFARX1 I_82526 (I680976,I3563,I1406533,I1406559,);
DFFARX1 I_82527 (I680958,I3563,I1406533,I1406576,);
not I_82528 (I1406584,I1406576);
nor I_82529 (I1406501,I1406559,I1406584);
DFFARX1 I_82530 (I1406584,I3563,I1406533,I1406516,);
nor I_82531 (I1406629,I680964,I680967);
and I_82532 (I1406646,I1406629,I680955);
nor I_82533 (I1406663,I1406646,I680964);
not I_82534 (I1406680,I680964);
and I_82535 (I1406697,I1406680,I680973);
nand I_82536 (I1406714,I1406697,I680961);
nor I_82537 (I1406731,I1406680,I1406714);
DFFARX1 I_82538 (I1406731,I3563,I1406533,I1406498,);
not I_82539 (I1406762,I1406714);
nand I_82540 (I1406779,I1406584,I1406762);
nand I_82541 (I1406510,I1406646,I1406762);
DFFARX1 I_82542 (I1406680,I3563,I1406533,I1406525,);
not I_82543 (I1406824,I680958);
nor I_82544 (I1406841,I1406824,I680973);
nor I_82545 (I1406858,I1406841,I1406663);
DFFARX1 I_82546 (I1406858,I3563,I1406533,I1406522,);
not I_82547 (I1406889,I1406841);
DFFARX1 I_82548 (I1406889,I3563,I1406533,I1406915,);
not I_82549 (I1406923,I1406915);
nor I_82550 (I1406519,I1406923,I1406841);
nor I_82551 (I1406954,I1406824,I680970);
and I_82552 (I1406971,I1406954,I680979);
or I_82553 (I1406988,I1406971,I680955);
DFFARX1 I_82554 (I1406988,I3563,I1406533,I1407014,);
not I_82555 (I1407022,I1407014);
nand I_82556 (I1407039,I1407022,I1406762);
not I_82557 (I1406513,I1407039);
nand I_82558 (I1406507,I1407039,I1406779);
nand I_82559 (I1406504,I1407022,I1406646);
not I_82560 (I1407128,I3570);
DFFARX1 I_82561 (I176803,I3563,I1407128,I1407154,);
DFFARX1 I_82562 (I176806,I3563,I1407128,I1407171,);
not I_82563 (I1407179,I1407171);
nor I_82564 (I1407096,I1407154,I1407179);
DFFARX1 I_82565 (I1407179,I3563,I1407128,I1407111,);
nor I_82566 (I1407224,I176812,I176806);
and I_82567 (I1407241,I1407224,I176809);
nor I_82568 (I1407258,I1407241,I176812);
not I_82569 (I1407275,I176812);
and I_82570 (I1407292,I1407275,I176803);
nand I_82571 (I1407309,I1407292,I176821);
nor I_82572 (I1407326,I1407275,I1407309);
DFFARX1 I_82573 (I1407326,I3563,I1407128,I1407093,);
not I_82574 (I1407357,I1407309);
nand I_82575 (I1407374,I1407179,I1407357);
nand I_82576 (I1407105,I1407241,I1407357);
DFFARX1 I_82577 (I1407275,I3563,I1407128,I1407120,);
not I_82578 (I1407419,I176815);
nor I_82579 (I1407436,I1407419,I176803);
nor I_82580 (I1407453,I1407436,I1407258);
DFFARX1 I_82581 (I1407453,I3563,I1407128,I1407117,);
not I_82582 (I1407484,I1407436);
DFFARX1 I_82583 (I1407484,I3563,I1407128,I1407510,);
not I_82584 (I1407518,I1407510);
nor I_82585 (I1407114,I1407518,I1407436);
nor I_82586 (I1407549,I1407419,I176818);
and I_82587 (I1407566,I1407549,I176824);
or I_82588 (I1407583,I1407566,I176827);
DFFARX1 I_82589 (I1407583,I3563,I1407128,I1407609,);
not I_82590 (I1407617,I1407609);
nand I_82591 (I1407634,I1407617,I1407357);
not I_82592 (I1407108,I1407634);
nand I_82593 (I1407102,I1407634,I1407374);
nand I_82594 (I1407099,I1407617,I1407241);
not I_82595 (I1407723,I3570);
DFFARX1 I_82596 (I1018887,I3563,I1407723,I1407749,);
DFFARX1 I_82597 (I1018905,I3563,I1407723,I1407766,);
not I_82598 (I1407774,I1407766);
nor I_82599 (I1407691,I1407749,I1407774);
DFFARX1 I_82600 (I1407774,I3563,I1407723,I1407706,);
nor I_82601 (I1407819,I1018884,I1018896);
and I_82602 (I1407836,I1407819,I1018881);
nor I_82603 (I1407853,I1407836,I1018884);
not I_82604 (I1407870,I1018884);
and I_82605 (I1407887,I1407870,I1018890);
nand I_82606 (I1407904,I1407887,I1018902);
nor I_82607 (I1407921,I1407870,I1407904);
DFFARX1 I_82608 (I1407921,I3563,I1407723,I1407688,);
not I_82609 (I1407952,I1407904);
nand I_82610 (I1407969,I1407774,I1407952);
nand I_82611 (I1407700,I1407836,I1407952);
DFFARX1 I_82612 (I1407870,I3563,I1407723,I1407715,);
not I_82613 (I1408014,I1018893);
nor I_82614 (I1408031,I1408014,I1018890);
nor I_82615 (I1408048,I1408031,I1407853);
DFFARX1 I_82616 (I1408048,I3563,I1407723,I1407712,);
not I_82617 (I1408079,I1408031);
DFFARX1 I_82618 (I1408079,I3563,I1407723,I1408105,);
not I_82619 (I1408113,I1408105);
nor I_82620 (I1407709,I1408113,I1408031);
nor I_82621 (I1408144,I1408014,I1018881);
and I_82622 (I1408161,I1408144,I1018908);
or I_82623 (I1408178,I1408161,I1018899);
DFFARX1 I_82624 (I1408178,I3563,I1407723,I1408204,);
not I_82625 (I1408212,I1408204);
nand I_82626 (I1408229,I1408212,I1407952);
not I_82627 (I1407703,I1408229);
nand I_82628 (I1407697,I1408229,I1407969);
nand I_82629 (I1407694,I1408212,I1407836);
endmodule


