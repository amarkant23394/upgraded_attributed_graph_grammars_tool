module test_I3362(I1637,I1383,I1477,I1470,I3362);
input I1637,I1383,I1477,I1470;
output I3362;
wire I1518,I3388,I3422,I1480,I1976,I1880,I1483,I1959;
not I_0(I1518,I1477);
not I_1(I3388,I1477);
or I_2(I3422,I1483,I1480);
DFFARX1 I_3(I3422,I1470,I3388,,,I3362,);
DFFARX1 I_4(I1976,I1470,I1518,,,I1480,);
and I_5(I1976,I1637,I1959);
DFFARX1 I_6(I1383,I1470,I1518,,,I1880,);
DFFARX1 I_7(I1880,I1470,I1518,,,I1483,);
nand I_8(I1959,I1880);
endmodule


