module test_I14945(I1477,I1470,I14945);
input I1477,I1470;
output I14945;
wire I12602,I12670,I12584,I12913,I15109,I12930,I12783,I15126,I14965,I15372,I10609;
not I_0(I12602,I12930);
DFFARX1 I_1(I1470,,,I12670,);
and I_2(I12584,I12670,I12783);
DFFARX1 I_3(I1470,,,I12913,);
not I_4(I15109,I12584);
and I_5(I12930,I12913,I10609);
DFFARX1 I_6(I1470,,,I12783,);
nand I_7(I14945,I15372,I15126);
not I_8(I15126,I15109);
not I_9(I14965,I1477);
DFFARX1 I_10(I12602,I1470,I14965,,,I15372,);
DFFARX1 I_11(I1470,,,I10609,);
endmodule


