module test_final(IN_1_0_l_6,IN_2_0_l_6,IN_3_0_l_6,IN_4_0_l_6,IN_1_1_l_6,IN_2_1_l_6,IN_3_1_l_6,IN_1_10_l_6,IN_2_10_l_6,IN_3_10_l_6,IN_4_10_l_6,blif_clk_net_5_r_2,blif_reset_net_5_r_2,N1371_0_r_2,N6147_3_r_2,G78_5_r_2,n_576_5_r_2,n_547_5_r_2,N1372_10_r_2,N1508_10_r_2);
input IN_1_0_l_6,IN_2_0_l_6,IN_3_0_l_6,IN_4_0_l_6,IN_1_1_l_6,IN_2_1_l_6,IN_3_1_l_6,IN_1_10_l_6,IN_2_10_l_6,IN_3_10_l_6,IN_4_10_l_6,blif_clk_net_5_r_2,blif_reset_net_5_r_2;
output N1371_0_r_2,N6147_3_r_2,G78_5_r_2,n_576_5_r_2,n_547_5_r_2,N1372_10_r_2,N1508_10_r_2;
wire N1371_0_r_6,N1508_0_r_6,N6147_3_r_6,n_429_or_0_5_r_6,G78_5_r_6,n_576_5_r_6,n_102_5_r_6,n_547_5_r_6,N1372_10_r_6,N1508_10_r_6,n_431_5_r_6,n24_6,n25_6,n26_6,n27_6,n28_6,n29_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,N1508_0_r_2,n_429_or_0_5_r_2,n_102_5_r_2,n_431_5_r_2,n6_2,n21_2,n22_2,n23_2,n24_2,n25_2,n26_2,n27_2,n28_2,n29_2,n30_2,n31_2,n32_2;
nor I_0(N1371_0_r_6,n26_6,n38_6);
not I_1(N1508_0_r_6,n38_6);
nor I_2(N6147_3_r_6,n30_6,n35_6);
nand I_3(n_429_or_0_5_r_6,n30_6,n32_6);
DFFARX1 I_4(n_431_5_r_6,blif_clk_net_5_r_2,n6_2,G78_5_r_6,);
nand I_5(n_576_5_r_6,n24_6,n25_6);
not I_6(n_102_5_r_6,n26_6);
or I_7(n_547_5_r_6,n_429_or_0_5_r_6,n26_6);
not I_8(N1372_10_r_6,n37_6);
nor I_9(N1508_10_r_6,n36_6,n37_6);
nand I_10(n_431_5_r_6,n_102_5_r_6,n28_6);
nor I_11(n24_6,n33_6,n34_6);
nor I_12(n25_6,n26_6,n27_6);
nor I_13(n26_6,IN_2_0_l_6,n40_6);
nand I_14(n27_6,IN_1_1_l_6,IN_2_1_l_6);
nand I_15(n28_6,n29_6,n30_6);
nor I_16(n29_6,IN_3_1_l_6,n31_6);
not I_17(n30_6,n27_6);
nor I_18(n31_6,n39_6,n40_6);
nor I_19(n32_6,IN_3_1_l_6,n24_6);
not I_20(n33_6,IN_1_10_l_6);
not I_21(n34_6,IN_2_10_l_6);
or I_22(n35_6,n26_6,n31_6);
and I_23(n36_6,IN_3_1_l_6,n38_6);
nand I_24(n37_6,n30_6,n31_6);
nand I_25(n38_6,IN_2_10_l_6,n41_6);
nor I_26(n39_6,IN_3_0_l_6,IN_4_0_l_6);
not I_27(n40_6,IN_1_0_l_6);
nor I_28(n41_6,n33_6,n42_6);
nor I_29(n42_6,IN_3_10_l_6,IN_4_10_l_6);
nor I_30(N1371_0_r_2,n23_2,n24_2);
not I_31(N1508_0_r_2,n24_2);
nor I_32(N6147_3_r_2,n22_2,n26_2);
nand I_33(n_429_or_0_5_r_2,n22_2,N1508_10_r_6);
DFFARX1 I_34(n_431_5_r_2,blif_clk_net_5_r_2,n6_2,G78_5_r_2,);
nand I_35(n_576_5_r_2,n21_2,n22_2);
not I_36(n_102_5_r_2,n23_2);
nand I_37(n_547_5_r_2,n22_2,n24_2);
not I_38(N1372_10_r_2,n29_2);
nor I_39(N1508_10_r_2,n28_2,n29_2);
nand I_40(n_431_5_r_2,n_102_5_r_2,n25_2);
not I_41(n6_2,blif_reset_net_5_r_2);
nor I_42(n21_2,n23_2,N1508_10_r_6);
and I_43(n22_2,G78_5_r_6,n_576_5_r_6);
nor I_44(n23_2,n24_2,n31_2);
nand I_45(n24_2,N1371_0_r_6,n_547_5_r_6);
nand I_46(n25_2,n26_2,n27_2);
nor I_47(n26_2,n30_2,N1371_0_r_6);
not I_48(n27_2,n_429_or_0_5_r_2);
nor I_49(n28_2,n22_2,n23_2);
nand I_50(n29_2,N1508_0_r_2,n26_2);
or I_51(n30_2,N1508_0_r_6,N6147_3_r_6);
nor I_52(n31_2,n32_2,N6147_3_r_6);
and I_53(n32_2,N1372_10_r_6,N1508_0_r_6);
endmodule


