module test_I10185(I6321,I1477,I6309,I7799,I7652,I1470,I6318,I10185);
input I6321,I1477,I6309,I7799,I7652,I1470,I6318;
output I10185;
wire I8107,I7562,I8090,I7547,I7570,I7816,I8059,I7833,I7977,I7669;
not I_0(I8107,I8090);
nand I_1(I7562,I8107,I7833);
DFFARX1 I_2(I6309,I1470,I7570,,,I8090,);
not I_3(I7547,I8059);
not I_4(I7570,I1477);
DFFARX1 I_5(I7799,I1470,I7570,,,I7816,);
DFFARX1 I_6(I7977,I1470,I7570,,,I8059,);
nor I_7(I7833,I7816,I7669);
nand I_8(I10185,I7547,I7562);
DFFARX1 I_9(I6321,I1470,I7570,,,I7977,);
nand I_10(I7669,I7652,I6318);
endmodule


