module test_I3815(I1477,I1849,I1637,I1928,I2038,I1470,I1959,I3815);
input I1477,I1849,I1637,I1928,I2038,I1470,I1959;
output I3815;
wire I3422,I3781,I1507,I1495,I3764,I3685,I3747,I1483,I3388,I3668,I3405,I1518,I1480,I1498,I3798,I1976,I2103;
or I_0(I3422,I1483,I1480);
nor I_1(I3781,I3422,I3764);
nor I_2(I1507,I1637);
DFFARX1 I_3(I2103,I1470,I1518,,,I1495,);
not I_4(I3764,I3747);
or I_5(I3815,I3405,I3798);
and I_6(I3685,I3668,I1498);
DFFARX1 I_7(I1470,I3388,,,I3747,);
DFFARX1 I_8(I1470,I1518,,,I1483,);
not I_9(I3388,I1477);
DFFARX1 I_10(I1507,I1470,I3388,,,I3668,);
or I_11(I3405,I1480,I1495);
not I_12(I1518,I1477);
DFFARX1 I_13(I1976,I1470,I1518,,,I1480,);
nand I_14(I1498,I2038,I1928);
and I_15(I3798,I3685,I3781);
and I_16(I1976,I1637,I1959);
or I_17(I2103,I2038,I1849);
endmodule


