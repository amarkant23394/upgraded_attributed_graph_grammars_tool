module test_final(G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_17,blif_reset_net_1_r_17,G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17);
input G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_17,blif_reset_net_1_r_17;
output G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17;
wire G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16,n4_1_l_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16,n_431_0_l_17,n6_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17;
DFFARX1 I_0(n4_1_r_16,blif_clk_net_1_r_17,n6_17,G42_1_r_16,);
nor I_1(n_572_1_r_16,n20_16,n21_16);
nand I_2(n_573_1_r_16,n18_16,n19_16);
nor I_3(n_549_1_r_16,n23_16,n24_16);
nand I_4(n_569_1_r_16,n18_16,n22_16);
nor I_5(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_6(N1_4_r_16,blif_clk_net_1_r_17,n6_17,G199_4_r_16,);
DFFARX1 I_7(n6_16,blif_clk_net_1_r_17,n6_17,G214_4_r_16,);
DFFARX1 I_8(n_573_1_l_16,blif_clk_net_1_r_17,n6_17,ACVQN1_5_r_16,);
not I_9(P6_5_r_16,P6_5_r_internal_16);
nor I_10(n4_1_l_16,G18_1_l_16,IN_1_1_l_16);
DFFARX1 I_11(n4_1_l_16,blif_clk_net_1_r_17,n6_17,n29_16,);
DFFARX1 I_12(IN_1_3_l_16,blif_clk_net_1_r_17,n6_17,n16_internal_16,);
not I_13(n16_16,n16_internal_16);
DFFARX1 I_14(IN_2_3_l_16,blif_clk_net_1_r_17,n6_17,ACVQN1_3_l_16,);
nor I_15(n4_1_r_16,n29_16,n21_16);
nor I_16(N1_4_r_16,n27_16,n28_16);
not I_17(n6_16,n19_16);
or I_18(n_573_1_l_16,IN_5_1_l_16,IN_9_1_l_16);
nor I_19(n_452_1_l_16,G18_1_l_16,IN_5_1_l_16);
DFFARX1 I_20(n_452_1_l_16,blif_clk_net_1_r_17,n6_17,P6_5_r_internal_16,);
not I_21(n18_16,n20_16);
nor I_22(n19_16,IN_9_1_l_16,IN_10_1_l_16);
nor I_23(n20_16,G15_1_l_16,IN_7_1_l_16);
nor I_24(n21_16,IN_10_1_l_16,n25_16);
nand I_25(n22_16,IN_4_3_l_16,ACVQN1_3_l_16);
not I_26(n23_16,n22_16);
nor I_27(n24_16,n16_16,n20_16);
nor I_28(n25_16,G15_1_l_16,n26_16);
not I_29(n26_16,IN_4_1_l_16);
and I_30(n27_16,IN_9_1_l_16,n29_16);
not I_31(n28_16,n_452_1_l_16);
DFFARX1 I_32(n4_1_r_17,blif_clk_net_1_r_17,n6_17,G42_1_r_17,);
nor I_33(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_34(n_573_1_r_17,n20_17,n21_17);
nand I_35(n_549_1_r_17,n23_17,n24_17);
nand I_36(n_569_1_r_17,n21_17,n22_17);
not I_37(n_452_1_r_17,n23_17);
DFFARX1 I_38(n19_17,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_17,);
nor I_39(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_40(N1_4_r_17,blif_clk_net_1_r_17,n6_17,G199_4_r_17,);
DFFARX1 I_41(n5_17,blif_clk_net_1_r_17,n6_17,G214_4_r_17,);
or I_42(n_431_0_l_17,n26_17,n_572_1_r_16);
not I_43(n6_17,blif_reset_net_1_r_17);
DFFARX1 I_44(n_431_0_l_17,blif_clk_net_1_r_17,n6_17,n20_internal_17,);
not I_45(n20_17,n20_internal_17);
DFFARX1 I_46(P6_5_r_16,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_17,);
DFFARX1 I_47(n_569_1_r_16,blif_clk_net_1_r_17,n6_17,n19_internal_17,);
not I_48(n19_17,n19_internal_17);
nor I_49(n4_1_r_17,n5_17,n25_17);
not I_50(n2_17,n29_17);
DFFARX1 I_51(n2_17,blif_clk_net_1_r_17,n6_17,n17_internal_17,);
not I_52(n17_17,n17_internal_17);
nor I_53(N1_4_r_17,n29_17,n31_17);
not I_54(n5_17,n_549_1_r_16);
and I_55(n21_17,n32_17,ACVQN1_5_r_16);
not I_56(n22_17,n25_17);
nand I_57(n23_17,n20_17,n22_17);
nand I_58(n24_17,n19_17,n22_17);
nand I_59(n25_17,n30_17,G42_1_r_16);
and I_60(n26_17,n27_17,G214_4_r_16);
nor I_61(n27_17,n28_17,n_452_1_r_16);
not I_62(n28_17,G42_1_r_16);
nor I_63(n29_17,n28_17,n_573_1_r_16);
and I_64(n30_17,n5_17,n_573_1_r_16);
nor I_65(n31_17,n21_17,n_549_1_r_16);
nor I_66(n32_17,n_549_1_r_16,G199_4_r_16);
endmodule


