module test_final(IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_3_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_4_4_l_2,IN_5_4_l_2,blif_clk_net_5_r_4,blif_reset_net_5_r_4,N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4);
input IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_3_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_4_4_l_2,IN_5_4_l_2,blif_clk_net_5_r_4,blif_reset_net_5_r_4;
output N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4;
wire N1371_0_r_2,N1508_0_r_2,N6147_3_r_2,n_429_or_0_5_r_2,G78_5_r_2,n_576_5_r_2,n_102_5_r_2,n_547_5_r_2,N1372_10_r_2,N1508_10_r_2,n_431_5_r_2,n21_2,n22_2,n23_2,n24_2,n25_2,n26_2,n27_2,n28_2,n29_2,n30_2,n31_2,n32_2,N1371_0_r_4,n_102_5_r_4,n_431_5_r_4,n4_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4;
nor I_0(N1371_0_r_2,n23_2,n24_2);
not I_1(N1508_0_r_2,n24_2);
nor I_2(N6147_3_r_2,n22_2,n26_2);
nand I_3(n_429_or_0_5_r_2,IN_3_1_l_2,n22_2);
DFFARX1 I_4(n_431_5_r_2,blif_clk_net_5_r_4,n4_4,G78_5_r_2,);
nand I_5(n_576_5_r_2,n21_2,n22_2);
not I_6(n_102_5_r_2,n23_2);
nand I_7(n_547_5_r_2,n22_2,n24_2);
not I_8(N1372_10_r_2,n29_2);
nor I_9(N1508_10_r_2,n28_2,n29_2);
nand I_10(n_431_5_r_2,n_102_5_r_2,n25_2);
nor I_11(n21_2,IN_3_1_l_2,n23_2);
and I_12(n22_2,IN_1_1_l_2,IN_2_1_l_2);
nor I_13(n23_2,n24_2,n31_2);
nand I_14(n24_2,IN_1_4_l_2,IN_2_4_l_2);
nand I_15(n25_2,n26_2,n27_2);
nor I_16(n26_2,IN_1_3_l_2,n30_2);
not I_17(n27_2,n_429_or_0_5_r_2);
nor I_18(n28_2,n22_2,n23_2);
nand I_19(n29_2,N1508_0_r_2,n26_2);
or I_20(n30_2,IN_2_3_l_2,IN_3_3_l_2);
nor I_21(n31_2,IN_5_4_l_2,n32_2);
and I_22(n32_2,IN_3_4_l_2,IN_4_4_l_2);
nor I_23(N1371_0_r_4,n25_4,n29_4);
nor I_24(N1508_0_r_4,n25_4,n32_4);
nor I_25(N6147_2_r_4,n24_4,n31_4);
or I_26(n_429_or_0_5_r_4,n23_4,n30_4);
DFFARX1 I_27(n_431_5_r_4,blif_clk_net_5_r_4,n4_4,G78_5_r_4,);
nand I_28(n_576_5_r_4,n22_4,n23_4);
nand I_29(n_102_5_r_4,n34_4,n35_4);
nand I_30(n_547_5_r_4,n26_4,n27_4);
nor I_31(N1507_6_r_4,n27_4,n30_4);
nor I_32(N1508_6_r_4,n30_4,n33_4);
nand I_33(n_431_5_r_4,n_102_5_r_4,n28_4);
not I_34(n4_4,blif_reset_net_5_r_4);
nor I_35(n22_4,n24_4,n25_4);
nor I_36(n23_4,n37_4,N1371_0_r_2);
not I_37(n24_4,n_102_5_r_4);
nand I_38(n25_4,n_547_5_r_2,G78_5_r_2);
nor I_39(n26_4,n23_4,n24_4);
not I_40(n27_4,n25_4);
nand I_41(n28_4,n23_4,n29_4);
nor I_42(n29_4,n25_4,n_576_5_r_2);
not I_43(n30_4,n29_4);
nor I_44(n31_4,N1371_0_r_4,n32_4);
nor I_45(n32_4,n23_4,n29_4);
nand I_46(n33_4,n23_4,n24_4);
nor I_47(n34_4,N6147_3_r_2,N1508_10_r_2);
or I_48(n35_4,n36_4,N1372_10_r_2);
nor I_49(n36_4,G78_5_r_2,n_576_5_r_2);
or I_50(n37_4,N1371_0_r_2,N6147_3_r_2);
endmodule


