module test_I6045(I4512,I4578,I4917,I4506,I4629,I1470_clk,I1477_rst,I6045);
input I4512,I4578,I4917,I4506,I4629,I1470_clk,I1477_rst;
output I6045;
wire I5932,I5994,I6028,I5915,I4595,I4544_rst,I6011,I4527,I5751_rst,I4521;
not I_0(I5932,I5915);
nand I_1(I5994,I4512,I4506);
DFFARX1 I_2 (I6011,I1470_clk,I5751_rst,I6028);
DFFARX1 I_3 (I4527,I1470_clk,I5751_rst,I5915);
DFFARX1 I_4 (I4578,I1470_clk,I4544_rst,I4595);
not I_5(I4544_rst,I1477_rst);
nor I_6(I6045,I6028,I5932);
and I_7(I6011,I5994,I4521);
or I_8(I4527,I4629,I4595);
not I_9(I5751_rst,I1477_rst);
DFFARX1 I_10 (I4917,I1470_clk,I4544_rst,I4521);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule