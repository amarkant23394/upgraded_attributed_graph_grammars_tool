module test_I17413(I1477,I17413);
input I1477;
output I17413;
wire ;
not I_0(I17413,I1477);
endmodule


