module test_I10120(I6843,I6705,I7587,I7799,I1470_clk,I1477_rst,I10120);
input I6843,I6705,I7587,I7799,I1470_clk,I1477_rst;
output I10120;
wire I6291,I7816,I7535,I7881,I7946,I7570_rst,I7538,I7898,I6329_rst,I6297,I7915,I7714;
DFFARX1 I_0 (I6705,I1470_clk,I6329_rst,I6291);
nor I_1(I10120,I7538,I7535);
DFFARX1 I_2 (I7799,I1470_clk,I7570_rst,I7816);
and I_3(I7535,I7714,I7946);
nand I_4(I7881,I7587,I6291);
DFFARX1 I_5 (I7881,I1470_clk,I7570_rst,I7946);
not I_6(I7570_rst,I1477_rst);
DFFARX1 I_7 (I7915,I1470_clk,I7570_rst,I7538);
nand I_8(I7898,I7881,I7816);
not I_9(I6329_rst,I1477_rst);
DFFARX1 I_10 (I6843,I1470_clk,I6329_rst,I6297);
and I_11(I7915,I7881,I7898);
not I_12(I7714,I6297);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule