module test_final(IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_7_r_2,blif_reset_net_7_r_2,N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2);
input IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_7_r_2,blif_reset_net_7_r_2;
output N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2;
wire N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_549_7_r_5,n_569_7_r_5,n_452_7_r_5,n4_7_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5,n4_7_l_2,n10_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2;
nor I_0(N1371_0_r_5,n28_5,n46_5);
nand I_1(N1508_0_r_5,n26_5,n43_5);
not I_2(N1372_1_r_5,n43_5);
nor I_3(N1508_1_r_5,n30_5,n43_5);
nor I_4(N6147_2_r_5,n29_5,n32_5);
nor I_5(N1507_6_r_5,n26_5,n44_5);
nor I_6(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_7(n4_7_r_5,blif_clk_net_7_r_2,n10_2,G42_7_r_5,);
and I_8(n_572_7_r_5,n27_5,n28_5);
nand I_9(n_573_7_r_5,n26_5,n27_5);
nand I_10(n_549_7_r_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_11(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_12(n_452_7_r_5,n29_5);
nor I_13(n4_7_r_5,n30_5,n31_5);
not I_14(n26_5,n35_5);
nand I_15(n27_5,n40_5,n41_5);
nand I_16(n28_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_17(n29_5,n27_5,n33_5);
nor I_18(n30_5,IN_1_3_l_5,n45_5);
not I_19(n31_5,n_549_7_r_5);
nor I_20(n32_5,n34_5,n35_5);
not I_21(n33_5,n30_5);
nor I_22(n34_5,n31_5,n36_5);
nor I_23(n35_5,IN_3_1_l_5,n28_5);
not I_24(n36_5,n28_5);
nand I_25(n37_5,n36_5,n38_5);
nand I_26(n38_5,n26_5,n39_5);
nand I_27(n39_5,n30_5,n31_5);
nor I_28(n40_5,IN_1_2_l_5,IN_2_2_l_5);
or I_29(n41_5,IN_5_2_l_5,n42_5);
nor I_30(n42_5,IN_3_2_l_5,IN_4_2_l_5);
nand I_31(n43_5,n36_5,n46_5);
nor I_32(n44_5,n_549_7_r_5,n33_5);
or I_33(n45_5,IN_2_3_l_5,IN_3_3_l_5);
and I_34(n46_5,n31_5,n47_5);
or I_35(n47_5,IN_3_10_l_5,IN_4_10_l_5);
nor I_36(N1371_0_r_2,n32_2,n35_2);
nor I_37(N1508_0_r_2,n32_2,n55_2);
not I_38(N1372_1_r_2,n54_2);
nor I_39(N1508_1_r_2,n59_2,n54_2);
nor I_40(N6147_2_r_2,n42_2,n43_2);
nor I_41(N1507_6_r_2,n40_2,n53_2);
nor I_42(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_43(n4_7_r_2,blif_clk_net_7_r_2,n10_2,G42_7_r_2,);
nor I_44(n_572_7_r_2,n36_2,n37_2);
or I_45(n_573_7_r_2,n34_2,n35_2);
nor I_46(n_549_7_r_2,n40_2,n41_2);
nand I_47(n_569_7_r_2,n38_2,n39_2);
nor I_48(n_452_7_r_2,n59_2,n35_2);
nor I_49(n4_7_l_2,N1508_6_r_5,N1372_1_r_5);
not I_50(n10_2,blif_reset_net_7_r_2);
DFFARX1 I_51(n4_7_l_2,blif_clk_net_7_r_2,n10_2,n59_2,);
not I_52(n33_2,n59_2);
and I_53(N3_8_l_2,n49_2,n_573_7_r_5);
DFFARX1 I_54(N3_8_l_2,blif_clk_net_7_r_2,n10_2,n32_internal_2,);
not I_55(n32_2,n32_internal_2);
nor I_56(n4_7_r_2,n59_2,n36_2);
not I_57(n34_2,n39_2);
nor I_58(n35_2,N1508_0_r_5,N6147_2_r_5);
nor I_59(n36_2,G42_7_r_5,N1372_1_r_5);
or I_60(n37_2,N1371_0_r_5,N1507_6_r_5);
not I_61(n38_2,n40_2);
nand I_62(n39_2,n45_2,n57_2);
nor I_63(n40_2,n47_2,N1372_1_r_5);
nor I_64(n41_2,n32_2,n36_2);
not I_65(n42_2,n53_2);
nand I_66(n43_2,n44_2,n45_2);
nand I_67(n44_2,n38_2,n46_2);
not I_68(n45_2,N1371_0_r_5);
nand I_69(n46_2,n47_2,n48_2);
nand I_70(n47_2,n_569_7_r_5,N1371_0_r_5);
or I_71(n48_2,N1508_1_r_5,n_452_7_r_5);
nand I_72(n49_2,N6147_2_r_5,n_572_7_r_5);
nand I_73(n50_2,n51_2,n52_2);
not I_74(n51_2,n47_2);
nand I_75(n52_2,n38_2,n53_2);
nor I_76(n53_2,N1507_6_r_5,G42_7_r_5);
nand I_77(n54_2,n42_2,n56_2);
nor I_78(n55_2,n34_2,n56_2);
nor I_79(n56_2,N1508_1_r_5,n_452_7_r_5);
nand I_80(n57_2,n58_2,N1508_0_r_5);
not I_81(n58_2,n_452_7_r_5);
endmodule


