module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_8,blif_reset_net_1_r_8,G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_8,blif_reset_net_1_r_8;
output G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8;
wire G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6,N3_2_l_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6,n_431_0_l_8,n8_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8;
DFFARX1 I_0(n4_1_r_6,blif_clk_net_1_r_8,n8_8,G42_1_r_6,);
nor I_1(n_572_1_r_6,n27_6,n28_6);
nand I_2(n_573_1_r_6,n18_6,n19_6);
nor I_3(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_4(n_569_1_r_6,n19_6,n20_6);
nor I_5(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_6(N1_4_r_6,blif_clk_net_1_r_8,n8_8,G199_4_r_6,);
DFFARX1 I_7(n_42_2_l_6,blif_clk_net_1_r_8,n8_8,G214_4_r_6,);
DFFARX1 I_8(n_42_2_l_6,blif_clk_net_1_r_8,n8_8,ACVQN1_5_r_6,);
not I_9(P6_5_r_6,P6_5_r_internal_6);
and I_10(N3_2_l_6,IN_6_2_l_6,n23_6);
DFFARX1 I_11(N3_2_l_6,blif_clk_net_1_r_8,n8_8,n27_6,);
not I_12(n17_6,n27_6);
DFFARX1 I_13(IN_1_3_l_6,blif_clk_net_1_r_8,n8_8,n28_6,);
DFFARX1 I_14(IN_2_3_l_6,blif_clk_net_1_r_8,n8_8,n26_6,);
and I_15(N1_4_l_6,IN_6_4_l_6,n25_6);
DFFARX1 I_16(N1_4_l_6,blif_clk_net_1_r_8,n8_8,n29_6,);
not I_17(n18_6,n29_6);
DFFARX1 I_18(IN_3_4_l_6,blif_clk_net_1_r_8,n8_8,G214_4_l_6,);
not I_19(n12_6,G214_4_l_6);
nor I_20(n4_1_r_6,n28_6,n22_6);
nor I_21(N1_4_r_6,n12_6,n24_6);
nor I_22(n_42_2_l_6,IN_1_2_l_6,IN_3_2_l_6);
DFFARX1 I_23(G214_4_l_6,blif_clk_net_1_r_8,n8_8,P6_5_r_internal_6,);
nand I_24(n19_6,IN_4_3_l_6,n26_6);
not I_25(n20_6,n_42_2_l_6);
nor I_26(n21_6,n17_6,n28_6);
and I_27(n22_6,IN_4_3_l_6,n26_6);
nand I_28(n23_6,IN_2_2_l_6,IN_3_2_l_6);
nor I_29(n24_6,n17_6,n18_6);
nand I_30(n25_6,IN_1_4_l_6,IN_2_4_l_6);
DFFARX1 I_31(n4_1_r_8,blif_clk_net_1_r_8,n8_8,G42_1_r_8,);
nor I_32(n_572_1_r_8,n39_8,n23_8);
and I_33(n_549_1_r_8,n38_8,n23_8);
nand I_34(n_569_1_r_8,n38_8,n24_8);
nor I_35(n_452_1_r_8,n25_8,n26_8);
nor I_36(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_37(N3_2_r_8,blif_clk_net_1_r_8,n8_8,G199_2_r_8,);
DFFARX1 I_38(N1_4_r_8,blif_clk_net_1_r_8,n8_8,G199_4_r_8,);
DFFARX1 I_39(G78_0_l_8,blif_clk_net_1_r_8,n8_8,G214_4_r_8,);
or I_40(n_431_0_l_8,n29_8,G199_4_r_6);
not I_41(n8_8,blif_reset_net_1_r_8);
DFFARX1 I_42(n_431_0_l_8,blif_clk_net_1_r_8,n8_8,G78_0_l_8,);
not I_43(n19_8,G78_0_l_8);
DFFARX1 I_44(G214_4_r_6,blif_clk_net_1_r_8,n8_8,n39_8,);
not I_45(n22_8,n39_8);
DFFARX1 I_46(G42_1_r_6,blif_clk_net_1_r_8,n8_8,n38_8,);
nor I_47(n4_1_r_8,G78_0_l_8,n33_8);
nor I_48(N3_2_r_8,n22_8,n35_8);
nor I_49(N1_4_r_8,n27_8,n37_8);
nand I_50(n23_8,n32_8,n_452_1_r_6);
not I_51(n24_8,n23_8);
nand I_52(n25_8,n36_8,G42_1_r_6);
nand I_53(n26_8,n27_8,n28_8);
nor I_54(n27_8,n31_8,ACVQN1_5_r_6);
not I_55(n28_8,n_549_1_r_6);
and I_56(n29_8,n30_8,n_569_1_r_6);
nor I_57(n30_8,n31_8,n_572_1_r_6);
not I_58(n31_8,n_573_1_r_6);
and I_59(n32_8,n28_8,ACVQN1_5_r_6);
nand I_60(n33_8,n28_8,n34_8);
not I_61(n34_8,n25_8);
nor I_62(n35_8,n34_8,n_549_1_r_6);
not I_63(n36_8,P6_5_r_6);
nor I_64(n37_8,n19_8,n38_8);
endmodule


