module test_I13809(I12287,I1477,I1470,I10287,I13809);
input I12287,I1477,I1470,I10287;
output I13809;
wire I11947,I12541,I12442,I12304,I12425,I11953,I12349,I10052,I13792,I10020,I12106,I12524,I11965,I11973;
nand I_0(I11947,I12106,I12524);
nor I_1(I12541,I12349,I12524);
not I_2(I12442,I12425);
and I_3(I12304,I12106,I12287);
DFFARX1 I_4(I1470,I11973,,,I12425,);
nand I_5(I11953,I12442,I12541);
DFFARX1 I_6(I1470,I11973,,,I12349,);
not I_7(I10052,I1477);
nand I_8(I13792,I11953,I11965);
DFFARX1 I_9(I10287,I1470,I10052,,,I10020,);
and I_10(I13809,I13792,I11947);
not I_11(I12106,I10020);
not I_12(I12524,I12442);
DFFARX1 I_13(I12304,I1470,I11973,,,I11965,);
not I_14(I11973,I1477);
endmodule


