module test_I10044(I7550,I7621,I1477,I7850,I1470,I10202,I10044);
input I7550,I7621,I1477,I7850,I1470,I10202;
output I10044;
wire I7556,I10349,I10219,I10507,I10490,I10052,I10366,I10332;
nand I_0(I7556,I7621,I7850);
and I_1(I10349,I10332,I7550);
DFFARX1 I_2(I10202,I1470,I10052,,,I10219,);
and I_3(I10507,I10490,I10366);
DFFARX1 I_4(I10507,I1470,I10052,,,I10044,);
DFFARX1 I_5(I7556,I1470,I10052,,,I10490,);
not I_6(I10052,I1477);
nand I_7(I10366,I10349,I10219);
DFFARX1 I_8(I1470,I10052,,,I10332,);
endmodule


