module Benchmark_testing1000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458,I2515,I2527,I2536,I2539,I2524,I2533,I2521,I2530,I2518);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458;
output I2515,I2527,I2536,I2539,I2524,I2533,I2521,I2530,I2518;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458,I1493,I14897,I1519,I1527,I1544,I14912,I14891,I1561,I14894,I1587,I14915,I1604,I1612,I1629,I1461,I1660,I1677,I1473,I1717,I1482,I1739,I14903,I14900,I1756,I14906,I1782,I1799,I1485,I1821,I1470,I1852,I14909,I1869,I1886,I1903,I1479,I1934,I1467,I1476,I1464,I2020,I11588,I2046,I2054,I2071,I11579,I11597,I2088,I11576,I2114,I2131,I2139,I11582,I2156,I1988,I2187,I2204,I2000,I2244,I2009,I2266,I11594,I11585,I2283,I11600,I2309,I2326,I2012,I2348,I1997,I2379,I11591,I2396,I2413,I2430,I2006,I2461,I1994,I2003,I1991,I2547,I3649,I2573,I2581,I2598,I3643,I3637,I2615,I3658,I2641,I3655,I2658,I2666,I3652,I2683,I2714,I2731,I2771,I2793,I3640,I2810,I3661,I2836,I2853,I2875,I2906,I3646,I2923,I2940,I2957,I2988,I3074,I3100,I3117,I3066,I3139,I3165,I3173,I3190,I3207,I3224,I3241,I3258,I3275,I3292,I3042,I3323,I3340,I3357,I3374,I3054,I3048,I3419,I3063,I3057,I3464,I3481,I3498,I3515,I3541,I3549,I3051,I3045,I3603,I3611,I3060,I3669,I5422,I3695,I3712,I3734,I5437,I3760,I3768,I3785,I5434,I3802,I3819,I3836,I5431,I3853,I5446,I3870,I5443,I3887,I3918,I3935,I3952,I3969,I4014,I5440,I4059,I4076,I5428,I4093,I5449,I4110,I5425,I4136,I4144,I4198,I4206,I4264,I8123,I4290,I4307,I4256,I4329,I8114,I4355,I4363,I4380,I8132,I4397,I8129,I4414,I4431,I8108,I4448,I8111,I4465,I8120,I4482,I4232,I4513,I4530,I4547,I4564,I4244,I4238,I4609,I8126,I4253,I4247,I4654,I4671,I4688,I8117,I4705,I4731,I4739,I4241,I4235,I4793,I4801,I4250,I4859,I4885,I4902,I4851,I4924,I4950,I4958,I4975,I4992,I5009,I5026,I5043,I5060,I5077,I4827,I5108,I5125,I5142,I5159,I4839,I4833,I5204,I4848,I4842,I5249,I5266,I5283,I5300,I5326,I5334,I4836,I4830,I5388,I5396,I4845,I5457,I17150,I5483,I5491,I17147,I17138,I5508,I17135,I5534,I5556,I17144,I5582,I5590,I17153,I5607,I5633,I5655,I17156,I5695,I5712,I5720,I5737,I5768,I17141,I5785,I17159,I5811,I5819,I5864,I5881,I5984,I7032,I6010,I6018,I7044,I7023,I6035,I7047,I6061,I5952,I6083,I7038,I6109,I6117,I7020,I6134,I6160,I5976,I6182,I5958,I7035,I6222,I6239,I6247,I6264,I5961,I6295,I7026,I6312,I7029,I6338,I6346,I5949,I5967,I6391,I7041,I6408,I5970,I5955,I5964,I5973,I6511,I9267,I6537,I6554,I6503,I6576,I6593,I9288,I9279,I6610,I6636,I6644,I9273,I6670,I6678,I9270,I6695,I6482,I9264,I6735,I6743,I6476,I6491,I6788,I9276,I6805,I9285,I6831,I6479,I6853,I6870,I6887,I6494,I6918,I6935,I9282,I6485,I6966,I6488,I6500,I6497,I7055,I11001,I7081,I7098,I7120,I7137,I11022,I11013,I7154,I7180,I7188,I11007,I7214,I7222,I11004,I7239,I10998,I7279,I7287,I7332,I11010,I7349,I11019,I7375,I7397,I7414,I7431,I7462,I7479,I11016,I7510,I7599,I16050,I7625,I7642,I7591,I7664,I7681,I16062,I16065,I7698,I16068,I7724,I7732,I16053,I7758,I7766,I16059,I7783,I7570,I16047,I7823,I7831,I7564,I7579,I7876,I16071,I7893,I16056,I7919,I7567,I7941,I7958,I7975,I7582,I8006,I8023,I7573,I8054,I7576,I7588,I7585,I8140,I9842,I8166,I8174,I9854,I8200,I8208,I9845,I8225,I9848,I8242,I8259,I9851,I8276,I8307,I8324,I8341,I8358,I9857,I8403,I8448,I9863,I8465,I8482,I8513,I8530,I9860,I8547,I9866,I8573,I8581,I8626,I8643,I8660,I8718,I12169,I8744,I8752,I8769,I12157,I12175,I8786,I12172,I8812,I8820,I12163,I12160,I8846,I8854,I8871,I8888,I8905,I8701,I12154,I8945,I8953,I8970,I8987,I9004,I8704,I9035,I9052,I9078,I9086,I8686,I9117,I8695,I9148,I9165,I8707,I9196,I12166,I8698,I8689,I8692,I8710,I9296,I9322,I9330,I9347,I9364,I9390,I9398,I9424,I9432,I9449,I9466,I9483,I9523,I9531,I9548,I9565,I9582,I9613,I9630,I9656,I9664,I9695,I9726,I9743,I9774,I9874,I9900,I9908,I9925,I9942,I9968,I9976,I10002,I10010,I10027,I10044,I10061,I10101,I10109,I10126,I10143,I10160,I10191,I10208,I10234,I10242,I10273,I10304,I10321,I10352,I10452,I10478,I10486,I10503,I10520,I10546,I10554,I10580,I10588,I10605,I10622,I10639,I10435,I10679,I10687,I10704,I10721,I10738,I10438,I10769,I10786,I10812,I10820,I10420,I10851,I10429,I10882,I10899,I10441,I10930,I10432,I10423,I10426,I10444,I11030,I11056,I11064,I11081,I11098,I11124,I11132,I11158,I11166,I11183,I11200,I11217,I11257,I11265,I11282,I11299,I11316,I11347,I11364,I11390,I11398,I11429,I11460,I11477,I11508,I11608,I15487,I11634,I11642,I11659,I15469,I15481,I11676,I15484,I11702,I11710,I15478,I15475,I11736,I11744,I11761,I11778,I11795,I15493,I11835,I11843,I11860,I11877,I11894,I11925,I15472,I11942,I11968,I11976,I12007,I12038,I12055,I12086,I15490,I12183,I14331,I12209,I12217,I12234,I14313,I12251,I14319,I12277,I14316,I12308,I12316,I14325,I12333,I12359,I12367,I14337,I12407,I12443,I14328,I14322,I12460,I12486,I12494,I12511,I12542,I14334,I12559,I12576,I12607,I12638,I12655,I12710,I12736,I12744,I12761,I12778,I12804,I12699,I12835,I12843,I12860,I12886,I12894,I12702,I12934,I12693,I12684,I12970,I12987,I13013,I13021,I13038,I12687,I13069,I13086,I13103,I12696,I13134,I12681,I13165,I13182,I12690,I13237,I13753,I13263,I13271,I13288,I13735,I13305,I13741,I13331,I13226,I13738,I13362,I13370,I13747,I13387,I13413,I13421,I13229,I13759,I13461,I13220,I13211,I13497,I13750,I13744,I13514,I13540,I13548,I13565,I13214,I13596,I13756,I13613,I13630,I13223,I13661,I13208,I13692,I13709,I13217,I13767,I13793,I13801,I13841,I13849,I13866,I13883,I13923,I13945,I13962,I13988,I13996,I14013,I14030,I14047,I14064,I14109,I14140,I14157,I14183,I14191,I14222,I14239,I14256,I14273,I14345,I14371,I14379,I14419,I14427,I14444,I14461,I14501,I14523,I14540,I14566,I14574,I14591,I14608,I14625,I14642,I14687,I14718,I14735,I14761,I14769,I14800,I14817,I14834,I14851,I14923,I14949,I14957,I14997,I15005,I15022,I15039,I15079,I15101,I15118,I15144,I15152,I15169,I15186,I15203,I15220,I15265,I15296,I15313,I15339,I15347,I15378,I15395,I15412,I15429,I15501,I16612,I15527,I15535,I16606,I16591,I15575,I15583,I16597,I15600,I16609,I15617,I15657,I15679,I15696,I15722,I15730,I15747,I16615,I15764,I16603,I15781,I15798,I15843,I16594,I15874,I15891,I16600,I15917,I15925,I15956,I15973,I15990,I16007,I16079,I16105,I16113,I16139,I16156,I16178,I16195,I16212,I16229,I16246,I16277,I16294,I16311,I16328,I16373,I16390,I16407,I16466,I16492,I16500,I16517,I16534,I16565,I16623,I16649,I16657,I16683,I16700,I16722,I16739,I16756,I16773,I16790,I16821,I16838,I16855,I16872,I16917,I16934,I16951,I17010,I17036,I17044,I17061,I17078,I17109,I17167,I17193,I17201,I17218,I17244,I17252,I17269,I17286,I17303,I17320,I17351,I17368,I17385,I17416,I17433,I17473,I17481,I17512,I17529,I17546,I17563,I17594,I17625,I17651,I17673;
not I_0 (I1493,I1458);
DFFARX1 I_1 (I14897,I1451,I1493,I1519,);
not I_2 (I1527,I1519);
nand I_3 (I1544,I14912,I14891);
and I_4 (I1561,I1544,I14894);
DFFARX1 I_5 (I1561,I1451,I1493,I1587,);
DFFARX1 I_6 (I14915,I1451,I1493,I1604,);
and I_7 (I1612,I1604,I14894);
nor I_8 (I1629,I1587,I1612);
DFFARX1 I_9 (I1629,I1451,I1493,I1461,);
nand I_10 (I1660,I1604,I14894);
nand I_11 (I1677,I1527,I1660);
not I_12 (I1473,I1677);
DFFARX1 I_13 (I14891,I1451,I1493,I1717,);
DFFARX1 I_14 (I1717,I1451,I1493,I1482,);
nand I_15 (I1739,I14903,I14900);
and I_16 (I1756,I1739,I14906);
DFFARX1 I_17 (I1756,I1451,I1493,I1782,);
DFFARX1 I_18 (I1782,I1451,I1493,I1799,);
not I_19 (I1485,I1799);
not I_20 (I1821,I1782);
nand I_21 (I1470,I1821,I1660);
nor I_22 (I1852,I14909,I14900);
not I_23 (I1869,I1852);
nor I_24 (I1886,I1821,I1869);
nor I_25 (I1903,I1527,I1886);
DFFARX1 I_26 (I1903,I1451,I1493,I1479,);
nor I_27 (I1934,I1587,I1869);
nor I_28 (I1467,I1782,I1934);
nor I_29 (I1476,I1717,I1852);
nor I_30 (I1464,I1587,I1852);
not I_31 (I2020,I1458);
DFFARX1 I_32 (I11588,I1451,I2020,I2046,);
not I_33 (I2054,I2046);
nand I_34 (I2071,I11579,I11597);
and I_35 (I2088,I2071,I11576);
DFFARX1 I_36 (I2088,I1451,I2020,I2114,);
DFFARX1 I_37 (I11579,I1451,I2020,I2131,);
and I_38 (I2139,I2131,I11582);
nor I_39 (I2156,I2114,I2139);
DFFARX1 I_40 (I2156,I1451,I2020,I1988,);
nand I_41 (I2187,I2131,I11582);
nand I_42 (I2204,I2054,I2187);
not I_43 (I2000,I2204);
DFFARX1 I_44 (I11576,I1451,I2020,I2244,);
DFFARX1 I_45 (I2244,I1451,I2020,I2009,);
nand I_46 (I2266,I11594,I11585);
and I_47 (I2283,I2266,I11600);
DFFARX1 I_48 (I2283,I1451,I2020,I2309,);
DFFARX1 I_49 (I2309,I1451,I2020,I2326,);
not I_50 (I2012,I2326);
not I_51 (I2348,I2309);
nand I_52 (I1997,I2348,I2187);
nor I_53 (I2379,I11591,I11585);
not I_54 (I2396,I2379);
nor I_55 (I2413,I2348,I2396);
nor I_56 (I2430,I2054,I2413);
DFFARX1 I_57 (I2430,I1451,I2020,I2006,);
nor I_58 (I2461,I2114,I2396);
nor I_59 (I1994,I2309,I2461);
nor I_60 (I2003,I2244,I2379);
nor I_61 (I1991,I2114,I2379);
not I_62 (I2547,I1458);
DFFARX1 I_63 (I3649,I1451,I2547,I2573,);
not I_64 (I2581,I2573);
nand I_65 (I2598,I3643,I3637);
and I_66 (I2615,I2598,I3658);
DFFARX1 I_67 (I2615,I1451,I2547,I2641,);
DFFARX1 I_68 (I3655,I1451,I2547,I2658,);
and I_69 (I2666,I2658,I3652);
nor I_70 (I2683,I2641,I2666);
DFFARX1 I_71 (I2683,I1451,I2547,I2515,);
nand I_72 (I2714,I2658,I3652);
nand I_73 (I2731,I2581,I2714);
not I_74 (I2527,I2731);
DFFARX1 I_75 (I3637,I1451,I2547,I2771,);
DFFARX1 I_76 (I2771,I1451,I2547,I2536,);
nand I_77 (I2793,I3640,I3640);
and I_78 (I2810,I2793,I3661);
DFFARX1 I_79 (I2810,I1451,I2547,I2836,);
DFFARX1 I_80 (I2836,I1451,I2547,I2853,);
not I_81 (I2539,I2853);
not I_82 (I2875,I2836);
nand I_83 (I2524,I2875,I2714);
nor I_84 (I2906,I3646,I3640);
not I_85 (I2923,I2906);
nor I_86 (I2940,I2875,I2923);
nor I_87 (I2957,I2581,I2940);
DFFARX1 I_88 (I2957,I1451,I2547,I2533,);
nor I_89 (I2988,I2641,I2923);
nor I_90 (I2521,I2836,I2988);
nor I_91 (I2530,I2771,I2906);
nor I_92 (I2518,I2641,I2906);
not I_93 (I3074,I1458);
DFFARX1 I_94 (I1997,I1451,I3074,I3100,);
DFFARX1 I_95 (I3100,I1451,I3074,I3117,);
not I_96 (I3066,I3117);
not I_97 (I3139,I3100);
DFFARX1 I_98 (I1991,I1451,I3074,I3165,);
not I_99 (I3173,I3165);
and I_100 (I3190,I3139,I1988);
not I_101 (I3207,I2009);
nand I_102 (I3224,I3207,I1988);
not I_103 (I3241,I2003);
nor I_104 (I3258,I3241,I1994);
nand I_105 (I3275,I3258,I2000);
nor I_106 (I3292,I3275,I3224);
DFFARX1 I_107 (I3292,I1451,I3074,I3042,);
not I_108 (I3323,I3275);
not I_109 (I3340,I1994);
nand I_110 (I3357,I3340,I1988);
nor I_111 (I3374,I1994,I2009);
nand I_112 (I3054,I3190,I3374);
nand I_113 (I3048,I3139,I1994);
nand I_114 (I3419,I3241,I1988);
DFFARX1 I_115 (I3419,I1451,I3074,I3063,);
DFFARX1 I_116 (I3419,I1451,I3074,I3057,);
not I_117 (I3464,I1988);
nor I_118 (I3481,I3464,I2006);
and I_119 (I3498,I3481,I2012);
or I_120 (I3515,I3498,I1991);
DFFARX1 I_121 (I3515,I1451,I3074,I3541,);
nand I_122 (I3549,I3541,I3207);
nor I_123 (I3051,I3549,I3357);
nor I_124 (I3045,I3541,I3173);
DFFARX1 I_125 (I3541,I1451,I3074,I3603,);
not I_126 (I3611,I3603);
nor I_127 (I3060,I3611,I3323);
not I_128 (I3669,I1458);
DFFARX1 I_129 (I5422,I1451,I3669,I3695,);
DFFARX1 I_130 (I3695,I1451,I3669,I3712,);
not I_131 (I3661,I3712);
not I_132 (I3734,I3695);
DFFARX1 I_133 (I5437,I1451,I3669,I3760,);
not I_134 (I3768,I3760);
and I_135 (I3785,I3734,I5434);
not I_136 (I3802,I5422);
nand I_137 (I3819,I3802,I5434);
not I_138 (I3836,I5431);
nor I_139 (I3853,I3836,I5446);
nand I_140 (I3870,I3853,I5443);
nor I_141 (I3887,I3870,I3819);
DFFARX1 I_142 (I3887,I1451,I3669,I3637,);
not I_143 (I3918,I3870);
not I_144 (I3935,I5446);
nand I_145 (I3952,I3935,I5434);
nor I_146 (I3969,I5446,I5422);
nand I_147 (I3649,I3785,I3969);
nand I_148 (I3643,I3734,I5446);
nand I_149 (I4014,I3836,I5440);
DFFARX1 I_150 (I4014,I1451,I3669,I3658,);
DFFARX1 I_151 (I4014,I1451,I3669,I3652,);
not I_152 (I4059,I5440);
nor I_153 (I4076,I4059,I5428);
and I_154 (I4093,I4076,I5449);
or I_155 (I4110,I4093,I5425);
DFFARX1 I_156 (I4110,I1451,I3669,I4136,);
nand I_157 (I4144,I4136,I3802);
nor I_158 (I3646,I4144,I3952);
nor I_159 (I3640,I4136,I3768);
DFFARX1 I_160 (I4136,I1451,I3669,I4198,);
not I_161 (I4206,I4198);
nor I_162 (I3655,I4206,I3918);
not I_163 (I4264,I1458);
DFFARX1 I_164 (I8123,I1451,I4264,I4290,);
DFFARX1 I_165 (I4290,I1451,I4264,I4307,);
not I_166 (I4256,I4307);
not I_167 (I4329,I4290);
DFFARX1 I_168 (I8114,I1451,I4264,I4355,);
not I_169 (I4363,I4355);
and I_170 (I4380,I4329,I8132);
not I_171 (I4397,I8129);
nand I_172 (I4414,I4397,I8132);
not I_173 (I4431,I8108);
nor I_174 (I4448,I4431,I8111);
nand I_175 (I4465,I4448,I8120);
nor I_176 (I4482,I4465,I4414);
DFFARX1 I_177 (I4482,I1451,I4264,I4232,);
not I_178 (I4513,I4465);
not I_179 (I4530,I8111);
nand I_180 (I4547,I4530,I8132);
nor I_181 (I4564,I8111,I8129);
nand I_182 (I4244,I4380,I4564);
nand I_183 (I4238,I4329,I8111);
nand I_184 (I4609,I4431,I8126);
DFFARX1 I_185 (I4609,I1451,I4264,I4253,);
DFFARX1 I_186 (I4609,I1451,I4264,I4247,);
not I_187 (I4654,I8126);
nor I_188 (I4671,I4654,I8108);
and I_189 (I4688,I4671,I8117);
or I_190 (I4705,I4688,I8111);
DFFARX1 I_191 (I4705,I1451,I4264,I4731,);
nand I_192 (I4739,I4731,I4397);
nor I_193 (I4241,I4739,I4547);
nor I_194 (I4235,I4731,I4363);
DFFARX1 I_195 (I4731,I1451,I4264,I4793,);
not I_196 (I4801,I4793);
nor I_197 (I4250,I4801,I4513);
not I_198 (I4859,I1458);
DFFARX1 I_199 (I1470,I1451,I4859,I4885,);
DFFARX1 I_200 (I4885,I1451,I4859,I4902,);
not I_201 (I4851,I4902);
not I_202 (I4924,I4885);
DFFARX1 I_203 (I1464,I1451,I4859,I4950,);
not I_204 (I4958,I4950);
and I_205 (I4975,I4924,I1461);
not I_206 (I4992,I1482);
nand I_207 (I5009,I4992,I1461);
not I_208 (I5026,I1476);
nor I_209 (I5043,I5026,I1467);
nand I_210 (I5060,I5043,I1473);
nor I_211 (I5077,I5060,I5009);
DFFARX1 I_212 (I5077,I1451,I4859,I4827,);
not I_213 (I5108,I5060);
not I_214 (I5125,I1467);
nand I_215 (I5142,I5125,I1461);
nor I_216 (I5159,I1467,I1482);
nand I_217 (I4839,I4975,I5159);
nand I_218 (I4833,I4924,I1467);
nand I_219 (I5204,I5026,I1461);
DFFARX1 I_220 (I5204,I1451,I4859,I4848,);
DFFARX1 I_221 (I5204,I1451,I4859,I4842,);
not I_222 (I5249,I1461);
nor I_223 (I5266,I5249,I1479);
and I_224 (I5283,I5266,I1485);
or I_225 (I5300,I5283,I1464);
DFFARX1 I_226 (I5300,I1451,I4859,I5326,);
nand I_227 (I5334,I5326,I4992);
nor I_228 (I4836,I5334,I5142);
nor I_229 (I4830,I5326,I4958);
DFFARX1 I_230 (I5326,I1451,I4859,I5388,);
not I_231 (I5396,I5388);
nor I_232 (I4845,I5396,I5108);
not I_233 (I5457,I1458);
DFFARX1 I_234 (I17150,I1451,I5457,I5483,);
nand I_235 (I5491,I17147,I17138);
and I_236 (I5508,I5491,I17135);
DFFARX1 I_237 (I5508,I1451,I5457,I5534,);
nor I_238 (I5425,I5534,I5483);
not I_239 (I5556,I5534);
DFFARX1 I_240 (I17144,I1451,I5457,I5582,);
nand I_241 (I5590,I5582,I17153);
not I_242 (I5607,I5590);
DFFARX1 I_243 (I5607,I1451,I5457,I5633,);
not I_244 (I5449,I5633);
nor I_245 (I5655,I5483,I5590);
nor I_246 (I5431,I5534,I5655);
DFFARX1 I_247 (I17156,I1451,I5457,I5695,);
DFFARX1 I_248 (I5695,I1451,I5457,I5712,);
not I_249 (I5720,I5712);
not I_250 (I5737,I5695);
nand I_251 (I5434,I5737,I5556);
nand I_252 (I5768,I17135,I17141);
and I_253 (I5785,I5768,I17159);
DFFARX1 I_254 (I5785,I1451,I5457,I5811,);
nor I_255 (I5819,I5811,I5483);
DFFARX1 I_256 (I5819,I1451,I5457,I5422,);
DFFARX1 I_257 (I5811,I1451,I5457,I5440,);
nor I_258 (I5864,I17138,I17141);
not I_259 (I5881,I5864);
nor I_260 (I5443,I5720,I5881);
nand I_261 (I5428,I5737,I5881);
nor I_262 (I5437,I5483,I5864);
DFFARX1 I_263 (I5864,I1451,I5457,I5446,);
not I_264 (I5984,I1458);
DFFARX1 I_265 (I7032,I1451,I5984,I6010,);
nand I_266 (I6018,I7044,I7023);
and I_267 (I6035,I6018,I7047);
DFFARX1 I_268 (I6035,I1451,I5984,I6061,);
nor I_269 (I5952,I6061,I6010);
not I_270 (I6083,I6061);
DFFARX1 I_271 (I7038,I1451,I5984,I6109,);
nand I_272 (I6117,I6109,I7020);
not I_273 (I6134,I6117);
DFFARX1 I_274 (I6134,I1451,I5984,I6160,);
not I_275 (I5976,I6160);
nor I_276 (I6182,I6010,I6117);
nor I_277 (I5958,I6061,I6182);
DFFARX1 I_278 (I7035,I1451,I5984,I6222,);
DFFARX1 I_279 (I6222,I1451,I5984,I6239,);
not I_280 (I6247,I6239);
not I_281 (I6264,I6222);
nand I_282 (I5961,I6264,I6083);
nand I_283 (I6295,I7020,I7026);
and I_284 (I6312,I6295,I7029);
DFFARX1 I_285 (I6312,I1451,I5984,I6338,);
nor I_286 (I6346,I6338,I6010);
DFFARX1 I_287 (I6346,I1451,I5984,I5949,);
DFFARX1 I_288 (I6338,I1451,I5984,I5967,);
nor I_289 (I6391,I7041,I7026);
not I_290 (I6408,I6391);
nor I_291 (I5970,I6247,I6408);
nand I_292 (I5955,I6264,I6408);
nor I_293 (I5964,I6010,I6391);
DFFARX1 I_294 (I6391,I1451,I5984,I5973,);
not I_295 (I6511,I1458);
DFFARX1 I_296 (I9267,I1451,I6511,I6537,);
DFFARX1 I_297 (I6537,I1451,I6511,I6554,);
not I_298 (I6503,I6554);
not I_299 (I6576,I6537);
nand I_300 (I6593,I9288,I9279);
and I_301 (I6610,I6593,I9267);
DFFARX1 I_302 (I6610,I1451,I6511,I6636,);
not I_303 (I6644,I6636);
DFFARX1 I_304 (I9273,I1451,I6511,I6670,);
and I_305 (I6678,I6670,I9270);
nand I_306 (I6695,I6670,I9270);
nand I_307 (I6482,I6644,I6695);
DFFARX1 I_308 (I9264,I1451,I6511,I6735,);
nor I_309 (I6743,I6735,I6678);
DFFARX1 I_310 (I6743,I1451,I6511,I6476,);
nor I_311 (I6491,I6735,I6636);
nand I_312 (I6788,I9264,I9276);
and I_313 (I6805,I6788,I9285);
DFFARX1 I_314 (I6805,I1451,I6511,I6831,);
nor I_315 (I6479,I6831,I6735);
not I_316 (I6853,I6831);
nor I_317 (I6870,I6853,I6644);
nor I_318 (I6887,I6576,I6870);
DFFARX1 I_319 (I6887,I1451,I6511,I6494,);
nor I_320 (I6918,I6853,I6735);
nor I_321 (I6935,I9282,I9276);
nor I_322 (I6485,I6935,I6918);
not I_323 (I6966,I6935);
nand I_324 (I6488,I6695,I6966);
DFFARX1 I_325 (I6935,I1451,I6511,I6500,);
DFFARX1 I_326 (I6935,I1451,I6511,I6497,);
not I_327 (I7055,I1458);
DFFARX1 I_328 (I11001,I1451,I7055,I7081,);
DFFARX1 I_329 (I7081,I1451,I7055,I7098,);
not I_330 (I7047,I7098);
not I_331 (I7120,I7081);
nand I_332 (I7137,I11022,I11013);
and I_333 (I7154,I7137,I11001);
DFFARX1 I_334 (I7154,I1451,I7055,I7180,);
not I_335 (I7188,I7180);
DFFARX1 I_336 (I11007,I1451,I7055,I7214,);
and I_337 (I7222,I7214,I11004);
nand I_338 (I7239,I7214,I11004);
nand I_339 (I7026,I7188,I7239);
DFFARX1 I_340 (I10998,I1451,I7055,I7279,);
nor I_341 (I7287,I7279,I7222);
DFFARX1 I_342 (I7287,I1451,I7055,I7020,);
nor I_343 (I7035,I7279,I7180);
nand I_344 (I7332,I10998,I11010);
and I_345 (I7349,I7332,I11019);
DFFARX1 I_346 (I7349,I1451,I7055,I7375,);
nor I_347 (I7023,I7375,I7279);
not I_348 (I7397,I7375);
nor I_349 (I7414,I7397,I7188);
nor I_350 (I7431,I7120,I7414);
DFFARX1 I_351 (I7431,I1451,I7055,I7038,);
nor I_352 (I7462,I7397,I7279);
nor I_353 (I7479,I11016,I11010);
nor I_354 (I7029,I7479,I7462);
not I_355 (I7510,I7479);
nand I_356 (I7032,I7239,I7510);
DFFARX1 I_357 (I7479,I1451,I7055,I7044,);
DFFARX1 I_358 (I7479,I1451,I7055,I7041,);
not I_359 (I7599,I1458);
DFFARX1 I_360 (I16050,I1451,I7599,I7625,);
DFFARX1 I_361 (I7625,I1451,I7599,I7642,);
not I_362 (I7591,I7642);
not I_363 (I7664,I7625);
nand I_364 (I7681,I16062,I16065);
and I_365 (I7698,I7681,I16068);
DFFARX1 I_366 (I7698,I1451,I7599,I7724,);
not I_367 (I7732,I7724);
DFFARX1 I_368 (I16053,I1451,I7599,I7758,);
and I_369 (I7766,I7758,I16059);
nand I_370 (I7783,I7758,I16059);
nand I_371 (I7570,I7732,I7783);
DFFARX1 I_372 (I16047,I1451,I7599,I7823,);
nor I_373 (I7831,I7823,I7766);
DFFARX1 I_374 (I7831,I1451,I7599,I7564,);
nor I_375 (I7579,I7823,I7724);
nand I_376 (I7876,I16050,I16071);
and I_377 (I7893,I7876,I16056);
DFFARX1 I_378 (I7893,I1451,I7599,I7919,);
nor I_379 (I7567,I7919,I7823);
not I_380 (I7941,I7919);
nor I_381 (I7958,I7941,I7732);
nor I_382 (I7975,I7664,I7958);
DFFARX1 I_383 (I7975,I1451,I7599,I7582,);
nor I_384 (I8006,I7941,I7823);
nor I_385 (I8023,I16047,I16071);
nor I_386 (I7573,I8023,I8006);
not I_387 (I8054,I8023);
nand I_388 (I7576,I7783,I8054);
DFFARX1 I_389 (I8023,I1451,I7599,I7588,);
DFFARX1 I_390 (I8023,I1451,I7599,I7585,);
not I_391 (I8140,I1458);
DFFARX1 I_392 (I9842,I1451,I8140,I8166,);
not I_393 (I8174,I8166);
DFFARX1 I_394 (I9854,I1451,I8140,I8200,);
not I_395 (I8208,I9845);
nand I_396 (I8225,I8208,I9848);
not I_397 (I8242,I8225);
nor I_398 (I8259,I8242,I9851);
nor I_399 (I8276,I8174,I8259);
DFFARX1 I_400 (I8276,I1451,I8140,I8126,);
not I_401 (I8307,I9851);
nand I_402 (I8324,I8307,I8242);
and I_403 (I8341,I8307,I9845);
nand I_404 (I8358,I8341,I9857);
nor I_405 (I8123,I8358,I8307);
and I_406 (I8114,I8200,I8358);
not I_407 (I8403,I8358);
nand I_408 (I8117,I8200,I8403);
nor I_409 (I8111,I8166,I8358);
not I_410 (I8448,I9863);
nor I_411 (I8465,I8448,I9845);
nand I_412 (I8482,I8465,I8307);
nor I_413 (I8120,I8225,I8482);
nor I_414 (I8513,I8448,I9842);
and I_415 (I8530,I8513,I9860);
or I_416 (I8547,I8530,I9866);
DFFARX1 I_417 (I8547,I1451,I8140,I8573,);
nor I_418 (I8581,I8573,I8324);
DFFARX1 I_419 (I8581,I1451,I8140,I8108,);
DFFARX1 I_420 (I8573,I1451,I8140,I8132,);
not I_421 (I8626,I8573);
nor I_422 (I8643,I8626,I8200);
nor I_423 (I8660,I8465,I8643);
DFFARX1 I_424 (I8660,I1451,I8140,I8129,);
not I_425 (I8718,I1458);
DFFARX1 I_426 (I12169,I1451,I8718,I8744,);
not I_427 (I8752,I8744);
nand I_428 (I8769,I12157,I12175);
and I_429 (I8786,I8769,I12172);
DFFARX1 I_430 (I8786,I1451,I8718,I8812,);
not I_431 (I8820,I12163);
DFFARX1 I_432 (I12160,I1451,I8718,I8846,);
not I_433 (I8854,I8846);
nor I_434 (I8871,I8854,I8752);
and I_435 (I8888,I8871,I12163);
nor I_436 (I8905,I8854,I8820);
nor I_437 (I8701,I8812,I8905);
DFFARX1 I_438 (I12154,I1451,I8718,I8945,);
nor I_439 (I8953,I8945,I8812);
not I_440 (I8970,I8953);
not I_441 (I8987,I8945);
nor I_442 (I9004,I8987,I8888);
DFFARX1 I_443 (I9004,I1451,I8718,I8704,);
nand I_444 (I9035,I12154,I12157);
and I_445 (I9052,I9035,I12160);
DFFARX1 I_446 (I9052,I1451,I8718,I9078,);
nor I_447 (I9086,I9078,I8945);
DFFARX1 I_448 (I9086,I1451,I8718,I8686,);
nand I_449 (I9117,I9078,I8987);
nand I_450 (I8695,I8970,I9117);
not I_451 (I9148,I9078);
nor I_452 (I9165,I9148,I8888);
DFFARX1 I_453 (I9165,I1451,I8718,I8707,);
nor I_454 (I9196,I12166,I12157);
or I_455 (I8698,I8945,I9196);
nor I_456 (I8689,I9078,I9196);
or I_457 (I8692,I8812,I9196);
DFFARX1 I_458 (I9196,I1451,I8718,I8710,);
not I_459 (I9296,I1458);
DFFARX1 I_460 (I7573,I1451,I9296,I9322,);
not I_461 (I9330,I9322);
nand I_462 (I9347,I7564,I7582);
and I_463 (I9364,I9347,I7585);
DFFARX1 I_464 (I9364,I1451,I9296,I9390,);
not I_465 (I9398,I7579);
DFFARX1 I_466 (I7567,I1451,I9296,I9424,);
not I_467 (I9432,I9424);
nor I_468 (I9449,I9432,I9330);
and I_469 (I9466,I9449,I7579);
nor I_470 (I9483,I9432,I9398);
nor I_471 (I9279,I9390,I9483);
DFFARX1 I_472 (I7576,I1451,I9296,I9523,);
nor I_473 (I9531,I9523,I9390);
not I_474 (I9548,I9531);
not I_475 (I9565,I9523);
nor I_476 (I9582,I9565,I9466);
DFFARX1 I_477 (I9582,I1451,I9296,I9282,);
nand I_478 (I9613,I7591,I7588);
and I_479 (I9630,I9613,I7570);
DFFARX1 I_480 (I9630,I1451,I9296,I9656,);
nor I_481 (I9664,I9656,I9523);
DFFARX1 I_482 (I9664,I1451,I9296,I9264,);
nand I_483 (I9695,I9656,I9565);
nand I_484 (I9273,I9548,I9695);
not I_485 (I9726,I9656);
nor I_486 (I9743,I9726,I9466);
DFFARX1 I_487 (I9743,I1451,I9296,I9285,);
nor I_488 (I9774,I7564,I7588);
or I_489 (I9276,I9523,I9774);
nor I_490 (I9267,I9656,I9774);
or I_491 (I9270,I9390,I9774);
DFFARX1 I_492 (I9774,I1451,I9296,I9288,);
not I_493 (I9874,I1458);
DFFARX1 I_494 (I1364,I1451,I9874,I9900,);
not I_495 (I9908,I9900);
nand I_496 (I9925,I1396,I1404);
and I_497 (I9942,I9925,I1380);
DFFARX1 I_498 (I9942,I1451,I9874,I9968,);
not I_499 (I9976,I1388);
DFFARX1 I_500 (I1428,I1451,I9874,I10002,);
not I_501 (I10010,I10002);
nor I_502 (I10027,I10010,I9908);
and I_503 (I10044,I10027,I1388);
nor I_504 (I10061,I10010,I9976);
nor I_505 (I9857,I9968,I10061);
DFFARX1 I_506 (I1412,I1451,I9874,I10101,);
nor I_507 (I10109,I10101,I9968);
not I_508 (I10126,I10109);
not I_509 (I10143,I10101);
nor I_510 (I10160,I10143,I10044);
DFFARX1 I_511 (I10160,I1451,I9874,I9860,);
nand I_512 (I10191,I1444,I1436);
and I_513 (I10208,I10191,I1420);
DFFARX1 I_514 (I10208,I1451,I9874,I10234,);
nor I_515 (I10242,I10234,I10101);
DFFARX1 I_516 (I10242,I1451,I9874,I9842,);
nand I_517 (I10273,I10234,I10143);
nand I_518 (I9851,I10126,I10273);
not I_519 (I10304,I10234);
nor I_520 (I10321,I10304,I10044);
DFFARX1 I_521 (I10321,I1451,I9874,I9863,);
nor I_522 (I10352,I1372,I1436);
or I_523 (I9854,I10101,I10352);
nor I_524 (I9845,I10234,I10352);
or I_525 (I9848,I9968,I10352);
DFFARX1 I_526 (I10352,I1451,I9874,I9866,);
not I_527 (I10452,I1458);
DFFARX1 I_528 (I4232,I1451,I10452,I10478,);
not I_529 (I10486,I10478);
nand I_530 (I10503,I4235,I4256);
and I_531 (I10520,I10503,I4244);
DFFARX1 I_532 (I10520,I1451,I10452,I10546,);
not I_533 (I10554,I4241);
DFFARX1 I_534 (I4232,I1451,I10452,I10580,);
not I_535 (I10588,I10580);
nor I_536 (I10605,I10588,I10486);
and I_537 (I10622,I10605,I4241);
nor I_538 (I10639,I10588,I10554);
nor I_539 (I10435,I10546,I10639);
DFFARX1 I_540 (I4250,I1451,I10452,I10679,);
nor I_541 (I10687,I10679,I10546);
not I_542 (I10704,I10687);
not I_543 (I10721,I10679);
nor I_544 (I10738,I10721,I10622);
DFFARX1 I_545 (I10738,I1451,I10452,I10438,);
nand I_546 (I10769,I4235,I4238);
and I_547 (I10786,I10769,I4247);
DFFARX1 I_548 (I10786,I1451,I10452,I10812,);
nor I_549 (I10820,I10812,I10679);
DFFARX1 I_550 (I10820,I1451,I10452,I10420,);
nand I_551 (I10851,I10812,I10721);
nand I_552 (I10429,I10704,I10851);
not I_553 (I10882,I10812);
nor I_554 (I10899,I10882,I10622);
DFFARX1 I_555 (I10899,I1451,I10452,I10441,);
nor I_556 (I10930,I4253,I4238);
or I_557 (I10432,I10679,I10930);
nor I_558 (I10423,I10812,I10930);
or I_559 (I10426,I10546,I10930);
DFFARX1 I_560 (I10930,I1451,I10452,I10444,);
not I_561 (I11030,I1458);
DFFARX1 I_562 (I4827,I1451,I11030,I11056,);
not I_563 (I11064,I11056);
nand I_564 (I11081,I4830,I4851);
and I_565 (I11098,I11081,I4839);
DFFARX1 I_566 (I11098,I1451,I11030,I11124,);
not I_567 (I11132,I4836);
DFFARX1 I_568 (I4827,I1451,I11030,I11158,);
not I_569 (I11166,I11158);
nor I_570 (I11183,I11166,I11064);
and I_571 (I11200,I11183,I4836);
nor I_572 (I11217,I11166,I11132);
nor I_573 (I11013,I11124,I11217);
DFFARX1 I_574 (I4845,I1451,I11030,I11257,);
nor I_575 (I11265,I11257,I11124);
not I_576 (I11282,I11265);
not I_577 (I11299,I11257);
nor I_578 (I11316,I11299,I11200);
DFFARX1 I_579 (I11316,I1451,I11030,I11016,);
nand I_580 (I11347,I4830,I4833);
and I_581 (I11364,I11347,I4842);
DFFARX1 I_582 (I11364,I1451,I11030,I11390,);
nor I_583 (I11398,I11390,I11257);
DFFARX1 I_584 (I11398,I1451,I11030,I10998,);
nand I_585 (I11429,I11390,I11299);
nand I_586 (I11007,I11282,I11429);
not I_587 (I11460,I11390);
nor I_588 (I11477,I11460,I11200);
DFFARX1 I_589 (I11477,I1451,I11030,I11019,);
nor I_590 (I11508,I4848,I4833);
or I_591 (I11010,I11257,I11508);
nor I_592 (I11001,I11390,I11508);
or I_593 (I11004,I11124,I11508);
DFFARX1 I_594 (I11508,I1451,I11030,I11022,);
not I_595 (I11608,I1458);
DFFARX1 I_596 (I15487,I1451,I11608,I11634,);
not I_597 (I11642,I11634);
nand I_598 (I11659,I15469,I15481);
and I_599 (I11676,I11659,I15484);
DFFARX1 I_600 (I11676,I1451,I11608,I11702,);
not I_601 (I11710,I15478);
DFFARX1 I_602 (I15475,I1451,I11608,I11736,);
not I_603 (I11744,I11736);
nor I_604 (I11761,I11744,I11642);
and I_605 (I11778,I11761,I15478);
nor I_606 (I11795,I11744,I11710);
nor I_607 (I11591,I11702,I11795);
DFFARX1 I_608 (I15493,I1451,I11608,I11835,);
nor I_609 (I11843,I11835,I11702);
not I_610 (I11860,I11843);
not I_611 (I11877,I11835);
nor I_612 (I11894,I11877,I11778);
DFFARX1 I_613 (I11894,I1451,I11608,I11594,);
nand I_614 (I11925,I15472,I15472);
and I_615 (I11942,I11925,I15469);
DFFARX1 I_616 (I11942,I1451,I11608,I11968,);
nor I_617 (I11976,I11968,I11835);
DFFARX1 I_618 (I11976,I1451,I11608,I11576,);
nand I_619 (I12007,I11968,I11877);
nand I_620 (I11585,I11860,I12007);
not I_621 (I12038,I11968);
nor I_622 (I12055,I12038,I11778);
DFFARX1 I_623 (I12055,I1451,I11608,I11597,);
nor I_624 (I12086,I15490,I15472);
or I_625 (I11588,I11835,I12086);
nor I_626 (I11579,I11968,I12086);
or I_627 (I11582,I11702,I12086);
DFFARX1 I_628 (I12086,I1451,I11608,I11600,);
not I_629 (I12183,I1458);
DFFARX1 I_630 (I14331,I1451,I12183,I12209,);
not I_631 (I12217,I12209);
nand I_632 (I12234,I14313,I14313);
and I_633 (I12251,I12234,I14319);
DFFARX1 I_634 (I12251,I1451,I12183,I12277,);
DFFARX1 I_635 (I12277,I1451,I12183,I12172,);
DFFARX1 I_636 (I14316,I1451,I12183,I12308,);
nand I_637 (I12316,I12308,I14325);
not I_638 (I12333,I12316);
DFFARX1 I_639 (I12333,I1451,I12183,I12359,);
not I_640 (I12367,I12359);
nor I_641 (I12175,I12217,I12367);
DFFARX1 I_642 (I14337,I1451,I12183,I12407,);
nor I_643 (I12166,I12407,I12277);
nor I_644 (I12157,I12407,I12333);
nand I_645 (I12443,I14328,I14322);
and I_646 (I12460,I12443,I14316);
DFFARX1 I_647 (I12460,I1451,I12183,I12486,);
not I_648 (I12494,I12486);
nand I_649 (I12511,I12494,I12407);
nand I_650 (I12160,I12494,I12316);
nor I_651 (I12542,I14334,I14322);
and I_652 (I12559,I12407,I12542);
nor I_653 (I12576,I12494,I12559);
DFFARX1 I_654 (I12576,I1451,I12183,I12169,);
nor I_655 (I12607,I12209,I12542);
DFFARX1 I_656 (I12607,I1451,I12183,I12154,);
nor I_657 (I12638,I12486,I12542);
not I_658 (I12655,I12638);
nand I_659 (I12163,I12655,I12511);
not I_660 (I12710,I1458);
DFFARX1 I_661 (I3048,I1451,I12710,I12736,);
not I_662 (I12744,I12736);
nand I_663 (I12761,I3045,I3063);
and I_664 (I12778,I12761,I3054);
DFFARX1 I_665 (I12778,I1451,I12710,I12804,);
DFFARX1 I_666 (I12804,I1451,I12710,I12699,);
DFFARX1 I_667 (I3060,I1451,I12710,I12835,);
nand I_668 (I12843,I12835,I3057);
not I_669 (I12860,I12843);
DFFARX1 I_670 (I12860,I1451,I12710,I12886,);
not I_671 (I12894,I12886);
nor I_672 (I12702,I12744,I12894);
DFFARX1 I_673 (I3051,I1451,I12710,I12934,);
nor I_674 (I12693,I12934,I12804);
nor I_675 (I12684,I12934,I12860);
nand I_676 (I12970,I3042,I3066);
and I_677 (I12987,I12970,I3045);
DFFARX1 I_678 (I12987,I1451,I12710,I13013,);
not I_679 (I13021,I13013);
nand I_680 (I13038,I13021,I12934);
nand I_681 (I12687,I13021,I12843);
nor I_682 (I13069,I3042,I3066);
and I_683 (I13086,I12934,I13069);
nor I_684 (I13103,I13021,I13086);
DFFARX1 I_685 (I13103,I1451,I12710,I12696,);
nor I_686 (I13134,I12736,I13069);
DFFARX1 I_687 (I13134,I1451,I12710,I12681,);
nor I_688 (I13165,I13013,I13069);
not I_689 (I13182,I13165);
nand I_690 (I12690,I13182,I13038);
not I_691 (I13237,I1458);
DFFARX1 I_692 (I13753,I1451,I13237,I13263,);
not I_693 (I13271,I13263);
nand I_694 (I13288,I13735,I13735);
and I_695 (I13305,I13288,I13741);
DFFARX1 I_696 (I13305,I1451,I13237,I13331,);
DFFARX1 I_697 (I13331,I1451,I13237,I13226,);
DFFARX1 I_698 (I13738,I1451,I13237,I13362,);
nand I_699 (I13370,I13362,I13747);
not I_700 (I13387,I13370);
DFFARX1 I_701 (I13387,I1451,I13237,I13413,);
not I_702 (I13421,I13413);
nor I_703 (I13229,I13271,I13421);
DFFARX1 I_704 (I13759,I1451,I13237,I13461,);
nor I_705 (I13220,I13461,I13331);
nor I_706 (I13211,I13461,I13387);
nand I_707 (I13497,I13750,I13744);
and I_708 (I13514,I13497,I13738);
DFFARX1 I_709 (I13514,I1451,I13237,I13540,);
not I_710 (I13548,I13540);
nand I_711 (I13565,I13548,I13461);
nand I_712 (I13214,I13548,I13370);
nor I_713 (I13596,I13756,I13744);
and I_714 (I13613,I13461,I13596);
nor I_715 (I13630,I13548,I13613);
DFFARX1 I_716 (I13630,I1451,I13237,I13223,);
nor I_717 (I13661,I13263,I13596);
DFFARX1 I_718 (I13661,I1451,I13237,I13208,);
nor I_719 (I13692,I13540,I13596);
not I_720 (I13709,I13692);
nand I_721 (I13217,I13709,I13565);
not I_722 (I13767,I1458);
DFFARX1 I_723 (I6476,I1451,I13767,I13793,);
and I_724 (I13801,I13793,I6491);
DFFARX1 I_725 (I13801,I1451,I13767,I13750,);
DFFARX1 I_726 (I6494,I1451,I13767,I13841,);
not I_727 (I13849,I6488);
not I_728 (I13866,I6503);
nand I_729 (I13883,I13866,I13849);
nor I_730 (I13738,I13841,I13883);
DFFARX1 I_731 (I13883,I1451,I13767,I13923,);
not I_732 (I13759,I13923);
not I_733 (I13945,I6479);
nand I_734 (I13962,I13866,I13945);
DFFARX1 I_735 (I13962,I1451,I13767,I13988,);
not I_736 (I13996,I13988);
not I_737 (I14013,I6482);
nand I_738 (I14030,I14013,I6476);
and I_739 (I14047,I13849,I14030);
nor I_740 (I14064,I13962,I14047);
DFFARX1 I_741 (I14064,I1451,I13767,I13735,);
DFFARX1 I_742 (I14047,I1451,I13767,I13756,);
nor I_743 (I14109,I6482,I6485);
nor I_744 (I13747,I13962,I14109);
or I_745 (I14140,I6482,I6485);
nor I_746 (I14157,I6500,I6497);
DFFARX1 I_747 (I14157,I1451,I13767,I14183,);
not I_748 (I14191,I14183);
nor I_749 (I13753,I14191,I13996);
nand I_750 (I14222,I14191,I13841);
not I_751 (I14239,I6500);
nand I_752 (I14256,I14239,I13945);
nand I_753 (I14273,I14191,I14256);
nand I_754 (I13744,I14273,I14222);
nand I_755 (I13741,I14256,I14140);
not I_756 (I14345,I1458);
DFFARX1 I_757 (I13211,I1451,I14345,I14371,);
and I_758 (I14379,I14371,I13217);
DFFARX1 I_759 (I14379,I1451,I14345,I14328,);
DFFARX1 I_760 (I13223,I1451,I14345,I14419,);
not I_761 (I14427,I13208);
not I_762 (I14444,I13208);
nand I_763 (I14461,I14444,I14427);
nor I_764 (I14316,I14419,I14461);
DFFARX1 I_765 (I14461,I1451,I14345,I14501,);
not I_766 (I14337,I14501);
not I_767 (I14523,I13226);
nand I_768 (I14540,I14444,I14523);
DFFARX1 I_769 (I14540,I1451,I14345,I14566,);
not I_770 (I14574,I14566);
not I_771 (I14591,I13220);
nand I_772 (I14608,I14591,I13211);
and I_773 (I14625,I14427,I14608);
nor I_774 (I14642,I14540,I14625);
DFFARX1 I_775 (I14642,I1451,I14345,I14313,);
DFFARX1 I_776 (I14625,I1451,I14345,I14334,);
nor I_777 (I14687,I13220,I13229);
nor I_778 (I14325,I14540,I14687);
or I_779 (I14718,I13220,I13229);
nor I_780 (I14735,I13214,I13214);
DFFARX1 I_781 (I14735,I1451,I14345,I14761,);
not I_782 (I14769,I14761);
nor I_783 (I14331,I14769,I14574);
nand I_784 (I14800,I14769,I14419);
not I_785 (I14817,I13214);
nand I_786 (I14834,I14817,I14523);
nand I_787 (I14851,I14769,I14834);
nand I_788 (I14322,I14851,I14800);
nand I_789 (I14319,I14834,I14718);
not I_790 (I14923,I1458);
DFFARX1 I_791 (I12684,I1451,I14923,I14949,);
and I_792 (I14957,I14949,I12690);
DFFARX1 I_793 (I14957,I1451,I14923,I14906,);
DFFARX1 I_794 (I12696,I1451,I14923,I14997,);
not I_795 (I15005,I12681);
not I_796 (I15022,I12681);
nand I_797 (I15039,I15022,I15005);
nor I_798 (I14894,I14997,I15039);
DFFARX1 I_799 (I15039,I1451,I14923,I15079,);
not I_800 (I14915,I15079);
not I_801 (I15101,I12699);
nand I_802 (I15118,I15022,I15101);
DFFARX1 I_803 (I15118,I1451,I14923,I15144,);
not I_804 (I15152,I15144);
not I_805 (I15169,I12693);
nand I_806 (I15186,I15169,I12684);
and I_807 (I15203,I15005,I15186);
nor I_808 (I15220,I15118,I15203);
DFFARX1 I_809 (I15220,I1451,I14923,I14891,);
DFFARX1 I_810 (I15203,I1451,I14923,I14912,);
nor I_811 (I15265,I12693,I12702);
nor I_812 (I14903,I15118,I15265);
or I_813 (I15296,I12693,I12702);
nor I_814 (I15313,I12687,I12687);
DFFARX1 I_815 (I15313,I1451,I14923,I15339,);
not I_816 (I15347,I15339);
nor I_817 (I14909,I15347,I15152);
nand I_818 (I15378,I15347,I14997);
not I_819 (I15395,I12687);
nand I_820 (I15412,I15395,I15101);
nand I_821 (I15429,I15347,I15412);
nand I_822 (I14900,I15429,I15378);
nand I_823 (I14897,I15412,I15296);
not I_824 (I15501,I1458);
DFFARX1 I_825 (I16612,I1451,I15501,I15527,);
and I_826 (I15535,I15527,I16606);
DFFARX1 I_827 (I15535,I1451,I15501,I15484,);
DFFARX1 I_828 (I16591,I1451,I15501,I15575,);
not I_829 (I15583,I16597);
not I_830 (I15600,I16609);
nand I_831 (I15617,I15600,I15583);
nor I_832 (I15472,I15575,I15617);
DFFARX1 I_833 (I15617,I1451,I15501,I15657,);
not I_834 (I15493,I15657);
not I_835 (I15679,I16591);
nand I_836 (I15696,I15600,I15679);
DFFARX1 I_837 (I15696,I1451,I15501,I15722,);
not I_838 (I15730,I15722);
not I_839 (I15747,I16615);
nand I_840 (I15764,I15747,I16603);
and I_841 (I15781,I15583,I15764);
nor I_842 (I15798,I15696,I15781);
DFFARX1 I_843 (I15798,I1451,I15501,I15469,);
DFFARX1 I_844 (I15781,I1451,I15501,I15490,);
nor I_845 (I15843,I16615,I16594);
nor I_846 (I15481,I15696,I15843);
or I_847 (I15874,I16615,I16594);
nor I_848 (I15891,I16600,I16594);
DFFARX1 I_849 (I15891,I1451,I15501,I15917,);
not I_850 (I15925,I15917);
nor I_851 (I15487,I15925,I15730);
nand I_852 (I15956,I15925,I15575);
not I_853 (I15973,I16600);
nand I_854 (I15990,I15973,I15679);
nand I_855 (I16007,I15925,I15990);
nand I_856 (I15478,I16007,I15956);
nand I_857 (I15475,I15990,I15874);
not I_858 (I16079,I1458);
DFFARX1 I_859 (I10423,I1451,I16079,I16105,);
nand I_860 (I16113,I16105,I10438);
DFFARX1 I_861 (I10432,I1451,I16079,I16139,);
DFFARX1 I_862 (I16139,I1451,I16079,I16156,);
not I_863 (I16071,I16156);
not I_864 (I16178,I10435);
nor I_865 (I16195,I10435,I10441);
not I_866 (I16212,I10423);
nand I_867 (I16229,I16178,I16212);
nor I_868 (I16246,I10423,I10435);
and I_869 (I16050,I16246,I16113);
not I_870 (I16277,I10420);
nand I_871 (I16294,I16277,I10426);
nor I_872 (I16311,I10420,I10420);
not I_873 (I16328,I16311);
nand I_874 (I16053,I16195,I16328);
DFFARX1 I_875 (I16311,I1451,I16079,I16068,);
nor I_876 (I16373,I10429,I10423);
nor I_877 (I16390,I16373,I10441);
and I_878 (I16407,I16390,I16294);
DFFARX1 I_879 (I16407,I1451,I16079,I16065,);
nor I_880 (I16062,I16373,I16229);
or I_881 (I16059,I16311,I16373);
nor I_882 (I16466,I10429,I10444);
DFFARX1 I_883 (I16466,I1451,I16079,I16492,);
not I_884 (I16500,I16492);
nand I_885 (I16517,I16500,I16178);
nor I_886 (I16534,I16517,I10441);
DFFARX1 I_887 (I16534,I1451,I16079,I16047,);
nor I_888 (I16565,I16500,I16229);
nor I_889 (I16056,I16373,I16565);
not I_890 (I16623,I1458);
DFFARX1 I_891 (I8689,I1451,I16623,I16649,);
nand I_892 (I16657,I16649,I8704);
DFFARX1 I_893 (I8698,I1451,I16623,I16683,);
DFFARX1 I_894 (I16683,I1451,I16623,I16700,);
not I_895 (I16615,I16700);
not I_896 (I16722,I8701);
nor I_897 (I16739,I8701,I8707);
not I_898 (I16756,I8689);
nand I_899 (I16773,I16722,I16756);
nor I_900 (I16790,I8689,I8701);
and I_901 (I16594,I16790,I16657);
not I_902 (I16821,I8686);
nand I_903 (I16838,I16821,I8692);
nor I_904 (I16855,I8686,I8686);
not I_905 (I16872,I16855);
nand I_906 (I16597,I16739,I16872);
DFFARX1 I_907 (I16855,I1451,I16623,I16612,);
nor I_908 (I16917,I8695,I8689);
nor I_909 (I16934,I16917,I8707);
and I_910 (I16951,I16934,I16838);
DFFARX1 I_911 (I16951,I1451,I16623,I16609,);
nor I_912 (I16606,I16917,I16773);
or I_913 (I16603,I16855,I16917);
nor I_914 (I17010,I8695,I8710);
DFFARX1 I_915 (I17010,I1451,I16623,I17036,);
not I_916 (I17044,I17036);
nand I_917 (I17061,I17044,I16722);
nor I_918 (I17078,I17061,I8707);
DFFARX1 I_919 (I17078,I1451,I16623,I16591,);
nor I_920 (I17109,I17044,I16773);
nor I_921 (I16600,I16917,I17109);
not I_922 (I17167,I1458);
DFFARX1 I_923 (I5955,I1451,I17167,I17193,);
nand I_924 (I17201,I17193,I5976);
not I_925 (I17218,I17201);
DFFARX1 I_926 (I5970,I1451,I17167,I17244,);
not I_927 (I17252,I17244);
not I_928 (I17269,I5958);
or I_929 (I17286,I5973,I5958);
nor I_930 (I17303,I5973,I5958);
or I_931 (I17320,I5964,I5973);
DFFARX1 I_932 (I17320,I1451,I17167,I17159,);
not I_933 (I17351,I5952);
nand I_934 (I17368,I17351,I5949);
nand I_935 (I17385,I17269,I17368);
and I_936 (I17138,I17252,I17385);
nor I_937 (I17416,I5952,I5961);
and I_938 (I17433,I17252,I17416);
nor I_939 (I17144,I17218,I17433);
DFFARX1 I_940 (I17416,I1451,I17167,I17473,);
not I_941 (I17481,I17473);
nor I_942 (I17153,I17252,I17481);
or I_943 (I17512,I17320,I5967);
nor I_944 (I17529,I5967,I5964);
nand I_945 (I17546,I17385,I17529);
nand I_946 (I17563,I17512,I17546);
DFFARX1 I_947 (I17563,I1451,I17167,I17156,);
nor I_948 (I17594,I17529,I17286);
DFFARX1 I_949 (I17594,I1451,I17167,I17135,);
nor I_950 (I17625,I5967,I5949);
DFFARX1 I_951 (I17625,I1451,I17167,I17651,);
DFFARX1 I_952 (I17651,I1451,I17167,I17150,);
not I_953 (I17673,I17651);
nand I_954 (I17147,I17673,I17201);
nand I_955 (I17141,I17673,I17303);
endmodule


