module test_I17174(I1477,I14954,I15310,I17013,I15228,I14930,I1470,I15502,I17174);
input I1477,I14954,I15310,I17013,I15228,I14930,I1470,I15502;
output I17174;
wire I14948,I14965,I17157,I17047,I16835,I16852,I17030,I14957,I14933,I17092,I16818,I17109,I14936,I16869;
DFFARX1 I_0(I1470,I14965,,,I14948,);
not I_1(I14965,I1477);
nand I_2(I17157,I17109,I17047);
DFFARX1 I_3(I17030,I1470,I16818,,,I17047,);
nand I_4(I16835,I14936,I14948);
and I_5(I16852,I16835,I14957);
and I_6(I17030,I17013,I14930);
nand I_7(I14957,I15502,I15228);
DFFARX1 I_8(I15310,I1470,I14965,,,I14933,);
DFFARX1 I_9(I14954,I1470,I16818,,,I17092,);
not I_10(I16818,I1477);
and I_11(I17109,I17092,I14933);
DFFARX1 I_12(I1470,I14965,,,I14936,);
and I_13(I17174,I16869,I17157);
DFFARX1 I_14(I16852,I1470,I16818,,,I16869,);
endmodule


