module test_I9453(I1477,I1470,I9655,I8208,I9453);
input I1477,I1470,I9655,I8208;
output I9453;
wire I8216,I9672,I9720,I8623,I9816,I8705,I9689,I8193,I9491;
not I_0(I8216,I1477);
and I_1(I9672,I9655,I8208);
not I_2(I9720,I9689);
DFFARX1 I_3(I1470,I8216,,,I8623,);
DFFARX1 I_4(I8193,I1470,I9491,,,I9816,);
DFFARX1 I_5(I8623,I1470,I8216,,,I8705,);
nand I_6(I9453,I9816,I9720);
DFFARX1 I_7(I9672,I1470,I9491,,,I9689,);
not I_8(I8193,I8705);
not I_9(I9491,I1477);
endmodule


