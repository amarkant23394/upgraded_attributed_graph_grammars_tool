module test_I16968(I1477,I15126,I14999,I1470,I15502,I16968);
input I1477,I15126,I14999,I1470,I15502;
output I16968;
wire I15245,I14948,I14951,I14965,I12581,I15423,I14945,I16818,I15211,I15016,I16934,I16951,I15519,I15372,I16886;
nor I_0(I15245,I15211,I15126);
DFFARX1 I_1(I15519,I1470,I14965,,,I14948,);
nand I_2(I14951,I15016,I15245);
not I_3(I14965,I1477);
DFFARX1 I_4(I1470,,,I12581,);
and I_5(I15423,I15372);
nand I_6(I14945,I15372,I15126);
nor I_7(I16968,I16886,I16951);
not I_8(I16818,I1477);
DFFARX1 I_9(I1470,I14965,,,I15211,);
nand I_10(I15016,I14999,I12581);
DFFARX1 I_11(I14945,I1470,I16818,,,I16934,);
not I_12(I16951,I16934);
or I_13(I15519,I15502,I15423);
DFFARX1 I_14(I1470,I14965,,,I15372,);
nor I_15(I16886,I14951,I14948);
endmodule


