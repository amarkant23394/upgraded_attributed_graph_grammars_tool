module test_I1495(I1477,I1295,I1470,I1535,I1207,I1620,I1495);
input I1477,I1295,I1470,I1535,I1207,I1620;
output I1495;
wire I1518,I1784,I2038,I2021,I2103,I1832,I1849,I1767;
not I_0(I1518,I1477);
nor I_1(I1784,I1767,I1620);
not I_2(I2038,I2021);
DFFARX1 I_3(I1295,I1470,I1518,,,I2021,);
DFFARX1 I_4(I2103,I1470,I1518,,,I1495,);
or I_5(I2103,I2038,I1849);
nand I_6(I1832,I1535,I1207);
and I_7(I1849,I1832,I1784);
DFFARX1 I_8(I1470,I1518,,,I1767,);
endmodule


