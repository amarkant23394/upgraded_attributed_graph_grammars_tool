module test_I6510(I2742,I4017,I1477,I1470,I6510);
input I2742,I4017,I1477,I1470;
output I6510;
wire I3966,I6329,I6493,I4068,I4034,I2724,I3983;
not I_0(I6510,I6493);
or I_1(I3966,I4068,I4034);
not I_2(I6329,I1477);
DFFARX1 I_3(I3966,I1470,I6329,,,I6493,);
nor I_4(I4068,I2742,I2724);
DFFARX1 I_5(I4017,I1470,I3983,,,I4034,);
DFFARX1 I_6(I1470,,,I2724,);
not I_7(I3983,I1477);
endmodule


