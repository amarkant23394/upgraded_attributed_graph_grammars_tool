module test_I10490(I6476,I7799,I1477,I1470,I6294,I10490);
input I6476,I7799,I1477,I1470,I6294;
output I10490;
wire I6781,I7556,I6297,I7621,I7816,I7570,I7714,I7850,I7604,I7731,I10052,I6315;
DFFARX1 I_0(I1470,,,I6781,);
nand I_1(I7556,I7621,I7850);
DFFARX1 I_2(I1470,,,I6297,);
nand I_3(I7621,I7604,I6315);
DFFARX1 I_4(I7799,I1470,I7570,,,I7816,);
not I_5(I7570,I1477);
not I_6(I7714,I6297);
nor I_7(I7850,I7816,I7731);
nor I_8(I7604,I6297,I6294);
not I_9(I7731,I7714);
DFFARX1 I_10(I7556,I1470,I10052,,,I10490,);
not I_11(I10052,I1477);
nand I_12(I6315,I6781,I6476);
endmodule


