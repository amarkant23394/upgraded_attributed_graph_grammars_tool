module test_final(G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_3,blif_reset_net_1_r_3,G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3);
input G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_3,blif_reset_net_1_r_3;
output G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3;
wire G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16,n4_1_l_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16,n4_1_l_3,n9_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3;
DFFARX1 I_0(n4_1_r_16,blif_clk_net_1_r_3,n9_3,G42_1_r_16,);
nor I_1(n_572_1_r_16,n20_16,n21_16);
nand I_2(n_573_1_r_16,n18_16,n19_16);
nor I_3(n_549_1_r_16,n23_16,n24_16);
nand I_4(n_569_1_r_16,n18_16,n22_16);
nor I_5(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_6(N1_4_r_16,blif_clk_net_1_r_3,n9_3,G199_4_r_16,);
DFFARX1 I_7(n6_16,blif_clk_net_1_r_3,n9_3,G214_4_r_16,);
DFFARX1 I_8(n_573_1_l_16,blif_clk_net_1_r_3,n9_3,ACVQN1_5_r_16,);
not I_9(P6_5_r_16,P6_5_r_internal_16);
nor I_10(n4_1_l_16,G18_1_l_16,IN_1_1_l_16);
DFFARX1 I_11(n4_1_l_16,blif_clk_net_1_r_3,n9_3,n29_16,);
DFFARX1 I_12(IN_1_3_l_16,blif_clk_net_1_r_3,n9_3,n16_internal_16,);
not I_13(n16_16,n16_internal_16);
DFFARX1 I_14(IN_2_3_l_16,blif_clk_net_1_r_3,n9_3,ACVQN1_3_l_16,);
nor I_15(n4_1_r_16,n29_16,n21_16);
nor I_16(N1_4_r_16,n27_16,n28_16);
not I_17(n6_16,n19_16);
or I_18(n_573_1_l_16,IN_5_1_l_16,IN_9_1_l_16);
nor I_19(n_452_1_l_16,G18_1_l_16,IN_5_1_l_16);
DFFARX1 I_20(n_452_1_l_16,blif_clk_net_1_r_3,n9_3,P6_5_r_internal_16,);
not I_21(n18_16,n20_16);
nor I_22(n19_16,IN_9_1_l_16,IN_10_1_l_16);
nor I_23(n20_16,G15_1_l_16,IN_7_1_l_16);
nor I_24(n21_16,IN_10_1_l_16,n25_16);
nand I_25(n22_16,IN_4_3_l_16,ACVQN1_3_l_16);
not I_26(n23_16,n22_16);
nor I_27(n24_16,n16_16,n20_16);
nor I_28(n25_16,G15_1_l_16,n26_16);
not I_29(n26_16,IN_4_1_l_16);
and I_30(n27_16,IN_9_1_l_16,n29_16);
not I_31(n28_16,n_452_1_l_16);
DFFARX1 I_32(n4_1_r_3,blif_clk_net_1_r_3,n9_3,G42_1_r_3,);
nor I_33(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_34(n_573_1_r_3,n26_3,n27_3);
nor I_35(n_549_1_r_3,n40_3,n32_3);
nand I_36(n_569_1_r_3,n27_3,n31_3);
and I_37(n_452_1_r_3,n26_3,n_549_1_r_16);
nor I_38(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_39(N3_2_r_3,blif_clk_net_1_r_3,n9_3,G199_2_r_3,);
DFFARX1 I_40(n_572_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_3,);
nor I_41(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_42(n4_1_l_3,n_549_1_r_16,G199_4_r_16);
not I_43(n9_3,blif_reset_net_1_r_3);
DFFARX1 I_44(n4_1_l_3,blif_clk_net_1_r_3,n9_3,G42_1_l_3,);
not I_45(n22_3,G42_1_l_3);
DFFARX1 I_46(n_572_1_r_16,blif_clk_net_1_r_3,n9_3,n40_3,);
DFFARX1 I_47(ACVQN1_5_r_16,blif_clk_net_1_r_3,n9_3,n25_internal_3,);
not I_48(n25_3,n25_internal_3);
nor I_49(n4_1_r_3,n40_3,n36_3);
nor I_50(N3_2_r_3,n26_3,n37_3);
nor I_51(n_572_1_l_3,G42_1_r_16,P6_5_r_16);
DFFARX1 I_52(G42_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN1_3_r_3,);
nor I_53(n26_3,n_573_1_r_16,G42_1_r_16);
not I_54(n27_3,G214_4_r_16);
nor I_55(n28_3,n29_3,G214_4_r_16);
nor I_56(n29_3,n30_3,P6_5_r_16);
not I_57(n30_3,n_569_1_r_16);
nor I_58(n31_3,n40_3,n_573_1_r_16);
nor I_59(n32_3,n25_3,n33_3);
nand I_60(n33_3,n22_3,n_452_1_r_16);
or I_61(n34_3,n_573_1_r_16,G214_4_r_16);
nand I_62(n35_3,ACVQN1_3_r_3,n_452_1_r_16);
nor I_63(n36_3,n_549_1_r_16,G42_1_r_16);
nor I_64(n37_3,n38_3,n39_3);
not I_65(n38_3,n_572_1_l_3);
nand I_66(n39_3,n27_3,n30_3);
endmodule


