module test_final(IN_1_0_l_9,IN_2_0_l_9,IN_4_0_l_9,G18_4_l_9,G15_4_l_9,IN_1_4_l_9,IN_4_4_l_9,IN_5_4_l_9,IN_7_4_l_9,IN_9_4_l_9,IN_10_4_l_9,blif_clk_net_3_r_10,blif_reset_net_3_r_10,n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10);
input IN_1_0_l_9,IN_2_0_l_9,IN_4_0_l_9,G18_4_l_9,G15_4_l_9,IN_1_4_l_9,IN_4_4_l_9,IN_5_4_l_9,IN_7_4_l_9,IN_9_4_l_9,IN_10_4_l_9,blif_clk_net_3_r_10,blif_reset_net_3_r_10;
output n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10;
wire G199_1_r_9,G214_1_r_9,ACVQN1_2_r_9,P6_2_r_9,n_429_or_0_3_r_9,G78_3_r_9,n_576_3_r_9,n_102_3_r_9,n_547_3_r_9,n_42_5_r_9,G199_5_r_9,ACVQN2_0_l_9,n_266_and_0_0_l_9,ACVQN1_0_l_9,n4_4_l_9,G42_4_l_9,n_87_4_l_9,n_572_4_l_9,n_573_4_l_9,n_549_4_l_9,n7_4_l_9,n_569_4_l_9,n_452_4_l_9,N1_1_r_9,n3_1_r_9,P6_internal_2_r_9,n12_3_r_9,n_431_3_r_9,n11_3_r_9,n13_3_r_9,n14_3_r_9,n15_3_r_9,n16_3_r_9,N3_5_r_9,n3_5_r_9,n2_3_r_10,ACVQN2_0_l_10,n_266_and_0_0_l_10,ACVQN1_0_l_10,n4_4_l_10,G42_4_l_10,n_87_4_l_10,n_572_4_l_10,n_573_4_l_10,n_549_4_l_10,n7_4_l_10,n_569_4_l_10,n_452_4_l_10,n12_3_r_10,n_431_3_r_10,n11_3_r_10,n13_3_r_10,n14_3_r_10,n15_3_r_10,n16_3_r_10,n4_4_r_10,n_87_4_r_10,n7_4_r_10;
DFFARX1 I_0(N1_1_r_9,blif_clk_net_3_r_10,n2_3_r_10,G199_1_r_9,);
DFFARX1 I_1(G42_4_l_9,blif_clk_net_3_r_10,n2_3_r_10,G214_1_r_9,);
DFFARX1 I_2(n_572_4_l_9,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_2_r_9,);
not I_3(P6_2_r_9,P6_internal_2_r_9);
nand I_4(n_429_or_0_3_r_9,n_572_4_l_9,n12_3_r_9);
DFFARX1 I_5(n_431_3_r_9,blif_clk_net_3_r_10,n2_3_r_10,G78_3_r_9,);
nand I_6(n_576_3_r_9,n_573_4_l_9,n11_3_r_9);
not I_7(n_102_3_r_9,n_266_and_0_0_l_9);
nand I_8(n_547_3_r_9,n_549_4_l_9,n13_3_r_9);
nor I_9(n_42_5_r_9,n_569_4_l_9,n_452_4_l_9);
DFFARX1 I_10(N3_5_r_9,blif_clk_net_3_r_10,n2_3_r_10,G199_5_r_9,);
DFFARX1 I_11(IN_1_0_l_9,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_l_9,);
and I_12(n_266_and_0_0_l_9,IN_4_0_l_9,ACVQN1_0_l_9);
DFFARX1 I_13(IN_2_0_l_9,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_l_9,);
nor I_14(n4_4_l_9,G18_4_l_9,IN_1_4_l_9);
DFFARX1 I_15(n4_4_l_9,blif_clk_net_3_r_10,n2_3_r_10,G42_4_l_9,);
not I_16(n_87_4_l_9,G15_4_l_9);
nor I_17(n_572_4_l_9,G15_4_l_9,IN_7_4_l_9);
or I_18(n_573_4_l_9,IN_5_4_l_9,IN_9_4_l_9);
nor I_19(n_549_4_l_9,IN_10_4_l_9,n7_4_l_9);
and I_20(n7_4_l_9,IN_4_4_l_9,n_87_4_l_9);
or I_21(n_569_4_l_9,IN_9_4_l_9,IN_10_4_l_9);
nor I_22(n_452_4_l_9,G18_4_l_9,IN_5_4_l_9);
and I_23(N1_1_r_9,n_266_and_0_0_l_9,n3_1_r_9);
nand I_24(n3_1_r_9,n_572_4_l_9,n_569_4_l_9);
DFFARX1 I_25(n_266_and_0_0_l_9,blif_clk_net_3_r_10,n2_3_r_10,P6_internal_2_r_9,);
not I_26(n12_3_r_9,G42_4_l_9);
or I_27(n_431_3_r_9,n_549_4_l_9,n14_3_r_9);
nor I_28(n11_3_r_9,ACVQN2_0_l_9,n12_3_r_9);
nor I_29(n13_3_r_9,ACVQN2_0_l_9,n_266_and_0_0_l_9);
and I_30(n14_3_r_9,n_452_4_l_9,n15_3_r_9);
nor I_31(n15_3_r_9,G42_4_l_9,n16_3_r_9);
not I_32(n16_3_r_9,n_572_4_l_9);
and I_33(N3_5_r_9,ACVQN2_0_l_9,n3_5_r_9);
nand I_34(n3_5_r_9,n_573_4_l_9,n_452_4_l_9);
nand I_35(n_429_or_0_3_r_10,n_266_and_0_0_l_10,n12_3_r_10);
DFFARX1 I_36(n_431_3_r_10,blif_clk_net_3_r_10,n2_3_r_10,G78_3_r_10,);
nand I_37(n_576_3_r_10,ACVQN2_0_l_10,n11_3_r_10);
not I_38(n_102_3_r_10,G42_4_l_10);
nand I_39(n_547_3_r_10,n_569_4_l_10,n13_3_r_10);
DFFARX1 I_40(n4_4_r_10,blif_clk_net_3_r_10,n2_3_r_10,G42_4_r_10,);
nor I_41(n_572_4_r_10,ACVQN2_0_l_10,n_573_4_l_10);
or I_42(n_573_4_r_10,n_569_4_l_10,n_452_4_l_10);
nor I_43(n_549_4_r_10,n_572_4_l_10,n7_4_r_10);
or I_44(n_569_4_r_10,n_572_4_l_10,n_569_4_l_10);
nor I_45(n_452_4_r_10,n_266_and_0_0_l_10,n_452_4_l_10);
not I_46(n2_3_r_10,blif_reset_net_3_r_10);
DFFARX1 I_47(ACVQN1_2_r_9,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_l_10,);
and I_48(n_266_and_0_0_l_10,ACVQN1_0_l_10,n_547_3_r_9);
DFFARX1 I_49(n_576_3_r_9,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_l_10,);
nor I_50(n4_4_l_10,G78_3_r_9,n_42_5_r_9);
DFFARX1 I_51(n4_4_l_10,blif_clk_net_3_r_10,n2_3_r_10,G42_4_l_10,);
not I_52(n_87_4_l_10,G214_1_r_9);
nor I_53(n_572_4_l_10,G214_1_r_9,G199_5_r_9);
or I_54(n_573_4_l_10,G199_1_r_9,n_102_3_r_9);
nor I_55(n_549_4_l_10,n7_4_l_10,P6_2_r_9);
and I_56(n7_4_l_10,n_87_4_l_10,n_429_or_0_3_r_9);
or I_57(n_569_4_l_10,P6_2_r_9,n_102_3_r_9);
nor I_58(n_452_4_l_10,G199_1_r_9,G78_3_r_9);
not I_59(n12_3_r_10,n_549_4_l_10);
or I_60(n_431_3_r_10,n_572_4_l_10,n14_3_r_10);
nor I_61(n11_3_r_10,G42_4_l_10,n12_3_r_10);
nor I_62(n13_3_r_10,G42_4_l_10,n_549_4_l_10);
and I_63(n14_3_r_10,ACVQN2_0_l_10,n15_3_r_10);
nor I_64(n15_3_r_10,n_573_4_l_10,n16_3_r_10);
not I_65(n16_3_r_10,n_266_and_0_0_l_10);
nor I_66(n4_4_r_10,n_266_and_0_0_l_10,G42_4_l_10);
not I_67(n_87_4_r_10,ACVQN2_0_l_10);
and I_68(n7_4_r_10,n_452_4_l_10,n_87_4_r_10);
endmodule


