module test_I15597(I11938,I1470,I13775,I13843,I15597);
input I11938,I1470,I13775,I13843;
output I15597;
wire I13908,I13761,I15696,I13743,I15832,I16145,I14162,I15628,I15679,I13749,I13891,I16052,I13758,I16162,I16069;
not I_0(I13908,I13891);
nand I_1(I13761,I13891);
nor I_2(I15597,I15832,I16162);
nand I_3(I15696,I15679,I13758);
DFFARX1 I_4(I13891,I1470,I13775,,,I13743,);
nand I_5(I15832,I15628,I13749);
not I_6(I16145,I16069);
DFFARX1 I_7(I11938,I1470,I13775,,,I14162,);
not I_8(I15628,I13743);
nor I_9(I15679,I15628,I13761);
nand I_10(I13749,I14162,I13908);
DFFARX1 I_11(I1470,I13775,,,I13891,);
DFFARX1 I_12(I1470,,,I16052,);
not I_13(I13758,I13843);
and I_14(I16162,I15696,I16145);
not I_15(I16069,I16052);
endmodule


