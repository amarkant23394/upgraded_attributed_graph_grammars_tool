module test_final(G1_0_l_8,G2_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_5_0_l_8,IN_7_0_l_8,IN_8_0_l_8,IN_10_0_l_8,IN_11_0_l_8,IN_1_5_l_8,IN_2_5_l_8,blif_clk_net_1_r_4,blif_reset_net_1_r_4,G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4);
input G1_0_l_8,G2_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_5_0_l_8,IN_7_0_l_8,IN_8_0_l_8,IN_10_0_l_8,IN_11_0_l_8,IN_1_5_l_8,IN_2_5_l_8,blif_clk_net_1_r_4,blif_reset_net_1_r_4;
output G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4;
wire G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8,n_431_0_l_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n_431_0_l_4,n6_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4;
DFFARX1 I_0(n4_1_r_8,blif_clk_net_1_r_4,n6_4,G42_1_r_8,);
nor I_1(n_572_1_r_8,n39_8,n23_8);
and I_2(n_549_1_r_8,n38_8,n23_8);
nand I_3(n_569_1_r_8,n38_8,n24_8);
nor I_4(n_452_1_r_8,n25_8,n26_8);
nor I_5(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_6(N3_2_r_8,blif_clk_net_1_r_4,n6_4,G199_2_r_8,);
DFFARX1 I_7(N1_4_r_8,blif_clk_net_1_r_4,n6_4,G199_4_r_8,);
DFFARX1 I_8(G78_0_l_8,blif_clk_net_1_r_4,n6_4,G214_4_r_8,);
or I_9(n_431_0_l_8,IN_8_0_l_8,n29_8);
DFFARX1 I_10(n_431_0_l_8,blif_clk_net_1_r_4,n6_4,G78_0_l_8,);
not I_11(n19_8,G78_0_l_8);
DFFARX1 I_12(IN_2_5_l_8,blif_clk_net_1_r_4,n6_4,n39_8,);
not I_13(n22_8,n39_8);
DFFARX1 I_14(IN_1_5_l_8,blif_clk_net_1_r_4,n6_4,n38_8,);
nor I_15(n4_1_r_8,G78_0_l_8,n33_8);
nor I_16(N3_2_r_8,n22_8,n35_8);
nor I_17(N1_4_r_8,n27_8,n37_8);
nand I_18(n23_8,IN_7_0_l_8,n32_8);
not I_19(n24_8,n23_8);
nand I_20(n25_8,IN_11_0_l_8,n36_8);
nand I_21(n26_8,n27_8,n28_8);
nor I_22(n27_8,IN_5_0_l_8,n31_8);
not I_23(n28_8,G2_0_l_8);
and I_24(n29_8,IN_2_0_l_8,n30_8);
nor I_25(n30_8,IN_4_0_l_8,n31_8);
not I_26(n31_8,G1_0_l_8);
and I_27(n32_8,IN_5_0_l_8,n28_8);
nand I_28(n33_8,n28_8,n34_8);
not I_29(n34_8,n25_8);
nor I_30(n35_8,G2_0_l_8,n34_8);
not I_31(n36_8,IN_10_0_l_8);
nor I_32(n37_8,n19_8,n38_8);
DFFARX1 I_33(n4_1_r_4,blif_clk_net_1_r_4,n6_4,G42_1_r_4,);
nor I_34(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_35(n_573_1_r_4,n16_4,n_572_1_r_8);
nor I_36(n_549_1_r_4,n22_4,n23_4);
nand I_37(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_38(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_4,);
nor I_39(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_40(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_4,);
not I_41(P6_5_r_4,P6_5_r_internal_4);
or I_42(n_431_0_l_4,n26_4,n_42_2_r_8);
not I_43(n6_4,blif_reset_net_1_r_4);
DFFARX1 I_44(n_431_0_l_4,blif_clk_net_1_r_4,n6_4,G78_0_l_4,);
DFFARX1 I_45(G199_2_r_8,blif_clk_net_1_r_4,n6_4,ACVQN1_5_l_4,);
not I_46(n16_4,ACVQN1_5_l_4);
DFFARX1 I_47(G42_1_r_8,blif_clk_net_1_r_4,n6_4,n17_internal_4,);
not I_48(n17_4,n17_internal_4);
nor I_49(n4_1_r_4,n30_4,n31_4);
nand I_50(n19_4,n33_4,n_452_1_r_8);
DFFARX1 I_51(G78_0_l_4,blif_clk_net_1_r_4,n6_4,n15_internal_4,);
not I_52(n15_4,n15_internal_4);
DFFARX1 I_53(ACVQN1_5_l_4,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_4,);
and I_54(n20_4,n16_4,G199_4_r_8);
nor I_55(n21_4,n_569_1_r_8,n_572_1_r_8);
nand I_56(n22_4,G78_0_l_4,n25_4);
nand I_57(n23_4,n24_4,G199_4_r_8);
not I_58(n24_4,n_572_1_r_8);
not I_59(n25_4,n_569_1_r_8);
and I_60(n26_4,n27_4,G214_4_r_8);
nor I_61(n27_4,n28_4,n_549_1_r_8);
not I_62(n28_4,n_452_1_r_8);
not I_63(n29_4,n30_4);
nand I_64(n30_4,n32_4,G42_1_r_8);
nand I_65(n31_4,n25_4,G199_4_r_8);
nor I_66(n32_4,n33_4,n_572_1_r_8);
not I_67(n33_4,n_572_1_r_8);
endmodule


