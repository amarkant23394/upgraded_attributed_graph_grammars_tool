module test_I3983_rst(I1477_rst,I3983_rst);
,I3983_rst);
input I1477_rst;
output I3983_rst;
wire ;
not I_0(I3983_rst,I1477_rst);
endmodule


