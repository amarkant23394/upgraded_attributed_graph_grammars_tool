module test_I11281(I1477,I11525,I8833,I1470,I11281);
input I1477,I11525,I8833,I1470;
output I11281;
wire I11542,I11593,I11559,I11310;
or I_0(I11542,I11525,I8833);
not I_1(I11281,I11593);
DFFARX1 I_2(I11559,I1470,I11310,,,I11593,);
DFFARX1 I_3(I11542,I1470,I11310,,,I11559,);
not I_4(I11310,I1477);
endmodule


