module test_I17792(I1477,I13749,I15579,I15696,I15628,I1470,I15798,I17792);
input I1477,I13749,I15579,I15696,I15628,I1470,I15798;
output I17792;
wire I17413,I15585,I15600,I15832,I15815,I16052,I15611,I15959,I17498,I15928,I15597,I17775,I16162,I16069,I17430,I17481;
not I_0(I17413,I1477);
nand I_1(I15585,I16069,I15959);
nor I_2(I17792,I17775,I17498);
or I_3(I15600,I15832,I15815);
nand I_4(I15832,I15628,I13749);
DFFARX1 I_5(I15798,I1470,I15611,,,I15815,);
DFFARX1 I_6(I1470,I15611,,,I16052,);
not I_7(I15611,I1477);
nor I_8(I15959,I15928,I15696);
nand I_9(I17498,I17481,I15600);
DFFARX1 I_10(I1470,I15611,,,I15928,);
nor I_11(I15597,I15832,I16162);
DFFARX1 I_12(I15585,I1470,I17413,,,I17775,);
and I_13(I16162,I15696);
not I_14(I16069,I16052);
not I_15(I17430,I15579);
nor I_16(I17481,I17430,I15597);
endmodule


