module test_I10017(I1477,I7604,I7731,I1470,I6315,I10017);
input I1477,I7604,I7731,I1470,I6315;
output I10017;
wire I7556,I7621,I7816,I10583,I7850,I10052,I10490;
nand I_0(I7556,I7621,I7850);
nand I_1(I7621,I7604,I6315);
DFFARX1 I_2(I1470,,,I7816,);
DFFARX1 I_3(I10490,I1470,I10052,,,I10583,);
nor I_4(I7850,I7816,I7731);
not I_5(I10052,I1477);
DFFARX1 I_6(I7556,I1470,I10052,,,I10490,);
and I_7(I10017,I10490,I10583);
endmodule


