module test_I12541(I7550,I1477,I7535,I1470,I12541);
input I7550,I1477,I7535,I1470;
output I12541;
wire I10349,I7538,I12442,I10038,I10041,I12349,I12425,I12524,I11973,I10120,I10332;
and I_0(I10349,I10332,I7550);
nor I_1(I12541,I12349,I12524);
DFFARX1 I_2(I1470,,,I7538,);
not I_3(I12442,I12425);
nand I_4(I10038,I10349);
nor I_5(I10041,I10349,I10120);
DFFARX1 I_6(I10041,I1470,I11973,,,I12349,);
DFFARX1 I_7(I10038,I1470,I11973,,,I12425,);
not I_8(I12524,I12442);
not I_9(I11973,I1477);
nor I_10(I10120,I7538,I7535);
DFFARX1 I_11(I1470,,,I10332,);
endmodule


