module test_I2895(I1415,I2895);
input I1415;
output I2895;
wire ;
not I_0(I2895,I1415);
endmodule


