module test_final(IN_1_1_l_3,IN_2_1_l_3,IN_3_1_l_3,IN_1_8_l_3,IN_2_8_l_3,IN_3_8_l_3,IN_6_8_l_3,IN_1_10_l_3,IN_2_10_l_3,IN_3_10_l_3,IN_4_10_l_3,blif_clk_net_5_r_5,blif_reset_net_5_r_5,N1371_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1508_6_r_5);
input IN_1_1_l_3,IN_2_1_l_3,IN_3_1_l_3,IN_1_8_l_3,IN_2_8_l_3,IN_3_8_l_3,IN_6_8_l_3,IN_1_10_l_3,IN_2_10_l_3,IN_3_10_l_3,IN_4_10_l_3,blif_clk_net_5_r_5,blif_reset_net_5_r_5;
output N1371_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1508_6_r_5;
wire N1371_0_r_3,N1508_0_r_3,N6147_3_r_3,n_429_or_0_5_r_3,G78_5_r_3,n_576_5_r_3,n_102_5_r_3,n_547_5_r_3,N1372_10_r_3,N1508_10_r_3,N3_8_l_3,n39_3,n_431_5_r_3,n22_3,n23_3,n24_3,n25_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,N1508_0_r_5,N1507_6_r_5,n_431_5_r_5,n6_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5;
nor I_0(N1371_0_r_3,n39_3,n37_3);
nor I_1(N1508_0_r_3,n25_3,n37_3);
nor I_2(N6147_3_r_3,N1372_10_r_3,n33_3);
nand I_3(n_429_or_0_5_r_3,N1372_10_r_3,n30_3);
DFFARX1 I_4(n_431_5_r_3,blif_clk_net_5_r_5,n6_5,G78_5_r_3,);
nand I_5(n_576_5_r_3,n22_3,n23_3);
not I_6(n_102_5_r_3,n39_3);
nand I_7(n_547_5_r_3,n26_3,n27_3);
not I_8(N1372_10_r_3,n36_3);
nor I_9(N1508_10_r_3,n35_3,n36_3);
and I_10(N3_8_l_3,IN_6_8_l_3,n34_3);
DFFARX1 I_11(N3_8_l_3,blif_clk_net_5_r_5,n6_5,n39_3,);
nand I_12(n_431_5_r_3,n29_3,n30_3);
nor I_13(n22_3,n24_3,n25_3);
nor I_14(n23_3,IN_3_1_l_3,n39_3);
not I_15(n24_3,n27_3);
nand I_16(n25_3,IN_1_1_l_3,IN_2_1_l_3);
nor I_17(n26_3,n39_3,n28_3);
nor I_18(n27_3,IN_1_8_l_3,IN_3_8_l_3);
not I_19(n28_3,n37_3);
nand I_20(n29_3,N1372_10_r_3,n39_3);
nand I_21(n30_3,n31_3,n32_3);
not I_22(n31_3,n25_3);
not I_23(n32_3,IN_3_1_l_3);
nand I_24(n33_3,n24_3,n25_3);
nand I_25(n34_3,IN_2_8_l_3,IN_3_8_l_3);
nor I_26(n35_3,n27_3,n31_3);
nand I_27(n36_3,n28_3,n38_3);
nand I_28(n37_3,IN_1_10_l_3,IN_2_10_l_3);
or I_29(n38_3,IN_3_10_l_3,IN_4_10_l_3);
nor I_30(N1371_0_r_5,n28_5,n39_5);
not I_31(N1508_0_r_5,n39_5);
nor I_32(N6147_2_r_5,n28_5,n37_5);
nand I_33(n_429_or_0_5_r_5,n30_5,n32_5);
DFFARX1 I_34(n_431_5_r_5,blif_clk_net_5_r_5,n6_5,G78_5_r_5,);
nand I_35(n_576_5_r_5,n26_5,n27_5);
not I_36(n_102_5_r_5,n28_5);
nand I_37(n_547_5_r_5,n31_5,n32_5);
nor I_38(N1507_6_r_5,n30_5,n32_5);
nor I_39(N1508_6_r_5,n39_5,n41_5);
nand I_40(n_431_5_r_5,n34_5,n35_5);
not I_41(n6_5,blif_reset_net_5_r_5);
nor I_42(n26_5,n29_5,n30_5);
nor I_43(n27_5,n28_5,N1508_0_r_3);
nor I_44(n28_5,n29_5,n44_5);
not I_45(n29_5,N1371_0_r_3);
nand I_46(n30_5,N1508_0_r_5,n43_5);
nor I_47(n31_5,n28_5,n33_5);
nor I_48(n32_5,n40_5,n_429_or_0_5_r_3);
nor I_49(n33_5,n29_5,N1508_0_r_3);
or I_50(n34_5,n29_5,N1508_0_r_3);
nand I_51(n35_5,n32_5,n36_5);
not I_52(n36_5,n30_5);
nor I_53(n37_5,N1507_6_r_5,n38_5);
and I_54(n38_5,n39_5,n40_5);
nand I_55(n39_5,N1371_0_r_3,N6147_3_r_3);
nand I_56(n40_5,n_576_5_r_3,n_102_5_r_3);
nand I_57(n41_5,n28_5,n42_5);
or I_58(n42_5,n32_5,n36_5);
or I_59(n43_5,G78_5_r_3,N1508_10_r_3);
nor I_60(n44_5,N1508_0_r_3,n_547_5_r_3);
endmodule


