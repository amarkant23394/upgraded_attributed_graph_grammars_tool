module test_final(G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_3,blif_reset_net_1_r_3,G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3);
input G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_3,blif_reset_net_1_r_3;
output G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3;
wire G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,n_452_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15,n4_1_l_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15,n4_1_l_3,n9_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3;
DFFARX1 I_0(n_452_1_r_15,blif_clk_net_1_r_3,n9_3,G42_1_r_15,);
and I_1(n_572_1_r_15,n17_15,n19_15);
nand I_2(n_573_1_r_15,n15_15,n18_15);
nor I_3(n_549_1_r_15,n21_15,n22_15);
nand I_4(n_569_1_r_15,n15_15,n20_15);
nor I_5(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_6(G42_1_l_15,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_15,);
nor I_7(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_8(N1_4_r_15,blif_clk_net_1_r_3,n9_3,G199_4_r_15,);
DFFARX1 I_9(n_573_1_l_15,blif_clk_net_1_r_3,n9_3,G214_4_r_15,);
nor I_10(n4_1_l_15,G18_1_l_15,IN_1_1_l_15);
DFFARX1 I_11(n4_1_l_15,blif_clk_net_1_r_3,n9_3,G42_1_l_15,);
not I_12(n15_15,G42_1_l_15);
DFFARX1 I_13(IN_1_3_l_15,blif_clk_net_1_r_3,n9_3,n17_internal_15,);
not I_14(n17_15,n17_internal_15);
DFFARX1 I_15(IN_2_3_l_15,blif_clk_net_1_r_3,n9_3,n30_15,);
nor I_16(n_572_1_l_15,G15_1_l_15,IN_7_1_l_15);
DFFARX1 I_17(n_572_1_l_15,blif_clk_net_1_r_3,n9_3,n14_internal_15,);
not I_18(n14_15,n14_internal_15);
nand I_19(N1_4_r_15,n25_15,n26_15);
or I_20(n_573_1_l_15,IN_5_1_l_15,IN_9_1_l_15);
nor I_21(n18_15,IN_9_1_l_15,IN_10_1_l_15);
nand I_22(n19_15,n27_15,n28_15);
nand I_23(n20_15,IN_4_3_l_15,n30_15);
not I_24(n21_15,n20_15);
and I_25(n22_15,n17_15,n_572_1_l_15);
nor I_26(n23_15,G18_1_l_15,IN_5_1_l_15);
or I_27(n24_15,IN_9_1_l_15,IN_10_1_l_15);
or I_28(n25_15,G18_1_l_15,n_573_1_l_15);
nand I_29(n26_15,n19_15,n23_15);
not I_30(n27_15,IN_10_1_l_15);
nand I_31(n28_15,IN_4_1_l_15,n29_15);
not I_32(n29_15,G15_1_l_15);
DFFARX1 I_33(n4_1_r_3,blif_clk_net_1_r_3,n9_3,G42_1_r_3,);
nor I_34(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_35(n_573_1_r_3,n26_3,n27_3);
nor I_36(n_549_1_r_3,n40_3,n32_3);
nand I_37(n_569_1_r_3,n27_3,n31_3);
and I_38(n_452_1_r_3,n26_3,G199_4_r_15);
nor I_39(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_40(N3_2_r_3,blif_clk_net_1_r_3,n9_3,G199_2_r_3,);
DFFARX1 I_41(n_572_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_3,);
nor I_42(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_43(n4_1_l_3,G199_4_r_15,G42_1_r_15);
not I_44(n9_3,blif_reset_net_1_r_3);
DFFARX1 I_45(n4_1_l_3,blif_clk_net_1_r_3,n9_3,G42_1_l_3,);
not I_46(n22_3,G42_1_l_3);
DFFARX1 I_47(G42_1_r_15,blif_clk_net_1_r_3,n9_3,n40_3,);
DFFARX1 I_48(n_572_1_r_15,blif_clk_net_1_r_3,n9_3,n25_internal_3,);
not I_49(n25_3,n25_internal_3);
nor I_50(n4_1_r_3,n40_3,n36_3);
nor I_51(N3_2_r_3,n26_3,n37_3);
nor I_52(n_572_1_l_3,n_549_1_r_15,ACVQN2_3_r_15);
DFFARX1 I_53(G42_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN1_3_r_3,);
nor I_54(n26_3,n_573_1_r_15,n_569_1_r_15);
not I_55(n27_3,n_266_and_0_3_r_15);
nor I_56(n28_3,n29_3,n_266_and_0_3_r_15);
nor I_57(n29_3,n30_3,n_549_1_r_15);
not I_58(n30_3,n_572_1_r_15);
nor I_59(n31_3,n40_3,n_569_1_r_15);
nor I_60(n32_3,n25_3,n33_3);
nand I_61(n33_3,n22_3,G214_4_r_15);
or I_62(n34_3,n_569_1_r_15,n_266_and_0_3_r_15);
nand I_63(n35_3,ACVQN1_3_r_3,G214_4_r_15);
nor I_64(n36_3,n_573_1_r_15,G199_4_r_15);
nor I_65(n37_3,n38_3,n39_3);
not I_66(n38_3,n_572_1_l_3);
nand I_67(n39_3,n27_3,n30_3);
endmodule


