module test_I13231(I8854,I11429,I8836,I1477,I1470,I11624,I13231);
input I8854,I11429,I8836,I1477,I1470,I11624;
output I13231;
wire I13214,I11672,I11290,I11720,I11813,I11830,I11275,I11302,I11847,I11460,I11310,I11864;
nand I_0(I13214,I11275,I11302);
DFFARX1 I_1(I8836,I1470,I11310,,,I11672,);
and I_2(I13231,I13214,I11290);
nand I_3(I11290,I11830,I11720);
nor I_4(I11720,I11672,I11460);
DFFARX1 I_5(I8854,I1470,I11310,,,I11813,);
not I_6(I11830,I11813);
DFFARX1 I_7(I11672,I1470,I11310,,,I11275,);
DFFARX1 I_8(I11864,I1470,I11310,,,I11302,);
nand I_9(I11847,I11830);
not I_10(I11460,I11429);
not I_11(I11310,I1477);
and I_12(I11864,I11624,I11847);
endmodule


