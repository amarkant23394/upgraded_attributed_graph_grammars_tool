module test_I1376(I1215,I1223,I1376);
input I1215,I1223;
output I1376;
wire ;
nor I_0(I1376,I1215,I1223);
endmodule


