module test_I13057(I10664,I1477,I10766,I9459,I10732,I1470,I13057);
input I10664,I1477,I10766,I9459,I10732,I1470;
output I13057;
wire I10647,I10961,I10639,I11009,I13040,I13023,I12718,I11184,I10636,I12619,I12735,I10615,I11201,I10630;
not I_0(I10647,I1477);
nand I_1(I10961,I10664,I9459);
DFFARX1 I_2(I11201,I1470,I10647,,,I10639,);
DFFARX1 I_3(I1470,I10647,,,I11009,);
nand I_4(I13040,I13023,I12735);
DFFARX1 I_5(I10636,I1470,I12619,,,I13023,);
nor I_6(I12718,I10615,I10639);
nand I_7(I11184,I10732);
nor I_8(I10636,I10732,I10766);
not I_9(I12619,I1477);
DFFARX1 I_10(I10630,I1470,I12619,,,I12735,);
DFFARX1 I_11(I10961,I1470,I10647,,,I10615,);
and I_12(I13057,I12718,I13040);
and I_13(I11201,I10961,I11184);
not I_14(I10630,I11009);
endmodule


