module test_I13775_rst(I1477_rst,I13775_rst);
,I13775_rst);
input I1477_rst;
output I13775_rst;
wire ;
not I_0(I13775_rst,I1477_rst);
endmodule


