module test_I13792(I12270,I10038,I1477,I10041,I1470,I12024,I13792);
input I12270,I10038,I1477,I10041,I1470,I12024;
output I13792;
wire I12541,I12287,I12304,I12425,I11953,I12349,I10020,I12106,I11973,I12442,I12524,I11965;
nor I_0(I12541,I12349,I12524);
nand I_1(I12287,I12270,I12024);
and I_2(I12304,I12106,I12287);
DFFARX1 I_3(I10038,I1470,I11973,,,I12425,);
nand I_4(I11953,I12442,I12541);
DFFARX1 I_5(I10041,I1470,I11973,,,I12349,);
nand I_6(I13792,I11953,I11965);
DFFARX1 I_7(I1470,,,I10020,);
not I_8(I12106,I10020);
not I_9(I11973,I1477);
not I_10(I12442,I12425);
not I_11(I12524,I12442);
DFFARX1 I_12(I12304,I1470,I11973,,,I11965,);
endmodule


