module test_I7538(I7799,I1477,I1470,I6705,I7538);
input I7799,I1477,I1470,I6705;
output I7538;
wire I7898,I6300,I7816,I7570,I7881,I7587,I6329,I7915,I6291;
nand I_0(I7898,I7881,I7816);
DFFARX1 I_1(I7915,I1470,I7570,,,I7538,);
DFFARX1 I_2(I1470,I6329,,,I6300,);
DFFARX1 I_3(I7799,I1470,I7570,,,I7816,);
not I_4(I7570,I1477);
nand I_5(I7881,I7587,I6291);
not I_6(I7587,I6300);
not I_7(I6329,I1477);
and I_8(I7915,I7881,I7898);
DFFARX1 I_9(I6705,I1470,I6329,,,I6291,);
endmodule


