module test_I6079(I4917,I1477,I4512,I4506,I1470,I4515,I4530,I6079);
input I4917,I1477,I4512,I4506,I1470,I4515,I4530;
output I6079;
wire I4595,I5994,I5751,I6028,I6011,I4521,I4524,I5785,I4742,I5802,I5768,I4544;
DFFARX1 I_0(I1470,I4544,,,I4595,);
nand I_1(I5994,I4512,I4506);
not I_2(I5751,I1477);
DFFARX1 I_3(I6011,I1470,I5751,,,I6028,);
and I_4(I6011,I5994,I4521);
DFFARX1 I_5(I4917,I1470,I4544,,,I4521,);
nor I_6(I4524,I4742,I4595);
nor I_7(I6079,I6028,I5802);
and I_8(I5785,I5768,I4524);
DFFARX1 I_9(I1470,I4544,,,I4742,);
DFFARX1 I_10(I5785,I1470,I5751,,,I5802,);
nand I_11(I5768,I4530,I4515);
not I_12(I4544,I1477);
endmodule


