module test_I16217(I16308,I1477,I1470,I14605,I16217);
input I16308,I1477,I1470,I14605;
output I16217;
wire I14338,I16740,I16339,I16486,I16469,I16240,I16723,I14347,I14353,I14808,I16644,I14370;
DFFARX1 I_0(I14605,I1470,I14370,,,I14338,);
or I_1(I16740,I16339,I16723);
DFFARX1 I_2(I16740,I1470,I16240,,,I16217,);
nor I_3(I16339,I14353,I14338);
nor I_4(I16486,I16469,I16308);
DFFARX1 I_5(I1470,I16240,,,I16469,);
not I_6(I16240,I1477);
and I_7(I16723,I16644,I16486);
DFFARX1 I_8(I1470,I14370,,,I14347,);
not I_9(I14353,I14808);
DFFARX1 I_10(I1470,I14370,,,I14808,);
DFFARX1 I_11(I14347,I1470,I16240,,,I16644,);
not I_12(I14370,I1477);
endmodule


