module test_I15310(I12930,I1477,I15177,I12882,I1470,I15310);
input I12930,I1477,I15177,I12882,I1470;
output I15310;
wire I12596,I10639,I15276,I14965,I12718,I12608,I13119,I15194,I12964,I12619,I14982,I12599,I15211,I10615,I15293;
DFFARX1 I_0(I13119,I1470,I12619,,,I12596,);
DFFARX1 I_1(I1470,,,I10639,);
nand I_2(I15276,I14982,I12599);
and I_3(I15310,I15276,I15293);
not I_4(I14965,I1477);
nor I_5(I12718,I10615,I10639);
nor I_6(I12608,I12930);
or I_7(I13119,I12718);
or I_8(I15194,I15177,I12608);
nor I_9(I12964,I12930,I12882);
not I_10(I12619,I1477);
not I_11(I14982,I12596);
nand I_12(I12599,I12718,I12964);
DFFARX1 I_13(I15194,I1470,I14965,,,I15211,);
DFFARX1 I_14(I1470,,,I10615,);
nand I_15(I15293,I15276,I15211);
endmodule


