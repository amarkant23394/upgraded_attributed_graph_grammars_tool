module test_I11965(I1477,I1470,I11990,I10287,I11965);
input I1477,I1470,I11990,I10287;
output I11965;
wire I12270,I12287,I12304,I10014,I12007,I10020,I10044,I12106,I12024,I11973,I10052;
nand I_0(I12270,I11990,I10014);
nand I_1(I12287,I12270,I12024);
and I_2(I12304,I12106,I12287);
DFFARX1 I_3(I1470,I10052,,,I10014,);
nor I_4(I12007,I10020);
DFFARX1 I_5(I10287,I1470,I10052,,,I10020,);
DFFARX1 I_6(I1470,I10052,,,I10044,);
not I_7(I12106,I10020);
nand I_8(I12024,I12007,I10044);
not I_9(I11973,I1477);
DFFARX1 I_10(I12304,I1470,I11973,,,I11965,);
not I_11(I10052,I1477);
endmodule


