module test_I2070(I1410,I1294,I1492,I1301,I2070);
input I1410,I1294,I1492,I1301;
output I2070;
wire I1444,I1342,I1427,I1509,I1310,I1577;
nand I_0(I1444,I1427,I1410);
not I_1(I1342,I1301);
DFFARX1 I_2(I1294,I1342,,,I1427,);
not I_3(I2070,I1310);
DFFARX1 I_4(I1492,I1294,I1342,,,I1509,);
DFFARX1 I_5(I1577,I1294,I1342,,,I1310,);
and I_6(I1577,I1509,I1444);
endmodule


