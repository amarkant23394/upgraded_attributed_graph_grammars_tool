module test_I11460(I8947,I6881,I9396,I8879,I11460);
input I8947,I6881,I9396,I8879;
output I11460;
wire I9413,I9083,I8848,I11429;
and I_0(I9413,I8947,I9396);
nand I_1(I9083,I8879,I6881);
not I_2(I11460,I11429);
nor I_3(I8848,I9083,I9413);
not I_4(I11429,I8848);
endmodule


