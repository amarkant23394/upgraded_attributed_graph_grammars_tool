module test_I15177(I13040,I12831,I12718,I1477,I10627,I1470,I12636,I15177);
input I13040,I12831,I12718,I1477,I10627,I1470,I12636;
output I15177;
wire I12619,I12670,I15160,I15143,I12599,I13057,I12593,I12653,I12964,I12882,I12848,I12611;
not I_0(I12619,I1477);
DFFARX1 I_1(I12653,I1470,I12619,,,I12670,);
and I_2(I15177,I15160,I12593);
nor I_3(I15160,I15143,I12611);
not I_4(I15143,I12599);
nand I_5(I12599,I12718,I12964);
and I_6(I13057,I12718,I13040);
nand I_7(I12593,I12670,I12882);
and I_8(I12653,I12636,I10627);
nor I_9(I12964,I12882);
not I_10(I12882,I12848);
DFFARX1 I_11(I12831,I1470,I12619,,,I12848,);
DFFARX1 I_12(I13057,I1470,I12619,,,I12611,);
endmodule


