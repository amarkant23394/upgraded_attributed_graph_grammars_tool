module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_4,blif_reset_net_1_r_4,G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_4,blif_reset_net_1_r_4;
output G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4;
wire G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6,N3_2_l_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6,n_431_0_l_4,n6_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4;
DFFARX1 I_0(n4_1_r_6,blif_clk_net_1_r_4,n6_4,G42_1_r_6,);
nor I_1(n_572_1_r_6,n27_6,n28_6);
nand I_2(n_573_1_r_6,n18_6,n19_6);
nor I_3(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_4(n_569_1_r_6,n19_6,n20_6);
nor I_5(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_6(N1_4_r_6,blif_clk_net_1_r_4,n6_4,G199_4_r_6,);
DFFARX1 I_7(n_42_2_l_6,blif_clk_net_1_r_4,n6_4,G214_4_r_6,);
DFFARX1 I_8(n_42_2_l_6,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_6,);
not I_9(P6_5_r_6,P6_5_r_internal_6);
and I_10(N3_2_l_6,IN_6_2_l_6,n23_6);
DFFARX1 I_11(N3_2_l_6,blif_clk_net_1_r_4,n6_4,n27_6,);
not I_12(n17_6,n27_6);
DFFARX1 I_13(IN_1_3_l_6,blif_clk_net_1_r_4,n6_4,n28_6,);
DFFARX1 I_14(IN_2_3_l_6,blif_clk_net_1_r_4,n6_4,n26_6,);
and I_15(N1_4_l_6,IN_6_4_l_6,n25_6);
DFFARX1 I_16(N1_4_l_6,blif_clk_net_1_r_4,n6_4,n29_6,);
not I_17(n18_6,n29_6);
DFFARX1 I_18(IN_3_4_l_6,blif_clk_net_1_r_4,n6_4,G214_4_l_6,);
not I_19(n12_6,G214_4_l_6);
nor I_20(n4_1_r_6,n28_6,n22_6);
nor I_21(N1_4_r_6,n12_6,n24_6);
nor I_22(n_42_2_l_6,IN_1_2_l_6,IN_3_2_l_6);
DFFARX1 I_23(G214_4_l_6,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_6,);
nand I_24(n19_6,IN_4_3_l_6,n26_6);
not I_25(n20_6,n_42_2_l_6);
nor I_26(n21_6,n17_6,n28_6);
and I_27(n22_6,IN_4_3_l_6,n26_6);
nand I_28(n23_6,IN_2_2_l_6,IN_3_2_l_6);
nor I_29(n24_6,n17_6,n18_6);
nand I_30(n25_6,IN_1_4_l_6,IN_2_4_l_6);
DFFARX1 I_31(n4_1_r_4,blif_clk_net_1_r_4,n6_4,G42_1_r_4,);
nor I_32(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_33(n_573_1_r_4,n16_4,n_452_1_r_6);
nor I_34(n_549_1_r_4,n22_4,n23_4);
nand I_35(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_36(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_4,);
nor I_37(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_38(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_4,);
not I_39(P6_5_r_4,P6_5_r_internal_4);
or I_40(n_431_0_l_4,n26_4,P6_5_r_6);
not I_41(n6_4,blif_reset_net_1_r_4);
DFFARX1 I_42(n_431_0_l_4,blif_clk_net_1_r_4,n6_4,G78_0_l_4,);
DFFARX1 I_43(ACVQN1_5_r_6,blif_clk_net_1_r_4,n6_4,ACVQN1_5_l_4,);
not I_44(n16_4,ACVQN1_5_l_4);
DFFARX1 I_45(n_569_1_r_6,blif_clk_net_1_r_4,n6_4,n17_internal_4,);
not I_46(n17_4,n17_internal_4);
nor I_47(n4_1_r_4,n30_4,n31_4);
nand I_48(n19_4,n33_4,G42_1_r_6);
DFFARX1 I_49(G78_0_l_4,blif_clk_net_1_r_4,n6_4,n15_internal_4,);
not I_50(n15_4,n15_internal_4);
DFFARX1 I_51(ACVQN1_5_l_4,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_4,);
and I_52(n20_4,n16_4,G214_4_r_6);
nor I_53(n21_4,n_452_1_r_6,G199_4_r_6);
nand I_54(n22_4,G78_0_l_4,n25_4);
nand I_55(n23_4,n24_4,G214_4_r_6);
not I_56(n24_4,n_452_1_r_6);
not I_57(n25_4,G199_4_r_6);
and I_58(n26_4,n27_4,n_572_1_r_6);
nor I_59(n27_4,n28_4,n_573_1_r_6);
not I_60(n28_4,G42_1_r_6);
not I_61(n29_4,n30_4);
nand I_62(n30_4,n32_4,G42_1_r_6);
nand I_63(n31_4,n25_4,G214_4_r_6);
nor I_64(n32_4,n33_4,n_452_1_r_6);
not I_65(n33_4,n_549_1_r_6);
endmodule


