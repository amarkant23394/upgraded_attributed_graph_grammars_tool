module test_final(G1_0_l_11,G2_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_5_0_l_11,IN_7_0_l_11,IN_8_0_l_11,IN_10_0_l_11,IN_11_0_l_11,IN_1_5_l_11,IN_2_5_l_11,blif_clk_net_1_r_1,blif_reset_net_1_r_1,G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1);
input G1_0_l_11,G2_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_5_0_l_11,IN_7_0_l_11,IN_8_0_l_11,IN_10_0_l_11,IN_11_0_l_11,IN_1_5_l_11,IN_2_5_l_11,blif_clk_net_1_r_1,blif_reset_net_1_r_1;
output G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1;
wire G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11,n_431_0_l_11,n43_11,n26_11,n44_11,n45_11,n27_11,n4_1_r_11,N3_2_r_11,n24_11,n25_11,n20_internal_11,n20_11,n28_11,n29_11,n30_11,n31_11,n32_11,n33_11,n34_11,n35_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,N3_2_l_1,n5_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1;
DFFARX1 I_0(n4_1_r_11,blif_clk_net_1_r_1,n5_1,G42_1_r_11,);
nor I_1(n_572_1_r_11,n29_11,n30_11);
nand I_2(n_573_1_r_11,n26_11,n28_11);
nor I_3(n_549_1_r_11,n27_11,n32_11);
nand I_4(n_569_1_r_11,n45_11,n28_11);
nor I_5(n_452_1_r_11,n43_11,n44_11);
nor I_6(n_42_2_r_11,n35_11,n36_11);
DFFARX1 I_7(N3_2_r_11,blif_clk_net_1_r_1,n5_1,G199_2_r_11,);
DFFARX1 I_8(n24_11,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_11,);
nor I_9(n_266_and_0_3_r_11,n20_11,n37_11);
or I_10(n_431_0_l_11,IN_8_0_l_11,n33_11);
DFFARX1 I_11(n_431_0_l_11,blif_clk_net_1_r_1,n5_1,n43_11,);
not I_12(n26_11,n43_11);
DFFARX1 I_13(IN_2_5_l_11,blif_clk_net_1_r_1,n5_1,n44_11,);
DFFARX1 I_14(IN_1_5_l_11,blif_clk_net_1_r_1,n5_1,n45_11,);
not I_15(n27_11,n45_11);
nor I_16(n4_1_r_11,n44_11,n25_11);
nor I_17(N3_2_r_11,n45_11,n40_11);
nand I_18(n24_11,IN_11_0_l_11,n39_11);
nand I_19(n25_11,IN_7_0_l_11,n38_11);
DFFARX1 I_20(n25_11,blif_clk_net_1_r_1,n5_1,n20_internal_11,);
not I_21(n20_11,n20_internal_11);
not I_22(n28_11,n25_11);
not I_23(n29_11,G1_0_l_11);
nand I_24(n30_11,n26_11,n31_11);
not I_25(n31_11,IN_5_0_l_11);
and I_26(n32_11,n26_11,n44_11);
and I_27(n33_11,IN_2_0_l_11,n34_11);
nor I_28(n34_11,IN_4_0_l_11,n29_11);
not I_29(n35_11,G2_0_l_11);
nand I_30(n36_11,G1_0_l_11,n31_11);
nor I_31(n37_11,IN_5_0_l_11,n29_11);
nor I_32(n38_11,G2_0_l_11,n31_11);
nor I_33(n39_11,G2_0_l_11,IN_10_0_l_11);
nor I_34(n40_11,G2_0_l_11,n41_11);
nor I_35(n41_11,IN_10_0_l_11,n42_11);
not I_36(n42_11,IN_11_0_l_11);
DFFARX1 I_37(n4_1_r_1,blif_clk_net_1_r_1,n5_1,G42_1_r_1,);
nor I_38(n_572_1_r_1,n26_1,n19_1);
nand I_39(n_573_1_r_1,n16_1,n18_1);
nor I_40(n_549_1_r_1,n20_1,n21_1);
nor I_41(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_42(G199_4_l_1,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_1,);
nor I_43(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_44(N1_4_r_1,blif_clk_net_1_r_1,n5_1,G199_4_r_1,);
DFFARX1 I_45(G199_4_l_1,blif_clk_net_1_r_1,n5_1,G214_4_r_1,);
and I_46(N3_2_l_1,n23_1,G199_2_r_11);
not I_47(n5_1,blif_reset_net_1_r_1);
DFFARX1 I_48(N3_2_l_1,blif_clk_net_1_r_1,n5_1,n26_1,);
not I_49(n17_1,n26_1);
DFFARX1 I_50(n_573_1_r_11,blif_clk_net_1_r_1,n5_1,n16_internal_1,);
not I_51(n16_1,n16_internal_1);
DFFARX1 I_52(ACVQN2_3_r_11,blif_clk_net_1_r_1,n5_1,ACVQN1_3_l_1,);
and I_53(N1_4_l_1,n25_1,n_549_1_r_11);
DFFARX1 I_54(N1_4_l_1,blif_clk_net_1_r_1,n5_1,G199_4_l_1,);
DFFARX1 I_55(n_572_1_r_11,blif_clk_net_1_r_1,n5_1,G214_4_l_1,);
nor I_56(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_57(G214_4_l_1,blif_clk_net_1_r_1,n5_1,n14_internal_1,);
not I_58(n14_1,n14_internal_1);
nor I_59(N1_4_r_1,n17_1,n24_1);
nand I_60(n18_1,ACVQN1_3_l_1,n_266_and_0_3_r_11);
nor I_61(n19_1,n_569_1_r_11,n_42_2_r_11);
not I_62(n20_1,n18_1);
nor I_63(n21_1,n26_1,n22_1);
not I_64(n22_1,n19_1);
nand I_65(n23_1,n_42_2_r_11,G42_1_r_11);
nor I_66(n24_1,n18_1,n22_1);
nand I_67(n25_1,G42_1_r_11,n_452_1_r_11);
endmodule


