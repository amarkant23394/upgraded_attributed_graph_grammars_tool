module test_I15293(I12930,I1477,I12882,I15160,I1470,I15293);
input I12930,I1477,I12882,I15160,I1470;
output I15293;
wire I12596,I10639,I15276,I14965,I13023,I12718,I12608,I13119,I15194,I12593,I12964,I12619,I14982,I15177,I12599,I15211,I10615;
DFFARX1 I_0(I13119,I1470,I12619,,,I12596,);
DFFARX1 I_1(I1470,,,I10639,);
nand I_2(I15276,I14982,I12599);
not I_3(I14965,I1477);
DFFARX1 I_4(I1470,I12619,,,I13023,);
nor I_5(I12718,I10615,I10639);
nor I_6(I12608,I13023,I12930);
or I_7(I13119,I12718);
or I_8(I15194,I15177,I12608);
nand I_9(I12593,I12882);
nor I_10(I12964,I12930,I12882);
not I_11(I12619,I1477);
not I_12(I14982,I12596);
and I_13(I15177,I15160,I12593);
nand I_14(I12599,I12718,I12964);
DFFARX1 I_15(I15194,I1470,I14965,,,I15211,);
DFFARX1 I_16(I1470,,,I10615,);
nand I_17(I15293,I15276,I15211);
endmodule


