module test_final(IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_7_r_3,blif_reset_net_7_r_3,N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3);
input IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_7_r_3,blif_reset_net_7_r_3;
output N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3;
wire N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_102_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7,n_452_7_r_7,n4_7_l_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7,n_572_7_r_3,N6147_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n10_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3;
nor I_0(N1371_0_r_7,n53_7,n52_7);
nor I_1(N1508_0_r_7,n51_7,n52_7);
nand I_2(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_3(n_431_5_r_7,blif_clk_net_7_r_3,n10_3,G78_5_r_7,);
nand I_4(n_576_5_r_7,n31_7,n32_7);
nor I_5(n_102_5_r_7,IN_5_7_l_7,IN_9_7_l_7);
nand I_6(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_7(n4_7_r_7,blif_clk_net_7_r_3,n10_3,G42_7_r_7,);
nor I_8(n_572_7_r_7,n54_7,n33_7);
nand I_9(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_10(n_549_7_r_7,n53_7,n36_7);
nand I_11(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_12(n_452_7_r_7,IN_1_1_l_7,IN_2_1_l_7);
nor I_13(n4_7_l_7,G18_7_l_7,IN_1_7_l_7);
DFFARX1 I_14(n4_7_l_7,blif_clk_net_7_r_3,n10_3,n53_7,);
not I_15(n30_7,n53_7);
and I_16(N3_8_l_7,IN_6_8_l_7,n50_7);
DFFARX1 I_17(N3_8_l_7,blif_clk_net_7_r_3,n10_3,n54_7,);
nand I_18(n_431_5_r_7,n40_7,n41_7);
nor I_19(n4_7_r_7,n54_7,n49_7);
and I_20(n31_7,n_102_5_r_7,n39_7);
not I_21(n32_7,G18_7_l_7);
nor I_22(n33_7,IN_10_7_l_7,n34_7);
and I_23(n34_7,IN_4_7_l_7,n35_7);
not I_24(n35_7,G15_7_l_7);
nor I_25(n36_7,G18_7_l_7,n37_7);
or I_26(n37_7,IN_5_7_l_7,n54_7);
or I_27(n38_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_28(n39_7,IN_3_1_l_7,n_452_7_r_7);
nand I_29(n40_7,n46_7,n47_7);
nand I_30(n41_7,n42_7,n43_7);
nor I_31(n42_7,n44_7,n45_7);
nor I_32(n43_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_33(n44_7,G15_7_l_7,IN_7_7_l_7);
nor I_34(n45_7,IN_9_7_l_7,IN_10_7_l_7);
nand I_35(n46_7,IN_4_7_l_7,n35_7);
not I_36(n47_7,IN_10_7_l_7);
or I_37(n48_7,IN_3_1_l_7,n_452_7_r_7);
not I_38(n49_7,n_452_7_r_7);
nand I_39(n50_7,IN_2_8_l_7,IN_3_8_l_7);
and I_40(n51_7,n_452_7_r_7,n45_7);
not I_41(n52_7,n44_7);
not I_42(N1372_1_r_3,n40_3);
nor I_43(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_44(N1507_6_r_3,n31_3,n42_3);
nor I_45(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_46(n4_7_r_3,blif_clk_net_7_r_3,n10_3,G42_7_r_3,);
nor I_47(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_48(n_573_7_r_3,n30_3,n31_3);
nor I_49(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_50(n_569_7_r_3,n30_3,n32_3);
nor I_51(n_452_7_r_3,n35_3,N1371_0_r_7);
not I_52(N6147_9_r_3,n32_3);
nor I_53(N6134_9_r_3,n36_3,n37_3);
not I_54(I_BUFF_1_9_r_3,n45_3);
nor I_55(n4_7_r_3,I_BUFF_1_9_r_3,N1371_0_r_7);
not I_56(n10_3,blif_reset_net_7_r_3);
not I_57(n30_3,n39_3);
not I_58(n31_3,n35_3);
nand I_59(n32_3,n41_3,G78_5_r_7);
nor I_60(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_61(n34_3,n46_3,n_429_or_0_5_r_7);
nor I_62(n35_3,n43_3,n44_3);
not I_63(n36_3,n34_3);
nor I_64(n37_3,N6147_9_r_3,N1371_0_r_7);
or I_65(n38_3,n_572_7_r_3,n34_3);
nor I_66(n39_3,n44_3,n_547_5_r_7);
nand I_67(n40_3,n39_3,N1371_0_r_7);
nand I_68(n41_3,N1508_0_r_7,n_549_7_r_7);
nor I_69(n42_3,n34_3,n45_3);
not I_70(n43_3,n_572_7_r_7);
nor I_71(n44_3,G78_5_r_7,n_576_5_r_7);
nand I_72(n45_3,n49_3,n50_3);
and I_73(n46_3,n47_3,n_569_7_r_7);
nand I_74(n47_3,n41_3,n48_3);
not I_75(n48_3,G78_5_r_7);
nor I_76(n49_3,N1371_0_r_7,n_429_or_0_5_r_7);
or I_77(n50_3,n51_3,n_573_7_r_7);
nor I_78(n51_3,G42_7_r_7,N1508_0_r_7);
endmodule


