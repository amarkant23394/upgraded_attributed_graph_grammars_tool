module test_I1586(I1455,I1215,I1586);
input I1455,I1215;
output I1586;
wire I1535;
nor I_0(I1586,I1535,I1215);
not I_1(I1535,I1455);
endmodule


