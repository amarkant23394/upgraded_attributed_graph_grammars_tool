module test_I3103(I1301,I1294,I1331,I3103);
input I1301,I1294,I1331;
output I3103;
wire I2583,I2313,I1937,I3086,I1920;
not I_0(I2583,I1301);
DFFARX1 I_1(I1331,I1294,I1937,,,I2313,);
not I_2(I1937,I1301);
DFFARX1 I_3(I1920,I1294,I2583,,,I3086,);
not I_4(I3103,I3086);
not I_5(I1920,I2313);
endmodule


