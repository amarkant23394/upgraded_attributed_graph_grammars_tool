module test_I14588(I1477,I11299,I14520,I1470,I14588);
input I1477,I11299,I14520,I1470;
output I14588;
wire I14554,I13183,I14421,I13601,I13186,I14537,I14387,I14370,I13197,I13159,I14438,I14571,I11272,I14404,I13508,I13491;
not I_0(I14554,I14537);
nand I_1(I13183,I13601);
DFFARX1 I_2(I14404,I1470,I14370,,,I14421,);
DFFARX1 I_3(I11299,I1470,I13197,,,I13601,);
nor I_4(I13186,I13601,I13508);
DFFARX1 I_5(I14520,I1470,I14370,,,I14537,);
nand I_6(I14387,I13186);
not I_7(I14370,I1477);
not I_8(I13197,I1477);
DFFARX1 I_9(I13508,I1470,I13197,,,I13159,);
nor I_10(I14438,I13159,I13186);
nor I_11(I14571,I14421,I14554);
DFFARX1 I_12(I1470,,,I11272,);
and I_13(I14404,I14387,I13183);
and I_14(I13508,I13491,I11272);
and I_15(I14588,I14438,I14571);
DFFARX1 I_16(I1470,I13197,,,I13491,);
endmodule


