module test_I1552(I1215,I1399,I1552);
input I1215,I1399;
output I1552;
wire ;
nor I_0(I1552,I1215,I1399);
endmodule


