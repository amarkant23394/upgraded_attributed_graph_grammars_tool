module test_final(IN_1_1_l_3,IN_2_1_l_3,IN_3_1_l_3,IN_1_8_l_3,IN_2_8_l_3,IN_3_8_l_3,IN_6_8_l_3,IN_1_10_l_3,IN_2_10_l_3,IN_3_10_l_3,IN_4_10_l_3,blif_clk_net_5_r_6,blif_reset_net_5_r_6,N1371_0_r_6,N1508_0_r_6,N6147_3_r_6,G78_5_r_6,n_576_5_r_6,n_547_5_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_1_l_3,IN_2_1_l_3,IN_3_1_l_3,IN_1_8_l_3,IN_2_8_l_3,IN_3_8_l_3,IN_6_8_l_3,IN_1_10_l_3,IN_2_10_l_3,IN_3_10_l_3,IN_4_10_l_3,blif_clk_net_5_r_6,blif_reset_net_5_r_6;
output N1371_0_r_6,N1508_0_r_6,N6147_3_r_6,G78_5_r_6,n_576_5_r_6,n_547_5_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_3,N1508_0_r_3,N6147_3_r_3,n_429_or_0_5_r_3,G78_5_r_3,n_576_5_r_3,n_102_5_r_3,n_547_5_r_3,N1372_10_r_3,N1508_10_r_3,N3_8_l_3,n39_3,n_431_5_r_3,n22_3,n23_3,n24_3,n25_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n_429_or_0_5_r_6,n_102_5_r_6,n_431_5_r_6,n6_6,n24_6,n25_6,n26_6,n27_6,n28_6,n29_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6;
nor I_0(N1371_0_r_3,n39_3,n37_3);
nor I_1(N1508_0_r_3,n25_3,n37_3);
nor I_2(N6147_3_r_3,N1372_10_r_3,n33_3);
nand I_3(n_429_or_0_5_r_3,N1372_10_r_3,n30_3);
DFFARX1 I_4(n_431_5_r_3,blif_clk_net_5_r_6,n6_6,G78_5_r_3,);
nand I_5(n_576_5_r_3,n22_3,n23_3);
not I_6(n_102_5_r_3,n39_3);
nand I_7(n_547_5_r_3,n26_3,n27_3);
not I_8(N1372_10_r_3,n36_3);
nor I_9(N1508_10_r_3,n35_3,n36_3);
and I_10(N3_8_l_3,IN_6_8_l_3,n34_3);
DFFARX1 I_11(N3_8_l_3,blif_clk_net_5_r_6,n6_6,n39_3,);
nand I_12(n_431_5_r_3,n29_3,n30_3);
nor I_13(n22_3,n24_3,n25_3);
nor I_14(n23_3,IN_3_1_l_3,n39_3);
not I_15(n24_3,n27_3);
nand I_16(n25_3,IN_1_1_l_3,IN_2_1_l_3);
nor I_17(n26_3,n39_3,n28_3);
nor I_18(n27_3,IN_1_8_l_3,IN_3_8_l_3);
not I_19(n28_3,n37_3);
nand I_20(n29_3,N1372_10_r_3,n39_3);
nand I_21(n30_3,n31_3,n32_3);
not I_22(n31_3,n25_3);
not I_23(n32_3,IN_3_1_l_3);
nand I_24(n33_3,n24_3,n25_3);
nand I_25(n34_3,IN_2_8_l_3,IN_3_8_l_3);
nor I_26(n35_3,n27_3,n31_3);
nand I_27(n36_3,n28_3,n38_3);
nand I_28(n37_3,IN_1_10_l_3,IN_2_10_l_3);
or I_29(n38_3,IN_3_10_l_3,IN_4_10_l_3);
nor I_30(N1371_0_r_6,n26_6,n38_6);
not I_31(N1508_0_r_6,n38_6);
nor I_32(N6147_3_r_6,n30_6,n35_6);
nand I_33(n_429_or_0_5_r_6,n30_6,n32_6);
DFFARX1 I_34(n_431_5_r_6,blif_clk_net_5_r_6,n6_6,G78_5_r_6,);
nand I_35(n_576_5_r_6,n24_6,n25_6);
not I_36(n_102_5_r_6,n26_6);
or I_37(n_547_5_r_6,n_429_or_0_5_r_6,n26_6);
not I_38(N1372_10_r_6,n37_6);
nor I_39(N1508_10_r_6,n36_6,n37_6);
nand I_40(n_431_5_r_6,n_102_5_r_6,n28_6);
not I_41(n6_6,blif_reset_net_5_r_6);
nor I_42(n24_6,n33_6,n34_6);
nor I_43(n25_6,n26_6,n27_6);
nor I_44(n26_6,n40_6,N6147_3_r_3);
nand I_45(n27_6,N1508_0_r_3,n_547_5_r_3);
nand I_46(n28_6,n29_6,n30_6);
nor I_47(n29_6,n31_6,n_429_or_0_5_r_3);
not I_48(n30_6,n27_6);
nor I_49(n31_6,n39_6,n40_6);
nor I_50(n32_6,n24_6,n_429_or_0_5_r_3);
not I_51(n33_6,G78_5_r_3);
not I_52(n34_6,N1508_0_r_3);
or I_53(n35_6,n26_6,n31_6);
and I_54(n36_6,n38_6,n_429_or_0_5_r_3);
nand I_55(n37_6,n30_6,n31_6);
nand I_56(n38_6,n41_6,N1508_0_r_3);
nor I_57(n39_6,N1371_0_r_3,N1508_10_r_3);
not I_58(n40_6,N1371_0_r_3);
nor I_59(n41_6,n33_6,n42_6);
nor I_60(n42_6,n_576_5_r_3,n_102_5_r_3);
endmodule


