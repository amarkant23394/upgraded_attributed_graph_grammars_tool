module test_I15611_rst(I1477_rst,I15611_rst);
,I15611_rst);
input I1477_rst;
output I15611_rst;
wire ;
not I_0(I15611_rst,I1477_rst);
endmodule


