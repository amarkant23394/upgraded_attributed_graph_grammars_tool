module test_final(IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_7_r_3,blif_reset_net_7_r_3,N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3);
input IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_7_r_3,blif_reset_net_7_r_3;
output N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3;
wire N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,n_429_or_0_5_r_9,G78_5_r_9,n_576_5_r_9,n_102_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9,n_572_7_r_3,N6147_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n10_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3;
nor I_0(N6147_2_r_9,n62_9,n46_9);
not I_1(N1372_4_r_9,n59_9);
nor I_2(N1508_4_r_9,n58_9,n59_9);
nand I_3(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_4(n_431_5_r_9,blif_clk_net_7_r_3,n10_3,G78_5_r_9,);
nand I_5(n_576_5_r_9,n39_9,n40_9);
not I_6(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_7(n_547_5_r_9,IN_3_1_l_9,n43_9);
and I_8(n_42_8_r_9,G18_7_l_9,n44_9);
DFFARX1 I_9(N3_8_r_9,blif_clk_net_7_r_3,n10_3,G199_8_r_9,);
nor I_10(N6147_9_r_9,n41_9,n45_9);
nor I_11(N6134_9_r_9,n45_9,n51_9);
nor I_12(I_BUFF_1_9_r_9,IN_3_1_l_9,n41_9);
nor I_13(n4_7_l_9,G18_7_l_9,IN_1_7_l_9);
DFFARX1 I_14(n4_7_l_9,blif_clk_net_7_r_3,n10_3,n62_9,);
and I_15(N3_8_l_9,IN_6_8_l_9,n57_9);
DFFARX1 I_16(N3_8_l_9,blif_clk_net_7_r_3,n10_3,n63_9,);
not I_17(n38_9,n63_9);
nor I_18(n_431_5_r_9,G15_7_l_9,IN_7_7_l_9);
nor I_19(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_20(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_21(n40_9,n41_9);
nand I_22(n41_9,IN_1_1_l_9,IN_2_1_l_9);
nor I_23(n42_9,IN_9_7_l_9,IN_10_7_l_9);
nor I_24(n43_9,n63_9,n41_9);
nor I_25(n44_9,IN_5_7_l_9,IN_9_7_l_9);
and I_26(n45_9,IN_4_7_l_9,n52_9);
nor I_27(n46_9,n47_9,n48_9);
nor I_28(n47_9,n49_9,n50_9);
not I_29(n48_9,n_429_or_0_5_r_9);
not I_30(n49_9,n42_9);
or I_31(n50_9,n63_9,n51_9);
nor I_32(n51_9,IN_1_8_l_9,IN_3_8_l_9);
nor I_33(n52_9,G15_7_l_9,n49_9);
nor I_34(n53_9,n54_9,n55_9);
nor I_35(n54_9,G15_7_l_9,n56_9);
or I_36(n55_9,IN_10_7_l_9,n44_9);
not I_37(n56_9,IN_4_7_l_9);
nand I_38(n57_9,IN_2_8_l_9,IN_3_8_l_9);
nor I_39(n58_9,n62_9,n60_9);
nand I_40(n59_9,n51_9,n61_9);
nor I_41(n60_9,n38_9,n44_9);
nor I_42(n61_9,G18_7_l_9,IN_5_7_l_9);
not I_43(N1372_1_r_3,n40_3);
nor I_44(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_45(N1507_6_r_3,n31_3,n42_3);
nor I_46(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_47(n4_7_r_3,blif_clk_net_7_r_3,n10_3,G42_7_r_3,);
nor I_48(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_49(n_573_7_r_3,n30_3,n31_3);
nor I_50(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_51(n_569_7_r_3,n30_3,n32_3);
nor I_52(n_452_7_r_3,n35_3,n_547_5_r_9);
not I_53(N6147_9_r_3,n32_3);
nor I_54(N6134_9_r_3,n36_3,n37_3);
not I_55(I_BUFF_1_9_r_3,n45_3);
nor I_56(n4_7_r_3,I_BUFF_1_9_r_3,n_547_5_r_9);
not I_57(n10_3,blif_reset_net_7_r_3);
not I_58(n30_3,n39_3);
not I_59(n31_3,n35_3);
nand I_60(n32_3,n41_3,N1508_4_r_9);
nor I_61(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_62(n34_3,n46_3,N6147_2_r_9);
nor I_63(n35_3,n43_3,n44_3);
not I_64(n36_3,n34_3);
nor I_65(n37_3,N6147_9_r_3,n_547_5_r_9);
or I_66(n38_3,n_572_7_r_3,n34_3);
nor I_67(n39_3,n44_3,n_42_8_r_9);
nand I_68(n40_3,n39_3,n_547_5_r_9);
nand I_69(n41_3,N1372_4_r_9,n_576_5_r_9);
nor I_70(n42_3,n34_3,n45_3);
not I_71(n43_3,N6147_2_r_9);
nor I_72(n44_3,N6147_9_r_9,N1372_4_r_9);
nand I_73(n45_3,n49_3,n50_3);
and I_74(n46_3,n47_3,G199_8_r_9);
nand I_75(n47_3,n41_3,n48_3);
not I_76(n48_3,N1508_4_r_9);
nor I_77(n49_3,G78_5_r_9,N6134_9_r_9);
or I_78(n50_3,n51_3,n_576_5_r_9);
nor I_79(n51_3,N1508_4_r_9,G78_5_r_9);
endmodule


