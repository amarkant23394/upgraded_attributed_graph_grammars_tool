module test_I1518(I1477,I1518);
input I1477;
output I1518;
wire ;
not I_0(I1518,I1477);
endmodule


