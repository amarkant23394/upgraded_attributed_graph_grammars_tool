module test_final(IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_549_7_r_5,n_569_7_r_5,n_452_7_r_5,n4_7_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
nor I_0(N1371_0_r_5,n28_5,n46_5);
nand I_1(N1508_0_r_5,n26_5,n43_5);
not I_2(N1372_1_r_5,n43_5);
nor I_3(N1508_1_r_5,n30_5,n43_5);
nor I_4(N6147_2_r_5,n29_5,n32_5);
nor I_5(N1507_6_r_5,n26_5,n44_5);
nor I_6(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_7(n4_7_r_5,blif_clk_net_7_r_1,n9_1,G42_7_r_5,);
and I_8(n_572_7_r_5,n27_5,n28_5);
nand I_9(n_573_7_r_5,n26_5,n27_5);
nand I_10(n_549_7_r_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_11(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_12(n_452_7_r_5,n29_5);
nor I_13(n4_7_r_5,n30_5,n31_5);
not I_14(n26_5,n35_5);
nand I_15(n27_5,n40_5,n41_5);
nand I_16(n28_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_17(n29_5,n27_5,n33_5);
nor I_18(n30_5,IN_1_3_l_5,n45_5);
not I_19(n31_5,n_549_7_r_5);
nor I_20(n32_5,n34_5,n35_5);
not I_21(n33_5,n30_5);
nor I_22(n34_5,n31_5,n36_5);
nor I_23(n35_5,IN_3_1_l_5,n28_5);
not I_24(n36_5,n28_5);
nand I_25(n37_5,n36_5,n38_5);
nand I_26(n38_5,n26_5,n39_5);
nand I_27(n39_5,n30_5,n31_5);
nor I_28(n40_5,IN_1_2_l_5,IN_2_2_l_5);
or I_29(n41_5,IN_5_2_l_5,n42_5);
nor I_30(n42_5,IN_3_2_l_5,IN_4_2_l_5);
nand I_31(n43_5,n36_5,n46_5);
nor I_32(n44_5,n_549_7_r_5,n33_5);
or I_33(n45_5,IN_2_3_l_5,IN_3_3_l_5);
and I_34(n46_5,n31_5,n47_5);
or I_35(n47_5,IN_3_10_l_5,IN_4_10_l_5);
and I_36(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_37(N1508_0_r_1,n40_1,n44_1);
nor I_38(N1507_6_r_1,n43_1,n49_1);
nor I_39(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_40(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_41(n_572_7_r_1,n29_1,n30_1);
not I_42(n_573_7_r_1,n_452_7_r_1);
nor I_43(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_44(n_569_7_r_1,n30_1,n31_1);
nor I_45(n_452_7_r_1,n30_1,n32_1);
nor I_46(N6147_9_r_1,n35_1,n36_1);
nand I_47(N6134_9_r_1,n38_1,n39_1);
not I_48(I_BUFF_1_9_r_1,n40_1);
nor I_49(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_50(n9_1,blif_reset_net_7_r_1);
nor I_51(n29_1,n34_1,n_569_7_r_5);
nor I_52(n30_1,n33_1,n34_1);
nor I_53(n31_1,n54_1,N1371_0_r_5);
not I_54(n32_1,n48_1);
nor I_55(n33_1,N6147_2_r_5,N1372_1_r_5);
not I_56(n34_1,N1508_0_r_5);
nor I_57(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_58(n36_1,n29_1);
not I_59(n37_1,n41_1);
nand I_60(n38_1,I_BUFF_1_9_r_1,N1371_0_r_5);
nand I_61(n39_1,n37_1,n40_1);
nand I_62(n40_1,N1508_1_r_5,N1508_0_r_5);
nand I_63(n41_1,n52_1,n_572_7_r_5);
or I_64(n42_1,n36_1,n43_1);
nor I_65(n43_1,n32_1,n49_1);
nand I_66(n44_1,n45_1,n46_1);
nand I_67(n45_1,n47_1,n48_1);
not I_68(n46_1,N1371_0_r_5);
not I_69(n47_1,n31_1);
nand I_70(n48_1,n50_1,N1507_6_r_5);
nor I_71(n49_1,n41_1,n47_1);
and I_72(n50_1,n51_1,N1372_1_r_5);
nand I_73(n51_1,n52_1,n53_1);
nand I_74(n52_1,N1508_6_r_5,n_573_7_r_5);
not I_75(n53_1,n_572_7_r_5);
or I_76(n54_1,G42_7_r_5,n_452_7_r_5);
nor I_77(n55_1,n29_1,N1371_0_r_5);
endmodule


