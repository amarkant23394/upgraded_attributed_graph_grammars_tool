module test_I16644(I14571,I1477,I1470,I14438,I16644);
input I14571,I1477,I1470,I14438;
output I16644;
wire I14667,I13189,I14777,I14347,I16240,I14588,I14650,I14370;
and I_0(I14667,I14650,I13189);
DFFARX1 I_1(I1470,,,I13189,);
or I_2(I14777,I14667,I14588);
DFFARX1 I_3(I14777,I1470,I14370,,,I14347,);
not I_4(I16240,I1477);
and I_5(I14588,I14438,I14571);
DFFARX1 I_6(I14347,I1470,I16240,,,I16644,);
DFFARX1 I_7(I1470,I14370,,,I14650,);
not I_8(I14370,I1477);
endmodule


