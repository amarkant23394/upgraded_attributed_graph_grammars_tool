module test_I13542(I11751,I11429,I13392,I1477,I11281,I1470,I11689,I13542);
input I11751,I11429,I13392,I1477,I11281,I1470,I11689;
output I13542;
wire I11559,I11296,I13197,I13426,I11768,I11272,I13409,I13508,I13460,I11310,I13491;
DFFARX1 I_0(I1470,I11310,,,I11559,);
nand I_1(I11296,I11559,I11689);
not I_2(I13197,I1477);
nor I_3(I13542,I13508,I13460);
DFFARX1 I_4(I13409,I1470,I13197,,,I13426,);
and I_5(I11768,I11429,I11751);
DFFARX1 I_6(I11768,I1470,I11310,,,I11272,);
and I_7(I13409,I13392,I11281);
and I_8(I13508,I13491,I11272);
not I_9(I13460,I13426);
not I_10(I11310,I1477);
DFFARX1 I_11(I11296,I1470,I13197,,,I13491,);
endmodule


