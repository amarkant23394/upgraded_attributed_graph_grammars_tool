module test_I2569(I2600,I2781,I2234,I1908,I1294,I2406,I1301,I2505,I2569);
input I2600,I2781,I2234,I1908,I1294,I2406,I1301,I2505;
output I2569;
wire I2668,I1914,I2583,I1902,I2945,I2798,I1899,I2962,I2832,I2651,I2203,I2815,I1917,I1937,I2457;
nand I_0(I2668,I2651,I1914);
DFFARX1 I_1(I2457,I1294,I1937,,,I1914,);
not I_2(I2583,I1301);
and I_3(I1902,I2234,I2203);
DFFARX1 I_4(I1902,I1294,I2583,,,I2945,);
and I_5(I2798,I2781,I1899);
DFFARX1 I_6(I1294,I1937,,,I1899,);
nor I_7(I2962,I2945,I2668);
DFFARX1 I_8(I2815,I1294,I2583,,,I2832,);
nor I_9(I2651,I2600,I1908);
DFFARX1 I_10(I1294,I1937,,,I2203,);
or I_11(I2815,I2798,I1917);
nand I_12(I1917,I2406,I2505);
not I_13(I1937,I1301);
nand I_14(I2569,I2832,I2962);
or I_15(I2457,I2234);
endmodule


