module test_final(IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,IN_1_3_l_7,IN_2_3_l_7,IN_3_3_l_7,IN_1_4_l_7,IN_2_4_l_7,IN_3_4_l_7,IN_4_4_l_7,IN_5_4_l_7,blif_clk_net_5_r_3,blif_reset_net_5_r_3,N1371_0_r_3,N1508_0_r_3,N6147_3_r_3,n_429_or_0_5_r_3,G78_5_r_3,n_576_5_r_3,n_102_5_r_3,n_547_5_r_3,N1508_10_r_3);
input IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,IN_1_3_l_7,IN_2_3_l_7,IN_3_3_l_7,IN_1_4_l_7,IN_2_4_l_7,IN_3_4_l_7,IN_4_4_l_7,IN_5_4_l_7,blif_clk_net_5_r_3,blif_reset_net_5_r_3;
output N1371_0_r_3,N1508_0_r_3,N6147_3_r_3,n_429_or_0_5_r_3,G78_5_r_3,n_576_5_r_3,n_102_5_r_3,n_547_5_r_3,N1508_10_r_3;
wire N1371_0_r_7,N1508_0_r_7,N6147_2_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_102_5_r_7,n_547_5_r_7,N1507_6_r_7,N1508_6_r_7,n_431_5_r_7,n19_7,n20_7,n21_7,n22_7,n23_7,n24_7,n25_7,n26_7,n27_7,n28_7,n29_7,n30_7,n31_7,n32_7,N1372_10_r_3,N3_8_l_3,n5_3,n39_3,n_431_5_r_3,n22_3,n23_3,n24_3,n25_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3;
nor I_0(N1371_0_r_7,n22_7,n24_7);
nor I_1(N1508_0_r_7,n24_7,n28_7);
nor I_2(N6147_2_r_7,n21_7,n26_7);
nand I_3(n_429_or_0_5_r_7,n19_7,n24_7);
DFFARX1 I_4(n_431_5_r_7,blif_clk_net_5_r_3,n5_3,G78_5_r_7,);
nand I_5(n_576_5_r_7,N1371_0_r_7,n19_7);
not I_6(n_102_5_r_7,n22_7);
nand I_7(n_547_5_r_7,n20_7,n21_7);
nor I_8(N1507_6_r_7,n22_7,n27_7);
nor I_9(N1508_6_r_7,IN_3_1_l_7,n27_7);
nand I_10(n_431_5_r_7,n24_7,n25_7);
nor I_11(n19_7,IN_1_3_l_7,n30_7);
nor I_12(n20_7,n22_7,n23_7);
not I_13(n21_7,n29_7);
nor I_14(n22_7,n29_7,n31_7);
not I_15(n23_7,n27_7);
not I_16(n24_7,N1508_6_r_7);
nand I_17(n25_7,N1507_6_r_7,n19_7);
or I_18(n26_7,n19_7,n23_7);
nand I_19(n27_7,IN_1_1_l_7,IN_2_1_l_7);
nor I_20(n28_7,n19_7,n21_7);
nand I_21(n29_7,IN_1_4_l_7,IN_2_4_l_7);
or I_22(n30_7,IN_2_3_l_7,IN_3_3_l_7);
nor I_23(n31_7,IN_5_4_l_7,n32_7);
and I_24(n32_7,IN_3_4_l_7,IN_4_4_l_7);
nor I_25(N1371_0_r_3,n39_3,n37_3);
nor I_26(N1508_0_r_3,n25_3,n37_3);
nor I_27(N6147_3_r_3,N1372_10_r_3,n33_3);
nand I_28(n_429_or_0_5_r_3,N1372_10_r_3,n30_3);
DFFARX1 I_29(n_431_5_r_3,blif_clk_net_5_r_3,n5_3,G78_5_r_3,);
nand I_30(n_576_5_r_3,n22_3,n23_3);
not I_31(n_102_5_r_3,n39_3);
nand I_32(n_547_5_r_3,n26_3,n27_3);
not I_33(N1372_10_r_3,n36_3);
nor I_34(N1508_10_r_3,n35_3,n36_3);
and I_35(N3_8_l_3,n34_3,N1508_0_r_7);
not I_36(n5_3,blif_reset_net_5_r_3);
DFFARX1 I_37(N3_8_l_3,blif_clk_net_5_r_3,n5_3,n39_3,);
nand I_38(n_431_5_r_3,n29_3,n30_3);
nor I_39(n22_3,n24_3,n25_3);
nor I_40(n23_3,n39_3,n_429_or_0_5_r_7);
not I_41(n24_3,n27_3);
nand I_42(n25_3,G78_5_r_7,n_576_5_r_7);
nor I_43(n26_3,n39_3,n28_3);
nor I_44(n27_3,N1508_0_r_7,N6147_2_r_7);
not I_45(n28_3,n37_3);
nand I_46(n29_3,N1372_10_r_3,n39_3);
nand I_47(n30_3,n31_3,n32_3);
not I_48(n31_3,n25_3);
not I_49(n32_3,n_429_or_0_5_r_7);
nand I_50(n33_3,n24_3,n25_3);
nand I_51(n34_3,N1508_0_r_7,G78_5_r_7);
nor I_52(n35_3,n27_3,n31_3);
nand I_53(n36_3,n28_3,n38_3);
nand I_54(n37_3,n_102_5_r_7,n_547_5_r_7);
or I_55(n38_3,N6147_2_r_7,n_429_or_0_5_r_7);
endmodule


