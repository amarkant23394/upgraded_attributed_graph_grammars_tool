module test_I2313(I1223,I1255,I1294,I1239,I1207,I1301,I2313);
input I1223,I1255,I1294,I1239,I1207,I1301;
output I2313;
wire I1410,I1622,I1937,I1342,I1331,I1639;
nor I_0(I1410,I1223,I1239);
DFFARX1 I_1(I1255,I1294,I1342,,,I1622,);
DFFARX1 I_2(I1331,I1294,I1937,,,I2313,);
not I_3(I1937,I1301);
not I_4(I1342,I1301);
nor I_5(I1331,I1639,I1410);
and I_6(I1639,I1622,I1207);
endmodule


