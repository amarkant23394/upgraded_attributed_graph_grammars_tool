module test_I10879(I8496,I9459,I8193,I9491,I8360,I8267,I1470,I10879);
input I8496,I9459,I8193,I9491,I8360,I8267,I1470;
output I10879;
wire I8202,I9720,I10845,I9542,I10862,I9816,I9453,I8181,I8592,I10828,I9462,I9576,I9483,I9689;
or I_0(I10879,I10862,I9462);
nand I_1(I8202,I8267,I8496);
not I_2(I9720,I9689);
nor I_3(I10845,I10828,I9483);
DFFARX1 I_4(I1470,I9491,,,I9542,);
and I_5(I10862,I10845,I9453);
DFFARX1 I_6(I8193,I1470,I9491,,,I9816,);
nand I_7(I9453,I9816,I9720);
and I_8(I8181,I8360,I8592);
DFFARX1 I_9(I1470,,,I8592,);
not I_10(I10828,I9459);
not I_11(I9462,I9576);
nor I_12(I9576,I8181,I8202);
nor I_13(I9483,I9816,I9542);
DFFARX1 I_14(I1470,I9491,,,I9689,);
endmodule


