module test_I4595(I1477,I2557,I2294,I1470,I1375,I4595);
input I1477,I2557,I2294,I1470,I1375;
output I4595;
wire I2173,I2181,I4544,I4561,I2458,I2509,I2152,I2345,I4578,I2311,I2161;
nand I_0(I2173,I2557,I2509);
not I_1(I2181,I1477);
DFFARX1 I_2(I4578,I1470,I4544,,,I4595,);
not I_3(I4544,I1477);
nand I_4(I4561,I2152,I2173);
DFFARX1 I_5(I1470,I2181,,,I2458,);
nor I_6(I2509,I2458);
DFFARX1 I_7(I2458,I1470,I2181,,,I2152,);
DFFARX1 I_8(I1375,I1470,I2181,,,I2345,);
and I_9(I4578,I4561,I2161);
not I_10(I2311,I2294);
nand I_11(I2161,I2345,I2311);
endmodule


