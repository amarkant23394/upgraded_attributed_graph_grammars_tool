module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_7_r_16,blif_reset_net_7_r_16,N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_7_r_16,blif_reset_net_7_r_16;
output N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,n_549_7_r_16,N3_8_l_16,n8_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_7_r_16,n8_16,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
nor I_35(N1371_0_r_16,n35_16,n39_16);
nor I_36(N1508_0_r_16,n39_16,n46_16);
not I_37(N1372_1_r_16,n45_16);
nor I_38(N1508_1_r_16,n53_16,n45_16);
nor I_39(N6147_2_r_16,n37_16,n38_16);
nor I_40(N1507_6_r_16,n44_16,n49_16);
nor I_41(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_42(n4_7_r_16,blif_clk_net_7_r_16,n8_16,G42_7_r_16,);
nor I_43(n_572_7_r_16,n32_16,n33_16);
nand I_44(n_573_7_r_16,n30_16,n31_16);
nand I_45(n_549_7_r_16,n47_16,N1371_0_r_4);
nand I_46(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_47(n_452_7_r_16,n34_16,n35_16);
and I_48(N3_8_l_16,n41_16,N1508_6_r_4);
not I_49(n8_16,blif_reset_net_7_r_16);
DFFARX1 I_50(N3_8_l_16,blif_clk_net_7_r_16,n8_16,n53_16,);
not I_51(n29_16,n53_16);
nor I_52(n4_7_r_16,n35_16,n36_16);
nand I_53(n30_16,n_549_7_r_4,N1371_0_r_4);
not I_54(n31_16,n34_16);
nor I_55(n32_16,n30_16,n_572_7_r_4);
not I_56(n33_16,n_549_7_r_16);
nor I_57(n34_16,n48_16,N1507_6_r_4);
and I_58(n35_16,n50_16,n_452_7_r_4);
not I_59(n36_16,n30_16);
nor I_60(n37_16,n31_16,n40_16);
nand I_61(n38_16,n29_16,n39_16);
not I_62(n39_16,n32_16);
nor I_63(n40_16,N1507_6_r_4,G42_7_r_4);
nand I_64(n41_16,N1507_6_r_4,n_549_7_r_4);
nand I_65(n42_16,n35_16,n43_16);
not I_66(n43_16,n44_16);
nor I_67(n44_16,n32_16,n49_16);
nand I_68(n45_16,n36_16,n40_16);
nor I_69(n46_16,n33_16,n34_16);
nand I_70(n47_16,n_569_7_r_4,n_572_7_r_4);
or I_71(n48_16,N1508_6_r_4,N6134_9_r_4);
and I_72(n49_16,n35_16,n36_16);
and I_73(n50_16,n51_16,G42_7_r_4);
nand I_74(n51_16,n47_16,n52_16);
not I_75(n52_16,N1371_0_r_4);
endmodule


