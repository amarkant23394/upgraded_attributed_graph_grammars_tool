module test_I2424(I1255,I1223,I2424);
input I1255,I1223;
output I2424;
wire ;
nand I_0(I2424,I1223,I1255);
endmodule


