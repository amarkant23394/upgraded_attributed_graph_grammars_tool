module test_I13987(I12270,I12476,I1477,I1470,I12174,I13987);
input I12270,I12476,I1477,I1470,I12174;
output I13987;
wire I11935,I11950,I12208,I10023,I12493,I11973,I13970,I12191,I11941;
DFFARX1 I_0(I12208,I1470,I11973,,,I11935,);
DFFARX1 I_1(I12493,I1470,I11973,,,I11950,);
DFFARX1 I_2(I12191,I1470,I11973,,,I12208,);
DFFARX1 I_3(I1470,,,I10023,);
or I_4(I12493,I12270,I12476);
and I_5(I13987,I13970,I11941);
not I_6(I11973,I1477);
nand I_7(I13970,I11935,I11950);
or I_8(I12191,I12174,I10023);
DFFARX1 I_9(I12208,I1470,I11973,,,I11941,);
endmodule


