module test_final(G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_10,blif_reset_net_1_r_10,G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10);
input G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_10,blif_reset_net_1_r_10;
output G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10;
wire G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,n_452_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15,n4_1_l_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15,n_452_1_r_10,N3_2_l_10,n4_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10;
DFFARX1 I_0(n_452_1_r_15,blif_clk_net_1_r_10,n4_10,G42_1_r_15,);
and I_1(n_572_1_r_15,n17_15,n19_15);
nand I_2(n_573_1_r_15,n15_15,n18_15);
nor I_3(n_549_1_r_15,n21_15,n22_15);
nand I_4(n_569_1_r_15,n15_15,n20_15);
nor I_5(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_6(G42_1_l_15,blif_clk_net_1_r_10,n4_10,ACVQN2_3_r_15,);
nor I_7(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_8(N1_4_r_15,blif_clk_net_1_r_10,n4_10,G199_4_r_15,);
DFFARX1 I_9(n_573_1_l_15,blif_clk_net_1_r_10,n4_10,G214_4_r_15,);
nor I_10(n4_1_l_15,G18_1_l_15,IN_1_1_l_15);
DFFARX1 I_11(n4_1_l_15,blif_clk_net_1_r_10,n4_10,G42_1_l_15,);
not I_12(n15_15,G42_1_l_15);
DFFARX1 I_13(IN_1_3_l_15,blif_clk_net_1_r_10,n4_10,n17_internal_15,);
not I_14(n17_15,n17_internal_15);
DFFARX1 I_15(IN_2_3_l_15,blif_clk_net_1_r_10,n4_10,n30_15,);
nor I_16(n_572_1_l_15,G15_1_l_15,IN_7_1_l_15);
DFFARX1 I_17(n_572_1_l_15,blif_clk_net_1_r_10,n4_10,n14_internal_15,);
not I_18(n14_15,n14_internal_15);
nand I_19(N1_4_r_15,n25_15,n26_15);
or I_20(n_573_1_l_15,IN_5_1_l_15,IN_9_1_l_15);
nor I_21(n18_15,IN_9_1_l_15,IN_10_1_l_15);
nand I_22(n19_15,n27_15,n28_15);
nand I_23(n20_15,IN_4_3_l_15,n30_15);
not I_24(n21_15,n20_15);
and I_25(n22_15,n17_15,n_572_1_l_15);
nor I_26(n23_15,G18_1_l_15,IN_5_1_l_15);
or I_27(n24_15,IN_9_1_l_15,IN_10_1_l_15);
or I_28(n25_15,G18_1_l_15,n_573_1_l_15);
nand I_29(n26_15,n19_15,n23_15);
not I_30(n27_15,IN_10_1_l_15);
nand I_31(n28_15,IN_4_1_l_15,n29_15);
not I_32(n29_15,G15_1_l_15);
DFFARX1 I_33(n4_1_r_10,blif_clk_net_1_r_10,n4_10,G42_1_r_10,);
nor I_34(n_572_1_r_10,n26_10,n3_10);
nand I_35(n_573_1_r_10,n16_10,n18_10);
nand I_36(n_549_1_r_10,n19_10,n20_10);
nor I_37(n_452_1_r_10,n25_10,n21_10);
nor I_38(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_39(N3_2_r_10,blif_clk_net_1_r_10,n4_10,G199_2_r_10,);
DFFARX1 I_40(G199_4_l_10,blif_clk_net_1_r_10,n4_10,ACVQN2_3_r_10,);
nor I_41(n_266_and_0_3_r_10,n17_10,n13_10);
and I_42(N3_2_l_10,n23_10,G42_1_r_15);
not I_43(n4_10,blif_reset_net_1_r_10);
DFFARX1 I_44(N3_2_l_10,blif_clk_net_1_r_10,n4_10,n25_10,);
not I_45(n16_10,n25_10);
DFFARX1 I_46(G199_4_r_15,blif_clk_net_1_r_10,n4_10,n26_10,);
DFFARX1 I_47(G214_4_r_15,blif_clk_net_1_r_10,n4_10,ACVQN1_3_l_10,);
and I_48(N1_4_l_10,n24_10,ACVQN2_3_r_15);
DFFARX1 I_49(N1_4_l_10,blif_clk_net_1_r_10,n4_10,G199_4_l_10,);
DFFARX1 I_50(n_266_and_0_3_r_15,blif_clk_net_1_r_10,n4_10,n27_10,);
not I_51(n17_10,n27_10);
nor I_52(n4_1_r_10,n27_10,n21_10);
nor I_53(N3_2_r_10,n16_10,n22_10);
not I_54(n3_10,n18_10);
DFFARX1 I_55(n3_10,blif_clk_net_1_r_10,n4_10,n13_internal_10,);
not I_56(n13_10,n13_internal_10);
nand I_57(n18_10,ACVQN1_3_l_10,n_549_1_r_15);
not I_58(n19_10,n_452_1_r_10);
nand I_59(n20_10,n16_10,n26_10);
nor I_60(n21_10,n_573_1_r_15,n_572_1_r_15);
and I_61(n22_10,n26_10,n21_10);
nand I_62(n23_10,n_573_1_r_15,n_569_1_r_15);
nand I_63(n24_10,G42_1_r_15,n_572_1_r_15);
endmodule


