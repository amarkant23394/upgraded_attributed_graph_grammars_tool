module test_I8930(I7122,I5085,I1477,I5097,I6975,I7057,I1470,I8930);
input I7122,I5085,I1477,I5097,I6975,I7057,I1470;
output I8930;
wire I6893,I7317,I5067,I6907,I6887,I7139,I7410,I7269,I6992,I7286,I7156,I7427,I8879;
nand I_0(I6893,I7156,I7286);
nor I_1(I7317,I7269,I7057);
DFFARX1 I_2(I1470,,,I5067,);
not I_3(I6907,I1477);
nand I_4(I6887,I7427,I7317);
or I_5(I7139,I7122,I5085);
nor I_6(I8930,I8879,I6893);
DFFARX1 I_7(I1470,I6907,,,I7410,);
DFFARX1 I_8(I5067,I1470,I6907,,,I7269,);
nand I_9(I6992,I6975,I5097);
nor I_10(I7286,I7269,I6992);
DFFARX1 I_11(I7139,I1470,I6907,,,I7156,);
not I_12(I7427,I7410);
not I_13(I8879,I6887);
endmodule


