module test_final(G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_1,blif_reset_net_1_r_1,G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1);
input G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_1,blif_reset_net_1_r_1;
output G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1;
wire G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_452_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14,n4_1_l_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14,N3_2_l_1,n5_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1;
DFFARX1 I_0(n_452_1_r_14,blif_clk_net_1_r_1,n5_1,G42_1_r_14,);
and I_1(n_572_1_r_14,n18_14,n19_14);
nand I_2(n_573_1_r_14,n16_14,n17_14);
nor I_3(n_549_1_r_14,n20_14,n21_14);
or I_4(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_5(n_452_1_r_14,IN_10_1_l_14,n23_14);
nor I_6(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_7(N3_2_r_14,blif_clk_net_1_r_1,n5_1,G199_2_r_14,);
DFFARX1 I_8(n_572_1_l_14,blif_clk_net_1_r_1,n5_1,ACVQN1_5_r_14,);
not I_9(P6_5_r_14,P6_5_r_internal_14);
nor I_10(n4_1_l_14,G18_1_l_14,IN_1_1_l_14);
DFFARX1 I_11(n4_1_l_14,blif_clk_net_1_r_1,n5_1,n15_internal_14,);
not I_12(n15_14,n15_internal_14);
DFFARX1 I_13(IN_1_3_l_14,blif_clk_net_1_r_1,n5_1,ACVQN2_3_l_14,);
DFFARX1 I_14(IN_2_3_l_14,blif_clk_net_1_r_1,n5_1,ACVQN1_3_l_14,);
and I_15(N3_2_r_14,n26_14,n27_14);
nor I_16(n_572_1_l_14,G15_1_l_14,IN_7_1_l_14);
DFFARX1 I_17(ACVQN2_3_l_14,blif_clk_net_1_r_1,n5_1,P6_5_r_internal_14,);
nor I_18(n16_14,IN_9_1_l_14,IN_10_1_l_14);
not I_19(n17_14,n_572_1_l_14);
nor I_20(n18_14,IN_5_1_l_14,IN_9_1_l_14);
nand I_21(n19_14,IN_4_3_l_14,ACVQN1_3_l_14);
nor I_22(n20_14,G18_1_l_14,IN_5_1_l_14);
nor I_23(n21_14,n15_14,n22_14);
nand I_24(n22_14,n24_14,n25_14);
nand I_25(n23_14,n15_14,n24_14);
not I_26(n24_14,IN_9_1_l_14);
not I_27(n25_14,IN_5_1_l_14);
nor I_28(n26_14,IN_10_1_l_14,n20_14);
nand I_29(n27_14,IN_4_1_l_14,n28_14);
not I_30(n28_14,G15_1_l_14);
DFFARX1 I_31(n4_1_r_1,blif_clk_net_1_r_1,n5_1,G42_1_r_1,);
nor I_32(n_572_1_r_1,n26_1,n19_1);
nand I_33(n_573_1_r_1,n16_1,n18_1);
nor I_34(n_549_1_r_1,n20_1,n21_1);
nor I_35(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_36(G199_4_l_1,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_1,);
nor I_37(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_38(N1_4_r_1,blif_clk_net_1_r_1,n5_1,G199_4_r_1,);
DFFARX1 I_39(G199_4_l_1,blif_clk_net_1_r_1,n5_1,G214_4_r_1,);
and I_40(N3_2_l_1,n23_1,P6_5_r_14);
not I_41(n5_1,blif_reset_net_1_r_1);
DFFARX1 I_42(N3_2_l_1,blif_clk_net_1_r_1,n5_1,n26_1,);
not I_43(n17_1,n26_1);
DFFARX1 I_44(G42_1_r_14,blif_clk_net_1_r_1,n5_1,n16_internal_1,);
not I_45(n16_1,n16_internal_1);
DFFARX1 I_46(n_573_1_r_14,blif_clk_net_1_r_1,n5_1,ACVQN1_3_l_1,);
and I_47(N1_4_l_1,n25_1,n_549_1_r_14);
DFFARX1 I_48(N1_4_l_1,blif_clk_net_1_r_1,n5_1,G199_4_l_1,);
DFFARX1 I_49(n_42_2_r_14,blif_clk_net_1_r_1,n5_1,G214_4_l_1,);
nor I_50(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_51(G214_4_l_1,blif_clk_net_1_r_1,n5_1,n14_internal_1,);
not I_52(n14_1,n14_internal_1);
nor I_53(N1_4_r_1,n17_1,n24_1);
nand I_54(n18_1,ACVQN1_3_l_1,n_569_1_r_14);
nor I_55(n19_1,G199_2_r_14,G42_1_r_14);
not I_56(n20_1,n18_1);
nor I_57(n21_1,n26_1,n22_1);
not I_58(n22_1,n19_1);
nand I_59(n23_1,n_572_1_r_14,G42_1_r_14);
nor I_60(n24_1,n18_1,n22_1);
nand I_61(n25_1,ACVQN1_5_r_14,n_572_1_r_14);
endmodule


