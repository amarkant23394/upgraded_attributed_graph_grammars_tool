module test_I10618(I9462,I10862,I1470_clk,I1477_rst,I10618);
input I9462,I10862,I1470_clk,I1477_rst;
output I10618;
wire I10930,I10879,I10647,I10896;
DFFARX1 I_0 (I10896,I10647,I1470_clk,);
or I_1(I10879,I10862,I9462);
not I_2(I10647,I1477_rst);
not I_3(I10618,I10930);
DFFARX1 I_4 (I10879,I10647,I1470_clk,);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule