module test_I7714(I3966,I1477,I6442,I1470,I7714);
input I3966,I1477,I6442,I1470;
output I7714;
wire I6781,I6297,I6826,I6329,I6493,I6843;
DFFARX1 I_0(I1470,I6329,,,I6781,);
DFFARX1 I_1(I6843,I1470,I6329,,,I6297,);
not I_2(I7714,I6297);
nand I_3(I6826,I6781,I6442);
not I_4(I6329,I1477);
DFFARX1 I_5(I3966,I1470,I6329,,,I6493,);
and I_6(I6843,I6493,I6826);
endmodule


