module test_final(G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_1,blif_reset_net_1_r_1,G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1);
input G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_1,blif_reset_net_1_r_1;
output G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1;
wire G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,n_452_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15,n4_1_l_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15,N3_2_l_1,n5_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1;
DFFARX1 I_0(n_452_1_r_15,blif_clk_net_1_r_1,n5_1,G42_1_r_15,);
and I_1(n_572_1_r_15,n17_15,n19_15);
nand I_2(n_573_1_r_15,n15_15,n18_15);
nor I_3(n_549_1_r_15,n21_15,n22_15);
nand I_4(n_569_1_r_15,n15_15,n20_15);
nor I_5(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_6(G42_1_l_15,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_15,);
nor I_7(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_8(N1_4_r_15,blif_clk_net_1_r_1,n5_1,G199_4_r_15,);
DFFARX1 I_9(n_573_1_l_15,blif_clk_net_1_r_1,n5_1,G214_4_r_15,);
nor I_10(n4_1_l_15,G18_1_l_15,IN_1_1_l_15);
DFFARX1 I_11(n4_1_l_15,blif_clk_net_1_r_1,n5_1,G42_1_l_15,);
not I_12(n15_15,G42_1_l_15);
DFFARX1 I_13(IN_1_3_l_15,blif_clk_net_1_r_1,n5_1,n17_internal_15,);
not I_14(n17_15,n17_internal_15);
DFFARX1 I_15(IN_2_3_l_15,blif_clk_net_1_r_1,n5_1,n30_15,);
nor I_16(n_572_1_l_15,G15_1_l_15,IN_7_1_l_15);
DFFARX1 I_17(n_572_1_l_15,blif_clk_net_1_r_1,n5_1,n14_internal_15,);
not I_18(n14_15,n14_internal_15);
nand I_19(N1_4_r_15,n25_15,n26_15);
or I_20(n_573_1_l_15,IN_5_1_l_15,IN_9_1_l_15);
nor I_21(n18_15,IN_9_1_l_15,IN_10_1_l_15);
nand I_22(n19_15,n27_15,n28_15);
nand I_23(n20_15,IN_4_3_l_15,n30_15);
not I_24(n21_15,n20_15);
and I_25(n22_15,n17_15,n_572_1_l_15);
nor I_26(n23_15,G18_1_l_15,IN_5_1_l_15);
or I_27(n24_15,IN_9_1_l_15,IN_10_1_l_15);
or I_28(n25_15,G18_1_l_15,n_573_1_l_15);
nand I_29(n26_15,n19_15,n23_15);
not I_30(n27_15,IN_10_1_l_15);
nand I_31(n28_15,IN_4_1_l_15,n29_15);
not I_32(n29_15,G15_1_l_15);
DFFARX1 I_33(n4_1_r_1,blif_clk_net_1_r_1,n5_1,G42_1_r_1,);
nor I_34(n_572_1_r_1,n26_1,n19_1);
nand I_35(n_573_1_r_1,n16_1,n18_1);
nor I_36(n_549_1_r_1,n20_1,n21_1);
nor I_37(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_38(G199_4_l_1,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_1,);
nor I_39(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_40(N1_4_r_1,blif_clk_net_1_r_1,n5_1,G199_4_r_1,);
DFFARX1 I_41(G199_4_l_1,blif_clk_net_1_r_1,n5_1,G214_4_r_1,);
and I_42(N3_2_l_1,n23_1,n_266_and_0_3_r_15);
not I_43(n5_1,blif_reset_net_1_r_1);
DFFARX1 I_44(N3_2_l_1,blif_clk_net_1_r_1,n5_1,n26_1,);
not I_45(n17_1,n26_1);
DFFARX1 I_46(ACVQN2_3_r_15,blif_clk_net_1_r_1,n5_1,n16_internal_1,);
not I_47(n16_1,n16_internal_1);
DFFARX1 I_48(G199_4_r_15,blif_clk_net_1_r_1,n5_1,ACVQN1_3_l_1,);
and I_49(N1_4_l_1,n25_1,n_573_1_r_15);
DFFARX1 I_50(N1_4_l_1,blif_clk_net_1_r_1,n5_1,G199_4_l_1,);
DFFARX1 I_51(n_549_1_r_15,blif_clk_net_1_r_1,n5_1,G214_4_l_1,);
nor I_52(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_53(G214_4_l_1,blif_clk_net_1_r_1,n5_1,n14_internal_1,);
not I_54(n14_1,n14_internal_1);
nor I_55(N1_4_r_1,n17_1,n24_1);
nand I_56(n18_1,ACVQN1_3_l_1,G214_4_r_15);
nor I_57(n19_1,n_569_1_r_15,G42_1_r_15);
not I_58(n20_1,n18_1);
nor I_59(n21_1,n26_1,n22_1);
not I_60(n22_1,n19_1);
nand I_61(n23_1,n_572_1_r_15,n_569_1_r_15);
nor I_62(n24_1,n18_1,n22_1);
nand I_63(n25_1,G42_1_r_15,n_572_1_r_15);
endmodule


