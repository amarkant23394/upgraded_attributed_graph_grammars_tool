module test_final(IN_1_0_l,IN_2_0_l,IN_3_0_l,IN_4_0_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,IN_1_8_l,IN_2_8_l,IN_3_8_l,IN_6_8_l,IN_1_10_l,IN_2_10_l,IN_3_10_l,IN_4_10_l,blif_clk_net_5_r,blif_reset_net_5_r,N1372_1_r,N1508_1_r,N6147_2_r,N6147_3_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,N1507_6_r,N1508_6_r,N1372_10_r,N1508_10_r);
input IN_1_0_l,IN_2_0_l,IN_3_0_l,IN_4_0_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,IN_1_8_l,IN_2_8_l,IN_3_8_l,IN_6_8_l,IN_1_10_l,IN_2_10_l,IN_3_10_l,IN_4_10_l,blif_clk_net_5_r,blif_reset_net_5_r;
output N1372_1_r,N1508_1_r,N6147_2_r,N6147_3_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,N1507_6_r,N1508_6_r,N1372_10_r,N1508_10_r;
wire N1371_0_l,N1508_0_l,n3_0_l,n4_0_l,N6147_3_l,n3_3_l,N6138_3_l,n_42_8_l,G199_8_l,N3_8_l,n3_8_l,N1372_10_l,N1508_10_l,n5_10_l,n6_10_l,n4_1_r,n5_2_r,n6_2_r,N6138_2_r,n7_2_r,n3_3_r,N6138_3_r,n_431_5_r,n2_5_r,n11_5_r,n12_5_r,n13_5_r,n14_5_r,n15_5_r,n16_5_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,n5_10_r,n6_10_r;
nor I_0(N1371_0_l,IN_2_0_l,n4_0_l);
nor I_1(N1508_0_l,n3_0_l,n4_0_l);
nor I_2(n3_0_l,IN_3_0_l,IN_4_0_l);
not I_3(n4_0_l,IN_1_0_l);
nor I_4(N6147_3_l,IN_3_3_l,n3_3_l);
not I_5(n3_3_l,N6138_3_l);
nor I_6(N6138_3_l,IN_1_3_l,IN_2_3_l);
nor I_7(n_42_8_l,IN_1_8_l,IN_3_8_l);
DFFARX1 I_8(N3_8_l,blif_clk_net_5_r,n2_5_r,G199_8_l,);
and I_9(N3_8_l,IN_6_8_l,n3_8_l);
nand I_10(n3_8_l,IN_2_8_l,IN_3_8_l);
not I_11(N1372_10_l,n6_10_l);
nor I_12(N1508_10_l,n5_10_l,n6_10_l);
nor I_13(n5_10_l,IN_3_10_l,IN_4_10_l);
nand I_14(n6_10_l,IN_1_10_l,IN_2_10_l);
not I_15(N1372_1_r,n4_1_r);
nor I_16(N1508_1_r,n4_1_r,N1372_10_l);
nand I_17(n4_1_r,N1508_0_l,n_42_8_l);
nor I_18(N6147_2_r,n5_2_r,n6_2_r);
nor I_19(n5_2_r,n7_2_r,N1372_10_l);
not I_20(n6_2_r,N6138_2_r);
nor I_21(N6138_2_r,n_42_8_l,N6147_3_l);
nor I_22(n7_2_r,N1508_0_l,N6147_3_l);
nor I_23(N6147_3_r,n3_3_r,N1508_10_l);
not I_24(n3_3_r,N6138_3_r);
nor I_25(N6138_3_r,N1508_0_l,N1371_0_l);
nand I_26(n_429_or_0_5_r,n12_5_r,n_42_8_l);
DFFARX1 I_27(n_431_5_r,blif_clk_net_5_r,n2_5_r,G78_5_r,);
nand I_28(n_576_5_r,n11_5_r,G199_8_l);
not I_29(n_102_5_r,N1508_0_l);
nand I_30(n_547_5_r,n13_5_r,N1371_0_l);
or I_31(n_431_5_r,n14_5_r,N1508_10_l);
not I_32(n2_5_r,blif_reset_net_5_r);
nor I_33(n11_5_r,n12_5_r,N1508_0_l);
not I_34(n12_5_r,N1372_10_l);
nor I_35(n13_5_r,N1508_0_l,G199_8_l);
and I_36(n14_5_r,n15_5_r,N1371_0_l);
nor I_37(n15_5_r,n16_5_r,N1371_0_l);
not I_38(n16_5_r,n_42_8_l);
nor I_39(N1507_6_r,n8_6_r,n9_6_r);
and I_40(N1508_6_r,n6_6_r,N6147_3_l);
nor I_41(n6_6_r,n7_6_r,n8_6_r);
not I_42(n7_6_r,N1371_0_l);
nor I_43(n8_6_r,n9_6_r,G199_8_l);
and I_44(n9_6_r,N1372_10_l,N1508_10_l);
not I_45(N1372_10_r,n6_10_r);
nor I_46(N1508_10_r,n5_10_r,n6_10_r);
nor I_47(n5_10_r,G199_8_l,N1508_10_l);
nand I_48(n6_10_r,N6147_3_l,n_42_8_l);
endmodule


