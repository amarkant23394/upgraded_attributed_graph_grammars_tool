module test_I8202(I8428,I1477,I5728,I4518,I5881,I6265,I1470,I8202);
input I8428,I1477,I5728,I4518,I5881,I6265,I1470;
output I8202;
wire I5963,I8496,I5898,I5802,I5716,I8216,I5719,I8377,I8250,I5737,I8360,I6203,I5751,I8445,I8462,I8267;
nand I_0(I8202,I8267,I8496);
DFFARX1 I_1(I1470,I5751,,,I5963,);
nor I_2(I8496,I8462,I8377);
nor I_3(I5898,I5802,I5881);
DFFARX1 I_4(I1470,I5751,,,I5802,);
and I_5(I5716,I5802,I5963);
not I_6(I8216,I1477);
DFFARX1 I_7(I6265,I1470,I5751,,,I5719,);
not I_8(I8377,I8360);
nor I_9(I8250,I5719,I5716);
nand I_10(I5737,I6203,I5898);
not I_11(I8360,I5719);
DFFARX1 I_12(I4518,I1470,I5751,,,I6203,);
not I_13(I5751,I1477);
or I_14(I8445,I8428,I5728);
DFFARX1 I_15(I8445,I1470,I8216,,,I8462,);
nand I_16(I8267,I8250,I5737);
endmodule


