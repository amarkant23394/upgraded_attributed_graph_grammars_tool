module test_final(G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_7,blif_reset_net_1_r_7,G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7);
input G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_7,blif_reset_net_1_r_7;
output G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7;
wire G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4,n_431_0_l_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n_431_0_l_7,n8_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7;
DFFARX1 I_0(n4_1_r_4,blif_clk_net_1_r_7,n8_7,G42_1_r_4,);
nor I_1(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_2(n_573_1_r_4,G2_0_l_4,n16_4);
nor I_3(n_549_1_r_4,n22_4,n23_4);
nand I_4(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_5(n19_4,blif_clk_net_1_r_7,n8_7,ACVQN2_3_r_4,);
nor I_6(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_7(n19_4,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_4,);
not I_8(P6_5_r_4,P6_5_r_internal_4);
or I_9(n_431_0_l_4,IN_8_0_l_4,n26_4);
DFFARX1 I_10(n_431_0_l_4,blif_clk_net_1_r_7,n8_7,G78_0_l_4,);
DFFARX1 I_11(IN_2_5_l_4,blif_clk_net_1_r_7,n8_7,ACVQN1_5_l_4,);
not I_12(n16_4,ACVQN1_5_l_4);
DFFARX1 I_13(IN_1_5_l_4,blif_clk_net_1_r_7,n8_7,n17_internal_4,);
not I_14(n17_4,n17_internal_4);
nor I_15(n4_1_r_4,n30_4,n31_4);
nand I_16(n19_4,G1_0_l_4,n33_4);
DFFARX1 I_17(G78_0_l_4,blif_clk_net_1_r_7,n8_7,n15_internal_4,);
not I_18(n15_4,n15_internal_4);
DFFARX1 I_19(ACVQN1_5_l_4,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_4,);
and I_20(n20_4,IN_11_0_l_4,n16_4);
nor I_21(n21_4,G2_0_l_4,IN_10_0_l_4);
nand I_22(n22_4,G78_0_l_4,n25_4);
nand I_23(n23_4,IN_11_0_l_4,n24_4);
not I_24(n24_4,G2_0_l_4);
not I_25(n25_4,IN_10_0_l_4);
and I_26(n26_4,IN_2_0_l_4,n27_4);
nor I_27(n27_4,IN_4_0_l_4,n28_4);
not I_28(n28_4,G1_0_l_4);
not I_29(n29_4,n30_4);
nand I_30(n30_4,IN_7_0_l_4,n32_4);
nand I_31(n31_4,IN_11_0_l_4,n25_4);
nor I_32(n32_4,G2_0_l_4,n33_4);
not I_33(n33_4,IN_5_0_l_4);
DFFARX1 I_34(n4_1_r_7,blif_clk_net_1_r_7,n8_7,G42_1_r_7,);
nor I_35(n_572_1_r_7,n30_7,n31_7);
nand I_36(n_573_1_r_7,n28_7,n_266_and_0_3_r_4);
nor I_37(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_38(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_39(N1_4_r_7,blif_clk_net_1_r_7,n8_7,G199_4_r_7,);
DFFARX1 I_40(n26_7,blif_clk_net_1_r_7,n8_7,G214_4_r_7,);
DFFARX1 I_41(n5_7,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_7,);
not I_42(P6_5_r_7,P6_5_r_internal_7);
or I_43(n_431_0_l_7,n36_7,n_572_1_r_4);
not I_44(n8_7,blif_reset_net_1_r_7);
DFFARX1 I_45(n_431_0_l_7,blif_clk_net_1_r_7,n8_7,n43_7,);
not I_46(n27_7,n43_7);
DFFARX1 I_47(G42_1_r_4,blif_clk_net_1_r_7,n8_7,ACVQN1_5_l_7,);
DFFARX1 I_48(P6_5_r_4,blif_clk_net_1_r_7,n8_7,n44_7,);
nor I_49(n4_1_r_7,n30_7,n38_7);
nor I_50(N1_4_r_7,n27_7,n40_7);
nand I_51(n26_7,n39_7,ACVQN1_5_r_4);
not I_52(n5_7,n_549_1_r_4);
DFFARX1 I_53(ACVQN1_5_l_7,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_7,);
nor I_54(n28_7,n26_7,n29_7);
not I_55(n29_7,n_569_1_r_4);
not I_56(n30_7,ACVQN2_3_r_4);
nand I_57(n31_7,n27_7,n29_7);
nor I_58(n32_7,ACVQN1_5_l_7,n34_7);
nor I_59(n33_7,n29_7,n_549_1_r_4);
not I_60(n34_7,n_266_and_0_3_r_4);
nor I_61(n35_7,n43_7,n44_7);
and I_62(n36_7,n37_7,n_573_1_r_4);
nor I_63(n37_7,n30_7,G42_1_r_4);
nand I_64(n38_7,n29_7,n_549_1_r_4);
nor I_65(n39_7,n_549_1_r_4,n_572_1_r_4);
nor I_66(n40_7,n44_7,n41_7);
nor I_67(n41_7,n34_7,n42_7);
nand I_68(n42_7,n5_7,n_569_1_r_4);
endmodule


