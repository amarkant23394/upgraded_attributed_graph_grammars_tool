module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_8_r_10,n11_10,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_8_r_10,n11_10,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
nor I_35(N1371_0_r_10,n37_10,n38_10);
nor I_36(N1508_0_r_10,n37_10,n58_10);
nand I_37(N6147_2_r_10,n39_10,n40_10);
not I_38(N6147_3_r_10,n39_10);
nor I_39(N1372_4_r_10,n46_10,n49_10);
nor I_40(N1508_4_r_10,n51_10,n52_10);
nor I_41(N1507_6_r_10,n49_10,n60_10);
nor I_42(N1508_6_r_10,n49_10,n50_10);
nor I_43(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_44(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_45(N6147_9_r_10,n36_10,n37_10);
nor I_46(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_47(I_BUFF_1_9_r_10,n48_10);
nor I_48(N3_8_r_10,n44_10,n47_10);
not I_49(n11_10,blif_reset_net_8_r_10);
not I_50(n35_10,n49_10);
nor I_51(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_52(n37_10,n_549_7_r_0);
not I_53(n38_10,n46_10);
nand I_54(n39_10,n43_10,n44_10);
nand I_55(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_56(n41_10,n42_10,n_549_7_r_0);
not I_57(n42_10,n44_10);
nor I_58(n43_10,n45_10,n_549_7_r_0);
nand I_59(n44_10,n54_10,G78_5_r_0);
nor I_60(n45_10,n59_10,N1508_0_r_0);
nand I_61(n46_10,n61_10,G78_5_r_0);
nor I_62(n47_10,n46_10,n48_10);
nand I_63(n48_10,n62_10,n63_10);
nand I_64(n49_10,n56_10,n_429_or_0_5_r_0);
not I_65(n50_10,n45_10);
nor I_66(n51_10,n42_10,n53_10);
not I_67(n52_10,N1372_4_r_10);
nor I_68(n53_10,n48_10,n50_10);
and I_69(n54_10,n55_10,G42_7_r_0);
nand I_70(n55_10,n56_10,n57_10);
nand I_71(n56_10,N1371_0_r_0,n_429_or_0_5_r_0);
not I_72(n57_10,n_429_or_0_5_r_0);
nor I_73(n58_10,n35_10,n45_10);
nor I_74(n59_10,n_576_5_r_0,n_573_7_r_0);
nor I_75(n60_10,n37_10,n46_10);
or I_76(n61_10,n_576_5_r_0,n_573_7_r_0);
nor I_77(n62_10,n_572_7_r_0,N1508_0_r_0);
or I_78(n63_10,n64_10,n_547_5_r_0);
nor I_79(n64_10,n_569_7_r_0,N1371_0_r_0);
endmodule


