module test_I5898(I4629,I1477,I1470,I4530,I5898);
input I4629,I1477,I1470,I4530;
output I5898;
wire I5864,I5751,I5768,I4536,I4524,I4515,I4595,I4869,I5785,I5881,I4742,I5802;
nor I_0(I5864,I4536,I4515);
not I_1(I5751,I1477);
nand I_2(I5768,I4530,I4515);
nor I_3(I4536,I4869,I4595);
nor I_4(I4524,I4742,I4595);
not I_5(I4515,I4629);
DFFARX1 I_6(I1470,,,I4595,);
DFFARX1 I_7(I1470,,,I4869,);
and I_8(I5785,I5768,I4524);
not I_9(I5881,I5864);
DFFARX1 I_10(I1470,,,I4742,);
nor I_11(I5898,I5802,I5881);
DFFARX1 I_12(I5785,I1470,I5751,,,I5802,);
endmodule


