module test_I10627(I9477,I9576,I1477,I1470,I9864,I10627);
input I9477,I9576,I1477,I1470,I9864;
output I10627;
wire I10647,I9542,I9491,I10797,I11167,I11057,I9474,I9468,I10766,I11150,I11009;
not I_0(I10647,I1477);
DFFARX1 I_1(I1470,I9491,,,I9542,);
not I_2(I9491,I1477);
not I_3(I10797,I10766);
not I_4(I11167,I11150);
nor I_5(I11057,I11009,I10797);
or I_6(I9474,I9576,I9542);
nand I_7(I10627,I11167,I11057);
DFFARX1 I_8(I9864,I1470,I9491,,,I9468,);
not I_9(I10766,I9477);
DFFARX1 I_10(I9474,I1470,I10647,,,I11150,);
DFFARX1 I_11(I9468,I1470,I10647,,,I11009,);
endmodule


