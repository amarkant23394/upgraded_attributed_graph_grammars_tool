module test_final(IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_7_r_2,blif_reset_net_7_r_2,N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2);
input IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_7_r_2,blif_reset_net_7_r_2;
output N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2;
wire N1371_0_r_8,N1508_0_r_8,N1372_1_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N1508_10_r_8,N3_8_l_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8,n4_7_l_2,n10_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2;
nor I_0(N1371_0_r_8,n46_8,n51_8);
not I_1(N1508_0_r_8,n46_8);
nor I_2(N1372_1_r_8,n37_8,n49_8);
and I_3(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_4(N1507_6_r_8,n47_8,n48_8);
nor I_5(N1508_6_r_8,n37_8,n38_8);
nor I_6(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_7(N3_8_r_8,blif_clk_net_7_r_2,n10_2,G199_8_r_8,);
nor I_8(N6147_9_r_8,n29_8,n30_8);
nor I_9(N6134_9_r_8,n30_8,n31_8);
not I_10(I_BUFF_1_9_r_8,n35_8);
nor I_11(N1372_10_r_8,n46_8,n49_8);
nor I_12(N1508_10_r_8,n40_8,n41_8);
and I_13(N3_8_l_8,IN_6_8_l_8,n36_8);
DFFARX1 I_14(N3_8_l_8,blif_clk_net_7_r_2,n10_2,n53_8,);
not I_15(n29_8,n53_8);
nor I_16(N3_8_r_8,n33_8,n34_8);
and I_17(n30_8,n32_8,n33_8);
nor I_18(n31_8,IN_1_8_l_8,IN_3_8_l_8);
nand I_19(n32_8,IN_2_6_l_8,n42_8);
or I_20(n33_8,IN_3_1_l_8,n46_8);
nor I_21(n34_8,n32_8,n35_8);
nand I_22(n35_8,IN_5_6_l_8,n44_8);
nand I_23(n36_8,IN_2_8_l_8,IN_3_8_l_8);
not I_24(n37_8,n31_8);
nand I_25(n38_8,N1508_0_r_8,n39_8);
nand I_26(n39_8,n33_8,n50_8);
and I_27(n40_8,n32_8,n35_8);
not I_28(n41_8,N1372_10_r_8);
and I_29(n42_8,IN_1_6_l_8,n43_8);
nand I_30(n43_8,n44_8,n45_8);
nand I_31(n44_8,IN_3_6_l_8,IN_4_6_l_8);
not I_32(n45_8,IN_5_6_l_8);
nand I_33(n46_8,IN_1_1_l_8,IN_2_1_l_8);
not I_34(n47_8,n39_8);
nor I_35(n48_8,n35_8,n49_8);
not I_36(n49_8,n51_8);
nand I_37(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_38(n51_8,IN_1_3_l_8,n52_8);
or I_39(n52_8,IN_2_3_l_8,IN_3_3_l_8);
nor I_40(N1371_0_r_2,n32_2,n35_2);
nor I_41(N1508_0_r_2,n32_2,n55_2);
not I_42(N1372_1_r_2,n54_2);
nor I_43(N1508_1_r_2,n59_2,n54_2);
nor I_44(N6147_2_r_2,n42_2,n43_2);
nor I_45(N1507_6_r_2,n40_2,n53_2);
nor I_46(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_47(n4_7_r_2,blif_clk_net_7_r_2,n10_2,G42_7_r_2,);
nor I_48(n_572_7_r_2,n36_2,n37_2);
or I_49(n_573_7_r_2,n34_2,n35_2);
nor I_50(n_549_7_r_2,n40_2,n41_2);
nand I_51(n_569_7_r_2,n38_2,n39_2);
nor I_52(n_452_7_r_2,n59_2,n35_2);
nor I_53(n4_7_l_2,N1508_1_r_8,N6147_9_r_8);
not I_54(n10_2,blif_reset_net_7_r_2);
DFFARX1 I_55(n4_7_l_2,blif_clk_net_7_r_2,n10_2,n59_2,);
not I_56(n33_2,n59_2);
and I_57(N3_8_l_2,n49_2,N1508_6_r_8);
DFFARX1 I_58(N3_8_l_2,blif_clk_net_7_r_2,n10_2,n32_internal_2,);
not I_59(n32_2,n32_internal_2);
nor I_60(n4_7_r_2,n59_2,n36_2);
not I_61(n34_2,n39_2);
nor I_62(n35_2,n_42_8_r_8,N1507_6_r_8);
nor I_63(n36_2,N1508_1_r_8,N1508_6_r_8);
or I_64(n37_2,N1371_0_r_8,G199_8_r_8);
not I_65(n38_2,n40_2);
nand I_66(n39_2,n45_2,n57_2);
nor I_67(n40_2,n47_2,N1507_6_r_8);
nor I_68(n41_2,n32_2,n36_2);
not I_69(n42_2,n53_2);
nand I_70(n43_2,n44_2,n45_2);
nand I_71(n44_2,n38_2,n46_2);
not I_72(n45_2,N1371_0_r_8);
nand I_73(n46_2,n47_2,n48_2);
nand I_74(n47_2,N6134_9_r_8,n_42_8_r_8);
or I_75(n48_2,N1508_10_r_8,N1508_1_r_8);
nand I_76(n49_2,n_42_8_r_8,G199_8_r_8);
nand I_77(n50_2,n51_2,n52_2);
not I_78(n51_2,n47_2);
nand I_79(n52_2,n38_2,n53_2);
nor I_80(n53_2,N1508_6_r_8,G199_8_r_8);
nand I_81(n54_2,n42_2,n56_2);
nor I_82(n55_2,n34_2,n56_2);
nor I_83(n56_2,N1508_10_r_8,N1508_1_r_8);
nand I_84(n57_2,n58_2,N1371_0_r_8);
not I_85(n58_2,N1508_10_r_8);
endmodule


