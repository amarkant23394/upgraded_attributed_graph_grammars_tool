module test_final(G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_11,blif_reset_net_1_r_11,G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11);
input G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_11,blif_reset_net_1_r_11;
output G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11;
wire G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_569_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13,n4_1_l_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13,n_431_0_l_11,n9_11,n43_11,n26_11,n44_11,n45_11,n27_11,n4_1_r_11,N3_2_r_11,n24_11,n25_11,n20_internal_11,n20_11,n28_11,n29_11,n30_11,n31_11,n32_11,n33_11,n34_11,n35_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11;
DFFARX1 I_0(n4_1_r_13,blif_clk_net_1_r_11,n9_11,G42_1_r_13,);
nor I_1(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_2(n_573_1_r_13,n18_13,n19_13);
nand I_3(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_4(n_569_1_r_13,n17_13,n18_13);
nor I_5(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_6(n_266_and_0_3_l_13,blif_clk_net_1_r_11,n9_11,ACVQN2_3_r_13,);
nor I_7(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_8(n_549_1_l_13,blif_clk_net_1_r_11,n9_11,ACVQN1_5_r_13,);
not I_9(P6_5_r_13,P6_5_r_internal_13);
nor I_10(n4_1_l_13,G18_1_l_13,IN_1_1_l_13);
DFFARX1 I_11(n4_1_l_13,blif_clk_net_1_r_11,n9_11,n17_internal_13,);
not I_12(n17_13,n17_internal_13);
DFFARX1 I_13(IN_1_3_l_13,blif_clk_net_1_r_11,n9_11,n28_13,);
DFFARX1 I_14(IN_2_3_l_13,blif_clk_net_1_r_11,n9_11,ACVQN1_3_l_13,);
nor I_15(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_16(n_266_and_0_3_l_13,IN_4_3_l_13,ACVQN1_3_l_13);
nand I_17(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_18(n_573_1_l_13,blif_clk_net_1_r_11,n9_11,n14_internal_13,);
not I_19(n14_13,n14_internal_13);
and I_20(n_549_1_l_13,n21_13,n26_13);
nand I_21(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_22(n_569_1_l_13,blif_clk_net_1_r_11,n9_11,P6_5_r_internal_13,);
nand I_23(n18_13,n23_13,n24_13);
or I_24(n19_13,G15_1_l_13,IN_7_1_l_13);
not I_25(n20_13,IN_9_1_l_13);
not I_26(n21_13,IN_10_1_l_13);
nand I_27(n22_13,n17_13,n28_13);
not I_28(n23_13,G18_1_l_13);
not I_29(n24_13,IN_5_1_l_13);
nor I_30(n25_13,G15_1_l_13,IN_7_1_l_13);
nand I_31(n26_13,IN_4_1_l_13,n27_13);
not I_32(n27_13,G15_1_l_13);
DFFARX1 I_33(n4_1_r_11,blif_clk_net_1_r_11,n9_11,G42_1_r_11,);
nor I_34(n_572_1_r_11,n29_11,n30_11);
nand I_35(n_573_1_r_11,n26_11,n28_11);
nor I_36(n_549_1_r_11,n27_11,n32_11);
nand I_37(n_569_1_r_11,n45_11,n28_11);
nor I_38(n_452_1_r_11,n43_11,n44_11);
nor I_39(n_42_2_r_11,n35_11,n36_11);
DFFARX1 I_40(N3_2_r_11,blif_clk_net_1_r_11,n9_11,G199_2_r_11,);
DFFARX1 I_41(n24_11,blif_clk_net_1_r_11,n9_11,ACVQN2_3_r_11,);
nor I_42(n_266_and_0_3_r_11,n20_11,n37_11);
or I_43(n_431_0_l_11,n33_11,n_572_1_r_13);
not I_44(n9_11,blif_reset_net_1_r_11);
DFFARX1 I_45(n_431_0_l_11,blif_clk_net_1_r_11,n9_11,n43_11,);
not I_46(n26_11,n43_11);
DFFARX1 I_47(n_266_and_0_3_r_13,blif_clk_net_1_r_11,n9_11,n44_11,);
DFFARX1 I_48(G42_1_r_13,blif_clk_net_1_r_11,n9_11,n45_11,);
not I_49(n27_11,n45_11);
nor I_50(n4_1_r_11,n44_11,n25_11);
nor I_51(N3_2_r_11,n45_11,n40_11);
nand I_52(n24_11,n39_11,n_549_1_r_13);
nand I_53(n25_11,n38_11,P6_5_r_13);
DFFARX1 I_54(n25_11,blif_clk_net_1_r_11,n9_11,n20_internal_11,);
not I_55(n20_11,n20_internal_11);
not I_56(n28_11,n25_11);
not I_57(n29_11,G42_1_r_13);
nand I_58(n30_11,n26_11,n31_11);
not I_59(n31_11,n_572_1_r_13);
and I_60(n32_11,n26_11,n44_11);
and I_61(n33_11,n34_11,ACVQN2_3_r_13);
nor I_62(n34_11,n29_11,n_573_1_r_13);
not I_63(n35_11,n_452_1_r_13);
nand I_64(n36_11,n31_11,G42_1_r_13);
nor I_65(n37_11,n29_11,n_572_1_r_13);
nor I_66(n38_11,n31_11,n_452_1_r_13);
nor I_67(n39_11,n_452_1_r_13,ACVQN1_5_r_13);
nor I_68(n40_11,n41_11,n_452_1_r_13);
nor I_69(n41_11,n42_11,ACVQN1_5_r_13);
not I_70(n42_11,n_549_1_r_13);
endmodule


