module test_final(IN_1_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_6_1_l_12,IN_1_5_l_12,IN_2_5_l_12,IN_3_5_l_12,IN_6_5_l_12,blif_reset_net_0_r_2,blif_clk_net_0_r_2,ACVQN2_0_r_2,n_266_and_0_0_r_2,G199_1_r_2,G214_1_r_2,n_429_or_0_3_r_2,G78_3_r_2,n_576_3_r_2,n_102_3_r_2,n_547_3_r_2,n_42_5_r_2,G199_5_r_2);
input IN_1_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_6_1_l_12,IN_1_5_l_12,IN_2_5_l_12,IN_3_5_l_12,IN_6_5_l_12,blif_reset_net_0_r_2,blif_clk_net_0_r_2;
output ACVQN2_0_r_2,n_266_and_0_0_r_2,G199_1_r_2,G214_1_r_2,n_429_or_0_3_r_2,G78_3_r_2,n_576_3_r_2,n_102_3_r_2,n_547_3_r_2,n_42_5_r_2,G199_5_r_2;
wire ACVQN2_0_r_12,n_266_and_0_0_r_12,G199_1_r_12,G214_1_r_12,n_429_or_0_3_r_12,G78_3_r_12,n_576_3_r_12,n_102_3_r_12,n_547_3_r_12,n_42_5_r_12,G199_5_r_12,ACVQN2_0_l_12,n_266_and_0_0_l_12,ACVQN1_0_l_12,N1_1_l_12,G199_1_l_12,G214_1_l_12,n3_1_l_12,n_42_5_l_12,N3_5_l_12,G199_5_l_12,n3_5_l_12,ACVQN1_0_r_12,N1_1_r_12,n3_1_r_12,n12_3_r_12,n_431_3_r_12,n11_3_r_12,n13_3_r_12,n14_3_r_12,n15_3_r_12,n16_3_r_12,N3_5_r_12,n3_5_r_12,n1_0_r_2,ACVQN1_2_l_2,P6_2_l_2,P6_internal_2_l_2,n_429_or_0_3_l_2,n12_3_l_2,n_431_3_l_2,G78_3_l_2,n_576_3_l_2,n11_3_l_2,n_102_3_l_2,n_547_3_l_2,n13_3_l_2,n14_3_l_2,n15_3_l_2,n16_3_l_2,ACVQN1_0_r_2,N1_1_r_2,n3_1_r_2,n12_3_r_2,n_431_3_r_2,n11_3_r_2,n13_3_r_2,n14_3_r_2,n15_3_r_2,n16_3_r_2,N3_5_r_2,n3_5_r_2;
DFFARX1 I_0(G199_1_l_12,blif_clk_net_0_r_2,n1_0_r_2,ACVQN2_0_r_12,);
and I_1(n_266_and_0_0_r_12,ACVQN2_0_l_12,ACVQN1_0_r_12);
DFFARX1 I_2(N1_1_r_12,blif_clk_net_0_r_2,n1_0_r_2,G199_1_r_12,);
DFFARX1 I_3(G214_1_l_12,blif_clk_net_0_r_2,n1_0_r_2,G214_1_r_12,);
nand I_4(n_429_or_0_3_r_12,G199_1_l_12,n12_3_r_12);
DFFARX1 I_5(n_431_3_r_12,blif_clk_net_0_r_2,n1_0_r_2,G78_3_r_12,);
nand I_6(n_576_3_r_12,G214_1_l_12,n11_3_r_12);
not I_7(n_102_3_r_12,ACVQN2_0_l_12);
nand I_8(n_547_3_r_12,n_266_and_0_0_l_12,n13_3_r_12);
nor I_9(n_42_5_r_12,n_266_and_0_0_l_12,n_42_5_l_12);
DFFARX1 I_10(N3_5_r_12,blif_clk_net_0_r_2,n1_0_r_2,G199_5_r_12,);
DFFARX1 I_11(IN_1_0_l_12,blif_clk_net_0_r_2,n1_0_r_2,ACVQN2_0_l_12,);
and I_12(n_266_and_0_0_l_12,IN_4_0_l_12,ACVQN1_0_l_12);
DFFARX1 I_13(IN_2_0_l_12,blif_clk_net_0_r_2,n1_0_r_2,ACVQN1_0_l_12,);
and I_14(N1_1_l_12,IN_6_1_l_12,n3_1_l_12);
DFFARX1 I_15(N1_1_l_12,blif_clk_net_0_r_2,n1_0_r_2,G199_1_l_12,);
DFFARX1 I_16(IN_3_1_l_12,blif_clk_net_0_r_2,n1_0_r_2,G214_1_l_12,);
nand I_17(n3_1_l_12,IN_1_1_l_12,IN_2_1_l_12);
nor I_18(n_42_5_l_12,IN_1_5_l_12,IN_3_5_l_12);
and I_19(N3_5_l_12,IN_6_5_l_12,n3_5_l_12);
DFFARX1 I_20(N3_5_l_12,blif_clk_net_0_r_2,n1_0_r_2,G199_5_l_12,);
nand I_21(n3_5_l_12,IN_2_5_l_12,IN_3_5_l_12);
DFFARX1 I_22(ACVQN2_0_l_12,blif_clk_net_0_r_2,n1_0_r_2,ACVQN1_0_r_12,);
and I_23(N1_1_r_12,G199_1_l_12,n3_1_r_12);
nand I_24(n3_1_r_12,G214_1_l_12,n_42_5_l_12);
not I_25(n12_3_r_12,n_266_and_0_0_l_12);
or I_26(n_431_3_r_12,n_266_and_0_0_l_12,n14_3_r_12);
nor I_27(n11_3_r_12,G199_5_l_12,n12_3_r_12);
nor I_28(n13_3_r_12,ACVQN2_0_l_12,G199_5_l_12);
and I_29(n14_3_r_12,n_42_5_l_12,n15_3_r_12);
nor I_30(n15_3_r_12,G199_5_l_12,n16_3_r_12);
not I_31(n16_3_r_12,G199_1_l_12);
and I_32(N3_5_r_12,ACVQN2_0_l_12,n3_5_r_12);
nand I_33(n3_5_r_12,n_266_and_0_0_l_12,G199_1_l_12);
DFFARX1 I_34(P6_2_l_2,blif_clk_net_0_r_2,n1_0_r_2,ACVQN2_0_r_2,);
and I_35(n_266_and_0_0_r_2,n_102_3_l_2,ACVQN1_0_r_2);
DFFARX1 I_36(N1_1_r_2,blif_clk_net_0_r_2,n1_0_r_2,G199_1_r_2,);
DFFARX1 I_37(n_547_3_l_2,blif_clk_net_0_r_2,n1_0_r_2,G214_1_r_2,);
nand I_38(n_429_or_0_3_r_2,ACVQN1_2_l_2,n12_3_r_2);
DFFARX1 I_39(n_431_3_r_2,blif_clk_net_0_r_2,n1_0_r_2,G78_3_r_2,);
nand I_40(n_576_3_r_2,ACVQN1_2_l_2,n11_3_r_2);
not I_41(n_102_3_r_2,G78_3_l_2);
nand I_42(n_547_3_r_2,n_102_3_l_2,n13_3_r_2);
nor I_43(n_42_5_r_2,ACVQN1_2_l_2,P6_2_l_2);
DFFARX1 I_44(N3_5_r_2,blif_clk_net_0_r_2,n1_0_r_2,G199_5_r_2,);
not I_45(n1_0_r_2,blif_reset_net_0_r_2);
DFFARX1 I_46(n_576_3_r_12,blif_clk_net_0_r_2,n1_0_r_2,ACVQN1_2_l_2,);
not I_47(P6_2_l_2,P6_internal_2_l_2);
DFFARX1 I_48(n_547_3_r_12,blif_clk_net_0_r_2,n1_0_r_2,P6_internal_2_l_2,);
nand I_49(n_429_or_0_3_l_2,n12_3_l_2,G199_5_r_12);
not I_50(n12_3_l_2,G199_1_r_12);
or I_51(n_431_3_l_2,n14_3_l_2,n_42_5_r_12);
DFFARX1 I_52(n_431_3_l_2,blif_clk_net_0_r_2,n1_0_r_2,G78_3_l_2,);
nand I_53(n_576_3_l_2,n11_3_l_2,n_429_or_0_3_r_12);
nor I_54(n11_3_l_2,n12_3_l_2,n_102_3_r_12);
not I_55(n_102_3_l_2,n_102_3_r_12);
nand I_56(n_547_3_l_2,n13_3_l_2,G78_3_r_12);
nor I_57(n13_3_l_2,n_266_and_0_0_r_12,n_102_3_r_12);
and I_58(n14_3_l_2,n15_3_l_2,G214_1_r_12);
nor I_59(n15_3_l_2,n16_3_l_2,ACVQN2_0_r_12);
not I_60(n16_3_l_2,G199_5_r_12);
DFFARX1 I_61(G78_3_l_2,blif_clk_net_0_r_2,n1_0_r_2,ACVQN1_0_r_2,);
and I_62(N1_1_r_2,G78_3_l_2,n3_1_r_2);
nand I_63(n3_1_r_2,n_576_3_l_2,n_547_3_l_2);
not I_64(n12_3_r_2,n_429_or_0_3_l_2);
or I_65(n_431_3_r_2,n_429_or_0_3_l_2,n14_3_r_2);
nor I_66(n11_3_r_2,G78_3_l_2,n12_3_r_2);
nor I_67(n13_3_r_2,G78_3_l_2,n_576_3_l_2);
and I_68(n14_3_r_2,n_576_3_l_2,n15_3_r_2);
nor I_69(n15_3_r_2,P6_2_l_2,n16_3_r_2);
not I_70(n16_3_r_2,ACVQN1_2_l_2);
and I_71(N3_5_r_2,n_102_3_l_2,n3_5_r_2);
nand I_72(n3_5_r_2,ACVQN1_2_l_2,n_429_or_0_3_l_2);
endmodule


