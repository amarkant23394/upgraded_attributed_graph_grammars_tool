module test_I7547(I6657,I6705,I1470_clk,I1477_rst,I7547);
input I6657,I6705,I1470_clk,I1477_rst;
output I7547;
wire I7977,I6321,I7570_rst,I8059;
not I_0(I7547,I8059);
DFFARX1 I_1 (I6321,I1470_clk,I7570_rst,I7977);
nand I_2(I6321,I6705,I6657);
not I_3(I7570_rst,I1477_rst);
DFFARX1 I_4 (I7977,I1470_clk,I7570_rst,I8059);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule