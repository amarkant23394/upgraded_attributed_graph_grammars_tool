module test_I12783(I1477,I1470,I12783);
input I1477,I1470;
output I12783;
wire I12619,I10647,I9468,I12735,I10630,I11009;
not I_0(I12619,I1477);
not I_1(I10647,I1477);
DFFARX1 I_2(I12735,I1470,I12619,,,I12783,);
DFFARX1 I_3(I1470,,,I9468,);
DFFARX1 I_4(I10630,I1470,I12619,,,I12735,);
not I_5(I10630,I11009);
DFFARX1 I_6(I9468,I1470,I10647,,,I11009,);
endmodule


