module test_I3405(I1784,I1477,I1215,I1470,I1569,I1832,I3405);
input I1784,I1477,I1215,I1470,I1569,I1832;
output I3405;
wire I1518,I1637,I1480,I2038,I1976,I1880,I1495,I2103,I2021,I1849,I1959;
not I_0(I1518,I1477);
not I_1(I1637,I1215);
DFFARX1 I_2(I1976,I1470,I1518,,,I1480,);
not I_3(I2038,I2021);
or I_4(I3405,I1480,I1495);
and I_5(I1976,I1637,I1959);
DFFARX1 I_6(I1470,I1518,,,I1880,);
DFFARX1 I_7(I2103,I1470,I1518,,,I1495,);
or I_8(I2103,I2038,I1849);
DFFARX1 I_9(I1470,I1518,,,I2021,);
and I_10(I1849,I1832,I1784);
nand I_11(I1959,I1880,I1569);
endmodule


