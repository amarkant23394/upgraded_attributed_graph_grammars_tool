module test_I11272(I8845,I8836,I1477,I1470,I9083,I9413,I11272);
input I8845,I8836,I1477,I1470,I9083,I9413;
output I11272;
wire I11672,I11361,I11429,I11344,I11768,I8848,I11310,I11751;
DFFARX1 I_0(I8836,I1470,I11310,,,I11672,);
nand I_1(I11361,I11344,I8845);
not I_2(I11429,I8848);
nor I_3(I11344,I8848);
and I_4(I11768,I11429,I11751);
DFFARX1 I_5(I11768,I1470,I11310,,,I11272,);
nor I_6(I8848,I9083,I9413);
not I_7(I11310,I1477);
nand I_8(I11751,I11672,I11361);
endmodule


