module test_I8445(I6062,I6127,I1477,I5785,I1470,I8445);
input I6062,I6127,I1477,I5785,I1470;
output I8445;
wire I8394,I5728,I8428,I5751,I5713,I6203,I8411,I5833,I5725,I5802,I5734,I6144;
not I_0(I8394,I5713);
not I_1(I5728,I5833);
and I_2(I8428,I8411,I5734);
not I_3(I5751,I1477);
DFFARX1 I_4(I6127,I1470,I5751,,,I5713,);
DFFARX1 I_5(I1470,I5751,,,I6203,);
nor I_6(I8411,I8394,I5725);
DFFARX1 I_7(I5802,I1470,I5751,,,I5833,);
or I_8(I8445,I8428,I5728);
DFFARX1 I_9(I6203,I1470,I5751,,,I5725,);
DFFARX1 I_10(I5785,I1470,I5751,,,I5802,);
DFFARX1 I_11(I6144,I1470,I5751,,,I5734,);
or I_12(I6144,I6127,I6062);
endmodule


