module test_I9491(I1477,I9491);
input I1477;
output I9491;
wire ;
not I_0(I9491,I1477);
endmodule


