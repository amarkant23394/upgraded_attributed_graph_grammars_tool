module test_final(IN_1_0_l_3,IN_2_0_l_3,IN_4_0_l_3,G18_4_l_3,G15_4_l_3,IN_1_4_l_3,IN_4_4_l_3,IN_5_4_l_3,IN_7_4_l_3,IN_9_4_l_3,IN_10_4_l_3,blif_reset_net_0_r_12,blif_clk_net_0_r_12,ACVQN2_0_r_12,n_266_and_0_0_r_12,G199_1_r_12,G214_1_r_12,n_429_or_0_3_r_12,G78_3_r_12,n_576_3_r_12,n_102_3_r_12,n_547_3_r_12,n_42_5_r_12,G199_5_r_12);
input IN_1_0_l_3,IN_2_0_l_3,IN_4_0_l_3,G18_4_l_3,G15_4_l_3,IN_1_4_l_3,IN_4_4_l_3,IN_5_4_l_3,IN_7_4_l_3,IN_9_4_l_3,IN_10_4_l_3,blif_reset_net_0_r_12,blif_clk_net_0_r_12;
output ACVQN2_0_r_12,n_266_and_0_0_r_12,G199_1_r_12,G214_1_r_12,n_429_or_0_3_r_12,G78_3_r_12,n_576_3_r_12,n_102_3_r_12,n_547_3_r_12,n_42_5_r_12,G199_5_r_12;
wire ACVQN2_0_r_3,n_266_and_0_0_r_3,G199_1_r_3,G214_1_r_3,ACVQN1_2_r_3,P6_2_r_3,n_429_or_0_3_r_3,G78_3_r_3,n_576_3_r_3,n_102_3_r_3,n_547_3_r_3,ACVQN2_0_l_3,n_266_and_0_0_l_3,ACVQN1_0_l_3,n4_4_l_3,G42_4_l_3,n_87_4_l_3,n_572_4_l_3,n_573_4_l_3,n_549_4_l_3,n7_4_l_3,n_569_4_l_3,n_452_4_l_3,ACVQN1_0_r_3,N1_1_r_3,n3_1_r_3,P6_internal_2_r_3,n12_3_r_3,n_431_3_r_3,n11_3_r_3,n13_3_r_3,n14_3_r_3,n15_3_r_3,n16_3_r_3,n1_0_r_12,ACVQN2_0_l_12,n_266_and_0_0_l_12,ACVQN1_0_l_12,N1_1_l_12,G199_1_l_12,G214_1_l_12,n3_1_l_12,n_42_5_l_12,N3_5_l_12,G199_5_l_12,n3_5_l_12,ACVQN1_0_r_12,N1_1_r_12,n3_1_r_12,n12_3_r_12,n_431_3_r_12,n11_3_r_12,n13_3_r_12,n14_3_r_12,n15_3_r_12,n16_3_r_12,N3_5_r_12,n3_5_r_12;
DFFARX1 I_0(n_266_and_0_0_l_3,blif_clk_net_0_r_12,n1_0_r_12,ACVQN2_0_r_3,);
and I_1(n_266_and_0_0_r_3,n_572_4_l_3,ACVQN1_0_r_3);
DFFARX1 I_2(N1_1_r_3,blif_clk_net_0_r_12,n1_0_r_12,G199_1_r_3,);
DFFARX1 I_3(ACVQN2_0_l_3,blif_clk_net_0_r_12,n1_0_r_12,G214_1_r_3,);
DFFARX1 I_4(n_573_4_l_3,blif_clk_net_0_r_12,n1_0_r_12,ACVQN1_2_r_3,);
not I_5(P6_2_r_3,P6_internal_2_r_3);
nand I_6(n_429_or_0_3_r_3,ACVQN2_0_l_3,n12_3_r_3);
DFFARX1 I_7(n_431_3_r_3,blif_clk_net_0_r_12,n1_0_r_12,G78_3_r_3,);
nand I_8(n_576_3_r_3,n_452_4_l_3,n11_3_r_3);
not I_9(n_102_3_r_3,ACVQN2_0_l_3);
nand I_10(n_547_3_r_3,n_549_4_l_3,n13_3_r_3);
DFFARX1 I_11(IN_1_0_l_3,blif_clk_net_0_r_12,n1_0_r_12,ACVQN2_0_l_3,);
and I_12(n_266_and_0_0_l_3,IN_4_0_l_3,ACVQN1_0_l_3);
DFFARX1 I_13(IN_2_0_l_3,blif_clk_net_0_r_12,n1_0_r_12,ACVQN1_0_l_3,);
nor I_14(n4_4_l_3,G18_4_l_3,IN_1_4_l_3);
DFFARX1 I_15(n4_4_l_3,blif_clk_net_0_r_12,n1_0_r_12,G42_4_l_3,);
not I_16(n_87_4_l_3,G15_4_l_3);
nor I_17(n_572_4_l_3,G15_4_l_3,IN_7_4_l_3);
or I_18(n_573_4_l_3,IN_5_4_l_3,IN_9_4_l_3);
nor I_19(n_549_4_l_3,IN_10_4_l_3,n7_4_l_3);
and I_20(n7_4_l_3,IN_4_4_l_3,n_87_4_l_3);
or I_21(n_569_4_l_3,IN_9_4_l_3,IN_10_4_l_3);
nor I_22(n_452_4_l_3,G18_4_l_3,IN_5_4_l_3);
DFFARX1 I_23(n_452_4_l_3,blif_clk_net_0_r_12,n1_0_r_12,ACVQN1_0_r_3,);
and I_24(N1_1_r_3,n_549_4_l_3,n3_1_r_3);
nand I_25(n3_1_r_3,G42_4_l_3,n_569_4_l_3);
DFFARX1 I_26(n_266_and_0_0_l_3,blif_clk_net_0_r_12,n1_0_r_12,P6_internal_2_r_3,);
not I_27(n12_3_r_3,n_572_4_l_3);
or I_28(n_431_3_r_3,n_569_4_l_3,n14_3_r_3);
nor I_29(n11_3_r_3,ACVQN2_0_l_3,n12_3_r_3);
nor I_30(n13_3_r_3,ACVQN2_0_l_3,G42_4_l_3);
and I_31(n14_3_r_3,n_266_and_0_0_l_3,n15_3_r_3);
nor I_32(n15_3_r_3,n_573_4_l_3,n16_3_r_3);
not I_33(n16_3_r_3,ACVQN2_0_l_3);
DFFARX1 I_34(G199_1_l_12,blif_clk_net_0_r_12,n1_0_r_12,ACVQN2_0_r_12,);
and I_35(n_266_and_0_0_r_12,ACVQN2_0_l_12,ACVQN1_0_r_12);
DFFARX1 I_36(N1_1_r_12,blif_clk_net_0_r_12,n1_0_r_12,G199_1_r_12,);
DFFARX1 I_37(G214_1_l_12,blif_clk_net_0_r_12,n1_0_r_12,G214_1_r_12,);
nand I_38(n_429_or_0_3_r_12,G199_1_l_12,n12_3_r_12);
DFFARX1 I_39(n_431_3_r_12,blif_clk_net_0_r_12,n1_0_r_12,G78_3_r_12,);
nand I_40(n_576_3_r_12,G214_1_l_12,n11_3_r_12);
not I_41(n_102_3_r_12,ACVQN2_0_l_12);
nand I_42(n_547_3_r_12,n_266_and_0_0_l_12,n13_3_r_12);
nor I_43(n_42_5_r_12,n_266_and_0_0_l_12,n_42_5_l_12);
DFFARX1 I_44(N3_5_r_12,blif_clk_net_0_r_12,n1_0_r_12,G199_5_r_12,);
not I_45(n1_0_r_12,blif_reset_net_0_r_12);
DFFARX1 I_46(ACVQN1_2_r_3,blif_clk_net_0_r_12,n1_0_r_12,ACVQN2_0_l_12,);
and I_47(n_266_and_0_0_l_12,ACVQN1_0_l_12,G199_1_r_3);
DFFARX1 I_48(G78_3_r_3,blif_clk_net_0_r_12,n1_0_r_12,ACVQN1_0_l_12,);
and I_49(N1_1_l_12,n3_1_l_12,n_266_and_0_0_r_3);
DFFARX1 I_50(N1_1_l_12,blif_clk_net_0_r_12,n1_0_r_12,G199_1_l_12,);
DFFARX1 I_51(G214_1_r_3,blif_clk_net_0_r_12,n1_0_r_12,G214_1_l_12,);
nand I_52(n3_1_l_12,ACVQN2_0_r_3,n_576_3_r_3);
nor I_53(n_42_5_l_12,P6_2_r_3,n_429_or_0_3_r_3);
and I_54(N3_5_l_12,n3_5_l_12,n_102_3_r_3);
DFFARX1 I_55(N3_5_l_12,blif_clk_net_0_r_12,n1_0_r_12,G199_5_l_12,);
nand I_56(n3_5_l_12,P6_2_r_3,n_547_3_r_3);
DFFARX1 I_57(ACVQN2_0_l_12,blif_clk_net_0_r_12,n1_0_r_12,ACVQN1_0_r_12,);
and I_58(N1_1_r_12,G199_1_l_12,n3_1_r_12);
nand I_59(n3_1_r_12,G214_1_l_12,n_42_5_l_12);
not I_60(n12_3_r_12,n_266_and_0_0_l_12);
or I_61(n_431_3_r_12,n_266_and_0_0_l_12,n14_3_r_12);
nor I_62(n11_3_r_12,G199_5_l_12,n12_3_r_12);
nor I_63(n13_3_r_12,ACVQN2_0_l_12,G199_5_l_12);
and I_64(n14_3_r_12,n_42_5_l_12,n15_3_r_12);
nor I_65(n15_3_r_12,G199_5_l_12,n16_3_r_12);
not I_66(n16_3_r_12,G199_1_l_12);
and I_67(N3_5_r_12,ACVQN2_0_l_12,n3_5_r_12);
nand I_68(n3_5_r_12,n_266_and_0_0_l_12,G199_1_l_12);
endmodule


