module test_I14162(I10032,I1477,I1470,I12191,I14162);
input I10032,I1477,I1470,I12191;
output I14162;
wire I12270,I10219,I12239,I10014,I11938,I12208,I13775,I11990,I11973,I10052;
nand I_0(I12270,I11990,I10014);
DFFARX1 I_1(I1470,I10052,,,I10219,);
DFFARX1 I_2(I12208,I1470,I11973,,,I12239,);
DFFARX1 I_3(I11938,I1470,I13775,,,I14162,);
DFFARX1 I_4(I10219,I1470,I10052,,,I10014,);
and I_5(I11938,I12270,I12239);
DFFARX1 I_6(I12191,I1470,I11973,,,I12208,);
not I_7(I13775,I1477);
not I_8(I11990,I10032);
not I_9(I11973,I1477);
not I_10(I10052,I1477);
endmodule


