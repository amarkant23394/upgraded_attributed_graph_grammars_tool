module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_4_0_l_14,IN_1_1_l_14,IN_2_1_l_14,IN_3_1_l_14,IN_6_1_l_14,IN_1_5_l_14,IN_2_5_l_14,IN_3_5_l_14,IN_6_5_l_14,blif_clk_net_3_r_0,blif_reset_net_3_r_0,n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0);
input IN_1_0_l_14,IN_2_0_l_14,IN_4_0_l_14,IN_1_1_l_14,IN_2_1_l_14,IN_3_1_l_14,IN_6_1_l_14,IN_1_5_l_14,IN_2_5_l_14,IN_3_5_l_14,IN_6_5_l_14,blif_clk_net_3_r_0,blif_reset_net_3_r_0;
output n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0;
wire ACVQN2_0_r_14,n_266_and_0_0_r_14,G199_1_r_14,G214_1_r_14,ACVQN1_2_r_14,P6_2_r_14,n_429_or_0_3_r_14,G78_3_r_14,n_576_3_r_14,n_102_3_r_14,n_547_3_r_14,ACVQN2_0_l_14,n_266_and_0_0_l_14,ACVQN1_0_l_14,N1_1_l_14,G199_1_l_14,G214_1_l_14,n3_1_l_14,n_42_5_l_14,N3_5_l_14,G199_5_l_14,n3_5_l_14,ACVQN1_0_r_14,N1_1_r_14,n3_1_r_14,P6_internal_2_r_14,n12_3_r_14,n_431_3_r_14,n11_3_r_14,n13_3_r_14,n14_3_r_14,n15_3_r_14,n16_3_r_14,n2_3_r_0,ACVQN2_0_l_0,n_266_and_0_0_l_0,ACVQN1_0_l_0,N1_1_l_0,G199_1_l_0,G214_1_l_0,n3_1_l_0,n_42_5_l_0,N3_5_l_0,G199_5_l_0,n3_5_l_0,n12_3_r_0,n_431_3_r_0,n11_3_r_0,n13_3_r_0,n14_3_r_0,n15_3_r_0,n16_3_r_0,n4_4_r_0,n_87_4_r_0,n7_4_r_0;
DFFARX1 I_0(n_266_and_0_0_l_14,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_r_14,);
and I_1(n_266_and_0_0_r_14,G199_5_l_14,ACVQN1_0_r_14);
DFFARX1 I_2(N1_1_r_14,blif_clk_net_3_r_0,n2_3_r_0,G199_1_r_14,);
DFFARX1 I_3(G199_1_l_14,blif_clk_net_3_r_0,n2_3_r_0,G214_1_r_14,);
DFFARX1 I_4(ACVQN2_0_l_14,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_2_r_14,);
not I_5(P6_2_r_14,P6_internal_2_r_14);
nand I_6(n_429_or_0_3_r_14,G214_1_l_14,n12_3_r_14);
DFFARX1 I_7(n_431_3_r_14,blif_clk_net_3_r_0,n2_3_r_0,G78_3_r_14,);
nand I_8(n_576_3_r_14,ACVQN2_0_l_14,n11_3_r_14);
not I_9(n_102_3_r_14,G199_5_l_14);
nand I_10(n_547_3_r_14,n_266_and_0_0_l_14,n13_3_r_14);
DFFARX1 I_11(IN_1_0_l_14,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_l_14,);
and I_12(n_266_and_0_0_l_14,IN_4_0_l_14,ACVQN1_0_l_14);
DFFARX1 I_13(IN_2_0_l_14,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_l_14,);
and I_14(N1_1_l_14,IN_6_1_l_14,n3_1_l_14);
DFFARX1 I_15(N1_1_l_14,blif_clk_net_3_r_0,n2_3_r_0,G199_1_l_14,);
DFFARX1 I_16(IN_3_1_l_14,blif_clk_net_3_r_0,n2_3_r_0,G214_1_l_14,);
nand I_17(n3_1_l_14,IN_1_1_l_14,IN_2_1_l_14);
nor I_18(n_42_5_l_14,IN_1_5_l_14,IN_3_5_l_14);
and I_19(N3_5_l_14,IN_6_5_l_14,n3_5_l_14);
DFFARX1 I_20(N3_5_l_14,blif_clk_net_3_r_0,n2_3_r_0,G199_5_l_14,);
nand I_21(n3_5_l_14,IN_2_5_l_14,IN_3_5_l_14);
DFFARX1 I_22(G214_1_l_14,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_r_14,);
and I_23(N1_1_r_14,G214_1_l_14,n3_1_r_14);
nand I_24(n3_1_r_14,ACVQN2_0_l_14,n_42_5_l_14);
DFFARX1 I_25(G199_5_l_14,blif_clk_net_3_r_0,n2_3_r_0,P6_internal_2_r_14,);
not I_26(n12_3_r_14,n_42_5_l_14);
or I_27(n_431_3_r_14,n_266_and_0_0_l_14,n14_3_r_14);
nor I_28(n11_3_r_14,G199_5_l_14,n12_3_r_14);
nor I_29(n13_3_r_14,G199_1_l_14,G199_5_l_14);
and I_30(n14_3_r_14,n_42_5_l_14,n15_3_r_14);
nor I_31(n15_3_r_14,G199_1_l_14,n16_3_r_14);
not I_32(n16_3_r_14,G214_1_l_14);
nand I_33(n_429_or_0_3_r_0,ACVQN2_0_l_0,n12_3_r_0);
DFFARX1 I_34(n_431_3_r_0,blif_clk_net_3_r_0,n2_3_r_0,G78_3_r_0,);
nand I_35(n_576_3_r_0,n_266_and_0_0_l_0,n11_3_r_0);
not I_36(n_102_3_r_0,n_42_5_l_0);
nand I_37(n_547_3_r_0,ACVQN2_0_l_0,n13_3_r_0);
DFFARX1 I_38(n4_4_r_0,blif_clk_net_3_r_0,n2_3_r_0,G42_4_r_0,);
nor I_39(n_572_4_r_0,G199_1_l_0,G199_5_l_0);
or I_40(n_573_4_r_0,n_42_5_l_0,G199_5_l_0);
nor I_41(n_549_4_r_0,n_266_and_0_0_l_0,n7_4_r_0);
or I_42(n_569_4_r_0,n_266_and_0_0_l_0,n_42_5_l_0);
nor I_43(n_452_4_r_0,ACVQN2_0_l_0,G199_5_l_0);
not I_44(n2_3_r_0,blif_reset_net_3_r_0);
DFFARX1 I_45(G199_1_r_14,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_l_0,);
and I_46(n_266_and_0_0_l_0,ACVQN1_0_l_0,ACVQN2_0_r_14);
DFFARX1 I_47(n_102_3_r_14,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_l_0,);
and I_48(N1_1_l_0,n3_1_l_0,P6_2_r_14);
DFFARX1 I_49(N1_1_l_0,blif_clk_net_3_r_0,n2_3_r_0,G199_1_l_0,);
DFFARX1 I_50(ACVQN1_2_r_14,blif_clk_net_3_r_0,n2_3_r_0,G214_1_l_0,);
nand I_51(n3_1_l_0,n_266_and_0_0_r_14,G78_3_r_14);
nor I_52(n_42_5_l_0,n_576_3_r_14,n_547_3_r_14);
and I_53(N3_5_l_0,n3_5_l_0,n_429_or_0_3_r_14);
DFFARX1 I_54(N3_5_l_0,blif_clk_net_3_r_0,n2_3_r_0,G199_5_l_0,);
nand I_55(n3_5_l_0,G214_1_r_14,n_547_3_r_14);
not I_56(n12_3_r_0,G199_1_l_0);
or I_57(n_431_3_r_0,n_266_and_0_0_l_0,n14_3_r_0);
nor I_58(n11_3_r_0,G214_1_l_0,n12_3_r_0);
nor I_59(n13_3_r_0,G214_1_l_0,n_42_5_l_0);
and I_60(n14_3_r_0,n_42_5_l_0,n15_3_r_0);
nor I_61(n15_3_r_0,G199_1_l_0,n16_3_r_0);
not I_62(n16_3_r_0,ACVQN2_0_l_0);
nor I_63(n4_4_r_0,ACVQN2_0_l_0,G214_1_l_0);
not I_64(n_87_4_r_0,G199_5_l_0);
and I_65(n7_4_r_0,ACVQN2_0_l_0,n_87_4_r_0);
endmodule


