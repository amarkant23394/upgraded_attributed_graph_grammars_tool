module test_I10154(I8107,I7881,I1477,I1470,I8028,I10154);
input I8107,I7881,I1477,I1470,I8028;
output I10154;
wire I7898,I6297,I7538,I7714,I7570,I7946,I7535,I7915,I10137,I7553,I10052,I8124,I10120;
nand I_0(I7898,I7881);
DFFARX1 I_1(I1470,,,I6297,);
DFFARX1 I_2(I7915,I1470,I7570,,,I7538,);
not I_3(I7714,I6297);
nand I_4(I10154,I10137,I10120);
not I_5(I7570,I1477);
DFFARX1 I_6(I7881,I1470,I7570,,,I7946,);
and I_7(I7535,I7714,I7946);
and I_8(I7915,I7881,I7898);
DFFARX1 I_9(I7553,I1470,I10052,,,I10137,);
DFFARX1 I_10(I8124,I1470,I7570,,,I7553,);
not I_11(I10052,I1477);
or I_12(I8124,I8107,I8028);
nor I_13(I10120,I7538,I7535);
endmodule


