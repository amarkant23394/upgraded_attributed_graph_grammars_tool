module test_I12735(I1477,I1470,I9864,I12735);
input I1477,I1470,I9864;
output I12735;
wire I12619,I10647,I9491,I9468,I10630,I11009;
not I_0(I12619,I1477);
not I_1(I10647,I1477);
not I_2(I9491,I1477);
DFFARX1 I_3(I9864,I1470,I9491,,,I9468,);
DFFARX1 I_4(I10630,I1470,I12619,,,I12735,);
not I_5(I10630,I11009);
DFFARX1 I_6(I9468,I1470,I10647,,,I11009,);
endmodule


