module test_I10032(I8107,I7550,I1477,I8028,I1470,I10069,I10032);
input I8107,I7550,I1477,I8028,I1470,I10069;
output I10032;
wire I10349,I10086,I7570,I10414,I10397,I7553,I10137,I7544,I10052,I8124,I10103,I10332;
and I_0(I10349,I10332,I7550);
nand I_1(I10032,I10137,I10414);
and I_2(I10086,I10069,I7544);
not I_3(I7570,I1477);
nor I_4(I10414,I10103,I10397);
not I_5(I10397,I10349);
DFFARX1 I_6(I8124,I1470,I7570,,,I7553,);
DFFARX1 I_7(I7553,I1470,I10052,,,I10137,);
DFFARX1 I_8(I1470,I7570,,,I7544,);
not I_9(I10052,I1477);
or I_10(I8124,I8107,I8028);
DFFARX1 I_11(I10086,I1470,I10052,,,I10103,);
DFFARX1 I_12(I1470,I10052,,,I10332,);
endmodule


