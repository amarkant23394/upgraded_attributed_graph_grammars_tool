module test_I12602(I1477,I10766,I1470,I11088,I11026,I12602);
input I1477,I10766,I1470,I11088,I11026;
output I12602;
wire I12619,I11105,I12913,I10647,I12930,I10633,I10896,I10609;
not I_0(I12619,I1477);
not I_1(I12602,I12930);
and I_2(I11105,I10766,I11088);
DFFARX1 I_3(I10633,I1470,I12619,,,I12913,);
not I_4(I10647,I1477);
and I_5(I12930,I12913,I10609);
nand I_6(I10633,I10896,I11026);
DFFARX1 I_7(I1470,I10647,,,I10896,);
DFFARX1 I_8(I11105,I1470,I10647,,,I10609,);
endmodule


