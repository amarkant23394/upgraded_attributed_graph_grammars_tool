module test_I7550(I1477,I6843,I1470,I3972,I7550);
input I1477,I6843,I1470,I3972;
output I7550;
wire I6606,I6297,I6321,I7714,I7570,I6688,I6380,I7731,I6329,I6705,I7977,I6657;
DFFARX1 I_0(I1470,I6329,,,I6606,);
DFFARX1 I_1(I6843,I1470,I6329,,,I6297,);
nand I_2(I7550,I7977,I7731);
nand I_3(I6321,I6705,I6657);
not I_4(I7714,I6297);
not I_5(I7570,I1477);
DFFARX1 I_6(I1470,I6329,,,I6688,);
DFFARX1 I_7(I1470,I6329,,,I6380,);
not I_8(I7731,I7714);
not I_9(I6329,I1477);
and I_10(I6705,I6688,I3972);
DFFARX1 I_11(I6321,I1470,I7570,,,I7977,);
nor I_12(I6657,I6606,I6380);
endmodule


