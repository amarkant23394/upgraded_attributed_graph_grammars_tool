module test_I10103(I7714,I1477,I7604,I1470,I6315,I7669,I10103);
input I7714,I1477,I7604,I1470,I6315,I7669;
output I10103;
wire I10086,I7621,I7570,I7946,I7559,I7535,I7544,I10052,I10069;
and I_0(I10086,I10069,I7544);
nand I_1(I7621,I7604,I6315);
not I_2(I7570,I1477);
DFFARX1 I_3(I1470,I7570,,,I7946,);
not I_4(I7559,I7669);
and I_5(I7535,I7714,I7946);
DFFARX1 I_6(I7621,I1470,I7570,,,I7544,);
not I_7(I10052,I1477);
DFFARX1 I_8(I10086,I1470,I10052,,,I10103,);
nand I_9(I10069,I7559,I7535);
endmodule


