module test_final(IN_1_0_l_5,IN_2_0_l_5,IN_3_0_l_5,IN_4_0_l_5,IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_8_r_1,blif_reset_net_8_r_1,N6147_3_r_1,N1372_4_r_1,N1508_4_r_1,n_42_8_r_1,G199_8_r_1,N6147_9_r_1,N6134_9_r_1,N1372_10_r_1,N1508_10_r_1);
input IN_1_0_l_5,IN_2_0_l_5,IN_3_0_l_5,IN_4_0_l_5,IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_8_r_1,blif_reset_net_8_r_1;
output N6147_3_r_1,N1372_4_r_1,N1508_4_r_1,n_42_8_r_1,G199_8_r_1,N6147_9_r_1,N6134_9_r_1,N1372_10_r_1,N1508_10_r_1;
wire N1371_0_r_5,N1508_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1507_6_r_5,N1508_6_r_5,n_431_5_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,I_BUFF_1_9_r_1,N3_8_l_1,n7_1,n38_1,n22_1,N3_8_r_1,n23_1,n24_1,n25_1,n26_1,n27_1,n28_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1;
nor I_0(N1371_0_r_5,n28_5,n39_5);
not I_1(N1508_0_r_5,n39_5);
nor I_2(N6147_2_r_5,n28_5,n37_5);
nand I_3(n_429_or_0_5_r_5,n30_5,n32_5);
DFFARX1 I_4(n_431_5_r_5,blif_clk_net_8_r_1,n7_1,G78_5_r_5,);
nand I_5(n_576_5_r_5,n26_5,n27_5);
not I_6(n_102_5_r_5,n28_5);
nand I_7(n_547_5_r_5,n31_5,n32_5);
nor I_8(N1507_6_r_5,n30_5,n32_5);
nor I_9(N1508_6_r_5,n39_5,n41_5);
nand I_10(n_431_5_r_5,n34_5,n35_5);
nor I_11(n26_5,n29_5,n30_5);
nor I_12(n27_5,IN_2_0_l_5,n28_5);
nor I_13(n28_5,n29_5,n44_5);
not I_14(n29_5,IN_1_0_l_5);
nand I_15(n30_5,N1508_0_r_5,n43_5);
nor I_16(n31_5,n28_5,n33_5);
nor I_17(n32_5,IN_3_1_l_5,n40_5);
nor I_18(n33_5,IN_2_0_l_5,n29_5);
or I_19(n34_5,IN_2_0_l_5,n29_5);
nand I_20(n35_5,n32_5,n36_5);
not I_21(n36_5,n30_5);
nor I_22(n37_5,N1507_6_r_5,n38_5);
and I_23(n38_5,n39_5,n40_5);
nand I_24(n39_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_25(n40_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_26(n41_5,n28_5,n42_5);
or I_27(n42_5,n32_5,n36_5);
or I_28(n43_5,IN_3_10_l_5,IN_4_10_l_5);
nor I_29(n44_5,IN_3_0_l_5,IN_4_0_l_5);
nor I_30(N6147_3_r_1,n26_1,n27_1);
not I_31(N1372_4_r_1,n34_1);
nor I_32(N1508_4_r_1,n30_1,n34_1);
nor I_33(n_42_8_r_1,n23_1,n24_1);
DFFARX1 I_34(N3_8_r_1,blif_clk_net_8_r_1,n7_1,G199_8_r_1,);
nor I_35(N6147_9_r_1,n22_1,n25_1);
nor I_36(N6134_9_r_1,n29_1,n30_1);
not I_37(I_BUFF_1_9_r_1,n32_1);
not I_38(N1372_10_r_1,n36_1);
nor I_39(N1508_10_r_1,n35_1,n36_1);
and I_40(N3_8_l_1,n33_1,n_102_5_r_5);
not I_41(n7_1,blif_reset_net_8_r_1);
DFFARX1 I_42(N3_8_l_1,blif_clk_net_8_r_1,n7_1,n38_1,);
not I_43(n22_1,n38_1);
nor I_44(N3_8_r_1,n31_1,n32_1);
nor I_45(n23_1,n28_1,N1371_0_r_5);
nor I_46(n24_1,G78_5_r_5,N1508_6_r_5);
nor I_47(n25_1,n23_1,n26_1);
not I_48(n26_1,n30_1);
nand I_49(n27_1,n22_1,n28_1);
nand I_50(n28_1,n_576_5_r_5,n_429_or_0_5_r_5);
not I_51(n29_1,n28_1);
nand I_52(n30_1,n_429_or_0_5_r_5,n_547_5_r_5);
and I_53(n31_1,n38_1,n24_1);
nand I_54(n32_1,n26_1,n37_1);
nand I_55(n33_1,N6147_2_r_5,G78_5_r_5);
nand I_56(n34_1,n24_1,n29_1);
nor I_57(n35_1,n38_1,n24_1);
nand I_58(n36_1,I_BUFF_1_9_r_1,n23_1);
or I_59(n37_1,N1371_0_r_5,N6147_2_r_5);
endmodule


