module Benchmark_testing25000(I631,I639,I647,I655,I663,I671,I679,I687,I695,I703,I711,I719,I727,I735,I743,I751,I759,I767,I775,I783,I791,I799,I807,I815,I823,I831,I839,I847,I855,I863,I871,I879,I887,I895,I903,I911,I919,I927,I935,I943,I951,I959,I967,I975,I983,I991,I999,I1007,I1015,I1023,I1031,I1039,I1047,I1055,I1063,I1071,I1079,I1087,I1095,I1103,I1111,I1119,I1127,I1135,I1143,I1151,I1159,I1167,I1175,I1183,I1191,I1199,I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1862,I1869,I36445,I36454,I36457,I36448,I36442,I36436,I36439,I36451,I36433,I44095,I44104,I44107,I44098,I44092,I44086,I44089,I44101,I44083,I45625,I45634,I45637,I45628,I45622,I45616,I45619,I45631,I45613,I82345,I82354,I82357,I82348,I82342,I82336,I82339,I82351,I82333,I89995,I90004,I90007,I89998,I89992,I89986,I89989,I90001,I89983,I179505,I179523,I179526,I179508,I179529,I179514,I179517,I179511,I179520,I185302,I185320,I185323,I185305,I185326,I185311,I185314,I185308,I185317,I201558,I201543,I201537,I201540,I201546,I201555,I201552,I201549,I241542,I241527,I241521,I241524,I241530,I241539,I241536,I241533,I243446,I243431,I243425,I243428,I243434,I243443,I243440,I243437,I257726,I257711,I257705,I257708,I257714,I257723,I257720,I257717,I264866,I264851,I264845,I264848,I264854,I264863,I264860,I264857,I285810,I285795,I285789,I285792,I285798,I285807,I285804,I285801,I368135,I368132,I368120,I368126,I368129,I368123,I368138);
input I631,I639,I647,I655,I663,I671,I679,I687,I695,I703,I711,I719,I727,I735,I743,I751,I759,I767,I775,I783,I791,I799,I807,I815,I823,I831,I839,I847,I855,I863,I871,I879,I887,I895,I903,I911,I919,I927,I935,I943,I951,I959,I967,I975,I983,I991,I999,I1007,I1015,I1023,I1031,I1039,I1047,I1055,I1063,I1071,I1079,I1087,I1095,I1103,I1111,I1119,I1127,I1135,I1143,I1151,I1159,I1167,I1175,I1183,I1191,I1199,I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1862,I1869;
output I36445,I36454,I36457,I36448,I36442,I36436,I36439,I36451,I36433,I44095,I44104,I44107,I44098,I44092,I44086,I44089,I44101,I44083,I45625,I45634,I45637,I45628,I45622,I45616,I45619,I45631,I45613,I82345,I82354,I82357,I82348,I82342,I82336,I82339,I82351,I82333,I89995,I90004,I90007,I89998,I89992,I89986,I89989,I90001,I89983,I179505,I179523,I179526,I179508,I179529,I179514,I179517,I179511,I179520,I185302,I185320,I185323,I185305,I185326,I185311,I185314,I185308,I185317,I201558,I201543,I201537,I201540,I201546,I201555,I201552,I201549,I241542,I241527,I241521,I241524,I241530,I241539,I241536,I241533,I243446,I243431,I243425,I243428,I243434,I243443,I243440,I243437,I257726,I257711,I257705,I257708,I257714,I257723,I257720,I257717,I264866,I264851,I264845,I264848,I264854,I264863,I264860,I264857,I285810,I285795,I285789,I285792,I285798,I285807,I285804,I285801,I368135,I368132,I368120,I368126,I368129,I368123,I368138;
wire I631,I639,I647,I655,I663,I671,I679,I687,I695,I703,I711,I719,I727,I735,I743,I751,I759,I767,I775,I783,I791,I799,I807,I815,I823,I831,I839,I847,I855,I863,I871,I879,I887,I895,I903,I911,I919,I927,I935,I943,I951,I959,I967,I975,I983,I991,I999,I1007,I1015,I1023,I1031,I1039,I1047,I1055,I1063,I1071,I1079,I1087,I1095,I1103,I1111,I1119,I1127,I1135,I1143,I1151,I1159,I1167,I1175,I1183,I1191,I1199,I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1862,I1869,I1901,I1918,I145780,I145798,I1935,I145783,I145777,I1952,I1969,I1881,I2000,I145801,I2017,I145792,I2043,I2051,I2068,I2085,I2102,I2119,I2136,I2153,I1887,I2184,I145786,I2201,I2218,I145795,I145789,I1872,I2249,I2266,I2283,I1890,I1893,I2328,I1875,I1878,I2373,I1884,I2428,I2445,I2462,I2479,I2496,I2408,I2527,I2544,I2570,I2578,I2595,I2612,I2629,I2646,I2663,I2680,I2414,I2711,I2728,I2745,I2399,I2776,I2793,I2810,I2417,I2420,I2855,I2402,I2405,I2900,I2411,I2955,I2972,I337869,I337881,I2989,I337860,I337863,I3006,I3023,I2935,I3054,I337872,I3071,I337875,I3097,I3105,I3122,I3139,I337866,I3156,I3173,I3190,I3207,I2941,I3238,I3255,I3272,I337878,I2926,I3303,I3320,I3337,I2944,I2947,I3382,I2929,I2932,I3427,I2938,I3482,I3499,I363712,I363706,I3516,I363703,I3533,I3550,I3462,I3581,I363709,I363715,I3598,I3624,I3632,I3649,I3666,I363700,I3683,I3700,I3717,I3734,I3468,I3765,I3782,I3799,I363718,I3453,I3830,I3847,I3864,I3471,I3474,I3909,I3456,I3459,I3954,I3465,I4009,I4026,I18586,I4043,I18607,I18604,I4060,I4077,I3989,I4108,I18583,I18595,I4125,I18592,I4151,I4159,I4176,I4193,I18601,I4210,I4227,I4244,I4261,I3995,I4292,I4309,I4326,I18598,I18589,I3980,I4357,I4374,I4391,I3998,I4001,I4436,I3983,I3986,I4481,I3992,I4536,I4553,I384044,I384038,I4570,I384035,I4587,I4604,I4516,I4635,I384041,I384047,I4652,I4678,I4686,I4703,I4720,I384032,I4737,I4754,I4771,I4788,I4522,I4819,I4836,I4853,I384050,I4507,I4884,I4901,I4918,I4525,I4528,I4963,I4510,I4513,I5008,I4519,I5063,I5080,I355787,I355799,I5097,I355778,I355781,I5114,I5131,I5043,I5162,I355790,I5179,I355793,I5205,I5213,I5230,I5247,I355784,I5264,I5281,I5298,I5315,I5049,I5346,I5363,I5380,I355796,I5034,I5411,I5428,I5445,I5052,I5055,I5490,I5037,I5040,I5535,I5046,I5590,I5607,I272479,I272461,I5624,I272467,I272482,I5641,I5658,I5570,I5689,I272464,I272470,I5706,I5732,I5740,I5757,I5774,I272473,I5791,I5808,I5825,I5842,I5576,I5873,I5890,I5907,I272476,I5561,I5938,I5955,I5972,I5579,I5582,I6017,I5564,I5567,I6062,I5573,I6117,I6134,I184251,I184269,I6151,I184254,I184248,I6168,I6185,I6097,I6216,I184272,I6233,I184263,I6259,I6267,I6284,I6301,I6318,I6335,I6352,I6369,I6103,I6400,I184257,I6417,I6434,I184266,I184260,I6088,I6465,I6482,I6499,I6106,I6109,I6544,I6091,I6094,I6589,I6100,I6644,I6661,I64486,I6678,I64507,I64504,I6695,I6712,I6624,I6743,I64483,I64495,I6760,I64492,I6786,I6794,I6811,I6828,I64501,I6845,I6862,I6879,I6896,I6630,I6927,I6944,I6961,I64498,I64489,I6615,I6992,I7009,I7026,I6633,I6636,I7071,I6618,I6621,I7116,I6627,I7171,I7188,I175819,I175837,I7205,I175822,I175816,I7222,I7239,I7151,I7270,I175840,I7287,I175831,I7313,I7321,I7338,I7355,I7372,I7389,I7406,I7423,I7157,I7454,I175825,I7471,I7488,I175834,I175828,I7142,I7519,I7536,I7553,I7160,I7163,I7598,I7145,I7148,I7643,I7154,I7698,I7715,I38476,I7732,I38497,I38494,I7749,I7766,I7678,I7797,I38473,I38485,I7814,I38482,I7840,I7848,I7865,I7882,I38491,I7899,I7916,I7933,I7950,I7684,I7981,I7998,I8015,I38488,I38479,I7669,I8046,I8063,I8080,I7687,I7690,I8125,I7672,I7675,I8170,I7681,I8225,I8242,I169495,I169513,I8259,I169498,I169492,I8276,I8293,I8205,I8324,I169516,I8341,I169507,I8367,I8375,I8392,I8409,I8426,I8443,I8460,I8477,I8211,I8508,I169501,I8525,I8542,I169510,I169504,I8196,I8573,I8590,I8607,I8214,I8217,I8652,I8199,I8202,I8697,I8208,I8752,I8769,I219643,I219625,I8786,I219631,I219646,I8803,I8820,I8732,I8851,I219628,I219634,I8868,I8894,I8902,I8919,I8936,I219637,I8953,I8970,I8987,I9004,I8738,I9035,I9052,I9069,I219640,I8723,I9100,I9117,I9134,I8741,I8744,I9179,I8726,I8729,I9224,I8735,I9279,I9296,I134186,I134204,I9313,I134189,I134183,I9330,I9347,I9259,I9378,I134207,I9395,I134198,I9421,I9429,I9446,I9463,I9480,I9497,I9514,I9531,I9265,I9562,I134192,I9579,I9596,I134201,I134195,I9250,I9627,I9644,I9661,I9268,I9271,I9706,I9253,I9256,I9751,I9262,I9806,I9823,I291490,I291484,I9840,I291499,I291502,I9857,I9874,I9786,I9905,I291487,I9922,I9948,I9956,I9973,I9990,I291505,I10007,I10024,I10041,I10058,I9792,I10089,I10106,I10123,I291496,I291493,I9777,I10154,I10171,I10188,I9795,I9798,I10233,I9780,I9783,I10278,I9789,I10333,I10350,I246299,I246281,I10367,I246287,I246302,I10384,I10401,I10313,I10432,I246284,I246290,I10449,I10475,I10483,I10500,I10517,I246293,I10534,I10551,I10568,I10585,I10319,I10616,I10633,I10650,I246296,I10304,I10681,I10698,I10715,I10322,I10325,I10760,I10307,I10310,I10805,I10316,I10860,I10877,I332599,I332611,I10894,I332590,I332593,I10911,I10928,I10840,I10959,I332602,I10976,I332605,I11002,I11010,I11027,I11044,I332596,I11061,I11078,I11095,I11112,I10846,I11143,I11160,I11177,I332608,I10831,I11208,I11225,I11242,I10849,I10852,I11287,I10834,I10837,I11332,I10843,I11387,I11404,I71626,I11421,I71647,I71644,I11438,I11455,I11367,I11486,I71623,I71635,I11503,I71632,I11529,I11537,I11554,I11571,I71641,I11588,I11605,I11622,I11639,I11373,I11670,I11687,I11704,I71638,I71629,I11358,I11735,I11752,I11769,I11376,I11379,I11814,I11361,I11364,I11859,I11370,I11914,I11931,I121011,I121029,I11948,I121014,I121008,I11965,I11982,I11894,I12013,I121032,I12030,I121023,I12056,I12064,I12081,I12098,I12115,I12132,I12149,I12166,I11900,I12197,I121017,I12214,I12231,I121026,I121020,I11885,I12262,I12279,I12296,I11903,I11906,I12341,I11888,I11891,I12386,I11897,I12441,I12458,I142618,I142636,I12475,I142621,I142615,I12492,I12509,I12421,I12540,I142639,I12557,I142630,I12583,I12591,I12608,I12625,I12642,I12659,I12676,I12693,I12427,I12724,I142624,I12741,I12758,I142633,I142627,I12412,I12789,I12806,I12823,I12430,I12433,I12868,I12415,I12418,I12913,I12424,I12968,I12985,I129443,I129461,I13002,I129446,I129440,I13019,I13036,I12948,I13067,I129464,I13084,I129455,I13110,I13118,I13135,I13152,I13169,I13186,I13203,I13220,I12954,I13251,I129449,I13268,I13285,I129458,I129452,I12939,I13316,I13333,I13350,I12957,I12960,I13395,I12942,I12945,I13440,I12951,I13495,I13512,I39496,I13529,I39517,I39514,I13546,I13563,I13475,I13594,I39493,I39505,I13611,I39502,I13637,I13645,I13662,I13679,I39511,I13696,I13713,I13730,I13747,I13481,I13778,I13795,I13812,I39508,I39499,I13466,I13843,I13860,I13877,I13484,I13487,I13922,I13469,I13472,I13967,I13478,I14025,I14042,I202492,I202495,I14059,I202501,I202489,I14076,I14093,I14110,I14127,I202507,I202510,I14144,I202504,I14170,I14178,I14195,I14212,I14229,I14246,I14005,I14277,I202498,I14294,I14311,I14014,I14017,I14356,I14008,I14002,I14401,I14418,I13996,I13999,I14011,I14477,I13993,I14535,I14552,I388010,I14569,I388025,I388028,I14586,I14603,I14620,I14637,I388016,I388019,I14654,I388013,I14680,I14688,I14705,I14722,I14739,I14756,I14515,I14787,I388022,I14804,I14821,I14524,I14527,I14866,I14518,I14512,I14911,I14928,I14506,I14509,I14521,I14987,I14503,I15045,I15062,I109165,I109159,I15079,I109177,I15096,I15113,I15130,I15147,I109171,I109162,I15164,I15190,I15198,I15215,I109174,I15232,I15249,I15266,I15025,I15297,I109168,I15314,I15331,I15034,I15037,I15376,I15028,I15022,I15421,I15438,I15016,I15019,I15031,I15497,I15013,I15555,I15572,I335758,I335752,I15589,I335761,I335764,I15606,I15623,I15640,I15657,I335755,I15674,I15700,I15708,I15725,I335770,I15742,I15759,I15776,I15535,I15807,I335767,I15824,I335773,I15841,I15544,I15547,I15886,I15538,I15532,I15931,I15948,I15526,I15529,I15541,I16007,I15523,I16065,I16082,I374750,I16099,I374765,I374768,I16116,I16133,I16150,I16167,I374756,I374759,I16184,I374753,I16210,I16218,I16235,I16252,I16269,I16286,I16045,I16317,I374762,I16334,I16351,I16054,I16057,I16396,I16048,I16042,I16441,I16458,I16036,I16039,I16051,I16517,I16033,I16575,I16592,I281032,I281035,I16609,I281041,I281029,I16626,I16643,I16660,I16677,I281047,I281050,I16694,I281044,I16720,I16728,I16745,I16762,I16779,I16796,I16555,I16827,I281038,I16844,I16861,I16564,I16567,I16906,I16558,I16552,I16951,I16968,I16546,I16549,I16561,I17027,I16543,I17085,I17102,I265800,I265803,I17119,I265809,I265797,I17136,I17153,I17170,I17187,I265815,I265818,I17204,I265812,I17230,I17238,I17255,I17272,I17289,I17306,I17065,I17337,I265806,I17354,I17371,I17074,I17077,I17416,I17068,I17062,I17461,I17478,I17056,I17059,I17071,I17537,I17053,I17595,I17612,I17629,I17646,I17663,I17680,I17697,I17714,I17740,I17748,I17765,I17782,I17799,I17816,I17575,I17847,I17864,I17881,I17584,I17587,I17926,I17578,I17572,I17971,I17988,I17566,I17569,I17581,I18047,I17563,I18105,I18122,I228672,I228675,I18139,I228681,I228669,I18156,I18173,I18190,I18207,I228687,I228690,I18224,I228684,I18250,I18258,I18275,I18292,I18309,I18326,I18085,I18357,I228678,I18374,I18391,I18094,I18097,I18436,I18088,I18082,I18481,I18498,I18076,I18079,I18091,I18557,I18073,I18615,I18632,I333123,I333117,I18649,I333126,I333129,I18666,I18683,I18700,I18717,I333120,I18734,I18760,I18768,I18785,I333135,I18802,I18819,I18836,I18867,I333132,I18884,I333138,I18901,I18946,I18991,I19008,I19067,I19125,I19142,I224864,I224867,I19159,I224873,I224861,I19176,I19193,I19210,I19227,I224879,I224882,I19244,I224876,I19270,I19278,I19295,I19312,I19329,I19346,I19105,I19377,I224870,I19394,I19411,I19114,I19117,I19456,I19108,I19102,I19501,I19518,I19096,I19099,I19111,I19577,I19093,I19635,I19652,I331542,I331536,I19669,I331545,I331548,I19686,I19703,I19720,I19737,I331539,I19754,I19780,I19788,I19805,I331554,I19822,I19839,I19856,I19615,I19887,I331551,I19904,I331557,I19921,I19624,I19627,I19966,I19618,I19612,I20011,I20028,I19606,I19609,I19621,I20087,I19603,I20145,I20162,I257232,I257235,I20179,I257241,I257229,I20196,I20213,I20230,I20247,I257247,I257250,I20264,I257244,I20290,I20298,I20315,I20332,I20349,I20366,I20125,I20397,I257238,I20414,I20431,I20134,I20137,I20476,I20128,I20122,I20521,I20538,I20116,I20119,I20131,I20597,I20113,I20655,I20672,I238192,I238195,I20689,I238201,I238189,I20706,I20723,I20740,I20757,I238207,I238210,I20774,I238204,I20800,I20808,I20825,I20842,I20859,I20876,I20635,I20907,I238198,I20924,I20941,I20644,I20647,I20986,I20638,I20632,I21031,I21048,I20626,I20629,I20641,I21107,I20623,I21165,I21182,I331015,I331009,I21199,I331018,I331021,I21216,I21233,I21250,I21267,I331012,I21284,I21310,I21318,I21335,I331027,I21352,I21369,I21386,I21145,I21417,I331024,I21434,I331030,I21451,I21154,I21157,I21496,I21148,I21142,I21541,I21558,I21136,I21139,I21151,I21617,I21133,I21675,I21692,I21709,I21726,I21743,I21760,I21777,I21794,I21820,I21828,I21845,I21862,I21879,I21896,I21655,I21927,I21944,I21961,I21664,I21667,I22006,I21658,I21652,I22051,I22068,I21646,I21649,I21661,I22127,I21643,I22185,I22202,I176894,I176873,I22219,I176882,I176891,I22236,I22253,I22270,I22287,I176888,I22304,I176879,I22330,I22338,I22355,I176870,I22372,I22389,I22406,I22165,I22437,I176885,I22454,I176876,I22471,I22174,I22177,I22516,I22168,I22162,I22561,I22578,I22156,I22159,I22171,I22637,I22153,I22695,I22712,I282460,I282463,I22729,I282469,I282457,I22746,I22763,I22780,I22797,I282475,I282478,I22814,I282472,I22840,I22848,I22865,I22882,I22899,I22916,I22675,I22947,I282466,I22964,I22981,I22684,I22687,I23026,I22678,I22672,I23071,I23088,I22666,I22669,I22681,I23147,I22663,I23205,I23222,I369446,I23239,I369461,I369464,I23256,I23273,I23290,I23307,I369452,I369455,I23324,I369449,I23350,I23358,I23375,I23392,I23409,I23426,I23185,I23457,I369458,I23474,I23491,I23194,I23197,I23536,I23188,I23182,I23581,I23598,I23176,I23179,I23191,I23657,I23173,I23715,I23732,I214392,I214395,I23749,I214401,I214389,I23766,I23783,I23800,I23817,I214407,I214410,I23834,I214404,I23860,I23868,I23885,I23902,I23919,I23936,I23695,I23967,I214398,I23984,I24001,I23704,I23707,I24046,I23698,I23692,I24091,I24108,I23686,I23689,I23701,I24167,I23683,I24225,I24242,I105085,I105079,I24259,I105097,I24276,I24293,I24310,I24327,I105091,I105082,I24344,I24370,I24378,I24395,I105094,I24412,I24429,I24446,I24205,I24477,I105088,I24494,I24511,I24214,I24217,I24556,I24208,I24202,I24601,I24618,I24196,I24199,I24211,I24677,I24193,I24735,I24752,I312043,I312037,I24769,I312046,I312049,I24786,I24803,I24820,I24837,I312040,I24854,I24880,I24888,I24905,I312055,I24922,I24939,I24956,I24715,I24987,I312052,I25004,I312058,I25021,I24724,I24727,I25066,I24718,I24712,I25111,I25128,I24706,I24709,I24721,I25187,I24703,I25245,I25262,I346825,I346819,I25279,I346828,I346831,I25296,I25313,I25330,I25347,I346822,I25364,I25390,I25398,I25415,I346837,I25432,I25449,I25466,I25225,I25497,I346834,I25514,I346840,I25531,I25234,I25237,I25576,I25228,I25222,I25621,I25638,I25216,I25219,I25231,I25697,I25213,I25755,I25772,I126829,I126808,I25789,I126817,I126826,I25806,I25823,I25840,I25857,I126823,I25874,I126814,I25900,I25908,I25925,I126805,I25942,I25959,I25976,I25735,I26007,I126820,I26024,I126811,I26041,I25744,I25747,I26086,I25738,I25732,I26131,I26148,I25726,I25729,I25741,I26207,I25723,I26265,I26282,I189015,I188994,I26299,I189003,I189012,I26316,I26333,I26350,I26367,I189009,I26384,I189000,I26410,I26418,I26435,I188991,I26452,I26469,I26486,I26245,I26517,I189006,I26534,I188997,I26551,I26254,I26257,I26596,I26248,I26242,I26641,I26658,I26236,I26239,I26251,I26717,I26233,I26775,I26792,I107125,I107119,I26809,I107137,I26826,I26843,I26860,I26877,I107131,I107122,I26894,I26920,I26928,I26945,I107134,I26962,I26979,I26996,I26755,I27027,I107128,I27044,I27061,I26764,I26767,I27106,I26758,I26752,I27151,I27168,I26746,I26749,I26761,I27227,I26743,I27285,I27302,I182164,I182143,I27319,I182152,I182161,I27336,I27353,I27370,I27387,I182158,I27404,I182149,I27430,I27438,I27455,I182140,I27472,I27489,I27506,I27265,I27537,I182155,I27554,I182146,I27571,I27274,I27277,I27616,I27268,I27262,I27661,I27678,I27256,I27259,I27271,I27737,I27253,I27795,I27812,I107533,I107527,I27829,I107545,I27846,I27863,I27880,I27897,I107539,I107530,I27914,I27940,I27948,I27965,I107542,I27982,I27999,I28016,I27775,I28047,I107536,I28064,I28081,I27784,I27787,I28126,I27778,I27772,I28171,I28188,I27766,I27769,I27781,I28247,I27763,I28305,I28322,I276748,I276751,I28339,I276757,I276745,I28356,I28373,I28390,I28407,I276763,I276766,I28424,I276760,I28450,I28458,I28475,I28492,I28509,I28526,I28285,I28557,I276754,I28574,I28591,I28294,I28297,I28636,I28288,I28282,I28681,I28698,I28276,I28279,I28291,I28757,I28273,I28815,I28832,I159503,I159482,I28849,I159491,I159500,I28866,I28883,I28900,I28917,I159497,I28934,I159488,I28960,I28968,I28985,I159479,I29002,I29019,I29036,I28795,I29067,I159494,I29084,I159485,I29101,I28804,I28807,I29146,I28798,I28792,I29191,I29208,I28786,I28789,I28801,I29267,I28783,I29325,I29342,I296757,I296754,I29359,I296760,I296772,I29376,I29393,I29410,I29427,I296763,I29444,I296769,I29470,I29478,I29495,I296775,I29512,I29529,I29546,I29305,I29577,I296766,I29594,I29611,I29314,I29317,I29656,I29308,I29302,I29701,I29718,I29296,I29299,I29311,I29777,I29293,I29835,I29852,I361932,I29869,I361947,I361950,I29886,I29903,I29920,I29937,I361938,I361941,I29954,I361935,I29980,I29988,I30005,I30022,I30039,I30056,I29815,I30087,I361944,I30104,I30121,I29824,I29827,I30166,I29818,I29812,I30211,I30228,I29806,I29809,I29821,I30287,I29803,I30345,I30362,I134734,I134713,I30379,I134722,I134731,I30396,I30413,I30430,I30447,I134728,I30464,I134719,I30490,I30498,I30515,I134710,I30532,I30549,I30566,I30325,I30597,I134725,I30614,I134716,I30631,I30334,I30337,I30676,I30328,I30322,I30721,I30738,I30316,I30319,I30331,I30797,I30313,I30855,I30872,I251044,I251047,I30889,I251053,I251041,I30906,I30923,I30940,I30957,I251059,I251062,I30974,I251056,I31000,I31008,I31025,I31042,I31059,I31076,I30835,I31107,I251050,I31124,I31141,I30844,I30847,I31186,I30838,I30832,I31231,I31248,I30826,I30829,I30841,I31307,I30823,I31365,I31382,I170570,I170549,I31399,I170558,I170567,I31416,I31433,I31450,I31467,I170564,I31484,I170555,I31510,I31518,I31535,I170546,I31552,I31569,I31586,I31345,I31617,I170561,I31634,I170552,I31651,I31354,I31357,I31696,I31348,I31342,I31741,I31758,I31336,I31339,I31351,I31817,I31333,I31875,I31892,I161611,I161590,I31909,I161599,I161608,I31926,I31943,I31960,I31977,I161605,I31994,I161596,I32020,I32028,I32045,I161587,I32062,I32079,I32096,I31855,I32127,I161602,I32144,I161593,I32161,I31864,I31867,I32206,I31858,I31852,I32251,I32268,I31846,I31849,I31861,I32327,I31843,I32385,I32402,I161084,I161063,I32419,I161072,I161081,I32436,I32453,I32470,I32487,I161078,I32504,I161069,I32530,I32538,I32555,I161060,I32572,I32589,I32606,I32365,I32637,I161075,I32654,I161066,I32671,I32374,I32377,I32716,I32368,I32362,I32761,I32778,I32356,I32359,I32371,I32837,I32353,I32895,I32912,I402154,I32929,I402169,I402172,I32946,I32963,I32980,I32997,I402160,I402163,I33014,I402157,I33040,I33048,I33065,I33082,I33099,I33116,I32875,I33147,I402166,I33164,I33181,I32884,I32887,I33226,I32878,I32872,I33271,I33288,I32866,I32869,I32881,I33347,I32863,I33405,I33422,I124721,I124700,I33439,I124709,I124718,I33456,I33473,I33490,I33507,I124715,I33524,I124706,I33550,I33558,I33575,I124697,I33592,I33609,I33626,I33385,I33657,I124712,I33674,I124703,I33691,I33394,I33397,I33736,I33388,I33382,I33781,I33798,I33376,I33379,I33391,I33857,I33373,I33915,I33932,I305719,I305713,I33949,I305722,I305725,I33966,I33983,I34000,I34017,I305716,I34034,I34060,I34068,I34085,I305731,I34102,I34119,I34136,I33895,I34167,I305728,I34184,I305734,I34201,I33904,I33907,I34246,I33898,I33892,I34291,I34308,I33886,I33889,I33901,I34367,I33883,I34425,I34442,I370330,I34459,I370345,I370348,I34476,I34493,I34510,I34527,I370336,I370339,I34544,I370333,I34570,I34578,I34595,I34612,I34629,I34646,I34405,I34677,I370342,I34694,I34711,I34414,I34417,I34756,I34408,I34402,I34801,I34818,I34396,I34399,I34411,I34877,I34393,I34935,I34952,I303084,I303078,I34969,I303087,I303090,I34986,I35003,I35020,I35037,I303081,I35054,I35080,I35088,I35105,I303096,I35122,I35139,I35156,I34915,I35187,I303093,I35204,I303099,I35221,I34924,I34927,I35266,I34918,I34912,I35311,I35328,I34906,I34909,I34921,I35387,I34903,I35445,I35462,I212012,I212015,I35479,I212021,I212009,I35496,I35513,I35530,I35547,I212027,I212030,I35564,I212024,I35590,I35598,I35615,I35632,I35649,I35666,I35425,I35697,I212018,I35714,I35731,I35434,I35437,I35776,I35428,I35422,I35821,I35838,I35416,I35419,I35431,I35897,I35413,I35955,I35972,I195866,I195845,I35989,I195854,I195863,I36006,I36023,I36040,I36057,I195860,I36074,I195851,I36100,I36108,I36125,I195842,I36142,I36159,I36176,I35935,I36207,I195857,I36224,I195848,I36241,I35944,I35947,I36286,I35938,I35932,I36331,I36348,I35926,I35929,I35941,I36407,I35923,I36465,I36482,I210584,I210587,I36499,I210593,I210581,I36516,I36533,I36550,I36567,I210599,I210602,I36584,I210596,I36610,I36618,I36635,I36652,I36669,I36686,I36717,I210590,I36734,I36751,I36796,I36841,I36858,I36917,I36975,I36992,I225340,I225343,I37009,I225349,I225337,I37026,I37043,I37060,I37077,I225355,I225358,I37094,I225352,I37120,I37128,I37145,I37162,I37179,I37196,I36955,I37227,I225346,I37244,I37261,I36964,I36967,I37306,I36958,I36952,I37351,I37368,I36946,I36949,I36961,I37427,I36943,I37485,I37502,I175313,I175292,I37519,I175301,I175310,I37536,I37553,I37570,I37587,I175307,I37604,I175298,I37630,I37638,I37655,I175289,I37672,I37689,I37706,I37465,I37737,I175304,I37754,I175295,I37771,I37474,I37477,I37816,I37468,I37462,I37861,I37878,I37456,I37459,I37471,I37937,I37453,I37995,I38012,I402596,I38029,I402611,I402614,I38046,I38063,I38080,I38097,I402602,I402605,I38114,I402599,I38140,I38148,I38165,I38182,I38199,I38216,I37975,I38247,I402608,I38264,I38281,I37984,I37987,I38326,I37978,I37972,I38371,I38388,I37966,I37969,I37981,I38447,I37963,I38505,I38522,I281508,I281511,I38539,I281517,I281505,I38556,I38573,I38590,I38607,I281523,I281526,I38624,I281520,I38650,I38658,I38675,I38692,I38709,I38726,I38757,I281514,I38774,I38791,I38836,I38881,I38898,I38957,I39015,I39032,I407016,I39049,I407031,I407034,I39066,I39083,I39100,I39117,I407022,I407025,I39134,I407019,I39160,I39168,I39185,I39202,I39219,I39236,I38995,I39267,I407028,I39284,I39301,I39004,I39007,I39346,I38998,I38992,I39391,I39408,I38986,I38989,I39001,I39467,I38983,I39525,I39542,I410552,I39559,I410567,I410570,I39576,I39593,I39610,I39627,I410558,I410561,I39644,I410555,I39670,I39678,I39695,I39712,I39729,I39746,I39777,I410564,I39794,I39811,I39856,I39901,I39918,I39977,I40035,I40052,I216296,I216299,I40069,I216305,I216293,I40086,I40103,I40120,I40137,I216311,I216314,I40154,I216308,I40180,I40188,I40205,I40222,I40239,I40256,I40015,I40287,I216302,I40304,I40321,I40024,I40027,I40366,I40018,I40012,I40411,I40428,I40006,I40009,I40021,I40487,I40003,I40545,I40562,I232480,I232483,I40579,I232489,I232477,I40596,I40613,I40630,I40647,I232495,I232498,I40664,I232492,I40690,I40698,I40715,I40732,I40749,I40766,I40525,I40797,I232486,I40814,I40831,I40534,I40537,I40876,I40528,I40522,I40921,I40938,I40516,I40519,I40531,I40997,I40513,I41055,I41072,I163192,I163171,I41089,I163180,I163189,I41106,I41123,I41140,I41157,I163186,I41174,I163177,I41200,I41208,I41225,I163168,I41242,I41259,I41276,I41035,I41307,I163183,I41324,I163174,I41341,I41044,I41047,I41386,I41038,I41032,I41431,I41448,I41026,I41029,I41041,I41507,I41023,I41565,I41582,I368562,I41599,I368577,I368580,I41616,I41633,I41650,I41667,I368568,I368571,I41684,I368565,I41710,I41718,I41735,I41752,I41769,I41786,I41545,I41817,I368574,I41834,I41851,I41554,I41557,I41896,I41548,I41542,I41941,I41958,I41536,I41539,I41551,I42017,I41533,I42075,I42092,I329434,I329428,I42109,I329437,I329440,I42126,I42143,I42160,I42177,I329431,I42194,I42220,I42228,I42245,I329446,I42262,I42279,I42296,I42055,I42327,I329443,I42344,I329449,I42361,I42064,I42067,I42406,I42058,I42052,I42451,I42468,I42046,I42049,I42061,I42527,I42043,I42585,I42602,I186380,I186359,I42619,I186368,I186377,I42636,I42653,I42670,I42687,I186374,I42704,I186365,I42730,I42738,I42755,I186356,I42772,I42789,I42806,I42565,I42837,I186371,I42854,I186362,I42871,I42574,I42577,I42916,I42568,I42562,I42961,I42978,I42556,I42559,I42571,I43037,I42553,I43095,I43112,I43129,I43146,I43163,I43180,I43197,I43214,I43240,I43248,I43265,I43282,I43299,I43316,I43075,I43347,I43364,I43381,I43084,I43087,I43426,I43078,I43072,I43471,I43488,I43066,I43069,I43081,I43547,I43063,I43605,I43622,I248188,I248191,I43639,I248197,I248185,I43656,I43673,I43690,I43707,I248203,I248206,I43724,I248200,I43750,I43758,I43775,I43792,I43809,I43826,I43585,I43857,I248194,I43874,I43891,I43594,I43597,I43936,I43588,I43582,I43981,I43998,I43576,I43579,I43591,I44057,I43573,I44115,I44132,I299919,I299916,I44149,I299922,I299934,I44166,I44183,I44200,I44217,I299925,I44234,I299931,I44260,I44268,I44285,I299937,I44302,I44319,I44336,I44367,I299928,I44384,I44401,I44446,I44491,I44508,I44567,I44625,I44642,I206776,I206779,I44659,I206785,I206773,I44676,I44693,I44710,I44727,I206791,I206794,I44744,I206788,I44770,I44778,I44795,I44812,I44829,I44846,I44605,I44877,I206782,I44894,I44911,I44614,I44617,I44956,I44608,I44602,I45001,I45018,I44596,I44599,I44611,I45077,I44593,I45135,I45152,I201064,I201067,I45169,I201073,I201061,I45186,I45203,I45220,I45237,I201079,I201082,I45254,I201076,I45280,I45288,I45305,I45322,I45339,I45356,I45115,I45387,I201070,I45404,I45421,I45124,I45127,I45466,I45118,I45112,I45511,I45528,I45106,I45109,I45121,I45587,I45103,I45645,I45662,I325745,I325739,I45679,I325748,I325751,I45696,I45713,I45730,I45747,I325742,I45764,I45790,I45798,I45815,I325757,I45832,I45849,I45866,I45897,I325754,I45914,I325760,I45931,I45976,I46021,I46038,I46097,I46155,I46172,I256280,I256283,I46189,I256289,I256277,I46206,I46223,I46240,I46257,I256295,I256298,I46274,I256292,I46300,I46308,I46325,I46342,I46359,I46376,I46135,I46407,I256286,I46424,I46441,I46144,I46147,I46486,I46138,I46132,I46531,I46548,I46126,I46129,I46141,I46607,I46123,I46665,I46682,I383590,I46699,I383605,I383608,I46716,I46733,I46750,I46767,I383596,I383599,I46784,I383593,I46810,I46818,I46835,I46852,I46869,I46886,I46645,I46917,I383602,I46934,I46951,I46654,I46657,I46996,I46648,I46642,I47041,I47058,I46636,I46639,I46651,I47117,I46633,I47175,I47192,I208204,I208207,I47209,I208213,I208201,I47226,I47243,I47260,I47277,I208219,I208222,I47294,I208216,I47320,I47328,I47345,I47362,I47379,I47396,I47155,I47427,I208210,I47444,I47461,I47164,I47167,I47506,I47158,I47152,I47551,I47568,I47146,I47149,I47161,I47627,I47143,I47685,I47702,I268656,I268659,I47719,I268665,I268653,I47736,I47753,I47770,I47787,I268671,I268674,I47804,I268668,I47830,I47838,I47855,I47872,I47889,I47906,I47665,I47937,I268662,I47954,I47971,I47674,I47677,I48016,I47668,I47662,I48061,I48078,I47656,I47659,I47671,I48137,I47653,I48195,I48212,I308354,I308348,I48229,I308357,I308360,I48246,I48263,I48280,I48297,I308351,I48314,I48340,I48348,I48365,I308366,I48382,I48399,I48416,I48175,I48447,I308363,I48464,I308369,I48481,I48184,I48187,I48526,I48178,I48172,I48571,I48588,I48166,I48169,I48181,I48647,I48163,I48705,I48722,I234860,I234863,I48739,I234869,I234857,I48756,I48773,I48790,I48807,I234875,I234878,I48824,I234872,I48850,I48858,I48875,I48892,I48909,I48926,I48685,I48957,I234866,I48974,I48991,I48694,I48697,I49036,I48688,I48682,I49081,I49098,I48676,I48679,I48691,I49157,I48673,I49215,I49232,I208680,I208683,I49249,I208689,I208677,I49266,I49283,I49300,I49317,I208695,I208698,I49334,I208692,I49360,I49368,I49385,I49402,I49419,I49436,I49195,I49467,I208686,I49484,I49501,I49204,I49207,I49546,I49198,I49192,I49591,I49608,I49186,I49189,I49201,I49667,I49183,I49725,I49742,I280556,I280559,I49759,I280565,I280553,I49776,I49793,I49810,I49827,I280571,I280574,I49844,I280568,I49870,I49878,I49895,I49912,I49929,I49946,I49705,I49977,I280562,I49994,I50011,I49714,I49717,I50056,I49708,I49702,I50101,I50118,I49696,I49699,I49711,I50177,I49693,I50235,I50252,I298865,I298862,I50269,I298868,I298880,I50286,I50303,I50320,I50337,I298871,I50354,I298877,I50380,I50388,I50405,I298883,I50422,I50439,I50456,I50215,I50487,I298874,I50504,I50521,I50224,I50227,I50566,I50218,I50212,I50611,I50628,I50206,I50209,I50221,I50687,I50203,I50745,I50762,I105493,I105487,I50779,I105505,I50796,I50813,I50830,I50847,I105499,I105490,I50864,I50890,I50898,I50915,I105502,I50932,I50949,I50966,I50725,I50997,I105496,I51014,I51031,I50734,I50737,I51076,I50728,I50722,I51121,I51138,I50716,I50719,I50731,I51197,I50713,I51255,I51272,I251520,I251523,I51289,I251529,I251517,I51306,I51323,I51340,I51357,I251535,I251538,I51374,I251532,I51400,I51408,I51425,I51442,I51459,I51476,I51235,I51507,I251526,I51524,I51541,I51244,I51247,I51586,I51238,I51232,I51631,I51648,I51226,I51229,I51241,I51707,I51223,I51765,I51782,I336812,I336806,I51799,I336815,I336818,I51816,I51833,I51850,I51867,I336809,I51884,I51910,I51918,I51935,I336824,I51952,I51969,I51986,I51745,I52017,I336821,I52034,I336827,I52051,I51754,I51757,I52096,I51748,I51742,I52141,I52158,I51736,I51739,I51751,I52217,I51733,I52275,I52292,I199555,I199534,I52309,I199543,I199552,I52326,I52343,I52360,I52377,I199549,I52394,I199540,I52420,I52428,I52445,I199531,I52462,I52479,I52496,I52255,I52527,I199546,I52544,I199537,I52561,I52264,I52267,I52606,I52258,I52252,I52651,I52668,I52246,I52249,I52261,I52727,I52243,I52785,I52802,I147909,I147888,I52819,I147897,I147906,I52836,I52853,I52870,I52887,I147903,I52904,I147894,I52930,I52938,I52955,I147885,I52972,I52989,I53006,I52765,I53037,I147900,I53054,I147891,I53071,I52774,I52777,I53116,I52768,I52762,I53161,I53178,I52756,I52759,I52771,I53237,I52753,I53295,I53312,I324691,I324685,I53329,I324694,I324697,I53346,I53363,I53380,I53397,I324688,I53414,I53440,I53448,I53465,I324703,I53482,I53499,I53516,I53275,I53547,I324700,I53564,I324706,I53581,I53284,I53287,I53626,I53278,I53272,I53671,I53688,I53266,I53269,I53281,I53747,I53263,I53805,I53822,I381380,I53839,I381395,I381398,I53856,I53873,I53890,I53907,I381386,I381389,I53924,I381383,I53950,I53958,I53975,I53992,I54009,I54026,I53785,I54057,I381392,I54074,I54091,I53794,I53797,I54136,I53788,I53782,I54181,I54198,I53776,I53779,I53791,I54257,I53773,I54315,I54332,I247712,I247715,I54349,I247721,I247709,I54366,I54383,I54400,I54417,I247727,I247730,I54434,I247724,I54460,I54468,I54485,I54502,I54519,I54536,I54295,I54567,I247718,I54584,I54601,I54304,I54307,I54646,I54298,I54292,I54691,I54708,I54286,I54289,I54301,I54767,I54283,I54825,I54842,I54859,I54876,I54893,I54910,I54927,I54944,I54970,I54978,I54995,I55012,I55029,I55046,I54805,I55077,I55094,I55111,I54814,I54817,I55156,I54808,I54802,I55201,I55218,I54796,I54799,I54811,I55277,I54793,I55335,I55352,I217248,I217251,I55369,I217257,I217245,I55386,I55403,I55420,I55437,I217263,I217266,I55454,I217260,I55480,I55488,I55505,I55522,I55539,I55556,I55315,I55587,I217254,I55604,I55621,I55324,I55327,I55666,I55318,I55312,I55711,I55728,I55306,I55309,I55321,I55787,I55303,I55845,I55862,I230576,I230579,I55879,I230585,I230573,I55896,I55913,I55930,I55947,I230591,I230594,I55964,I230588,I55990,I55998,I56015,I56032,I56049,I56066,I55825,I56097,I230582,I56114,I56131,I55834,I55837,I56176,I55828,I55822,I56221,I56238,I55816,I55819,I55831,I56297,I55813,I56355,I56372,I191123,I191102,I56389,I191111,I191120,I56406,I56423,I56440,I56457,I191117,I56474,I191108,I56500,I56508,I56525,I191099,I56542,I56559,I56576,I56335,I56607,I191114,I56624,I191105,I56641,I56344,I56347,I56686,I56338,I56332,I56731,I56748,I56326,I56329,I56341,I56807,I56323,I56865,I56882,I121559,I121538,I56899,I121547,I121556,I56916,I56933,I56950,I56967,I121553,I56984,I121544,I57010,I57018,I57035,I121535,I57052,I57069,I57086,I56845,I57117,I121550,I57134,I121541,I57151,I56854,I56857,I57196,I56848,I56842,I57241,I57258,I56836,I56839,I56851,I57317,I56833,I57375,I57392,I341028,I341022,I57409,I341031,I341034,I57426,I57443,I57460,I57477,I341025,I57494,I57520,I57528,I57545,I341040,I57562,I57579,I57596,I57355,I57627,I341037,I57644,I341043,I57661,I57364,I57367,I57706,I57358,I57352,I57751,I57768,I57346,I57349,I57361,I57827,I57343,I57885,I57902,I379170,I57919,I379185,I379188,I57936,I57953,I57970,I57987,I379176,I379179,I58004,I379173,I58030,I58038,I58055,I58072,I58089,I58106,I57865,I58137,I379182,I58154,I58171,I57874,I57877,I58216,I57868,I57862,I58261,I58278,I57856,I57859,I57871,I58337,I57853,I58395,I58412,I233908,I233911,I58429,I233917,I233905,I58446,I58463,I58480,I58497,I233923,I233926,I58514,I233920,I58540,I58548,I58565,I58582,I58599,I58616,I58375,I58647,I233914,I58664,I58681,I58384,I58387,I58726,I58378,I58372,I58771,I58788,I58366,I58369,I58381,I58847,I58363,I58905,I58922,I260564,I260567,I58939,I260573,I260561,I58956,I58973,I58990,I59007,I260579,I260582,I59024,I260576,I59050,I59058,I59075,I59092,I59109,I59126,I58885,I59157,I260570,I59174,I59191,I58894,I58897,I59236,I58888,I58882,I59281,I59298,I58876,I58879,I58891,I59357,I58873,I59415,I59432,I131045,I131024,I59449,I131033,I131042,I59466,I59483,I59500,I59517,I131039,I59534,I131030,I59560,I59568,I59585,I131021,I59602,I59619,I59636,I59395,I59667,I131036,I59684,I131027,I59701,I59404,I59407,I59746,I59398,I59392,I59791,I59808,I59386,I59389,I59401,I59867,I59383,I59925,I59942,I215820,I215823,I59959,I215829,I215817,I59976,I59993,I60010,I60027,I215835,I215838,I60044,I215832,I60070,I60078,I60095,I60112,I60129,I60146,I59905,I60177,I215826,I60194,I60211,I59914,I59917,I60256,I59908,I59902,I60301,I60318,I59896,I59899,I59911,I60377,I59893,I60435,I60452,I250568,I250571,I60469,I250577,I250565,I60486,I60503,I60520,I60537,I250583,I250586,I60554,I250580,I60580,I60588,I60605,I60622,I60639,I60656,I60415,I60687,I250574,I60704,I60721,I60424,I60427,I60766,I60418,I60412,I60811,I60828,I60406,I60409,I60421,I60887,I60403,I60945,I60962,I60979,I60996,I61013,I61030,I61047,I61064,I61090,I61098,I61115,I61132,I61149,I61166,I60925,I61197,I61214,I61231,I60934,I60937,I61276,I60928,I60922,I61321,I61338,I60916,I60919,I60931,I61397,I60913,I61455,I61472,I61489,I61506,I61523,I61540,I61557,I61574,I61600,I61608,I61625,I61642,I61659,I61676,I61435,I61707,I61724,I61741,I61444,I61447,I61786,I61438,I61432,I61831,I61848,I61426,I61429,I61441,I61907,I61423,I61965,I61982,I126302,I126281,I61999,I126290,I126299,I62016,I62033,I62050,I62067,I126296,I62084,I126287,I62110,I62118,I62135,I126278,I62152,I62169,I62186,I61945,I62217,I126293,I62234,I126284,I62251,I61954,I61957,I62296,I61948,I61942,I62341,I62358,I61936,I61939,I61951,I62417,I61933,I62475,I62492,I116101,I116095,I62509,I116113,I62526,I62543,I62560,I62577,I116107,I116098,I62594,I62620,I62628,I62645,I116110,I62662,I62679,I62696,I62455,I62727,I116104,I62744,I62761,I62464,I62467,I62806,I62458,I62452,I62851,I62868,I62446,I62449,I62461,I62927,I62443,I62985,I63002,I155814,I155793,I63019,I155802,I155811,I63036,I63053,I63070,I63087,I155808,I63104,I155799,I63130,I63138,I63155,I155790,I63172,I63189,I63206,I62965,I63237,I155805,I63254,I155796,I63271,I62974,I62977,I63316,I62968,I62962,I63361,I63378,I62956,I62959,I62971,I63437,I62953,I63495,I63512,I261516,I261519,I63529,I261525,I261513,I63546,I63563,I63580,I63597,I261531,I261534,I63614,I261528,I63640,I63648,I63665,I63682,I63699,I63716,I63475,I63747,I261522,I63764,I63781,I63484,I63487,I63826,I63478,I63472,I63871,I63888,I63466,I63469,I63481,I63947,I63463,I64005,I64022,I395966,I64039,I395981,I395984,I64056,I64073,I64090,I64107,I395972,I395975,I64124,I395969,I64150,I64158,I64175,I64192,I64209,I64226,I63985,I64257,I395978,I64274,I64291,I63994,I63997,I64336,I63988,I63982,I64381,I64398,I63976,I63979,I63991,I64457,I63973,I64515,I64532,I251996,I251999,I64549,I252005,I251993,I64566,I64583,I64600,I64617,I252011,I252014,I64634,I252008,I64660,I64668,I64685,I64702,I64719,I64736,I64767,I252002,I64784,I64801,I64846,I64891,I64908,I64967,I65025,I65042,I394640,I65059,I394655,I394658,I65076,I65093,I65110,I65127,I394646,I394649,I65144,I394643,I65170,I65178,I65195,I65212,I65229,I65246,I65005,I65277,I394652,I65294,I65311,I65014,I65017,I65356,I65008,I65002,I65401,I65418,I64996,I64999,I65011,I65477,I64993,I65535,I65552,I304138,I304132,I65569,I304141,I304144,I65586,I65603,I65620,I65637,I304135,I65654,I65680,I65688,I65705,I304150,I65722,I65739,I65756,I65515,I65787,I304147,I65804,I304153,I65821,I65524,I65527,I65866,I65518,I65512,I65911,I65928,I65506,I65509,I65521,I65987,I65503,I66045,I66062,I408342,I66079,I408357,I408360,I66096,I66113,I66130,I66147,I408348,I408351,I66164,I408345,I66190,I66198,I66215,I66232,I66249,I66266,I66025,I66297,I408354,I66314,I66331,I66034,I66037,I66376,I66028,I66022,I66421,I66438,I66016,I66019,I66031,I66497,I66013,I66555,I66572,I117343,I117322,I66589,I117331,I117340,I66606,I66623,I66640,I66657,I117337,I66674,I117328,I66700,I66708,I66725,I117319,I66742,I66759,I66776,I66535,I66807,I117334,I66824,I117325,I66841,I66544,I66547,I66886,I66538,I66532,I66931,I66948,I66526,I66529,I66541,I67007,I66523,I67065,I67082,I114877,I114871,I67099,I114889,I67116,I67133,I67150,I67167,I114883,I114874,I67184,I67210,I67218,I67235,I114886,I67252,I67269,I67286,I67045,I67317,I114880,I67334,I67351,I67054,I67057,I67396,I67048,I67042,I67441,I67458,I67036,I67039,I67051,I67517,I67033,I67575,I67592,I192177,I192156,I67609,I192165,I192174,I67626,I67643,I67660,I67677,I192171,I67694,I192162,I67720,I67728,I67745,I192153,I67762,I67779,I67796,I67555,I67827,I192168,I67844,I192159,I67861,I67564,I67567,I67906,I67558,I67552,I67951,I67968,I67546,I67549,I67561,I68027,I67543,I68085,I68102,I230100,I230103,I68119,I230109,I230097,I68136,I68153,I68170,I68187,I230115,I230118,I68204,I230112,I68230,I68238,I68255,I68272,I68289,I68306,I68065,I68337,I230106,I68354,I68371,I68074,I68077,I68416,I68068,I68062,I68461,I68478,I68056,I68059,I68071,I68537,I68053,I68595,I68612,I221532,I221535,I68629,I221541,I221529,I68646,I68663,I68680,I68697,I221547,I221550,I68714,I221544,I68740,I68748,I68765,I68782,I68799,I68816,I68575,I68847,I221538,I68864,I68881,I68584,I68587,I68926,I68578,I68572,I68971,I68988,I68566,I68569,I68581,I69047,I68563,I69105,I69122,I162665,I162644,I69139,I162653,I162662,I69156,I69173,I69190,I69207,I162659,I69224,I162650,I69250,I69258,I69275,I162641,I69292,I69309,I69326,I69085,I69357,I162656,I69374,I162647,I69391,I69094,I69097,I69436,I69088,I69082,I69481,I69498,I69076,I69079,I69091,I69557,I69073,I69615,I69632,I231052,I231055,I69649,I231061,I231049,I69666,I69683,I69700,I69717,I231067,I231070,I69734,I231064,I69760,I69768,I69785,I69802,I69819,I69836,I69595,I69867,I231058,I69884,I69901,I69604,I69607,I69946,I69598,I69592,I69991,I70008,I69586,I69589,I69601,I70067,I69583,I70125,I70142,I148436,I148415,I70159,I148424,I148433,I70176,I70193,I70210,I70227,I148430,I70244,I148421,I70270,I70278,I70295,I148412,I70312,I70329,I70346,I70105,I70377,I148427,I70394,I148418,I70411,I70114,I70117,I70456,I70108,I70102,I70501,I70518,I70096,I70099,I70111,I70577,I70093,I70635,I70652,I168989,I168968,I70669,I168977,I168986,I70686,I70703,I70720,I70737,I168983,I70754,I168974,I70780,I70788,I70805,I168965,I70822,I70839,I70856,I70615,I70887,I168980,I70904,I168971,I70921,I70624,I70627,I70966,I70618,I70612,I71011,I71028,I70606,I70609,I70621,I71087,I70603,I71145,I71162,I71179,I71196,I71213,I71230,I71247,I71264,I71290,I71298,I71315,I71332,I71349,I71366,I71125,I71397,I71414,I71431,I71134,I71137,I71476,I71128,I71122,I71521,I71538,I71116,I71119,I71131,I71597,I71113,I71655,I71672,I183218,I183197,I71689,I183206,I183215,I71706,I71723,I71740,I71757,I183212,I71774,I183203,I71800,I71808,I71825,I183194,I71842,I71859,I71876,I71907,I183209,I71924,I183200,I71941,I71986,I72031,I72048,I72107,I72165,I72182,I342609,I342603,I72199,I342612,I342615,I72216,I72233,I72250,I72267,I342606,I72284,I72310,I72318,I72335,I342621,I72352,I72369,I72386,I72145,I72417,I342618,I72434,I342624,I72451,I72154,I72157,I72496,I72148,I72142,I72541,I72558,I72136,I72139,I72151,I72617,I72133,I72675,I72692,I177948,I177927,I72709,I177936,I177945,I72726,I72743,I72760,I72777,I177942,I72794,I177933,I72820,I72828,I72845,I177924,I72862,I72879,I72896,I72655,I72927,I177939,I72944,I177930,I72961,I72664,I72667,I73006,I72658,I72652,I73051,I73068,I72646,I72649,I72661,I73127,I72643,I73185,I73202,I317840,I317834,I73219,I317843,I317846,I73236,I73253,I73270,I73287,I317837,I73304,I73330,I73338,I73355,I317852,I73372,I73389,I73406,I73165,I73437,I317849,I73454,I317855,I73471,I73174,I73177,I73516,I73168,I73162,I73561,I73578,I73156,I73159,I73171,I73637,I73153,I73695,I73712,I294649,I294646,I73729,I294652,I294664,I73746,I73763,I73780,I73797,I294655,I73814,I294661,I73840,I73848,I73865,I294667,I73882,I73899,I73916,I73675,I73947,I294658,I73964,I73981,I73684,I73687,I74026,I73678,I73672,I74071,I74088,I73666,I73669,I73681,I74147,I73663,I74205,I74222,I261040,I261043,I74239,I261049,I261037,I74256,I74273,I74290,I74307,I261055,I261058,I74324,I261052,I74350,I74358,I74375,I74392,I74409,I74426,I74185,I74457,I261046,I74474,I74491,I74194,I74197,I74536,I74188,I74182,I74581,I74598,I74176,I74179,I74191,I74657,I74173,I74715,I74732,I268180,I268183,I74749,I268189,I268177,I74766,I74783,I74800,I74817,I268195,I268198,I74834,I268192,I74860,I74868,I74885,I74902,I74919,I74936,I74695,I74967,I268186,I74984,I75001,I74704,I74707,I75046,I74698,I74692,I75091,I75108,I74686,I74689,I74701,I75167,I74683,I75225,I75242,I202968,I202971,I75259,I202977,I202965,I75276,I75293,I75310,I75327,I202983,I202986,I75344,I202980,I75370,I75378,I75395,I75412,I75429,I75446,I75205,I75477,I202974,I75494,I75511,I75214,I75217,I75556,I75208,I75202,I75601,I75618,I75196,I75199,I75211,I75677,I75193,I75735,I75752,I120505,I120484,I75769,I120493,I120502,I75786,I75803,I75820,I75837,I120499,I75854,I120490,I75880,I75888,I75905,I120481,I75922,I75939,I75956,I75715,I75987,I120496,I76004,I120487,I76021,I75724,I75727,I76066,I75718,I75712,I76111,I76128,I75706,I75709,I75721,I76187,I75703,I76245,I76262,I152652,I152631,I76279,I152640,I152649,I76296,I76313,I76330,I76347,I152646,I76364,I152637,I76390,I76398,I76415,I152628,I76432,I76449,I76466,I76225,I76497,I152643,I76514,I152634,I76531,I76234,I76237,I76576,I76228,I76222,I76621,I76638,I76216,I76219,I76231,I76697,I76213,I76755,I76772,I267704,I267707,I76789,I267713,I267701,I76806,I76823,I76840,I76857,I267719,I267722,I76874,I267716,I76900,I76908,I76925,I76942,I76959,I76976,I76735,I77007,I267710,I77024,I77041,I76744,I76747,I77086,I76738,I76732,I77131,I77148,I76726,I76729,I76741,I77207,I76723,I77265,I77282,I290433,I290430,I77299,I290436,I290448,I77316,I77333,I77350,I77367,I290439,I77384,I290445,I77410,I77418,I77435,I290451,I77452,I77469,I77486,I77245,I77517,I290442,I77534,I77551,I77254,I77257,I77596,I77248,I77242,I77641,I77658,I77236,I77239,I77251,I77717,I77233,I77775,I77792,I196393,I196372,I77809,I196381,I196390,I77826,I77843,I77860,I77877,I196387,I77894,I196378,I77920,I77928,I77945,I196369,I77962,I77979,I77996,I77755,I78027,I196384,I78044,I196375,I78061,I77764,I77767,I78106,I77758,I77752,I78151,I78168,I77746,I77749,I77761,I78227,I77743,I78285,I78302,I215344,I215347,I78319,I215353,I215341,I78336,I78353,I78370,I78387,I215359,I215362,I78404,I215356,I78430,I78438,I78455,I78472,I78489,I78506,I78265,I78537,I215350,I78554,I78571,I78274,I78277,I78616,I78268,I78262,I78661,I78678,I78256,I78259,I78271,I78737,I78253,I78795,I78812,I166881,I166860,I78829,I166869,I166878,I78846,I78863,I78880,I78897,I166875,I78914,I166866,I78940,I78948,I78965,I166857,I78982,I78999,I79016,I78775,I79047,I166872,I79064,I166863,I79081,I78784,I78787,I79126,I78778,I78772,I79171,I79188,I78766,I78769,I78781,I79247,I78763,I79305,I79322,I384916,I79339,I384931,I384934,I79356,I79373,I79390,I79407,I384922,I384925,I79424,I384919,I79450,I79458,I79475,I79492,I79509,I79526,I79285,I79557,I384928,I79574,I79591,I79294,I79297,I79636,I79288,I79282,I79681,I79698,I79276,I79279,I79291,I79757,I79273,I79815,I79832,I156868,I156847,I79849,I156856,I156865,I79866,I79883,I79900,I79917,I156862,I79934,I156853,I79960,I79968,I79985,I156844,I80002,I80019,I80036,I79795,I80067,I156859,I80084,I156850,I80101,I79804,I79807,I80146,I79798,I79792,I80191,I80208,I79786,I79789,I79801,I80267,I79783,I80325,I80342,I393314,I80359,I393329,I393332,I80376,I80393,I80410,I80427,I393320,I393323,I80444,I393317,I80470,I80478,I80495,I80512,I80529,I80546,I80305,I80577,I393326,I80594,I80611,I80314,I80317,I80656,I80308,I80302,I80701,I80718,I80296,I80299,I80311,I80777,I80293,I80835,I80852,I313624,I313618,I80869,I313627,I313630,I80886,I80903,I80920,I80937,I313621,I80954,I80980,I80988,I81005,I313636,I81022,I81039,I81056,I80815,I81087,I313633,I81104,I313639,I81121,I80824,I80827,I81166,I80818,I80812,I81211,I81228,I80806,I80809,I80821,I81287,I80803,I81345,I81362,I333650,I333644,I81379,I333653,I333656,I81396,I81413,I81430,I81447,I333647,I81464,I81490,I81498,I81515,I333662,I81532,I81549,I81566,I81325,I81597,I333659,I81614,I333665,I81631,I81334,I81337,I81676,I81328,I81322,I81721,I81738,I81316,I81319,I81331,I81797,I81313,I81855,I81872,I160030,I160009,I81889,I160018,I160027,I81906,I81923,I81940,I81957,I160024,I81974,I160015,I82000,I82008,I82025,I160006,I82042,I82059,I82076,I81835,I82107,I160021,I82124,I160012,I82141,I81844,I81847,I82186,I81838,I81832,I82231,I82248,I81826,I81829,I81841,I82307,I81823,I82365,I82382,I307300,I307294,I82399,I307303,I307306,I82416,I82433,I82450,I82467,I307297,I82484,I82510,I82518,I82535,I307312,I82552,I82569,I82586,I82617,I307309,I82634,I307315,I82651,I82696,I82741,I82758,I82817,I82875,I82892,I315205,I315199,I82909,I315208,I315211,I82926,I82943,I82960,I82977,I315202,I82994,I83020,I83028,I83045,I315217,I83062,I83079,I83096,I82855,I83127,I315214,I83144,I315220,I83161,I82864,I82867,I83206,I82858,I82852,I83251,I83268,I82846,I82849,I82861,I83327,I82843,I83385,I83402,I185853,I185832,I83419,I185841,I185850,I83436,I83453,I83470,I83487,I185847,I83504,I185838,I83530,I83538,I83555,I185829,I83572,I83589,I83606,I83365,I83637,I185844,I83654,I185835,I83671,I83374,I83377,I83716,I83368,I83362,I83761,I83778,I83356,I83359,I83371,I83837,I83353,I83895,I83912,I360527,I360521,I83929,I360530,I360533,I83946,I83963,I83980,I83997,I360524,I84014,I84040,I84048,I84065,I360539,I84082,I84099,I84116,I83875,I84147,I360536,I84164,I360542,I84181,I83884,I83887,I84226,I83878,I83872,I84271,I84288,I83866,I83869,I83881,I84347,I83863,I84405,I84422,I276272,I276275,I84439,I276281,I276269,I84456,I84473,I84490,I84507,I276287,I276290,I84524,I276284,I84550,I84558,I84575,I84592,I84609,I84626,I84385,I84657,I276278,I84674,I84691,I84394,I84397,I84736,I84388,I84382,I84781,I84798,I84376,I84379,I84391,I84857,I84373,I84915,I84932,I245332,I245335,I84949,I245341,I245329,I84966,I84983,I85000,I85017,I245347,I245350,I85034,I245344,I85060,I85068,I85085,I85102,I85119,I85136,I84895,I85167,I245338,I85184,I85201,I84904,I84907,I85246,I84898,I84892,I85291,I85308,I84886,I84889,I84901,I85367,I84883,I85425,I85442,I135261,I135240,I85459,I135249,I135258,I85476,I85493,I85510,I85527,I135255,I85544,I135246,I85570,I85578,I85595,I135237,I85612,I85629,I85646,I85405,I85677,I135252,I85694,I135243,I85711,I85414,I85417,I85756,I85408,I85402,I85801,I85818,I85396,I85399,I85411,I85877,I85393,I85935,I85952,I193231,I193210,I85969,I193219,I193228,I85986,I86003,I86020,I86037,I193225,I86054,I193216,I86080,I86088,I86105,I193207,I86122,I86139,I86156,I85915,I86187,I193222,I86204,I193213,I86221,I85924,I85927,I86266,I85918,I85912,I86311,I86328,I85906,I85909,I85921,I86387,I85903,I86445,I86462,I380496,I86479,I380511,I380514,I86496,I86513,I86530,I86547,I380502,I380505,I86564,I380499,I86590,I86598,I86615,I86632,I86649,I86666,I86425,I86697,I380508,I86714,I86731,I86434,I86437,I86776,I86428,I86422,I86821,I86838,I86416,I86419,I86431,I86897,I86413,I86955,I86972,I117870,I117849,I86989,I117858,I117867,I87006,I87023,I87040,I87057,I117864,I87074,I117855,I87100,I87108,I87125,I117846,I87142,I87159,I87176,I86935,I87207,I117861,I87224,I117852,I87241,I86944,I86947,I87286,I86938,I86932,I87331,I87348,I86926,I86929,I86941,I87407,I86923,I87465,I87482,I209156,I209159,I87499,I209165,I209153,I87516,I87533,I87550,I87567,I209171,I209174,I87584,I209168,I87610,I87618,I87635,I87652,I87669,I87686,I87445,I87717,I209162,I87734,I87751,I87454,I87457,I87796,I87448,I87442,I87841,I87858,I87436,I87439,I87451,I87917,I87433,I87975,I87992,I375192,I88009,I375207,I375210,I88026,I88043,I88060,I88077,I375198,I375201,I88094,I375195,I88120,I88128,I88145,I88162,I88179,I88196,I87955,I88227,I375204,I88244,I88261,I87964,I87967,I88306,I87958,I87952,I88351,I88368,I87946,I87949,I87961,I88427,I87943,I88485,I88502,I283888,I283891,I88519,I283897,I283885,I88536,I88553,I88570,I88587,I283903,I283906,I88604,I283900,I88630,I88638,I88655,I88672,I88689,I88706,I88465,I88737,I283894,I88754,I88771,I88474,I88477,I88816,I88468,I88462,I88861,I88878,I88456,I88459,I88471,I88937,I88453,I88995,I89012,I372540,I89029,I372555,I372558,I89046,I89063,I89080,I89097,I372546,I372549,I89114,I372543,I89140,I89148,I89165,I89182,I89199,I89216,I88975,I89247,I372552,I89264,I89281,I88984,I88987,I89326,I88978,I88972,I89371,I89388,I88966,I88969,I88981,I89447,I88963,I89505,I89522,I114061,I114055,I89539,I114073,I89556,I89573,I89590,I89607,I114067,I114058,I89624,I89650,I89658,I89675,I114070,I89692,I89709,I89726,I89485,I89757,I114064,I89774,I89791,I89494,I89497,I89836,I89488,I89482,I89881,I89898,I89476,I89479,I89491,I89957,I89473,I90015,I90032,I275796,I275799,I90049,I275805,I275793,I90066,I90083,I90100,I90117,I275811,I275814,I90134,I275808,I90160,I90168,I90185,I90202,I90219,I90236,I90267,I275802,I90284,I90301,I90346,I90391,I90408,I90467,I90525,I90542,I143166,I143145,I90559,I143154,I143163,I90576,I90593,I90610,I90627,I143160,I90644,I143151,I90670,I90678,I90695,I143142,I90712,I90729,I90746,I90505,I90777,I143157,I90794,I143148,I90811,I90514,I90517,I90856,I90508,I90502,I90901,I90918,I90496,I90499,I90511,I90977,I90493,I91035,I91052,I214868,I214871,I91069,I214877,I214865,I91086,I91103,I91120,I91137,I214883,I214886,I91154,I214880,I91180,I91188,I91205,I91222,I91239,I91256,I91015,I91287,I214874,I91304,I91321,I91024,I91027,I91366,I91018,I91012,I91411,I91428,I91006,I91009,I91021,I91487,I91003,I91545,I91562,I129991,I129970,I91579,I129979,I129988,I91596,I91613,I91630,I91647,I129985,I91664,I129976,I91690,I91698,I91715,I129967,I91732,I91749,I91766,I91525,I91797,I129982,I91814,I129973,I91831,I91534,I91537,I91876,I91528,I91522,I91921,I91938,I91516,I91519,I91531,I91997,I91513,I92055,I92072,I128410,I128389,I92089,I128398,I128407,I92106,I92123,I92140,I92157,I128404,I92174,I128395,I92200,I92208,I92225,I128386,I92242,I92259,I92276,I92035,I92307,I128401,I92324,I128392,I92341,I92044,I92047,I92386,I92038,I92032,I92431,I92448,I92026,I92029,I92041,I92507,I92023,I92565,I92582,I319948,I319942,I92599,I319951,I319954,I92616,I92633,I92650,I92667,I319945,I92684,I92710,I92718,I92735,I319960,I92752,I92769,I92786,I92545,I92817,I319957,I92834,I319963,I92851,I92554,I92557,I92896,I92548,I92542,I92941,I92958,I92536,I92539,I92551,I93017,I92533,I93075,I93092,I372098,I93109,I372113,I372116,I93126,I93143,I93160,I93177,I372104,I372107,I93194,I372101,I93220,I93228,I93245,I93262,I93279,I93296,I93055,I93327,I372110,I93344,I93361,I93064,I93067,I93406,I93058,I93052,I93451,I93468,I93046,I93049,I93061,I93527,I93043,I93585,I93602,I397292,I93619,I397307,I397310,I93636,I93653,I93670,I93687,I397298,I397301,I93704,I397295,I93730,I93738,I93755,I93772,I93789,I93806,I93565,I93837,I397304,I93854,I93871,I93574,I93577,I93916,I93568,I93562,I93961,I93978,I93556,I93559,I93571,I94037,I93553,I94095,I94112,I393756,I94129,I393771,I393774,I94146,I94163,I94180,I94197,I393762,I393765,I94214,I393759,I94240,I94248,I94265,I94282,I94299,I94316,I94075,I94347,I393768,I94364,I94381,I94084,I94087,I94426,I94078,I94072,I94471,I94488,I94066,I94069,I94081,I94547,I94063,I94605,I94622,I246760,I246763,I94639,I246769,I246757,I94656,I94673,I94690,I94707,I246775,I246778,I94724,I246772,I94750,I94758,I94775,I94792,I94809,I94826,I94585,I94857,I246766,I94874,I94891,I94594,I94597,I94936,I94588,I94582,I94981,I94998,I94576,I94579,I94591,I95057,I94573,I95115,I95132,I313097,I313091,I95149,I313100,I313103,I95166,I95183,I95200,I95217,I313094,I95234,I95260,I95268,I95285,I313109,I95302,I95319,I95336,I95095,I95367,I313106,I95384,I313112,I95401,I95104,I95107,I95446,I95098,I95092,I95491,I95508,I95086,I95089,I95101,I95567,I95083,I95625,I95642,I167408,I167387,I95659,I167396,I167405,I95676,I95693,I95710,I95727,I167402,I95744,I167393,I95770,I95778,I95795,I167384,I95812,I95829,I95846,I95605,I95877,I167399,I95894,I167390,I95911,I95614,I95617,I95956,I95608,I95602,I96001,I96018,I95596,I95599,I95611,I96077,I95593,I96135,I96152,I353149,I353143,I96169,I353152,I353155,I96186,I96203,I96220,I96237,I353146,I96254,I96280,I96288,I96305,I353161,I96322,I96339,I96356,I96115,I96387,I353158,I96404,I353164,I96421,I96124,I96127,I96466,I96118,I96112,I96511,I96528,I96106,I96109,I96121,I96587,I96103,I96645,I96662,I118397,I118376,I96679,I118385,I118394,I96696,I96713,I96730,I96747,I118391,I96764,I118382,I96790,I96798,I96815,I118373,I96832,I96849,I96866,I96625,I96897,I118388,I96914,I118379,I96931,I96634,I96637,I96976,I96628,I96622,I97021,I97038,I96616,I96619,I96631,I97097,I96613,I97155,I97172,I396408,I97189,I396423,I396426,I97206,I97223,I97240,I97257,I396414,I396417,I97274,I396411,I97300,I97308,I97325,I97342,I97359,I97376,I97135,I97407,I396420,I97424,I97441,I97144,I97147,I97486,I97138,I97132,I97531,I97548,I97126,I97129,I97141,I97607,I97123,I97665,I97682,I133153,I133132,I97699,I133141,I133150,I97716,I97733,I97750,I97767,I133147,I97784,I133138,I97810,I97818,I97835,I133129,I97852,I97869,I97886,I97645,I97917,I133144,I97934,I133135,I97951,I97654,I97657,I97996,I97648,I97642,I98041,I98058,I97636,I97639,I97651,I98117,I97633,I98175,I98192,I178475,I178454,I98209,I178463,I178472,I98226,I98243,I98260,I98277,I178469,I98294,I178460,I98320,I98328,I98345,I178451,I98362,I98379,I98396,I98155,I98427,I178466,I98444,I178457,I98461,I98164,I98167,I98506,I98158,I98152,I98551,I98568,I98146,I98149,I98161,I98627,I98143,I98685,I98702,I213440,I213443,I98719,I213449,I213437,I98736,I98753,I98770,I98787,I213455,I213458,I98804,I213452,I98830,I98838,I98855,I98872,I98889,I98906,I98665,I98937,I213446,I98954,I98971,I98674,I98677,I99016,I98668,I98662,I99061,I99078,I98656,I98659,I98671,I99137,I98653,I99195,I99212,I166354,I166333,I99229,I166342,I166351,I99246,I99263,I99280,I99297,I166348,I99314,I166339,I99340,I99348,I99365,I166330,I99382,I99399,I99416,I99175,I99447,I166345,I99464,I166336,I99481,I99184,I99187,I99526,I99178,I99172,I99571,I99588,I99166,I99169,I99181,I99647,I99163,I99705,I99722,I170043,I170022,I99739,I170031,I170040,I99756,I99773,I99790,I99807,I170037,I99824,I170028,I99850,I99858,I99875,I170019,I99892,I99909,I99926,I99685,I99957,I170034,I99974,I170025,I99991,I99694,I99697,I100036,I99688,I99682,I100081,I100098,I99676,I99679,I99691,I100157,I99673,I100215,I100232,I205824,I205827,I100249,I205833,I205821,I100266,I100283,I100300,I100317,I205839,I205842,I100334,I205836,I100360,I100368,I100385,I100402,I100419,I100436,I100195,I100467,I205830,I100484,I100501,I100204,I100207,I100546,I100198,I100192,I100591,I100608,I100186,I100189,I100201,I100667,I100183,I100725,I100742,I380938,I100759,I380953,I380956,I100776,I100793,I100810,I100827,I380944,I380947,I100844,I380941,I100870,I100878,I100895,I100912,I100929,I100946,I100705,I100977,I380950,I100994,I101011,I100714,I100717,I101056,I100708,I100702,I101101,I101118,I100696,I100699,I100711,I101177,I100693,I101235,I101252,I270560,I270563,I101269,I270569,I270557,I101286,I101303,I101320,I101337,I270575,I270578,I101354,I270572,I101380,I101388,I101405,I101422,I101439,I101456,I101215,I101487,I270566,I101504,I101521,I101224,I101227,I101566,I101218,I101212,I101611,I101628,I101206,I101209,I101221,I101687,I101203,I101745,I101762,I315732,I315726,I101779,I315735,I315738,I101796,I101813,I101830,I101847,I315729,I101864,I101890,I101898,I101915,I315744,I101932,I101949,I101966,I101725,I101997,I315741,I102014,I315747,I102031,I101734,I101737,I102076,I101728,I101722,I102121,I102138,I101716,I101719,I101731,I102197,I101713,I102249,I102266,I180053,I180035,I102283,I180056,I102300,I180032,I180047,I102317,I102223,I102348,I102365,I102382,I180050,I102399,I180038,I102416,I102238,I102447,I180044,I102464,I180041,I102481,I102241,I102226,I102526,I102543,I102560,I102577,I102229,I102235,I102232,I102657,I102674,I240093,I102691,I240114,I102708,I240096,I240099,I102725,I102631,I102756,I102773,I102790,I240102,I240111,I102807,I240108,I102824,I102646,I102855,I102872,I240105,I102889,I102649,I102634,I102934,I102951,I102968,I102985,I102637,I102643,I102640,I103065,I103082,I269605,I103099,I269626,I103116,I269608,I269611,I103133,I103039,I103164,I103181,I103198,I269614,I269623,I103215,I269620,I103232,I103054,I103263,I103280,I269617,I103297,I103057,I103042,I103342,I103359,I103376,I103393,I103045,I103051,I103048,I103473,I103490,I223909,I103507,I223930,I103524,I223912,I223915,I103541,I103447,I103572,I103589,I103606,I223918,I223927,I103623,I223924,I103640,I103462,I103671,I103688,I223921,I103705,I103465,I103450,I103750,I103767,I103784,I103801,I103453,I103459,I103456,I103881,I103898,I178999,I178981,I103915,I179002,I103932,I178978,I178993,I103949,I103855,I103980,I103997,I104014,I178996,I104031,I178984,I104048,I103870,I104079,I178990,I104096,I178987,I104113,I103873,I103858,I104158,I104175,I104192,I104209,I103861,I103867,I103864,I104289,I104306,I104323,I104340,I104357,I104263,I104388,I104405,I104422,I104439,I104456,I104278,I104487,I104504,I104521,I104281,I104266,I104566,I104583,I104600,I104617,I104269,I104275,I104272,I104697,I104714,I289388,I289397,I104731,I289379,I104748,I289394,I289382,I104765,I104671,I104796,I104813,I104830,I289376,I104847,I104864,I104686,I104895,I104912,I289385,I289391,I104929,I104689,I104674,I104974,I104991,I105008,I105025,I104677,I104683,I104680,I105105,I105122,I388909,I388903,I105139,I388906,I105156,I388900,I105173,I105204,I105221,I105238,I388897,I388894,I105255,I105272,I105303,I105320,I388912,I105337,I105382,I105399,I105416,I105433,I105513,I105530,I405705,I405699,I105547,I405702,I105564,I405696,I105581,I105612,I105629,I105646,I405693,I405690,I105663,I105680,I105711,I105728,I405708,I105745,I105790,I105807,I105824,I105841,I105921,I105938,I345256,I345241,I105955,I345244,I105972,I345238,I345253,I105989,I105895,I106020,I106037,I106054,I106071,I106088,I105910,I106119,I345259,I106136,I345250,I345247,I106153,I105913,I105898,I106198,I106215,I106232,I106249,I105901,I105907,I105904,I106329,I106346,I378743,I378737,I106363,I378740,I106380,I378734,I106397,I106303,I106428,I106445,I106462,I378731,I378728,I106479,I106496,I106318,I106527,I106544,I378746,I106561,I106321,I106306,I106606,I106623,I106640,I106657,I106309,I106315,I106312,I106737,I106754,I350526,I350511,I106771,I350514,I106788,I350508,I350523,I106805,I106711,I106836,I106853,I106870,I106887,I106904,I106726,I106935,I350529,I106952,I350520,I350517,I106969,I106729,I106714,I107014,I107031,I107048,I107065,I106717,I106723,I106720,I107145,I107162,I309420,I309405,I107179,I309408,I107196,I309402,I309417,I107213,I107244,I107261,I107278,I107295,I107312,I107343,I309423,I107360,I309414,I309411,I107377,I107422,I107439,I107456,I107473,I107553,I107570,I323649,I323634,I107587,I323637,I107604,I323631,I323646,I107621,I107652,I107669,I107686,I107703,I107720,I107751,I323652,I107768,I323643,I323640,I107785,I107830,I107847,I107864,I107881,I107961,I107978,I292550,I292559,I107995,I292541,I108012,I292556,I292544,I108029,I107935,I108060,I108077,I108094,I292538,I108111,I108128,I107950,I108159,I108176,I292547,I292553,I108193,I107953,I107938,I108238,I108255,I108272,I108289,I107941,I107947,I107944,I108369,I108386,I192701,I192683,I108403,I192704,I108420,I192680,I192695,I108437,I108343,I108468,I108485,I108502,I192698,I108519,I192686,I108536,I108358,I108567,I192692,I108584,I192689,I108601,I108361,I108346,I108646,I108663,I108680,I108697,I108349,I108355,I108352,I108777,I108794,I235333,I108811,I235354,I108828,I235336,I235339,I108845,I108751,I108876,I108893,I108910,I235342,I235351,I108927,I235348,I108944,I108766,I108975,I108992,I235345,I109009,I108769,I108754,I109054,I109071,I109088,I109105,I108757,I108763,I108760,I109185,I109202,I109219,I109236,I109253,I109284,I109301,I109318,I109335,I109352,I109383,I109400,I109417,I109462,I109479,I109496,I109513,I109593,I109610,I109627,I109644,I109661,I109567,I109692,I109709,I109726,I109743,I109760,I109582,I109791,I109808,I109825,I109585,I109570,I109870,I109887,I109904,I109921,I109573,I109579,I109576,I110001,I110018,I356323,I356308,I110035,I356311,I110052,I356305,I356320,I110069,I109975,I110100,I110117,I110134,I110151,I110168,I109990,I110199,I356326,I110216,I356317,I356314,I110233,I109993,I109978,I110278,I110295,I110312,I110329,I109981,I109987,I109984,I110409,I110426,I195336,I195318,I110443,I195339,I110460,I195315,I195330,I110477,I110383,I110508,I110525,I110542,I195333,I110559,I195321,I110576,I110398,I110607,I195327,I110624,I195324,I110641,I110401,I110386,I110686,I110703,I110720,I110737,I110389,I110395,I110392,I110817,I110834,I171094,I171076,I110851,I171097,I110868,I171073,I171088,I110885,I110791,I110916,I110933,I110950,I171091,I110967,I171079,I110984,I110806,I111015,I171085,I111032,I171082,I111049,I110809,I110794,I111094,I111111,I111128,I111145,I110797,I110803,I110800,I111225,I111242,I311528,I311513,I111259,I311516,I111276,I311510,I311525,I111293,I111199,I111324,I111341,I111358,I111375,I111392,I111214,I111423,I311531,I111440,I311522,I311519,I111457,I111217,I111202,I111502,I111519,I111536,I111553,I111205,I111211,I111208,I111633,I111650,I111667,I111684,I111701,I111607,I111732,I111749,I111766,I111783,I111800,I111622,I111831,I111848,I111865,I111625,I111610,I111910,I111927,I111944,I111961,I111613,I111619,I111616,I112041,I112058,I145271,I145253,I112075,I145274,I112092,I145250,I145265,I112109,I112015,I112140,I112157,I112174,I145268,I112191,I145256,I112208,I112030,I112239,I145262,I112256,I145259,I112273,I112033,I112018,I112318,I112335,I112352,I112369,I112021,I112027,I112024,I112449,I112466,I137366,I137348,I112483,I137369,I112500,I137345,I137360,I112517,I112423,I112548,I112565,I112582,I137363,I112599,I137351,I112616,I112438,I112647,I137357,I112664,I137354,I112681,I112441,I112426,I112726,I112743,I112760,I112777,I112429,I112435,I112432,I112857,I112874,I395097,I395091,I112891,I395094,I112908,I395088,I112925,I112831,I112956,I112973,I112990,I395085,I395082,I113007,I113024,I112846,I113055,I113072,I395100,I113089,I112849,I112834,I113134,I113151,I113168,I113185,I112837,I112843,I112840,I113265,I113282,I125772,I125754,I113299,I125775,I113316,I125751,I125766,I113333,I113239,I113364,I113381,I113398,I125769,I113415,I125757,I113432,I113254,I113463,I125763,I113480,I125760,I113497,I113257,I113242,I113542,I113559,I113576,I113593,I113245,I113251,I113248,I113673,I113690,I113707,I113724,I113741,I113647,I113772,I113789,I113806,I113823,I113840,I113662,I113871,I113888,I113905,I113665,I113650,I113950,I113967,I113984,I114001,I113653,I113659,I113656,I114081,I114098,I366809,I366803,I114115,I366806,I114132,I366800,I114149,I114180,I114197,I114214,I366797,I366794,I114231,I114248,I114279,I114296,I366812,I114313,I114358,I114375,I114392,I114409,I114489,I114506,I253897,I114523,I253918,I114540,I253900,I253903,I114557,I114463,I114588,I114605,I114622,I253906,I253915,I114639,I253912,I114656,I114478,I114687,I114704,I253909,I114721,I114481,I114466,I114766,I114783,I114800,I114817,I114469,I114475,I114472,I114897,I114914,I249137,I114931,I249158,I114948,I249140,I249143,I114965,I114996,I115013,I115030,I249146,I249155,I115047,I249152,I115064,I115095,I115112,I249149,I115129,I115174,I115191,I115208,I115225,I115305,I115322,I137893,I137875,I115339,I137896,I115356,I137872,I137887,I115373,I115279,I115404,I115421,I115438,I137890,I115455,I137878,I115472,I115294,I115503,I137884,I115520,I137881,I115537,I115297,I115282,I115582,I115599,I115616,I115633,I115285,I115291,I115288,I115713,I115730,I115747,I115764,I115781,I115687,I115812,I115829,I115846,I115863,I115880,I115702,I115911,I115928,I115945,I115705,I115690,I115990,I116007,I116024,I116041,I115693,I115699,I115696,I116121,I116138,I274365,I116155,I274386,I116172,I274368,I274371,I116189,I116220,I116237,I116254,I274374,I274383,I116271,I274380,I116288,I116319,I116336,I274377,I116353,I116398,I116415,I116432,I116449,I116529,I116546,I116563,I116580,I116597,I116503,I116628,I116645,I116662,I116679,I116696,I116518,I116727,I116744,I116761,I116521,I116506,I116806,I116823,I116840,I116857,I116509,I116515,I116512,I116937,I116954,I144744,I144726,I116971,I144747,I116988,I144723,I144738,I117005,I116911,I117036,I117053,I117070,I144741,I117087,I144729,I117104,I116926,I117135,I144735,I117152,I144732,I117169,I116929,I116914,I117214,I117231,I117248,I117265,I116917,I116923,I116920,I117351,I117368,I322595,I322583,I117385,I322577,I117402,I117419,I117436,I117453,I322580,I117470,I322586,I117496,I117518,I117535,I117566,I322592,I117583,I117614,I322598,I117631,I117648,I322589,I117679,I117696,I117727,I117758,I117789,I117820,I117878,I117895,I363264,I363261,I117912,I363273,I363276,I117929,I117946,I117963,I117980,I363267,I363258,I117997,I118023,I118045,I118062,I118093,I118110,I118141,I118158,I118175,I363270,I118206,I118223,I118254,I118285,I118316,I118347,I118405,I118422,I118439,I118456,I118473,I118490,I118507,I118524,I118550,I118572,I118589,I118620,I118637,I118668,I118685,I118702,I118733,I118750,I118781,I118812,I118843,I118874,I118932,I118949,I233429,I233432,I118966,I233435,I233444,I118983,I119000,I119017,I119034,I233441,I233447,I119051,I119077,I118900,I119099,I119116,I118918,I119147,I119164,I118921,I119195,I233450,I119212,I119229,I233438,I118903,I119260,I119277,I118924,I119308,I118909,I119339,I118912,I119370,I118906,I119401,I118915,I119459,I119476,I244377,I244380,I119493,I244383,I244392,I119510,I119527,I119544,I119561,I244389,I244395,I119578,I119604,I119427,I119626,I119643,I119445,I119674,I119691,I119448,I119722,I244398,I119739,I119756,I244386,I119430,I119787,I119804,I119451,I119835,I119436,I119866,I119439,I119897,I119433,I119928,I119442,I119986,I120003,I348945,I348933,I120020,I348927,I120037,I120054,I120071,I120088,I348930,I120105,I348936,I120131,I119954,I120153,I120170,I119972,I120201,I348942,I120218,I119975,I120249,I348948,I120266,I120283,I348939,I119957,I120314,I120331,I119978,I120362,I119963,I120393,I119966,I120424,I119960,I120455,I119969,I120513,I120530,I120547,I120564,I120581,I120598,I120615,I120632,I120658,I120680,I120697,I120728,I120745,I120776,I120793,I120810,I120841,I120858,I120889,I120920,I120951,I120982,I121040,I121057,I121074,I121091,I121108,I121125,I121142,I121159,I121185,I121207,I121224,I121255,I121272,I121303,I121320,I121337,I121368,I121385,I121416,I121447,I121478,I121509,I121567,I121584,I203441,I203444,I121601,I203447,I203456,I121618,I121635,I121652,I121669,I203453,I203459,I121686,I121712,I121734,I121751,I121782,I121799,I121830,I203462,I121847,I121864,I203450,I121895,I121912,I121943,I121974,I122005,I122036,I122094,I122111,I358958,I358946,I122128,I358940,I122145,I122162,I122179,I122196,I358943,I122213,I358949,I122239,I122062,I122261,I122278,I122080,I122309,I358955,I122326,I122083,I122357,I358961,I122374,I122391,I358952,I122065,I122422,I122439,I122086,I122470,I122071,I122501,I122074,I122532,I122068,I122563,I122077,I122621,I122638,I238665,I238668,I122655,I238671,I238680,I122672,I122689,I122706,I122723,I238677,I238683,I122740,I122766,I122589,I122788,I122805,I122607,I122836,I122853,I122610,I122884,I238686,I122901,I122918,I238674,I122592,I122949,I122966,I122613,I122997,I122598,I123028,I122601,I123059,I122595,I123090,I122604,I123148,I123165,I355269,I355257,I123182,I355251,I123199,I123216,I123233,I123250,I355254,I123267,I355260,I123293,I123116,I123315,I123332,I123134,I123363,I355266,I123380,I123137,I123411,I355272,I123428,I123445,I355263,I123119,I123476,I123493,I123140,I123524,I123125,I123555,I123128,I123586,I123122,I123617,I123131,I123675,I123692,I123709,I123726,I123743,I123760,I123777,I123794,I123820,I123643,I123842,I123859,I123661,I123890,I123907,I123664,I123938,I123955,I123972,I123646,I124003,I124020,I123667,I124051,I123652,I124082,I123655,I124113,I123649,I124144,I123658,I124202,I124219,I227717,I227720,I124236,I227723,I227732,I124253,I124270,I124287,I124304,I227729,I227735,I124321,I124347,I124170,I124369,I124386,I124188,I124417,I124434,I124191,I124465,I227738,I124482,I124499,I227726,I124173,I124530,I124547,I124194,I124578,I124179,I124609,I124182,I124640,I124176,I124671,I124185,I124729,I124746,I124763,I124780,I124797,I124814,I124831,I124848,I124874,I124896,I124913,I124944,I124961,I124992,I125009,I125026,I125057,I125074,I125105,I125136,I125167,I125198,I125256,I125273,I377408,I377405,I125290,I377417,I377420,I125307,I125324,I125341,I125358,I377411,I377402,I125375,I125401,I125224,I125423,I125440,I125242,I125471,I125488,I125245,I125519,I125536,I125553,I377414,I125227,I125584,I125601,I125248,I125632,I125233,I125663,I125236,I125694,I125230,I125725,I125239,I125783,I125800,I244853,I244856,I125817,I244859,I244868,I125834,I125851,I125868,I125885,I244865,I244871,I125902,I125928,I125950,I125967,I125998,I126015,I126046,I244874,I126063,I126080,I244862,I126111,I126128,I126159,I126190,I126221,I126252,I126310,I126327,I126344,I126361,I126378,I126395,I126412,I126429,I126455,I126477,I126494,I126525,I126542,I126573,I126590,I126607,I126638,I126655,I126686,I126717,I126748,I126779,I126837,I126854,I249613,I249616,I126871,I249619,I249628,I126888,I126905,I126922,I126939,I249625,I249631,I126956,I126982,I127004,I127021,I127052,I127069,I127100,I249634,I127117,I127134,I249622,I127165,I127182,I127213,I127244,I127275,I127306,I127364,I127381,I127398,I127415,I127432,I127449,I127466,I127483,I127509,I127332,I127531,I127548,I127350,I127579,I127596,I127353,I127627,I127644,I127661,I127335,I127692,I127709,I127356,I127740,I127341,I127771,I127344,I127802,I127338,I127833,I127347,I127891,I127908,I383154,I383151,I127925,I383163,I383166,I127942,I127959,I127976,I127993,I383157,I383148,I128010,I128036,I127859,I128058,I128075,I127877,I128106,I128123,I127880,I128154,I128171,I128188,I383160,I127862,I128219,I128236,I127883,I128267,I127868,I128298,I127871,I128329,I127865,I128360,I127874,I128418,I128435,I128452,I128469,I128486,I128503,I128520,I128537,I128563,I128585,I128602,I128633,I128650,I128681,I128698,I128715,I128746,I128763,I128794,I128825,I128856,I128887,I128945,I128962,I128979,I128996,I129013,I129030,I129047,I129064,I129090,I128913,I129112,I129129,I128931,I129160,I129177,I128934,I129208,I129225,I129242,I128916,I129273,I129290,I128937,I129321,I128922,I129352,I128925,I129383,I128919,I129414,I128928,I129472,I129489,I322068,I322056,I129506,I322050,I129523,I129540,I129557,I129574,I322053,I129591,I322059,I129617,I129639,I129656,I129687,I322065,I129704,I129735,I322071,I129752,I129769,I322062,I129800,I129817,I129848,I129879,I129910,I129941,I129999,I130016,I130033,I130050,I130067,I130084,I130101,I130118,I130144,I130166,I130183,I130214,I130231,I130262,I130279,I130296,I130327,I130344,I130375,I130406,I130437,I130468,I130526,I130543,I130560,I130577,I130594,I130611,I130628,I130645,I130671,I130494,I130693,I130710,I130512,I130741,I130758,I130515,I130789,I130806,I130823,I130497,I130854,I130871,I130518,I130902,I130503,I130933,I130506,I130964,I130500,I130995,I130509,I131053,I131070,I229145,I229148,I131087,I229151,I229160,I131104,I131121,I131138,I131155,I229157,I229163,I131172,I131198,I131220,I131237,I131268,I131285,I131316,I229166,I131333,I131350,I229154,I131381,I131398,I131429,I131460,I131491,I131522,I131580,I131597,I385806,I385803,I131614,I385815,I385818,I131631,I131648,I131665,I131682,I385809,I385800,I131699,I131725,I131548,I131747,I131764,I131566,I131795,I131812,I131569,I131843,I131860,I131877,I385812,I131551,I131908,I131925,I131572,I131956,I131557,I131987,I131560,I132018,I131554,I132049,I131563,I132107,I132124,I334716,I334704,I132141,I334698,I132158,I132175,I132192,I132209,I334701,I132226,I334707,I132252,I132075,I132274,I132291,I132093,I132322,I334713,I132339,I132096,I132370,I334719,I132387,I132404,I334710,I132078,I132435,I132452,I132099,I132483,I132084,I132514,I132087,I132545,I132081,I132576,I132090,I132634,I132651,I231525,I231528,I132668,I231531,I231540,I132685,I132702,I132719,I132736,I231537,I231543,I132753,I132779,I132602,I132801,I132818,I132620,I132849,I132866,I132623,I132897,I231546,I132914,I132931,I231534,I132605,I132962,I132979,I132626,I133010,I132611,I133041,I132614,I133072,I132608,I133103,I132617,I133161,I133178,I218197,I218200,I133195,I218203,I218212,I133212,I133229,I133246,I133263,I218209,I218215,I133280,I133306,I133328,I133345,I133376,I133393,I133424,I218218,I133441,I133458,I218206,I133489,I133506,I133537,I133568,I133599,I133630,I133688,I133705,I212961,I212964,I133722,I212967,I212976,I133739,I133756,I133773,I133790,I212973,I212979,I133807,I133833,I133656,I133855,I133872,I133674,I133903,I133920,I133677,I133951,I212982,I133968,I133985,I212970,I133659,I134016,I134033,I133680,I134064,I133665,I134095,I133668,I134126,I133662,I134157,I133671,I134215,I134232,I222957,I222960,I134249,I222963,I222972,I134266,I134283,I134300,I134317,I222969,I222975,I134334,I134360,I134382,I134399,I134430,I134447,I134478,I222978,I134495,I134512,I222966,I134543,I134560,I134591,I134622,I134653,I134684,I134742,I134759,I304677,I304665,I134776,I304659,I134793,I134810,I134827,I134844,I304662,I134861,I304668,I134887,I134909,I134926,I134957,I304674,I134974,I135005,I304680,I135022,I135039,I304671,I135070,I135087,I135118,I135149,I135180,I135211,I135269,I135286,I135303,I135320,I135337,I135354,I135371,I135388,I135414,I135436,I135453,I135484,I135501,I135532,I135549,I135566,I135597,I135614,I135645,I135676,I135707,I135738,I135796,I135813,I135830,I135847,I135864,I135881,I135898,I135915,I135941,I135764,I135963,I135980,I135782,I136011,I136028,I135785,I136059,I136076,I136093,I135767,I136124,I136141,I135788,I136172,I135773,I136203,I135776,I136234,I135770,I136265,I135779,I136323,I136340,I362380,I362377,I136357,I362389,I362392,I136374,I136391,I136408,I136425,I362383,I362374,I136442,I136468,I136291,I136490,I136507,I136309,I136538,I136555,I136312,I136586,I136603,I136620,I362386,I136294,I136651,I136668,I136315,I136699,I136300,I136730,I136303,I136761,I136297,I136792,I136306,I136850,I136867,I406580,I406577,I136884,I406589,I406592,I136901,I136918,I136935,I136952,I406583,I406574,I136969,I136995,I136818,I137017,I137034,I136836,I137065,I137082,I136839,I137113,I137130,I137147,I406586,I136821,I137178,I137195,I136842,I137226,I136827,I137257,I136830,I137288,I136824,I137319,I136833,I137377,I137394,I137411,I137428,I137445,I137462,I137479,I137496,I137522,I137544,I137561,I137592,I137609,I137640,I137657,I137674,I137705,I137722,I137753,I137784,I137815,I137846,I137904,I137921,I137938,I137955,I137972,I137989,I138006,I138023,I138049,I138071,I138088,I138119,I138136,I138167,I138184,I138201,I138232,I138249,I138280,I138311,I138342,I138373,I138431,I138448,I138465,I138482,I138499,I138516,I138533,I138550,I138576,I138399,I138598,I138615,I138417,I138646,I138663,I138420,I138694,I138711,I138728,I138402,I138759,I138776,I138423,I138807,I138408,I138838,I138411,I138869,I138405,I138900,I138414,I138958,I138975,I255325,I255328,I138992,I255331,I255340,I139009,I139026,I139043,I139060,I255337,I255343,I139077,I139103,I138926,I139125,I139142,I138944,I139173,I139190,I138947,I139221,I255346,I139238,I139255,I255334,I138929,I139286,I139303,I138950,I139334,I138935,I139365,I138938,I139396,I138932,I139427,I138941,I139485,I139502,I205345,I205348,I139519,I205351,I205360,I139536,I139553,I139570,I139587,I205357,I205363,I139604,I139630,I139453,I139652,I139669,I139471,I139700,I139717,I139474,I139748,I205366,I139765,I139782,I205354,I139456,I139813,I139830,I139477,I139861,I139462,I139892,I139465,I139923,I139459,I139954,I139468,I140012,I140029,I140046,I140063,I140080,I140097,I140114,I140131,I140157,I139980,I140179,I140196,I139998,I140227,I140244,I140001,I140275,I140292,I140309,I139983,I140340,I140357,I140004,I140388,I139989,I140419,I139992,I140450,I139986,I140481,I139995,I140539,I140556,I140573,I140590,I140607,I140624,I140641,I140658,I140684,I140507,I140706,I140723,I140525,I140754,I140771,I140528,I140802,I140819,I140836,I140510,I140867,I140884,I140531,I140915,I140516,I140946,I140519,I140977,I140513,I141008,I140522,I141066,I141083,I294140,I294128,I141100,I294131,I294125,I141117,I141134,I141151,I141168,I294122,I141185,I294119,I141211,I141034,I141233,I141250,I141052,I141281,I141298,I141055,I141329,I141346,I141363,I294137,I294134,I141037,I141394,I141411,I141058,I141442,I141043,I141473,I141046,I141504,I141040,I141535,I141049,I141593,I141610,I227241,I227244,I141627,I227247,I227256,I141644,I141661,I141678,I141695,I227253,I227259,I141712,I141738,I141561,I141760,I141777,I141579,I141808,I141825,I141582,I141856,I227262,I141873,I141890,I227250,I141564,I141921,I141938,I141585,I141969,I141570,I142000,I141573,I142031,I141567,I142062,I141576,I142120,I142137,I309947,I309935,I142154,I309929,I142171,I142188,I142205,I142222,I309932,I142239,I309938,I142265,I142088,I142287,I142304,I142106,I142335,I309944,I142352,I142109,I142383,I309950,I142400,I142417,I309941,I142091,I142448,I142465,I142112,I142496,I142097,I142527,I142100,I142558,I142094,I142589,I142103,I142647,I142664,I142681,I142698,I142715,I142732,I142749,I142766,I142792,I142814,I142831,I142862,I142879,I142910,I142927,I142944,I142975,I142992,I143023,I143054,I143085,I143116,I143174,I143191,I143208,I143225,I143242,I143259,I143276,I143293,I143319,I143341,I143358,I143389,I143406,I143437,I143454,I143471,I143502,I143519,I143550,I143581,I143612,I143643,I143701,I143718,I143735,I143752,I143769,I143786,I143803,I143820,I143846,I143669,I143868,I143885,I143687,I143916,I143933,I143690,I143964,I143981,I143998,I143672,I144029,I144046,I143693,I144077,I143678,I144108,I143681,I144139,I143675,I144170,I143684,I144228,I144245,I353688,I353676,I144262,I353670,I144279,I144296,I144313,I144330,I353673,I144347,I353679,I144373,I144196,I144395,I144412,I144214,I144443,I353685,I144460,I144217,I144491,I353691,I144508,I144525,I353682,I144199,I144556,I144573,I144220,I144604,I144205,I144635,I144208,I144666,I144202,I144697,I144211,I144755,I144772,I204869,I204872,I144789,I204875,I204884,I144806,I144823,I144840,I144857,I204881,I204887,I144874,I144900,I144922,I144939,I144970,I144987,I145018,I204890,I145035,I145052,I204878,I145083,I145100,I145131,I145162,I145193,I145224,I145282,I145299,I282933,I282936,I145316,I282939,I282948,I145333,I145350,I145367,I145384,I282945,I282951,I145401,I145427,I145449,I145466,I145497,I145514,I145545,I282954,I145562,I145579,I282942,I145610,I145627,I145658,I145689,I145720,I145751,I145809,I145826,I299410,I299398,I145843,I299401,I299395,I145860,I145877,I145894,I145911,I299392,I145928,I299389,I145954,I145976,I145993,I146024,I146041,I146072,I146089,I146106,I299407,I299404,I146137,I146154,I146185,I146216,I146247,I146278,I146336,I146353,I146370,I146387,I146404,I146421,I146438,I146455,I146481,I146304,I146503,I146520,I146322,I146551,I146568,I146325,I146599,I146616,I146633,I146307,I146664,I146681,I146328,I146712,I146313,I146743,I146316,I146774,I146310,I146805,I146319,I146863,I146880,I258657,I258660,I146897,I258663,I258672,I146914,I146931,I146948,I146965,I258669,I258675,I146982,I147008,I146831,I147030,I147047,I146849,I147078,I147095,I146852,I147126,I258678,I147143,I147160,I258666,I146834,I147191,I147208,I146855,I147239,I146840,I147270,I146843,I147301,I146837,I147332,I146846,I147390,I147407,I147424,I147441,I147458,I147475,I147492,I147509,I147535,I147358,I147557,I147574,I147376,I147605,I147622,I147379,I147653,I147670,I147687,I147361,I147718,I147735,I147382,I147766,I147367,I147797,I147370,I147828,I147364,I147859,I147373,I147917,I147934,I147951,I147968,I147985,I148002,I148019,I148036,I148062,I148084,I148101,I148132,I148149,I148180,I148197,I148214,I148245,I148262,I148293,I148324,I148355,I148386,I148444,I148461,I148478,I148495,I148512,I148529,I148546,I148563,I148589,I148611,I148628,I148659,I148676,I148707,I148724,I148741,I148772,I148789,I148820,I148851,I148882,I148913,I148971,I148988,I200585,I200588,I149005,I200591,I200600,I149022,I149039,I149056,I149073,I200597,I200603,I149090,I149116,I148939,I149138,I149155,I148957,I149186,I149203,I148960,I149234,I200606,I149251,I149268,I200594,I148942,I149299,I149316,I148963,I149347,I148948,I149378,I148951,I149409,I148945,I149440,I148954,I149498,I149515,I387132,I387129,I149532,I387141,I387144,I149549,I149566,I149583,I149600,I387135,I387126,I149617,I149643,I149466,I149665,I149682,I149484,I149713,I149730,I149487,I149761,I149778,I149795,I387138,I149469,I149826,I149843,I149490,I149874,I149475,I149905,I149478,I149936,I149472,I149967,I149481,I150025,I150042,I150059,I150076,I150093,I150110,I150127,I150144,I150170,I149993,I150192,I150209,I150011,I150240,I150257,I150014,I150288,I150305,I150322,I149996,I150353,I150370,I150017,I150401,I150002,I150432,I150005,I150463,I149999,I150494,I150008,I150552,I150569,I382270,I382267,I150586,I382279,I382282,I150603,I150620,I150637,I150654,I382273,I382264,I150671,I150697,I150520,I150719,I150736,I150538,I150767,I150784,I150541,I150815,I150832,I150849,I382276,I150523,I150880,I150897,I150544,I150928,I150529,I150959,I150532,I150990,I150526,I151021,I150535,I151079,I151096,I151113,I151130,I151147,I151164,I151181,I151198,I151224,I151047,I151246,I151263,I151065,I151294,I151311,I151068,I151342,I151359,I151376,I151050,I151407,I151424,I151071,I151455,I151056,I151486,I151059,I151517,I151053,I151548,I151062,I151606,I151623,I151640,I151657,I151674,I151691,I151708,I151725,I151751,I151574,I151773,I151790,I151592,I151821,I151838,I151595,I151869,I151886,I151903,I151577,I151934,I151951,I151598,I151982,I151583,I152013,I151586,I152044,I151580,I152075,I151589,I152133,I152150,I403928,I403925,I152167,I403937,I403940,I152184,I152201,I152218,I152235,I403931,I403922,I152252,I152278,I152101,I152300,I152317,I152119,I152348,I152365,I152122,I152396,I152413,I152430,I403934,I152104,I152461,I152478,I152125,I152509,I152110,I152540,I152113,I152571,I152107,I152602,I152116,I152660,I152677,I306258,I306246,I152694,I306240,I152711,I152728,I152745,I152762,I306243,I152779,I306249,I152805,I152827,I152844,I152875,I306255,I152892,I152923,I306261,I152940,I152957,I306252,I152988,I153005,I153036,I153067,I153098,I153129,I153187,I153204,I302045,I302033,I153221,I302036,I302030,I153238,I153255,I153272,I153289,I302027,I153306,I302024,I153332,I153155,I153354,I153371,I153173,I153402,I153419,I153176,I153450,I153467,I153484,I302042,I302039,I153158,I153515,I153532,I153179,I153563,I153164,I153594,I153167,I153625,I153161,I153656,I153170,I153714,I153731,I153748,I153765,I153782,I153799,I153816,I153833,I153859,I153682,I153881,I153898,I153700,I153929,I153946,I153703,I153977,I153994,I154011,I153685,I154042,I154059,I153706,I154090,I153691,I154121,I153694,I154152,I153688,I154183,I153697,I154241,I154258,I154275,I154292,I154309,I154326,I154343,I154360,I154386,I154209,I154408,I154425,I154227,I154456,I154473,I154230,I154504,I154521,I154538,I154212,I154569,I154586,I154233,I154617,I154218,I154648,I154221,I154679,I154215,I154710,I154224,I154768,I154785,I154802,I154819,I154836,I154853,I154870,I154887,I154913,I154736,I154935,I154952,I154754,I154983,I155000,I154757,I155031,I155048,I155065,I154739,I155096,I155113,I154760,I155144,I154745,I155175,I154748,I155206,I154742,I155237,I154751,I155295,I155312,I155329,I155346,I155363,I155380,I155397,I155414,I155440,I155263,I155462,I155479,I155281,I155510,I155527,I155284,I155558,I155575,I155592,I155266,I155623,I155640,I155287,I155671,I155272,I155702,I155275,I155733,I155269,I155764,I155278,I155822,I155839,I278173,I278176,I155856,I278179,I278188,I155873,I155890,I155907,I155924,I278185,I278191,I155941,I155967,I155989,I156006,I156037,I156054,I156085,I278194,I156102,I156119,I278182,I156150,I156167,I156198,I156229,I156260,I156291,I156349,I156366,I367684,I367681,I156383,I367693,I367696,I156400,I156417,I156434,I156451,I367687,I367678,I156468,I156494,I156317,I156516,I156533,I156335,I156564,I156581,I156338,I156612,I156629,I156646,I367690,I156320,I156677,I156694,I156341,I156725,I156326,I156756,I156329,I156787,I156323,I156818,I156332,I156876,I156893,I254849,I254852,I156910,I254855,I254864,I156927,I156944,I156961,I156978,I254861,I254867,I156995,I157021,I157043,I157060,I157091,I157108,I157139,I254870,I157156,I157173,I254858,I157204,I157221,I157252,I157283,I157314,I157345,I157403,I157420,I225813,I225816,I157437,I225819,I225828,I157454,I157471,I157488,I157505,I225825,I225831,I157522,I157548,I157371,I157570,I157587,I157389,I157618,I157635,I157392,I157666,I225834,I157683,I157700,I225822,I157374,I157731,I157748,I157395,I157779,I157380,I157810,I157383,I157841,I157377,I157872,I157386,I157930,I157947,I376082,I376079,I157964,I376091,I376094,I157981,I157998,I158015,I158032,I376085,I376076,I158049,I158075,I157898,I158097,I158114,I157916,I158145,I158162,I157919,I158193,I158210,I158227,I376088,I157901,I158258,I158275,I157922,I158306,I157907,I158337,I157910,I158368,I157904,I158399,I157913,I158457,I158474,I158491,I158508,I158525,I158542,I158559,I158576,I158602,I158425,I158624,I158641,I158443,I158672,I158689,I158446,I158720,I158737,I158754,I158428,I158785,I158802,I158449,I158833,I158434,I158864,I158437,I158895,I158431,I158926,I158440,I158984,I159001,I366358,I366355,I159018,I366367,I366370,I159035,I159052,I159069,I159086,I366361,I366352,I159103,I159129,I158952,I159151,I159168,I158970,I159199,I159216,I158973,I159247,I159264,I159281,I366364,I158955,I159312,I159329,I158976,I159360,I158961,I159391,I158964,I159422,I158958,I159453,I158967,I159511,I159528,I303623,I303611,I159545,I303605,I159562,I159579,I159596,I159613,I303608,I159630,I303614,I159656,I159678,I159695,I159726,I303620,I159743,I159774,I303626,I159791,I159808,I303617,I159839,I159856,I159887,I159918,I159949,I159980,I160038,I160055,I241997,I242000,I160072,I242003,I242012,I160089,I160106,I160123,I160140,I242009,I242015,I160157,I160183,I160205,I160222,I160253,I160270,I160301,I242018,I160318,I160335,I242006,I160366,I160383,I160414,I160445,I160476,I160507,I160565,I160582,I160599,I160616,I160633,I160650,I160667,I160684,I160710,I160533,I160732,I160749,I160551,I160780,I160797,I160554,I160828,I160845,I160862,I160536,I160893,I160910,I160557,I160941,I160542,I160972,I160545,I161003,I160539,I161034,I160548,I161092,I161109,I361054,I361051,I161126,I361063,I361066,I161143,I161160,I161177,I161194,I361057,I361048,I161211,I161237,I161259,I161276,I161307,I161324,I161355,I161372,I161389,I361060,I161420,I161437,I161468,I161499,I161530,I161561,I161619,I161636,I161653,I161670,I161687,I161704,I161721,I161738,I161764,I161786,I161803,I161834,I161851,I161882,I161899,I161916,I161947,I161964,I161995,I162026,I162057,I162088,I162146,I162163,I248661,I248664,I162180,I248667,I248676,I162197,I162214,I162231,I162248,I248673,I248679,I162265,I162291,I162114,I162313,I162330,I162132,I162361,I162378,I162135,I162409,I248682,I162426,I162443,I248670,I162117,I162474,I162491,I162138,I162522,I162123,I162553,I162126,I162584,I162120,I162615,I162129,I162673,I162690,I371220,I371217,I162707,I371229,I371232,I162724,I162741,I162758,I162775,I371223,I371214,I162792,I162818,I162840,I162857,I162888,I162905,I162936,I162953,I162970,I371226,I163001,I163018,I163049,I163080,I163111,I163142,I163200,I163217,I369010,I369007,I163234,I369019,I369022,I163251,I163268,I163285,I163302,I369013,I369004,I163319,I163345,I163367,I163384,I163415,I163432,I163463,I163480,I163497,I369016,I163528,I163545,I163576,I163607,I163638,I163669,I163727,I163744,I271985,I271988,I163761,I271991,I272000,I163778,I163795,I163812,I163829,I271997,I272003,I163846,I163872,I163695,I163894,I163911,I163713,I163942,I163959,I163716,I163990,I272006,I164007,I164024,I271994,I163698,I164055,I164072,I163719,I164103,I163704,I164134,I163707,I164165,I163701,I164196,I163710,I164254,I164271,I209629,I209632,I164288,I209635,I209644,I164305,I164322,I164339,I164356,I209641,I209647,I164373,I164399,I164222,I164421,I164438,I164240,I164469,I164486,I164243,I164517,I209650,I164534,I164551,I209638,I164225,I164582,I164599,I164246,I164630,I164231,I164661,I164234,I164692,I164228,I164723,I164237,I164781,I164798,I164815,I164832,I164849,I164866,I164883,I164900,I164926,I164749,I164948,I164965,I164767,I164996,I165013,I164770,I165044,I165061,I165078,I164752,I165109,I165126,I164773,I165157,I164758,I165188,I164761,I165219,I164755,I165250,I164764,I165308,I165325,I165342,I165359,I165376,I165393,I165410,I165427,I165453,I165276,I165475,I165492,I165294,I165523,I165540,I165297,I165571,I165588,I165605,I165279,I165636,I165653,I165300,I165684,I165285,I165715,I165288,I165746,I165282,I165777,I165291,I165835,I165852,I277697,I277700,I165869,I277703,I277712,I165886,I165903,I165920,I165937,I277709,I277715,I165954,I165980,I165803,I166002,I166019,I165821,I166050,I166067,I165824,I166098,I277718,I166115,I166132,I277706,I165806,I166163,I166180,I165827,I166211,I165812,I166242,I165815,I166273,I165809,I166304,I165818,I166362,I166379,I357377,I357365,I166396,I357359,I166413,I166430,I166447,I166464,I357362,I166481,I357368,I166507,I166529,I166546,I166577,I357374,I166594,I166625,I357380,I166642,I166659,I357371,I166690,I166707,I166738,I166769,I166800,I166831,I166889,I166906,I259133,I259136,I166923,I259139,I259148,I166940,I166957,I166974,I166991,I259145,I259151,I167008,I167034,I167056,I167073,I167104,I167121,I167152,I259154,I167169,I167186,I259142,I167217,I167234,I167265,I167296,I167327,I167358,I167416,I167433,I266273,I266276,I167450,I266279,I266288,I167467,I167484,I167501,I167518,I266285,I266291,I167535,I167561,I167583,I167600,I167631,I167648,I167679,I266294,I167696,I167713,I266282,I167744,I167761,I167792,I167823,I167854,I167885,I167943,I167960,I378292,I378289,I167977,I378301,I378304,I167994,I168011,I168028,I168045,I378295,I378286,I168062,I168088,I167911,I168110,I168127,I167929,I168158,I168175,I167932,I168206,I168223,I168240,I378298,I167914,I168271,I168288,I167935,I168319,I167920,I168350,I167923,I168381,I167917,I168412,I167926,I168470,I168487,I168504,I168521,I168538,I168555,I168572,I168589,I168615,I168438,I168637,I168654,I168456,I168685,I168702,I168459,I168733,I168750,I168767,I168441,I168798,I168815,I168462,I168846,I168447,I168877,I168450,I168908,I168444,I168939,I168453,I168997,I169014,I169031,I169048,I169065,I169082,I169099,I169116,I169142,I169164,I169181,I169212,I169229,I169260,I169277,I169294,I169325,I169342,I169373,I169404,I169435,I169466,I169524,I169541,I298356,I298344,I169558,I298347,I298341,I169575,I169592,I169609,I169626,I298338,I169643,I298335,I169669,I169691,I169708,I169739,I169756,I169787,I169804,I169821,I298353,I298350,I169852,I169869,I169900,I169931,I169962,I169993,I170051,I170068,I239141,I239144,I170085,I239147,I239156,I170102,I170119,I170136,I170153,I239153,I239159,I170170,I170196,I170218,I170235,I170266,I170283,I170314,I239162,I170331,I170348,I239150,I170379,I170396,I170427,I170458,I170489,I170520,I170578,I170595,I170612,I170629,I170646,I170663,I170680,I170697,I170723,I170745,I170762,I170793,I170810,I170841,I170858,I170875,I170906,I170923,I170954,I170985,I171016,I171047,I171105,I171122,I241045,I241048,I171139,I241051,I241060,I171156,I171173,I171190,I171207,I241057,I241063,I171224,I171250,I171272,I171289,I171320,I171337,I171368,I241066,I171385,I171402,I241054,I171433,I171450,I171481,I171512,I171543,I171574,I171632,I171649,I365032,I365029,I171666,I365041,I365044,I171683,I171700,I171717,I171734,I365035,I365026,I171751,I171777,I171600,I171799,I171816,I171618,I171847,I171864,I171621,I171895,I171912,I171929,I365038,I171603,I171960,I171977,I171624,I172008,I171609,I172039,I171612,I172070,I171606,I172101,I171615,I172159,I172176,I259609,I259612,I172193,I259615,I259624,I172210,I172227,I172244,I172261,I259621,I259627,I172278,I172304,I172127,I172326,I172343,I172145,I172374,I172391,I172148,I172422,I259630,I172439,I172456,I259618,I172130,I172487,I172504,I172151,I172535,I172136,I172566,I172139,I172597,I172133,I172628,I172142,I172686,I172703,I326811,I326799,I172720,I326793,I172737,I172754,I172771,I172788,I326796,I172805,I326802,I172831,I172654,I172853,I172870,I172672,I172901,I326808,I172918,I172675,I172949,I326814,I172966,I172983,I326805,I172657,I173014,I173031,I172678,I173062,I172663,I173093,I172666,I173124,I172660,I173155,I172669,I173213,I173230,I389784,I389781,I173247,I389793,I389796,I173264,I173281,I173298,I173315,I389787,I389778,I173332,I173358,I173181,I173380,I173397,I173199,I173428,I173445,I173202,I173476,I173493,I173510,I389790,I173184,I173541,I173558,I173205,I173589,I173190,I173620,I173193,I173651,I173187,I173682,I173196,I173740,I173757,I407464,I407461,I173774,I407473,I407476,I173791,I173808,I173825,I173842,I407467,I407458,I173859,I173885,I173708,I173907,I173924,I173726,I173955,I173972,I173729,I174003,I174020,I174037,I407470,I173711,I174068,I174085,I173732,I174116,I173717,I174147,I173720,I174178,I173714,I174209,I173723,I174267,I174284,I338932,I338920,I174301,I338914,I174318,I174335,I174352,I174369,I338917,I174386,I338923,I174412,I174235,I174434,I174451,I174253,I174482,I338929,I174499,I174256,I174530,I338935,I174547,I174564,I338926,I174238,I174595,I174612,I174259,I174643,I174244,I174674,I174247,I174705,I174241,I174736,I174250,I174794,I174811,I174828,I174845,I174862,I174879,I174896,I174913,I174939,I174762,I174961,I174978,I174780,I175009,I175026,I174783,I175057,I175074,I175091,I174765,I175122,I175139,I174786,I175170,I174771,I175201,I174774,I175232,I174768,I175263,I174777,I175321,I175338,I352634,I352622,I175355,I352616,I175372,I175389,I175406,I175423,I352619,I175440,I352625,I175466,I175488,I175505,I175536,I352631,I175553,I175584,I352637,I175601,I175618,I352628,I175649,I175666,I175697,I175728,I175759,I175790,I175848,I175865,I262465,I262468,I175882,I262471,I262480,I175899,I175916,I175933,I175950,I262477,I262483,I175967,I175993,I176015,I176032,I176063,I176080,I176111,I262486,I176128,I176145,I262474,I176176,I176193,I176224,I176255,I176286,I176317,I176375,I176392,I221053,I221056,I176409,I221059,I221068,I176426,I176443,I176460,I176477,I221065,I221071,I176494,I176520,I176343,I176542,I176559,I176361,I176590,I176607,I176364,I176638,I221074,I176655,I176672,I221062,I176346,I176703,I176720,I176367,I176751,I176352,I176782,I176355,I176813,I176349,I176844,I176358,I176902,I176919,I176936,I176953,I176970,I176987,I177004,I177021,I177047,I177069,I177086,I177117,I177134,I177165,I177182,I177199,I177230,I177247,I177278,I177309,I177340,I177371,I177429,I177446,I177463,I177480,I177497,I177514,I177531,I177548,I177574,I177397,I177596,I177613,I177415,I177644,I177661,I177418,I177692,I177709,I177726,I177400,I177757,I177774,I177421,I177805,I177406,I177836,I177409,I177867,I177403,I177898,I177412,I177956,I177973,I177990,I178007,I178024,I178041,I178058,I178075,I178101,I178123,I178140,I178171,I178188,I178219,I178236,I178253,I178284,I178301,I178332,I178363,I178394,I178425,I178483,I178500,I178517,I178534,I178551,I178568,I178585,I178602,I178628,I178650,I178667,I178698,I178715,I178746,I178763,I178780,I178811,I178828,I178859,I178890,I178921,I178952,I179010,I179027,I254373,I254376,I179044,I254379,I254388,I179061,I179078,I179095,I179112,I254385,I254391,I179129,I179155,I179177,I179194,I179225,I179242,I179273,I254394,I179290,I179307,I254382,I179338,I179355,I179386,I179417,I179448,I179479,I179537,I179554,I307839,I307827,I179571,I307821,I179588,I179605,I179622,I179639,I307824,I179656,I307830,I179682,I179704,I179721,I179752,I307836,I179769,I179800,I307842,I179817,I179834,I307833,I179865,I179882,I179913,I179944,I179975,I180006,I180064,I180081,I277221,I277224,I180098,I277227,I277236,I180115,I180132,I180149,I180166,I277233,I277239,I180183,I180209,I180231,I180248,I180279,I180296,I180327,I277242,I180344,I180361,I277230,I180392,I180409,I180440,I180471,I180502,I180533,I180591,I180608,I180625,I180642,I180659,I180676,I180693,I180710,I180736,I180559,I180758,I180775,I180577,I180806,I180823,I180580,I180854,I180871,I180888,I180562,I180919,I180936,I180583,I180967,I180568,I180998,I180571,I181029,I180565,I181060,I180574,I181118,I181135,I377850,I377847,I181152,I377859,I377862,I181169,I181186,I181203,I181220,I377853,I377844,I181237,I181263,I181086,I181285,I181302,I181104,I181333,I181350,I181107,I181381,I181398,I181415,I377856,I181089,I181446,I181463,I181110,I181494,I181095,I181525,I181098,I181556,I181092,I181587,I181101,I181645,I181662,I287289,I287277,I181679,I287280,I287274,I181696,I181713,I181730,I181747,I287271,I181764,I287268,I181790,I181613,I181812,I181829,I181631,I181860,I181877,I181634,I181908,I181925,I181942,I287286,I287283,I181616,I181973,I181990,I181637,I182021,I181622,I182052,I181625,I182083,I181619,I182114,I181628,I182172,I182189,I346310,I346298,I182206,I346292,I182223,I182240,I182257,I182274,I346295,I182291,I346301,I182317,I182339,I182356,I182387,I346307,I182404,I182435,I346313,I182452,I182469,I346304,I182500,I182517,I182548,I182579,I182610,I182641,I182699,I182716,I300464,I300452,I182733,I300455,I300449,I182750,I182767,I182784,I182801,I300446,I182818,I300443,I182844,I182667,I182866,I182883,I182685,I182914,I182931,I182688,I182962,I182979,I182996,I300461,I300458,I182670,I183027,I183044,I182691,I183075,I182676,I183106,I182679,I183137,I182673,I183168,I182682,I183226,I183243,I183260,I183277,I183294,I183311,I183328,I183345,I183371,I183393,I183410,I183441,I183458,I183489,I183506,I183523,I183554,I183571,I183602,I183633,I183664,I183695,I183753,I183770,I183787,I183804,I183821,I183838,I183855,I183872,I183898,I183721,I183920,I183937,I183739,I183968,I183985,I183742,I184016,I184033,I184050,I183724,I184081,I184098,I183745,I184129,I183730,I184160,I183733,I184191,I183727,I184222,I183736,I184280,I184297,I273413,I273416,I184314,I273419,I273428,I184331,I184348,I184365,I184382,I273425,I273431,I184399,I184425,I184447,I184464,I184495,I184512,I184543,I273434,I184560,I184577,I273422,I184608,I184625,I184656,I184687,I184718,I184749,I184807,I184824,I339459,I339447,I184841,I339441,I184858,I184875,I184892,I184909,I339444,I184926,I339450,I184952,I184775,I184974,I184991,I184793,I185022,I339456,I185039,I184796,I185070,I339462,I185087,I185104,I339453,I184778,I185135,I185152,I184799,I185183,I184784,I185214,I184787,I185245,I184781,I185276,I184790,I185334,I185351,I305204,I305192,I185368,I305186,I185385,I185402,I185419,I185436,I305189,I185453,I305195,I185479,I185501,I185518,I185549,I305201,I185566,I185597,I305207,I185614,I185631,I305198,I185662,I185679,I185710,I185741,I185772,I185803,I185861,I185878,I352107,I352095,I185895,I352089,I185912,I185929,I185946,I185963,I352092,I185980,I352098,I186006,I186028,I186045,I186076,I352104,I186093,I186124,I352110,I186141,I186158,I352101,I186189,I186206,I186237,I186268,I186299,I186330,I186388,I186405,I186422,I186439,I186456,I186473,I186490,I186507,I186533,I186555,I186572,I186603,I186620,I186651,I186668,I186685,I186716,I186733,I186764,I186795,I186826,I186857,I186915,I186932,I357904,I357892,I186949,I357886,I186966,I186983,I187000,I187017,I357889,I187034,I357895,I187060,I186883,I187082,I187099,I186901,I187130,I357901,I187147,I186904,I187178,I357907,I187195,I187212,I357898,I186886,I187243,I187260,I186907,I187291,I186892,I187322,I186895,I187353,I186889,I187384,I186898,I187442,I187459,I187476,I187493,I187510,I187527,I187544,I187561,I187587,I187410,I187609,I187626,I187428,I187657,I187674,I187431,I187705,I187722,I187739,I187413,I187770,I187787,I187434,I187818,I187419,I187849,I187422,I187880,I187416,I187911,I187425,I187969,I187986,I188003,I188020,I188037,I188054,I188071,I188088,I188114,I187937,I188136,I188153,I187955,I188184,I188201,I187958,I188232,I188249,I188266,I187940,I188297,I188314,I187961,I188345,I187946,I188376,I187949,I188407,I187943,I188438,I187952,I188496,I188513,I188530,I188547,I188564,I188581,I188598,I188615,I188641,I188464,I188663,I188680,I188482,I188711,I188728,I188485,I188759,I188776,I188793,I188467,I188824,I188841,I188488,I188872,I188473,I188903,I188476,I188934,I188470,I188965,I188479,I189023,I189040,I189057,I189074,I189091,I189108,I189125,I189142,I189168,I189190,I189207,I189238,I189255,I189286,I189303,I189320,I189351,I189368,I189399,I189430,I189461,I189492,I189550,I189567,I318379,I318367,I189584,I318361,I189601,I189618,I189635,I189652,I318364,I189669,I318370,I189695,I189518,I189717,I189734,I189536,I189765,I318376,I189782,I189539,I189813,I318382,I189830,I189847,I318373,I189521,I189878,I189895,I189542,I189926,I189527,I189957,I189530,I189988,I189524,I190019,I189533,I190077,I190094,I400834,I400831,I190111,I400843,I400846,I190128,I190145,I190162,I190179,I400837,I400828,I190196,I190222,I190045,I190244,I190261,I190063,I190292,I190309,I190066,I190340,I190357,I190374,I400840,I190048,I190405,I190422,I190069,I190453,I190054,I190484,I190057,I190515,I190051,I190546,I190060,I190604,I190621,I190638,I190655,I190672,I190689,I190706,I190723,I190749,I190572,I190771,I190788,I190590,I190819,I190836,I190593,I190867,I190884,I190901,I190575,I190932,I190949,I190596,I190980,I190581,I191011,I190584,I191042,I190578,I191073,I190587,I191131,I191148,I263893,I263896,I191165,I263899,I263908,I191182,I191199,I191216,I191233,I263905,I263911,I191250,I191276,I191298,I191315,I191346,I191363,I191394,I263914,I191411,I191428,I263902,I191459,I191476,I191507,I191538,I191569,I191600,I191658,I191675,I204393,I204396,I191692,I204399,I204408,I191709,I191726,I191743,I191760,I204405,I204411,I191777,I191803,I191626,I191825,I191842,I191644,I191873,I191890,I191647,I191921,I204414,I191938,I191955,I204402,I191629,I191986,I192003,I191650,I192034,I191635,I192065,I191638,I192096,I191632,I192127,I191641,I192185,I192202,I316271,I316259,I192219,I316253,I192236,I192253,I192270,I192287,I316256,I192304,I316262,I192330,I192352,I192369,I192400,I316268,I192417,I192448,I316274,I192465,I192482,I316265,I192513,I192530,I192561,I192592,I192623,I192654,I192712,I192729,I192746,I192763,I192780,I192797,I192814,I192831,I192857,I192879,I192896,I192927,I192944,I192975,I192992,I193009,I193040,I193057,I193088,I193119,I193150,I193181,I193239,I193256,I203917,I203920,I193273,I203923,I203932,I193290,I193307,I193324,I193341,I203929,I203935,I193358,I193384,I193406,I193423,I193454,I193471,I193502,I203938,I193519,I193536,I203926,I193567,I193584,I193615,I193646,I193677,I193708,I193766,I193783,I275317,I275320,I193800,I275323,I275332,I193817,I193834,I193851,I193868,I275329,I275335,I193885,I193911,I193734,I193933,I193950,I193752,I193981,I193998,I193755,I194029,I275338,I194046,I194063,I275326,I193737,I194094,I194111,I193758,I194142,I193743,I194173,I193746,I194204,I193740,I194235,I193749,I194293,I194310,I232001,I232004,I194327,I232007,I232016,I194344,I194361,I194378,I194395,I232013,I232019,I194412,I194438,I194261,I194460,I194477,I194279,I194508,I194525,I194282,I194556,I232022,I194573,I194590,I232010,I194264,I194621,I194638,I194285,I194669,I194270,I194700,I194273,I194731,I194267,I194762,I194276,I194820,I194837,I194854,I194871,I194888,I194905,I194922,I194939,I194965,I194788,I194987,I195004,I194806,I195035,I195052,I194809,I195083,I195100,I195117,I194791,I195148,I195165,I194812,I195196,I194797,I195227,I194800,I195258,I194794,I195289,I194803,I195347,I195364,I195381,I195398,I195415,I195432,I195449,I195466,I195492,I195514,I195531,I195562,I195579,I195610,I195627,I195644,I195675,I195692,I195723,I195754,I195785,I195816,I195874,I195891,I401718,I401715,I195908,I401727,I401730,I195925,I195942,I195959,I195976,I401721,I401712,I195993,I196019,I196041,I196058,I196089,I196106,I196137,I196154,I196171,I401724,I196202,I196219,I196250,I196281,I196312,I196343,I196401,I196418,I348418,I348406,I196435,I348400,I196452,I196469,I196486,I196503,I348403,I196520,I348409,I196546,I196568,I196585,I196616,I348415,I196633,I196664,I348421,I196681,I196698,I348412,I196729,I196746,I196777,I196808,I196839,I196870,I196928,I196945,I196962,I196979,I196996,I197013,I197030,I197047,I197073,I196896,I197095,I197112,I196914,I197143,I197160,I196917,I197191,I197208,I197225,I196899,I197256,I197273,I196920,I197304,I196905,I197335,I196908,I197366,I196902,I197397,I196911,I197455,I197472,I286265,I286268,I197489,I286271,I286280,I197506,I197523,I197540,I197557,I286277,I286283,I197574,I197600,I197423,I197622,I197639,I197441,I197670,I197687,I197444,I197718,I286286,I197735,I197752,I286274,I197426,I197783,I197800,I197447,I197831,I197432,I197862,I197435,I197893,I197429,I197924,I197438,I197982,I197999,I354215,I354203,I198016,I354197,I198033,I198050,I198067,I198084,I354200,I198101,I354206,I198127,I197950,I198149,I198166,I197968,I198197,I354212,I198214,I197971,I198245,I354218,I198262,I198279,I354209,I197953,I198310,I198327,I197974,I198358,I197959,I198389,I197962,I198420,I197956,I198451,I197965,I198509,I198526,I329973,I329961,I198543,I329955,I198560,I198577,I198594,I198611,I329958,I198628,I329964,I198654,I198477,I198676,I198693,I198495,I198724,I329970,I198741,I198498,I198772,I329976,I198789,I198806,I329967,I198480,I198837,I198854,I198501,I198885,I198486,I198916,I198489,I198947,I198483,I198978,I198492,I199036,I199053,I364590,I364587,I199070,I364599,I364602,I199087,I199104,I199121,I199138,I364593,I364584,I199155,I199181,I199004,I199203,I199220,I199022,I199251,I199268,I199025,I199299,I199316,I199333,I364596,I199007,I199364,I199381,I199028,I199412,I199013,I199443,I199016,I199474,I199010,I199505,I199019,I199563,I199580,I396856,I396853,I199597,I396865,I396868,I199614,I199631,I199648,I199665,I396859,I396850,I199682,I199708,I199730,I199747,I199778,I199795,I199826,I199843,I199860,I396862,I199891,I199908,I199939,I199970,I200001,I200032,I200090,I200107,I364148,I364145,I200124,I364157,I364160,I200141,I200158,I200175,I200192,I364151,I364142,I200209,I200235,I200058,I200257,I200274,I200076,I200305,I200322,I200079,I200353,I200370,I200387,I364154,I200061,I200418,I200435,I200082,I200466,I200067,I200497,I200070,I200528,I200064,I200559,I200073,I200614,I200631,I200648,I200665,I200682,I200699,I200716,I200733,I200750,I200767,I200784,I200801,I200818,I200835,I200880,I200911,I200942,I200959,I200990,I201035,I201090,I201107,I201124,I201141,I201158,I201175,I201192,I201209,I201226,I201243,I201260,I201277,I201294,I201311,I201356,I201387,I201418,I201435,I201466,I201511,I201566,I201583,I201600,I201617,I201634,I201651,I201668,I201685,I201702,I201719,I201736,I201753,I201770,I201787,I201832,I201863,I201894,I201911,I201942,I201987,I202042,I202059,I202076,I202093,I202110,I202127,I202144,I202161,I202178,I202195,I202212,I202229,I202246,I202263,I202034,I202019,I202308,I202013,I202339,I202016,I202370,I202387,I202022,I202418,I202031,I202028,I202463,I202025,I202518,I202535,I202552,I202569,I202586,I202603,I202620,I202637,I202654,I202671,I202688,I202705,I202722,I202739,I202784,I202815,I202846,I202863,I202894,I202939,I202994,I203011,I203028,I203045,I203062,I203079,I203096,I203113,I203130,I203147,I203164,I203181,I203198,I203215,I203260,I203291,I203322,I203339,I203370,I203415,I203470,I203487,I203504,I203521,I203538,I203555,I203572,I203589,I203606,I203623,I203640,I203657,I203674,I203691,I203736,I203767,I203798,I203815,I203846,I203891,I203946,I203963,I399063,I399066,I203980,I203997,I399060,I399078,I204014,I204031,I399069,I204048,I204065,I204082,I204099,I204116,I399075,I399072,I204133,I204150,I204167,I204212,I204243,I204274,I204291,I204322,I204367,I204422,I204439,I204456,I204473,I204490,I204507,I204524,I204541,I204558,I204575,I204592,I204609,I204626,I204643,I204688,I204719,I204750,I204767,I204798,I204843,I204898,I204915,I204932,I204949,I204966,I204983,I205000,I205017,I205034,I205051,I205068,I205085,I205102,I205119,I205164,I205195,I205226,I205243,I205274,I205319,I205374,I205391,I384477,I384480,I205408,I205425,I384474,I384492,I205442,I205459,I384483,I205476,I205493,I205510,I205527,I205544,I384489,I384486,I205561,I205578,I205595,I205640,I205671,I205702,I205719,I205750,I205795,I205850,I205867,I205884,I205901,I205918,I205935,I205952,I205969,I205986,I206003,I206020,I206037,I206054,I206071,I206116,I206147,I206178,I206195,I206226,I206271,I206326,I206343,I206360,I206377,I206394,I206411,I206428,I206445,I206462,I206479,I206496,I206513,I206530,I206547,I206318,I206303,I206592,I206297,I206623,I206300,I206654,I206671,I206306,I206702,I206315,I206312,I206747,I206309,I206802,I206819,I206836,I206853,I206870,I206887,I206904,I206921,I206938,I206955,I206972,I206989,I207006,I207023,I207068,I207099,I207130,I207147,I207178,I207223,I207278,I207295,I403483,I403486,I207312,I207329,I403480,I403498,I207346,I207363,I403489,I207380,I207397,I207414,I207431,I207448,I403495,I403492,I207465,I207482,I207499,I207270,I207255,I207544,I207249,I207575,I207252,I207606,I207623,I207258,I207654,I207267,I207264,I207699,I207261,I207754,I207771,I345765,I345786,I207788,I345771,I207805,I345783,I207822,I345774,I207839,I345768,I207856,I207873,I207890,I207907,I207924,I345777,I345780,I207941,I207958,I207975,I207746,I207731,I208020,I207725,I208051,I207728,I208082,I208099,I207734,I208130,I207743,I207740,I208175,I207737,I208230,I208247,I338387,I338408,I208264,I338393,I208281,I338405,I208298,I338396,I208315,I338390,I208332,I208349,I208366,I208383,I208400,I338399,I338402,I208417,I208434,I208451,I208496,I208527,I208558,I208575,I208606,I208651,I208706,I208723,I208740,I208757,I208774,I208791,I208808,I208825,I208842,I208859,I208876,I208893,I208910,I208927,I208972,I209003,I209034,I209051,I209082,I209127,I209182,I209199,I209216,I209233,I209250,I209267,I209284,I209301,I209318,I209335,I209352,I209369,I209386,I209403,I209448,I209479,I209510,I209527,I209558,I209603,I209658,I209675,I209692,I209709,I209726,I209743,I209760,I209777,I209794,I209811,I209828,I209845,I209862,I209879,I209924,I209955,I209986,I210003,I210034,I210079,I210134,I210151,I347873,I347894,I210168,I347879,I210185,I347891,I210202,I347882,I210219,I347876,I210236,I210253,I210270,I210287,I210304,I347885,I347888,I210321,I210338,I210355,I210126,I210111,I210400,I210105,I210431,I210108,I210462,I210479,I210114,I210510,I210123,I210120,I210555,I210117,I210610,I210627,I289906,I289903,I210644,I289912,I210661,I289924,I289909,I210678,I210695,I289915,I210712,I210729,I210746,I210763,I210780,I289921,I210797,I289918,I210814,I210831,I210876,I210907,I210938,I210955,I210986,I211031,I211086,I211103,I211120,I211137,I211154,I211171,I211188,I211205,I211222,I211239,I211256,I211273,I211290,I211307,I211078,I211063,I211352,I211057,I211383,I211060,I211414,I211431,I211066,I211462,I211075,I211072,I211507,I211069,I211562,I211579,I211596,I211613,I211630,I211647,I211664,I211681,I211698,I211715,I211732,I211749,I211766,I211783,I211554,I211539,I211828,I211533,I211859,I211536,I211890,I211907,I211542,I211938,I211551,I211548,I211983,I211545,I212038,I212055,I212072,I212089,I212106,I212123,I212140,I212157,I212174,I212191,I212208,I212225,I212242,I212259,I212304,I212335,I212366,I212383,I212414,I212459,I212514,I212531,I319415,I319436,I212548,I319421,I212565,I319433,I212582,I319424,I212599,I319418,I212616,I212633,I212650,I212667,I212684,I319427,I319430,I212701,I212718,I212735,I212506,I212491,I212780,I212485,I212811,I212488,I212842,I212859,I212494,I212890,I212503,I212500,I212935,I212497,I212990,I213007,I390665,I390668,I213024,I213041,I390662,I390680,I213058,I213075,I390671,I213092,I213109,I213126,I213143,I213160,I390677,I390674,I213177,I213194,I213211,I213256,I213287,I213318,I213335,I213366,I213411,I213466,I213483,I213500,I213517,I213534,I213551,I213568,I213585,I213602,I213619,I213636,I213653,I213670,I213687,I213732,I213763,I213794,I213811,I213842,I213887,I213942,I213959,I213976,I213993,I214010,I214027,I214044,I214061,I214078,I214095,I214112,I214129,I214146,I214163,I213934,I213919,I214208,I213913,I214239,I213916,I214270,I214287,I213922,I214318,I213931,I213928,I214363,I213925,I214418,I214435,I214452,I214469,I214486,I214503,I214520,I214537,I214554,I214571,I214588,I214605,I214622,I214639,I214684,I214715,I214746,I214763,I214794,I214839,I214894,I214911,I321523,I321544,I214928,I321529,I214945,I321541,I214962,I321532,I214979,I321526,I214996,I215013,I215030,I215047,I215064,I321535,I321538,I215081,I215098,I215115,I215160,I215191,I215222,I215239,I215270,I215315,I215370,I215387,I215404,I215421,I215438,I215455,I215472,I215489,I215506,I215523,I215540,I215557,I215574,I215591,I215636,I215667,I215698,I215715,I215746,I215791,I215846,I215863,I358413,I358434,I215880,I358419,I215897,I358431,I215914,I358422,I215931,I358416,I215948,I215965,I215982,I215999,I216016,I358425,I358428,I216033,I216050,I216067,I216112,I216143,I216174,I216191,I216222,I216267,I216322,I216339,I216356,I216373,I216390,I216407,I216424,I216441,I216458,I216475,I216492,I216509,I216526,I216543,I216588,I216619,I216650,I216667,I216698,I216743,I216798,I216815,I369891,I369894,I216832,I216849,I369888,I369906,I216866,I216883,I369897,I216900,I216917,I216934,I216951,I216968,I369903,I369900,I216985,I217002,I217019,I216790,I216775,I217064,I216769,I217095,I216772,I217126,I217143,I216778,I217174,I216787,I216784,I217219,I216781,I217274,I217291,I217308,I217325,I217342,I217359,I217376,I217393,I217410,I217427,I217444,I217461,I217478,I217495,I217540,I217571,I217602,I217619,I217650,I217695,I217750,I217767,I217784,I217801,I217818,I217835,I217852,I217869,I217886,I217903,I217920,I217937,I217954,I217971,I217742,I217727,I218016,I217721,I218047,I217724,I218078,I218095,I217730,I218126,I217739,I217736,I218171,I217733,I218226,I218243,I218260,I218277,I218294,I218311,I218328,I218345,I218362,I218379,I218396,I218413,I218430,I218447,I218492,I218523,I218554,I218571,I218602,I218647,I218702,I218719,I394201,I394204,I218736,I218753,I394198,I394216,I218770,I218787,I394207,I218804,I218821,I218838,I218855,I218872,I394213,I394210,I218889,I218906,I218923,I218694,I218679,I218968,I218673,I218999,I218676,I219030,I219047,I218682,I219078,I218691,I218688,I219123,I218685,I219178,I219195,I219212,I219229,I219246,I219263,I219280,I219297,I219314,I219331,I219348,I219365,I219382,I219399,I219170,I219155,I219444,I219149,I219475,I219152,I219506,I219523,I219158,I219554,I219167,I219164,I219599,I219161,I219654,I219671,I219688,I219705,I219722,I219739,I219756,I219773,I219790,I219807,I219824,I219841,I219858,I219875,I219920,I219951,I219982,I219999,I220030,I220075,I220130,I220147,I301500,I301497,I220164,I301506,I220181,I301518,I301503,I220198,I220215,I301509,I220232,I220249,I220266,I220283,I220300,I301515,I220317,I301512,I220334,I220351,I220122,I220107,I220396,I220101,I220427,I220104,I220458,I220475,I220110,I220506,I220119,I220116,I220551,I220113,I220606,I220623,I408787,I408790,I220640,I220657,I408784,I408802,I220674,I220691,I408793,I220708,I220725,I220742,I220759,I220776,I408799,I408796,I220793,I220810,I220827,I220598,I220583,I220872,I220577,I220903,I220580,I220934,I220951,I220586,I220982,I220595,I220592,I221027,I220589,I221082,I221099,I290960,I290957,I221116,I290966,I221133,I290978,I290963,I221150,I221167,I290969,I221184,I221201,I221218,I221235,I221252,I290975,I221269,I290972,I221286,I221303,I221348,I221379,I221410,I221427,I221458,I221503,I221558,I221575,I221592,I221609,I221626,I221643,I221660,I221677,I221694,I221711,I221728,I221745,I221762,I221779,I221824,I221855,I221886,I221903,I221934,I221979,I222034,I222051,I222068,I222085,I222102,I222119,I222136,I222153,I222170,I222187,I222204,I222221,I222238,I222255,I222026,I222011,I222300,I222005,I222331,I222008,I222362,I222379,I222014,I222410,I222023,I222020,I222455,I222017,I222510,I222527,I327320,I327341,I222544,I327326,I222561,I327338,I222578,I327329,I222595,I327323,I222612,I222629,I222646,I222663,I222680,I327332,I327335,I222697,I222714,I222731,I222502,I222487,I222776,I222481,I222807,I222484,I222838,I222855,I222490,I222886,I222499,I222496,I222931,I222493,I222986,I223003,I223020,I223037,I223054,I223071,I223088,I223105,I223122,I223139,I223156,I223173,I223190,I223207,I223252,I223283,I223314,I223331,I223362,I223407,I223462,I223479,I223496,I223513,I223530,I223547,I223564,I223581,I223598,I223615,I223632,I223649,I223666,I223683,I223454,I223439,I223728,I223433,I223759,I223436,I223790,I223807,I223442,I223838,I223451,I223448,I223883,I223445,I223938,I223955,I325212,I325233,I223972,I325218,I223989,I325230,I224006,I325221,I224023,I325215,I224040,I224057,I224074,I224091,I224108,I325224,I325227,I224125,I224142,I224159,I224204,I224235,I224266,I224283,I224314,I224359,I224414,I224431,I404809,I404812,I224448,I224465,I404806,I404824,I224482,I224499,I404815,I224516,I224533,I224550,I224567,I224584,I404821,I404818,I224601,I224618,I224635,I224406,I224391,I224680,I224385,I224711,I224388,I224742,I224759,I224394,I224790,I224403,I224400,I224835,I224397,I224890,I224907,I336279,I336300,I224924,I336285,I224941,I336297,I224958,I336288,I224975,I336282,I224992,I225009,I225026,I225043,I225060,I336291,I336294,I225077,I225094,I225111,I225156,I225187,I225218,I225235,I225266,I225311,I225366,I225383,I380057,I380060,I225400,I225417,I380054,I380072,I225434,I225451,I380063,I225468,I225485,I225502,I225519,I225536,I380069,I380066,I225553,I225570,I225587,I225632,I225663,I225694,I225711,I225742,I225787,I225842,I225859,I225876,I225893,I225910,I225927,I225944,I225961,I225978,I225995,I226012,I226029,I226046,I226063,I226108,I226139,I226170,I226187,I226218,I226263,I226318,I226335,I226352,I226369,I226386,I226403,I226420,I226437,I226454,I226471,I226488,I226505,I226522,I226539,I226310,I226295,I226584,I226289,I226615,I226292,I226646,I226663,I226298,I226694,I226307,I226304,I226739,I226301,I226794,I226811,I398179,I398182,I226828,I226845,I398176,I398194,I226862,I226879,I398185,I226896,I226913,I226930,I226947,I226964,I398191,I398188,I226981,I226998,I227015,I226786,I226771,I227060,I226765,I227091,I226768,I227122,I227139,I226774,I227170,I226783,I226780,I227215,I226777,I227270,I227287,I334171,I334192,I227304,I334177,I227321,I334189,I227338,I334180,I227355,I334174,I227372,I227389,I227406,I227423,I227440,I334183,I334186,I227457,I227474,I227491,I227536,I227567,I227598,I227615,I227646,I227691,I227746,I227763,I227780,I227797,I227814,I227831,I227848,I227865,I227882,I227899,I227916,I227933,I227950,I227967,I228012,I228043,I228074,I228091,I228122,I228167,I228222,I228239,I351035,I351056,I228256,I351041,I228273,I351053,I228290,I351044,I228307,I351038,I228324,I228341,I228358,I228375,I228392,I351047,I351050,I228409,I228426,I228443,I228214,I228199,I228488,I228193,I228519,I228196,I228550,I228567,I228202,I228598,I228211,I228208,I228643,I228205,I228698,I228715,I228732,I228749,I228766,I228783,I228800,I228817,I228834,I228851,I228868,I228885,I228902,I228919,I228964,I228995,I229026,I229043,I229074,I229119,I229174,I229191,I359467,I359488,I229208,I359473,I229225,I359485,I229242,I359476,I229259,I359470,I229276,I229293,I229310,I229327,I229344,I359479,I359482,I229361,I229378,I229395,I229440,I229471,I229502,I229519,I229550,I229595,I229650,I229667,I229684,I229701,I229718,I229735,I229752,I229769,I229786,I229803,I229820,I229837,I229854,I229871,I229642,I229627,I229916,I229621,I229947,I229624,I229978,I229995,I229630,I230026,I229639,I229636,I230071,I229633,I230126,I230143,I230160,I230177,I230194,I230211,I230228,I230245,I230262,I230279,I230296,I230313,I230330,I230347,I230392,I230423,I230454,I230471,I230502,I230547,I230602,I230619,I372985,I372988,I230636,I230653,I372982,I373000,I230670,I230687,I372991,I230704,I230721,I230738,I230755,I230772,I372997,I372994,I230789,I230806,I230823,I230868,I230899,I230930,I230947,I230978,I231023,I231078,I231095,I231112,I231129,I231146,I231163,I231180,I231197,I231214,I231231,I231248,I231265,I231282,I231299,I231344,I231375,I231406,I231423,I231454,I231499,I231554,I231571,I231588,I231605,I231622,I231639,I231656,I231673,I231690,I231707,I231724,I231741,I231758,I231775,I231820,I231851,I231882,I231899,I231930,I231975,I232030,I232047,I324158,I324179,I232064,I324164,I232081,I324176,I232098,I324167,I232115,I324161,I232132,I232149,I232166,I232183,I232200,I324170,I324173,I232217,I232234,I232251,I232296,I232327,I232358,I232375,I232406,I232451,I232506,I232523,I232540,I232557,I232574,I232591,I232608,I232625,I232642,I232659,I232676,I232693,I232710,I232727,I232772,I232803,I232834,I232851,I232882,I232927,I232982,I232999,I233016,I233033,I233050,I233067,I233084,I233101,I233118,I233135,I233152,I233169,I233186,I233203,I232974,I232959,I233248,I232953,I233279,I232956,I233310,I233327,I232962,I233358,I232971,I232968,I233403,I232965,I233458,I233475,I233492,I233509,I233526,I233543,I233560,I233577,I233594,I233611,I233628,I233645,I233662,I233679,I233724,I233755,I233786,I233803,I233834,I233879,I233934,I233951,I233968,I233985,I234002,I234019,I234036,I234053,I234070,I234087,I234104,I234121,I234138,I234155,I234200,I234231,I234262,I234279,I234310,I234355,I234410,I234427,I234444,I234461,I234478,I234495,I234512,I234529,I234546,I234563,I234580,I234597,I234614,I234631,I234402,I234387,I234676,I234381,I234707,I234384,I234738,I234755,I234390,I234786,I234399,I234396,I234831,I234393,I234886,I234903,I409229,I409232,I234920,I234937,I409226,I409244,I234954,I234971,I409235,I234988,I235005,I235022,I235039,I235056,I409241,I409238,I235073,I235090,I235107,I235152,I235183,I235214,I235231,I235262,I235307,I235362,I235379,I235396,I235413,I235430,I235447,I235464,I235481,I235498,I235515,I235532,I235549,I235566,I235583,I235628,I235659,I235690,I235707,I235738,I235783,I235838,I235855,I235872,I235889,I235906,I235923,I235940,I235957,I235974,I235991,I236008,I236025,I236042,I236059,I235830,I235815,I236104,I235809,I236135,I235812,I236166,I236183,I235818,I236214,I235827,I235824,I236259,I235821,I236314,I236331,I236348,I236365,I236382,I236399,I236416,I236433,I236450,I236467,I236484,I236501,I236518,I236535,I236306,I236291,I236580,I236285,I236611,I236288,I236642,I236659,I236294,I236690,I236303,I236300,I236735,I236297,I236790,I236807,I236824,I236841,I236858,I236875,I236892,I236909,I236926,I236943,I236960,I236977,I236994,I237011,I236782,I236767,I237056,I236761,I237087,I236764,I237118,I237135,I236770,I237166,I236779,I236776,I237211,I236773,I237266,I237283,I237300,I237317,I237334,I237351,I237368,I237385,I237402,I237419,I237436,I237453,I237470,I237487,I237258,I237243,I237532,I237237,I237563,I237240,I237594,I237611,I237246,I237642,I237255,I237252,I237687,I237249,I237742,I237759,I237776,I237793,I237810,I237827,I237844,I237861,I237878,I237895,I237912,I237929,I237946,I237963,I237734,I237719,I238008,I237713,I238039,I237716,I238070,I238087,I237722,I238118,I237731,I237728,I238163,I237725,I238218,I238235,I238252,I238269,I238286,I238303,I238320,I238337,I238354,I238371,I238388,I238405,I238422,I238439,I238484,I238515,I238546,I238563,I238594,I238639,I238694,I238711,I238728,I238745,I238762,I238779,I238796,I238813,I238830,I238847,I238864,I238881,I238898,I238915,I238960,I238991,I239022,I239039,I239070,I239115,I239170,I239187,I239204,I239221,I239238,I239255,I239272,I239289,I239306,I239323,I239340,I239357,I239374,I239391,I239436,I239467,I239498,I239515,I239546,I239591,I239646,I239663,I239680,I239697,I239714,I239731,I239748,I239765,I239782,I239799,I239816,I239833,I239850,I239867,I239638,I239623,I239912,I239617,I239943,I239620,I239974,I239991,I239626,I240022,I239635,I239632,I240067,I239629,I240122,I240139,I240156,I240173,I240190,I240207,I240224,I240241,I240258,I240275,I240292,I240309,I240326,I240343,I240388,I240419,I240450,I240467,I240498,I240543,I240598,I240615,I386245,I386248,I240632,I240649,I386242,I386260,I240666,I240683,I386251,I240700,I240717,I240734,I240751,I240768,I386257,I386254,I240785,I240802,I240819,I240590,I240575,I240864,I240569,I240895,I240572,I240926,I240943,I240578,I240974,I240587,I240584,I241019,I240581,I241074,I241091,I381825,I381828,I241108,I241125,I381822,I381840,I241142,I241159,I381831,I241176,I241193,I241210,I241227,I241244,I381837,I381834,I241261,I241278,I241295,I241340,I241371,I241402,I241419,I241450,I241495,I241550,I241567,I391549,I391552,I241584,I241601,I391546,I391564,I241618,I241635,I391555,I241652,I241669,I241686,I241703,I241720,I391561,I391558,I241737,I241754,I241771,I241816,I241847,I241878,I241895,I241926,I241971,I242026,I242043,I242060,I242077,I242094,I242111,I242128,I242145,I242162,I242179,I242196,I242213,I242230,I242247,I242292,I242323,I242354,I242371,I242402,I242447,I242502,I242519,I242536,I242553,I242570,I242587,I242604,I242621,I242638,I242655,I242672,I242689,I242706,I242723,I242494,I242479,I242768,I242473,I242799,I242476,I242830,I242847,I242482,I242878,I242491,I242488,I242923,I242485,I242978,I242995,I292014,I292011,I243012,I292020,I243029,I292032,I292017,I243046,I243063,I292023,I243080,I243097,I243114,I243131,I243148,I292029,I243165,I292026,I243182,I243199,I242970,I242955,I243244,I242949,I243275,I242952,I243306,I243323,I242958,I243354,I242967,I242964,I243399,I242961,I243454,I243471,I243488,I243505,I243522,I243539,I243556,I243573,I243590,I243607,I243624,I243641,I243658,I243675,I243720,I243751,I243782,I243799,I243830,I243875,I243930,I243947,I335225,I335246,I243964,I335231,I243981,I335243,I243998,I335234,I244015,I335228,I244032,I244049,I244066,I244083,I244100,I335237,I335240,I244117,I244134,I244151,I243922,I243907,I244196,I243901,I244227,I243904,I244258,I244275,I243910,I244306,I243919,I243916,I244351,I243913,I244406,I244423,I244440,I244457,I244474,I244491,I244508,I244525,I244542,I244559,I244576,I244593,I244610,I244627,I244672,I244703,I244734,I244751,I244782,I244827,I244882,I244899,I244916,I244933,I244950,I244967,I244984,I245001,I245018,I245035,I245052,I245069,I245086,I245103,I245148,I245179,I245210,I245227,I245258,I245303,I245358,I245375,I245392,I245409,I245426,I245443,I245460,I245477,I245494,I245511,I245528,I245545,I245562,I245579,I245624,I245655,I245686,I245703,I245734,I245779,I245834,I245851,I245868,I245885,I245902,I245919,I245936,I245953,I245970,I245987,I246004,I246021,I246038,I246055,I245826,I245811,I246100,I245805,I246131,I245808,I246162,I246179,I245814,I246210,I245823,I245820,I246255,I245817,I246310,I246327,I246344,I246361,I246378,I246395,I246412,I246429,I246446,I246463,I246480,I246497,I246514,I246531,I246576,I246607,I246638,I246655,I246686,I246731,I246786,I246803,I246820,I246837,I246854,I246871,I246888,I246905,I246922,I246939,I246956,I246973,I246990,I247007,I247052,I247083,I247114,I247131,I247162,I247207,I247262,I247279,I247296,I247313,I247330,I247347,I247364,I247381,I247398,I247415,I247432,I247449,I247466,I247483,I247254,I247239,I247528,I247233,I247559,I247236,I247590,I247607,I247242,I247638,I247251,I247248,I247683,I247245,I247738,I247755,I247772,I247789,I247806,I247823,I247840,I247857,I247874,I247891,I247908,I247925,I247942,I247959,I248004,I248035,I248066,I248083,I248114,I248159,I248214,I248231,I359994,I360015,I248248,I360000,I248265,I360012,I248282,I360003,I248299,I359997,I248316,I248333,I248350,I248367,I248384,I360006,I360009,I248401,I248418,I248435,I248480,I248511,I248542,I248559,I248590,I248635,I248690,I248707,I410113,I410116,I248724,I248741,I410110,I410128,I248758,I248775,I410119,I248792,I248809,I248826,I248843,I248860,I410125,I410122,I248877,I248894,I248911,I248956,I248987,I249018,I249035,I249066,I249111,I249166,I249183,I297811,I297808,I249200,I297817,I249217,I297829,I297814,I249234,I249251,I297820,I249268,I249285,I249302,I249319,I249336,I297826,I249353,I297823,I249370,I249387,I249432,I249463,I249494,I249511,I249542,I249587,I249642,I249659,I249676,I249693,I249710,I249727,I249744,I249761,I249778,I249795,I249812,I249829,I249846,I249863,I249908,I249939,I249970,I249987,I250018,I250063,I250118,I250135,I370775,I370778,I250152,I250169,I370772,I370790,I250186,I250203,I370781,I250220,I250237,I250254,I250271,I250288,I370787,I370784,I250305,I250322,I250339,I250110,I250095,I250384,I250089,I250415,I250092,I250446,I250463,I250098,I250494,I250107,I250104,I250539,I250101,I250594,I250611,I250628,I250645,I250662,I250679,I250696,I250713,I250730,I250747,I250764,I250781,I250798,I250815,I250860,I250891,I250922,I250939,I250970,I251015,I251070,I251087,I251104,I251121,I251138,I251155,I251172,I251189,I251206,I251223,I251240,I251257,I251274,I251291,I251336,I251367,I251398,I251415,I251446,I251491,I251546,I251563,I308875,I308896,I251580,I308881,I251597,I308893,I251614,I308884,I251631,I308878,I251648,I251665,I251682,I251699,I251716,I308887,I308890,I251733,I251750,I251767,I251812,I251843,I251874,I251891,I251922,I251967,I252022,I252039,I252056,I252073,I252090,I252107,I252124,I252141,I252158,I252175,I252192,I252209,I252226,I252243,I252288,I252319,I252350,I252367,I252398,I252443,I252498,I252515,I404367,I404370,I252532,I252549,I404364,I404382,I252566,I252583,I404373,I252600,I252617,I252634,I252651,I252668,I404379,I404376,I252685,I252702,I252719,I252490,I252475,I252764,I252469,I252795,I252472,I252826,I252843,I252478,I252874,I252487,I252484,I252919,I252481,I252974,I252991,I253008,I253025,I253042,I253059,I253076,I253093,I253110,I253127,I253144,I253161,I253178,I253195,I252966,I252951,I253240,I252945,I253271,I252948,I253302,I253319,I252954,I253350,I252963,I252960,I253395,I252957,I253450,I253467,I253484,I253501,I253518,I253535,I253552,I253569,I253586,I253603,I253620,I253637,I253654,I253671,I253442,I253427,I253716,I253421,I253747,I253424,I253778,I253795,I253430,I253826,I253439,I253436,I253871,I253433,I253926,I253943,I306767,I306788,I253960,I306773,I253977,I306785,I253994,I306776,I254011,I306770,I254028,I254045,I254062,I254079,I254096,I306779,I306782,I254113,I254130,I254147,I254192,I254223,I254254,I254271,I254302,I254347,I254402,I254419,I390223,I390226,I254436,I254453,I390220,I390238,I254470,I254487,I390229,I254504,I254521,I254538,I254555,I254572,I390235,I390232,I254589,I254606,I254623,I254668,I254699,I254730,I254747,I254778,I254823,I254878,I254895,I406135,I406138,I254912,I254929,I406132,I406150,I254946,I254963,I406141,I254980,I254997,I255014,I255031,I255048,I406147,I406144,I255065,I255082,I255099,I255144,I255175,I255206,I255223,I255254,I255299,I255354,I255371,I320469,I320490,I255388,I320475,I255405,I320487,I255422,I320478,I255439,I320472,I255456,I255473,I255490,I255507,I255524,I320481,I320484,I255541,I255558,I255575,I255620,I255651,I255682,I255699,I255730,I255775,I255830,I255847,I255864,I255881,I255898,I255915,I255932,I255949,I255966,I255983,I256000,I256017,I256034,I256051,I255822,I255807,I256096,I255801,I256127,I255804,I256158,I256175,I255810,I256206,I255819,I255816,I256251,I255813,I256306,I256323,I286744,I286741,I256340,I286750,I256357,I286762,I286747,I256374,I256391,I286753,I256408,I256425,I256442,I256459,I256476,I286759,I256493,I286756,I256510,I256527,I256572,I256603,I256634,I256651,I256682,I256727,I256782,I256799,I314672,I314693,I256816,I314678,I256833,I314690,I256850,I314681,I256867,I314675,I256884,I256901,I256918,I256935,I256952,I314684,I314687,I256969,I256986,I257003,I256774,I256759,I257048,I256753,I257079,I256756,I257110,I257127,I256762,I257158,I256771,I256768,I257203,I256765,I257258,I257275,I257292,I257309,I257326,I257343,I257360,I257377,I257394,I257411,I257428,I257445,I257462,I257479,I257524,I257555,I257586,I257603,I257634,I257679,I257734,I257751,I373427,I373430,I257768,I257785,I373424,I373442,I257802,I257819,I373433,I257836,I257853,I257870,I257887,I257904,I373439,I373436,I257921,I257938,I257955,I258000,I258031,I258062,I258079,I258110,I258155,I258210,I258227,I258244,I258261,I258278,I258295,I258312,I258329,I258346,I258363,I258380,I258397,I258414,I258431,I258202,I258187,I258476,I258181,I258507,I258184,I258538,I258555,I258190,I258586,I258199,I258196,I258631,I258193,I258686,I258703,I258720,I258737,I258754,I258771,I258788,I258805,I258822,I258839,I258856,I258873,I258890,I258907,I258952,I258983,I259014,I259031,I259062,I259107,I259162,I259179,I317307,I317328,I259196,I317313,I259213,I317325,I259230,I317316,I259247,I317310,I259264,I259281,I259298,I259315,I259332,I317319,I317322,I259349,I259366,I259383,I259428,I259459,I259490,I259507,I259538,I259583,I259638,I259655,I259672,I259689,I259706,I259723,I259740,I259757,I259774,I259791,I259808,I259825,I259842,I259859,I259904,I259935,I259966,I259983,I260014,I260059,I260114,I260131,I374311,I374314,I260148,I260165,I374308,I374326,I260182,I260199,I374317,I260216,I260233,I260250,I260267,I260284,I374323,I374320,I260301,I260318,I260335,I260106,I260091,I260380,I260085,I260411,I260088,I260442,I260459,I260094,I260490,I260103,I260100,I260535,I260097,I260590,I260607,I260624,I260641,I260658,I260675,I260692,I260709,I260726,I260743,I260760,I260777,I260794,I260811,I260856,I260887,I260918,I260935,I260966,I261011,I261066,I261083,I376521,I376524,I261100,I261117,I376518,I376536,I261134,I261151,I376527,I261168,I261185,I261202,I261219,I261236,I376533,I376530,I261253,I261270,I261287,I261332,I261363,I261394,I261411,I261442,I261487,I261542,I261559,I261576,I261593,I261610,I261627,I261644,I261661,I261678,I261695,I261712,I261729,I261746,I261763,I261808,I261839,I261870,I261887,I261918,I261963,I262018,I262035,I262052,I262069,I262086,I262103,I262120,I262137,I262154,I262171,I262188,I262205,I262222,I262239,I262010,I261995,I262284,I261989,I262315,I261992,I262346,I262363,I261998,I262394,I262007,I262004,I262439,I262001,I262494,I262511,I262528,I262545,I262562,I262579,I262596,I262613,I262630,I262647,I262664,I262681,I262698,I262715,I262760,I262791,I262822,I262839,I262870,I262915,I262970,I262987,I263004,I263021,I263038,I263055,I263072,I263089,I263106,I263123,I263140,I263157,I263174,I263191,I262962,I262947,I263236,I262941,I263267,I262944,I263298,I263315,I262950,I263346,I262959,I262956,I263391,I262953,I263446,I263463,I263480,I263497,I263514,I263531,I263548,I263565,I263582,I263599,I263616,I263633,I263650,I263667,I263438,I263423,I263712,I263417,I263743,I263420,I263774,I263791,I263426,I263822,I263435,I263432,I263867,I263429,I263922,I263939,I263956,I263973,I263990,I264007,I264024,I264041,I264058,I264075,I264092,I264109,I264126,I264143,I264188,I264219,I264250,I264267,I264298,I264343,I264398,I264415,I264432,I264449,I264466,I264483,I264500,I264517,I264534,I264551,I264568,I264585,I264602,I264619,I264390,I264375,I264664,I264369,I264695,I264372,I264726,I264743,I264378,I264774,I264387,I264384,I264819,I264381,I264874,I264891,I264908,I264925,I264942,I264959,I264976,I264993,I265010,I265027,I265044,I265061,I265078,I265095,I265140,I265171,I265202,I265219,I265250,I265295,I265350,I265367,I265384,I265401,I265418,I265435,I265452,I265469,I265486,I265503,I265520,I265537,I265554,I265571,I265342,I265327,I265616,I265321,I265647,I265324,I265678,I265695,I265330,I265726,I265339,I265336,I265771,I265333,I265826,I265843,I265860,I265877,I265894,I265911,I265928,I265945,I265962,I265979,I265996,I266013,I266030,I266047,I266092,I266123,I266154,I266171,I266202,I266247,I266302,I266319,I266336,I266353,I266370,I266387,I266404,I266421,I266438,I266455,I266472,I266489,I266506,I266523,I266568,I266599,I266630,I266647,I266678,I266723,I266778,I266795,I266812,I266829,I266846,I266863,I266880,I266897,I266914,I266931,I266948,I266965,I266982,I266999,I266770,I266755,I267044,I266749,I267075,I266752,I267106,I267123,I266758,I267154,I266767,I266764,I267199,I266761,I267254,I267271,I267288,I267305,I267322,I267339,I267356,I267373,I267390,I267407,I267424,I267441,I267458,I267475,I267246,I267231,I267520,I267225,I267551,I267228,I267582,I267599,I267234,I267630,I267243,I267240,I267675,I267237,I267730,I267747,I293068,I293065,I267764,I293074,I267781,I293086,I293071,I267798,I267815,I293077,I267832,I267849,I267866,I267883,I267900,I293083,I267917,I293080,I267934,I267951,I267996,I268027,I268058,I268075,I268106,I268151,I268206,I268223,I268240,I268257,I268274,I268291,I268308,I268325,I268342,I268359,I268376,I268393,I268410,I268427,I268472,I268503,I268534,I268551,I268582,I268627,I268682,I268699,I343657,I343678,I268716,I343663,I268733,I343675,I268750,I343666,I268767,I343660,I268784,I268801,I268818,I268835,I268852,I343669,I343672,I268869,I268886,I268903,I268948,I268979,I269010,I269027,I269058,I269103,I269158,I269175,I269192,I269209,I269226,I269243,I269260,I269277,I269294,I269311,I269328,I269345,I269362,I269379,I269150,I269135,I269424,I269129,I269455,I269132,I269486,I269503,I269138,I269534,I269147,I269144,I269579,I269141,I269634,I269651,I269668,I269685,I269702,I269719,I269736,I269753,I269770,I269787,I269804,I269821,I269838,I269855,I269900,I269931,I269962,I269979,I270010,I270055,I270110,I270127,I365471,I365474,I270144,I270161,I365468,I365486,I270178,I270195,I365477,I270212,I270229,I270246,I270263,I270280,I365483,I365480,I270297,I270314,I270331,I270102,I270087,I270376,I270081,I270407,I270084,I270438,I270455,I270090,I270486,I270099,I270096,I270531,I270093,I270586,I270603,I270620,I270637,I270654,I270671,I270688,I270705,I270722,I270739,I270756,I270773,I270790,I270807,I270852,I270883,I270914,I270931,I270962,I271007,I271062,I271079,I385361,I385364,I271096,I271113,I385358,I385376,I271130,I271147,I385367,I271164,I271181,I271198,I271215,I271232,I385373,I385370,I271249,I271266,I271283,I271054,I271039,I271328,I271033,I271359,I271036,I271390,I271407,I271042,I271438,I271051,I271048,I271483,I271045,I271538,I271555,I271572,I271589,I271606,I271623,I271640,I271657,I271674,I271691,I271708,I271725,I271742,I271759,I271530,I271515,I271804,I271509,I271835,I271512,I271866,I271883,I271518,I271914,I271527,I271524,I271959,I271521,I272014,I272031,I272048,I272065,I272082,I272099,I272116,I272133,I272150,I272167,I272184,I272201,I272218,I272235,I272280,I272311,I272342,I272359,I272390,I272435,I272490,I272507,I272524,I272541,I272558,I272575,I272592,I272609,I272626,I272643,I272660,I272677,I272694,I272711,I272756,I272787,I272818,I272835,I272866,I272911,I272966,I272983,I273000,I273017,I273034,I273051,I273068,I273085,I273102,I273119,I273136,I273153,I273170,I273187,I272958,I272943,I273232,I272937,I273263,I272940,I273294,I273311,I272946,I273342,I272955,I272952,I273387,I272949,I273442,I273459,I310983,I311004,I273476,I310989,I273493,I311001,I273510,I310992,I273527,I310986,I273544,I273561,I273578,I273595,I273612,I310995,I310998,I273629,I273646,I273663,I273708,I273739,I273770,I273787,I273818,I273863,I273918,I273935,I401273,I401276,I273952,I273969,I401270,I401288,I273986,I274003,I401279,I274020,I274037,I274054,I274071,I274088,I401285,I401282,I274105,I274122,I274139,I273910,I273895,I274184,I273889,I274215,I273892,I274246,I274263,I273898,I274294,I273907,I273904,I274339,I273901,I274394,I274411,I274428,I274445,I274462,I274479,I274496,I274513,I274530,I274547,I274564,I274581,I274598,I274615,I274660,I274691,I274722,I274739,I274770,I274815,I274870,I274887,I274904,I274921,I274938,I274955,I274972,I274989,I275006,I275023,I275040,I275057,I275074,I275091,I274862,I274847,I275136,I274841,I275167,I274844,I275198,I275215,I274850,I275246,I274859,I274856,I275291,I274853,I275346,I275363,I275380,I275397,I275414,I275431,I275448,I275465,I275482,I275499,I275516,I275533,I275550,I275567,I275612,I275643,I275674,I275691,I275722,I275767,I275822,I275839,I275856,I275873,I275890,I275907,I275924,I275941,I275958,I275975,I275992,I276009,I276026,I276043,I276088,I276119,I276150,I276167,I276198,I276243,I276298,I276315,I276332,I276349,I276366,I276383,I276400,I276417,I276434,I276451,I276468,I276485,I276502,I276519,I276564,I276595,I276626,I276643,I276674,I276719,I276774,I276791,I276808,I276825,I276842,I276859,I276876,I276893,I276910,I276927,I276944,I276961,I276978,I276995,I277040,I277071,I277102,I277119,I277150,I277195,I277250,I277267,I277284,I277301,I277318,I277335,I277352,I277369,I277386,I277403,I277420,I277437,I277454,I277471,I277516,I277547,I277578,I277595,I277626,I277671,I277726,I277743,I310456,I310477,I277760,I310462,I277777,I310474,I277794,I310465,I277811,I310459,I277828,I277845,I277862,I277879,I277896,I310468,I310471,I277913,I277930,I277947,I277992,I278023,I278054,I278071,I278102,I278147,I278202,I278219,I314145,I314166,I278236,I314151,I278253,I314163,I278270,I314154,I278287,I314148,I278304,I278321,I278338,I278355,I278372,I314157,I314160,I278389,I278406,I278423,I278468,I278499,I278530,I278547,I278578,I278623,I278678,I278695,I403041,I403044,I278712,I278729,I403038,I403056,I278746,I278763,I403047,I278780,I278797,I278814,I278831,I278848,I403053,I403050,I278865,I278882,I278899,I278670,I278655,I278944,I278649,I278975,I278652,I279006,I279023,I278658,I279054,I278667,I278664,I279099,I278661,I279154,I279171,I399505,I399508,I279188,I279205,I399502,I399520,I279222,I279239,I399511,I279256,I279273,I279290,I279307,I279324,I399517,I399514,I279341,I279358,I279375,I279146,I279131,I279420,I279125,I279451,I279128,I279482,I279499,I279134,I279530,I279143,I279140,I279575,I279137,I279630,I279647,I327847,I327868,I279664,I327853,I279681,I327865,I279698,I327856,I279715,I327850,I279732,I279749,I279766,I279783,I279800,I327859,I327862,I279817,I279834,I279851,I279622,I279607,I279896,I279601,I279927,I279604,I279958,I279975,I279610,I280006,I279619,I279616,I280051,I279613,I280106,I280123,I387571,I387574,I280140,I280157,I387568,I387586,I280174,I280191,I387577,I280208,I280225,I280242,I280259,I280276,I387583,I387580,I280293,I280310,I280327,I280098,I280083,I280372,I280077,I280403,I280080,I280434,I280451,I280086,I280482,I280095,I280092,I280527,I280089,I280582,I280599,I280616,I280633,I280650,I280667,I280684,I280701,I280718,I280735,I280752,I280769,I280786,I280803,I280848,I280879,I280910,I280927,I280958,I281003,I281058,I281075,I407903,I407906,I281092,I281109,I407900,I407918,I281126,I281143,I407909,I281160,I281177,I281194,I281211,I281228,I407915,I407912,I281245,I281262,I281279,I281324,I281355,I281386,I281403,I281434,I281479,I281534,I281551,I281568,I281585,I281602,I281619,I281636,I281653,I281670,I281687,I281704,I281721,I281738,I281755,I281800,I281831,I281862,I281879,I281910,I281955,I282010,I282027,I388455,I388458,I282044,I282061,I388452,I388470,I282078,I282095,I388461,I282112,I282129,I282146,I282163,I282180,I388467,I388464,I282197,I282214,I282231,I282002,I281987,I282276,I281981,I282307,I281984,I282338,I282355,I281990,I282386,I281999,I281996,I282431,I281993,I282486,I282503,I382709,I382712,I282520,I282537,I382706,I382724,I282554,I282571,I382715,I282588,I282605,I282622,I282639,I282656,I382721,I382718,I282673,I282690,I282707,I282752,I282783,I282814,I282831,I282862,I282907,I282962,I282979,I297284,I297281,I282996,I297290,I283013,I297302,I297287,I283030,I283047,I297293,I283064,I283081,I283098,I283115,I283132,I297299,I283149,I297296,I283166,I283183,I283228,I283259,I283290,I283307,I283338,I283383,I283438,I283455,I283472,I283489,I283506,I283523,I283540,I283557,I283574,I283591,I283608,I283625,I283642,I283659,I283430,I283415,I283704,I283409,I283735,I283412,I283766,I283783,I283418,I283814,I283427,I283424,I283859,I283421,I283914,I283931,I283948,I283965,I283982,I283999,I284016,I284033,I284050,I284067,I284084,I284101,I284118,I284135,I284180,I284211,I284242,I284259,I284290,I284335,I284390,I284407,I284424,I284441,I284458,I284475,I284492,I284509,I284526,I284543,I284560,I284577,I284594,I284611,I284382,I284367,I284656,I284361,I284687,I284364,I284718,I284735,I284370,I284766,I284379,I284376,I284811,I284373,I284866,I284883,I391991,I391994,I284900,I284917,I391988,I392006,I284934,I284951,I391997,I284968,I284985,I285002,I285019,I285036,I392003,I392000,I285053,I285070,I285087,I284858,I284843,I285132,I284837,I285163,I284840,I285194,I285211,I284846,I285242,I284855,I284852,I285287,I284849,I285342,I285359,I285376,I285393,I285410,I285427,I285444,I285461,I285478,I285495,I285512,I285529,I285546,I285563,I285334,I285319,I285608,I285313,I285639,I285316,I285670,I285687,I285322,I285718,I285331,I285328,I285763,I285325,I285818,I285835,I285852,I285869,I285886,I285903,I285920,I285937,I285954,I285971,I285988,I286005,I286022,I286039,I286084,I286115,I286146,I286163,I286194,I286239,I286294,I286311,I286328,I286345,I286362,I286379,I286396,I286413,I286430,I286447,I286464,I286481,I286498,I286515,I286560,I286591,I286622,I286639,I286670,I286715,I286770,I286787,I286804,I286821,I286838,I286855,I286872,I286889,I286906,I286923,I286954,I286971,I286988,I287005,I287022,I287039,I287070,I287129,I287146,I287163,I287194,I287211,I287242,I287297,I287314,I287331,I287348,I287365,I287382,I287399,I287416,I287433,I287450,I287481,I287498,I287515,I287532,I287549,I287566,I287597,I287656,I287673,I287690,I287721,I287738,I287769,I287824,I287841,I287858,I287875,I287892,I287909,I287926,I287943,I287960,I287977,I287801,I288008,I288025,I288042,I288059,I288076,I288093,I287795,I288124,I287816,I287798,I287810,I288183,I288200,I288217,I287804,I288248,I288265,I287813,I288296,I287807,I288351,I288368,I337333,I337345,I288385,I337348,I337351,I288402,I288419,I288436,I288453,I337336,I288470,I337339,I288487,I288504,I288328,I288535,I288552,I288569,I288586,I337342,I288603,I337354,I288620,I288322,I288651,I288343,I288325,I288337,I288710,I288727,I288744,I288331,I288775,I288792,I288340,I288823,I288334,I288878,I288895,I349981,I349993,I288912,I349996,I349999,I288929,I288946,I288963,I288980,I349984,I288997,I349987,I289014,I289031,I288855,I289062,I289079,I289096,I289113,I349990,I289130,I350002,I289147,I288849,I289178,I288870,I288852,I288864,I289237,I289254,I289271,I288858,I289302,I289319,I288867,I289350,I288861,I289405,I289422,I289439,I289456,I289473,I289490,I289507,I289524,I289541,I289558,I289589,I289606,I289623,I289640,I289657,I289674,I289705,I289764,I289781,I289798,I289829,I289846,I289877,I289932,I289949,I389336,I389339,I289966,I389345,I389342,I289983,I290000,I290017,I290034,I389351,I290051,I290068,I290085,I290116,I290133,I290150,I290167,I290184,I389348,I290201,I290232,I290291,I389354,I290308,I290325,I290356,I290373,I290404,I290459,I290476,I290493,I290510,I290527,I290544,I290561,I290578,I290595,I290612,I290643,I290660,I290677,I290694,I290711,I290728,I290759,I290818,I290835,I290852,I290883,I290900,I290931,I290986,I291003,I291020,I291037,I291054,I291071,I291088,I291105,I291122,I291139,I291170,I291187,I291204,I291221,I291238,I291255,I291286,I291345,I291362,I291379,I291410,I291427,I291458,I291513,I291530,I291547,I291564,I291581,I291598,I291615,I291632,I291649,I291666,I291697,I291714,I291731,I291748,I291765,I291782,I291813,I291872,I291889,I291906,I291937,I291954,I291985,I292040,I292057,I292074,I292091,I292108,I292125,I292142,I292159,I292176,I292193,I292224,I292241,I292258,I292275,I292292,I292309,I292340,I292399,I292416,I292433,I292464,I292481,I292512,I292567,I292584,I292601,I292618,I292635,I292652,I292669,I292686,I292703,I292720,I292751,I292768,I292785,I292802,I292819,I292836,I292867,I292926,I292943,I292960,I292991,I293008,I293039,I293094,I293111,I293128,I293145,I293162,I293179,I293196,I293213,I293230,I293247,I293278,I293295,I293312,I293329,I293346,I293363,I293394,I293453,I293470,I293487,I293518,I293535,I293566,I293621,I293638,I293655,I293672,I293689,I293706,I293723,I293740,I293757,I293774,I293598,I293805,I293822,I293839,I293856,I293873,I293890,I293592,I293921,I293613,I293595,I293607,I293980,I293997,I294014,I293601,I294045,I294062,I293610,I294093,I293604,I294148,I294165,I294182,I294199,I294216,I294233,I294250,I294267,I294284,I294301,I294332,I294349,I294366,I294383,I294400,I294417,I294448,I294507,I294524,I294541,I294572,I294589,I294620,I294675,I294692,I294709,I294726,I294743,I294760,I294777,I294794,I294811,I294828,I294859,I294876,I294893,I294910,I294927,I294944,I294975,I295034,I295051,I295068,I295099,I295116,I295147,I295202,I295219,I295236,I295253,I295270,I295287,I295304,I295321,I295338,I295355,I295179,I295386,I295403,I295420,I295437,I295454,I295471,I295173,I295502,I295194,I295176,I295188,I295561,I295578,I295595,I295182,I295626,I295643,I295191,I295674,I295185,I295729,I295746,I295763,I295780,I295797,I295814,I295831,I295848,I295865,I295882,I295706,I295913,I295930,I295947,I295964,I295981,I295998,I295700,I296029,I295721,I295703,I295715,I296088,I296105,I296122,I295709,I296153,I296170,I295718,I296201,I295712,I296256,I296273,I365910,I365913,I296290,I365919,I365916,I296307,I296324,I296341,I296358,I365925,I296375,I296392,I296409,I296233,I296440,I296457,I296474,I296491,I296508,I365922,I296525,I296227,I296556,I296248,I296230,I296242,I296615,I365928,I296632,I296649,I296236,I296680,I296697,I296245,I296728,I296239,I296783,I296800,I409668,I409671,I296817,I409677,I409674,I296834,I296851,I296868,I296885,I409683,I296902,I296919,I296936,I296967,I296984,I297001,I297018,I297035,I409680,I297052,I297083,I297142,I409686,I297159,I297176,I297207,I297224,I297255,I297310,I297327,I297344,I297361,I297378,I297395,I297412,I297429,I297446,I297463,I297494,I297511,I297528,I297545,I297562,I297579,I297610,I297669,I297686,I297703,I297734,I297751,I297782,I297837,I297854,I297871,I297888,I297905,I297922,I297939,I297956,I297973,I297990,I298021,I298038,I298055,I298072,I298089,I298106,I298137,I298196,I298213,I298230,I298261,I298278,I298309,I298364,I298381,I340495,I340507,I298398,I340510,I340513,I298415,I298432,I298449,I298466,I340498,I298483,I340501,I298500,I298517,I298548,I298565,I298582,I298599,I340504,I298616,I340516,I298633,I298664,I298723,I298740,I298757,I298788,I298805,I298836,I298891,I298908,I298925,I298942,I298959,I298976,I298993,I299010,I299027,I299044,I299075,I299092,I299109,I299126,I299143,I299160,I299191,I299250,I299267,I299284,I299315,I299332,I299363,I299418,I299435,I375634,I375637,I299452,I375643,I375640,I299469,I299486,I299503,I299520,I375649,I299537,I299554,I299571,I299602,I299619,I299636,I299653,I299670,I375646,I299687,I299718,I299777,I375652,I299794,I299811,I299842,I299859,I299890,I299945,I299962,I299979,I299996,I300013,I300030,I300047,I300064,I300081,I300098,I300129,I300146,I300163,I300180,I300197,I300214,I300245,I300304,I300321,I300338,I300369,I300386,I300417,I300472,I300489,I300506,I300523,I300540,I300557,I300574,I300591,I300608,I300625,I300656,I300673,I300690,I300707,I300724,I300741,I300772,I300831,I300848,I300865,I300896,I300913,I300944,I300999,I301016,I392872,I392875,I301033,I392881,I392878,I301050,I301067,I301084,I301101,I392887,I301118,I301135,I301152,I300976,I301183,I301200,I301217,I301234,I301251,I392884,I301268,I300970,I301299,I300991,I300973,I300985,I301358,I392890,I301375,I301392,I300979,I301423,I301440,I300988,I301471,I300982,I301526,I301543,I301560,I301577,I301594,I301611,I301628,I301645,I301662,I301679,I301710,I301727,I301744,I301761,I301778,I301795,I301826,I301885,I301902,I301919,I301950,I301967,I301998,I302053,I302070,I302087,I302104,I302121,I302138,I302155,I302172,I302189,I302206,I302237,I302254,I302271,I302288,I302305,I302322,I302353,I302412,I302429,I302446,I302477,I302494,I302525,I302580,I302597,I302614,I302631,I302648,I302665,I302682,I302699,I302716,I302733,I302557,I302764,I302781,I302798,I302815,I302832,I302849,I302551,I302880,I302572,I302554,I302566,I302939,I302956,I302973,I302560,I303004,I303021,I302569,I303052,I302563,I303107,I303124,I303141,I303158,I303175,I303192,I303223,I303240,I303257,I303274,I303291,I303308,I303325,I303342,I303359,I303390,I303421,I303452,I303469,I303514,I303545,I303562,I303579,I303634,I303651,I303668,I303685,I303702,I303719,I303750,I303767,I303784,I303801,I303818,I303835,I303852,I303869,I303886,I303917,I303948,I303979,I303996,I304041,I304072,I304089,I304106,I304161,I304178,I304195,I304212,I304229,I304246,I304277,I304294,I304311,I304328,I304345,I304362,I304379,I304396,I304413,I304444,I304475,I304506,I304523,I304568,I304599,I304616,I304633,I304688,I304705,I397734,I397737,I304722,I397749,I304739,I397740,I304756,I304773,I304804,I304821,I397743,I304838,I304855,I397746,I304872,I304889,I304906,I397752,I304923,I304940,I304971,I305002,I305033,I305050,I305095,I305126,I305143,I305160,I305215,I305232,I305249,I305266,I305283,I305300,I305331,I305348,I305365,I305382,I305399,I305416,I305433,I305450,I305467,I305498,I305529,I305560,I305577,I305622,I305653,I305670,I305687,I305742,I305759,I305776,I305793,I305810,I305827,I305858,I305875,I305892,I305909,I305926,I305943,I305960,I305977,I305994,I306025,I306056,I306087,I306104,I306149,I306180,I306197,I306214,I306269,I306286,I362816,I362819,I306303,I362831,I306320,I362822,I306337,I306354,I306385,I306402,I362825,I306419,I306436,I362828,I306453,I306470,I306487,I362834,I306504,I306521,I306552,I306583,I306614,I306631,I306676,I306707,I306724,I306741,I306796,I306813,I306830,I306847,I306864,I306881,I306912,I306929,I306946,I306963,I306980,I306997,I307014,I307031,I307048,I307079,I307110,I307141,I307158,I307203,I307234,I307251,I307268,I307323,I307340,I307357,I307374,I307391,I307408,I307439,I307456,I307473,I307490,I307507,I307524,I307541,I307558,I307575,I307606,I307637,I307668,I307685,I307730,I307761,I307778,I307795,I307850,I307867,I307884,I307901,I307918,I307935,I307966,I307983,I308000,I308017,I308034,I308051,I308068,I308085,I308102,I308133,I308164,I308195,I308212,I308257,I308288,I308305,I308322,I308377,I308394,I308411,I308428,I308445,I308462,I308493,I308510,I308527,I308544,I308561,I308578,I308595,I308612,I308629,I308660,I308691,I308722,I308739,I308784,I308815,I308832,I308849,I308904,I308921,I308938,I308955,I308972,I308989,I309020,I309037,I309054,I309071,I309088,I309105,I309122,I309139,I309156,I309187,I309218,I309249,I309266,I309311,I309342,I309359,I309376,I309431,I309448,I309465,I309482,I309499,I309516,I309547,I309564,I309581,I309598,I309615,I309632,I309649,I309666,I309683,I309714,I309745,I309776,I309793,I309838,I309869,I309886,I309903,I309958,I309975,I309992,I310009,I310026,I310043,I310074,I310091,I310108,I310125,I310142,I310159,I310176,I310193,I310210,I310241,I310272,I310303,I310320,I310365,I310396,I310413,I310430,I310485,I310502,I371656,I371659,I310519,I371671,I310536,I371662,I310553,I310570,I310601,I310618,I371665,I310635,I310652,I371668,I310669,I310686,I310703,I371674,I310720,I310737,I310768,I310799,I310830,I310847,I310892,I310923,I310940,I310957,I311012,I311029,I311046,I311063,I311080,I311097,I311128,I311145,I311162,I311179,I311196,I311213,I311230,I311247,I311264,I311295,I311326,I311357,I311374,I311419,I311450,I311467,I311484,I311539,I311556,I311573,I311590,I311607,I311624,I311655,I311672,I311689,I311706,I311723,I311740,I311757,I311774,I311791,I311822,I311853,I311884,I311901,I311946,I311977,I311994,I312011,I312066,I312083,I312100,I312117,I312134,I312151,I312182,I312199,I312216,I312233,I312250,I312267,I312284,I312301,I312318,I312349,I312380,I312411,I312428,I312473,I312504,I312521,I312538,I312593,I312610,I312627,I312644,I312661,I312678,I312567,I312709,I312726,I312743,I312760,I312777,I312794,I312811,I312828,I312845,I312564,I312876,I312579,I312907,I312576,I312938,I312955,I312582,I312585,I313000,I312570,I313031,I313048,I313065,I312573,I313120,I313137,I313154,I313171,I313188,I313205,I313236,I313253,I313270,I313287,I313304,I313321,I313338,I313355,I313372,I313403,I313434,I313465,I313482,I313527,I313558,I313575,I313592,I313647,I313664,I313681,I313698,I313715,I313732,I313763,I313780,I313797,I313814,I313831,I313848,I313865,I313882,I313899,I313930,I313961,I313992,I314009,I314054,I314085,I314102,I314119,I314174,I314191,I314208,I314225,I314242,I314259,I314290,I314307,I314324,I314341,I314358,I314375,I314392,I314409,I314426,I314457,I314488,I314519,I314536,I314581,I314612,I314629,I314646,I314701,I314718,I314735,I314752,I314769,I314786,I314817,I314834,I314851,I314868,I314885,I314902,I314919,I314936,I314953,I314984,I315015,I315046,I315063,I315108,I315139,I315156,I315173,I315228,I315245,I379612,I379615,I315262,I379627,I315279,I379618,I315296,I315313,I315344,I315361,I379621,I315378,I315395,I379624,I315412,I315429,I315446,I379630,I315463,I315480,I315511,I315542,I315573,I315590,I315635,I315666,I315683,I315700,I315755,I315772,I315789,I315806,I315823,I315840,I315871,I315888,I315905,I315922,I315939,I315956,I315973,I315990,I316007,I316038,I316069,I316100,I316117,I316162,I316193,I316210,I316227,I316282,I316299,I316316,I316333,I316350,I316367,I316398,I316415,I316432,I316449,I316466,I316483,I316500,I316517,I316534,I316565,I316596,I316627,I316644,I316689,I316720,I316737,I316754,I316809,I316826,I316843,I316860,I316877,I316894,I316783,I316925,I316942,I316959,I316976,I316993,I317010,I317027,I317044,I317061,I316780,I317092,I316795,I317123,I316792,I317154,I317171,I316798,I316801,I317216,I316786,I317247,I317264,I317281,I316789,I317336,I317353,I317370,I317387,I317404,I317421,I317452,I317469,I317486,I317503,I317520,I317537,I317554,I317571,I317588,I317619,I317650,I317681,I317698,I317743,I317774,I317791,I317808,I317863,I317880,I317897,I317914,I317931,I317948,I317979,I317996,I318013,I318030,I318047,I318064,I318081,I318098,I318115,I318146,I318177,I318208,I318225,I318270,I318301,I318318,I318335,I318390,I318407,I318424,I318441,I318458,I318475,I318506,I318523,I318540,I318557,I318574,I318591,I318608,I318625,I318642,I318673,I318704,I318735,I318752,I318797,I318828,I318845,I318862,I318917,I318934,I318951,I318968,I318985,I319002,I318891,I319033,I319050,I319067,I319084,I319101,I319118,I319135,I319152,I319169,I318888,I319200,I318903,I319231,I318900,I319262,I319279,I318906,I318909,I319324,I318894,I319355,I319372,I319389,I318897,I319444,I319461,I319478,I319495,I319512,I319529,I319560,I319577,I319594,I319611,I319628,I319645,I319662,I319679,I319696,I319727,I319758,I319789,I319806,I319851,I319882,I319899,I319916,I319971,I319988,I320005,I320022,I320039,I320056,I320087,I320104,I320121,I320138,I320155,I320172,I320189,I320206,I320223,I320254,I320285,I320316,I320333,I320378,I320409,I320426,I320443,I320498,I320515,I320532,I320549,I320566,I320583,I320614,I320631,I320648,I320665,I320682,I320699,I320716,I320733,I320750,I320781,I320812,I320843,I320860,I320905,I320936,I320953,I320970,I321025,I321042,I321059,I321076,I321093,I321110,I320999,I321141,I321158,I321175,I321192,I321209,I321226,I321243,I321260,I321277,I320996,I321308,I321011,I321339,I321008,I321370,I321387,I321014,I321017,I321432,I321002,I321463,I321480,I321497,I321005,I321552,I321569,I321586,I321603,I321620,I321637,I321668,I321685,I321702,I321719,I321736,I321753,I321770,I321787,I321804,I321835,I321866,I321897,I321914,I321959,I321990,I322007,I322024,I322079,I322096,I322113,I322130,I322147,I322164,I322195,I322212,I322229,I322246,I322263,I322280,I322297,I322314,I322331,I322362,I322393,I322424,I322441,I322486,I322517,I322534,I322551,I322606,I322623,I322640,I322657,I322674,I322691,I322722,I322739,I322756,I322773,I322790,I322807,I322824,I322841,I322858,I322889,I322920,I322951,I322968,I323013,I323044,I323061,I323078,I323133,I323150,I392430,I392433,I323167,I392445,I323184,I392436,I323201,I323218,I323107,I323249,I323266,I392439,I323283,I323300,I392442,I323317,I323334,I323351,I392448,I323368,I323385,I323104,I323416,I323119,I323447,I323116,I323478,I323495,I323122,I323125,I323540,I323110,I323571,I323588,I323605,I323113,I323660,I323677,I323694,I323711,I323728,I323745,I323776,I323793,I323810,I323827,I323844,I323861,I323878,I323895,I323912,I323943,I323974,I324005,I324022,I324067,I324098,I324115,I324132,I324187,I324204,I391104,I391107,I324221,I391119,I324238,I391110,I324255,I324272,I324303,I324320,I391113,I324337,I324354,I391116,I324371,I324388,I324405,I391122,I324422,I324439,I324470,I324501,I324532,I324549,I324594,I324625,I324642,I324659,I324714,I324731,I324748,I324765,I324782,I324799,I324830,I324847,I324864,I324881,I324898,I324915,I324932,I324949,I324966,I324997,I325028,I325059,I325076,I325121,I325152,I325169,I325186,I325241,I325258,I325275,I325292,I325309,I325326,I325357,I325374,I325391,I325408,I325425,I325442,I325459,I325476,I325493,I325524,I325555,I325586,I325603,I325648,I325679,I325696,I325713,I325768,I325785,I325802,I325819,I325836,I325853,I325884,I325901,I325918,I325935,I325952,I325969,I325986,I326003,I326020,I326051,I326082,I326113,I326130,I326175,I326206,I326223,I326240,I326295,I326312,I367236,I367239,I326329,I367251,I326346,I367242,I326363,I326380,I326269,I326411,I326428,I367245,I326445,I326462,I367248,I326479,I326496,I326513,I367254,I326530,I326547,I326266,I326578,I326281,I326609,I326278,I326640,I326657,I326284,I326287,I326702,I326272,I326733,I326750,I326767,I326275,I326822,I326839,I326856,I326873,I326890,I326907,I326938,I326955,I326972,I326989,I327006,I327023,I327040,I327057,I327074,I327105,I327136,I327167,I327184,I327229,I327260,I327277,I327294,I327349,I327366,I327383,I327400,I327417,I327434,I327465,I327482,I327499,I327516,I327533,I327550,I327567,I327584,I327601,I327632,I327663,I327694,I327711,I327756,I327787,I327804,I327821,I327876,I327893,I327910,I327927,I327944,I327961,I327992,I328009,I328026,I328043,I328060,I328077,I328094,I328111,I328128,I328159,I328190,I328221,I328238,I328283,I328314,I328331,I328348,I328403,I328420,I328437,I328454,I328471,I328488,I328377,I328519,I328536,I328553,I328570,I328587,I328604,I328621,I328638,I328655,I328374,I328686,I328389,I328717,I328386,I328748,I328765,I328392,I328395,I328810,I328380,I328841,I328858,I328875,I328383,I328930,I328947,I386684,I386687,I328964,I386699,I328981,I386690,I328998,I329015,I328904,I329046,I329063,I386693,I329080,I329097,I386696,I329114,I329131,I329148,I386702,I329165,I329182,I328901,I329213,I328916,I329244,I328913,I329275,I329292,I328919,I328922,I329337,I328907,I329368,I329385,I329402,I328910,I329457,I329474,I329491,I329508,I329525,I329542,I329573,I329590,I329607,I329624,I329641,I329658,I329675,I329692,I329709,I329740,I329771,I329802,I329819,I329864,I329895,I329912,I329929,I329984,I330001,I330018,I330035,I330052,I330069,I330100,I330117,I330134,I330151,I330168,I330185,I330202,I330219,I330236,I330267,I330298,I330329,I330346,I330391,I330422,I330439,I330456,I330511,I330528,I330545,I330562,I330579,I330596,I330485,I330627,I330644,I330661,I330678,I330695,I330712,I330729,I330746,I330763,I330482,I330794,I330497,I330825,I330494,I330856,I330873,I330500,I330503,I330918,I330488,I330949,I330966,I330983,I330491,I331038,I331055,I331072,I331089,I331106,I331123,I331154,I331171,I331188,I331205,I331222,I331239,I331256,I331273,I331290,I331321,I331352,I331383,I331400,I331445,I331476,I331493,I331510,I331565,I331582,I331599,I331616,I331633,I331650,I331681,I331698,I331715,I331732,I331749,I331766,I331783,I331800,I331817,I331848,I331879,I331910,I331927,I331972,I332003,I332020,I332037,I332092,I332109,I332126,I332143,I332160,I332177,I332066,I332208,I332225,I332242,I332259,I332276,I332293,I332310,I332327,I332344,I332063,I332375,I332078,I332406,I332075,I332437,I332454,I332081,I332084,I332499,I332069,I332530,I332547,I332564,I332072,I332619,I332636,I332653,I332670,I332687,I332704,I332735,I332752,I332769,I332786,I332803,I332820,I332837,I332854,I332871,I332902,I332933,I332964,I332981,I333026,I333057,I333074,I333091,I333146,I333163,I333180,I333197,I333214,I333231,I333262,I333279,I333296,I333313,I333330,I333347,I333364,I333381,I333398,I333429,I333460,I333491,I333508,I333553,I333584,I333601,I333618,I333673,I333690,I333707,I333724,I333741,I333758,I333789,I333806,I333823,I333840,I333857,I333874,I333891,I333908,I333925,I333956,I333987,I334018,I334035,I334080,I334111,I334128,I334145,I334200,I334217,I334234,I334251,I334268,I334285,I334316,I334333,I334350,I334367,I334384,I334401,I334418,I334435,I334452,I334483,I334514,I334545,I334562,I334607,I334638,I334655,I334672,I334727,I334744,I334761,I334778,I334795,I334812,I334843,I334860,I334877,I334894,I334911,I334928,I334945,I334962,I334979,I335010,I335041,I335072,I335089,I335134,I335165,I335182,I335199,I335254,I335271,I335288,I335305,I335322,I335339,I335370,I335387,I335404,I335421,I335438,I335455,I335472,I335489,I335506,I335537,I335568,I335599,I335616,I335661,I335692,I335709,I335726,I335781,I335798,I335815,I335832,I335849,I335866,I335897,I335914,I335931,I335948,I335965,I335982,I335999,I336016,I336033,I336064,I336095,I336126,I336143,I336188,I336219,I336236,I336253,I336308,I336325,I336342,I336359,I336376,I336393,I336424,I336441,I336458,I336475,I336492,I336509,I336526,I336543,I336560,I336591,I336622,I336653,I336670,I336715,I336746,I336763,I336780,I336835,I336852,I336869,I336886,I336903,I336920,I336951,I336968,I336985,I337002,I337019,I337036,I337053,I337070,I337087,I337118,I337149,I337180,I337197,I337242,I337273,I337290,I337307,I337362,I337379,I337396,I337413,I337430,I337447,I337478,I337495,I337512,I337529,I337546,I337563,I337580,I337597,I337614,I337645,I337676,I337707,I337724,I337769,I337800,I337817,I337834,I337889,I337906,I337923,I337940,I337957,I337974,I338005,I338022,I338039,I338056,I338073,I338090,I338107,I338124,I338141,I338172,I338203,I338234,I338251,I338296,I338327,I338344,I338361,I338416,I338433,I338450,I338467,I338484,I338501,I338532,I338549,I338566,I338583,I338600,I338617,I338634,I338651,I338668,I338699,I338730,I338761,I338778,I338823,I338854,I338871,I338888,I338943,I338960,I338977,I338994,I339011,I339028,I339059,I339076,I339093,I339110,I339127,I339144,I339161,I339178,I339195,I339226,I339257,I339288,I339305,I339350,I339381,I339398,I339415,I339470,I339487,I395524,I395527,I339504,I395539,I339521,I395530,I339538,I339555,I339586,I339603,I395533,I339620,I339637,I395536,I339654,I339671,I339688,I395542,I339705,I339722,I339753,I339784,I339815,I339832,I339877,I339908,I339925,I339942,I339997,I340014,I340031,I340048,I340065,I340082,I339971,I340113,I340130,I340147,I340164,I340181,I340198,I340215,I340232,I340249,I339968,I340280,I339983,I340311,I339980,I340342,I340359,I339986,I339989,I340404,I339974,I340435,I340452,I340469,I339977,I340524,I340541,I340558,I340575,I340592,I340609,I340640,I340657,I340674,I340691,I340708,I340725,I340742,I340759,I340776,I340807,I340838,I340869,I340886,I340931,I340962,I340979,I340996,I341051,I341068,I405248,I405251,I341085,I405263,I341102,I405254,I341119,I341136,I341167,I341184,I405257,I341201,I341218,I405260,I341235,I341252,I341269,I405266,I341286,I341303,I341334,I341365,I341396,I341413,I341458,I341489,I341506,I341523,I341578,I341595,I341612,I341629,I341646,I341663,I341552,I341694,I341711,I341728,I341745,I341762,I341779,I341796,I341813,I341830,I341549,I341861,I341564,I341892,I341561,I341923,I341940,I341567,I341570,I341985,I341555,I342016,I342033,I342050,I341558,I342105,I342122,I342139,I342156,I342173,I342190,I342079,I342221,I342238,I342255,I342272,I342289,I342306,I342323,I342340,I342357,I342076,I342388,I342091,I342419,I342088,I342450,I342467,I342094,I342097,I342512,I342082,I342543,I342560,I342577,I342085,I342632,I342649,I342666,I342683,I342700,I342717,I342748,I342765,I342782,I342799,I342816,I342833,I342850,I342867,I342884,I342915,I342946,I342977,I342994,I343039,I343070,I343087,I343104,I343159,I343176,I343193,I343210,I343227,I343244,I343133,I343275,I343292,I343309,I343326,I343343,I343360,I343377,I343394,I343411,I343130,I343442,I343145,I343473,I343142,I343504,I343521,I343148,I343151,I343566,I343136,I343597,I343614,I343631,I343139,I343686,I343703,I343720,I343737,I343754,I343771,I343802,I343819,I343836,I343853,I343870,I343887,I343904,I343921,I343938,I343969,I344000,I344031,I344048,I344093,I344124,I344141,I344158,I344213,I344230,I344247,I344264,I344281,I344298,I344187,I344329,I344346,I344363,I344380,I344397,I344414,I344431,I344448,I344465,I344184,I344496,I344199,I344527,I344196,I344558,I344575,I344202,I344205,I344620,I344190,I344651,I344668,I344685,I344193,I344740,I344757,I344774,I344791,I344808,I344825,I344714,I344856,I344873,I344890,I344907,I344924,I344941,I344958,I344975,I344992,I344711,I345023,I344726,I345054,I344723,I345085,I345102,I344729,I344732,I345147,I344717,I345178,I345195,I345212,I344720,I345267,I345284,I345301,I345318,I345335,I345352,I345383,I345400,I345417,I345434,I345451,I345468,I345485,I345502,I345519,I345550,I345581,I345612,I345629,I345674,I345705,I345722,I345739,I345794,I345811,I345828,I345845,I345862,I345879,I345910,I345927,I345944,I345961,I345978,I345995,I346012,I346029,I346046,I346077,I346108,I346139,I346156,I346201,I346232,I346249,I346266,I346321,I346338,I398618,I398621,I346355,I398633,I346372,I398624,I346389,I346406,I346437,I346454,I398627,I346471,I346488,I398630,I346505,I346522,I346539,I398636,I346556,I346573,I346604,I346635,I346666,I346683,I346728,I346759,I346776,I346793,I346848,I346865,I346882,I346899,I346916,I346933,I346964,I346981,I346998,I347015,I347032,I347049,I347066,I347083,I347100,I347131,I347162,I347193,I347210,I347255,I347286,I347303,I347320,I347375,I347392,I347409,I347426,I347443,I347460,I347349,I347491,I347508,I347525,I347542,I347559,I347576,I347593,I347610,I347627,I347346,I347658,I347361,I347689,I347358,I347720,I347737,I347364,I347367,I347782,I347352,I347813,I347830,I347847,I347355,I347902,I347919,I347936,I347953,I347970,I347987,I348018,I348035,I348052,I348069,I348086,I348103,I348120,I348137,I348154,I348185,I348216,I348247,I348264,I348309,I348340,I348357,I348374,I348429,I348446,I348463,I348480,I348497,I348514,I348545,I348562,I348579,I348596,I348613,I348630,I348647,I348664,I348681,I348712,I348743,I348774,I348791,I348836,I348867,I348884,I348901,I348956,I348973,I361490,I361493,I348990,I361505,I349007,I361496,I349024,I349041,I349072,I349089,I361499,I349106,I349123,I361502,I349140,I349157,I349174,I361508,I349191,I349208,I349239,I349270,I349301,I349318,I349363,I349394,I349411,I349428,I349483,I349500,I349517,I349534,I349551,I349568,I349457,I349599,I349616,I349633,I349650,I349667,I349684,I349701,I349718,I349735,I349454,I349766,I349469,I349797,I349466,I349828,I349845,I349472,I349475,I349890,I349460,I349921,I349938,I349955,I349463,I350010,I350027,I350044,I350061,I350078,I350095,I350126,I350143,I350160,I350177,I350194,I350211,I350228,I350245,I350262,I350293,I350324,I350355,I350372,I350417,I350448,I350465,I350482,I350537,I350554,I350571,I350588,I350605,I350622,I350653,I350670,I350687,I350704,I350721,I350738,I350755,I350772,I350789,I350820,I350851,I350882,I350899,I350944,I350975,I350992,I351009,I351064,I351081,I351098,I351115,I351132,I351149,I351180,I351197,I351214,I351231,I351248,I351265,I351282,I351299,I351316,I351347,I351378,I351409,I351426,I351471,I351502,I351519,I351536,I351591,I351608,I351625,I351642,I351659,I351676,I351565,I351707,I351724,I351741,I351758,I351775,I351792,I351809,I351826,I351843,I351562,I351874,I351577,I351905,I351574,I351936,I351953,I351580,I351583,I351998,I351568,I352029,I352046,I352063,I351571,I352118,I352135,I352152,I352169,I352186,I352203,I352234,I352251,I352268,I352285,I352302,I352319,I352336,I352353,I352370,I352401,I352432,I352463,I352480,I352525,I352556,I352573,I352590,I352645,I352662,I352679,I352696,I352713,I352730,I352761,I352778,I352795,I352812,I352829,I352846,I352863,I352880,I352897,I352928,I352959,I352990,I353007,I353052,I353083,I353100,I353117,I353172,I353189,I353206,I353223,I353240,I353257,I353288,I353305,I353322,I353339,I353356,I353373,I353390,I353407,I353424,I353455,I353486,I353517,I353534,I353579,I353610,I353627,I353644,I353699,I353716,I353733,I353750,I353767,I353784,I353815,I353832,I353849,I353866,I353883,I353900,I353917,I353934,I353951,I353982,I354013,I354044,I354061,I354106,I354137,I354154,I354171,I354226,I354243,I354260,I354277,I354294,I354311,I354342,I354359,I354376,I354393,I354410,I354427,I354444,I354461,I354478,I354509,I354540,I354571,I354588,I354633,I354664,I354681,I354698,I354753,I354770,I376960,I376963,I354787,I376975,I354804,I376966,I354821,I354838,I354727,I354869,I354886,I376969,I354903,I354920,I376972,I354937,I354954,I354971,I376978,I354988,I355005,I354724,I355036,I354739,I355067,I354736,I355098,I355115,I354742,I354745,I355160,I354730,I355191,I355208,I355225,I354733,I355280,I355297,I355314,I355331,I355348,I355365,I355396,I355413,I355430,I355447,I355464,I355481,I355498,I355515,I355532,I355563,I355594,I355625,I355642,I355687,I355718,I355735,I355752,I355807,I355824,I355841,I355858,I355875,I355892,I355923,I355940,I355957,I355974,I355991,I356008,I356025,I356042,I356059,I356090,I356121,I356152,I356169,I356214,I356245,I356262,I356279,I356334,I356351,I399944,I399947,I356368,I399959,I356385,I399950,I356402,I356419,I356450,I356467,I399953,I356484,I356501,I399956,I356518,I356535,I356552,I399962,I356569,I356586,I356617,I356648,I356679,I356696,I356741,I356772,I356789,I356806,I356861,I356878,I400386,I400389,I356895,I400401,I356912,I400392,I356929,I356946,I356835,I356977,I356994,I400395,I357011,I357028,I400398,I357045,I357062,I357079,I400404,I357096,I357113,I356832,I357144,I356847,I357175,I356844,I357206,I357223,I356850,I356853,I357268,I356838,I357299,I357316,I357333,I356841,I357388,I357405,I357422,I357439,I357456,I357473,I357504,I357521,I357538,I357555,I357572,I357589,I357606,I357623,I357640,I357671,I357702,I357733,I357750,I357795,I357826,I357843,I357860,I357915,I357932,I357949,I357966,I357983,I358000,I358031,I358048,I358065,I358082,I358099,I358116,I358133,I358150,I358167,I358198,I358229,I358260,I358277,I358322,I358353,I358370,I358387,I358442,I358459,I358476,I358493,I358510,I358527,I358558,I358575,I358592,I358609,I358626,I358643,I358660,I358677,I358694,I358725,I358756,I358787,I358804,I358849,I358880,I358897,I358914,I358969,I358986,I373866,I373869,I359003,I373881,I359020,I373872,I359037,I359054,I359085,I359102,I373875,I359119,I359136,I373878,I359153,I359170,I359187,I373884,I359204,I359221,I359252,I359283,I359314,I359331,I359376,I359407,I359424,I359441,I359496,I359513,I359530,I359547,I359564,I359581,I359612,I359629,I359646,I359663,I359680,I359697,I359714,I359731,I359748,I359779,I359810,I359841,I359858,I359903,I359934,I359951,I359968,I360023,I360040,I360057,I360074,I360091,I360108,I360139,I360156,I360173,I360190,I360207,I360224,I360241,I360258,I360275,I360306,I360337,I360368,I360385,I360430,I360461,I360478,I360495,I360550,I360567,I360584,I360601,I360618,I360635,I360666,I360683,I360700,I360717,I360734,I360751,I360768,I360785,I360802,I360833,I360864,I360895,I360912,I360957,I360988,I361005,I361022,I361074,I361091,I361108,I361125,I361142,I361173,I361190,I361207,I361224,I361241,I361258,I361275,I361292,I361351,I361368,I361385,I361416,I361433,I361464,I361516,I361533,I361550,I361567,I361584,I361615,I361632,I361649,I361666,I361683,I361700,I361717,I361734,I361793,I361810,I361827,I361858,I361875,I361906,I361958,I361975,I361992,I362009,I362026,I362057,I362074,I362091,I362108,I362125,I362142,I362159,I362176,I362235,I362252,I362269,I362300,I362317,I362348,I362400,I362417,I362434,I362451,I362468,I362499,I362516,I362533,I362550,I362567,I362584,I362601,I362618,I362677,I362694,I362711,I362742,I362759,I362790,I362842,I362859,I362876,I362893,I362910,I362941,I362958,I362975,I362992,I363009,I363026,I363043,I363060,I363119,I363136,I363153,I363184,I363201,I363232,I363284,I363301,I363318,I363335,I363352,I363383,I363400,I363417,I363434,I363451,I363468,I363485,I363502,I363561,I363578,I363595,I363626,I363643,I363674,I363726,I363743,I363760,I363777,I363794,I363825,I363842,I363859,I363876,I363893,I363910,I363927,I363944,I364003,I364020,I364037,I364068,I364085,I364116,I364168,I364185,I364202,I364219,I364236,I364267,I364284,I364301,I364318,I364335,I364352,I364369,I364386,I364445,I364462,I364479,I364510,I364527,I364558,I364610,I364627,I364644,I364661,I364678,I364709,I364726,I364743,I364760,I364777,I364794,I364811,I364828,I364887,I364904,I364921,I364952,I364969,I365000,I365052,I365069,I365086,I365103,I365120,I365151,I365168,I365185,I365202,I365219,I365236,I365253,I365270,I365329,I365346,I365363,I365394,I365411,I365442,I365494,I365511,I365528,I365545,I365562,I365593,I365610,I365627,I365644,I365661,I365678,I365695,I365712,I365771,I365788,I365805,I365836,I365853,I365884,I365936,I365953,I365970,I365987,I366004,I366035,I366052,I366069,I366086,I366103,I366120,I366137,I366154,I366213,I366230,I366247,I366278,I366295,I366326,I366378,I366395,I366412,I366429,I366446,I366477,I366494,I366511,I366528,I366545,I366562,I366579,I366596,I366655,I366672,I366689,I366720,I366737,I366768,I366820,I366837,I366854,I366871,I366888,I366919,I366936,I366953,I366970,I366987,I367004,I367021,I367038,I367097,I367114,I367131,I367162,I367179,I367210,I367262,I367279,I367296,I367313,I367330,I367361,I367378,I367395,I367412,I367429,I367446,I367463,I367480,I367539,I367556,I367573,I367604,I367621,I367652,I367704,I367721,I367738,I367755,I367772,I367803,I367820,I367837,I367854,I367871,I367888,I367905,I367922,I367981,I367998,I368015,I368046,I368063,I368094,I368146,I368163,I368180,I368197,I368214,I368245,I368262,I368279,I368296,I368313,I368330,I368347,I368364,I368423,I368440,I368457,I368488,I368505,I368536,I368588,I368605,I368622,I368639,I368656,I368687,I368704,I368721,I368738,I368755,I368772,I368789,I368806,I368865,I368882,I368899,I368930,I368947,I368978,I369030,I369047,I369064,I369081,I369098,I369129,I369146,I369163,I369180,I369197,I369214,I369231,I369248,I369307,I369324,I369341,I369372,I369389,I369420,I369472,I369489,I369506,I369523,I369540,I369571,I369588,I369605,I369622,I369639,I369656,I369673,I369690,I369749,I369766,I369783,I369814,I369831,I369862,I369914,I369931,I369948,I369965,I369982,I370013,I370030,I370047,I370064,I370081,I370098,I370115,I370132,I370191,I370208,I370225,I370256,I370273,I370304,I370356,I370373,I370390,I370407,I370424,I370455,I370472,I370489,I370506,I370523,I370540,I370557,I370574,I370633,I370650,I370667,I370698,I370715,I370746,I370798,I370815,I370832,I370849,I370866,I370897,I370914,I370931,I370948,I370965,I370982,I370999,I371016,I371075,I371092,I371109,I371140,I371157,I371188,I371240,I371257,I371274,I371291,I371308,I371339,I371356,I371373,I371390,I371407,I371424,I371441,I371458,I371517,I371534,I371551,I371582,I371599,I371630,I371682,I371699,I371716,I371733,I371750,I371781,I371798,I371815,I371832,I371849,I371866,I371883,I371900,I371959,I371976,I371993,I372024,I372041,I372072,I372124,I372141,I372158,I372175,I372192,I372223,I372240,I372257,I372274,I372291,I372308,I372325,I372342,I372401,I372418,I372435,I372466,I372483,I372514,I372566,I372583,I372600,I372617,I372634,I372665,I372682,I372699,I372716,I372733,I372750,I372767,I372784,I372843,I372860,I372877,I372908,I372925,I372956,I373008,I373025,I373042,I373059,I373076,I373107,I373124,I373141,I373158,I373175,I373192,I373209,I373226,I373285,I373302,I373319,I373350,I373367,I373398,I373450,I373467,I373484,I373501,I373518,I373549,I373566,I373583,I373600,I373617,I373634,I373651,I373668,I373727,I373744,I373761,I373792,I373809,I373840,I373892,I373909,I373926,I373943,I373960,I373991,I374008,I374025,I374042,I374059,I374076,I374093,I374110,I374169,I374186,I374203,I374234,I374251,I374282,I374334,I374351,I374368,I374385,I374402,I374433,I374450,I374467,I374484,I374501,I374518,I374535,I374552,I374611,I374628,I374645,I374676,I374693,I374724,I374776,I374793,I374810,I374827,I374844,I374875,I374892,I374909,I374926,I374943,I374960,I374977,I374994,I375053,I375070,I375087,I375118,I375135,I375166,I375218,I375235,I375252,I375269,I375286,I375317,I375334,I375351,I375368,I375385,I375402,I375419,I375436,I375495,I375512,I375529,I375560,I375577,I375608,I375660,I375677,I375694,I375711,I375728,I375759,I375776,I375793,I375810,I375827,I375844,I375861,I375878,I375937,I375954,I375971,I376002,I376019,I376050,I376102,I376119,I376136,I376153,I376170,I376201,I376218,I376235,I376252,I376269,I376286,I376303,I376320,I376379,I376396,I376413,I376444,I376461,I376492,I376544,I376561,I376578,I376595,I376612,I376643,I376660,I376677,I376694,I376711,I376728,I376745,I376762,I376821,I376838,I376855,I376886,I376903,I376934,I376986,I377003,I377020,I377037,I377054,I377085,I377102,I377119,I377136,I377153,I377170,I377187,I377204,I377263,I377280,I377297,I377328,I377345,I377376,I377428,I377445,I377462,I377479,I377496,I377527,I377544,I377561,I377578,I377595,I377612,I377629,I377646,I377705,I377722,I377739,I377770,I377787,I377818,I377870,I377887,I377904,I377921,I377938,I377969,I377986,I378003,I378020,I378037,I378054,I378071,I378088,I378147,I378164,I378181,I378212,I378229,I378260,I378312,I378329,I378346,I378363,I378380,I378411,I378428,I378445,I378462,I378479,I378496,I378513,I378530,I378589,I378606,I378623,I378654,I378671,I378702,I378754,I378771,I378788,I378805,I378822,I378853,I378870,I378887,I378904,I378921,I378938,I378955,I378972,I379031,I379048,I379065,I379096,I379113,I379144,I379196,I379213,I379230,I379247,I379264,I379295,I379312,I379329,I379346,I379363,I379380,I379397,I379414,I379473,I379490,I379507,I379538,I379555,I379586,I379638,I379655,I379672,I379689,I379706,I379737,I379754,I379771,I379788,I379805,I379822,I379839,I379856,I379915,I379932,I379949,I379980,I379997,I380028,I380080,I380097,I380114,I380131,I380148,I380179,I380196,I380213,I380230,I380247,I380264,I380281,I380298,I380357,I380374,I380391,I380422,I380439,I380470,I380522,I380539,I380556,I380573,I380590,I380621,I380638,I380655,I380672,I380689,I380706,I380723,I380740,I380799,I380816,I380833,I380864,I380881,I380912,I380964,I380981,I380998,I381015,I381032,I381063,I381080,I381097,I381114,I381131,I381148,I381165,I381182,I381241,I381258,I381275,I381306,I381323,I381354,I381406,I381423,I381440,I381457,I381474,I381505,I381522,I381539,I381556,I381573,I381590,I381607,I381624,I381683,I381700,I381717,I381748,I381765,I381796,I381848,I381865,I381882,I381899,I381916,I381947,I381964,I381981,I381998,I382015,I382032,I382049,I382066,I382125,I382142,I382159,I382190,I382207,I382238,I382290,I382307,I382324,I382341,I382358,I382389,I382406,I382423,I382440,I382457,I382474,I382491,I382508,I382567,I382584,I382601,I382632,I382649,I382680,I382732,I382749,I382766,I382783,I382800,I382831,I382848,I382865,I382882,I382899,I382916,I382933,I382950,I383009,I383026,I383043,I383074,I383091,I383122,I383174,I383191,I383208,I383225,I383242,I383273,I383290,I383307,I383324,I383341,I383358,I383375,I383392,I383451,I383468,I383485,I383516,I383533,I383564,I383616,I383633,I383650,I383667,I383684,I383715,I383732,I383749,I383766,I383783,I383800,I383817,I383834,I383893,I383910,I383927,I383958,I383975,I384006,I384058,I384075,I384092,I384109,I384126,I384157,I384174,I384191,I384208,I384225,I384242,I384259,I384276,I384335,I384352,I384369,I384400,I384417,I384448,I384500,I384517,I384534,I384551,I384568,I384599,I384616,I384633,I384650,I384667,I384684,I384701,I384718,I384777,I384794,I384811,I384842,I384859,I384890,I384942,I384959,I384976,I384993,I385010,I385041,I385058,I385075,I385092,I385109,I385126,I385143,I385160,I385219,I385236,I385253,I385284,I385301,I385332,I385384,I385401,I385418,I385435,I385452,I385483,I385500,I385517,I385534,I385551,I385568,I385585,I385602,I385661,I385678,I385695,I385726,I385743,I385774,I385826,I385843,I385860,I385877,I385894,I385925,I385942,I385959,I385976,I385993,I386010,I386027,I386044,I386103,I386120,I386137,I386168,I386185,I386216,I386268,I386285,I386302,I386319,I386336,I386367,I386384,I386401,I386418,I386435,I386452,I386469,I386486,I386545,I386562,I386579,I386610,I386627,I386658,I386710,I386727,I386744,I386761,I386778,I386809,I386826,I386843,I386860,I386877,I386894,I386911,I386928,I386987,I387004,I387021,I387052,I387069,I387100,I387152,I387169,I387186,I387203,I387220,I387251,I387268,I387285,I387302,I387319,I387336,I387353,I387370,I387429,I387446,I387463,I387494,I387511,I387542,I387594,I387611,I387628,I387645,I387662,I387693,I387710,I387727,I387744,I387761,I387778,I387795,I387812,I387871,I387888,I387905,I387936,I387953,I387984,I388036,I388053,I388070,I388087,I388104,I388135,I388152,I388169,I388186,I388203,I388220,I388237,I388254,I388313,I388330,I388347,I388378,I388395,I388426,I388478,I388495,I388512,I388529,I388546,I388577,I388594,I388611,I388628,I388645,I388662,I388679,I388696,I388755,I388772,I388789,I388820,I388837,I388868,I388920,I388937,I388954,I388971,I388988,I389019,I389036,I389053,I389070,I389087,I389104,I389121,I389138,I389197,I389214,I389231,I389262,I389279,I389310,I389362,I389379,I389396,I389413,I389430,I389461,I389478,I389495,I389512,I389529,I389546,I389563,I389580,I389639,I389656,I389673,I389704,I389721,I389752,I389804,I389821,I389838,I389855,I389872,I389903,I389920,I389937,I389954,I389971,I389988,I390005,I390022,I390081,I390098,I390115,I390146,I390163,I390194,I390246,I390263,I390280,I390297,I390314,I390345,I390362,I390379,I390396,I390413,I390430,I390447,I390464,I390523,I390540,I390557,I390588,I390605,I390636,I390688,I390705,I390722,I390739,I390756,I390787,I390804,I390821,I390838,I390855,I390872,I390889,I390906,I390965,I390982,I390999,I391030,I391047,I391078,I391130,I391147,I391164,I391181,I391198,I391229,I391246,I391263,I391280,I391297,I391314,I391331,I391348,I391407,I391424,I391441,I391472,I391489,I391520,I391572,I391589,I391606,I391623,I391640,I391671,I391688,I391705,I391722,I391739,I391756,I391773,I391790,I391849,I391866,I391883,I391914,I391931,I391962,I392014,I392031,I392048,I392065,I392082,I392113,I392130,I392147,I392164,I392181,I392198,I392215,I392232,I392291,I392308,I392325,I392356,I392373,I392404,I392456,I392473,I392490,I392507,I392524,I392555,I392572,I392589,I392606,I392623,I392640,I392657,I392674,I392733,I392750,I392767,I392798,I392815,I392846,I392898,I392915,I392932,I392949,I392966,I392997,I393014,I393031,I393048,I393065,I393082,I393099,I393116,I393175,I393192,I393209,I393240,I393257,I393288,I393340,I393357,I393374,I393391,I393408,I393439,I393456,I393473,I393490,I393507,I393524,I393541,I393558,I393617,I393634,I393651,I393682,I393699,I393730,I393782,I393799,I393816,I393833,I393850,I393881,I393898,I393915,I393932,I393949,I393966,I393983,I394000,I394059,I394076,I394093,I394124,I394141,I394172,I394224,I394241,I394258,I394275,I394292,I394323,I394340,I394357,I394374,I394391,I394408,I394425,I394442,I394501,I394518,I394535,I394566,I394583,I394614,I394666,I394683,I394700,I394717,I394734,I394765,I394782,I394799,I394816,I394833,I394850,I394867,I394884,I394943,I394960,I394977,I395008,I395025,I395056,I395108,I395125,I395142,I395159,I395176,I395207,I395224,I395241,I395258,I395275,I395292,I395309,I395326,I395385,I395402,I395419,I395450,I395467,I395498,I395550,I395567,I395584,I395601,I395618,I395649,I395666,I395683,I395700,I395717,I395734,I395751,I395768,I395827,I395844,I395861,I395892,I395909,I395940,I395992,I396009,I396026,I396043,I396060,I396091,I396108,I396125,I396142,I396159,I396176,I396193,I396210,I396269,I396286,I396303,I396334,I396351,I396382,I396434,I396451,I396468,I396485,I396502,I396533,I396550,I396567,I396584,I396601,I396618,I396635,I396652,I396711,I396728,I396745,I396776,I396793,I396824,I396876,I396893,I396910,I396927,I396944,I396975,I396992,I397009,I397026,I397043,I397060,I397077,I397094,I397153,I397170,I397187,I397218,I397235,I397266,I397318,I397335,I397352,I397369,I397386,I397417,I397434,I397451,I397468,I397485,I397502,I397519,I397536,I397595,I397612,I397629,I397660,I397677,I397708,I397760,I397777,I397794,I397811,I397828,I397859,I397876,I397893,I397910,I397927,I397944,I397961,I397978,I398037,I398054,I398071,I398102,I398119,I398150,I398202,I398219,I398236,I398253,I398270,I398301,I398318,I398335,I398352,I398369,I398386,I398403,I398420,I398479,I398496,I398513,I398544,I398561,I398592,I398644,I398661,I398678,I398695,I398712,I398743,I398760,I398777,I398794,I398811,I398828,I398845,I398862,I398921,I398938,I398955,I398986,I399003,I399034,I399086,I399103,I399120,I399137,I399154,I399185,I399202,I399219,I399236,I399253,I399270,I399287,I399304,I399363,I399380,I399397,I399428,I399445,I399476,I399528,I399545,I399562,I399579,I399596,I399627,I399644,I399661,I399678,I399695,I399712,I399729,I399746,I399805,I399822,I399839,I399870,I399887,I399918,I399970,I399987,I400004,I400021,I400038,I400069,I400086,I400103,I400120,I400137,I400154,I400171,I400188,I400247,I400264,I400281,I400312,I400329,I400360,I400412,I400429,I400446,I400463,I400480,I400511,I400528,I400545,I400562,I400579,I400596,I400613,I400630,I400689,I400706,I400723,I400754,I400771,I400802,I400854,I400871,I400888,I400905,I400922,I400953,I400970,I400987,I401004,I401021,I401038,I401055,I401072,I401131,I401148,I401165,I401196,I401213,I401244,I401296,I401313,I401330,I401347,I401364,I401395,I401412,I401429,I401446,I401463,I401480,I401497,I401514,I401573,I401590,I401607,I401638,I401655,I401686,I401738,I401755,I401772,I401789,I401806,I401837,I401854,I401871,I401888,I401905,I401922,I401939,I401956,I402015,I402032,I402049,I402080,I402097,I402128,I402180,I402197,I402214,I402231,I402248,I402279,I402296,I402313,I402330,I402347,I402364,I402381,I402398,I402457,I402474,I402491,I402522,I402539,I402570,I402622,I402639,I402656,I402673,I402690,I402721,I402738,I402755,I402772,I402789,I402806,I402823,I402840,I402899,I402916,I402933,I402964,I402981,I403012,I403064,I403081,I403098,I403115,I403132,I403163,I403180,I403197,I403214,I403231,I403248,I403265,I403282,I403341,I403358,I403375,I403406,I403423,I403454,I403506,I403523,I403540,I403557,I403574,I403605,I403622,I403639,I403656,I403673,I403690,I403707,I403724,I403783,I403800,I403817,I403848,I403865,I403896,I403948,I403965,I403982,I403999,I404016,I404047,I404064,I404081,I404098,I404115,I404132,I404149,I404166,I404225,I404242,I404259,I404290,I404307,I404338,I404390,I404407,I404424,I404441,I404458,I404489,I404506,I404523,I404540,I404557,I404574,I404591,I404608,I404667,I404684,I404701,I404732,I404749,I404780,I404832,I404849,I404866,I404883,I404900,I404931,I404948,I404965,I404982,I404999,I405016,I405033,I405050,I405109,I405126,I405143,I405174,I405191,I405222,I405274,I405291,I405308,I405325,I405342,I405373,I405390,I405407,I405424,I405441,I405458,I405475,I405492,I405551,I405568,I405585,I405616,I405633,I405664,I405716,I405733,I405750,I405767,I405784,I405815,I405832,I405849,I405866,I405883,I405900,I405917,I405934,I405993,I406010,I406027,I406058,I406075,I406106,I406158,I406175,I406192,I406209,I406226,I406257,I406274,I406291,I406308,I406325,I406342,I406359,I406376,I406435,I406452,I406469,I406500,I406517,I406548,I406600,I406617,I406634,I406651,I406668,I406699,I406716,I406733,I406750,I406767,I406784,I406801,I406818,I406877,I406894,I406911,I406942,I406959,I406990,I407042,I407059,I407076,I407093,I407110,I407141,I407158,I407175,I407192,I407209,I407226,I407243,I407260,I407319,I407336,I407353,I407384,I407401,I407432,I407484,I407501,I407518,I407535,I407552,I407583,I407600,I407617,I407634,I407651,I407668,I407685,I407702,I407761,I407778,I407795,I407826,I407843,I407874,I407926,I407943,I407960,I407977,I407994,I408025,I408042,I408059,I408076,I408093,I408110,I408127,I408144,I408203,I408220,I408237,I408268,I408285,I408316,I408368,I408385,I408402,I408419,I408436,I408467,I408484,I408501,I408518,I408535,I408552,I408569,I408586,I408645,I408662,I408679,I408710,I408727,I408758,I408810,I408827,I408844,I408861,I408878,I408909,I408926,I408943,I408960,I408977,I408994,I409011,I409028,I409087,I409104,I409121,I409152,I409169,I409200,I409252,I409269,I409286,I409303,I409320,I409351,I409368,I409385,I409402,I409419,I409436,I409453,I409470,I409529,I409546,I409563,I409594,I409611,I409642,I409694,I409711,I409728,I409745,I409762,I409793,I409810,I409827,I409844,I409861,I409878,I409895,I409912,I409971,I409988,I410005,I410036,I410053,I410084,I410136,I410153,I410170,I410187,I410204,I410235,I410252,I410269,I410286,I410303,I410320,I410337,I410354,I410413,I410430,I410447,I410478,I410495,I410526,I410578,I410595,I410612,I410629,I410646,I410677,I410694,I410711,I410728,I410745,I410762,I410779,I410796,I410855,I410872,I410889,I410920,I410937,I410968;
not I_0 (I1901,I1869);
or I_1 (I1918,I145780,I145798);
nand I_2 (I1935,I145783,I145777);
not I_3 (I1952,I1935);
and I_4 (I1969,I1952,I1918);
DFFARX1 I_5 (I1952,I1862,I1901,I1881,);
nand I_6 (I2000,I145777,I145801);
and I_7 (I2017,I2000,I145792);
DFFARX1 I_8 (I2017,I1862,I1901,I2043,);
nor I_9 (I2051,I2043,I1969);
not I_10 (I2068,I2043);
nor I_11 (I2085,I145780,I145801);
not I_12 (I2102,I2085);
nand I_13 (I2119,I2068,I2102);
nand I_14 (I2136,I2085,I1935);
nand I_15 (I2153,I2068,I2136);
nand I_16 (I1887,I2051,I2085);
not I_17 (I2184,I145786);
nand I_18 (I2201,I2119,I2184);
nand I_19 (I2218,I145795,I145789);
nor I_20 (I1872,I1969,I2218);
not I_21 (I2249,I2218);
nand I_22 (I2266,I2249,I2184);
nor I_23 (I2283,I2102,I2266);
nor I_24 (I1890,I2068,I2283);
nor I_25 (I1893,I2218,I2201);
nor I_26 (I2328,I2218,I145786);
nor I_27 (I1875,I2328,I2153);
nand I_28 (I1878,I1952,I2218);
nor I_29 (I2373,I2043,I2218);
nand I_30 (I1884,I2373,I1969);
not I_31 (I2428,I1869);
or I_32 (I2445,I1503,I999);
nand I_33 (I2462,I1151,I1415);
not I_34 (I2479,I2462);
and I_35 (I2496,I2479,I2445);
DFFARX1 I_36 (I2479,I1862,I2428,I2408,);
nand I_37 (I2527,I1679,I1727);
and I_38 (I2544,I2527,I1687);
DFFARX1 I_39 (I2544,I1862,I2428,I2570,);
nor I_40 (I2578,I2570,I2496);
not I_41 (I2595,I2570);
nor I_42 (I2612,I1263,I1727);
not I_43 (I2629,I2612);
nand I_44 (I2646,I2595,I2629);
nand I_45 (I2663,I2612,I2462);
nand I_46 (I2680,I2595,I2663);
nand I_47 (I2414,I2578,I2612);
not I_48 (I2711,I1231);
nand I_49 (I2728,I2646,I2711);
nand I_50 (I2745,I1767,I1343);
nor I_51 (I2399,I2496,I2745);
not I_52 (I2776,I2745);
nand I_53 (I2793,I2776,I2711);
nor I_54 (I2810,I2629,I2793);
nor I_55 (I2417,I2595,I2810);
nor I_56 (I2420,I2745,I2728);
nor I_57 (I2855,I2745,I1231);
nor I_58 (I2402,I2855,I2680);
nand I_59 (I2405,I2479,I2745);
nor I_60 (I2900,I2570,I2745);
nand I_61 (I2411,I2900,I2496);
not I_62 (I2955,I1869);
or I_63 (I2972,I337869,I337881);
nand I_64 (I2989,I337860,I337863);
not I_65 (I3006,I2989);
and I_66 (I3023,I3006,I2972);
DFFARX1 I_67 (I3006,I1862,I2955,I2935,);
nand I_68 (I3054,I337860,I337872);
and I_69 (I3071,I3054,I337875);
DFFARX1 I_70 (I3071,I1862,I2955,I3097,);
nor I_71 (I3105,I3097,I3023);
not I_72 (I3122,I3097);
nor I_73 (I3139,I337866,I337872);
not I_74 (I3156,I3139);
nand I_75 (I3173,I3122,I3156);
nand I_76 (I3190,I3139,I2989);
nand I_77 (I3207,I3122,I3190);
nand I_78 (I2941,I3105,I3139);
not I_79 (I3238,I337866);
nand I_80 (I3255,I3173,I3238);
nand I_81 (I3272,I337863,I337878);
nor I_82 (I2926,I3023,I3272);
not I_83 (I3303,I3272);
nand I_84 (I3320,I3303,I3238);
nor I_85 (I3337,I3156,I3320);
nor I_86 (I2944,I3122,I3337);
nor I_87 (I2947,I3272,I3255);
nor I_88 (I3382,I3272,I337866);
nor I_89 (I2929,I3382,I3207);
nand I_90 (I2932,I3006,I3272);
nor I_91 (I3427,I3097,I3272);
nand I_92 (I2938,I3427,I3023);
not I_93 (I3482,I1869);
or I_94 (I3499,I363712,I363706);
nand I_95 (I3516,I363703,I363703);
not I_96 (I3533,I3516);
and I_97 (I3550,I3533,I3499);
DFFARX1 I_98 (I3533,I1862,I3482,I3462,);
nand I_99 (I3581,I363709,I363715);
and I_100 (I3598,I3581,I363709);
DFFARX1 I_101 (I3598,I1862,I3482,I3624,);
nor I_102 (I3632,I3624,I3550);
not I_103 (I3649,I3624);
nor I_104 (I3666,I363700,I363715);
not I_105 (I3683,I3666);
nand I_106 (I3700,I3649,I3683);
nand I_107 (I3717,I3666,I3516);
nand I_108 (I3734,I3649,I3717);
nand I_109 (I3468,I3632,I3666);
not I_110 (I3765,I363700);
nand I_111 (I3782,I3700,I3765);
nand I_112 (I3799,I363718,I363706);
nor I_113 (I3453,I3550,I3799);
not I_114 (I3830,I3799);
nand I_115 (I3847,I3830,I3765);
nor I_116 (I3864,I3683,I3847);
nor I_117 (I3471,I3649,I3864);
nor I_118 (I3474,I3799,I3782);
nor I_119 (I3909,I3799,I363700);
nor I_120 (I3456,I3909,I3734);
nand I_121 (I3459,I3533,I3799);
nor I_122 (I3954,I3624,I3799);
nand I_123 (I3465,I3954,I3550);
not I_124 (I4009,I1869);
or I_125 (I4026,I18586,I18586);
nand I_126 (I4043,I18607,I18604);
not I_127 (I4060,I4043);
and I_128 (I4077,I4060,I4026);
DFFARX1 I_129 (I4060,I1862,I4009,I3989,);
nand I_130 (I4108,I18583,I18595);
and I_131 (I4125,I4108,I18592);
DFFARX1 I_132 (I4125,I1862,I4009,I4151,);
nor I_133 (I4159,I4151,I4077);
not I_134 (I4176,I4151);
nor I_135 (I4193,I18601,I18595);
not I_136 (I4210,I4193);
nand I_137 (I4227,I4176,I4210);
nand I_138 (I4244,I4193,I4043);
nand I_139 (I4261,I4176,I4244);
nand I_140 (I3995,I4159,I4193);
not I_141 (I4292,I18583);
nand I_142 (I4309,I4227,I4292);
nand I_143 (I4326,I18598,I18589);
nor I_144 (I3980,I4077,I4326);
not I_145 (I4357,I4326);
nand I_146 (I4374,I4357,I4292);
nor I_147 (I4391,I4210,I4374);
nor I_148 (I3998,I4176,I4391);
nor I_149 (I4001,I4326,I4309);
nor I_150 (I4436,I4326,I18583);
nor I_151 (I3983,I4436,I4261);
nand I_152 (I3986,I4060,I4326);
nor I_153 (I4481,I4151,I4326);
nand I_154 (I3992,I4481,I4077);
not I_155 (I4536,I1869);
or I_156 (I4553,I384044,I384038);
nand I_157 (I4570,I384035,I384035);
not I_158 (I4587,I4570);
and I_159 (I4604,I4587,I4553);
DFFARX1 I_160 (I4587,I1862,I4536,I4516,);
nand I_161 (I4635,I384041,I384047);
and I_162 (I4652,I4635,I384041);
DFFARX1 I_163 (I4652,I1862,I4536,I4678,);
nor I_164 (I4686,I4678,I4604);
not I_165 (I4703,I4678);
nor I_166 (I4720,I384032,I384047);
not I_167 (I4737,I4720);
nand I_168 (I4754,I4703,I4737);
nand I_169 (I4771,I4720,I4570);
nand I_170 (I4788,I4703,I4771);
nand I_171 (I4522,I4686,I4720);
not I_172 (I4819,I384032);
nand I_173 (I4836,I4754,I4819);
nand I_174 (I4853,I384050,I384038);
nor I_175 (I4507,I4604,I4853);
not I_176 (I4884,I4853);
nand I_177 (I4901,I4884,I4819);
nor I_178 (I4918,I4737,I4901);
nor I_179 (I4525,I4703,I4918);
nor I_180 (I4528,I4853,I4836);
nor I_181 (I4963,I4853,I384032);
nor I_182 (I4510,I4963,I4788);
nand I_183 (I4513,I4587,I4853);
nor I_184 (I5008,I4678,I4853);
nand I_185 (I4519,I5008,I4604);
not I_186 (I5063,I1869);
or I_187 (I5080,I355787,I355799);
nand I_188 (I5097,I355778,I355781);
not I_189 (I5114,I5097);
and I_190 (I5131,I5114,I5080);
DFFARX1 I_191 (I5114,I1862,I5063,I5043,);
nand I_192 (I5162,I355778,I355790);
and I_193 (I5179,I5162,I355793);
DFFARX1 I_194 (I5179,I1862,I5063,I5205,);
nor I_195 (I5213,I5205,I5131);
not I_196 (I5230,I5205);
nor I_197 (I5247,I355784,I355790);
not I_198 (I5264,I5247);
nand I_199 (I5281,I5230,I5264);
nand I_200 (I5298,I5247,I5097);
nand I_201 (I5315,I5230,I5298);
nand I_202 (I5049,I5213,I5247);
not I_203 (I5346,I355784);
nand I_204 (I5363,I5281,I5346);
nand I_205 (I5380,I355781,I355796);
nor I_206 (I5034,I5131,I5380);
not I_207 (I5411,I5380);
nand I_208 (I5428,I5411,I5346);
nor I_209 (I5445,I5264,I5428);
nor I_210 (I5052,I5230,I5445);
nor I_211 (I5055,I5380,I5363);
nor I_212 (I5490,I5380,I355784);
nor I_213 (I5037,I5490,I5315);
nand I_214 (I5040,I5114,I5380);
nor I_215 (I5535,I5205,I5380);
nand I_216 (I5046,I5535,I5131);
not I_217 (I5590,I1869);
or I_218 (I5607,I272479,I272461);
nand I_219 (I5624,I272467,I272482);
not I_220 (I5641,I5624);
and I_221 (I5658,I5641,I5607);
DFFARX1 I_222 (I5641,I1862,I5590,I5570,);
nand I_223 (I5689,I272464,I272470);
and I_224 (I5706,I5689,I272467);
DFFARX1 I_225 (I5706,I1862,I5590,I5732,);
nor I_226 (I5740,I5732,I5658);
not I_227 (I5757,I5732);
nor I_228 (I5774,I272473,I272470);
not I_229 (I5791,I5774);
nand I_230 (I5808,I5757,I5791);
nand I_231 (I5825,I5774,I5624);
nand I_232 (I5842,I5757,I5825);
nand I_233 (I5576,I5740,I5774);
not I_234 (I5873,I272464);
nand I_235 (I5890,I5808,I5873);
nand I_236 (I5907,I272476,I272461);
nor I_237 (I5561,I5658,I5907);
not I_238 (I5938,I5907);
nand I_239 (I5955,I5938,I5873);
nor I_240 (I5972,I5791,I5955);
nor I_241 (I5579,I5757,I5972);
nor I_242 (I5582,I5907,I5890);
nor I_243 (I6017,I5907,I272464);
nor I_244 (I5564,I6017,I5842);
nand I_245 (I5567,I5641,I5907);
nor I_246 (I6062,I5732,I5907);
nand I_247 (I5573,I6062,I5658);
not I_248 (I6117,I1869);
or I_249 (I6134,I184251,I184269);
nand I_250 (I6151,I184254,I184248);
not I_251 (I6168,I6151);
and I_252 (I6185,I6168,I6134);
DFFARX1 I_253 (I6168,I1862,I6117,I6097,);
nand I_254 (I6216,I184248,I184272);
and I_255 (I6233,I6216,I184263);
DFFARX1 I_256 (I6233,I1862,I6117,I6259,);
nor I_257 (I6267,I6259,I6185);
not I_258 (I6284,I6259);
nor I_259 (I6301,I184251,I184272);
not I_260 (I6318,I6301);
nand I_261 (I6335,I6284,I6318);
nand I_262 (I6352,I6301,I6151);
nand I_263 (I6369,I6284,I6352);
nand I_264 (I6103,I6267,I6301);
not I_265 (I6400,I184257);
nand I_266 (I6417,I6335,I6400);
nand I_267 (I6434,I184266,I184260);
nor I_268 (I6088,I6185,I6434);
not I_269 (I6465,I6434);
nand I_270 (I6482,I6465,I6400);
nor I_271 (I6499,I6318,I6482);
nor I_272 (I6106,I6284,I6499);
nor I_273 (I6109,I6434,I6417);
nor I_274 (I6544,I6434,I184257);
nor I_275 (I6091,I6544,I6369);
nand I_276 (I6094,I6168,I6434);
nor I_277 (I6589,I6259,I6434);
nand I_278 (I6100,I6589,I6185);
not I_279 (I6644,I1869);
or I_280 (I6661,I64486,I64486);
nand I_281 (I6678,I64507,I64504);
not I_282 (I6695,I6678);
and I_283 (I6712,I6695,I6661);
DFFARX1 I_284 (I6695,I1862,I6644,I6624,);
nand I_285 (I6743,I64483,I64495);
and I_286 (I6760,I6743,I64492);
DFFARX1 I_287 (I6760,I1862,I6644,I6786,);
nor I_288 (I6794,I6786,I6712);
not I_289 (I6811,I6786);
nor I_290 (I6828,I64501,I64495);
not I_291 (I6845,I6828);
nand I_292 (I6862,I6811,I6845);
nand I_293 (I6879,I6828,I6678);
nand I_294 (I6896,I6811,I6879);
nand I_295 (I6630,I6794,I6828);
not I_296 (I6927,I64483);
nand I_297 (I6944,I6862,I6927);
nand I_298 (I6961,I64498,I64489);
nor I_299 (I6615,I6712,I6961);
not I_300 (I6992,I6961);
nand I_301 (I7009,I6992,I6927);
nor I_302 (I7026,I6845,I7009);
nor I_303 (I6633,I6811,I7026);
nor I_304 (I6636,I6961,I6944);
nor I_305 (I7071,I6961,I64483);
nor I_306 (I6618,I7071,I6896);
nand I_307 (I6621,I6695,I6961);
nor I_308 (I7116,I6786,I6961);
nand I_309 (I6627,I7116,I6712);
not I_310 (I7171,I1869);
or I_311 (I7188,I175819,I175837);
nand I_312 (I7205,I175822,I175816);
not I_313 (I7222,I7205);
and I_314 (I7239,I7222,I7188);
DFFARX1 I_315 (I7222,I1862,I7171,I7151,);
nand I_316 (I7270,I175816,I175840);
and I_317 (I7287,I7270,I175831);
DFFARX1 I_318 (I7287,I1862,I7171,I7313,);
nor I_319 (I7321,I7313,I7239);
not I_320 (I7338,I7313);
nor I_321 (I7355,I175819,I175840);
not I_322 (I7372,I7355);
nand I_323 (I7389,I7338,I7372);
nand I_324 (I7406,I7355,I7205);
nand I_325 (I7423,I7338,I7406);
nand I_326 (I7157,I7321,I7355);
not I_327 (I7454,I175825);
nand I_328 (I7471,I7389,I7454);
nand I_329 (I7488,I175834,I175828);
nor I_330 (I7142,I7239,I7488);
not I_331 (I7519,I7488);
nand I_332 (I7536,I7519,I7454);
nor I_333 (I7553,I7372,I7536);
nor I_334 (I7160,I7338,I7553);
nor I_335 (I7163,I7488,I7471);
nor I_336 (I7598,I7488,I175825);
nor I_337 (I7145,I7598,I7423);
nand I_338 (I7148,I7222,I7488);
nor I_339 (I7643,I7313,I7488);
nand I_340 (I7154,I7643,I7239);
not I_341 (I7698,I1869);
or I_342 (I7715,I38476,I38476);
nand I_343 (I7732,I38497,I38494);
not I_344 (I7749,I7732);
and I_345 (I7766,I7749,I7715);
DFFARX1 I_346 (I7749,I1862,I7698,I7678,);
nand I_347 (I7797,I38473,I38485);
and I_348 (I7814,I7797,I38482);
DFFARX1 I_349 (I7814,I1862,I7698,I7840,);
nor I_350 (I7848,I7840,I7766);
not I_351 (I7865,I7840);
nor I_352 (I7882,I38491,I38485);
not I_353 (I7899,I7882);
nand I_354 (I7916,I7865,I7899);
nand I_355 (I7933,I7882,I7732);
nand I_356 (I7950,I7865,I7933);
nand I_357 (I7684,I7848,I7882);
not I_358 (I7981,I38473);
nand I_359 (I7998,I7916,I7981);
nand I_360 (I8015,I38488,I38479);
nor I_361 (I7669,I7766,I8015);
not I_362 (I8046,I8015);
nand I_363 (I8063,I8046,I7981);
nor I_364 (I8080,I7899,I8063);
nor I_365 (I7687,I7865,I8080);
nor I_366 (I7690,I8015,I7998);
nor I_367 (I8125,I8015,I38473);
nor I_368 (I7672,I8125,I7950);
nand I_369 (I7675,I7749,I8015);
nor I_370 (I8170,I7840,I8015);
nand I_371 (I7681,I8170,I7766);
not I_372 (I8225,I1869);
or I_373 (I8242,I169495,I169513);
nand I_374 (I8259,I169498,I169492);
not I_375 (I8276,I8259);
and I_376 (I8293,I8276,I8242);
DFFARX1 I_377 (I8276,I1862,I8225,I8205,);
nand I_378 (I8324,I169492,I169516);
and I_379 (I8341,I8324,I169507);
DFFARX1 I_380 (I8341,I1862,I8225,I8367,);
nor I_381 (I8375,I8367,I8293);
not I_382 (I8392,I8367);
nor I_383 (I8409,I169495,I169516);
not I_384 (I8426,I8409);
nand I_385 (I8443,I8392,I8426);
nand I_386 (I8460,I8409,I8259);
nand I_387 (I8477,I8392,I8460);
nand I_388 (I8211,I8375,I8409);
not I_389 (I8508,I169501);
nand I_390 (I8525,I8443,I8508);
nand I_391 (I8542,I169510,I169504);
nor I_392 (I8196,I8293,I8542);
not I_393 (I8573,I8542);
nand I_394 (I8590,I8573,I8508);
nor I_395 (I8607,I8426,I8590);
nor I_396 (I8214,I8392,I8607);
nor I_397 (I8217,I8542,I8525);
nor I_398 (I8652,I8542,I169501);
nor I_399 (I8199,I8652,I8477);
nand I_400 (I8202,I8276,I8542);
nor I_401 (I8697,I8367,I8542);
nand I_402 (I8208,I8697,I8293);
not I_403 (I8752,I1869);
or I_404 (I8769,I219643,I219625);
nand I_405 (I8786,I219631,I219646);
not I_406 (I8803,I8786);
and I_407 (I8820,I8803,I8769);
DFFARX1 I_408 (I8803,I1862,I8752,I8732,);
nand I_409 (I8851,I219628,I219634);
and I_410 (I8868,I8851,I219631);
DFFARX1 I_411 (I8868,I1862,I8752,I8894,);
nor I_412 (I8902,I8894,I8820);
not I_413 (I8919,I8894);
nor I_414 (I8936,I219637,I219634);
not I_415 (I8953,I8936);
nand I_416 (I8970,I8919,I8953);
nand I_417 (I8987,I8936,I8786);
nand I_418 (I9004,I8919,I8987);
nand I_419 (I8738,I8902,I8936);
not I_420 (I9035,I219628);
nand I_421 (I9052,I8970,I9035);
nand I_422 (I9069,I219640,I219625);
nor I_423 (I8723,I8820,I9069);
not I_424 (I9100,I9069);
nand I_425 (I9117,I9100,I9035);
nor I_426 (I9134,I8953,I9117);
nor I_427 (I8741,I8919,I9134);
nor I_428 (I8744,I9069,I9052);
nor I_429 (I9179,I9069,I219628);
nor I_430 (I8726,I9179,I9004);
nand I_431 (I8729,I8803,I9069);
nor I_432 (I9224,I8894,I9069);
nand I_433 (I8735,I9224,I8820);
not I_434 (I9279,I1869);
or I_435 (I9296,I134186,I134204);
nand I_436 (I9313,I134189,I134183);
not I_437 (I9330,I9313);
and I_438 (I9347,I9330,I9296);
DFFARX1 I_439 (I9330,I1862,I9279,I9259,);
nand I_440 (I9378,I134183,I134207);
and I_441 (I9395,I9378,I134198);
DFFARX1 I_442 (I9395,I1862,I9279,I9421,);
nor I_443 (I9429,I9421,I9347);
not I_444 (I9446,I9421);
nor I_445 (I9463,I134186,I134207);
not I_446 (I9480,I9463);
nand I_447 (I9497,I9446,I9480);
nand I_448 (I9514,I9463,I9313);
nand I_449 (I9531,I9446,I9514);
nand I_450 (I9265,I9429,I9463);
not I_451 (I9562,I134192);
nand I_452 (I9579,I9497,I9562);
nand I_453 (I9596,I134201,I134195);
nor I_454 (I9250,I9347,I9596);
not I_455 (I9627,I9596);
nand I_456 (I9644,I9627,I9562);
nor I_457 (I9661,I9480,I9644);
nor I_458 (I9268,I9446,I9661);
nor I_459 (I9271,I9596,I9579);
nor I_460 (I9706,I9596,I134192);
nor I_461 (I9253,I9706,I9531);
nand I_462 (I9256,I9330,I9596);
nor I_463 (I9751,I9421,I9596);
nand I_464 (I9262,I9751,I9347);
not I_465 (I9806,I1869);
or I_466 (I9823,I291490,I291484);
nand I_467 (I9840,I291499,I291502);
not I_468 (I9857,I9840);
and I_469 (I9874,I9857,I9823);
DFFARX1 I_470 (I9857,I1862,I9806,I9786,);
nand I_471 (I9905,I291484,I291487);
and I_472 (I9922,I9905,I291490);
DFFARX1 I_473 (I9922,I1862,I9806,I9948,);
nor I_474 (I9956,I9948,I9874);
not I_475 (I9973,I9948);
nor I_476 (I9990,I291505,I291487);
not I_477 (I10007,I9990);
nand I_478 (I10024,I9973,I10007);
nand I_479 (I10041,I9990,I9840);
nand I_480 (I10058,I9973,I10041);
nand I_481 (I9792,I9956,I9990);
not I_482 (I10089,I291487);
nand I_483 (I10106,I10024,I10089);
nand I_484 (I10123,I291496,I291493);
nor I_485 (I9777,I9874,I10123);
not I_486 (I10154,I10123);
nand I_487 (I10171,I10154,I10089);
nor I_488 (I10188,I10007,I10171);
nor I_489 (I9795,I9973,I10188);
nor I_490 (I9798,I10123,I10106);
nor I_491 (I10233,I10123,I291487);
nor I_492 (I9780,I10233,I10058);
nand I_493 (I9783,I9857,I10123);
nor I_494 (I10278,I9948,I10123);
nand I_495 (I9789,I10278,I9874);
not I_496 (I10333,I1869);
or I_497 (I10350,I246299,I246281);
nand I_498 (I10367,I246287,I246302);
not I_499 (I10384,I10367);
and I_500 (I10401,I10384,I10350);
DFFARX1 I_501 (I10384,I1862,I10333,I10313,);
nand I_502 (I10432,I246284,I246290);
and I_503 (I10449,I10432,I246287);
DFFARX1 I_504 (I10449,I1862,I10333,I10475,);
nor I_505 (I10483,I10475,I10401);
not I_506 (I10500,I10475);
nor I_507 (I10517,I246293,I246290);
not I_508 (I10534,I10517);
nand I_509 (I10551,I10500,I10534);
nand I_510 (I10568,I10517,I10367);
nand I_511 (I10585,I10500,I10568);
nand I_512 (I10319,I10483,I10517);
not I_513 (I10616,I246284);
nand I_514 (I10633,I10551,I10616);
nand I_515 (I10650,I246296,I246281);
nor I_516 (I10304,I10401,I10650);
not I_517 (I10681,I10650);
nand I_518 (I10698,I10681,I10616);
nor I_519 (I10715,I10534,I10698);
nor I_520 (I10322,I10500,I10715);
nor I_521 (I10325,I10650,I10633);
nor I_522 (I10760,I10650,I246284);
nor I_523 (I10307,I10760,I10585);
nand I_524 (I10310,I10384,I10650);
nor I_525 (I10805,I10475,I10650);
nand I_526 (I10316,I10805,I10401);
not I_527 (I10860,I1869);
or I_528 (I10877,I332599,I332611);
nand I_529 (I10894,I332590,I332593);
not I_530 (I10911,I10894);
and I_531 (I10928,I10911,I10877);
DFFARX1 I_532 (I10911,I1862,I10860,I10840,);
nand I_533 (I10959,I332590,I332602);
and I_534 (I10976,I10959,I332605);
DFFARX1 I_535 (I10976,I1862,I10860,I11002,);
nor I_536 (I11010,I11002,I10928);
not I_537 (I11027,I11002);
nor I_538 (I11044,I332596,I332602);
not I_539 (I11061,I11044);
nand I_540 (I11078,I11027,I11061);
nand I_541 (I11095,I11044,I10894);
nand I_542 (I11112,I11027,I11095);
nand I_543 (I10846,I11010,I11044);
not I_544 (I11143,I332596);
nand I_545 (I11160,I11078,I11143);
nand I_546 (I11177,I332593,I332608);
nor I_547 (I10831,I10928,I11177);
not I_548 (I11208,I11177);
nand I_549 (I11225,I11208,I11143);
nor I_550 (I11242,I11061,I11225);
nor I_551 (I10849,I11027,I11242);
nor I_552 (I10852,I11177,I11160);
nor I_553 (I11287,I11177,I332596);
nor I_554 (I10834,I11287,I11112);
nand I_555 (I10837,I10911,I11177);
nor I_556 (I11332,I11002,I11177);
nand I_557 (I10843,I11332,I10928);
not I_558 (I11387,I1869);
or I_559 (I11404,I71626,I71626);
nand I_560 (I11421,I71647,I71644);
not I_561 (I11438,I11421);
and I_562 (I11455,I11438,I11404);
DFFARX1 I_563 (I11438,I1862,I11387,I11367,);
nand I_564 (I11486,I71623,I71635);
and I_565 (I11503,I11486,I71632);
DFFARX1 I_566 (I11503,I1862,I11387,I11529,);
nor I_567 (I11537,I11529,I11455);
not I_568 (I11554,I11529);
nor I_569 (I11571,I71641,I71635);
not I_570 (I11588,I11571);
nand I_571 (I11605,I11554,I11588);
nand I_572 (I11622,I11571,I11421);
nand I_573 (I11639,I11554,I11622);
nand I_574 (I11373,I11537,I11571);
not I_575 (I11670,I71623);
nand I_576 (I11687,I11605,I11670);
nand I_577 (I11704,I71638,I71629);
nor I_578 (I11358,I11455,I11704);
not I_579 (I11735,I11704);
nand I_580 (I11752,I11735,I11670);
nor I_581 (I11769,I11588,I11752);
nor I_582 (I11376,I11554,I11769);
nor I_583 (I11379,I11704,I11687);
nor I_584 (I11814,I11704,I71623);
nor I_585 (I11361,I11814,I11639);
nand I_586 (I11364,I11438,I11704);
nor I_587 (I11859,I11529,I11704);
nand I_588 (I11370,I11859,I11455);
not I_589 (I11914,I1869);
or I_590 (I11931,I121011,I121029);
nand I_591 (I11948,I121014,I121008);
not I_592 (I11965,I11948);
and I_593 (I11982,I11965,I11931);
DFFARX1 I_594 (I11965,I1862,I11914,I11894,);
nand I_595 (I12013,I121008,I121032);
and I_596 (I12030,I12013,I121023);
DFFARX1 I_597 (I12030,I1862,I11914,I12056,);
nor I_598 (I12064,I12056,I11982);
not I_599 (I12081,I12056);
nor I_600 (I12098,I121011,I121032);
not I_601 (I12115,I12098);
nand I_602 (I12132,I12081,I12115);
nand I_603 (I12149,I12098,I11948);
nand I_604 (I12166,I12081,I12149);
nand I_605 (I11900,I12064,I12098);
not I_606 (I12197,I121017);
nand I_607 (I12214,I12132,I12197);
nand I_608 (I12231,I121026,I121020);
nor I_609 (I11885,I11982,I12231);
not I_610 (I12262,I12231);
nand I_611 (I12279,I12262,I12197);
nor I_612 (I12296,I12115,I12279);
nor I_613 (I11903,I12081,I12296);
nor I_614 (I11906,I12231,I12214);
nor I_615 (I12341,I12231,I121017);
nor I_616 (I11888,I12341,I12166);
nand I_617 (I11891,I11965,I12231);
nor I_618 (I12386,I12056,I12231);
nand I_619 (I11897,I12386,I11982);
not I_620 (I12441,I1869);
or I_621 (I12458,I142618,I142636);
nand I_622 (I12475,I142621,I142615);
not I_623 (I12492,I12475);
and I_624 (I12509,I12492,I12458);
DFFARX1 I_625 (I12492,I1862,I12441,I12421,);
nand I_626 (I12540,I142615,I142639);
and I_627 (I12557,I12540,I142630);
DFFARX1 I_628 (I12557,I1862,I12441,I12583,);
nor I_629 (I12591,I12583,I12509);
not I_630 (I12608,I12583);
nor I_631 (I12625,I142618,I142639);
not I_632 (I12642,I12625);
nand I_633 (I12659,I12608,I12642);
nand I_634 (I12676,I12625,I12475);
nand I_635 (I12693,I12608,I12676);
nand I_636 (I12427,I12591,I12625);
not I_637 (I12724,I142624);
nand I_638 (I12741,I12659,I12724);
nand I_639 (I12758,I142633,I142627);
nor I_640 (I12412,I12509,I12758);
not I_641 (I12789,I12758);
nand I_642 (I12806,I12789,I12724);
nor I_643 (I12823,I12642,I12806);
nor I_644 (I12430,I12608,I12823);
nor I_645 (I12433,I12758,I12741);
nor I_646 (I12868,I12758,I142624);
nor I_647 (I12415,I12868,I12693);
nand I_648 (I12418,I12492,I12758);
nor I_649 (I12913,I12583,I12758);
nand I_650 (I12424,I12913,I12509);
not I_651 (I12968,I1869);
or I_652 (I12985,I129443,I129461);
nand I_653 (I13002,I129446,I129440);
not I_654 (I13019,I13002);
and I_655 (I13036,I13019,I12985);
DFFARX1 I_656 (I13019,I1862,I12968,I12948,);
nand I_657 (I13067,I129440,I129464);
and I_658 (I13084,I13067,I129455);
DFFARX1 I_659 (I13084,I1862,I12968,I13110,);
nor I_660 (I13118,I13110,I13036);
not I_661 (I13135,I13110);
nor I_662 (I13152,I129443,I129464);
not I_663 (I13169,I13152);
nand I_664 (I13186,I13135,I13169);
nand I_665 (I13203,I13152,I13002);
nand I_666 (I13220,I13135,I13203);
nand I_667 (I12954,I13118,I13152);
not I_668 (I13251,I129449);
nand I_669 (I13268,I13186,I13251);
nand I_670 (I13285,I129458,I129452);
nor I_671 (I12939,I13036,I13285);
not I_672 (I13316,I13285);
nand I_673 (I13333,I13316,I13251);
nor I_674 (I13350,I13169,I13333);
nor I_675 (I12957,I13135,I13350);
nor I_676 (I12960,I13285,I13268);
nor I_677 (I13395,I13285,I129449);
nor I_678 (I12942,I13395,I13220);
nand I_679 (I12945,I13019,I13285);
nor I_680 (I13440,I13110,I13285);
nand I_681 (I12951,I13440,I13036);
not I_682 (I13495,I1869);
or I_683 (I13512,I39496,I39496);
nand I_684 (I13529,I39517,I39514);
not I_685 (I13546,I13529);
and I_686 (I13563,I13546,I13512);
DFFARX1 I_687 (I13546,I1862,I13495,I13475,);
nand I_688 (I13594,I39493,I39505);
and I_689 (I13611,I13594,I39502);
DFFARX1 I_690 (I13611,I1862,I13495,I13637,);
nor I_691 (I13645,I13637,I13563);
not I_692 (I13662,I13637);
nor I_693 (I13679,I39511,I39505);
not I_694 (I13696,I13679);
nand I_695 (I13713,I13662,I13696);
nand I_696 (I13730,I13679,I13529);
nand I_697 (I13747,I13662,I13730);
nand I_698 (I13481,I13645,I13679);
not I_699 (I13778,I39493);
nand I_700 (I13795,I13713,I13778);
nand I_701 (I13812,I39508,I39499);
nor I_702 (I13466,I13563,I13812);
not I_703 (I13843,I13812);
nand I_704 (I13860,I13843,I13778);
nor I_705 (I13877,I13696,I13860);
nor I_706 (I13484,I13662,I13877);
nor I_707 (I13487,I13812,I13795);
nor I_708 (I13922,I13812,I39493);
nor I_709 (I13469,I13922,I13747);
nand I_710 (I13472,I13546,I13812);
nor I_711 (I13967,I13637,I13812);
nand I_712 (I13478,I13967,I13563);
not I_713 (I14025,I1869);
or I_714 (I14042,I202492,I202495);
nand I_715 (I14059,I202501,I202489);
not I_716 (I14076,I14059);
nand I_717 (I14093,I14076,I14042);
not I_718 (I14110,I14093);
nand I_719 (I14127,I202507,I202510);
and I_720 (I14144,I14127,I202504);
DFFARX1 I_721 (I14144,I1862,I14025,I14170,);
not I_722 (I14178,I14170);
nor I_723 (I14195,I202492,I202510);
nor I_724 (I14212,I14170,I14195);
and I_725 (I14229,I14170,I14195);
nor I_726 (I14246,I14229,I14093);
DFFARX1 I_727 (I14246,I1862,I14025,I14005,);
nand I_728 (I14277,I202495,I202498);
nor I_729 (I14294,I14277,I202489);
nand I_730 (I14311,I14110,I14294);
not I_731 (I14014,I14311);
nor I_732 (I14017,I14212,I14311);
nor I_733 (I14356,I14294,I14076);
nor I_734 (I14008,I14178,I14356);
nor I_735 (I14002,I14294,I14195);
not I_736 (I14401,I14277);
nand I_737 (I14418,I14195,I14401);
not I_738 (I13996,I14418);
nor I_739 (I13999,I14059,I14418);
nor I_740 (I14011,I14401,I14059);
nand I_741 (I14477,I14178,I14277);
nor I_742 (I13993,I14076,I14477);
not I_743 (I14535,I1869);
or I_744 (I14552,I388010,I388010);
nand I_745 (I14569,I388025,I388028);
not I_746 (I14586,I14569);
nand I_747 (I14603,I14586,I14552);
not I_748 (I14620,I14603);
nand I_749 (I14637,I388016,I388019);
and I_750 (I14654,I14637,I388013);
DFFARX1 I_751 (I14654,I1862,I14535,I14680,);
not I_752 (I14688,I14680);
nor I_753 (I14705,I388019,I388019);
nor I_754 (I14722,I14680,I14705);
and I_755 (I14739,I14680,I14705);
nor I_756 (I14756,I14739,I14603);
DFFARX1 I_757 (I14756,I1862,I14535,I14515,);
nand I_758 (I14787,I388022,I388016);
nor I_759 (I14804,I14787,I388013);
nand I_760 (I14821,I14620,I14804);
not I_761 (I14524,I14821);
nor I_762 (I14527,I14722,I14821);
nor I_763 (I14866,I14804,I14586);
nor I_764 (I14518,I14688,I14866);
nor I_765 (I14512,I14804,I14705);
not I_766 (I14911,I14787);
nand I_767 (I14928,I14705,I14911);
not I_768 (I14506,I14928);
nor I_769 (I14509,I14569,I14928);
nor I_770 (I14521,I14911,I14569);
nand I_771 (I14987,I14688,I14787);
nor I_772 (I14503,I14586,I14987);
not I_773 (I15045,I1869);
or I_774 (I15062,I109165,I109159);
nand I_775 (I15079,I109165,I109177);
not I_776 (I15096,I15079);
nand I_777 (I15113,I15096,I15062);
not I_778 (I15130,I15113);
nand I_779 (I15147,I109171,I109162);
and I_780 (I15164,I15147,I109159);
DFFARX1 I_781 (I15164,I1862,I15045,I15190,);
not I_782 (I15198,I15190);
nor I_783 (I15215,I109174,I109162);
nor I_784 (I15232,I15190,I15215);
and I_785 (I15249,I15190,I15215);
nor I_786 (I15266,I15249,I15113);
DFFARX1 I_787 (I15266,I1862,I15045,I15025,);
nand I_788 (I15297,I109168,I109168);
nor I_789 (I15314,I15297,I109162);
nand I_790 (I15331,I15130,I15314);
not I_791 (I15034,I15331);
nor I_792 (I15037,I15232,I15331);
nor I_793 (I15376,I15314,I15096);
nor I_794 (I15028,I15198,I15376);
nor I_795 (I15022,I15314,I15215);
not I_796 (I15421,I15297);
nand I_797 (I15438,I15215,I15421);
not I_798 (I15016,I15438);
nor I_799 (I15019,I15079,I15438);
nor I_800 (I15031,I15421,I15079);
nand I_801 (I15497,I15198,I15297);
nor I_802 (I15013,I15096,I15497);
not I_803 (I15555,I1869);
or I_804 (I15572,I335758,I335752);
nand I_805 (I15589,I335761,I335764);
not I_806 (I15606,I15589);
nand I_807 (I15623,I15606,I15572);
not I_808 (I15640,I15623);
nand I_809 (I15657,I335755,I335758);
and I_810 (I15674,I15657,I335752);
DFFARX1 I_811 (I15674,I1862,I15555,I15700,);
not I_812 (I15708,I15700);
nor I_813 (I15725,I335770,I335758);
nor I_814 (I15742,I15700,I15725);
and I_815 (I15759,I15700,I15725);
nor I_816 (I15776,I15759,I15623);
DFFARX1 I_817 (I15776,I1862,I15555,I15535,);
nand I_818 (I15807,I335767,I335755);
nor I_819 (I15824,I15807,I335773);
nand I_820 (I15841,I15640,I15824);
not I_821 (I15544,I15841);
nor I_822 (I15547,I15742,I15841);
nor I_823 (I15886,I15824,I15606);
nor I_824 (I15538,I15708,I15886);
nor I_825 (I15532,I15824,I15725);
not I_826 (I15931,I15807);
nand I_827 (I15948,I15725,I15931);
not I_828 (I15526,I15948);
nor I_829 (I15529,I15589,I15948);
nor I_830 (I15541,I15931,I15589);
nand I_831 (I16007,I15708,I15807);
nor I_832 (I15523,I15606,I16007);
not I_833 (I16065,I1869);
or I_834 (I16082,I374750,I374750);
nand I_835 (I16099,I374765,I374768);
not I_836 (I16116,I16099);
nand I_837 (I16133,I16116,I16082);
not I_838 (I16150,I16133);
nand I_839 (I16167,I374756,I374759);
and I_840 (I16184,I16167,I374753);
DFFARX1 I_841 (I16184,I1862,I16065,I16210,);
not I_842 (I16218,I16210);
nor I_843 (I16235,I374759,I374759);
nor I_844 (I16252,I16210,I16235);
and I_845 (I16269,I16210,I16235);
nor I_846 (I16286,I16269,I16133);
DFFARX1 I_847 (I16286,I1862,I16065,I16045,);
nand I_848 (I16317,I374762,I374756);
nor I_849 (I16334,I16317,I374753);
nand I_850 (I16351,I16150,I16334);
not I_851 (I16054,I16351);
nor I_852 (I16057,I16252,I16351);
nor I_853 (I16396,I16334,I16116);
nor I_854 (I16048,I16218,I16396);
nor I_855 (I16042,I16334,I16235);
not I_856 (I16441,I16317);
nand I_857 (I16458,I16235,I16441);
not I_858 (I16036,I16458);
nor I_859 (I16039,I16099,I16458);
nor I_860 (I16051,I16441,I16099);
nand I_861 (I16517,I16218,I16317);
nor I_862 (I16033,I16116,I16517);
not I_863 (I16575,I1869);
or I_864 (I16592,I281032,I281035);
nand I_865 (I16609,I281041,I281029);
not I_866 (I16626,I16609);
nand I_867 (I16643,I16626,I16592);
not I_868 (I16660,I16643);
nand I_869 (I16677,I281047,I281050);
and I_870 (I16694,I16677,I281044);
DFFARX1 I_871 (I16694,I1862,I16575,I16720,);
not I_872 (I16728,I16720);
nor I_873 (I16745,I281032,I281050);
nor I_874 (I16762,I16720,I16745);
and I_875 (I16779,I16720,I16745);
nor I_876 (I16796,I16779,I16643);
DFFARX1 I_877 (I16796,I1862,I16575,I16555,);
nand I_878 (I16827,I281035,I281038);
nor I_879 (I16844,I16827,I281029);
nand I_880 (I16861,I16660,I16844);
not I_881 (I16564,I16861);
nor I_882 (I16567,I16762,I16861);
nor I_883 (I16906,I16844,I16626);
nor I_884 (I16558,I16728,I16906);
nor I_885 (I16552,I16844,I16745);
not I_886 (I16951,I16827);
nand I_887 (I16968,I16745,I16951);
not I_888 (I16546,I16968);
nor I_889 (I16549,I16609,I16968);
nor I_890 (I16561,I16951,I16609);
nand I_891 (I17027,I16728,I16827);
nor I_892 (I16543,I16626,I17027);
not I_893 (I17085,I1869);
or I_894 (I17102,I265800,I265803);
nand I_895 (I17119,I265809,I265797);
not I_896 (I17136,I17119);
nand I_897 (I17153,I17136,I17102);
not I_898 (I17170,I17153);
nand I_899 (I17187,I265815,I265818);
and I_900 (I17204,I17187,I265812);
DFFARX1 I_901 (I17204,I1862,I17085,I17230,);
not I_902 (I17238,I17230);
nor I_903 (I17255,I265800,I265818);
nor I_904 (I17272,I17230,I17255);
and I_905 (I17289,I17230,I17255);
nor I_906 (I17306,I17289,I17153);
DFFARX1 I_907 (I17306,I1862,I17085,I17065,);
nand I_908 (I17337,I265803,I265806);
nor I_909 (I17354,I17337,I265797);
nand I_910 (I17371,I17170,I17354);
not I_911 (I17074,I17371);
nor I_912 (I17077,I17272,I17371);
nor I_913 (I17416,I17354,I17136);
nor I_914 (I17068,I17238,I17416);
nor I_915 (I17062,I17354,I17255);
not I_916 (I17461,I17337);
nand I_917 (I17478,I17255,I17461);
not I_918 (I17056,I17478);
nor I_919 (I17059,I17119,I17478);
nor I_920 (I17071,I17461,I17119);
nand I_921 (I17537,I17238,I17337);
nor I_922 (I17053,I17136,I17537);
not I_923 (I17595,I1869);
or I_924 (I17612,I1031,I1527);
nand I_925 (I17629,I807,I1591);
not I_926 (I17646,I17629);
nand I_927 (I17663,I17646,I17612);
not I_928 (I17680,I17663);
nand I_929 (I17697,I1559,I1271);
and I_930 (I17714,I17697,I1407);
DFFARX1 I_931 (I17714,I1862,I17595,I17740,);
not I_932 (I17748,I17740);
nor I_933 (I17765,I935,I1271);
nor I_934 (I17782,I17740,I17765);
and I_935 (I17799,I17740,I17765);
nor I_936 (I17816,I17799,I17663);
DFFARX1 I_937 (I17816,I1862,I17595,I17575,);
nand I_938 (I17847,I871,I1255);
nor I_939 (I17864,I17847,I1119);
nand I_940 (I17881,I17680,I17864);
not I_941 (I17584,I17881);
nor I_942 (I17587,I17782,I17881);
nor I_943 (I17926,I17864,I17646);
nor I_944 (I17578,I17748,I17926);
nor I_945 (I17572,I17864,I17765);
not I_946 (I17971,I17847);
nand I_947 (I17988,I17765,I17971);
not I_948 (I17566,I17988);
nor I_949 (I17569,I17629,I17988);
nor I_950 (I17581,I17971,I17629);
nand I_951 (I18047,I17748,I17847);
nor I_952 (I17563,I17646,I18047);
not I_953 (I18105,I1869);
or I_954 (I18122,I228672,I228675);
nand I_955 (I18139,I228681,I228669);
not I_956 (I18156,I18139);
nand I_957 (I18173,I18156,I18122);
not I_958 (I18190,I18173);
nand I_959 (I18207,I228687,I228690);
and I_960 (I18224,I18207,I228684);
DFFARX1 I_961 (I18224,I1862,I18105,I18250,);
not I_962 (I18258,I18250);
nor I_963 (I18275,I228672,I228690);
nor I_964 (I18292,I18250,I18275);
and I_965 (I18309,I18250,I18275);
nor I_966 (I18326,I18309,I18173);
DFFARX1 I_967 (I18326,I1862,I18105,I18085,);
nand I_968 (I18357,I228675,I228678);
nor I_969 (I18374,I18357,I228669);
nand I_970 (I18391,I18190,I18374);
not I_971 (I18094,I18391);
nor I_972 (I18097,I18292,I18391);
nor I_973 (I18436,I18374,I18156);
nor I_974 (I18088,I18258,I18436);
nor I_975 (I18082,I18374,I18275);
not I_976 (I18481,I18357);
nand I_977 (I18498,I18275,I18481);
not I_978 (I18076,I18498);
nor I_979 (I18079,I18139,I18498);
nor I_980 (I18091,I18481,I18139);
nand I_981 (I18557,I18258,I18357);
nor I_982 (I18073,I18156,I18557);
not I_983 (I18615,I1869);
or I_984 (I18632,I333123,I333117);
nand I_985 (I18649,I333126,I333129);
not I_986 (I18666,I18649);
nand I_987 (I18683,I18666,I18632);
not I_988 (I18700,I18683);
nand I_989 (I18717,I333120,I333123);
and I_990 (I18734,I18717,I333117);
DFFARX1 I_991 (I18734,I1862,I18615,I18760,);
not I_992 (I18768,I18760);
nor I_993 (I18785,I333135,I333123);
nor I_994 (I18802,I18760,I18785);
and I_995 (I18819,I18760,I18785);
nor I_996 (I18836,I18819,I18683);
DFFARX1 I_997 (I18836,I1862,I18615,I18595,);
nand I_998 (I18867,I333132,I333120);
nor I_999 (I18884,I18867,I333138);
nand I_1000 (I18901,I18700,I18884);
not I_1001 (I18604,I18901);
nor I_1002 (I18607,I18802,I18901);
nor I_1003 (I18946,I18884,I18666);
nor I_1004 (I18598,I18768,I18946);
nor I_1005 (I18592,I18884,I18785);
not I_1006 (I18991,I18867);
nand I_1007 (I19008,I18785,I18991);
not I_1008 (I18586,I19008);
nor I_1009 (I18589,I18649,I19008);
nor I_1010 (I18601,I18991,I18649);
nand I_1011 (I19067,I18768,I18867);
nor I_1012 (I18583,I18666,I19067);
not I_1013 (I19125,I1869);
or I_1014 (I19142,I224864,I224867);
nand I_1015 (I19159,I224873,I224861);
not I_1016 (I19176,I19159);
nand I_1017 (I19193,I19176,I19142);
not I_1018 (I19210,I19193);
nand I_1019 (I19227,I224879,I224882);
and I_1020 (I19244,I19227,I224876);
DFFARX1 I_1021 (I19244,I1862,I19125,I19270,);
not I_1022 (I19278,I19270);
nor I_1023 (I19295,I224864,I224882);
nor I_1024 (I19312,I19270,I19295);
and I_1025 (I19329,I19270,I19295);
nor I_1026 (I19346,I19329,I19193);
DFFARX1 I_1027 (I19346,I1862,I19125,I19105,);
nand I_1028 (I19377,I224867,I224870);
nor I_1029 (I19394,I19377,I224861);
nand I_1030 (I19411,I19210,I19394);
not I_1031 (I19114,I19411);
nor I_1032 (I19117,I19312,I19411);
nor I_1033 (I19456,I19394,I19176);
nor I_1034 (I19108,I19278,I19456);
nor I_1035 (I19102,I19394,I19295);
not I_1036 (I19501,I19377);
nand I_1037 (I19518,I19295,I19501);
not I_1038 (I19096,I19518);
nor I_1039 (I19099,I19159,I19518);
nor I_1040 (I19111,I19501,I19159);
nand I_1041 (I19577,I19278,I19377);
nor I_1042 (I19093,I19176,I19577);
not I_1043 (I19635,I1869);
or I_1044 (I19652,I331542,I331536);
nand I_1045 (I19669,I331545,I331548);
not I_1046 (I19686,I19669);
nand I_1047 (I19703,I19686,I19652);
not I_1048 (I19720,I19703);
nand I_1049 (I19737,I331539,I331542);
and I_1050 (I19754,I19737,I331536);
DFFARX1 I_1051 (I19754,I1862,I19635,I19780,);
not I_1052 (I19788,I19780);
nor I_1053 (I19805,I331554,I331542);
nor I_1054 (I19822,I19780,I19805);
and I_1055 (I19839,I19780,I19805);
nor I_1056 (I19856,I19839,I19703);
DFFARX1 I_1057 (I19856,I1862,I19635,I19615,);
nand I_1058 (I19887,I331551,I331539);
nor I_1059 (I19904,I19887,I331557);
nand I_1060 (I19921,I19720,I19904);
not I_1061 (I19624,I19921);
nor I_1062 (I19627,I19822,I19921);
nor I_1063 (I19966,I19904,I19686);
nor I_1064 (I19618,I19788,I19966);
nor I_1065 (I19612,I19904,I19805);
not I_1066 (I20011,I19887);
nand I_1067 (I20028,I19805,I20011);
not I_1068 (I19606,I20028);
nor I_1069 (I19609,I19669,I20028);
nor I_1070 (I19621,I20011,I19669);
nand I_1071 (I20087,I19788,I19887);
nor I_1072 (I19603,I19686,I20087);
not I_1073 (I20145,I1869);
or I_1074 (I20162,I257232,I257235);
nand I_1075 (I20179,I257241,I257229);
not I_1076 (I20196,I20179);
nand I_1077 (I20213,I20196,I20162);
not I_1078 (I20230,I20213);
nand I_1079 (I20247,I257247,I257250);
and I_1080 (I20264,I20247,I257244);
DFFARX1 I_1081 (I20264,I1862,I20145,I20290,);
not I_1082 (I20298,I20290);
nor I_1083 (I20315,I257232,I257250);
nor I_1084 (I20332,I20290,I20315);
and I_1085 (I20349,I20290,I20315);
nor I_1086 (I20366,I20349,I20213);
DFFARX1 I_1087 (I20366,I1862,I20145,I20125,);
nand I_1088 (I20397,I257235,I257238);
nor I_1089 (I20414,I20397,I257229);
nand I_1090 (I20431,I20230,I20414);
not I_1091 (I20134,I20431);
nor I_1092 (I20137,I20332,I20431);
nor I_1093 (I20476,I20414,I20196);
nor I_1094 (I20128,I20298,I20476);
nor I_1095 (I20122,I20414,I20315);
not I_1096 (I20521,I20397);
nand I_1097 (I20538,I20315,I20521);
not I_1098 (I20116,I20538);
nor I_1099 (I20119,I20179,I20538);
nor I_1100 (I20131,I20521,I20179);
nand I_1101 (I20597,I20298,I20397);
nor I_1102 (I20113,I20196,I20597);
not I_1103 (I20655,I1869);
or I_1104 (I20672,I238192,I238195);
nand I_1105 (I20689,I238201,I238189);
not I_1106 (I20706,I20689);
nand I_1107 (I20723,I20706,I20672);
not I_1108 (I20740,I20723);
nand I_1109 (I20757,I238207,I238210);
and I_1110 (I20774,I20757,I238204);
DFFARX1 I_1111 (I20774,I1862,I20655,I20800,);
not I_1112 (I20808,I20800);
nor I_1113 (I20825,I238192,I238210);
nor I_1114 (I20842,I20800,I20825);
and I_1115 (I20859,I20800,I20825);
nor I_1116 (I20876,I20859,I20723);
DFFARX1 I_1117 (I20876,I1862,I20655,I20635,);
nand I_1118 (I20907,I238195,I238198);
nor I_1119 (I20924,I20907,I238189);
nand I_1120 (I20941,I20740,I20924);
not I_1121 (I20644,I20941);
nor I_1122 (I20647,I20842,I20941);
nor I_1123 (I20986,I20924,I20706);
nor I_1124 (I20638,I20808,I20986);
nor I_1125 (I20632,I20924,I20825);
not I_1126 (I21031,I20907);
nand I_1127 (I21048,I20825,I21031);
not I_1128 (I20626,I21048);
nor I_1129 (I20629,I20689,I21048);
nor I_1130 (I20641,I21031,I20689);
nand I_1131 (I21107,I20808,I20907);
nor I_1132 (I20623,I20706,I21107);
not I_1133 (I21165,I1869);
or I_1134 (I21182,I331015,I331009);
nand I_1135 (I21199,I331018,I331021);
not I_1136 (I21216,I21199);
nand I_1137 (I21233,I21216,I21182);
not I_1138 (I21250,I21233);
nand I_1139 (I21267,I331012,I331015);
and I_1140 (I21284,I21267,I331009);
DFFARX1 I_1141 (I21284,I1862,I21165,I21310,);
not I_1142 (I21318,I21310);
nor I_1143 (I21335,I331027,I331015);
nor I_1144 (I21352,I21310,I21335);
and I_1145 (I21369,I21310,I21335);
nor I_1146 (I21386,I21369,I21233);
DFFARX1 I_1147 (I21386,I1862,I21165,I21145,);
nand I_1148 (I21417,I331024,I331012);
nor I_1149 (I21434,I21417,I331030);
nand I_1150 (I21451,I21250,I21434);
not I_1151 (I21154,I21451);
nor I_1152 (I21157,I21352,I21451);
nor I_1153 (I21496,I21434,I21216);
nor I_1154 (I21148,I21318,I21496);
nor I_1155 (I21142,I21434,I21335);
not I_1156 (I21541,I21417);
nand I_1157 (I21558,I21335,I21541);
not I_1158 (I21136,I21558);
nor I_1159 (I21139,I21199,I21558);
nor I_1160 (I21151,I21541,I21199);
nand I_1161 (I21617,I21318,I21417);
nor I_1162 (I21133,I21216,I21617);
not I_1163 (I21675,I1869);
or I_1164 (I21692,I1607,I991);
nand I_1165 (I21709,I1287,I1623);
not I_1166 (I21726,I21709);
nand I_1167 (I21743,I21726,I21692);
not I_1168 (I21760,I21743);
nand I_1169 (I21777,I1223,I1303);
and I_1170 (I21794,I21777,I1847);
DFFARX1 I_1171 (I21794,I1862,I21675,I21820,);
not I_1172 (I21828,I21820);
nor I_1173 (I21845,I1095,I1303);
nor I_1174 (I21862,I21820,I21845);
and I_1175 (I21879,I21820,I21845);
nor I_1176 (I21896,I21879,I21743);
DFFARX1 I_1177 (I21896,I1862,I21675,I21655,);
nand I_1178 (I21927,I639,I695);
nor I_1179 (I21944,I21927,I1799);
nand I_1180 (I21961,I21760,I21944);
not I_1181 (I21664,I21961);
nor I_1182 (I21667,I21862,I21961);
nor I_1183 (I22006,I21944,I21726);
nor I_1184 (I21658,I21828,I22006);
nor I_1185 (I21652,I21944,I21845);
not I_1186 (I22051,I21927);
nand I_1187 (I22068,I21845,I22051);
not I_1188 (I21646,I22068);
nor I_1189 (I21649,I21709,I22068);
nor I_1190 (I21661,I22051,I21709);
nand I_1191 (I22127,I21828,I21927);
nor I_1192 (I21643,I21726,I22127);
not I_1193 (I22185,I1869);
or I_1194 (I22202,I176894,I176873);
nand I_1195 (I22219,I176882,I176891);
not I_1196 (I22236,I22219);
nand I_1197 (I22253,I22236,I22202);
not I_1198 (I22270,I22253);
nand I_1199 (I22287,I176888,I176873);
and I_1200 (I22304,I22287,I176879);
DFFARX1 I_1201 (I22304,I1862,I22185,I22330,);
not I_1202 (I22338,I22330);
nor I_1203 (I22355,I176870,I176873);
nor I_1204 (I22372,I22330,I22355);
and I_1205 (I22389,I22330,I22355);
nor I_1206 (I22406,I22389,I22253);
DFFARX1 I_1207 (I22406,I1862,I22185,I22165,);
nand I_1208 (I22437,I176885,I176870);
nor I_1209 (I22454,I22437,I176876);
nand I_1210 (I22471,I22270,I22454);
not I_1211 (I22174,I22471);
nor I_1212 (I22177,I22372,I22471);
nor I_1213 (I22516,I22454,I22236);
nor I_1214 (I22168,I22338,I22516);
nor I_1215 (I22162,I22454,I22355);
not I_1216 (I22561,I22437);
nand I_1217 (I22578,I22355,I22561);
not I_1218 (I22156,I22578);
nor I_1219 (I22159,I22219,I22578);
nor I_1220 (I22171,I22561,I22219);
nand I_1221 (I22637,I22338,I22437);
nor I_1222 (I22153,I22236,I22637);
not I_1223 (I22695,I1869);
or I_1224 (I22712,I282460,I282463);
nand I_1225 (I22729,I282469,I282457);
not I_1226 (I22746,I22729);
nand I_1227 (I22763,I22746,I22712);
not I_1228 (I22780,I22763);
nand I_1229 (I22797,I282475,I282478);
and I_1230 (I22814,I22797,I282472);
DFFARX1 I_1231 (I22814,I1862,I22695,I22840,);
not I_1232 (I22848,I22840);
nor I_1233 (I22865,I282460,I282478);
nor I_1234 (I22882,I22840,I22865);
and I_1235 (I22899,I22840,I22865);
nor I_1236 (I22916,I22899,I22763);
DFFARX1 I_1237 (I22916,I1862,I22695,I22675,);
nand I_1238 (I22947,I282463,I282466);
nor I_1239 (I22964,I22947,I282457);
nand I_1240 (I22981,I22780,I22964);
not I_1241 (I22684,I22981);
nor I_1242 (I22687,I22882,I22981);
nor I_1243 (I23026,I22964,I22746);
nor I_1244 (I22678,I22848,I23026);
nor I_1245 (I22672,I22964,I22865);
not I_1246 (I23071,I22947);
nand I_1247 (I23088,I22865,I23071);
not I_1248 (I22666,I23088);
nor I_1249 (I22669,I22729,I23088);
nor I_1250 (I22681,I23071,I22729);
nand I_1251 (I23147,I22848,I22947);
nor I_1252 (I22663,I22746,I23147);
not I_1253 (I23205,I1869);
or I_1254 (I23222,I369446,I369446);
nand I_1255 (I23239,I369461,I369464);
not I_1256 (I23256,I23239);
nand I_1257 (I23273,I23256,I23222);
not I_1258 (I23290,I23273);
nand I_1259 (I23307,I369452,I369455);
and I_1260 (I23324,I23307,I369449);
DFFARX1 I_1261 (I23324,I1862,I23205,I23350,);
not I_1262 (I23358,I23350);
nor I_1263 (I23375,I369455,I369455);
nor I_1264 (I23392,I23350,I23375);
and I_1265 (I23409,I23350,I23375);
nor I_1266 (I23426,I23409,I23273);
DFFARX1 I_1267 (I23426,I1862,I23205,I23185,);
nand I_1268 (I23457,I369458,I369452);
nor I_1269 (I23474,I23457,I369449);
nand I_1270 (I23491,I23290,I23474);
not I_1271 (I23194,I23491);
nor I_1272 (I23197,I23392,I23491);
nor I_1273 (I23536,I23474,I23256);
nor I_1274 (I23188,I23358,I23536);
nor I_1275 (I23182,I23474,I23375);
not I_1276 (I23581,I23457);
nand I_1277 (I23598,I23375,I23581);
not I_1278 (I23176,I23598);
nor I_1279 (I23179,I23239,I23598);
nor I_1280 (I23191,I23581,I23239);
nand I_1281 (I23657,I23358,I23457);
nor I_1282 (I23173,I23256,I23657);
not I_1283 (I23715,I1869);
or I_1284 (I23732,I214392,I214395);
nand I_1285 (I23749,I214401,I214389);
not I_1286 (I23766,I23749);
nand I_1287 (I23783,I23766,I23732);
not I_1288 (I23800,I23783);
nand I_1289 (I23817,I214407,I214410);
and I_1290 (I23834,I23817,I214404);
DFFARX1 I_1291 (I23834,I1862,I23715,I23860,);
not I_1292 (I23868,I23860);
nor I_1293 (I23885,I214392,I214410);
nor I_1294 (I23902,I23860,I23885);
and I_1295 (I23919,I23860,I23885);
nor I_1296 (I23936,I23919,I23783);
DFFARX1 I_1297 (I23936,I1862,I23715,I23695,);
nand I_1298 (I23967,I214395,I214398);
nor I_1299 (I23984,I23967,I214389);
nand I_1300 (I24001,I23800,I23984);
not I_1301 (I23704,I24001);
nor I_1302 (I23707,I23902,I24001);
nor I_1303 (I24046,I23984,I23766);
nor I_1304 (I23698,I23868,I24046);
nor I_1305 (I23692,I23984,I23885);
not I_1306 (I24091,I23967);
nand I_1307 (I24108,I23885,I24091);
not I_1308 (I23686,I24108);
nor I_1309 (I23689,I23749,I24108);
nor I_1310 (I23701,I24091,I23749);
nand I_1311 (I24167,I23868,I23967);
nor I_1312 (I23683,I23766,I24167);
not I_1313 (I24225,I1869);
or I_1314 (I24242,I105085,I105079);
nand I_1315 (I24259,I105085,I105097);
not I_1316 (I24276,I24259);
nand I_1317 (I24293,I24276,I24242);
not I_1318 (I24310,I24293);
nand I_1319 (I24327,I105091,I105082);
and I_1320 (I24344,I24327,I105079);
DFFARX1 I_1321 (I24344,I1862,I24225,I24370,);
not I_1322 (I24378,I24370);
nor I_1323 (I24395,I105094,I105082);
nor I_1324 (I24412,I24370,I24395);
and I_1325 (I24429,I24370,I24395);
nor I_1326 (I24446,I24429,I24293);
DFFARX1 I_1327 (I24446,I1862,I24225,I24205,);
nand I_1328 (I24477,I105088,I105088);
nor I_1329 (I24494,I24477,I105082);
nand I_1330 (I24511,I24310,I24494);
not I_1331 (I24214,I24511);
nor I_1332 (I24217,I24412,I24511);
nor I_1333 (I24556,I24494,I24276);
nor I_1334 (I24208,I24378,I24556);
nor I_1335 (I24202,I24494,I24395);
not I_1336 (I24601,I24477);
nand I_1337 (I24618,I24395,I24601);
not I_1338 (I24196,I24618);
nor I_1339 (I24199,I24259,I24618);
nor I_1340 (I24211,I24601,I24259);
nand I_1341 (I24677,I24378,I24477);
nor I_1342 (I24193,I24276,I24677);
not I_1343 (I24735,I1869);
or I_1344 (I24752,I312043,I312037);
nand I_1345 (I24769,I312046,I312049);
not I_1346 (I24786,I24769);
nand I_1347 (I24803,I24786,I24752);
not I_1348 (I24820,I24803);
nand I_1349 (I24837,I312040,I312043);
and I_1350 (I24854,I24837,I312037);
DFFARX1 I_1351 (I24854,I1862,I24735,I24880,);
not I_1352 (I24888,I24880);
nor I_1353 (I24905,I312055,I312043);
nor I_1354 (I24922,I24880,I24905);
and I_1355 (I24939,I24880,I24905);
nor I_1356 (I24956,I24939,I24803);
DFFARX1 I_1357 (I24956,I1862,I24735,I24715,);
nand I_1358 (I24987,I312052,I312040);
nor I_1359 (I25004,I24987,I312058);
nand I_1360 (I25021,I24820,I25004);
not I_1361 (I24724,I25021);
nor I_1362 (I24727,I24922,I25021);
nor I_1363 (I25066,I25004,I24786);
nor I_1364 (I24718,I24888,I25066);
nor I_1365 (I24712,I25004,I24905);
not I_1366 (I25111,I24987);
nand I_1367 (I25128,I24905,I25111);
not I_1368 (I24706,I25128);
nor I_1369 (I24709,I24769,I25128);
nor I_1370 (I24721,I25111,I24769);
nand I_1371 (I25187,I24888,I24987);
nor I_1372 (I24703,I24786,I25187);
not I_1373 (I25245,I1869);
or I_1374 (I25262,I346825,I346819);
nand I_1375 (I25279,I346828,I346831);
not I_1376 (I25296,I25279);
nand I_1377 (I25313,I25296,I25262);
not I_1378 (I25330,I25313);
nand I_1379 (I25347,I346822,I346825);
and I_1380 (I25364,I25347,I346819);
DFFARX1 I_1381 (I25364,I1862,I25245,I25390,);
not I_1382 (I25398,I25390);
nor I_1383 (I25415,I346837,I346825);
nor I_1384 (I25432,I25390,I25415);
and I_1385 (I25449,I25390,I25415);
nor I_1386 (I25466,I25449,I25313);
DFFARX1 I_1387 (I25466,I1862,I25245,I25225,);
nand I_1388 (I25497,I346834,I346822);
nor I_1389 (I25514,I25497,I346840);
nand I_1390 (I25531,I25330,I25514);
not I_1391 (I25234,I25531);
nor I_1392 (I25237,I25432,I25531);
nor I_1393 (I25576,I25514,I25296);
nor I_1394 (I25228,I25398,I25576);
nor I_1395 (I25222,I25514,I25415);
not I_1396 (I25621,I25497);
nand I_1397 (I25638,I25415,I25621);
not I_1398 (I25216,I25638);
nor I_1399 (I25219,I25279,I25638);
nor I_1400 (I25231,I25621,I25279);
nand I_1401 (I25697,I25398,I25497);
nor I_1402 (I25213,I25296,I25697);
not I_1403 (I25755,I1869);
or I_1404 (I25772,I126829,I126808);
nand I_1405 (I25789,I126817,I126826);
not I_1406 (I25806,I25789);
nand I_1407 (I25823,I25806,I25772);
not I_1408 (I25840,I25823);
nand I_1409 (I25857,I126823,I126808);
and I_1410 (I25874,I25857,I126814);
DFFARX1 I_1411 (I25874,I1862,I25755,I25900,);
not I_1412 (I25908,I25900);
nor I_1413 (I25925,I126805,I126808);
nor I_1414 (I25942,I25900,I25925);
and I_1415 (I25959,I25900,I25925);
nor I_1416 (I25976,I25959,I25823);
DFFARX1 I_1417 (I25976,I1862,I25755,I25735,);
nand I_1418 (I26007,I126820,I126805);
nor I_1419 (I26024,I26007,I126811);
nand I_1420 (I26041,I25840,I26024);
not I_1421 (I25744,I26041);
nor I_1422 (I25747,I25942,I26041);
nor I_1423 (I26086,I26024,I25806);
nor I_1424 (I25738,I25908,I26086);
nor I_1425 (I25732,I26024,I25925);
not I_1426 (I26131,I26007);
nand I_1427 (I26148,I25925,I26131);
not I_1428 (I25726,I26148);
nor I_1429 (I25729,I25789,I26148);
nor I_1430 (I25741,I26131,I25789);
nand I_1431 (I26207,I25908,I26007);
nor I_1432 (I25723,I25806,I26207);
not I_1433 (I26265,I1869);
or I_1434 (I26282,I189015,I188994);
nand I_1435 (I26299,I189003,I189012);
not I_1436 (I26316,I26299);
nand I_1437 (I26333,I26316,I26282);
not I_1438 (I26350,I26333);
nand I_1439 (I26367,I189009,I188994);
and I_1440 (I26384,I26367,I189000);
DFFARX1 I_1441 (I26384,I1862,I26265,I26410,);
not I_1442 (I26418,I26410);
nor I_1443 (I26435,I188991,I188994);
nor I_1444 (I26452,I26410,I26435);
and I_1445 (I26469,I26410,I26435);
nor I_1446 (I26486,I26469,I26333);
DFFARX1 I_1447 (I26486,I1862,I26265,I26245,);
nand I_1448 (I26517,I189006,I188991);
nor I_1449 (I26534,I26517,I188997);
nand I_1450 (I26551,I26350,I26534);
not I_1451 (I26254,I26551);
nor I_1452 (I26257,I26452,I26551);
nor I_1453 (I26596,I26534,I26316);
nor I_1454 (I26248,I26418,I26596);
nor I_1455 (I26242,I26534,I26435);
not I_1456 (I26641,I26517);
nand I_1457 (I26658,I26435,I26641);
not I_1458 (I26236,I26658);
nor I_1459 (I26239,I26299,I26658);
nor I_1460 (I26251,I26641,I26299);
nand I_1461 (I26717,I26418,I26517);
nor I_1462 (I26233,I26316,I26717);
not I_1463 (I26775,I1869);
or I_1464 (I26792,I107125,I107119);
nand I_1465 (I26809,I107125,I107137);
not I_1466 (I26826,I26809);
nand I_1467 (I26843,I26826,I26792);
not I_1468 (I26860,I26843);
nand I_1469 (I26877,I107131,I107122);
and I_1470 (I26894,I26877,I107119);
DFFARX1 I_1471 (I26894,I1862,I26775,I26920,);
not I_1472 (I26928,I26920);
nor I_1473 (I26945,I107134,I107122);
nor I_1474 (I26962,I26920,I26945);
and I_1475 (I26979,I26920,I26945);
nor I_1476 (I26996,I26979,I26843);
DFFARX1 I_1477 (I26996,I1862,I26775,I26755,);
nand I_1478 (I27027,I107128,I107128);
nor I_1479 (I27044,I27027,I107122);
nand I_1480 (I27061,I26860,I27044);
not I_1481 (I26764,I27061);
nor I_1482 (I26767,I26962,I27061);
nor I_1483 (I27106,I27044,I26826);
nor I_1484 (I26758,I26928,I27106);
nor I_1485 (I26752,I27044,I26945);
not I_1486 (I27151,I27027);
nand I_1487 (I27168,I26945,I27151);
not I_1488 (I26746,I27168);
nor I_1489 (I26749,I26809,I27168);
nor I_1490 (I26761,I27151,I26809);
nand I_1491 (I27227,I26928,I27027);
nor I_1492 (I26743,I26826,I27227);
not I_1493 (I27285,I1869);
or I_1494 (I27302,I182164,I182143);
nand I_1495 (I27319,I182152,I182161);
not I_1496 (I27336,I27319);
nand I_1497 (I27353,I27336,I27302);
not I_1498 (I27370,I27353);
nand I_1499 (I27387,I182158,I182143);
and I_1500 (I27404,I27387,I182149);
DFFARX1 I_1501 (I27404,I1862,I27285,I27430,);
not I_1502 (I27438,I27430);
nor I_1503 (I27455,I182140,I182143);
nor I_1504 (I27472,I27430,I27455);
and I_1505 (I27489,I27430,I27455);
nor I_1506 (I27506,I27489,I27353);
DFFARX1 I_1507 (I27506,I1862,I27285,I27265,);
nand I_1508 (I27537,I182155,I182140);
nor I_1509 (I27554,I27537,I182146);
nand I_1510 (I27571,I27370,I27554);
not I_1511 (I27274,I27571);
nor I_1512 (I27277,I27472,I27571);
nor I_1513 (I27616,I27554,I27336);
nor I_1514 (I27268,I27438,I27616);
nor I_1515 (I27262,I27554,I27455);
not I_1516 (I27661,I27537);
nand I_1517 (I27678,I27455,I27661);
not I_1518 (I27256,I27678);
nor I_1519 (I27259,I27319,I27678);
nor I_1520 (I27271,I27661,I27319);
nand I_1521 (I27737,I27438,I27537);
nor I_1522 (I27253,I27336,I27737);
not I_1523 (I27795,I1869);
or I_1524 (I27812,I107533,I107527);
nand I_1525 (I27829,I107533,I107545);
not I_1526 (I27846,I27829);
nand I_1527 (I27863,I27846,I27812);
not I_1528 (I27880,I27863);
nand I_1529 (I27897,I107539,I107530);
and I_1530 (I27914,I27897,I107527);
DFFARX1 I_1531 (I27914,I1862,I27795,I27940,);
not I_1532 (I27948,I27940);
nor I_1533 (I27965,I107542,I107530);
nor I_1534 (I27982,I27940,I27965);
and I_1535 (I27999,I27940,I27965);
nor I_1536 (I28016,I27999,I27863);
DFFARX1 I_1537 (I28016,I1862,I27795,I27775,);
nand I_1538 (I28047,I107536,I107536);
nor I_1539 (I28064,I28047,I107530);
nand I_1540 (I28081,I27880,I28064);
not I_1541 (I27784,I28081);
nor I_1542 (I27787,I27982,I28081);
nor I_1543 (I28126,I28064,I27846);
nor I_1544 (I27778,I27948,I28126);
nor I_1545 (I27772,I28064,I27965);
not I_1546 (I28171,I28047);
nand I_1547 (I28188,I27965,I28171);
not I_1548 (I27766,I28188);
nor I_1549 (I27769,I27829,I28188);
nor I_1550 (I27781,I28171,I27829);
nand I_1551 (I28247,I27948,I28047);
nor I_1552 (I27763,I27846,I28247);
not I_1553 (I28305,I1869);
or I_1554 (I28322,I276748,I276751);
nand I_1555 (I28339,I276757,I276745);
not I_1556 (I28356,I28339);
nand I_1557 (I28373,I28356,I28322);
not I_1558 (I28390,I28373);
nand I_1559 (I28407,I276763,I276766);
and I_1560 (I28424,I28407,I276760);
DFFARX1 I_1561 (I28424,I1862,I28305,I28450,);
not I_1562 (I28458,I28450);
nor I_1563 (I28475,I276748,I276766);
nor I_1564 (I28492,I28450,I28475);
and I_1565 (I28509,I28450,I28475);
nor I_1566 (I28526,I28509,I28373);
DFFARX1 I_1567 (I28526,I1862,I28305,I28285,);
nand I_1568 (I28557,I276751,I276754);
nor I_1569 (I28574,I28557,I276745);
nand I_1570 (I28591,I28390,I28574);
not I_1571 (I28294,I28591);
nor I_1572 (I28297,I28492,I28591);
nor I_1573 (I28636,I28574,I28356);
nor I_1574 (I28288,I28458,I28636);
nor I_1575 (I28282,I28574,I28475);
not I_1576 (I28681,I28557);
nand I_1577 (I28698,I28475,I28681);
not I_1578 (I28276,I28698);
nor I_1579 (I28279,I28339,I28698);
nor I_1580 (I28291,I28681,I28339);
nand I_1581 (I28757,I28458,I28557);
nor I_1582 (I28273,I28356,I28757);
not I_1583 (I28815,I1869);
or I_1584 (I28832,I159503,I159482);
nand I_1585 (I28849,I159491,I159500);
not I_1586 (I28866,I28849);
nand I_1587 (I28883,I28866,I28832);
not I_1588 (I28900,I28883);
nand I_1589 (I28917,I159497,I159482);
and I_1590 (I28934,I28917,I159488);
DFFARX1 I_1591 (I28934,I1862,I28815,I28960,);
not I_1592 (I28968,I28960);
nor I_1593 (I28985,I159479,I159482);
nor I_1594 (I29002,I28960,I28985);
and I_1595 (I29019,I28960,I28985);
nor I_1596 (I29036,I29019,I28883);
DFFARX1 I_1597 (I29036,I1862,I28815,I28795,);
nand I_1598 (I29067,I159494,I159479);
nor I_1599 (I29084,I29067,I159485);
nand I_1600 (I29101,I28900,I29084);
not I_1601 (I28804,I29101);
nor I_1602 (I28807,I29002,I29101);
nor I_1603 (I29146,I29084,I28866);
nor I_1604 (I28798,I28968,I29146);
nor I_1605 (I28792,I29084,I28985);
not I_1606 (I29191,I29067);
nand I_1607 (I29208,I28985,I29191);
not I_1608 (I28786,I29208);
nor I_1609 (I28789,I28849,I29208);
nor I_1610 (I28801,I29191,I28849);
nand I_1611 (I29267,I28968,I29067);
nor I_1612 (I28783,I28866,I29267);
not I_1613 (I29325,I1869);
or I_1614 (I29342,I296757,I296754);
nand I_1615 (I29359,I296760,I296772);
not I_1616 (I29376,I29359);
nand I_1617 (I29393,I29376,I29342);
not I_1618 (I29410,I29393);
nand I_1619 (I29427,I296757,I296763);
and I_1620 (I29444,I29427,I296769);
DFFARX1 I_1621 (I29444,I1862,I29325,I29470,);
not I_1622 (I29478,I29470);
nor I_1623 (I29495,I296775,I296763);
nor I_1624 (I29512,I29470,I29495);
and I_1625 (I29529,I29470,I29495);
nor I_1626 (I29546,I29529,I29393);
DFFARX1 I_1627 (I29546,I1862,I29325,I29305,);
nand I_1628 (I29577,I296766,I296760);
nor I_1629 (I29594,I29577,I296754);
nand I_1630 (I29611,I29410,I29594);
not I_1631 (I29314,I29611);
nor I_1632 (I29317,I29512,I29611);
nor I_1633 (I29656,I29594,I29376);
nor I_1634 (I29308,I29478,I29656);
nor I_1635 (I29302,I29594,I29495);
not I_1636 (I29701,I29577);
nand I_1637 (I29718,I29495,I29701);
not I_1638 (I29296,I29718);
nor I_1639 (I29299,I29359,I29718);
nor I_1640 (I29311,I29701,I29359);
nand I_1641 (I29777,I29478,I29577);
nor I_1642 (I29293,I29376,I29777);
not I_1643 (I29835,I1869);
or I_1644 (I29852,I361932,I361932);
nand I_1645 (I29869,I361947,I361950);
not I_1646 (I29886,I29869);
nand I_1647 (I29903,I29886,I29852);
not I_1648 (I29920,I29903);
nand I_1649 (I29937,I361938,I361941);
and I_1650 (I29954,I29937,I361935);
DFFARX1 I_1651 (I29954,I1862,I29835,I29980,);
not I_1652 (I29988,I29980);
nor I_1653 (I30005,I361941,I361941);
nor I_1654 (I30022,I29980,I30005);
and I_1655 (I30039,I29980,I30005);
nor I_1656 (I30056,I30039,I29903);
DFFARX1 I_1657 (I30056,I1862,I29835,I29815,);
nand I_1658 (I30087,I361944,I361938);
nor I_1659 (I30104,I30087,I361935);
nand I_1660 (I30121,I29920,I30104);
not I_1661 (I29824,I30121);
nor I_1662 (I29827,I30022,I30121);
nor I_1663 (I30166,I30104,I29886);
nor I_1664 (I29818,I29988,I30166);
nor I_1665 (I29812,I30104,I30005);
not I_1666 (I30211,I30087);
nand I_1667 (I30228,I30005,I30211);
not I_1668 (I29806,I30228);
nor I_1669 (I29809,I29869,I30228);
nor I_1670 (I29821,I30211,I29869);
nand I_1671 (I30287,I29988,I30087);
nor I_1672 (I29803,I29886,I30287);
not I_1673 (I30345,I1869);
or I_1674 (I30362,I134734,I134713);
nand I_1675 (I30379,I134722,I134731);
not I_1676 (I30396,I30379);
nand I_1677 (I30413,I30396,I30362);
not I_1678 (I30430,I30413);
nand I_1679 (I30447,I134728,I134713);
and I_1680 (I30464,I30447,I134719);
DFFARX1 I_1681 (I30464,I1862,I30345,I30490,);
not I_1682 (I30498,I30490);
nor I_1683 (I30515,I134710,I134713);
nor I_1684 (I30532,I30490,I30515);
and I_1685 (I30549,I30490,I30515);
nor I_1686 (I30566,I30549,I30413);
DFFARX1 I_1687 (I30566,I1862,I30345,I30325,);
nand I_1688 (I30597,I134725,I134710);
nor I_1689 (I30614,I30597,I134716);
nand I_1690 (I30631,I30430,I30614);
not I_1691 (I30334,I30631);
nor I_1692 (I30337,I30532,I30631);
nor I_1693 (I30676,I30614,I30396);
nor I_1694 (I30328,I30498,I30676);
nor I_1695 (I30322,I30614,I30515);
not I_1696 (I30721,I30597);
nand I_1697 (I30738,I30515,I30721);
not I_1698 (I30316,I30738);
nor I_1699 (I30319,I30379,I30738);
nor I_1700 (I30331,I30721,I30379);
nand I_1701 (I30797,I30498,I30597);
nor I_1702 (I30313,I30396,I30797);
not I_1703 (I30855,I1869);
or I_1704 (I30872,I251044,I251047);
nand I_1705 (I30889,I251053,I251041);
not I_1706 (I30906,I30889);
nand I_1707 (I30923,I30906,I30872);
not I_1708 (I30940,I30923);
nand I_1709 (I30957,I251059,I251062);
and I_1710 (I30974,I30957,I251056);
DFFARX1 I_1711 (I30974,I1862,I30855,I31000,);
not I_1712 (I31008,I31000);
nor I_1713 (I31025,I251044,I251062);
nor I_1714 (I31042,I31000,I31025);
and I_1715 (I31059,I31000,I31025);
nor I_1716 (I31076,I31059,I30923);
DFFARX1 I_1717 (I31076,I1862,I30855,I30835,);
nand I_1718 (I31107,I251047,I251050);
nor I_1719 (I31124,I31107,I251041);
nand I_1720 (I31141,I30940,I31124);
not I_1721 (I30844,I31141);
nor I_1722 (I30847,I31042,I31141);
nor I_1723 (I31186,I31124,I30906);
nor I_1724 (I30838,I31008,I31186);
nor I_1725 (I30832,I31124,I31025);
not I_1726 (I31231,I31107);
nand I_1727 (I31248,I31025,I31231);
not I_1728 (I30826,I31248);
nor I_1729 (I30829,I30889,I31248);
nor I_1730 (I30841,I31231,I30889);
nand I_1731 (I31307,I31008,I31107);
nor I_1732 (I30823,I30906,I31307);
not I_1733 (I31365,I1869);
or I_1734 (I31382,I170570,I170549);
nand I_1735 (I31399,I170558,I170567);
not I_1736 (I31416,I31399);
nand I_1737 (I31433,I31416,I31382);
not I_1738 (I31450,I31433);
nand I_1739 (I31467,I170564,I170549);
and I_1740 (I31484,I31467,I170555);
DFFARX1 I_1741 (I31484,I1862,I31365,I31510,);
not I_1742 (I31518,I31510);
nor I_1743 (I31535,I170546,I170549);
nor I_1744 (I31552,I31510,I31535);
and I_1745 (I31569,I31510,I31535);
nor I_1746 (I31586,I31569,I31433);
DFFARX1 I_1747 (I31586,I1862,I31365,I31345,);
nand I_1748 (I31617,I170561,I170546);
nor I_1749 (I31634,I31617,I170552);
nand I_1750 (I31651,I31450,I31634);
not I_1751 (I31354,I31651);
nor I_1752 (I31357,I31552,I31651);
nor I_1753 (I31696,I31634,I31416);
nor I_1754 (I31348,I31518,I31696);
nor I_1755 (I31342,I31634,I31535);
not I_1756 (I31741,I31617);
nand I_1757 (I31758,I31535,I31741);
not I_1758 (I31336,I31758);
nor I_1759 (I31339,I31399,I31758);
nor I_1760 (I31351,I31741,I31399);
nand I_1761 (I31817,I31518,I31617);
nor I_1762 (I31333,I31416,I31817);
not I_1763 (I31875,I1869);
or I_1764 (I31892,I161611,I161590);
nand I_1765 (I31909,I161599,I161608);
not I_1766 (I31926,I31909);
nand I_1767 (I31943,I31926,I31892);
not I_1768 (I31960,I31943);
nand I_1769 (I31977,I161605,I161590);
and I_1770 (I31994,I31977,I161596);
DFFARX1 I_1771 (I31994,I1862,I31875,I32020,);
not I_1772 (I32028,I32020);
nor I_1773 (I32045,I161587,I161590);
nor I_1774 (I32062,I32020,I32045);
and I_1775 (I32079,I32020,I32045);
nor I_1776 (I32096,I32079,I31943);
DFFARX1 I_1777 (I32096,I1862,I31875,I31855,);
nand I_1778 (I32127,I161602,I161587);
nor I_1779 (I32144,I32127,I161593);
nand I_1780 (I32161,I31960,I32144);
not I_1781 (I31864,I32161);
nor I_1782 (I31867,I32062,I32161);
nor I_1783 (I32206,I32144,I31926);
nor I_1784 (I31858,I32028,I32206);
nor I_1785 (I31852,I32144,I32045);
not I_1786 (I32251,I32127);
nand I_1787 (I32268,I32045,I32251);
not I_1788 (I31846,I32268);
nor I_1789 (I31849,I31909,I32268);
nor I_1790 (I31861,I32251,I31909);
nand I_1791 (I32327,I32028,I32127);
nor I_1792 (I31843,I31926,I32327);
not I_1793 (I32385,I1869);
or I_1794 (I32402,I161084,I161063);
nand I_1795 (I32419,I161072,I161081);
not I_1796 (I32436,I32419);
nand I_1797 (I32453,I32436,I32402);
not I_1798 (I32470,I32453);
nand I_1799 (I32487,I161078,I161063);
and I_1800 (I32504,I32487,I161069);
DFFARX1 I_1801 (I32504,I1862,I32385,I32530,);
not I_1802 (I32538,I32530);
nor I_1803 (I32555,I161060,I161063);
nor I_1804 (I32572,I32530,I32555);
and I_1805 (I32589,I32530,I32555);
nor I_1806 (I32606,I32589,I32453);
DFFARX1 I_1807 (I32606,I1862,I32385,I32365,);
nand I_1808 (I32637,I161075,I161060);
nor I_1809 (I32654,I32637,I161066);
nand I_1810 (I32671,I32470,I32654);
not I_1811 (I32374,I32671);
nor I_1812 (I32377,I32572,I32671);
nor I_1813 (I32716,I32654,I32436);
nor I_1814 (I32368,I32538,I32716);
nor I_1815 (I32362,I32654,I32555);
not I_1816 (I32761,I32637);
nand I_1817 (I32778,I32555,I32761);
not I_1818 (I32356,I32778);
nor I_1819 (I32359,I32419,I32778);
nor I_1820 (I32371,I32761,I32419);
nand I_1821 (I32837,I32538,I32637);
nor I_1822 (I32353,I32436,I32837);
not I_1823 (I32895,I1869);
or I_1824 (I32912,I402154,I402154);
nand I_1825 (I32929,I402169,I402172);
not I_1826 (I32946,I32929);
nand I_1827 (I32963,I32946,I32912);
not I_1828 (I32980,I32963);
nand I_1829 (I32997,I402160,I402163);
and I_1830 (I33014,I32997,I402157);
DFFARX1 I_1831 (I33014,I1862,I32895,I33040,);
not I_1832 (I33048,I33040);
nor I_1833 (I33065,I402163,I402163);
nor I_1834 (I33082,I33040,I33065);
and I_1835 (I33099,I33040,I33065);
nor I_1836 (I33116,I33099,I32963);
DFFARX1 I_1837 (I33116,I1862,I32895,I32875,);
nand I_1838 (I33147,I402166,I402160);
nor I_1839 (I33164,I33147,I402157);
nand I_1840 (I33181,I32980,I33164);
not I_1841 (I32884,I33181);
nor I_1842 (I32887,I33082,I33181);
nor I_1843 (I33226,I33164,I32946);
nor I_1844 (I32878,I33048,I33226);
nor I_1845 (I32872,I33164,I33065);
not I_1846 (I33271,I33147);
nand I_1847 (I33288,I33065,I33271);
not I_1848 (I32866,I33288);
nor I_1849 (I32869,I32929,I33288);
nor I_1850 (I32881,I33271,I32929);
nand I_1851 (I33347,I33048,I33147);
nor I_1852 (I32863,I32946,I33347);
not I_1853 (I33405,I1869);
or I_1854 (I33422,I124721,I124700);
nand I_1855 (I33439,I124709,I124718);
not I_1856 (I33456,I33439);
nand I_1857 (I33473,I33456,I33422);
not I_1858 (I33490,I33473);
nand I_1859 (I33507,I124715,I124700);
and I_1860 (I33524,I33507,I124706);
DFFARX1 I_1861 (I33524,I1862,I33405,I33550,);
not I_1862 (I33558,I33550);
nor I_1863 (I33575,I124697,I124700);
nor I_1864 (I33592,I33550,I33575);
and I_1865 (I33609,I33550,I33575);
nor I_1866 (I33626,I33609,I33473);
DFFARX1 I_1867 (I33626,I1862,I33405,I33385,);
nand I_1868 (I33657,I124712,I124697);
nor I_1869 (I33674,I33657,I124703);
nand I_1870 (I33691,I33490,I33674);
not I_1871 (I33394,I33691);
nor I_1872 (I33397,I33592,I33691);
nor I_1873 (I33736,I33674,I33456);
nor I_1874 (I33388,I33558,I33736);
nor I_1875 (I33382,I33674,I33575);
not I_1876 (I33781,I33657);
nand I_1877 (I33798,I33575,I33781);
not I_1878 (I33376,I33798);
nor I_1879 (I33379,I33439,I33798);
nor I_1880 (I33391,I33781,I33439);
nand I_1881 (I33857,I33558,I33657);
nor I_1882 (I33373,I33456,I33857);
not I_1883 (I33915,I1869);
or I_1884 (I33932,I305719,I305713);
nand I_1885 (I33949,I305722,I305725);
not I_1886 (I33966,I33949);
nand I_1887 (I33983,I33966,I33932);
not I_1888 (I34000,I33983);
nand I_1889 (I34017,I305716,I305719);
and I_1890 (I34034,I34017,I305713);
DFFARX1 I_1891 (I34034,I1862,I33915,I34060,);
not I_1892 (I34068,I34060);
nor I_1893 (I34085,I305731,I305719);
nor I_1894 (I34102,I34060,I34085);
and I_1895 (I34119,I34060,I34085);
nor I_1896 (I34136,I34119,I33983);
DFFARX1 I_1897 (I34136,I1862,I33915,I33895,);
nand I_1898 (I34167,I305728,I305716);
nor I_1899 (I34184,I34167,I305734);
nand I_1900 (I34201,I34000,I34184);
not I_1901 (I33904,I34201);
nor I_1902 (I33907,I34102,I34201);
nor I_1903 (I34246,I34184,I33966);
nor I_1904 (I33898,I34068,I34246);
nor I_1905 (I33892,I34184,I34085);
not I_1906 (I34291,I34167);
nand I_1907 (I34308,I34085,I34291);
not I_1908 (I33886,I34308);
nor I_1909 (I33889,I33949,I34308);
nor I_1910 (I33901,I34291,I33949);
nand I_1911 (I34367,I34068,I34167);
nor I_1912 (I33883,I33966,I34367);
not I_1913 (I34425,I1869);
or I_1914 (I34442,I370330,I370330);
nand I_1915 (I34459,I370345,I370348);
not I_1916 (I34476,I34459);
nand I_1917 (I34493,I34476,I34442);
not I_1918 (I34510,I34493);
nand I_1919 (I34527,I370336,I370339);
and I_1920 (I34544,I34527,I370333);
DFFARX1 I_1921 (I34544,I1862,I34425,I34570,);
not I_1922 (I34578,I34570);
nor I_1923 (I34595,I370339,I370339);
nor I_1924 (I34612,I34570,I34595);
and I_1925 (I34629,I34570,I34595);
nor I_1926 (I34646,I34629,I34493);
DFFARX1 I_1927 (I34646,I1862,I34425,I34405,);
nand I_1928 (I34677,I370342,I370336);
nor I_1929 (I34694,I34677,I370333);
nand I_1930 (I34711,I34510,I34694);
not I_1931 (I34414,I34711);
nor I_1932 (I34417,I34612,I34711);
nor I_1933 (I34756,I34694,I34476);
nor I_1934 (I34408,I34578,I34756);
nor I_1935 (I34402,I34694,I34595);
not I_1936 (I34801,I34677);
nand I_1937 (I34818,I34595,I34801);
not I_1938 (I34396,I34818);
nor I_1939 (I34399,I34459,I34818);
nor I_1940 (I34411,I34801,I34459);
nand I_1941 (I34877,I34578,I34677);
nor I_1942 (I34393,I34476,I34877);
not I_1943 (I34935,I1869);
or I_1944 (I34952,I303084,I303078);
nand I_1945 (I34969,I303087,I303090);
not I_1946 (I34986,I34969);
nand I_1947 (I35003,I34986,I34952);
not I_1948 (I35020,I35003);
nand I_1949 (I35037,I303081,I303084);
and I_1950 (I35054,I35037,I303078);
DFFARX1 I_1951 (I35054,I1862,I34935,I35080,);
not I_1952 (I35088,I35080);
nor I_1953 (I35105,I303096,I303084);
nor I_1954 (I35122,I35080,I35105);
and I_1955 (I35139,I35080,I35105);
nor I_1956 (I35156,I35139,I35003);
DFFARX1 I_1957 (I35156,I1862,I34935,I34915,);
nand I_1958 (I35187,I303093,I303081);
nor I_1959 (I35204,I35187,I303099);
nand I_1960 (I35221,I35020,I35204);
not I_1961 (I34924,I35221);
nor I_1962 (I34927,I35122,I35221);
nor I_1963 (I35266,I35204,I34986);
nor I_1964 (I34918,I35088,I35266);
nor I_1965 (I34912,I35204,I35105);
not I_1966 (I35311,I35187);
nand I_1967 (I35328,I35105,I35311);
not I_1968 (I34906,I35328);
nor I_1969 (I34909,I34969,I35328);
nor I_1970 (I34921,I35311,I34969);
nand I_1971 (I35387,I35088,I35187);
nor I_1972 (I34903,I34986,I35387);
not I_1973 (I35445,I1869);
or I_1974 (I35462,I212012,I212015);
nand I_1975 (I35479,I212021,I212009);
not I_1976 (I35496,I35479);
nand I_1977 (I35513,I35496,I35462);
not I_1978 (I35530,I35513);
nand I_1979 (I35547,I212027,I212030);
and I_1980 (I35564,I35547,I212024);
DFFARX1 I_1981 (I35564,I1862,I35445,I35590,);
not I_1982 (I35598,I35590);
nor I_1983 (I35615,I212012,I212030);
nor I_1984 (I35632,I35590,I35615);
and I_1985 (I35649,I35590,I35615);
nor I_1986 (I35666,I35649,I35513);
DFFARX1 I_1987 (I35666,I1862,I35445,I35425,);
nand I_1988 (I35697,I212015,I212018);
nor I_1989 (I35714,I35697,I212009);
nand I_1990 (I35731,I35530,I35714);
not I_1991 (I35434,I35731);
nor I_1992 (I35437,I35632,I35731);
nor I_1993 (I35776,I35714,I35496);
nor I_1994 (I35428,I35598,I35776);
nor I_1995 (I35422,I35714,I35615);
not I_1996 (I35821,I35697);
nand I_1997 (I35838,I35615,I35821);
not I_1998 (I35416,I35838);
nor I_1999 (I35419,I35479,I35838);
nor I_2000 (I35431,I35821,I35479);
nand I_2001 (I35897,I35598,I35697);
nor I_2002 (I35413,I35496,I35897);
not I_2003 (I35955,I1869);
or I_2004 (I35972,I195866,I195845);
nand I_2005 (I35989,I195854,I195863);
not I_2006 (I36006,I35989);
nand I_2007 (I36023,I36006,I35972);
not I_2008 (I36040,I36023);
nand I_2009 (I36057,I195860,I195845);
and I_2010 (I36074,I36057,I195851);
DFFARX1 I_2011 (I36074,I1862,I35955,I36100,);
not I_2012 (I36108,I36100);
nor I_2013 (I36125,I195842,I195845);
nor I_2014 (I36142,I36100,I36125);
and I_2015 (I36159,I36100,I36125);
nor I_2016 (I36176,I36159,I36023);
DFFARX1 I_2017 (I36176,I1862,I35955,I35935,);
nand I_2018 (I36207,I195857,I195842);
nor I_2019 (I36224,I36207,I195848);
nand I_2020 (I36241,I36040,I36224);
not I_2021 (I35944,I36241);
nor I_2022 (I35947,I36142,I36241);
nor I_2023 (I36286,I36224,I36006);
nor I_2024 (I35938,I36108,I36286);
nor I_2025 (I35932,I36224,I36125);
not I_2026 (I36331,I36207);
nand I_2027 (I36348,I36125,I36331);
not I_2028 (I35926,I36348);
nor I_2029 (I35929,I35989,I36348);
nor I_2030 (I35941,I36331,I35989);
nand I_2031 (I36407,I36108,I36207);
nor I_2032 (I35923,I36006,I36407);
not I_2033 (I36465,I1869);
or I_2034 (I36482,I210584,I210587);
nand I_2035 (I36499,I210593,I210581);
not I_2036 (I36516,I36499);
nand I_2037 (I36533,I36516,I36482);
not I_2038 (I36550,I36533);
nand I_2039 (I36567,I210599,I210602);
and I_2040 (I36584,I36567,I210596);
DFFARX1 I_2041 (I36584,I1862,I36465,I36610,);
not I_2042 (I36618,I36610);
nor I_2043 (I36635,I210584,I210602);
nor I_2044 (I36652,I36610,I36635);
and I_2045 (I36669,I36610,I36635);
nor I_2046 (I36686,I36669,I36533);
DFFARX1 I_2047 (I36686,I1862,I36465,I36445,);
nand I_2048 (I36717,I210587,I210590);
nor I_2049 (I36734,I36717,I210581);
nand I_2050 (I36751,I36550,I36734);
not I_2051 (I36454,I36751);
nor I_2052 (I36457,I36652,I36751);
nor I_2053 (I36796,I36734,I36516);
nor I_2054 (I36448,I36618,I36796);
nor I_2055 (I36442,I36734,I36635);
not I_2056 (I36841,I36717);
nand I_2057 (I36858,I36635,I36841);
not I_2058 (I36436,I36858);
nor I_2059 (I36439,I36499,I36858);
nor I_2060 (I36451,I36841,I36499);
nand I_2061 (I36917,I36618,I36717);
nor I_2062 (I36433,I36516,I36917);
not I_2063 (I36975,I1869);
or I_2064 (I36992,I225340,I225343);
nand I_2065 (I37009,I225349,I225337);
not I_2066 (I37026,I37009);
nand I_2067 (I37043,I37026,I36992);
not I_2068 (I37060,I37043);
nand I_2069 (I37077,I225355,I225358);
and I_2070 (I37094,I37077,I225352);
DFFARX1 I_2071 (I37094,I1862,I36975,I37120,);
not I_2072 (I37128,I37120);
nor I_2073 (I37145,I225340,I225358);
nor I_2074 (I37162,I37120,I37145);
and I_2075 (I37179,I37120,I37145);
nor I_2076 (I37196,I37179,I37043);
DFFARX1 I_2077 (I37196,I1862,I36975,I36955,);
nand I_2078 (I37227,I225343,I225346);
nor I_2079 (I37244,I37227,I225337);
nand I_2080 (I37261,I37060,I37244);
not I_2081 (I36964,I37261);
nor I_2082 (I36967,I37162,I37261);
nor I_2083 (I37306,I37244,I37026);
nor I_2084 (I36958,I37128,I37306);
nor I_2085 (I36952,I37244,I37145);
not I_2086 (I37351,I37227);
nand I_2087 (I37368,I37145,I37351);
not I_2088 (I36946,I37368);
nor I_2089 (I36949,I37009,I37368);
nor I_2090 (I36961,I37351,I37009);
nand I_2091 (I37427,I37128,I37227);
nor I_2092 (I36943,I37026,I37427);
not I_2093 (I37485,I1869);
or I_2094 (I37502,I175313,I175292);
nand I_2095 (I37519,I175301,I175310);
not I_2096 (I37536,I37519);
nand I_2097 (I37553,I37536,I37502);
not I_2098 (I37570,I37553);
nand I_2099 (I37587,I175307,I175292);
and I_2100 (I37604,I37587,I175298);
DFFARX1 I_2101 (I37604,I1862,I37485,I37630,);
not I_2102 (I37638,I37630);
nor I_2103 (I37655,I175289,I175292);
nor I_2104 (I37672,I37630,I37655);
and I_2105 (I37689,I37630,I37655);
nor I_2106 (I37706,I37689,I37553);
DFFARX1 I_2107 (I37706,I1862,I37485,I37465,);
nand I_2108 (I37737,I175304,I175289);
nor I_2109 (I37754,I37737,I175295);
nand I_2110 (I37771,I37570,I37754);
not I_2111 (I37474,I37771);
nor I_2112 (I37477,I37672,I37771);
nor I_2113 (I37816,I37754,I37536);
nor I_2114 (I37468,I37638,I37816);
nor I_2115 (I37462,I37754,I37655);
not I_2116 (I37861,I37737);
nand I_2117 (I37878,I37655,I37861);
not I_2118 (I37456,I37878);
nor I_2119 (I37459,I37519,I37878);
nor I_2120 (I37471,I37861,I37519);
nand I_2121 (I37937,I37638,I37737);
nor I_2122 (I37453,I37536,I37937);
not I_2123 (I37995,I1869);
or I_2124 (I38012,I402596,I402596);
nand I_2125 (I38029,I402611,I402614);
not I_2126 (I38046,I38029);
nand I_2127 (I38063,I38046,I38012);
not I_2128 (I38080,I38063);
nand I_2129 (I38097,I402602,I402605);
and I_2130 (I38114,I38097,I402599);
DFFARX1 I_2131 (I38114,I1862,I37995,I38140,);
not I_2132 (I38148,I38140);
nor I_2133 (I38165,I402605,I402605);
nor I_2134 (I38182,I38140,I38165);
and I_2135 (I38199,I38140,I38165);
nor I_2136 (I38216,I38199,I38063);
DFFARX1 I_2137 (I38216,I1862,I37995,I37975,);
nand I_2138 (I38247,I402608,I402602);
nor I_2139 (I38264,I38247,I402599);
nand I_2140 (I38281,I38080,I38264);
not I_2141 (I37984,I38281);
nor I_2142 (I37987,I38182,I38281);
nor I_2143 (I38326,I38264,I38046);
nor I_2144 (I37978,I38148,I38326);
nor I_2145 (I37972,I38264,I38165);
not I_2146 (I38371,I38247);
nand I_2147 (I38388,I38165,I38371);
not I_2148 (I37966,I38388);
nor I_2149 (I37969,I38029,I38388);
nor I_2150 (I37981,I38371,I38029);
nand I_2151 (I38447,I38148,I38247);
nor I_2152 (I37963,I38046,I38447);
not I_2153 (I38505,I1869);
or I_2154 (I38522,I281508,I281511);
nand I_2155 (I38539,I281517,I281505);
not I_2156 (I38556,I38539);
nand I_2157 (I38573,I38556,I38522);
not I_2158 (I38590,I38573);
nand I_2159 (I38607,I281523,I281526);
and I_2160 (I38624,I38607,I281520);
DFFARX1 I_2161 (I38624,I1862,I38505,I38650,);
not I_2162 (I38658,I38650);
nor I_2163 (I38675,I281508,I281526);
nor I_2164 (I38692,I38650,I38675);
and I_2165 (I38709,I38650,I38675);
nor I_2166 (I38726,I38709,I38573);
DFFARX1 I_2167 (I38726,I1862,I38505,I38485,);
nand I_2168 (I38757,I281511,I281514);
nor I_2169 (I38774,I38757,I281505);
nand I_2170 (I38791,I38590,I38774);
not I_2171 (I38494,I38791);
nor I_2172 (I38497,I38692,I38791);
nor I_2173 (I38836,I38774,I38556);
nor I_2174 (I38488,I38658,I38836);
nor I_2175 (I38482,I38774,I38675);
not I_2176 (I38881,I38757);
nand I_2177 (I38898,I38675,I38881);
not I_2178 (I38476,I38898);
nor I_2179 (I38479,I38539,I38898);
nor I_2180 (I38491,I38881,I38539);
nand I_2181 (I38957,I38658,I38757);
nor I_2182 (I38473,I38556,I38957);
not I_2183 (I39015,I1869);
or I_2184 (I39032,I407016,I407016);
nand I_2185 (I39049,I407031,I407034);
not I_2186 (I39066,I39049);
nand I_2187 (I39083,I39066,I39032);
not I_2188 (I39100,I39083);
nand I_2189 (I39117,I407022,I407025);
and I_2190 (I39134,I39117,I407019);
DFFARX1 I_2191 (I39134,I1862,I39015,I39160,);
not I_2192 (I39168,I39160);
nor I_2193 (I39185,I407025,I407025);
nor I_2194 (I39202,I39160,I39185);
and I_2195 (I39219,I39160,I39185);
nor I_2196 (I39236,I39219,I39083);
DFFARX1 I_2197 (I39236,I1862,I39015,I38995,);
nand I_2198 (I39267,I407028,I407022);
nor I_2199 (I39284,I39267,I407019);
nand I_2200 (I39301,I39100,I39284);
not I_2201 (I39004,I39301);
nor I_2202 (I39007,I39202,I39301);
nor I_2203 (I39346,I39284,I39066);
nor I_2204 (I38998,I39168,I39346);
nor I_2205 (I38992,I39284,I39185);
not I_2206 (I39391,I39267);
nand I_2207 (I39408,I39185,I39391);
not I_2208 (I38986,I39408);
nor I_2209 (I38989,I39049,I39408);
nor I_2210 (I39001,I39391,I39049);
nand I_2211 (I39467,I39168,I39267);
nor I_2212 (I38983,I39066,I39467);
not I_2213 (I39525,I1869);
or I_2214 (I39542,I410552,I410552);
nand I_2215 (I39559,I410567,I410570);
not I_2216 (I39576,I39559);
nand I_2217 (I39593,I39576,I39542);
not I_2218 (I39610,I39593);
nand I_2219 (I39627,I410558,I410561);
and I_2220 (I39644,I39627,I410555);
DFFARX1 I_2221 (I39644,I1862,I39525,I39670,);
not I_2222 (I39678,I39670);
nor I_2223 (I39695,I410561,I410561);
nor I_2224 (I39712,I39670,I39695);
and I_2225 (I39729,I39670,I39695);
nor I_2226 (I39746,I39729,I39593);
DFFARX1 I_2227 (I39746,I1862,I39525,I39505,);
nand I_2228 (I39777,I410564,I410558);
nor I_2229 (I39794,I39777,I410555);
nand I_2230 (I39811,I39610,I39794);
not I_2231 (I39514,I39811);
nor I_2232 (I39517,I39712,I39811);
nor I_2233 (I39856,I39794,I39576);
nor I_2234 (I39508,I39678,I39856);
nor I_2235 (I39502,I39794,I39695);
not I_2236 (I39901,I39777);
nand I_2237 (I39918,I39695,I39901);
not I_2238 (I39496,I39918);
nor I_2239 (I39499,I39559,I39918);
nor I_2240 (I39511,I39901,I39559);
nand I_2241 (I39977,I39678,I39777);
nor I_2242 (I39493,I39576,I39977);
not I_2243 (I40035,I1869);
or I_2244 (I40052,I216296,I216299);
nand I_2245 (I40069,I216305,I216293);
not I_2246 (I40086,I40069);
nand I_2247 (I40103,I40086,I40052);
not I_2248 (I40120,I40103);
nand I_2249 (I40137,I216311,I216314);
and I_2250 (I40154,I40137,I216308);
DFFARX1 I_2251 (I40154,I1862,I40035,I40180,);
not I_2252 (I40188,I40180);
nor I_2253 (I40205,I216296,I216314);
nor I_2254 (I40222,I40180,I40205);
and I_2255 (I40239,I40180,I40205);
nor I_2256 (I40256,I40239,I40103);
DFFARX1 I_2257 (I40256,I1862,I40035,I40015,);
nand I_2258 (I40287,I216299,I216302);
nor I_2259 (I40304,I40287,I216293);
nand I_2260 (I40321,I40120,I40304);
not I_2261 (I40024,I40321);
nor I_2262 (I40027,I40222,I40321);
nor I_2263 (I40366,I40304,I40086);
nor I_2264 (I40018,I40188,I40366);
nor I_2265 (I40012,I40304,I40205);
not I_2266 (I40411,I40287);
nand I_2267 (I40428,I40205,I40411);
not I_2268 (I40006,I40428);
nor I_2269 (I40009,I40069,I40428);
nor I_2270 (I40021,I40411,I40069);
nand I_2271 (I40487,I40188,I40287);
nor I_2272 (I40003,I40086,I40487);
not I_2273 (I40545,I1869);
or I_2274 (I40562,I232480,I232483);
nand I_2275 (I40579,I232489,I232477);
not I_2276 (I40596,I40579);
nand I_2277 (I40613,I40596,I40562);
not I_2278 (I40630,I40613);
nand I_2279 (I40647,I232495,I232498);
and I_2280 (I40664,I40647,I232492);
DFFARX1 I_2281 (I40664,I1862,I40545,I40690,);
not I_2282 (I40698,I40690);
nor I_2283 (I40715,I232480,I232498);
nor I_2284 (I40732,I40690,I40715);
and I_2285 (I40749,I40690,I40715);
nor I_2286 (I40766,I40749,I40613);
DFFARX1 I_2287 (I40766,I1862,I40545,I40525,);
nand I_2288 (I40797,I232483,I232486);
nor I_2289 (I40814,I40797,I232477);
nand I_2290 (I40831,I40630,I40814);
not I_2291 (I40534,I40831);
nor I_2292 (I40537,I40732,I40831);
nor I_2293 (I40876,I40814,I40596);
nor I_2294 (I40528,I40698,I40876);
nor I_2295 (I40522,I40814,I40715);
not I_2296 (I40921,I40797);
nand I_2297 (I40938,I40715,I40921);
not I_2298 (I40516,I40938);
nor I_2299 (I40519,I40579,I40938);
nor I_2300 (I40531,I40921,I40579);
nand I_2301 (I40997,I40698,I40797);
nor I_2302 (I40513,I40596,I40997);
not I_2303 (I41055,I1869);
or I_2304 (I41072,I163192,I163171);
nand I_2305 (I41089,I163180,I163189);
not I_2306 (I41106,I41089);
nand I_2307 (I41123,I41106,I41072);
not I_2308 (I41140,I41123);
nand I_2309 (I41157,I163186,I163171);
and I_2310 (I41174,I41157,I163177);
DFFARX1 I_2311 (I41174,I1862,I41055,I41200,);
not I_2312 (I41208,I41200);
nor I_2313 (I41225,I163168,I163171);
nor I_2314 (I41242,I41200,I41225);
and I_2315 (I41259,I41200,I41225);
nor I_2316 (I41276,I41259,I41123);
DFFARX1 I_2317 (I41276,I1862,I41055,I41035,);
nand I_2318 (I41307,I163183,I163168);
nor I_2319 (I41324,I41307,I163174);
nand I_2320 (I41341,I41140,I41324);
not I_2321 (I41044,I41341);
nor I_2322 (I41047,I41242,I41341);
nor I_2323 (I41386,I41324,I41106);
nor I_2324 (I41038,I41208,I41386);
nor I_2325 (I41032,I41324,I41225);
not I_2326 (I41431,I41307);
nand I_2327 (I41448,I41225,I41431);
not I_2328 (I41026,I41448);
nor I_2329 (I41029,I41089,I41448);
nor I_2330 (I41041,I41431,I41089);
nand I_2331 (I41507,I41208,I41307);
nor I_2332 (I41023,I41106,I41507);
not I_2333 (I41565,I1869);
or I_2334 (I41582,I368562,I368562);
nand I_2335 (I41599,I368577,I368580);
not I_2336 (I41616,I41599);
nand I_2337 (I41633,I41616,I41582);
not I_2338 (I41650,I41633);
nand I_2339 (I41667,I368568,I368571);
and I_2340 (I41684,I41667,I368565);
DFFARX1 I_2341 (I41684,I1862,I41565,I41710,);
not I_2342 (I41718,I41710);
nor I_2343 (I41735,I368571,I368571);
nor I_2344 (I41752,I41710,I41735);
and I_2345 (I41769,I41710,I41735);
nor I_2346 (I41786,I41769,I41633);
DFFARX1 I_2347 (I41786,I1862,I41565,I41545,);
nand I_2348 (I41817,I368574,I368568);
nor I_2349 (I41834,I41817,I368565);
nand I_2350 (I41851,I41650,I41834);
not I_2351 (I41554,I41851);
nor I_2352 (I41557,I41752,I41851);
nor I_2353 (I41896,I41834,I41616);
nor I_2354 (I41548,I41718,I41896);
nor I_2355 (I41542,I41834,I41735);
not I_2356 (I41941,I41817);
nand I_2357 (I41958,I41735,I41941);
not I_2358 (I41536,I41958);
nor I_2359 (I41539,I41599,I41958);
nor I_2360 (I41551,I41941,I41599);
nand I_2361 (I42017,I41718,I41817);
nor I_2362 (I41533,I41616,I42017);
not I_2363 (I42075,I1869);
or I_2364 (I42092,I329434,I329428);
nand I_2365 (I42109,I329437,I329440);
not I_2366 (I42126,I42109);
nand I_2367 (I42143,I42126,I42092);
not I_2368 (I42160,I42143);
nand I_2369 (I42177,I329431,I329434);
and I_2370 (I42194,I42177,I329428);
DFFARX1 I_2371 (I42194,I1862,I42075,I42220,);
not I_2372 (I42228,I42220);
nor I_2373 (I42245,I329446,I329434);
nor I_2374 (I42262,I42220,I42245);
and I_2375 (I42279,I42220,I42245);
nor I_2376 (I42296,I42279,I42143);
DFFARX1 I_2377 (I42296,I1862,I42075,I42055,);
nand I_2378 (I42327,I329443,I329431);
nor I_2379 (I42344,I42327,I329449);
nand I_2380 (I42361,I42160,I42344);
not I_2381 (I42064,I42361);
nor I_2382 (I42067,I42262,I42361);
nor I_2383 (I42406,I42344,I42126);
nor I_2384 (I42058,I42228,I42406);
nor I_2385 (I42052,I42344,I42245);
not I_2386 (I42451,I42327);
nand I_2387 (I42468,I42245,I42451);
not I_2388 (I42046,I42468);
nor I_2389 (I42049,I42109,I42468);
nor I_2390 (I42061,I42451,I42109);
nand I_2391 (I42527,I42228,I42327);
nor I_2392 (I42043,I42126,I42527);
not I_2393 (I42585,I1869);
or I_2394 (I42602,I186380,I186359);
nand I_2395 (I42619,I186368,I186377);
not I_2396 (I42636,I42619);
nand I_2397 (I42653,I42636,I42602);
not I_2398 (I42670,I42653);
nand I_2399 (I42687,I186374,I186359);
and I_2400 (I42704,I42687,I186365);
DFFARX1 I_2401 (I42704,I1862,I42585,I42730,);
not I_2402 (I42738,I42730);
nor I_2403 (I42755,I186356,I186359);
nor I_2404 (I42772,I42730,I42755);
and I_2405 (I42789,I42730,I42755);
nor I_2406 (I42806,I42789,I42653);
DFFARX1 I_2407 (I42806,I1862,I42585,I42565,);
nand I_2408 (I42837,I186371,I186356);
nor I_2409 (I42854,I42837,I186362);
nand I_2410 (I42871,I42670,I42854);
not I_2411 (I42574,I42871);
nor I_2412 (I42577,I42772,I42871);
nor I_2413 (I42916,I42854,I42636);
nor I_2414 (I42568,I42738,I42916);
nor I_2415 (I42562,I42854,I42755);
not I_2416 (I42961,I42837);
nand I_2417 (I42978,I42755,I42961);
not I_2418 (I42556,I42978);
nor I_2419 (I42559,I42619,I42978);
nor I_2420 (I42571,I42961,I42619);
nand I_2421 (I43037,I42738,I42837);
nor I_2422 (I42553,I42636,I43037);
not I_2423 (I43095,I1869);
or I_2424 (I43112,I13466,I13466);
nand I_2425 (I43129,I13469,I13472);
not I_2426 (I43146,I43129);
nand I_2427 (I43163,I43146,I43112);
not I_2428 (I43180,I43163);
nand I_2429 (I43197,I13481,I13487);
and I_2430 (I43214,I43197,I13475);
DFFARX1 I_2431 (I43214,I1862,I43095,I43240,);
not I_2432 (I43248,I43240);
nor I_2433 (I43265,I13472,I13487);
nor I_2434 (I43282,I43240,I43265);
and I_2435 (I43299,I43240,I43265);
nor I_2436 (I43316,I43299,I43163);
DFFARX1 I_2437 (I43316,I1862,I43095,I43075,);
nand I_2438 (I43347,I13469,I13478);
nor I_2439 (I43364,I43347,I13484);
nand I_2440 (I43381,I43180,I43364);
not I_2441 (I43084,I43381);
nor I_2442 (I43087,I43282,I43381);
nor I_2443 (I43426,I43364,I43146);
nor I_2444 (I43078,I43248,I43426);
nor I_2445 (I43072,I43364,I43265);
not I_2446 (I43471,I43347);
nand I_2447 (I43488,I43265,I43471);
not I_2448 (I43066,I43488);
nor I_2449 (I43069,I43129,I43488);
nor I_2450 (I43081,I43471,I43129);
nand I_2451 (I43547,I43248,I43347);
nor I_2452 (I43063,I43146,I43547);
not I_2453 (I43605,I1869);
or I_2454 (I43622,I248188,I248191);
nand I_2455 (I43639,I248197,I248185);
not I_2456 (I43656,I43639);
nand I_2457 (I43673,I43656,I43622);
not I_2458 (I43690,I43673);
nand I_2459 (I43707,I248203,I248206);
and I_2460 (I43724,I43707,I248200);
DFFARX1 I_2461 (I43724,I1862,I43605,I43750,);
not I_2462 (I43758,I43750);
nor I_2463 (I43775,I248188,I248206);
nor I_2464 (I43792,I43750,I43775);
and I_2465 (I43809,I43750,I43775);
nor I_2466 (I43826,I43809,I43673);
DFFARX1 I_2467 (I43826,I1862,I43605,I43585,);
nand I_2468 (I43857,I248191,I248194);
nor I_2469 (I43874,I43857,I248185);
nand I_2470 (I43891,I43690,I43874);
not I_2471 (I43594,I43891);
nor I_2472 (I43597,I43792,I43891);
nor I_2473 (I43936,I43874,I43656);
nor I_2474 (I43588,I43758,I43936);
nor I_2475 (I43582,I43874,I43775);
not I_2476 (I43981,I43857);
nand I_2477 (I43998,I43775,I43981);
not I_2478 (I43576,I43998);
nor I_2479 (I43579,I43639,I43998);
nor I_2480 (I43591,I43981,I43639);
nand I_2481 (I44057,I43758,I43857);
nor I_2482 (I43573,I43656,I44057);
not I_2483 (I44115,I1869);
or I_2484 (I44132,I299919,I299916);
nand I_2485 (I44149,I299922,I299934);
not I_2486 (I44166,I44149);
nand I_2487 (I44183,I44166,I44132);
not I_2488 (I44200,I44183);
nand I_2489 (I44217,I299919,I299925);
and I_2490 (I44234,I44217,I299931);
DFFARX1 I_2491 (I44234,I1862,I44115,I44260,);
not I_2492 (I44268,I44260);
nor I_2493 (I44285,I299937,I299925);
nor I_2494 (I44302,I44260,I44285);
and I_2495 (I44319,I44260,I44285);
nor I_2496 (I44336,I44319,I44183);
DFFARX1 I_2497 (I44336,I1862,I44115,I44095,);
nand I_2498 (I44367,I299928,I299922);
nor I_2499 (I44384,I44367,I299916);
nand I_2500 (I44401,I44200,I44384);
not I_2501 (I44104,I44401);
nor I_2502 (I44107,I44302,I44401);
nor I_2503 (I44446,I44384,I44166);
nor I_2504 (I44098,I44268,I44446);
nor I_2505 (I44092,I44384,I44285);
not I_2506 (I44491,I44367);
nand I_2507 (I44508,I44285,I44491);
not I_2508 (I44086,I44508);
nor I_2509 (I44089,I44149,I44508);
nor I_2510 (I44101,I44491,I44149);
nand I_2511 (I44567,I44268,I44367);
nor I_2512 (I44083,I44166,I44567);
not I_2513 (I44625,I1869);
or I_2514 (I44642,I206776,I206779);
nand I_2515 (I44659,I206785,I206773);
not I_2516 (I44676,I44659);
nand I_2517 (I44693,I44676,I44642);
not I_2518 (I44710,I44693);
nand I_2519 (I44727,I206791,I206794);
and I_2520 (I44744,I44727,I206788);
DFFARX1 I_2521 (I44744,I1862,I44625,I44770,);
not I_2522 (I44778,I44770);
nor I_2523 (I44795,I206776,I206794);
nor I_2524 (I44812,I44770,I44795);
and I_2525 (I44829,I44770,I44795);
nor I_2526 (I44846,I44829,I44693);
DFFARX1 I_2527 (I44846,I1862,I44625,I44605,);
nand I_2528 (I44877,I206779,I206782);
nor I_2529 (I44894,I44877,I206773);
nand I_2530 (I44911,I44710,I44894);
not I_2531 (I44614,I44911);
nor I_2532 (I44617,I44812,I44911);
nor I_2533 (I44956,I44894,I44676);
nor I_2534 (I44608,I44778,I44956);
nor I_2535 (I44602,I44894,I44795);
not I_2536 (I45001,I44877);
nand I_2537 (I45018,I44795,I45001);
not I_2538 (I44596,I45018);
nor I_2539 (I44599,I44659,I45018);
nor I_2540 (I44611,I45001,I44659);
nand I_2541 (I45077,I44778,I44877);
nor I_2542 (I44593,I44676,I45077);
not I_2543 (I45135,I1869);
or I_2544 (I45152,I201064,I201067);
nand I_2545 (I45169,I201073,I201061);
not I_2546 (I45186,I45169);
nand I_2547 (I45203,I45186,I45152);
not I_2548 (I45220,I45203);
nand I_2549 (I45237,I201079,I201082);
and I_2550 (I45254,I45237,I201076);
DFFARX1 I_2551 (I45254,I1862,I45135,I45280,);
not I_2552 (I45288,I45280);
nor I_2553 (I45305,I201064,I201082);
nor I_2554 (I45322,I45280,I45305);
and I_2555 (I45339,I45280,I45305);
nor I_2556 (I45356,I45339,I45203);
DFFARX1 I_2557 (I45356,I1862,I45135,I45115,);
nand I_2558 (I45387,I201067,I201070);
nor I_2559 (I45404,I45387,I201061);
nand I_2560 (I45421,I45220,I45404);
not I_2561 (I45124,I45421);
nor I_2562 (I45127,I45322,I45421);
nor I_2563 (I45466,I45404,I45186);
nor I_2564 (I45118,I45288,I45466);
nor I_2565 (I45112,I45404,I45305);
not I_2566 (I45511,I45387);
nand I_2567 (I45528,I45305,I45511);
not I_2568 (I45106,I45528);
nor I_2569 (I45109,I45169,I45528);
nor I_2570 (I45121,I45511,I45169);
nand I_2571 (I45587,I45288,I45387);
nor I_2572 (I45103,I45186,I45587);
not I_2573 (I45645,I1869);
or I_2574 (I45662,I325745,I325739);
nand I_2575 (I45679,I325748,I325751);
not I_2576 (I45696,I45679);
nand I_2577 (I45713,I45696,I45662);
not I_2578 (I45730,I45713);
nand I_2579 (I45747,I325742,I325745);
and I_2580 (I45764,I45747,I325739);
DFFARX1 I_2581 (I45764,I1862,I45645,I45790,);
not I_2582 (I45798,I45790);
nor I_2583 (I45815,I325757,I325745);
nor I_2584 (I45832,I45790,I45815);
and I_2585 (I45849,I45790,I45815);
nor I_2586 (I45866,I45849,I45713);
DFFARX1 I_2587 (I45866,I1862,I45645,I45625,);
nand I_2588 (I45897,I325754,I325742);
nor I_2589 (I45914,I45897,I325760);
nand I_2590 (I45931,I45730,I45914);
not I_2591 (I45634,I45931);
nor I_2592 (I45637,I45832,I45931);
nor I_2593 (I45976,I45914,I45696);
nor I_2594 (I45628,I45798,I45976);
nor I_2595 (I45622,I45914,I45815);
not I_2596 (I46021,I45897);
nand I_2597 (I46038,I45815,I46021);
not I_2598 (I45616,I46038);
nor I_2599 (I45619,I45679,I46038);
nor I_2600 (I45631,I46021,I45679);
nand I_2601 (I46097,I45798,I45897);
nor I_2602 (I45613,I45696,I46097);
not I_2603 (I46155,I1869);
or I_2604 (I46172,I256280,I256283);
nand I_2605 (I46189,I256289,I256277);
not I_2606 (I46206,I46189);
nand I_2607 (I46223,I46206,I46172);
not I_2608 (I46240,I46223);
nand I_2609 (I46257,I256295,I256298);
and I_2610 (I46274,I46257,I256292);
DFFARX1 I_2611 (I46274,I1862,I46155,I46300,);
not I_2612 (I46308,I46300);
nor I_2613 (I46325,I256280,I256298);
nor I_2614 (I46342,I46300,I46325);
and I_2615 (I46359,I46300,I46325);
nor I_2616 (I46376,I46359,I46223);
DFFARX1 I_2617 (I46376,I1862,I46155,I46135,);
nand I_2618 (I46407,I256283,I256286);
nor I_2619 (I46424,I46407,I256277);
nand I_2620 (I46441,I46240,I46424);
not I_2621 (I46144,I46441);
nor I_2622 (I46147,I46342,I46441);
nor I_2623 (I46486,I46424,I46206);
nor I_2624 (I46138,I46308,I46486);
nor I_2625 (I46132,I46424,I46325);
not I_2626 (I46531,I46407);
nand I_2627 (I46548,I46325,I46531);
not I_2628 (I46126,I46548);
nor I_2629 (I46129,I46189,I46548);
nor I_2630 (I46141,I46531,I46189);
nand I_2631 (I46607,I46308,I46407);
nor I_2632 (I46123,I46206,I46607);
not I_2633 (I46665,I1869);
or I_2634 (I46682,I383590,I383590);
nand I_2635 (I46699,I383605,I383608);
not I_2636 (I46716,I46699);
nand I_2637 (I46733,I46716,I46682);
not I_2638 (I46750,I46733);
nand I_2639 (I46767,I383596,I383599);
and I_2640 (I46784,I46767,I383593);
DFFARX1 I_2641 (I46784,I1862,I46665,I46810,);
not I_2642 (I46818,I46810);
nor I_2643 (I46835,I383599,I383599);
nor I_2644 (I46852,I46810,I46835);
and I_2645 (I46869,I46810,I46835);
nor I_2646 (I46886,I46869,I46733);
DFFARX1 I_2647 (I46886,I1862,I46665,I46645,);
nand I_2648 (I46917,I383602,I383596);
nor I_2649 (I46934,I46917,I383593);
nand I_2650 (I46951,I46750,I46934);
not I_2651 (I46654,I46951);
nor I_2652 (I46657,I46852,I46951);
nor I_2653 (I46996,I46934,I46716);
nor I_2654 (I46648,I46818,I46996);
nor I_2655 (I46642,I46934,I46835);
not I_2656 (I47041,I46917);
nand I_2657 (I47058,I46835,I47041);
not I_2658 (I46636,I47058);
nor I_2659 (I46639,I46699,I47058);
nor I_2660 (I46651,I47041,I46699);
nand I_2661 (I47117,I46818,I46917);
nor I_2662 (I46633,I46716,I47117);
not I_2663 (I47175,I1869);
or I_2664 (I47192,I208204,I208207);
nand I_2665 (I47209,I208213,I208201);
not I_2666 (I47226,I47209);
nand I_2667 (I47243,I47226,I47192);
not I_2668 (I47260,I47243);
nand I_2669 (I47277,I208219,I208222);
and I_2670 (I47294,I47277,I208216);
DFFARX1 I_2671 (I47294,I1862,I47175,I47320,);
not I_2672 (I47328,I47320);
nor I_2673 (I47345,I208204,I208222);
nor I_2674 (I47362,I47320,I47345);
and I_2675 (I47379,I47320,I47345);
nor I_2676 (I47396,I47379,I47243);
DFFARX1 I_2677 (I47396,I1862,I47175,I47155,);
nand I_2678 (I47427,I208207,I208210);
nor I_2679 (I47444,I47427,I208201);
nand I_2680 (I47461,I47260,I47444);
not I_2681 (I47164,I47461);
nor I_2682 (I47167,I47362,I47461);
nor I_2683 (I47506,I47444,I47226);
nor I_2684 (I47158,I47328,I47506);
nor I_2685 (I47152,I47444,I47345);
not I_2686 (I47551,I47427);
nand I_2687 (I47568,I47345,I47551);
not I_2688 (I47146,I47568);
nor I_2689 (I47149,I47209,I47568);
nor I_2690 (I47161,I47551,I47209);
nand I_2691 (I47627,I47328,I47427);
nor I_2692 (I47143,I47226,I47627);
not I_2693 (I47685,I1869);
or I_2694 (I47702,I268656,I268659);
nand I_2695 (I47719,I268665,I268653);
not I_2696 (I47736,I47719);
nand I_2697 (I47753,I47736,I47702);
not I_2698 (I47770,I47753);
nand I_2699 (I47787,I268671,I268674);
and I_2700 (I47804,I47787,I268668);
DFFARX1 I_2701 (I47804,I1862,I47685,I47830,);
not I_2702 (I47838,I47830);
nor I_2703 (I47855,I268656,I268674);
nor I_2704 (I47872,I47830,I47855);
and I_2705 (I47889,I47830,I47855);
nor I_2706 (I47906,I47889,I47753);
DFFARX1 I_2707 (I47906,I1862,I47685,I47665,);
nand I_2708 (I47937,I268659,I268662);
nor I_2709 (I47954,I47937,I268653);
nand I_2710 (I47971,I47770,I47954);
not I_2711 (I47674,I47971);
nor I_2712 (I47677,I47872,I47971);
nor I_2713 (I48016,I47954,I47736);
nor I_2714 (I47668,I47838,I48016);
nor I_2715 (I47662,I47954,I47855);
not I_2716 (I48061,I47937);
nand I_2717 (I48078,I47855,I48061);
not I_2718 (I47656,I48078);
nor I_2719 (I47659,I47719,I48078);
nor I_2720 (I47671,I48061,I47719);
nand I_2721 (I48137,I47838,I47937);
nor I_2722 (I47653,I47736,I48137);
not I_2723 (I48195,I1869);
or I_2724 (I48212,I308354,I308348);
nand I_2725 (I48229,I308357,I308360);
not I_2726 (I48246,I48229);
nand I_2727 (I48263,I48246,I48212);
not I_2728 (I48280,I48263);
nand I_2729 (I48297,I308351,I308354);
and I_2730 (I48314,I48297,I308348);
DFFARX1 I_2731 (I48314,I1862,I48195,I48340,);
not I_2732 (I48348,I48340);
nor I_2733 (I48365,I308366,I308354);
nor I_2734 (I48382,I48340,I48365);
and I_2735 (I48399,I48340,I48365);
nor I_2736 (I48416,I48399,I48263);
DFFARX1 I_2737 (I48416,I1862,I48195,I48175,);
nand I_2738 (I48447,I308363,I308351);
nor I_2739 (I48464,I48447,I308369);
nand I_2740 (I48481,I48280,I48464);
not I_2741 (I48184,I48481);
nor I_2742 (I48187,I48382,I48481);
nor I_2743 (I48526,I48464,I48246);
nor I_2744 (I48178,I48348,I48526);
nor I_2745 (I48172,I48464,I48365);
not I_2746 (I48571,I48447);
nand I_2747 (I48588,I48365,I48571);
not I_2748 (I48166,I48588);
nor I_2749 (I48169,I48229,I48588);
nor I_2750 (I48181,I48571,I48229);
nand I_2751 (I48647,I48348,I48447);
nor I_2752 (I48163,I48246,I48647);
not I_2753 (I48705,I1869);
or I_2754 (I48722,I234860,I234863);
nand I_2755 (I48739,I234869,I234857);
not I_2756 (I48756,I48739);
nand I_2757 (I48773,I48756,I48722);
not I_2758 (I48790,I48773);
nand I_2759 (I48807,I234875,I234878);
and I_2760 (I48824,I48807,I234872);
DFFARX1 I_2761 (I48824,I1862,I48705,I48850,);
not I_2762 (I48858,I48850);
nor I_2763 (I48875,I234860,I234878);
nor I_2764 (I48892,I48850,I48875);
and I_2765 (I48909,I48850,I48875);
nor I_2766 (I48926,I48909,I48773);
DFFARX1 I_2767 (I48926,I1862,I48705,I48685,);
nand I_2768 (I48957,I234863,I234866);
nor I_2769 (I48974,I48957,I234857);
nand I_2770 (I48991,I48790,I48974);
not I_2771 (I48694,I48991);
nor I_2772 (I48697,I48892,I48991);
nor I_2773 (I49036,I48974,I48756);
nor I_2774 (I48688,I48858,I49036);
nor I_2775 (I48682,I48974,I48875);
not I_2776 (I49081,I48957);
nand I_2777 (I49098,I48875,I49081);
not I_2778 (I48676,I49098);
nor I_2779 (I48679,I48739,I49098);
nor I_2780 (I48691,I49081,I48739);
nand I_2781 (I49157,I48858,I48957);
nor I_2782 (I48673,I48756,I49157);
not I_2783 (I49215,I1869);
or I_2784 (I49232,I208680,I208683);
nand I_2785 (I49249,I208689,I208677);
not I_2786 (I49266,I49249);
nand I_2787 (I49283,I49266,I49232);
not I_2788 (I49300,I49283);
nand I_2789 (I49317,I208695,I208698);
and I_2790 (I49334,I49317,I208692);
DFFARX1 I_2791 (I49334,I1862,I49215,I49360,);
not I_2792 (I49368,I49360);
nor I_2793 (I49385,I208680,I208698);
nor I_2794 (I49402,I49360,I49385);
and I_2795 (I49419,I49360,I49385);
nor I_2796 (I49436,I49419,I49283);
DFFARX1 I_2797 (I49436,I1862,I49215,I49195,);
nand I_2798 (I49467,I208683,I208686);
nor I_2799 (I49484,I49467,I208677);
nand I_2800 (I49501,I49300,I49484);
not I_2801 (I49204,I49501);
nor I_2802 (I49207,I49402,I49501);
nor I_2803 (I49546,I49484,I49266);
nor I_2804 (I49198,I49368,I49546);
nor I_2805 (I49192,I49484,I49385);
not I_2806 (I49591,I49467);
nand I_2807 (I49608,I49385,I49591);
not I_2808 (I49186,I49608);
nor I_2809 (I49189,I49249,I49608);
nor I_2810 (I49201,I49591,I49249);
nand I_2811 (I49667,I49368,I49467);
nor I_2812 (I49183,I49266,I49667);
not I_2813 (I49725,I1869);
or I_2814 (I49742,I280556,I280559);
nand I_2815 (I49759,I280565,I280553);
not I_2816 (I49776,I49759);
nand I_2817 (I49793,I49776,I49742);
not I_2818 (I49810,I49793);
nand I_2819 (I49827,I280571,I280574);
and I_2820 (I49844,I49827,I280568);
DFFARX1 I_2821 (I49844,I1862,I49725,I49870,);
not I_2822 (I49878,I49870);
nor I_2823 (I49895,I280556,I280574);
nor I_2824 (I49912,I49870,I49895);
and I_2825 (I49929,I49870,I49895);
nor I_2826 (I49946,I49929,I49793);
DFFARX1 I_2827 (I49946,I1862,I49725,I49705,);
nand I_2828 (I49977,I280559,I280562);
nor I_2829 (I49994,I49977,I280553);
nand I_2830 (I50011,I49810,I49994);
not I_2831 (I49714,I50011);
nor I_2832 (I49717,I49912,I50011);
nor I_2833 (I50056,I49994,I49776);
nor I_2834 (I49708,I49878,I50056);
nor I_2835 (I49702,I49994,I49895);
not I_2836 (I50101,I49977);
nand I_2837 (I50118,I49895,I50101);
not I_2838 (I49696,I50118);
nor I_2839 (I49699,I49759,I50118);
nor I_2840 (I49711,I50101,I49759);
nand I_2841 (I50177,I49878,I49977);
nor I_2842 (I49693,I49776,I50177);
not I_2843 (I50235,I1869);
or I_2844 (I50252,I298865,I298862);
nand I_2845 (I50269,I298868,I298880);
not I_2846 (I50286,I50269);
nand I_2847 (I50303,I50286,I50252);
not I_2848 (I50320,I50303);
nand I_2849 (I50337,I298865,I298871);
and I_2850 (I50354,I50337,I298877);
DFFARX1 I_2851 (I50354,I1862,I50235,I50380,);
not I_2852 (I50388,I50380);
nor I_2853 (I50405,I298883,I298871);
nor I_2854 (I50422,I50380,I50405);
and I_2855 (I50439,I50380,I50405);
nor I_2856 (I50456,I50439,I50303);
DFFARX1 I_2857 (I50456,I1862,I50235,I50215,);
nand I_2858 (I50487,I298874,I298868);
nor I_2859 (I50504,I50487,I298862);
nand I_2860 (I50521,I50320,I50504);
not I_2861 (I50224,I50521);
nor I_2862 (I50227,I50422,I50521);
nor I_2863 (I50566,I50504,I50286);
nor I_2864 (I50218,I50388,I50566);
nor I_2865 (I50212,I50504,I50405);
not I_2866 (I50611,I50487);
nand I_2867 (I50628,I50405,I50611);
not I_2868 (I50206,I50628);
nor I_2869 (I50209,I50269,I50628);
nor I_2870 (I50221,I50611,I50269);
nand I_2871 (I50687,I50388,I50487);
nor I_2872 (I50203,I50286,I50687);
not I_2873 (I50745,I1869);
or I_2874 (I50762,I105493,I105487);
nand I_2875 (I50779,I105493,I105505);
not I_2876 (I50796,I50779);
nand I_2877 (I50813,I50796,I50762);
not I_2878 (I50830,I50813);
nand I_2879 (I50847,I105499,I105490);
and I_2880 (I50864,I50847,I105487);
DFFARX1 I_2881 (I50864,I1862,I50745,I50890,);
not I_2882 (I50898,I50890);
nor I_2883 (I50915,I105502,I105490);
nor I_2884 (I50932,I50890,I50915);
and I_2885 (I50949,I50890,I50915);
nor I_2886 (I50966,I50949,I50813);
DFFARX1 I_2887 (I50966,I1862,I50745,I50725,);
nand I_2888 (I50997,I105496,I105496);
nor I_2889 (I51014,I50997,I105490);
nand I_2890 (I51031,I50830,I51014);
not I_2891 (I50734,I51031);
nor I_2892 (I50737,I50932,I51031);
nor I_2893 (I51076,I51014,I50796);
nor I_2894 (I50728,I50898,I51076);
nor I_2895 (I50722,I51014,I50915);
not I_2896 (I51121,I50997);
nand I_2897 (I51138,I50915,I51121);
not I_2898 (I50716,I51138);
nor I_2899 (I50719,I50779,I51138);
nor I_2900 (I50731,I51121,I50779);
nand I_2901 (I51197,I50898,I50997);
nor I_2902 (I50713,I50796,I51197);
not I_2903 (I51255,I1869);
or I_2904 (I51272,I251520,I251523);
nand I_2905 (I51289,I251529,I251517);
not I_2906 (I51306,I51289);
nand I_2907 (I51323,I51306,I51272);
not I_2908 (I51340,I51323);
nand I_2909 (I51357,I251535,I251538);
and I_2910 (I51374,I51357,I251532);
DFFARX1 I_2911 (I51374,I1862,I51255,I51400,);
not I_2912 (I51408,I51400);
nor I_2913 (I51425,I251520,I251538);
nor I_2914 (I51442,I51400,I51425);
and I_2915 (I51459,I51400,I51425);
nor I_2916 (I51476,I51459,I51323);
DFFARX1 I_2917 (I51476,I1862,I51255,I51235,);
nand I_2918 (I51507,I251523,I251526);
nor I_2919 (I51524,I51507,I251517);
nand I_2920 (I51541,I51340,I51524);
not I_2921 (I51244,I51541);
nor I_2922 (I51247,I51442,I51541);
nor I_2923 (I51586,I51524,I51306);
nor I_2924 (I51238,I51408,I51586);
nor I_2925 (I51232,I51524,I51425);
not I_2926 (I51631,I51507);
nand I_2927 (I51648,I51425,I51631);
not I_2928 (I51226,I51648);
nor I_2929 (I51229,I51289,I51648);
nor I_2930 (I51241,I51631,I51289);
nand I_2931 (I51707,I51408,I51507);
nor I_2932 (I51223,I51306,I51707);
not I_2933 (I51765,I1869);
or I_2934 (I51782,I336812,I336806);
nand I_2935 (I51799,I336815,I336818);
not I_2936 (I51816,I51799);
nand I_2937 (I51833,I51816,I51782);
not I_2938 (I51850,I51833);
nand I_2939 (I51867,I336809,I336812);
and I_2940 (I51884,I51867,I336806);
DFFARX1 I_2941 (I51884,I1862,I51765,I51910,);
not I_2942 (I51918,I51910);
nor I_2943 (I51935,I336824,I336812);
nor I_2944 (I51952,I51910,I51935);
and I_2945 (I51969,I51910,I51935);
nor I_2946 (I51986,I51969,I51833);
DFFARX1 I_2947 (I51986,I1862,I51765,I51745,);
nand I_2948 (I52017,I336821,I336809);
nor I_2949 (I52034,I52017,I336827);
nand I_2950 (I52051,I51850,I52034);
not I_2951 (I51754,I52051);
nor I_2952 (I51757,I51952,I52051);
nor I_2953 (I52096,I52034,I51816);
nor I_2954 (I51748,I51918,I52096);
nor I_2955 (I51742,I52034,I51935);
not I_2956 (I52141,I52017);
nand I_2957 (I52158,I51935,I52141);
not I_2958 (I51736,I52158);
nor I_2959 (I51739,I51799,I52158);
nor I_2960 (I51751,I52141,I51799);
nand I_2961 (I52217,I51918,I52017);
nor I_2962 (I51733,I51816,I52217);
not I_2963 (I52275,I1869);
or I_2964 (I52292,I199555,I199534);
nand I_2965 (I52309,I199543,I199552);
not I_2966 (I52326,I52309);
nand I_2967 (I52343,I52326,I52292);
not I_2968 (I52360,I52343);
nand I_2969 (I52377,I199549,I199534);
and I_2970 (I52394,I52377,I199540);
DFFARX1 I_2971 (I52394,I1862,I52275,I52420,);
not I_2972 (I52428,I52420);
nor I_2973 (I52445,I199531,I199534);
nor I_2974 (I52462,I52420,I52445);
and I_2975 (I52479,I52420,I52445);
nor I_2976 (I52496,I52479,I52343);
DFFARX1 I_2977 (I52496,I1862,I52275,I52255,);
nand I_2978 (I52527,I199546,I199531);
nor I_2979 (I52544,I52527,I199537);
nand I_2980 (I52561,I52360,I52544);
not I_2981 (I52264,I52561);
nor I_2982 (I52267,I52462,I52561);
nor I_2983 (I52606,I52544,I52326);
nor I_2984 (I52258,I52428,I52606);
nor I_2985 (I52252,I52544,I52445);
not I_2986 (I52651,I52527);
nand I_2987 (I52668,I52445,I52651);
not I_2988 (I52246,I52668);
nor I_2989 (I52249,I52309,I52668);
nor I_2990 (I52261,I52651,I52309);
nand I_2991 (I52727,I52428,I52527);
nor I_2992 (I52243,I52326,I52727);
not I_2993 (I52785,I1869);
or I_2994 (I52802,I147909,I147888);
nand I_2995 (I52819,I147897,I147906);
not I_2996 (I52836,I52819);
nand I_2997 (I52853,I52836,I52802);
not I_2998 (I52870,I52853);
nand I_2999 (I52887,I147903,I147888);
and I_3000 (I52904,I52887,I147894);
DFFARX1 I_3001 (I52904,I1862,I52785,I52930,);
not I_3002 (I52938,I52930);
nor I_3003 (I52955,I147885,I147888);
nor I_3004 (I52972,I52930,I52955);
and I_3005 (I52989,I52930,I52955);
nor I_3006 (I53006,I52989,I52853);
DFFARX1 I_3007 (I53006,I1862,I52785,I52765,);
nand I_3008 (I53037,I147900,I147885);
nor I_3009 (I53054,I53037,I147891);
nand I_3010 (I53071,I52870,I53054);
not I_3011 (I52774,I53071);
nor I_3012 (I52777,I52972,I53071);
nor I_3013 (I53116,I53054,I52836);
nor I_3014 (I52768,I52938,I53116);
nor I_3015 (I52762,I53054,I52955);
not I_3016 (I53161,I53037);
nand I_3017 (I53178,I52955,I53161);
not I_3018 (I52756,I53178);
nor I_3019 (I52759,I52819,I53178);
nor I_3020 (I52771,I53161,I52819);
nand I_3021 (I53237,I52938,I53037);
nor I_3022 (I52753,I52836,I53237);
not I_3023 (I53295,I1869);
or I_3024 (I53312,I324691,I324685);
nand I_3025 (I53329,I324694,I324697);
not I_3026 (I53346,I53329);
nand I_3027 (I53363,I53346,I53312);
not I_3028 (I53380,I53363);
nand I_3029 (I53397,I324688,I324691);
and I_3030 (I53414,I53397,I324685);
DFFARX1 I_3031 (I53414,I1862,I53295,I53440,);
not I_3032 (I53448,I53440);
nor I_3033 (I53465,I324703,I324691);
nor I_3034 (I53482,I53440,I53465);
and I_3035 (I53499,I53440,I53465);
nor I_3036 (I53516,I53499,I53363);
DFFARX1 I_3037 (I53516,I1862,I53295,I53275,);
nand I_3038 (I53547,I324700,I324688);
nor I_3039 (I53564,I53547,I324706);
nand I_3040 (I53581,I53380,I53564);
not I_3041 (I53284,I53581);
nor I_3042 (I53287,I53482,I53581);
nor I_3043 (I53626,I53564,I53346);
nor I_3044 (I53278,I53448,I53626);
nor I_3045 (I53272,I53564,I53465);
not I_3046 (I53671,I53547);
nand I_3047 (I53688,I53465,I53671);
not I_3048 (I53266,I53688);
nor I_3049 (I53269,I53329,I53688);
nor I_3050 (I53281,I53671,I53329);
nand I_3051 (I53747,I53448,I53547);
nor I_3052 (I53263,I53346,I53747);
not I_3053 (I53805,I1869);
or I_3054 (I53822,I381380,I381380);
nand I_3055 (I53839,I381395,I381398);
not I_3056 (I53856,I53839);
nand I_3057 (I53873,I53856,I53822);
not I_3058 (I53890,I53873);
nand I_3059 (I53907,I381386,I381389);
and I_3060 (I53924,I53907,I381383);
DFFARX1 I_3061 (I53924,I1862,I53805,I53950,);
not I_3062 (I53958,I53950);
nor I_3063 (I53975,I381389,I381389);
nor I_3064 (I53992,I53950,I53975);
and I_3065 (I54009,I53950,I53975);
nor I_3066 (I54026,I54009,I53873);
DFFARX1 I_3067 (I54026,I1862,I53805,I53785,);
nand I_3068 (I54057,I381392,I381386);
nor I_3069 (I54074,I54057,I381383);
nand I_3070 (I54091,I53890,I54074);
not I_3071 (I53794,I54091);
nor I_3072 (I53797,I53992,I54091);
nor I_3073 (I54136,I54074,I53856);
nor I_3074 (I53788,I53958,I54136);
nor I_3075 (I53782,I54074,I53975);
not I_3076 (I54181,I54057);
nand I_3077 (I54198,I53975,I54181);
not I_3078 (I53776,I54198);
nor I_3079 (I53779,I53839,I54198);
nor I_3080 (I53791,I54181,I53839);
nand I_3081 (I54257,I53958,I54057);
nor I_3082 (I53773,I53856,I54257);
not I_3083 (I54315,I1869);
or I_3084 (I54332,I247712,I247715);
nand I_3085 (I54349,I247721,I247709);
not I_3086 (I54366,I54349);
nand I_3087 (I54383,I54366,I54332);
not I_3088 (I54400,I54383);
nand I_3089 (I54417,I247727,I247730);
and I_3090 (I54434,I54417,I247724);
DFFARX1 I_3091 (I54434,I1862,I54315,I54460,);
not I_3092 (I54468,I54460);
nor I_3093 (I54485,I247712,I247730);
nor I_3094 (I54502,I54460,I54485);
and I_3095 (I54519,I54460,I54485);
nor I_3096 (I54536,I54519,I54383);
DFFARX1 I_3097 (I54536,I1862,I54315,I54295,);
nand I_3098 (I54567,I247715,I247718);
nor I_3099 (I54584,I54567,I247709);
nand I_3100 (I54601,I54400,I54584);
not I_3101 (I54304,I54601);
nor I_3102 (I54307,I54502,I54601);
nor I_3103 (I54646,I54584,I54366);
nor I_3104 (I54298,I54468,I54646);
nor I_3105 (I54292,I54584,I54485);
not I_3106 (I54691,I54567);
nand I_3107 (I54708,I54485,I54691);
not I_3108 (I54286,I54708);
nor I_3109 (I54289,I54349,I54708);
nor I_3110 (I54301,I54691,I54349);
nand I_3111 (I54767,I54468,I54567);
nor I_3112 (I54283,I54366,I54767);
not I_3113 (I54825,I1869);
or I_3114 (I54842,I7142,I7142);
nand I_3115 (I54859,I7145,I7148);
not I_3116 (I54876,I54859);
nand I_3117 (I54893,I54876,I54842);
not I_3118 (I54910,I54893);
nand I_3119 (I54927,I7157,I7163);
and I_3120 (I54944,I54927,I7151);
DFFARX1 I_3121 (I54944,I1862,I54825,I54970,);
not I_3122 (I54978,I54970);
nor I_3123 (I54995,I7148,I7163);
nor I_3124 (I55012,I54970,I54995);
and I_3125 (I55029,I54970,I54995);
nor I_3126 (I55046,I55029,I54893);
DFFARX1 I_3127 (I55046,I1862,I54825,I54805,);
nand I_3128 (I55077,I7145,I7154);
nor I_3129 (I55094,I55077,I7160);
nand I_3130 (I55111,I54910,I55094);
not I_3131 (I54814,I55111);
nor I_3132 (I54817,I55012,I55111);
nor I_3133 (I55156,I55094,I54876);
nor I_3134 (I54808,I54978,I55156);
nor I_3135 (I54802,I55094,I54995);
not I_3136 (I55201,I55077);
nand I_3137 (I55218,I54995,I55201);
not I_3138 (I54796,I55218);
nor I_3139 (I54799,I54859,I55218);
nor I_3140 (I54811,I55201,I54859);
nand I_3141 (I55277,I54978,I55077);
nor I_3142 (I54793,I54876,I55277);
not I_3143 (I55335,I1869);
or I_3144 (I55352,I217248,I217251);
nand I_3145 (I55369,I217257,I217245);
not I_3146 (I55386,I55369);
nand I_3147 (I55403,I55386,I55352);
not I_3148 (I55420,I55403);
nand I_3149 (I55437,I217263,I217266);
and I_3150 (I55454,I55437,I217260);
DFFARX1 I_3151 (I55454,I1862,I55335,I55480,);
not I_3152 (I55488,I55480);
nor I_3153 (I55505,I217248,I217266);
nor I_3154 (I55522,I55480,I55505);
and I_3155 (I55539,I55480,I55505);
nor I_3156 (I55556,I55539,I55403);
DFFARX1 I_3157 (I55556,I1862,I55335,I55315,);
nand I_3158 (I55587,I217251,I217254);
nor I_3159 (I55604,I55587,I217245);
nand I_3160 (I55621,I55420,I55604);
not I_3161 (I55324,I55621);
nor I_3162 (I55327,I55522,I55621);
nor I_3163 (I55666,I55604,I55386);
nor I_3164 (I55318,I55488,I55666);
nor I_3165 (I55312,I55604,I55505);
not I_3166 (I55711,I55587);
nand I_3167 (I55728,I55505,I55711);
not I_3168 (I55306,I55728);
nor I_3169 (I55309,I55369,I55728);
nor I_3170 (I55321,I55711,I55369);
nand I_3171 (I55787,I55488,I55587);
nor I_3172 (I55303,I55386,I55787);
not I_3173 (I55845,I1869);
or I_3174 (I55862,I230576,I230579);
nand I_3175 (I55879,I230585,I230573);
not I_3176 (I55896,I55879);
nand I_3177 (I55913,I55896,I55862);
not I_3178 (I55930,I55913);
nand I_3179 (I55947,I230591,I230594);
and I_3180 (I55964,I55947,I230588);
DFFARX1 I_3181 (I55964,I1862,I55845,I55990,);
not I_3182 (I55998,I55990);
nor I_3183 (I56015,I230576,I230594);
nor I_3184 (I56032,I55990,I56015);
and I_3185 (I56049,I55990,I56015);
nor I_3186 (I56066,I56049,I55913);
DFFARX1 I_3187 (I56066,I1862,I55845,I55825,);
nand I_3188 (I56097,I230579,I230582);
nor I_3189 (I56114,I56097,I230573);
nand I_3190 (I56131,I55930,I56114);
not I_3191 (I55834,I56131);
nor I_3192 (I55837,I56032,I56131);
nor I_3193 (I56176,I56114,I55896);
nor I_3194 (I55828,I55998,I56176);
nor I_3195 (I55822,I56114,I56015);
not I_3196 (I56221,I56097);
nand I_3197 (I56238,I56015,I56221);
not I_3198 (I55816,I56238);
nor I_3199 (I55819,I55879,I56238);
nor I_3200 (I55831,I56221,I55879);
nand I_3201 (I56297,I55998,I56097);
nor I_3202 (I55813,I55896,I56297);
not I_3203 (I56355,I1869);
or I_3204 (I56372,I191123,I191102);
nand I_3205 (I56389,I191111,I191120);
not I_3206 (I56406,I56389);
nand I_3207 (I56423,I56406,I56372);
not I_3208 (I56440,I56423);
nand I_3209 (I56457,I191117,I191102);
and I_3210 (I56474,I56457,I191108);
DFFARX1 I_3211 (I56474,I1862,I56355,I56500,);
not I_3212 (I56508,I56500);
nor I_3213 (I56525,I191099,I191102);
nor I_3214 (I56542,I56500,I56525);
and I_3215 (I56559,I56500,I56525);
nor I_3216 (I56576,I56559,I56423);
DFFARX1 I_3217 (I56576,I1862,I56355,I56335,);
nand I_3218 (I56607,I191114,I191099);
nor I_3219 (I56624,I56607,I191105);
nand I_3220 (I56641,I56440,I56624);
not I_3221 (I56344,I56641);
nor I_3222 (I56347,I56542,I56641);
nor I_3223 (I56686,I56624,I56406);
nor I_3224 (I56338,I56508,I56686);
nor I_3225 (I56332,I56624,I56525);
not I_3226 (I56731,I56607);
nand I_3227 (I56748,I56525,I56731);
not I_3228 (I56326,I56748);
nor I_3229 (I56329,I56389,I56748);
nor I_3230 (I56341,I56731,I56389);
nand I_3231 (I56807,I56508,I56607);
nor I_3232 (I56323,I56406,I56807);
not I_3233 (I56865,I1869);
or I_3234 (I56882,I121559,I121538);
nand I_3235 (I56899,I121547,I121556);
not I_3236 (I56916,I56899);
nand I_3237 (I56933,I56916,I56882);
not I_3238 (I56950,I56933);
nand I_3239 (I56967,I121553,I121538);
and I_3240 (I56984,I56967,I121544);
DFFARX1 I_3241 (I56984,I1862,I56865,I57010,);
not I_3242 (I57018,I57010);
nor I_3243 (I57035,I121535,I121538);
nor I_3244 (I57052,I57010,I57035);
and I_3245 (I57069,I57010,I57035);
nor I_3246 (I57086,I57069,I56933);
DFFARX1 I_3247 (I57086,I1862,I56865,I56845,);
nand I_3248 (I57117,I121550,I121535);
nor I_3249 (I57134,I57117,I121541);
nand I_3250 (I57151,I56950,I57134);
not I_3251 (I56854,I57151);
nor I_3252 (I56857,I57052,I57151);
nor I_3253 (I57196,I57134,I56916);
nor I_3254 (I56848,I57018,I57196);
nor I_3255 (I56842,I57134,I57035);
not I_3256 (I57241,I57117);
nand I_3257 (I57258,I57035,I57241);
not I_3258 (I56836,I57258);
nor I_3259 (I56839,I56899,I57258);
nor I_3260 (I56851,I57241,I56899);
nand I_3261 (I57317,I57018,I57117);
nor I_3262 (I56833,I56916,I57317);
not I_3263 (I57375,I1869);
or I_3264 (I57392,I341028,I341022);
nand I_3265 (I57409,I341031,I341034);
not I_3266 (I57426,I57409);
nand I_3267 (I57443,I57426,I57392);
not I_3268 (I57460,I57443);
nand I_3269 (I57477,I341025,I341028);
and I_3270 (I57494,I57477,I341022);
DFFARX1 I_3271 (I57494,I1862,I57375,I57520,);
not I_3272 (I57528,I57520);
nor I_3273 (I57545,I341040,I341028);
nor I_3274 (I57562,I57520,I57545);
and I_3275 (I57579,I57520,I57545);
nor I_3276 (I57596,I57579,I57443);
DFFARX1 I_3277 (I57596,I1862,I57375,I57355,);
nand I_3278 (I57627,I341037,I341025);
nor I_3279 (I57644,I57627,I341043);
nand I_3280 (I57661,I57460,I57644);
not I_3281 (I57364,I57661);
nor I_3282 (I57367,I57562,I57661);
nor I_3283 (I57706,I57644,I57426);
nor I_3284 (I57358,I57528,I57706);
nor I_3285 (I57352,I57644,I57545);
not I_3286 (I57751,I57627);
nand I_3287 (I57768,I57545,I57751);
not I_3288 (I57346,I57768);
nor I_3289 (I57349,I57409,I57768);
nor I_3290 (I57361,I57751,I57409);
nand I_3291 (I57827,I57528,I57627);
nor I_3292 (I57343,I57426,I57827);
not I_3293 (I57885,I1869);
or I_3294 (I57902,I379170,I379170);
nand I_3295 (I57919,I379185,I379188);
not I_3296 (I57936,I57919);
nand I_3297 (I57953,I57936,I57902);
not I_3298 (I57970,I57953);
nand I_3299 (I57987,I379176,I379179);
and I_3300 (I58004,I57987,I379173);
DFFARX1 I_3301 (I58004,I1862,I57885,I58030,);
not I_3302 (I58038,I58030);
nor I_3303 (I58055,I379179,I379179);
nor I_3304 (I58072,I58030,I58055);
and I_3305 (I58089,I58030,I58055);
nor I_3306 (I58106,I58089,I57953);
DFFARX1 I_3307 (I58106,I1862,I57885,I57865,);
nand I_3308 (I58137,I379182,I379176);
nor I_3309 (I58154,I58137,I379173);
nand I_3310 (I58171,I57970,I58154);
not I_3311 (I57874,I58171);
nor I_3312 (I57877,I58072,I58171);
nor I_3313 (I58216,I58154,I57936);
nor I_3314 (I57868,I58038,I58216);
nor I_3315 (I57862,I58154,I58055);
not I_3316 (I58261,I58137);
nand I_3317 (I58278,I58055,I58261);
not I_3318 (I57856,I58278);
nor I_3319 (I57859,I57919,I58278);
nor I_3320 (I57871,I58261,I57919);
nand I_3321 (I58337,I58038,I58137);
nor I_3322 (I57853,I57936,I58337);
not I_3323 (I58395,I1869);
or I_3324 (I58412,I233908,I233911);
nand I_3325 (I58429,I233917,I233905);
not I_3326 (I58446,I58429);
nand I_3327 (I58463,I58446,I58412);
not I_3328 (I58480,I58463);
nand I_3329 (I58497,I233923,I233926);
and I_3330 (I58514,I58497,I233920);
DFFARX1 I_3331 (I58514,I1862,I58395,I58540,);
not I_3332 (I58548,I58540);
nor I_3333 (I58565,I233908,I233926);
nor I_3334 (I58582,I58540,I58565);
and I_3335 (I58599,I58540,I58565);
nor I_3336 (I58616,I58599,I58463);
DFFARX1 I_3337 (I58616,I1862,I58395,I58375,);
nand I_3338 (I58647,I233911,I233914);
nor I_3339 (I58664,I58647,I233905);
nand I_3340 (I58681,I58480,I58664);
not I_3341 (I58384,I58681);
nor I_3342 (I58387,I58582,I58681);
nor I_3343 (I58726,I58664,I58446);
nor I_3344 (I58378,I58548,I58726);
nor I_3345 (I58372,I58664,I58565);
not I_3346 (I58771,I58647);
nand I_3347 (I58788,I58565,I58771);
not I_3348 (I58366,I58788);
nor I_3349 (I58369,I58429,I58788);
nor I_3350 (I58381,I58771,I58429);
nand I_3351 (I58847,I58548,I58647);
nor I_3352 (I58363,I58446,I58847);
not I_3353 (I58905,I1869);
or I_3354 (I58922,I260564,I260567);
nand I_3355 (I58939,I260573,I260561);
not I_3356 (I58956,I58939);
nand I_3357 (I58973,I58956,I58922);
not I_3358 (I58990,I58973);
nand I_3359 (I59007,I260579,I260582);
and I_3360 (I59024,I59007,I260576);
DFFARX1 I_3361 (I59024,I1862,I58905,I59050,);
not I_3362 (I59058,I59050);
nor I_3363 (I59075,I260564,I260582);
nor I_3364 (I59092,I59050,I59075);
and I_3365 (I59109,I59050,I59075);
nor I_3366 (I59126,I59109,I58973);
DFFARX1 I_3367 (I59126,I1862,I58905,I58885,);
nand I_3368 (I59157,I260567,I260570);
nor I_3369 (I59174,I59157,I260561);
nand I_3370 (I59191,I58990,I59174);
not I_3371 (I58894,I59191);
nor I_3372 (I58897,I59092,I59191);
nor I_3373 (I59236,I59174,I58956);
nor I_3374 (I58888,I59058,I59236);
nor I_3375 (I58882,I59174,I59075);
not I_3376 (I59281,I59157);
nand I_3377 (I59298,I59075,I59281);
not I_3378 (I58876,I59298);
nor I_3379 (I58879,I58939,I59298);
nor I_3380 (I58891,I59281,I58939);
nand I_3381 (I59357,I59058,I59157);
nor I_3382 (I58873,I58956,I59357);
not I_3383 (I59415,I1869);
or I_3384 (I59432,I131045,I131024);
nand I_3385 (I59449,I131033,I131042);
not I_3386 (I59466,I59449);
nand I_3387 (I59483,I59466,I59432);
not I_3388 (I59500,I59483);
nand I_3389 (I59517,I131039,I131024);
and I_3390 (I59534,I59517,I131030);
DFFARX1 I_3391 (I59534,I1862,I59415,I59560,);
not I_3392 (I59568,I59560);
nor I_3393 (I59585,I131021,I131024);
nor I_3394 (I59602,I59560,I59585);
and I_3395 (I59619,I59560,I59585);
nor I_3396 (I59636,I59619,I59483);
DFFARX1 I_3397 (I59636,I1862,I59415,I59395,);
nand I_3398 (I59667,I131036,I131021);
nor I_3399 (I59684,I59667,I131027);
nand I_3400 (I59701,I59500,I59684);
not I_3401 (I59404,I59701);
nor I_3402 (I59407,I59602,I59701);
nor I_3403 (I59746,I59684,I59466);
nor I_3404 (I59398,I59568,I59746);
nor I_3405 (I59392,I59684,I59585);
not I_3406 (I59791,I59667);
nand I_3407 (I59808,I59585,I59791);
not I_3408 (I59386,I59808);
nor I_3409 (I59389,I59449,I59808);
nor I_3410 (I59401,I59791,I59449);
nand I_3411 (I59867,I59568,I59667);
nor I_3412 (I59383,I59466,I59867);
not I_3413 (I59925,I1869);
or I_3414 (I59942,I215820,I215823);
nand I_3415 (I59959,I215829,I215817);
not I_3416 (I59976,I59959);
nand I_3417 (I59993,I59976,I59942);
not I_3418 (I60010,I59993);
nand I_3419 (I60027,I215835,I215838);
and I_3420 (I60044,I60027,I215832);
DFFARX1 I_3421 (I60044,I1862,I59925,I60070,);
not I_3422 (I60078,I60070);
nor I_3423 (I60095,I215820,I215838);
nor I_3424 (I60112,I60070,I60095);
and I_3425 (I60129,I60070,I60095);
nor I_3426 (I60146,I60129,I59993);
DFFARX1 I_3427 (I60146,I1862,I59925,I59905,);
nand I_3428 (I60177,I215823,I215826);
nor I_3429 (I60194,I60177,I215817);
nand I_3430 (I60211,I60010,I60194);
not I_3431 (I59914,I60211);
nor I_3432 (I59917,I60112,I60211);
nor I_3433 (I60256,I60194,I59976);
nor I_3434 (I59908,I60078,I60256);
nor I_3435 (I59902,I60194,I60095);
not I_3436 (I60301,I60177);
nand I_3437 (I60318,I60095,I60301);
not I_3438 (I59896,I60318);
nor I_3439 (I59899,I59959,I60318);
nor I_3440 (I59911,I60301,I59959);
nand I_3441 (I60377,I60078,I60177);
nor I_3442 (I59893,I59976,I60377);
not I_3443 (I60435,I1869);
or I_3444 (I60452,I250568,I250571);
nand I_3445 (I60469,I250577,I250565);
not I_3446 (I60486,I60469);
nand I_3447 (I60503,I60486,I60452);
not I_3448 (I60520,I60503);
nand I_3449 (I60537,I250583,I250586);
and I_3450 (I60554,I60537,I250580);
DFFARX1 I_3451 (I60554,I1862,I60435,I60580,);
not I_3452 (I60588,I60580);
nor I_3453 (I60605,I250568,I250586);
nor I_3454 (I60622,I60580,I60605);
and I_3455 (I60639,I60580,I60605);
nor I_3456 (I60656,I60639,I60503);
DFFARX1 I_3457 (I60656,I1862,I60435,I60415,);
nand I_3458 (I60687,I250571,I250574);
nor I_3459 (I60704,I60687,I250565);
nand I_3460 (I60721,I60520,I60704);
not I_3461 (I60424,I60721);
nor I_3462 (I60427,I60622,I60721);
nor I_3463 (I60766,I60704,I60486);
nor I_3464 (I60418,I60588,I60766);
nor I_3465 (I60412,I60704,I60605);
not I_3466 (I60811,I60687);
nand I_3467 (I60828,I60605,I60811);
not I_3468 (I60406,I60828);
nor I_3469 (I60409,I60469,I60828);
nor I_3470 (I60421,I60811,I60469);
nand I_3471 (I60887,I60588,I60687);
nor I_3472 (I60403,I60486,I60887);
not I_3473 (I60945,I1869);
or I_3474 (I60962,I1047,I1839);
nand I_3475 (I60979,I679,I1575);
not I_3476 (I60996,I60979);
nand I_3477 (I61013,I60996,I60962);
not I_3478 (I61030,I61013);
nand I_3479 (I61047,I1455,I1279);
and I_3480 (I61064,I61047,I1247);
DFFARX1 I_3481 (I61064,I1862,I60945,I61090,);
not I_3482 (I61098,I61090);
nor I_3483 (I61115,I959,I1279);
nor I_3484 (I61132,I61090,I61115);
and I_3485 (I61149,I61090,I61115);
nor I_3486 (I61166,I61149,I61013);
DFFARX1 I_3487 (I61166,I1862,I60945,I60925,);
nand I_3488 (I61197,I775,I919);
nor I_3489 (I61214,I61197,I1359);
nand I_3490 (I61231,I61030,I61214);
not I_3491 (I60934,I61231);
nor I_3492 (I60937,I61132,I61231);
nor I_3493 (I61276,I61214,I60996);
nor I_3494 (I60928,I61098,I61276);
nor I_3495 (I60922,I61214,I61115);
not I_3496 (I61321,I61197);
nand I_3497 (I61338,I61115,I61321);
not I_3498 (I60916,I61338);
nor I_3499 (I60919,I60979,I61338);
nor I_3500 (I60931,I61321,I60979);
nand I_3501 (I61397,I61098,I61197);
nor I_3502 (I60913,I60996,I61397);
not I_3503 (I61455,I1869);
or I_3504 (I61472,I10304,I10304);
nand I_3505 (I61489,I10307,I10310);
not I_3506 (I61506,I61489);
nand I_3507 (I61523,I61506,I61472);
not I_3508 (I61540,I61523);
nand I_3509 (I61557,I10319,I10325);
and I_3510 (I61574,I61557,I10313);
DFFARX1 I_3511 (I61574,I1862,I61455,I61600,);
not I_3512 (I61608,I61600);
nor I_3513 (I61625,I10310,I10325);
nor I_3514 (I61642,I61600,I61625);
and I_3515 (I61659,I61600,I61625);
nor I_3516 (I61676,I61659,I61523);
DFFARX1 I_3517 (I61676,I1862,I61455,I61435,);
nand I_3518 (I61707,I10307,I10316);
nor I_3519 (I61724,I61707,I10322);
nand I_3520 (I61741,I61540,I61724);
not I_3521 (I61444,I61741);
nor I_3522 (I61447,I61642,I61741);
nor I_3523 (I61786,I61724,I61506);
nor I_3524 (I61438,I61608,I61786);
nor I_3525 (I61432,I61724,I61625);
not I_3526 (I61831,I61707);
nand I_3527 (I61848,I61625,I61831);
not I_3528 (I61426,I61848);
nor I_3529 (I61429,I61489,I61848);
nor I_3530 (I61441,I61831,I61489);
nand I_3531 (I61907,I61608,I61707);
nor I_3532 (I61423,I61506,I61907);
not I_3533 (I61965,I1869);
or I_3534 (I61982,I126302,I126281);
nand I_3535 (I61999,I126290,I126299);
not I_3536 (I62016,I61999);
nand I_3537 (I62033,I62016,I61982);
not I_3538 (I62050,I62033);
nand I_3539 (I62067,I126296,I126281);
and I_3540 (I62084,I62067,I126287);
DFFARX1 I_3541 (I62084,I1862,I61965,I62110,);
not I_3542 (I62118,I62110);
nor I_3543 (I62135,I126278,I126281);
nor I_3544 (I62152,I62110,I62135);
and I_3545 (I62169,I62110,I62135);
nor I_3546 (I62186,I62169,I62033);
DFFARX1 I_3547 (I62186,I1862,I61965,I61945,);
nand I_3548 (I62217,I126293,I126278);
nor I_3549 (I62234,I62217,I126284);
nand I_3550 (I62251,I62050,I62234);
not I_3551 (I61954,I62251);
nor I_3552 (I61957,I62152,I62251);
nor I_3553 (I62296,I62234,I62016);
nor I_3554 (I61948,I62118,I62296);
nor I_3555 (I61942,I62234,I62135);
not I_3556 (I62341,I62217);
nand I_3557 (I62358,I62135,I62341);
not I_3558 (I61936,I62358);
nor I_3559 (I61939,I61999,I62358);
nor I_3560 (I61951,I62341,I61999);
nand I_3561 (I62417,I62118,I62217);
nor I_3562 (I61933,I62016,I62417);
not I_3563 (I62475,I1869);
or I_3564 (I62492,I116101,I116095);
nand I_3565 (I62509,I116101,I116113);
not I_3566 (I62526,I62509);
nand I_3567 (I62543,I62526,I62492);
not I_3568 (I62560,I62543);
nand I_3569 (I62577,I116107,I116098);
and I_3570 (I62594,I62577,I116095);
DFFARX1 I_3571 (I62594,I1862,I62475,I62620,);
not I_3572 (I62628,I62620);
nor I_3573 (I62645,I116110,I116098);
nor I_3574 (I62662,I62620,I62645);
and I_3575 (I62679,I62620,I62645);
nor I_3576 (I62696,I62679,I62543);
DFFARX1 I_3577 (I62696,I1862,I62475,I62455,);
nand I_3578 (I62727,I116104,I116104);
nor I_3579 (I62744,I62727,I116098);
nand I_3580 (I62761,I62560,I62744);
not I_3581 (I62464,I62761);
nor I_3582 (I62467,I62662,I62761);
nor I_3583 (I62806,I62744,I62526);
nor I_3584 (I62458,I62628,I62806);
nor I_3585 (I62452,I62744,I62645);
not I_3586 (I62851,I62727);
nand I_3587 (I62868,I62645,I62851);
not I_3588 (I62446,I62868);
nor I_3589 (I62449,I62509,I62868);
nor I_3590 (I62461,I62851,I62509);
nand I_3591 (I62927,I62628,I62727);
nor I_3592 (I62443,I62526,I62927);
not I_3593 (I62985,I1869);
or I_3594 (I63002,I155814,I155793);
nand I_3595 (I63019,I155802,I155811);
not I_3596 (I63036,I63019);
nand I_3597 (I63053,I63036,I63002);
not I_3598 (I63070,I63053);
nand I_3599 (I63087,I155808,I155793);
and I_3600 (I63104,I63087,I155799);
DFFARX1 I_3601 (I63104,I1862,I62985,I63130,);
not I_3602 (I63138,I63130);
nor I_3603 (I63155,I155790,I155793);
nor I_3604 (I63172,I63130,I63155);
and I_3605 (I63189,I63130,I63155);
nor I_3606 (I63206,I63189,I63053);
DFFARX1 I_3607 (I63206,I1862,I62985,I62965,);
nand I_3608 (I63237,I155805,I155790);
nor I_3609 (I63254,I63237,I155796);
nand I_3610 (I63271,I63070,I63254);
not I_3611 (I62974,I63271);
nor I_3612 (I62977,I63172,I63271);
nor I_3613 (I63316,I63254,I63036);
nor I_3614 (I62968,I63138,I63316);
nor I_3615 (I62962,I63254,I63155);
not I_3616 (I63361,I63237);
nand I_3617 (I63378,I63155,I63361);
not I_3618 (I62956,I63378);
nor I_3619 (I62959,I63019,I63378);
nor I_3620 (I62971,I63361,I63019);
nand I_3621 (I63437,I63138,I63237);
nor I_3622 (I62953,I63036,I63437);
not I_3623 (I63495,I1869);
or I_3624 (I63512,I261516,I261519);
nand I_3625 (I63529,I261525,I261513);
not I_3626 (I63546,I63529);
nand I_3627 (I63563,I63546,I63512);
not I_3628 (I63580,I63563);
nand I_3629 (I63597,I261531,I261534);
and I_3630 (I63614,I63597,I261528);
DFFARX1 I_3631 (I63614,I1862,I63495,I63640,);
not I_3632 (I63648,I63640);
nor I_3633 (I63665,I261516,I261534);
nor I_3634 (I63682,I63640,I63665);
and I_3635 (I63699,I63640,I63665);
nor I_3636 (I63716,I63699,I63563);
DFFARX1 I_3637 (I63716,I1862,I63495,I63475,);
nand I_3638 (I63747,I261519,I261522);
nor I_3639 (I63764,I63747,I261513);
nand I_3640 (I63781,I63580,I63764);
not I_3641 (I63484,I63781);
nor I_3642 (I63487,I63682,I63781);
nor I_3643 (I63826,I63764,I63546);
nor I_3644 (I63478,I63648,I63826);
nor I_3645 (I63472,I63764,I63665);
not I_3646 (I63871,I63747);
nand I_3647 (I63888,I63665,I63871);
not I_3648 (I63466,I63888);
nor I_3649 (I63469,I63529,I63888);
nor I_3650 (I63481,I63871,I63529);
nand I_3651 (I63947,I63648,I63747);
nor I_3652 (I63463,I63546,I63947);
not I_3653 (I64005,I1869);
or I_3654 (I64022,I395966,I395966);
nand I_3655 (I64039,I395981,I395984);
not I_3656 (I64056,I64039);
nand I_3657 (I64073,I64056,I64022);
not I_3658 (I64090,I64073);
nand I_3659 (I64107,I395972,I395975);
and I_3660 (I64124,I64107,I395969);
DFFARX1 I_3661 (I64124,I1862,I64005,I64150,);
not I_3662 (I64158,I64150);
nor I_3663 (I64175,I395975,I395975);
nor I_3664 (I64192,I64150,I64175);
and I_3665 (I64209,I64150,I64175);
nor I_3666 (I64226,I64209,I64073);
DFFARX1 I_3667 (I64226,I1862,I64005,I63985,);
nand I_3668 (I64257,I395978,I395972);
nor I_3669 (I64274,I64257,I395969);
nand I_3670 (I64291,I64090,I64274);
not I_3671 (I63994,I64291);
nor I_3672 (I63997,I64192,I64291);
nor I_3673 (I64336,I64274,I64056);
nor I_3674 (I63988,I64158,I64336);
nor I_3675 (I63982,I64274,I64175);
not I_3676 (I64381,I64257);
nand I_3677 (I64398,I64175,I64381);
not I_3678 (I63976,I64398);
nor I_3679 (I63979,I64039,I64398);
nor I_3680 (I63991,I64381,I64039);
nand I_3681 (I64457,I64158,I64257);
nor I_3682 (I63973,I64056,I64457);
not I_3683 (I64515,I1869);
or I_3684 (I64532,I251996,I251999);
nand I_3685 (I64549,I252005,I251993);
not I_3686 (I64566,I64549);
nand I_3687 (I64583,I64566,I64532);
not I_3688 (I64600,I64583);
nand I_3689 (I64617,I252011,I252014);
and I_3690 (I64634,I64617,I252008);
DFFARX1 I_3691 (I64634,I1862,I64515,I64660,);
not I_3692 (I64668,I64660);
nor I_3693 (I64685,I251996,I252014);
nor I_3694 (I64702,I64660,I64685);
and I_3695 (I64719,I64660,I64685);
nor I_3696 (I64736,I64719,I64583);
DFFARX1 I_3697 (I64736,I1862,I64515,I64495,);
nand I_3698 (I64767,I251999,I252002);
nor I_3699 (I64784,I64767,I251993);
nand I_3700 (I64801,I64600,I64784);
not I_3701 (I64504,I64801);
nor I_3702 (I64507,I64702,I64801);
nor I_3703 (I64846,I64784,I64566);
nor I_3704 (I64498,I64668,I64846);
nor I_3705 (I64492,I64784,I64685);
not I_3706 (I64891,I64767);
nand I_3707 (I64908,I64685,I64891);
not I_3708 (I64486,I64908);
nor I_3709 (I64489,I64549,I64908);
nor I_3710 (I64501,I64891,I64549);
nand I_3711 (I64967,I64668,I64767);
nor I_3712 (I64483,I64566,I64967);
not I_3713 (I65025,I1869);
or I_3714 (I65042,I394640,I394640);
nand I_3715 (I65059,I394655,I394658);
not I_3716 (I65076,I65059);
nand I_3717 (I65093,I65076,I65042);
not I_3718 (I65110,I65093);
nand I_3719 (I65127,I394646,I394649);
and I_3720 (I65144,I65127,I394643);
DFFARX1 I_3721 (I65144,I1862,I65025,I65170,);
not I_3722 (I65178,I65170);
nor I_3723 (I65195,I394649,I394649);
nor I_3724 (I65212,I65170,I65195);
and I_3725 (I65229,I65170,I65195);
nor I_3726 (I65246,I65229,I65093);
DFFARX1 I_3727 (I65246,I1862,I65025,I65005,);
nand I_3728 (I65277,I394652,I394646);
nor I_3729 (I65294,I65277,I394643);
nand I_3730 (I65311,I65110,I65294);
not I_3731 (I65014,I65311);
nor I_3732 (I65017,I65212,I65311);
nor I_3733 (I65356,I65294,I65076);
nor I_3734 (I65008,I65178,I65356);
nor I_3735 (I65002,I65294,I65195);
not I_3736 (I65401,I65277);
nand I_3737 (I65418,I65195,I65401);
not I_3738 (I64996,I65418);
nor I_3739 (I64999,I65059,I65418);
nor I_3740 (I65011,I65401,I65059);
nand I_3741 (I65477,I65178,I65277);
nor I_3742 (I64993,I65076,I65477);
not I_3743 (I65535,I1869);
or I_3744 (I65552,I304138,I304132);
nand I_3745 (I65569,I304141,I304144);
not I_3746 (I65586,I65569);
nand I_3747 (I65603,I65586,I65552);
not I_3748 (I65620,I65603);
nand I_3749 (I65637,I304135,I304138);
and I_3750 (I65654,I65637,I304132);
DFFARX1 I_3751 (I65654,I1862,I65535,I65680,);
not I_3752 (I65688,I65680);
nor I_3753 (I65705,I304150,I304138);
nor I_3754 (I65722,I65680,I65705);
and I_3755 (I65739,I65680,I65705);
nor I_3756 (I65756,I65739,I65603);
DFFARX1 I_3757 (I65756,I1862,I65535,I65515,);
nand I_3758 (I65787,I304147,I304135);
nor I_3759 (I65804,I65787,I304153);
nand I_3760 (I65821,I65620,I65804);
not I_3761 (I65524,I65821);
nor I_3762 (I65527,I65722,I65821);
nor I_3763 (I65866,I65804,I65586);
nor I_3764 (I65518,I65688,I65866);
nor I_3765 (I65512,I65804,I65705);
not I_3766 (I65911,I65787);
nand I_3767 (I65928,I65705,I65911);
not I_3768 (I65506,I65928);
nor I_3769 (I65509,I65569,I65928);
nor I_3770 (I65521,I65911,I65569);
nand I_3771 (I65987,I65688,I65787);
nor I_3772 (I65503,I65586,I65987);
not I_3773 (I66045,I1869);
or I_3774 (I66062,I408342,I408342);
nand I_3775 (I66079,I408357,I408360);
not I_3776 (I66096,I66079);
nand I_3777 (I66113,I66096,I66062);
not I_3778 (I66130,I66113);
nand I_3779 (I66147,I408348,I408351);
and I_3780 (I66164,I66147,I408345);
DFFARX1 I_3781 (I66164,I1862,I66045,I66190,);
not I_3782 (I66198,I66190);
nor I_3783 (I66215,I408351,I408351);
nor I_3784 (I66232,I66190,I66215);
and I_3785 (I66249,I66190,I66215);
nor I_3786 (I66266,I66249,I66113);
DFFARX1 I_3787 (I66266,I1862,I66045,I66025,);
nand I_3788 (I66297,I408354,I408348);
nor I_3789 (I66314,I66297,I408345);
nand I_3790 (I66331,I66130,I66314);
not I_3791 (I66034,I66331);
nor I_3792 (I66037,I66232,I66331);
nor I_3793 (I66376,I66314,I66096);
nor I_3794 (I66028,I66198,I66376);
nor I_3795 (I66022,I66314,I66215);
not I_3796 (I66421,I66297);
nand I_3797 (I66438,I66215,I66421);
not I_3798 (I66016,I66438);
nor I_3799 (I66019,I66079,I66438);
nor I_3800 (I66031,I66421,I66079);
nand I_3801 (I66497,I66198,I66297);
nor I_3802 (I66013,I66096,I66497);
not I_3803 (I66555,I1869);
or I_3804 (I66572,I117343,I117322);
nand I_3805 (I66589,I117331,I117340);
not I_3806 (I66606,I66589);
nand I_3807 (I66623,I66606,I66572);
not I_3808 (I66640,I66623);
nand I_3809 (I66657,I117337,I117322);
and I_3810 (I66674,I66657,I117328);
DFFARX1 I_3811 (I66674,I1862,I66555,I66700,);
not I_3812 (I66708,I66700);
nor I_3813 (I66725,I117319,I117322);
nor I_3814 (I66742,I66700,I66725);
and I_3815 (I66759,I66700,I66725);
nor I_3816 (I66776,I66759,I66623);
DFFARX1 I_3817 (I66776,I1862,I66555,I66535,);
nand I_3818 (I66807,I117334,I117319);
nor I_3819 (I66824,I66807,I117325);
nand I_3820 (I66841,I66640,I66824);
not I_3821 (I66544,I66841);
nor I_3822 (I66547,I66742,I66841);
nor I_3823 (I66886,I66824,I66606);
nor I_3824 (I66538,I66708,I66886);
nor I_3825 (I66532,I66824,I66725);
not I_3826 (I66931,I66807);
nand I_3827 (I66948,I66725,I66931);
not I_3828 (I66526,I66948);
nor I_3829 (I66529,I66589,I66948);
nor I_3830 (I66541,I66931,I66589);
nand I_3831 (I67007,I66708,I66807);
nor I_3832 (I66523,I66606,I67007);
not I_3833 (I67065,I1869);
or I_3834 (I67082,I114877,I114871);
nand I_3835 (I67099,I114877,I114889);
not I_3836 (I67116,I67099);
nand I_3837 (I67133,I67116,I67082);
not I_3838 (I67150,I67133);
nand I_3839 (I67167,I114883,I114874);
and I_3840 (I67184,I67167,I114871);
DFFARX1 I_3841 (I67184,I1862,I67065,I67210,);
not I_3842 (I67218,I67210);
nor I_3843 (I67235,I114886,I114874);
nor I_3844 (I67252,I67210,I67235);
and I_3845 (I67269,I67210,I67235);
nor I_3846 (I67286,I67269,I67133);
DFFARX1 I_3847 (I67286,I1862,I67065,I67045,);
nand I_3848 (I67317,I114880,I114880);
nor I_3849 (I67334,I67317,I114874);
nand I_3850 (I67351,I67150,I67334);
not I_3851 (I67054,I67351);
nor I_3852 (I67057,I67252,I67351);
nor I_3853 (I67396,I67334,I67116);
nor I_3854 (I67048,I67218,I67396);
nor I_3855 (I67042,I67334,I67235);
not I_3856 (I67441,I67317);
nand I_3857 (I67458,I67235,I67441);
not I_3858 (I67036,I67458);
nor I_3859 (I67039,I67099,I67458);
nor I_3860 (I67051,I67441,I67099);
nand I_3861 (I67517,I67218,I67317);
nor I_3862 (I67033,I67116,I67517);
not I_3863 (I67575,I1869);
or I_3864 (I67592,I192177,I192156);
nand I_3865 (I67609,I192165,I192174);
not I_3866 (I67626,I67609);
nand I_3867 (I67643,I67626,I67592);
not I_3868 (I67660,I67643);
nand I_3869 (I67677,I192171,I192156);
and I_3870 (I67694,I67677,I192162);
DFFARX1 I_3871 (I67694,I1862,I67575,I67720,);
not I_3872 (I67728,I67720);
nor I_3873 (I67745,I192153,I192156);
nor I_3874 (I67762,I67720,I67745);
and I_3875 (I67779,I67720,I67745);
nor I_3876 (I67796,I67779,I67643);
DFFARX1 I_3877 (I67796,I1862,I67575,I67555,);
nand I_3878 (I67827,I192168,I192153);
nor I_3879 (I67844,I67827,I192159);
nand I_3880 (I67861,I67660,I67844);
not I_3881 (I67564,I67861);
nor I_3882 (I67567,I67762,I67861);
nor I_3883 (I67906,I67844,I67626);
nor I_3884 (I67558,I67728,I67906);
nor I_3885 (I67552,I67844,I67745);
not I_3886 (I67951,I67827);
nand I_3887 (I67968,I67745,I67951);
not I_3888 (I67546,I67968);
nor I_3889 (I67549,I67609,I67968);
nor I_3890 (I67561,I67951,I67609);
nand I_3891 (I68027,I67728,I67827);
nor I_3892 (I67543,I67626,I68027);
not I_3893 (I68085,I1869);
or I_3894 (I68102,I230100,I230103);
nand I_3895 (I68119,I230109,I230097);
not I_3896 (I68136,I68119);
nand I_3897 (I68153,I68136,I68102);
not I_3898 (I68170,I68153);
nand I_3899 (I68187,I230115,I230118);
and I_3900 (I68204,I68187,I230112);
DFFARX1 I_3901 (I68204,I1862,I68085,I68230,);
not I_3902 (I68238,I68230);
nor I_3903 (I68255,I230100,I230118);
nor I_3904 (I68272,I68230,I68255);
and I_3905 (I68289,I68230,I68255);
nor I_3906 (I68306,I68289,I68153);
DFFARX1 I_3907 (I68306,I1862,I68085,I68065,);
nand I_3908 (I68337,I230103,I230106);
nor I_3909 (I68354,I68337,I230097);
nand I_3910 (I68371,I68170,I68354);
not I_3911 (I68074,I68371);
nor I_3912 (I68077,I68272,I68371);
nor I_3913 (I68416,I68354,I68136);
nor I_3914 (I68068,I68238,I68416);
nor I_3915 (I68062,I68354,I68255);
not I_3916 (I68461,I68337);
nand I_3917 (I68478,I68255,I68461);
not I_3918 (I68056,I68478);
nor I_3919 (I68059,I68119,I68478);
nor I_3920 (I68071,I68461,I68119);
nand I_3921 (I68537,I68238,I68337);
nor I_3922 (I68053,I68136,I68537);
not I_3923 (I68595,I1869);
or I_3924 (I68612,I221532,I221535);
nand I_3925 (I68629,I221541,I221529);
not I_3926 (I68646,I68629);
nand I_3927 (I68663,I68646,I68612);
not I_3928 (I68680,I68663);
nand I_3929 (I68697,I221547,I221550);
and I_3930 (I68714,I68697,I221544);
DFFARX1 I_3931 (I68714,I1862,I68595,I68740,);
not I_3932 (I68748,I68740);
nor I_3933 (I68765,I221532,I221550);
nor I_3934 (I68782,I68740,I68765);
and I_3935 (I68799,I68740,I68765);
nor I_3936 (I68816,I68799,I68663);
DFFARX1 I_3937 (I68816,I1862,I68595,I68575,);
nand I_3938 (I68847,I221535,I221538);
nor I_3939 (I68864,I68847,I221529);
nand I_3940 (I68881,I68680,I68864);
not I_3941 (I68584,I68881);
nor I_3942 (I68587,I68782,I68881);
nor I_3943 (I68926,I68864,I68646);
nor I_3944 (I68578,I68748,I68926);
nor I_3945 (I68572,I68864,I68765);
not I_3946 (I68971,I68847);
nand I_3947 (I68988,I68765,I68971);
not I_3948 (I68566,I68988);
nor I_3949 (I68569,I68629,I68988);
nor I_3950 (I68581,I68971,I68629);
nand I_3951 (I69047,I68748,I68847);
nor I_3952 (I68563,I68646,I69047);
not I_3953 (I69105,I1869);
or I_3954 (I69122,I162665,I162644);
nand I_3955 (I69139,I162653,I162662);
not I_3956 (I69156,I69139);
nand I_3957 (I69173,I69156,I69122);
not I_3958 (I69190,I69173);
nand I_3959 (I69207,I162659,I162644);
and I_3960 (I69224,I69207,I162650);
DFFARX1 I_3961 (I69224,I1862,I69105,I69250,);
not I_3962 (I69258,I69250);
nor I_3963 (I69275,I162641,I162644);
nor I_3964 (I69292,I69250,I69275);
and I_3965 (I69309,I69250,I69275);
nor I_3966 (I69326,I69309,I69173);
DFFARX1 I_3967 (I69326,I1862,I69105,I69085,);
nand I_3968 (I69357,I162656,I162641);
nor I_3969 (I69374,I69357,I162647);
nand I_3970 (I69391,I69190,I69374);
not I_3971 (I69094,I69391);
nor I_3972 (I69097,I69292,I69391);
nor I_3973 (I69436,I69374,I69156);
nor I_3974 (I69088,I69258,I69436);
nor I_3975 (I69082,I69374,I69275);
not I_3976 (I69481,I69357);
nand I_3977 (I69498,I69275,I69481);
not I_3978 (I69076,I69498);
nor I_3979 (I69079,I69139,I69498);
nor I_3980 (I69091,I69481,I69139);
nand I_3981 (I69557,I69258,I69357);
nor I_3982 (I69073,I69156,I69557);
not I_3983 (I69615,I1869);
or I_3984 (I69632,I231052,I231055);
nand I_3985 (I69649,I231061,I231049);
not I_3986 (I69666,I69649);
nand I_3987 (I69683,I69666,I69632);
not I_3988 (I69700,I69683);
nand I_3989 (I69717,I231067,I231070);
and I_3990 (I69734,I69717,I231064);
DFFARX1 I_3991 (I69734,I1862,I69615,I69760,);
not I_3992 (I69768,I69760);
nor I_3993 (I69785,I231052,I231070);
nor I_3994 (I69802,I69760,I69785);
and I_3995 (I69819,I69760,I69785);
nor I_3996 (I69836,I69819,I69683);
DFFARX1 I_3997 (I69836,I1862,I69615,I69595,);
nand I_3998 (I69867,I231055,I231058);
nor I_3999 (I69884,I69867,I231049);
nand I_4000 (I69901,I69700,I69884);
not I_4001 (I69604,I69901);
nor I_4002 (I69607,I69802,I69901);
nor I_4003 (I69946,I69884,I69666);
nor I_4004 (I69598,I69768,I69946);
nor I_4005 (I69592,I69884,I69785);
not I_4006 (I69991,I69867);
nand I_4007 (I70008,I69785,I69991);
not I_4008 (I69586,I70008);
nor I_4009 (I69589,I69649,I70008);
nor I_4010 (I69601,I69991,I69649);
nand I_4011 (I70067,I69768,I69867);
nor I_4012 (I69583,I69666,I70067);
not I_4013 (I70125,I1869);
or I_4014 (I70142,I148436,I148415);
nand I_4015 (I70159,I148424,I148433);
not I_4016 (I70176,I70159);
nand I_4017 (I70193,I70176,I70142);
not I_4018 (I70210,I70193);
nand I_4019 (I70227,I148430,I148415);
and I_4020 (I70244,I70227,I148421);
DFFARX1 I_4021 (I70244,I1862,I70125,I70270,);
not I_4022 (I70278,I70270);
nor I_4023 (I70295,I148412,I148415);
nor I_4024 (I70312,I70270,I70295);
and I_4025 (I70329,I70270,I70295);
nor I_4026 (I70346,I70329,I70193);
DFFARX1 I_4027 (I70346,I1862,I70125,I70105,);
nand I_4028 (I70377,I148427,I148412);
nor I_4029 (I70394,I70377,I148418);
nand I_4030 (I70411,I70210,I70394);
not I_4031 (I70114,I70411);
nor I_4032 (I70117,I70312,I70411);
nor I_4033 (I70456,I70394,I70176);
nor I_4034 (I70108,I70278,I70456);
nor I_4035 (I70102,I70394,I70295);
not I_4036 (I70501,I70377);
nand I_4037 (I70518,I70295,I70501);
not I_4038 (I70096,I70518);
nor I_4039 (I70099,I70159,I70518);
nor I_4040 (I70111,I70501,I70159);
nand I_4041 (I70577,I70278,I70377);
nor I_4042 (I70093,I70176,I70577);
not I_4043 (I70635,I1869);
or I_4044 (I70652,I168989,I168968);
nand I_4045 (I70669,I168977,I168986);
not I_4046 (I70686,I70669);
nand I_4047 (I70703,I70686,I70652);
not I_4048 (I70720,I70703);
nand I_4049 (I70737,I168983,I168968);
and I_4050 (I70754,I70737,I168974);
DFFARX1 I_4051 (I70754,I1862,I70635,I70780,);
not I_4052 (I70788,I70780);
nor I_4053 (I70805,I168965,I168968);
nor I_4054 (I70822,I70780,I70805);
and I_4055 (I70839,I70780,I70805);
nor I_4056 (I70856,I70839,I70703);
DFFARX1 I_4057 (I70856,I1862,I70635,I70615,);
nand I_4058 (I70887,I168980,I168965);
nor I_4059 (I70904,I70887,I168971);
nand I_4060 (I70921,I70720,I70904);
not I_4061 (I70624,I70921);
nor I_4062 (I70627,I70822,I70921);
nor I_4063 (I70966,I70904,I70686);
nor I_4064 (I70618,I70788,I70966);
nor I_4065 (I70612,I70904,I70805);
not I_4066 (I71011,I70887);
nand I_4067 (I71028,I70805,I71011);
not I_4068 (I70606,I71028);
nor I_4069 (I70609,I70669,I71028);
nor I_4070 (I70621,I71011,I70669);
nand I_4071 (I71087,I70788,I70887);
nor I_4072 (I70603,I70686,I71087);
not I_4073 (I71145,I1869);
or I_4074 (I71162,I2926,I2926);
nand I_4075 (I71179,I2929,I2932);
not I_4076 (I71196,I71179);
nand I_4077 (I71213,I71196,I71162);
not I_4078 (I71230,I71213);
nand I_4079 (I71247,I2941,I2947);
and I_4080 (I71264,I71247,I2935);
DFFARX1 I_4081 (I71264,I1862,I71145,I71290,);
not I_4082 (I71298,I71290);
nor I_4083 (I71315,I2932,I2947);
nor I_4084 (I71332,I71290,I71315);
and I_4085 (I71349,I71290,I71315);
nor I_4086 (I71366,I71349,I71213);
DFFARX1 I_4087 (I71366,I1862,I71145,I71125,);
nand I_4088 (I71397,I2929,I2938);
nor I_4089 (I71414,I71397,I2944);
nand I_4090 (I71431,I71230,I71414);
not I_4091 (I71134,I71431);
nor I_4092 (I71137,I71332,I71431);
nor I_4093 (I71476,I71414,I71196);
nor I_4094 (I71128,I71298,I71476);
nor I_4095 (I71122,I71414,I71315);
not I_4096 (I71521,I71397);
nand I_4097 (I71538,I71315,I71521);
not I_4098 (I71116,I71538);
nor I_4099 (I71119,I71179,I71538);
nor I_4100 (I71131,I71521,I71179);
nand I_4101 (I71597,I71298,I71397);
nor I_4102 (I71113,I71196,I71597);
not I_4103 (I71655,I1869);
or I_4104 (I71672,I183218,I183197);
nand I_4105 (I71689,I183206,I183215);
not I_4106 (I71706,I71689);
nand I_4107 (I71723,I71706,I71672);
not I_4108 (I71740,I71723);
nand I_4109 (I71757,I183212,I183197);
and I_4110 (I71774,I71757,I183203);
DFFARX1 I_4111 (I71774,I1862,I71655,I71800,);
not I_4112 (I71808,I71800);
nor I_4113 (I71825,I183194,I183197);
nor I_4114 (I71842,I71800,I71825);
and I_4115 (I71859,I71800,I71825);
nor I_4116 (I71876,I71859,I71723);
DFFARX1 I_4117 (I71876,I1862,I71655,I71635,);
nand I_4118 (I71907,I183209,I183194);
nor I_4119 (I71924,I71907,I183200);
nand I_4120 (I71941,I71740,I71924);
not I_4121 (I71644,I71941);
nor I_4122 (I71647,I71842,I71941);
nor I_4123 (I71986,I71924,I71706);
nor I_4124 (I71638,I71808,I71986);
nor I_4125 (I71632,I71924,I71825);
not I_4126 (I72031,I71907);
nand I_4127 (I72048,I71825,I72031);
not I_4128 (I71626,I72048);
nor I_4129 (I71629,I71689,I72048);
nor I_4130 (I71641,I72031,I71689);
nand I_4131 (I72107,I71808,I71907);
nor I_4132 (I71623,I71706,I72107);
not I_4133 (I72165,I1869);
or I_4134 (I72182,I342609,I342603);
nand I_4135 (I72199,I342612,I342615);
not I_4136 (I72216,I72199);
nand I_4137 (I72233,I72216,I72182);
not I_4138 (I72250,I72233);
nand I_4139 (I72267,I342606,I342609);
and I_4140 (I72284,I72267,I342603);
DFFARX1 I_4141 (I72284,I1862,I72165,I72310,);
not I_4142 (I72318,I72310);
nor I_4143 (I72335,I342621,I342609);
nor I_4144 (I72352,I72310,I72335);
and I_4145 (I72369,I72310,I72335);
nor I_4146 (I72386,I72369,I72233);
DFFARX1 I_4147 (I72386,I1862,I72165,I72145,);
nand I_4148 (I72417,I342618,I342606);
nor I_4149 (I72434,I72417,I342624);
nand I_4150 (I72451,I72250,I72434);
not I_4151 (I72154,I72451);
nor I_4152 (I72157,I72352,I72451);
nor I_4153 (I72496,I72434,I72216);
nor I_4154 (I72148,I72318,I72496);
nor I_4155 (I72142,I72434,I72335);
not I_4156 (I72541,I72417);
nand I_4157 (I72558,I72335,I72541);
not I_4158 (I72136,I72558);
nor I_4159 (I72139,I72199,I72558);
nor I_4160 (I72151,I72541,I72199);
nand I_4161 (I72617,I72318,I72417);
nor I_4162 (I72133,I72216,I72617);
not I_4163 (I72675,I1869);
or I_4164 (I72692,I177948,I177927);
nand I_4165 (I72709,I177936,I177945);
not I_4166 (I72726,I72709);
nand I_4167 (I72743,I72726,I72692);
not I_4168 (I72760,I72743);
nand I_4169 (I72777,I177942,I177927);
and I_4170 (I72794,I72777,I177933);
DFFARX1 I_4171 (I72794,I1862,I72675,I72820,);
not I_4172 (I72828,I72820);
nor I_4173 (I72845,I177924,I177927);
nor I_4174 (I72862,I72820,I72845);
and I_4175 (I72879,I72820,I72845);
nor I_4176 (I72896,I72879,I72743);
DFFARX1 I_4177 (I72896,I1862,I72675,I72655,);
nand I_4178 (I72927,I177939,I177924);
nor I_4179 (I72944,I72927,I177930);
nand I_4180 (I72961,I72760,I72944);
not I_4181 (I72664,I72961);
nor I_4182 (I72667,I72862,I72961);
nor I_4183 (I73006,I72944,I72726);
nor I_4184 (I72658,I72828,I73006);
nor I_4185 (I72652,I72944,I72845);
not I_4186 (I73051,I72927);
nand I_4187 (I73068,I72845,I73051);
not I_4188 (I72646,I73068);
nor I_4189 (I72649,I72709,I73068);
nor I_4190 (I72661,I73051,I72709);
nand I_4191 (I73127,I72828,I72927);
nor I_4192 (I72643,I72726,I73127);
not I_4193 (I73185,I1869);
or I_4194 (I73202,I317840,I317834);
nand I_4195 (I73219,I317843,I317846);
not I_4196 (I73236,I73219);
nand I_4197 (I73253,I73236,I73202);
not I_4198 (I73270,I73253);
nand I_4199 (I73287,I317837,I317840);
and I_4200 (I73304,I73287,I317834);
DFFARX1 I_4201 (I73304,I1862,I73185,I73330,);
not I_4202 (I73338,I73330);
nor I_4203 (I73355,I317852,I317840);
nor I_4204 (I73372,I73330,I73355);
and I_4205 (I73389,I73330,I73355);
nor I_4206 (I73406,I73389,I73253);
DFFARX1 I_4207 (I73406,I1862,I73185,I73165,);
nand I_4208 (I73437,I317849,I317837);
nor I_4209 (I73454,I73437,I317855);
nand I_4210 (I73471,I73270,I73454);
not I_4211 (I73174,I73471);
nor I_4212 (I73177,I73372,I73471);
nor I_4213 (I73516,I73454,I73236);
nor I_4214 (I73168,I73338,I73516);
nor I_4215 (I73162,I73454,I73355);
not I_4216 (I73561,I73437);
nand I_4217 (I73578,I73355,I73561);
not I_4218 (I73156,I73578);
nor I_4219 (I73159,I73219,I73578);
nor I_4220 (I73171,I73561,I73219);
nand I_4221 (I73637,I73338,I73437);
nor I_4222 (I73153,I73236,I73637);
not I_4223 (I73695,I1869);
or I_4224 (I73712,I294649,I294646);
nand I_4225 (I73729,I294652,I294664);
not I_4226 (I73746,I73729);
nand I_4227 (I73763,I73746,I73712);
not I_4228 (I73780,I73763);
nand I_4229 (I73797,I294649,I294655);
and I_4230 (I73814,I73797,I294661);
DFFARX1 I_4231 (I73814,I1862,I73695,I73840,);
not I_4232 (I73848,I73840);
nor I_4233 (I73865,I294667,I294655);
nor I_4234 (I73882,I73840,I73865);
and I_4235 (I73899,I73840,I73865);
nor I_4236 (I73916,I73899,I73763);
DFFARX1 I_4237 (I73916,I1862,I73695,I73675,);
nand I_4238 (I73947,I294658,I294652);
nor I_4239 (I73964,I73947,I294646);
nand I_4240 (I73981,I73780,I73964);
not I_4241 (I73684,I73981);
nor I_4242 (I73687,I73882,I73981);
nor I_4243 (I74026,I73964,I73746);
nor I_4244 (I73678,I73848,I74026);
nor I_4245 (I73672,I73964,I73865);
not I_4246 (I74071,I73947);
nand I_4247 (I74088,I73865,I74071);
not I_4248 (I73666,I74088);
nor I_4249 (I73669,I73729,I74088);
nor I_4250 (I73681,I74071,I73729);
nand I_4251 (I74147,I73848,I73947);
nor I_4252 (I73663,I73746,I74147);
not I_4253 (I74205,I1869);
or I_4254 (I74222,I261040,I261043);
nand I_4255 (I74239,I261049,I261037);
not I_4256 (I74256,I74239);
nand I_4257 (I74273,I74256,I74222);
not I_4258 (I74290,I74273);
nand I_4259 (I74307,I261055,I261058);
and I_4260 (I74324,I74307,I261052);
DFFARX1 I_4261 (I74324,I1862,I74205,I74350,);
not I_4262 (I74358,I74350);
nor I_4263 (I74375,I261040,I261058);
nor I_4264 (I74392,I74350,I74375);
and I_4265 (I74409,I74350,I74375);
nor I_4266 (I74426,I74409,I74273);
DFFARX1 I_4267 (I74426,I1862,I74205,I74185,);
nand I_4268 (I74457,I261043,I261046);
nor I_4269 (I74474,I74457,I261037);
nand I_4270 (I74491,I74290,I74474);
not I_4271 (I74194,I74491);
nor I_4272 (I74197,I74392,I74491);
nor I_4273 (I74536,I74474,I74256);
nor I_4274 (I74188,I74358,I74536);
nor I_4275 (I74182,I74474,I74375);
not I_4276 (I74581,I74457);
nand I_4277 (I74598,I74375,I74581);
not I_4278 (I74176,I74598);
nor I_4279 (I74179,I74239,I74598);
nor I_4280 (I74191,I74581,I74239);
nand I_4281 (I74657,I74358,I74457);
nor I_4282 (I74173,I74256,I74657);
not I_4283 (I74715,I1869);
or I_4284 (I74732,I268180,I268183);
nand I_4285 (I74749,I268189,I268177);
not I_4286 (I74766,I74749);
nand I_4287 (I74783,I74766,I74732);
not I_4288 (I74800,I74783);
nand I_4289 (I74817,I268195,I268198);
and I_4290 (I74834,I74817,I268192);
DFFARX1 I_4291 (I74834,I1862,I74715,I74860,);
not I_4292 (I74868,I74860);
nor I_4293 (I74885,I268180,I268198);
nor I_4294 (I74902,I74860,I74885);
and I_4295 (I74919,I74860,I74885);
nor I_4296 (I74936,I74919,I74783);
DFFARX1 I_4297 (I74936,I1862,I74715,I74695,);
nand I_4298 (I74967,I268183,I268186);
nor I_4299 (I74984,I74967,I268177);
nand I_4300 (I75001,I74800,I74984);
not I_4301 (I74704,I75001);
nor I_4302 (I74707,I74902,I75001);
nor I_4303 (I75046,I74984,I74766);
nor I_4304 (I74698,I74868,I75046);
nor I_4305 (I74692,I74984,I74885);
not I_4306 (I75091,I74967);
nand I_4307 (I75108,I74885,I75091);
not I_4308 (I74686,I75108);
nor I_4309 (I74689,I74749,I75108);
nor I_4310 (I74701,I75091,I74749);
nand I_4311 (I75167,I74868,I74967);
nor I_4312 (I74683,I74766,I75167);
not I_4313 (I75225,I1869);
or I_4314 (I75242,I202968,I202971);
nand I_4315 (I75259,I202977,I202965);
not I_4316 (I75276,I75259);
nand I_4317 (I75293,I75276,I75242);
not I_4318 (I75310,I75293);
nand I_4319 (I75327,I202983,I202986);
and I_4320 (I75344,I75327,I202980);
DFFARX1 I_4321 (I75344,I1862,I75225,I75370,);
not I_4322 (I75378,I75370);
nor I_4323 (I75395,I202968,I202986);
nor I_4324 (I75412,I75370,I75395);
and I_4325 (I75429,I75370,I75395);
nor I_4326 (I75446,I75429,I75293);
DFFARX1 I_4327 (I75446,I1862,I75225,I75205,);
nand I_4328 (I75477,I202971,I202974);
nor I_4329 (I75494,I75477,I202965);
nand I_4330 (I75511,I75310,I75494);
not I_4331 (I75214,I75511);
nor I_4332 (I75217,I75412,I75511);
nor I_4333 (I75556,I75494,I75276);
nor I_4334 (I75208,I75378,I75556);
nor I_4335 (I75202,I75494,I75395);
not I_4336 (I75601,I75477);
nand I_4337 (I75618,I75395,I75601);
not I_4338 (I75196,I75618);
nor I_4339 (I75199,I75259,I75618);
nor I_4340 (I75211,I75601,I75259);
nand I_4341 (I75677,I75378,I75477);
nor I_4342 (I75193,I75276,I75677);
not I_4343 (I75735,I1869);
or I_4344 (I75752,I120505,I120484);
nand I_4345 (I75769,I120493,I120502);
not I_4346 (I75786,I75769);
nand I_4347 (I75803,I75786,I75752);
not I_4348 (I75820,I75803);
nand I_4349 (I75837,I120499,I120484);
and I_4350 (I75854,I75837,I120490);
DFFARX1 I_4351 (I75854,I1862,I75735,I75880,);
not I_4352 (I75888,I75880);
nor I_4353 (I75905,I120481,I120484);
nor I_4354 (I75922,I75880,I75905);
and I_4355 (I75939,I75880,I75905);
nor I_4356 (I75956,I75939,I75803);
DFFARX1 I_4357 (I75956,I1862,I75735,I75715,);
nand I_4358 (I75987,I120496,I120481);
nor I_4359 (I76004,I75987,I120487);
nand I_4360 (I76021,I75820,I76004);
not I_4361 (I75724,I76021);
nor I_4362 (I75727,I75922,I76021);
nor I_4363 (I76066,I76004,I75786);
nor I_4364 (I75718,I75888,I76066);
nor I_4365 (I75712,I76004,I75905);
not I_4366 (I76111,I75987);
nand I_4367 (I76128,I75905,I76111);
not I_4368 (I75706,I76128);
nor I_4369 (I75709,I75769,I76128);
nor I_4370 (I75721,I76111,I75769);
nand I_4371 (I76187,I75888,I75987);
nor I_4372 (I75703,I75786,I76187);
not I_4373 (I76245,I1869);
or I_4374 (I76262,I152652,I152631);
nand I_4375 (I76279,I152640,I152649);
not I_4376 (I76296,I76279);
nand I_4377 (I76313,I76296,I76262);
not I_4378 (I76330,I76313);
nand I_4379 (I76347,I152646,I152631);
and I_4380 (I76364,I76347,I152637);
DFFARX1 I_4381 (I76364,I1862,I76245,I76390,);
not I_4382 (I76398,I76390);
nor I_4383 (I76415,I152628,I152631);
nor I_4384 (I76432,I76390,I76415);
and I_4385 (I76449,I76390,I76415);
nor I_4386 (I76466,I76449,I76313);
DFFARX1 I_4387 (I76466,I1862,I76245,I76225,);
nand I_4388 (I76497,I152643,I152628);
nor I_4389 (I76514,I76497,I152634);
nand I_4390 (I76531,I76330,I76514);
not I_4391 (I76234,I76531);
nor I_4392 (I76237,I76432,I76531);
nor I_4393 (I76576,I76514,I76296);
nor I_4394 (I76228,I76398,I76576);
nor I_4395 (I76222,I76514,I76415);
not I_4396 (I76621,I76497);
nand I_4397 (I76638,I76415,I76621);
not I_4398 (I76216,I76638);
nor I_4399 (I76219,I76279,I76638);
nor I_4400 (I76231,I76621,I76279);
nand I_4401 (I76697,I76398,I76497);
nor I_4402 (I76213,I76296,I76697);
not I_4403 (I76755,I1869);
or I_4404 (I76772,I267704,I267707);
nand I_4405 (I76789,I267713,I267701);
not I_4406 (I76806,I76789);
nand I_4407 (I76823,I76806,I76772);
not I_4408 (I76840,I76823);
nand I_4409 (I76857,I267719,I267722);
and I_4410 (I76874,I76857,I267716);
DFFARX1 I_4411 (I76874,I1862,I76755,I76900,);
not I_4412 (I76908,I76900);
nor I_4413 (I76925,I267704,I267722);
nor I_4414 (I76942,I76900,I76925);
and I_4415 (I76959,I76900,I76925);
nor I_4416 (I76976,I76959,I76823);
DFFARX1 I_4417 (I76976,I1862,I76755,I76735,);
nand I_4418 (I77007,I267707,I267710);
nor I_4419 (I77024,I77007,I267701);
nand I_4420 (I77041,I76840,I77024);
not I_4421 (I76744,I77041);
nor I_4422 (I76747,I76942,I77041);
nor I_4423 (I77086,I77024,I76806);
nor I_4424 (I76738,I76908,I77086);
nor I_4425 (I76732,I77024,I76925);
not I_4426 (I77131,I77007);
nand I_4427 (I77148,I76925,I77131);
not I_4428 (I76726,I77148);
nor I_4429 (I76729,I76789,I77148);
nor I_4430 (I76741,I77131,I76789);
nand I_4431 (I77207,I76908,I77007);
nor I_4432 (I76723,I76806,I77207);
not I_4433 (I77265,I1869);
or I_4434 (I77282,I290433,I290430);
nand I_4435 (I77299,I290436,I290448);
not I_4436 (I77316,I77299);
nand I_4437 (I77333,I77316,I77282);
not I_4438 (I77350,I77333);
nand I_4439 (I77367,I290433,I290439);
and I_4440 (I77384,I77367,I290445);
DFFARX1 I_4441 (I77384,I1862,I77265,I77410,);
not I_4442 (I77418,I77410);
nor I_4443 (I77435,I290451,I290439);
nor I_4444 (I77452,I77410,I77435);
and I_4445 (I77469,I77410,I77435);
nor I_4446 (I77486,I77469,I77333);
DFFARX1 I_4447 (I77486,I1862,I77265,I77245,);
nand I_4448 (I77517,I290442,I290436);
nor I_4449 (I77534,I77517,I290430);
nand I_4450 (I77551,I77350,I77534);
not I_4451 (I77254,I77551);
nor I_4452 (I77257,I77452,I77551);
nor I_4453 (I77596,I77534,I77316);
nor I_4454 (I77248,I77418,I77596);
nor I_4455 (I77242,I77534,I77435);
not I_4456 (I77641,I77517);
nand I_4457 (I77658,I77435,I77641);
not I_4458 (I77236,I77658);
nor I_4459 (I77239,I77299,I77658);
nor I_4460 (I77251,I77641,I77299);
nand I_4461 (I77717,I77418,I77517);
nor I_4462 (I77233,I77316,I77717);
not I_4463 (I77775,I1869);
or I_4464 (I77792,I196393,I196372);
nand I_4465 (I77809,I196381,I196390);
not I_4466 (I77826,I77809);
nand I_4467 (I77843,I77826,I77792);
not I_4468 (I77860,I77843);
nand I_4469 (I77877,I196387,I196372);
and I_4470 (I77894,I77877,I196378);
DFFARX1 I_4471 (I77894,I1862,I77775,I77920,);
not I_4472 (I77928,I77920);
nor I_4473 (I77945,I196369,I196372);
nor I_4474 (I77962,I77920,I77945);
and I_4475 (I77979,I77920,I77945);
nor I_4476 (I77996,I77979,I77843);
DFFARX1 I_4477 (I77996,I1862,I77775,I77755,);
nand I_4478 (I78027,I196384,I196369);
nor I_4479 (I78044,I78027,I196375);
nand I_4480 (I78061,I77860,I78044);
not I_4481 (I77764,I78061);
nor I_4482 (I77767,I77962,I78061);
nor I_4483 (I78106,I78044,I77826);
nor I_4484 (I77758,I77928,I78106);
nor I_4485 (I77752,I78044,I77945);
not I_4486 (I78151,I78027);
nand I_4487 (I78168,I77945,I78151);
not I_4488 (I77746,I78168);
nor I_4489 (I77749,I77809,I78168);
nor I_4490 (I77761,I78151,I77809);
nand I_4491 (I78227,I77928,I78027);
nor I_4492 (I77743,I77826,I78227);
not I_4493 (I78285,I1869);
or I_4494 (I78302,I215344,I215347);
nand I_4495 (I78319,I215353,I215341);
not I_4496 (I78336,I78319);
nand I_4497 (I78353,I78336,I78302);
not I_4498 (I78370,I78353);
nand I_4499 (I78387,I215359,I215362);
and I_4500 (I78404,I78387,I215356);
DFFARX1 I_4501 (I78404,I1862,I78285,I78430,);
not I_4502 (I78438,I78430);
nor I_4503 (I78455,I215344,I215362);
nor I_4504 (I78472,I78430,I78455);
and I_4505 (I78489,I78430,I78455);
nor I_4506 (I78506,I78489,I78353);
DFFARX1 I_4507 (I78506,I1862,I78285,I78265,);
nand I_4508 (I78537,I215347,I215350);
nor I_4509 (I78554,I78537,I215341);
nand I_4510 (I78571,I78370,I78554);
not I_4511 (I78274,I78571);
nor I_4512 (I78277,I78472,I78571);
nor I_4513 (I78616,I78554,I78336);
nor I_4514 (I78268,I78438,I78616);
nor I_4515 (I78262,I78554,I78455);
not I_4516 (I78661,I78537);
nand I_4517 (I78678,I78455,I78661);
not I_4518 (I78256,I78678);
nor I_4519 (I78259,I78319,I78678);
nor I_4520 (I78271,I78661,I78319);
nand I_4521 (I78737,I78438,I78537);
nor I_4522 (I78253,I78336,I78737);
not I_4523 (I78795,I1869);
or I_4524 (I78812,I166881,I166860);
nand I_4525 (I78829,I166869,I166878);
not I_4526 (I78846,I78829);
nand I_4527 (I78863,I78846,I78812);
not I_4528 (I78880,I78863);
nand I_4529 (I78897,I166875,I166860);
and I_4530 (I78914,I78897,I166866);
DFFARX1 I_4531 (I78914,I1862,I78795,I78940,);
not I_4532 (I78948,I78940);
nor I_4533 (I78965,I166857,I166860);
nor I_4534 (I78982,I78940,I78965);
and I_4535 (I78999,I78940,I78965);
nor I_4536 (I79016,I78999,I78863);
DFFARX1 I_4537 (I79016,I1862,I78795,I78775,);
nand I_4538 (I79047,I166872,I166857);
nor I_4539 (I79064,I79047,I166863);
nand I_4540 (I79081,I78880,I79064);
not I_4541 (I78784,I79081);
nor I_4542 (I78787,I78982,I79081);
nor I_4543 (I79126,I79064,I78846);
nor I_4544 (I78778,I78948,I79126);
nor I_4545 (I78772,I79064,I78965);
not I_4546 (I79171,I79047);
nand I_4547 (I79188,I78965,I79171);
not I_4548 (I78766,I79188);
nor I_4549 (I78769,I78829,I79188);
nor I_4550 (I78781,I79171,I78829);
nand I_4551 (I79247,I78948,I79047);
nor I_4552 (I78763,I78846,I79247);
not I_4553 (I79305,I1869);
or I_4554 (I79322,I384916,I384916);
nand I_4555 (I79339,I384931,I384934);
not I_4556 (I79356,I79339);
nand I_4557 (I79373,I79356,I79322);
not I_4558 (I79390,I79373);
nand I_4559 (I79407,I384922,I384925);
and I_4560 (I79424,I79407,I384919);
DFFARX1 I_4561 (I79424,I1862,I79305,I79450,);
not I_4562 (I79458,I79450);
nor I_4563 (I79475,I384925,I384925);
nor I_4564 (I79492,I79450,I79475);
and I_4565 (I79509,I79450,I79475);
nor I_4566 (I79526,I79509,I79373);
DFFARX1 I_4567 (I79526,I1862,I79305,I79285,);
nand I_4568 (I79557,I384928,I384922);
nor I_4569 (I79574,I79557,I384919);
nand I_4570 (I79591,I79390,I79574);
not I_4571 (I79294,I79591);
nor I_4572 (I79297,I79492,I79591);
nor I_4573 (I79636,I79574,I79356);
nor I_4574 (I79288,I79458,I79636);
nor I_4575 (I79282,I79574,I79475);
not I_4576 (I79681,I79557);
nand I_4577 (I79698,I79475,I79681);
not I_4578 (I79276,I79698);
nor I_4579 (I79279,I79339,I79698);
nor I_4580 (I79291,I79681,I79339);
nand I_4581 (I79757,I79458,I79557);
nor I_4582 (I79273,I79356,I79757);
not I_4583 (I79815,I1869);
or I_4584 (I79832,I156868,I156847);
nand I_4585 (I79849,I156856,I156865);
not I_4586 (I79866,I79849);
nand I_4587 (I79883,I79866,I79832);
not I_4588 (I79900,I79883);
nand I_4589 (I79917,I156862,I156847);
and I_4590 (I79934,I79917,I156853);
DFFARX1 I_4591 (I79934,I1862,I79815,I79960,);
not I_4592 (I79968,I79960);
nor I_4593 (I79985,I156844,I156847);
nor I_4594 (I80002,I79960,I79985);
and I_4595 (I80019,I79960,I79985);
nor I_4596 (I80036,I80019,I79883);
DFFARX1 I_4597 (I80036,I1862,I79815,I79795,);
nand I_4598 (I80067,I156859,I156844);
nor I_4599 (I80084,I80067,I156850);
nand I_4600 (I80101,I79900,I80084);
not I_4601 (I79804,I80101);
nor I_4602 (I79807,I80002,I80101);
nor I_4603 (I80146,I80084,I79866);
nor I_4604 (I79798,I79968,I80146);
nor I_4605 (I79792,I80084,I79985);
not I_4606 (I80191,I80067);
nand I_4607 (I80208,I79985,I80191);
not I_4608 (I79786,I80208);
nor I_4609 (I79789,I79849,I80208);
nor I_4610 (I79801,I80191,I79849);
nand I_4611 (I80267,I79968,I80067);
nor I_4612 (I79783,I79866,I80267);
not I_4613 (I80325,I1869);
or I_4614 (I80342,I393314,I393314);
nand I_4615 (I80359,I393329,I393332);
not I_4616 (I80376,I80359);
nand I_4617 (I80393,I80376,I80342);
not I_4618 (I80410,I80393);
nand I_4619 (I80427,I393320,I393323);
and I_4620 (I80444,I80427,I393317);
DFFARX1 I_4621 (I80444,I1862,I80325,I80470,);
not I_4622 (I80478,I80470);
nor I_4623 (I80495,I393323,I393323);
nor I_4624 (I80512,I80470,I80495);
and I_4625 (I80529,I80470,I80495);
nor I_4626 (I80546,I80529,I80393);
DFFARX1 I_4627 (I80546,I1862,I80325,I80305,);
nand I_4628 (I80577,I393326,I393320);
nor I_4629 (I80594,I80577,I393317);
nand I_4630 (I80611,I80410,I80594);
not I_4631 (I80314,I80611);
nor I_4632 (I80317,I80512,I80611);
nor I_4633 (I80656,I80594,I80376);
nor I_4634 (I80308,I80478,I80656);
nor I_4635 (I80302,I80594,I80495);
not I_4636 (I80701,I80577);
nand I_4637 (I80718,I80495,I80701);
not I_4638 (I80296,I80718);
nor I_4639 (I80299,I80359,I80718);
nor I_4640 (I80311,I80701,I80359);
nand I_4641 (I80777,I80478,I80577);
nor I_4642 (I80293,I80376,I80777);
not I_4643 (I80835,I1869);
or I_4644 (I80852,I313624,I313618);
nand I_4645 (I80869,I313627,I313630);
not I_4646 (I80886,I80869);
nand I_4647 (I80903,I80886,I80852);
not I_4648 (I80920,I80903);
nand I_4649 (I80937,I313621,I313624);
and I_4650 (I80954,I80937,I313618);
DFFARX1 I_4651 (I80954,I1862,I80835,I80980,);
not I_4652 (I80988,I80980);
nor I_4653 (I81005,I313636,I313624);
nor I_4654 (I81022,I80980,I81005);
and I_4655 (I81039,I80980,I81005);
nor I_4656 (I81056,I81039,I80903);
DFFARX1 I_4657 (I81056,I1862,I80835,I80815,);
nand I_4658 (I81087,I313633,I313621);
nor I_4659 (I81104,I81087,I313639);
nand I_4660 (I81121,I80920,I81104);
not I_4661 (I80824,I81121);
nor I_4662 (I80827,I81022,I81121);
nor I_4663 (I81166,I81104,I80886);
nor I_4664 (I80818,I80988,I81166);
nor I_4665 (I80812,I81104,I81005);
not I_4666 (I81211,I81087);
nand I_4667 (I81228,I81005,I81211);
not I_4668 (I80806,I81228);
nor I_4669 (I80809,I80869,I81228);
nor I_4670 (I80821,I81211,I80869);
nand I_4671 (I81287,I80988,I81087);
nor I_4672 (I80803,I80886,I81287);
not I_4673 (I81345,I1869);
or I_4674 (I81362,I333650,I333644);
nand I_4675 (I81379,I333653,I333656);
not I_4676 (I81396,I81379);
nand I_4677 (I81413,I81396,I81362);
not I_4678 (I81430,I81413);
nand I_4679 (I81447,I333647,I333650);
and I_4680 (I81464,I81447,I333644);
DFFARX1 I_4681 (I81464,I1862,I81345,I81490,);
not I_4682 (I81498,I81490);
nor I_4683 (I81515,I333662,I333650);
nor I_4684 (I81532,I81490,I81515);
and I_4685 (I81549,I81490,I81515);
nor I_4686 (I81566,I81549,I81413);
DFFARX1 I_4687 (I81566,I1862,I81345,I81325,);
nand I_4688 (I81597,I333659,I333647);
nor I_4689 (I81614,I81597,I333665);
nand I_4690 (I81631,I81430,I81614);
not I_4691 (I81334,I81631);
nor I_4692 (I81337,I81532,I81631);
nor I_4693 (I81676,I81614,I81396);
nor I_4694 (I81328,I81498,I81676);
nor I_4695 (I81322,I81614,I81515);
not I_4696 (I81721,I81597);
nand I_4697 (I81738,I81515,I81721);
not I_4698 (I81316,I81738);
nor I_4699 (I81319,I81379,I81738);
nor I_4700 (I81331,I81721,I81379);
nand I_4701 (I81797,I81498,I81597);
nor I_4702 (I81313,I81396,I81797);
not I_4703 (I81855,I1869);
or I_4704 (I81872,I160030,I160009);
nand I_4705 (I81889,I160018,I160027);
not I_4706 (I81906,I81889);
nand I_4707 (I81923,I81906,I81872);
not I_4708 (I81940,I81923);
nand I_4709 (I81957,I160024,I160009);
and I_4710 (I81974,I81957,I160015);
DFFARX1 I_4711 (I81974,I1862,I81855,I82000,);
not I_4712 (I82008,I82000);
nor I_4713 (I82025,I160006,I160009);
nor I_4714 (I82042,I82000,I82025);
and I_4715 (I82059,I82000,I82025);
nor I_4716 (I82076,I82059,I81923);
DFFARX1 I_4717 (I82076,I1862,I81855,I81835,);
nand I_4718 (I82107,I160021,I160006);
nor I_4719 (I82124,I82107,I160012);
nand I_4720 (I82141,I81940,I82124);
not I_4721 (I81844,I82141);
nor I_4722 (I81847,I82042,I82141);
nor I_4723 (I82186,I82124,I81906);
nor I_4724 (I81838,I82008,I82186);
nor I_4725 (I81832,I82124,I82025);
not I_4726 (I82231,I82107);
nand I_4727 (I82248,I82025,I82231);
not I_4728 (I81826,I82248);
nor I_4729 (I81829,I81889,I82248);
nor I_4730 (I81841,I82231,I81889);
nand I_4731 (I82307,I82008,I82107);
nor I_4732 (I81823,I81906,I82307);
not I_4733 (I82365,I1869);
or I_4734 (I82382,I307300,I307294);
nand I_4735 (I82399,I307303,I307306);
not I_4736 (I82416,I82399);
nand I_4737 (I82433,I82416,I82382);
not I_4738 (I82450,I82433);
nand I_4739 (I82467,I307297,I307300);
and I_4740 (I82484,I82467,I307294);
DFFARX1 I_4741 (I82484,I1862,I82365,I82510,);
not I_4742 (I82518,I82510);
nor I_4743 (I82535,I307312,I307300);
nor I_4744 (I82552,I82510,I82535);
and I_4745 (I82569,I82510,I82535);
nor I_4746 (I82586,I82569,I82433);
DFFARX1 I_4747 (I82586,I1862,I82365,I82345,);
nand I_4748 (I82617,I307309,I307297);
nor I_4749 (I82634,I82617,I307315);
nand I_4750 (I82651,I82450,I82634);
not I_4751 (I82354,I82651);
nor I_4752 (I82357,I82552,I82651);
nor I_4753 (I82696,I82634,I82416);
nor I_4754 (I82348,I82518,I82696);
nor I_4755 (I82342,I82634,I82535);
not I_4756 (I82741,I82617);
nand I_4757 (I82758,I82535,I82741);
not I_4758 (I82336,I82758);
nor I_4759 (I82339,I82399,I82758);
nor I_4760 (I82351,I82741,I82399);
nand I_4761 (I82817,I82518,I82617);
nor I_4762 (I82333,I82416,I82817);
not I_4763 (I82875,I1869);
or I_4764 (I82892,I315205,I315199);
nand I_4765 (I82909,I315208,I315211);
not I_4766 (I82926,I82909);
nand I_4767 (I82943,I82926,I82892);
not I_4768 (I82960,I82943);
nand I_4769 (I82977,I315202,I315205);
and I_4770 (I82994,I82977,I315199);
DFFARX1 I_4771 (I82994,I1862,I82875,I83020,);
not I_4772 (I83028,I83020);
nor I_4773 (I83045,I315217,I315205);
nor I_4774 (I83062,I83020,I83045);
and I_4775 (I83079,I83020,I83045);
nor I_4776 (I83096,I83079,I82943);
DFFARX1 I_4777 (I83096,I1862,I82875,I82855,);
nand I_4778 (I83127,I315214,I315202);
nor I_4779 (I83144,I83127,I315220);
nand I_4780 (I83161,I82960,I83144);
not I_4781 (I82864,I83161);
nor I_4782 (I82867,I83062,I83161);
nor I_4783 (I83206,I83144,I82926);
nor I_4784 (I82858,I83028,I83206);
nor I_4785 (I82852,I83144,I83045);
not I_4786 (I83251,I83127);
nand I_4787 (I83268,I83045,I83251);
not I_4788 (I82846,I83268);
nor I_4789 (I82849,I82909,I83268);
nor I_4790 (I82861,I83251,I82909);
nand I_4791 (I83327,I83028,I83127);
nor I_4792 (I82843,I82926,I83327);
not I_4793 (I83385,I1869);
or I_4794 (I83402,I185853,I185832);
nand I_4795 (I83419,I185841,I185850);
not I_4796 (I83436,I83419);
nand I_4797 (I83453,I83436,I83402);
not I_4798 (I83470,I83453);
nand I_4799 (I83487,I185847,I185832);
and I_4800 (I83504,I83487,I185838);
DFFARX1 I_4801 (I83504,I1862,I83385,I83530,);
not I_4802 (I83538,I83530);
nor I_4803 (I83555,I185829,I185832);
nor I_4804 (I83572,I83530,I83555);
and I_4805 (I83589,I83530,I83555);
nor I_4806 (I83606,I83589,I83453);
DFFARX1 I_4807 (I83606,I1862,I83385,I83365,);
nand I_4808 (I83637,I185844,I185829);
nor I_4809 (I83654,I83637,I185835);
nand I_4810 (I83671,I83470,I83654);
not I_4811 (I83374,I83671);
nor I_4812 (I83377,I83572,I83671);
nor I_4813 (I83716,I83654,I83436);
nor I_4814 (I83368,I83538,I83716);
nor I_4815 (I83362,I83654,I83555);
not I_4816 (I83761,I83637);
nand I_4817 (I83778,I83555,I83761);
not I_4818 (I83356,I83778);
nor I_4819 (I83359,I83419,I83778);
nor I_4820 (I83371,I83761,I83419);
nand I_4821 (I83837,I83538,I83637);
nor I_4822 (I83353,I83436,I83837);
not I_4823 (I83895,I1869);
or I_4824 (I83912,I360527,I360521);
nand I_4825 (I83929,I360530,I360533);
not I_4826 (I83946,I83929);
nand I_4827 (I83963,I83946,I83912);
not I_4828 (I83980,I83963);
nand I_4829 (I83997,I360524,I360527);
and I_4830 (I84014,I83997,I360521);
DFFARX1 I_4831 (I84014,I1862,I83895,I84040,);
not I_4832 (I84048,I84040);
nor I_4833 (I84065,I360539,I360527);
nor I_4834 (I84082,I84040,I84065);
and I_4835 (I84099,I84040,I84065);
nor I_4836 (I84116,I84099,I83963);
DFFARX1 I_4837 (I84116,I1862,I83895,I83875,);
nand I_4838 (I84147,I360536,I360524);
nor I_4839 (I84164,I84147,I360542);
nand I_4840 (I84181,I83980,I84164);
not I_4841 (I83884,I84181);
nor I_4842 (I83887,I84082,I84181);
nor I_4843 (I84226,I84164,I83946);
nor I_4844 (I83878,I84048,I84226);
nor I_4845 (I83872,I84164,I84065);
not I_4846 (I84271,I84147);
nand I_4847 (I84288,I84065,I84271);
not I_4848 (I83866,I84288);
nor I_4849 (I83869,I83929,I84288);
nor I_4850 (I83881,I84271,I83929);
nand I_4851 (I84347,I84048,I84147);
nor I_4852 (I83863,I83946,I84347);
not I_4853 (I84405,I1869);
or I_4854 (I84422,I276272,I276275);
nand I_4855 (I84439,I276281,I276269);
not I_4856 (I84456,I84439);
nand I_4857 (I84473,I84456,I84422);
not I_4858 (I84490,I84473);
nand I_4859 (I84507,I276287,I276290);
and I_4860 (I84524,I84507,I276284);
DFFARX1 I_4861 (I84524,I1862,I84405,I84550,);
not I_4862 (I84558,I84550);
nor I_4863 (I84575,I276272,I276290);
nor I_4864 (I84592,I84550,I84575);
and I_4865 (I84609,I84550,I84575);
nor I_4866 (I84626,I84609,I84473);
DFFARX1 I_4867 (I84626,I1862,I84405,I84385,);
nand I_4868 (I84657,I276275,I276278);
nor I_4869 (I84674,I84657,I276269);
nand I_4870 (I84691,I84490,I84674);
not I_4871 (I84394,I84691);
nor I_4872 (I84397,I84592,I84691);
nor I_4873 (I84736,I84674,I84456);
nor I_4874 (I84388,I84558,I84736);
nor I_4875 (I84382,I84674,I84575);
not I_4876 (I84781,I84657);
nand I_4877 (I84798,I84575,I84781);
not I_4878 (I84376,I84798);
nor I_4879 (I84379,I84439,I84798);
nor I_4880 (I84391,I84781,I84439);
nand I_4881 (I84857,I84558,I84657);
nor I_4882 (I84373,I84456,I84857);
not I_4883 (I84915,I1869);
or I_4884 (I84932,I245332,I245335);
nand I_4885 (I84949,I245341,I245329);
not I_4886 (I84966,I84949);
nand I_4887 (I84983,I84966,I84932);
not I_4888 (I85000,I84983);
nand I_4889 (I85017,I245347,I245350);
and I_4890 (I85034,I85017,I245344);
DFFARX1 I_4891 (I85034,I1862,I84915,I85060,);
not I_4892 (I85068,I85060);
nor I_4893 (I85085,I245332,I245350);
nor I_4894 (I85102,I85060,I85085);
and I_4895 (I85119,I85060,I85085);
nor I_4896 (I85136,I85119,I84983);
DFFARX1 I_4897 (I85136,I1862,I84915,I84895,);
nand I_4898 (I85167,I245335,I245338);
nor I_4899 (I85184,I85167,I245329);
nand I_4900 (I85201,I85000,I85184);
not I_4901 (I84904,I85201);
nor I_4902 (I84907,I85102,I85201);
nor I_4903 (I85246,I85184,I84966);
nor I_4904 (I84898,I85068,I85246);
nor I_4905 (I84892,I85184,I85085);
not I_4906 (I85291,I85167);
nand I_4907 (I85308,I85085,I85291);
not I_4908 (I84886,I85308);
nor I_4909 (I84889,I84949,I85308);
nor I_4910 (I84901,I85291,I84949);
nand I_4911 (I85367,I85068,I85167);
nor I_4912 (I84883,I84966,I85367);
not I_4913 (I85425,I1869);
or I_4914 (I85442,I135261,I135240);
nand I_4915 (I85459,I135249,I135258);
not I_4916 (I85476,I85459);
nand I_4917 (I85493,I85476,I85442);
not I_4918 (I85510,I85493);
nand I_4919 (I85527,I135255,I135240);
and I_4920 (I85544,I85527,I135246);
DFFARX1 I_4921 (I85544,I1862,I85425,I85570,);
not I_4922 (I85578,I85570);
nor I_4923 (I85595,I135237,I135240);
nor I_4924 (I85612,I85570,I85595);
and I_4925 (I85629,I85570,I85595);
nor I_4926 (I85646,I85629,I85493);
DFFARX1 I_4927 (I85646,I1862,I85425,I85405,);
nand I_4928 (I85677,I135252,I135237);
nor I_4929 (I85694,I85677,I135243);
nand I_4930 (I85711,I85510,I85694);
not I_4931 (I85414,I85711);
nor I_4932 (I85417,I85612,I85711);
nor I_4933 (I85756,I85694,I85476);
nor I_4934 (I85408,I85578,I85756);
nor I_4935 (I85402,I85694,I85595);
not I_4936 (I85801,I85677);
nand I_4937 (I85818,I85595,I85801);
not I_4938 (I85396,I85818);
nor I_4939 (I85399,I85459,I85818);
nor I_4940 (I85411,I85801,I85459);
nand I_4941 (I85877,I85578,I85677);
nor I_4942 (I85393,I85476,I85877);
not I_4943 (I85935,I1869);
or I_4944 (I85952,I193231,I193210);
nand I_4945 (I85969,I193219,I193228);
not I_4946 (I85986,I85969);
nand I_4947 (I86003,I85986,I85952);
not I_4948 (I86020,I86003);
nand I_4949 (I86037,I193225,I193210);
and I_4950 (I86054,I86037,I193216);
DFFARX1 I_4951 (I86054,I1862,I85935,I86080,);
not I_4952 (I86088,I86080);
nor I_4953 (I86105,I193207,I193210);
nor I_4954 (I86122,I86080,I86105);
and I_4955 (I86139,I86080,I86105);
nor I_4956 (I86156,I86139,I86003);
DFFARX1 I_4957 (I86156,I1862,I85935,I85915,);
nand I_4958 (I86187,I193222,I193207);
nor I_4959 (I86204,I86187,I193213);
nand I_4960 (I86221,I86020,I86204);
not I_4961 (I85924,I86221);
nor I_4962 (I85927,I86122,I86221);
nor I_4963 (I86266,I86204,I85986);
nor I_4964 (I85918,I86088,I86266);
nor I_4965 (I85912,I86204,I86105);
not I_4966 (I86311,I86187);
nand I_4967 (I86328,I86105,I86311);
not I_4968 (I85906,I86328);
nor I_4969 (I85909,I85969,I86328);
nor I_4970 (I85921,I86311,I85969);
nand I_4971 (I86387,I86088,I86187);
nor I_4972 (I85903,I85986,I86387);
not I_4973 (I86445,I1869);
or I_4974 (I86462,I380496,I380496);
nand I_4975 (I86479,I380511,I380514);
not I_4976 (I86496,I86479);
nand I_4977 (I86513,I86496,I86462);
not I_4978 (I86530,I86513);
nand I_4979 (I86547,I380502,I380505);
and I_4980 (I86564,I86547,I380499);
DFFARX1 I_4981 (I86564,I1862,I86445,I86590,);
not I_4982 (I86598,I86590);
nor I_4983 (I86615,I380505,I380505);
nor I_4984 (I86632,I86590,I86615);
and I_4985 (I86649,I86590,I86615);
nor I_4986 (I86666,I86649,I86513);
DFFARX1 I_4987 (I86666,I1862,I86445,I86425,);
nand I_4988 (I86697,I380508,I380502);
nor I_4989 (I86714,I86697,I380499);
nand I_4990 (I86731,I86530,I86714);
not I_4991 (I86434,I86731);
nor I_4992 (I86437,I86632,I86731);
nor I_4993 (I86776,I86714,I86496);
nor I_4994 (I86428,I86598,I86776);
nor I_4995 (I86422,I86714,I86615);
not I_4996 (I86821,I86697);
nand I_4997 (I86838,I86615,I86821);
not I_4998 (I86416,I86838);
nor I_4999 (I86419,I86479,I86838);
nor I_5000 (I86431,I86821,I86479);
nand I_5001 (I86897,I86598,I86697);
nor I_5002 (I86413,I86496,I86897);
not I_5003 (I86955,I1869);
or I_5004 (I86972,I117870,I117849);
nand I_5005 (I86989,I117858,I117867);
not I_5006 (I87006,I86989);
nand I_5007 (I87023,I87006,I86972);
not I_5008 (I87040,I87023);
nand I_5009 (I87057,I117864,I117849);
and I_5010 (I87074,I87057,I117855);
DFFARX1 I_5011 (I87074,I1862,I86955,I87100,);
not I_5012 (I87108,I87100);
nor I_5013 (I87125,I117846,I117849);
nor I_5014 (I87142,I87100,I87125);
and I_5015 (I87159,I87100,I87125);
nor I_5016 (I87176,I87159,I87023);
DFFARX1 I_5017 (I87176,I1862,I86955,I86935,);
nand I_5018 (I87207,I117861,I117846);
nor I_5019 (I87224,I87207,I117852);
nand I_5020 (I87241,I87040,I87224);
not I_5021 (I86944,I87241);
nor I_5022 (I86947,I87142,I87241);
nor I_5023 (I87286,I87224,I87006);
nor I_5024 (I86938,I87108,I87286);
nor I_5025 (I86932,I87224,I87125);
not I_5026 (I87331,I87207);
nand I_5027 (I87348,I87125,I87331);
not I_5028 (I86926,I87348);
nor I_5029 (I86929,I86989,I87348);
nor I_5030 (I86941,I87331,I86989);
nand I_5031 (I87407,I87108,I87207);
nor I_5032 (I86923,I87006,I87407);
not I_5033 (I87465,I1869);
or I_5034 (I87482,I209156,I209159);
nand I_5035 (I87499,I209165,I209153);
not I_5036 (I87516,I87499);
nand I_5037 (I87533,I87516,I87482);
not I_5038 (I87550,I87533);
nand I_5039 (I87567,I209171,I209174);
and I_5040 (I87584,I87567,I209168);
DFFARX1 I_5041 (I87584,I1862,I87465,I87610,);
not I_5042 (I87618,I87610);
nor I_5043 (I87635,I209156,I209174);
nor I_5044 (I87652,I87610,I87635);
and I_5045 (I87669,I87610,I87635);
nor I_5046 (I87686,I87669,I87533);
DFFARX1 I_5047 (I87686,I1862,I87465,I87445,);
nand I_5048 (I87717,I209159,I209162);
nor I_5049 (I87734,I87717,I209153);
nand I_5050 (I87751,I87550,I87734);
not I_5051 (I87454,I87751);
nor I_5052 (I87457,I87652,I87751);
nor I_5053 (I87796,I87734,I87516);
nor I_5054 (I87448,I87618,I87796);
nor I_5055 (I87442,I87734,I87635);
not I_5056 (I87841,I87717);
nand I_5057 (I87858,I87635,I87841);
not I_5058 (I87436,I87858);
nor I_5059 (I87439,I87499,I87858);
nor I_5060 (I87451,I87841,I87499);
nand I_5061 (I87917,I87618,I87717);
nor I_5062 (I87433,I87516,I87917);
not I_5063 (I87975,I1869);
or I_5064 (I87992,I375192,I375192);
nand I_5065 (I88009,I375207,I375210);
not I_5066 (I88026,I88009);
nand I_5067 (I88043,I88026,I87992);
not I_5068 (I88060,I88043);
nand I_5069 (I88077,I375198,I375201);
and I_5070 (I88094,I88077,I375195);
DFFARX1 I_5071 (I88094,I1862,I87975,I88120,);
not I_5072 (I88128,I88120);
nor I_5073 (I88145,I375201,I375201);
nor I_5074 (I88162,I88120,I88145);
and I_5075 (I88179,I88120,I88145);
nor I_5076 (I88196,I88179,I88043);
DFFARX1 I_5077 (I88196,I1862,I87975,I87955,);
nand I_5078 (I88227,I375204,I375198);
nor I_5079 (I88244,I88227,I375195);
nand I_5080 (I88261,I88060,I88244);
not I_5081 (I87964,I88261);
nor I_5082 (I87967,I88162,I88261);
nor I_5083 (I88306,I88244,I88026);
nor I_5084 (I87958,I88128,I88306);
nor I_5085 (I87952,I88244,I88145);
not I_5086 (I88351,I88227);
nand I_5087 (I88368,I88145,I88351);
not I_5088 (I87946,I88368);
nor I_5089 (I87949,I88009,I88368);
nor I_5090 (I87961,I88351,I88009);
nand I_5091 (I88427,I88128,I88227);
nor I_5092 (I87943,I88026,I88427);
not I_5093 (I88485,I1869);
or I_5094 (I88502,I283888,I283891);
nand I_5095 (I88519,I283897,I283885);
not I_5096 (I88536,I88519);
nand I_5097 (I88553,I88536,I88502);
not I_5098 (I88570,I88553);
nand I_5099 (I88587,I283903,I283906);
and I_5100 (I88604,I88587,I283900);
DFFARX1 I_5101 (I88604,I1862,I88485,I88630,);
not I_5102 (I88638,I88630);
nor I_5103 (I88655,I283888,I283906);
nor I_5104 (I88672,I88630,I88655);
and I_5105 (I88689,I88630,I88655);
nor I_5106 (I88706,I88689,I88553);
DFFARX1 I_5107 (I88706,I1862,I88485,I88465,);
nand I_5108 (I88737,I283891,I283894);
nor I_5109 (I88754,I88737,I283885);
nand I_5110 (I88771,I88570,I88754);
not I_5111 (I88474,I88771);
nor I_5112 (I88477,I88672,I88771);
nor I_5113 (I88816,I88754,I88536);
nor I_5114 (I88468,I88638,I88816);
nor I_5115 (I88462,I88754,I88655);
not I_5116 (I88861,I88737);
nand I_5117 (I88878,I88655,I88861);
not I_5118 (I88456,I88878);
nor I_5119 (I88459,I88519,I88878);
nor I_5120 (I88471,I88861,I88519);
nand I_5121 (I88937,I88638,I88737);
nor I_5122 (I88453,I88536,I88937);
not I_5123 (I88995,I1869);
or I_5124 (I89012,I372540,I372540);
nand I_5125 (I89029,I372555,I372558);
not I_5126 (I89046,I89029);
nand I_5127 (I89063,I89046,I89012);
not I_5128 (I89080,I89063);
nand I_5129 (I89097,I372546,I372549);
and I_5130 (I89114,I89097,I372543);
DFFARX1 I_5131 (I89114,I1862,I88995,I89140,);
not I_5132 (I89148,I89140);
nor I_5133 (I89165,I372549,I372549);
nor I_5134 (I89182,I89140,I89165);
and I_5135 (I89199,I89140,I89165);
nor I_5136 (I89216,I89199,I89063);
DFFARX1 I_5137 (I89216,I1862,I88995,I88975,);
nand I_5138 (I89247,I372552,I372546);
nor I_5139 (I89264,I89247,I372543);
nand I_5140 (I89281,I89080,I89264);
not I_5141 (I88984,I89281);
nor I_5142 (I88987,I89182,I89281);
nor I_5143 (I89326,I89264,I89046);
nor I_5144 (I88978,I89148,I89326);
nor I_5145 (I88972,I89264,I89165);
not I_5146 (I89371,I89247);
nand I_5147 (I89388,I89165,I89371);
not I_5148 (I88966,I89388);
nor I_5149 (I88969,I89029,I89388);
nor I_5150 (I88981,I89371,I89029);
nand I_5151 (I89447,I89148,I89247);
nor I_5152 (I88963,I89046,I89447);
not I_5153 (I89505,I1869);
or I_5154 (I89522,I114061,I114055);
nand I_5155 (I89539,I114061,I114073);
not I_5156 (I89556,I89539);
nand I_5157 (I89573,I89556,I89522);
not I_5158 (I89590,I89573);
nand I_5159 (I89607,I114067,I114058);
and I_5160 (I89624,I89607,I114055);
DFFARX1 I_5161 (I89624,I1862,I89505,I89650,);
not I_5162 (I89658,I89650);
nor I_5163 (I89675,I114070,I114058);
nor I_5164 (I89692,I89650,I89675);
and I_5165 (I89709,I89650,I89675);
nor I_5166 (I89726,I89709,I89573);
DFFARX1 I_5167 (I89726,I1862,I89505,I89485,);
nand I_5168 (I89757,I114064,I114064);
nor I_5169 (I89774,I89757,I114058);
nand I_5170 (I89791,I89590,I89774);
not I_5171 (I89494,I89791);
nor I_5172 (I89497,I89692,I89791);
nor I_5173 (I89836,I89774,I89556);
nor I_5174 (I89488,I89658,I89836);
nor I_5175 (I89482,I89774,I89675);
not I_5176 (I89881,I89757);
nand I_5177 (I89898,I89675,I89881);
not I_5178 (I89476,I89898);
nor I_5179 (I89479,I89539,I89898);
nor I_5180 (I89491,I89881,I89539);
nand I_5181 (I89957,I89658,I89757);
nor I_5182 (I89473,I89556,I89957);
not I_5183 (I90015,I1869);
or I_5184 (I90032,I275796,I275799);
nand I_5185 (I90049,I275805,I275793);
not I_5186 (I90066,I90049);
nand I_5187 (I90083,I90066,I90032);
not I_5188 (I90100,I90083);
nand I_5189 (I90117,I275811,I275814);
and I_5190 (I90134,I90117,I275808);
DFFARX1 I_5191 (I90134,I1862,I90015,I90160,);
not I_5192 (I90168,I90160);
nor I_5193 (I90185,I275796,I275814);
nor I_5194 (I90202,I90160,I90185);
and I_5195 (I90219,I90160,I90185);
nor I_5196 (I90236,I90219,I90083);
DFFARX1 I_5197 (I90236,I1862,I90015,I89995,);
nand I_5198 (I90267,I275799,I275802);
nor I_5199 (I90284,I90267,I275793);
nand I_5200 (I90301,I90100,I90284);
not I_5201 (I90004,I90301);
nor I_5202 (I90007,I90202,I90301);
nor I_5203 (I90346,I90284,I90066);
nor I_5204 (I89998,I90168,I90346);
nor I_5205 (I89992,I90284,I90185);
not I_5206 (I90391,I90267);
nand I_5207 (I90408,I90185,I90391);
not I_5208 (I89986,I90408);
nor I_5209 (I89989,I90049,I90408);
nor I_5210 (I90001,I90391,I90049);
nand I_5211 (I90467,I90168,I90267);
nor I_5212 (I89983,I90066,I90467);
not I_5213 (I90525,I1869);
or I_5214 (I90542,I143166,I143145);
nand I_5215 (I90559,I143154,I143163);
not I_5216 (I90576,I90559);
nand I_5217 (I90593,I90576,I90542);
not I_5218 (I90610,I90593);
nand I_5219 (I90627,I143160,I143145);
and I_5220 (I90644,I90627,I143151);
DFFARX1 I_5221 (I90644,I1862,I90525,I90670,);
not I_5222 (I90678,I90670);
nor I_5223 (I90695,I143142,I143145);
nor I_5224 (I90712,I90670,I90695);
and I_5225 (I90729,I90670,I90695);
nor I_5226 (I90746,I90729,I90593);
DFFARX1 I_5227 (I90746,I1862,I90525,I90505,);
nand I_5228 (I90777,I143157,I143142);
nor I_5229 (I90794,I90777,I143148);
nand I_5230 (I90811,I90610,I90794);
not I_5231 (I90514,I90811);
nor I_5232 (I90517,I90712,I90811);
nor I_5233 (I90856,I90794,I90576);
nor I_5234 (I90508,I90678,I90856);
nor I_5235 (I90502,I90794,I90695);
not I_5236 (I90901,I90777);
nand I_5237 (I90918,I90695,I90901);
not I_5238 (I90496,I90918);
nor I_5239 (I90499,I90559,I90918);
nor I_5240 (I90511,I90901,I90559);
nand I_5241 (I90977,I90678,I90777);
nor I_5242 (I90493,I90576,I90977);
not I_5243 (I91035,I1869);
or I_5244 (I91052,I214868,I214871);
nand I_5245 (I91069,I214877,I214865);
not I_5246 (I91086,I91069);
nand I_5247 (I91103,I91086,I91052);
not I_5248 (I91120,I91103);
nand I_5249 (I91137,I214883,I214886);
and I_5250 (I91154,I91137,I214880);
DFFARX1 I_5251 (I91154,I1862,I91035,I91180,);
not I_5252 (I91188,I91180);
nor I_5253 (I91205,I214868,I214886);
nor I_5254 (I91222,I91180,I91205);
and I_5255 (I91239,I91180,I91205);
nor I_5256 (I91256,I91239,I91103);
DFFARX1 I_5257 (I91256,I1862,I91035,I91015,);
nand I_5258 (I91287,I214871,I214874);
nor I_5259 (I91304,I91287,I214865);
nand I_5260 (I91321,I91120,I91304);
not I_5261 (I91024,I91321);
nor I_5262 (I91027,I91222,I91321);
nor I_5263 (I91366,I91304,I91086);
nor I_5264 (I91018,I91188,I91366);
nor I_5265 (I91012,I91304,I91205);
not I_5266 (I91411,I91287);
nand I_5267 (I91428,I91205,I91411);
not I_5268 (I91006,I91428);
nor I_5269 (I91009,I91069,I91428);
nor I_5270 (I91021,I91411,I91069);
nand I_5271 (I91487,I91188,I91287);
nor I_5272 (I91003,I91086,I91487);
not I_5273 (I91545,I1869);
or I_5274 (I91562,I129991,I129970);
nand I_5275 (I91579,I129979,I129988);
not I_5276 (I91596,I91579);
nand I_5277 (I91613,I91596,I91562);
not I_5278 (I91630,I91613);
nand I_5279 (I91647,I129985,I129970);
and I_5280 (I91664,I91647,I129976);
DFFARX1 I_5281 (I91664,I1862,I91545,I91690,);
not I_5282 (I91698,I91690);
nor I_5283 (I91715,I129967,I129970);
nor I_5284 (I91732,I91690,I91715);
and I_5285 (I91749,I91690,I91715);
nor I_5286 (I91766,I91749,I91613);
DFFARX1 I_5287 (I91766,I1862,I91545,I91525,);
nand I_5288 (I91797,I129982,I129967);
nor I_5289 (I91814,I91797,I129973);
nand I_5290 (I91831,I91630,I91814);
not I_5291 (I91534,I91831);
nor I_5292 (I91537,I91732,I91831);
nor I_5293 (I91876,I91814,I91596);
nor I_5294 (I91528,I91698,I91876);
nor I_5295 (I91522,I91814,I91715);
not I_5296 (I91921,I91797);
nand I_5297 (I91938,I91715,I91921);
not I_5298 (I91516,I91938);
nor I_5299 (I91519,I91579,I91938);
nor I_5300 (I91531,I91921,I91579);
nand I_5301 (I91997,I91698,I91797);
nor I_5302 (I91513,I91596,I91997);
not I_5303 (I92055,I1869);
or I_5304 (I92072,I128410,I128389);
nand I_5305 (I92089,I128398,I128407);
not I_5306 (I92106,I92089);
nand I_5307 (I92123,I92106,I92072);
not I_5308 (I92140,I92123);
nand I_5309 (I92157,I128404,I128389);
and I_5310 (I92174,I92157,I128395);
DFFARX1 I_5311 (I92174,I1862,I92055,I92200,);
not I_5312 (I92208,I92200);
nor I_5313 (I92225,I128386,I128389);
nor I_5314 (I92242,I92200,I92225);
and I_5315 (I92259,I92200,I92225);
nor I_5316 (I92276,I92259,I92123);
DFFARX1 I_5317 (I92276,I1862,I92055,I92035,);
nand I_5318 (I92307,I128401,I128386);
nor I_5319 (I92324,I92307,I128392);
nand I_5320 (I92341,I92140,I92324);
not I_5321 (I92044,I92341);
nor I_5322 (I92047,I92242,I92341);
nor I_5323 (I92386,I92324,I92106);
nor I_5324 (I92038,I92208,I92386);
nor I_5325 (I92032,I92324,I92225);
not I_5326 (I92431,I92307);
nand I_5327 (I92448,I92225,I92431);
not I_5328 (I92026,I92448);
nor I_5329 (I92029,I92089,I92448);
nor I_5330 (I92041,I92431,I92089);
nand I_5331 (I92507,I92208,I92307);
nor I_5332 (I92023,I92106,I92507);
not I_5333 (I92565,I1869);
or I_5334 (I92582,I319948,I319942);
nand I_5335 (I92599,I319951,I319954);
not I_5336 (I92616,I92599);
nand I_5337 (I92633,I92616,I92582);
not I_5338 (I92650,I92633);
nand I_5339 (I92667,I319945,I319948);
and I_5340 (I92684,I92667,I319942);
DFFARX1 I_5341 (I92684,I1862,I92565,I92710,);
not I_5342 (I92718,I92710);
nor I_5343 (I92735,I319960,I319948);
nor I_5344 (I92752,I92710,I92735);
and I_5345 (I92769,I92710,I92735);
nor I_5346 (I92786,I92769,I92633);
DFFARX1 I_5347 (I92786,I1862,I92565,I92545,);
nand I_5348 (I92817,I319957,I319945);
nor I_5349 (I92834,I92817,I319963);
nand I_5350 (I92851,I92650,I92834);
not I_5351 (I92554,I92851);
nor I_5352 (I92557,I92752,I92851);
nor I_5353 (I92896,I92834,I92616);
nor I_5354 (I92548,I92718,I92896);
nor I_5355 (I92542,I92834,I92735);
not I_5356 (I92941,I92817);
nand I_5357 (I92958,I92735,I92941);
not I_5358 (I92536,I92958);
nor I_5359 (I92539,I92599,I92958);
nor I_5360 (I92551,I92941,I92599);
nand I_5361 (I93017,I92718,I92817);
nor I_5362 (I92533,I92616,I93017);
not I_5363 (I93075,I1869);
or I_5364 (I93092,I372098,I372098);
nand I_5365 (I93109,I372113,I372116);
not I_5366 (I93126,I93109);
nand I_5367 (I93143,I93126,I93092);
not I_5368 (I93160,I93143);
nand I_5369 (I93177,I372104,I372107);
and I_5370 (I93194,I93177,I372101);
DFFARX1 I_5371 (I93194,I1862,I93075,I93220,);
not I_5372 (I93228,I93220);
nor I_5373 (I93245,I372107,I372107);
nor I_5374 (I93262,I93220,I93245);
and I_5375 (I93279,I93220,I93245);
nor I_5376 (I93296,I93279,I93143);
DFFARX1 I_5377 (I93296,I1862,I93075,I93055,);
nand I_5378 (I93327,I372110,I372104);
nor I_5379 (I93344,I93327,I372101);
nand I_5380 (I93361,I93160,I93344);
not I_5381 (I93064,I93361);
nor I_5382 (I93067,I93262,I93361);
nor I_5383 (I93406,I93344,I93126);
nor I_5384 (I93058,I93228,I93406);
nor I_5385 (I93052,I93344,I93245);
not I_5386 (I93451,I93327);
nand I_5387 (I93468,I93245,I93451);
not I_5388 (I93046,I93468);
nor I_5389 (I93049,I93109,I93468);
nor I_5390 (I93061,I93451,I93109);
nand I_5391 (I93527,I93228,I93327);
nor I_5392 (I93043,I93126,I93527);
not I_5393 (I93585,I1869);
or I_5394 (I93602,I397292,I397292);
nand I_5395 (I93619,I397307,I397310);
not I_5396 (I93636,I93619);
nand I_5397 (I93653,I93636,I93602);
not I_5398 (I93670,I93653);
nand I_5399 (I93687,I397298,I397301);
and I_5400 (I93704,I93687,I397295);
DFFARX1 I_5401 (I93704,I1862,I93585,I93730,);
not I_5402 (I93738,I93730);
nor I_5403 (I93755,I397301,I397301);
nor I_5404 (I93772,I93730,I93755);
and I_5405 (I93789,I93730,I93755);
nor I_5406 (I93806,I93789,I93653);
DFFARX1 I_5407 (I93806,I1862,I93585,I93565,);
nand I_5408 (I93837,I397304,I397298);
nor I_5409 (I93854,I93837,I397295);
nand I_5410 (I93871,I93670,I93854);
not I_5411 (I93574,I93871);
nor I_5412 (I93577,I93772,I93871);
nor I_5413 (I93916,I93854,I93636);
nor I_5414 (I93568,I93738,I93916);
nor I_5415 (I93562,I93854,I93755);
not I_5416 (I93961,I93837);
nand I_5417 (I93978,I93755,I93961);
not I_5418 (I93556,I93978);
nor I_5419 (I93559,I93619,I93978);
nor I_5420 (I93571,I93961,I93619);
nand I_5421 (I94037,I93738,I93837);
nor I_5422 (I93553,I93636,I94037);
not I_5423 (I94095,I1869);
or I_5424 (I94112,I393756,I393756);
nand I_5425 (I94129,I393771,I393774);
not I_5426 (I94146,I94129);
nand I_5427 (I94163,I94146,I94112);
not I_5428 (I94180,I94163);
nand I_5429 (I94197,I393762,I393765);
and I_5430 (I94214,I94197,I393759);
DFFARX1 I_5431 (I94214,I1862,I94095,I94240,);
not I_5432 (I94248,I94240);
nor I_5433 (I94265,I393765,I393765);
nor I_5434 (I94282,I94240,I94265);
and I_5435 (I94299,I94240,I94265);
nor I_5436 (I94316,I94299,I94163);
DFFARX1 I_5437 (I94316,I1862,I94095,I94075,);
nand I_5438 (I94347,I393768,I393762);
nor I_5439 (I94364,I94347,I393759);
nand I_5440 (I94381,I94180,I94364);
not I_5441 (I94084,I94381);
nor I_5442 (I94087,I94282,I94381);
nor I_5443 (I94426,I94364,I94146);
nor I_5444 (I94078,I94248,I94426);
nor I_5445 (I94072,I94364,I94265);
not I_5446 (I94471,I94347);
nand I_5447 (I94488,I94265,I94471);
not I_5448 (I94066,I94488);
nor I_5449 (I94069,I94129,I94488);
nor I_5450 (I94081,I94471,I94129);
nand I_5451 (I94547,I94248,I94347);
nor I_5452 (I94063,I94146,I94547);
not I_5453 (I94605,I1869);
or I_5454 (I94622,I246760,I246763);
nand I_5455 (I94639,I246769,I246757);
not I_5456 (I94656,I94639);
nand I_5457 (I94673,I94656,I94622);
not I_5458 (I94690,I94673);
nand I_5459 (I94707,I246775,I246778);
and I_5460 (I94724,I94707,I246772);
DFFARX1 I_5461 (I94724,I1862,I94605,I94750,);
not I_5462 (I94758,I94750);
nor I_5463 (I94775,I246760,I246778);
nor I_5464 (I94792,I94750,I94775);
and I_5465 (I94809,I94750,I94775);
nor I_5466 (I94826,I94809,I94673);
DFFARX1 I_5467 (I94826,I1862,I94605,I94585,);
nand I_5468 (I94857,I246763,I246766);
nor I_5469 (I94874,I94857,I246757);
nand I_5470 (I94891,I94690,I94874);
not I_5471 (I94594,I94891);
nor I_5472 (I94597,I94792,I94891);
nor I_5473 (I94936,I94874,I94656);
nor I_5474 (I94588,I94758,I94936);
nor I_5475 (I94582,I94874,I94775);
not I_5476 (I94981,I94857);
nand I_5477 (I94998,I94775,I94981);
not I_5478 (I94576,I94998);
nor I_5479 (I94579,I94639,I94998);
nor I_5480 (I94591,I94981,I94639);
nand I_5481 (I95057,I94758,I94857);
nor I_5482 (I94573,I94656,I95057);
not I_5483 (I95115,I1869);
or I_5484 (I95132,I313097,I313091);
nand I_5485 (I95149,I313100,I313103);
not I_5486 (I95166,I95149);
nand I_5487 (I95183,I95166,I95132);
not I_5488 (I95200,I95183);
nand I_5489 (I95217,I313094,I313097);
and I_5490 (I95234,I95217,I313091);
DFFARX1 I_5491 (I95234,I1862,I95115,I95260,);
not I_5492 (I95268,I95260);
nor I_5493 (I95285,I313109,I313097);
nor I_5494 (I95302,I95260,I95285);
and I_5495 (I95319,I95260,I95285);
nor I_5496 (I95336,I95319,I95183);
DFFARX1 I_5497 (I95336,I1862,I95115,I95095,);
nand I_5498 (I95367,I313106,I313094);
nor I_5499 (I95384,I95367,I313112);
nand I_5500 (I95401,I95200,I95384);
not I_5501 (I95104,I95401);
nor I_5502 (I95107,I95302,I95401);
nor I_5503 (I95446,I95384,I95166);
nor I_5504 (I95098,I95268,I95446);
nor I_5505 (I95092,I95384,I95285);
not I_5506 (I95491,I95367);
nand I_5507 (I95508,I95285,I95491);
not I_5508 (I95086,I95508);
nor I_5509 (I95089,I95149,I95508);
nor I_5510 (I95101,I95491,I95149);
nand I_5511 (I95567,I95268,I95367);
nor I_5512 (I95083,I95166,I95567);
not I_5513 (I95625,I1869);
or I_5514 (I95642,I167408,I167387);
nand I_5515 (I95659,I167396,I167405);
not I_5516 (I95676,I95659);
nand I_5517 (I95693,I95676,I95642);
not I_5518 (I95710,I95693);
nand I_5519 (I95727,I167402,I167387);
and I_5520 (I95744,I95727,I167393);
DFFARX1 I_5521 (I95744,I1862,I95625,I95770,);
not I_5522 (I95778,I95770);
nor I_5523 (I95795,I167384,I167387);
nor I_5524 (I95812,I95770,I95795);
and I_5525 (I95829,I95770,I95795);
nor I_5526 (I95846,I95829,I95693);
DFFARX1 I_5527 (I95846,I1862,I95625,I95605,);
nand I_5528 (I95877,I167399,I167384);
nor I_5529 (I95894,I95877,I167390);
nand I_5530 (I95911,I95710,I95894);
not I_5531 (I95614,I95911);
nor I_5532 (I95617,I95812,I95911);
nor I_5533 (I95956,I95894,I95676);
nor I_5534 (I95608,I95778,I95956);
nor I_5535 (I95602,I95894,I95795);
not I_5536 (I96001,I95877);
nand I_5537 (I96018,I95795,I96001);
not I_5538 (I95596,I96018);
nor I_5539 (I95599,I95659,I96018);
nor I_5540 (I95611,I96001,I95659);
nand I_5541 (I96077,I95778,I95877);
nor I_5542 (I95593,I95676,I96077);
not I_5543 (I96135,I1869);
or I_5544 (I96152,I353149,I353143);
nand I_5545 (I96169,I353152,I353155);
not I_5546 (I96186,I96169);
nand I_5547 (I96203,I96186,I96152);
not I_5548 (I96220,I96203);
nand I_5549 (I96237,I353146,I353149);
and I_5550 (I96254,I96237,I353143);
DFFARX1 I_5551 (I96254,I1862,I96135,I96280,);
not I_5552 (I96288,I96280);
nor I_5553 (I96305,I353161,I353149);
nor I_5554 (I96322,I96280,I96305);
and I_5555 (I96339,I96280,I96305);
nor I_5556 (I96356,I96339,I96203);
DFFARX1 I_5557 (I96356,I1862,I96135,I96115,);
nand I_5558 (I96387,I353158,I353146);
nor I_5559 (I96404,I96387,I353164);
nand I_5560 (I96421,I96220,I96404);
not I_5561 (I96124,I96421);
nor I_5562 (I96127,I96322,I96421);
nor I_5563 (I96466,I96404,I96186);
nor I_5564 (I96118,I96288,I96466);
nor I_5565 (I96112,I96404,I96305);
not I_5566 (I96511,I96387);
nand I_5567 (I96528,I96305,I96511);
not I_5568 (I96106,I96528);
nor I_5569 (I96109,I96169,I96528);
nor I_5570 (I96121,I96511,I96169);
nand I_5571 (I96587,I96288,I96387);
nor I_5572 (I96103,I96186,I96587);
not I_5573 (I96645,I1869);
or I_5574 (I96662,I118397,I118376);
nand I_5575 (I96679,I118385,I118394);
not I_5576 (I96696,I96679);
nand I_5577 (I96713,I96696,I96662);
not I_5578 (I96730,I96713);
nand I_5579 (I96747,I118391,I118376);
and I_5580 (I96764,I96747,I118382);
DFFARX1 I_5581 (I96764,I1862,I96645,I96790,);
not I_5582 (I96798,I96790);
nor I_5583 (I96815,I118373,I118376);
nor I_5584 (I96832,I96790,I96815);
and I_5585 (I96849,I96790,I96815);
nor I_5586 (I96866,I96849,I96713);
DFFARX1 I_5587 (I96866,I1862,I96645,I96625,);
nand I_5588 (I96897,I118388,I118373);
nor I_5589 (I96914,I96897,I118379);
nand I_5590 (I96931,I96730,I96914);
not I_5591 (I96634,I96931);
nor I_5592 (I96637,I96832,I96931);
nor I_5593 (I96976,I96914,I96696);
nor I_5594 (I96628,I96798,I96976);
nor I_5595 (I96622,I96914,I96815);
not I_5596 (I97021,I96897);
nand I_5597 (I97038,I96815,I97021);
not I_5598 (I96616,I97038);
nor I_5599 (I96619,I96679,I97038);
nor I_5600 (I96631,I97021,I96679);
nand I_5601 (I97097,I96798,I96897);
nor I_5602 (I96613,I96696,I97097);
not I_5603 (I97155,I1869);
or I_5604 (I97172,I396408,I396408);
nand I_5605 (I97189,I396423,I396426);
not I_5606 (I97206,I97189);
nand I_5607 (I97223,I97206,I97172);
not I_5608 (I97240,I97223);
nand I_5609 (I97257,I396414,I396417);
and I_5610 (I97274,I97257,I396411);
DFFARX1 I_5611 (I97274,I1862,I97155,I97300,);
not I_5612 (I97308,I97300);
nor I_5613 (I97325,I396417,I396417);
nor I_5614 (I97342,I97300,I97325);
and I_5615 (I97359,I97300,I97325);
nor I_5616 (I97376,I97359,I97223);
DFFARX1 I_5617 (I97376,I1862,I97155,I97135,);
nand I_5618 (I97407,I396420,I396414);
nor I_5619 (I97424,I97407,I396411);
nand I_5620 (I97441,I97240,I97424);
not I_5621 (I97144,I97441);
nor I_5622 (I97147,I97342,I97441);
nor I_5623 (I97486,I97424,I97206);
nor I_5624 (I97138,I97308,I97486);
nor I_5625 (I97132,I97424,I97325);
not I_5626 (I97531,I97407);
nand I_5627 (I97548,I97325,I97531);
not I_5628 (I97126,I97548);
nor I_5629 (I97129,I97189,I97548);
nor I_5630 (I97141,I97531,I97189);
nand I_5631 (I97607,I97308,I97407);
nor I_5632 (I97123,I97206,I97607);
not I_5633 (I97665,I1869);
or I_5634 (I97682,I133153,I133132);
nand I_5635 (I97699,I133141,I133150);
not I_5636 (I97716,I97699);
nand I_5637 (I97733,I97716,I97682);
not I_5638 (I97750,I97733);
nand I_5639 (I97767,I133147,I133132);
and I_5640 (I97784,I97767,I133138);
DFFARX1 I_5641 (I97784,I1862,I97665,I97810,);
not I_5642 (I97818,I97810);
nor I_5643 (I97835,I133129,I133132);
nor I_5644 (I97852,I97810,I97835);
and I_5645 (I97869,I97810,I97835);
nor I_5646 (I97886,I97869,I97733);
DFFARX1 I_5647 (I97886,I1862,I97665,I97645,);
nand I_5648 (I97917,I133144,I133129);
nor I_5649 (I97934,I97917,I133135);
nand I_5650 (I97951,I97750,I97934);
not I_5651 (I97654,I97951);
nor I_5652 (I97657,I97852,I97951);
nor I_5653 (I97996,I97934,I97716);
nor I_5654 (I97648,I97818,I97996);
nor I_5655 (I97642,I97934,I97835);
not I_5656 (I98041,I97917);
nand I_5657 (I98058,I97835,I98041);
not I_5658 (I97636,I98058);
nor I_5659 (I97639,I97699,I98058);
nor I_5660 (I97651,I98041,I97699);
nand I_5661 (I98117,I97818,I97917);
nor I_5662 (I97633,I97716,I98117);
not I_5663 (I98175,I1869);
or I_5664 (I98192,I178475,I178454);
nand I_5665 (I98209,I178463,I178472);
not I_5666 (I98226,I98209);
nand I_5667 (I98243,I98226,I98192);
not I_5668 (I98260,I98243);
nand I_5669 (I98277,I178469,I178454);
and I_5670 (I98294,I98277,I178460);
DFFARX1 I_5671 (I98294,I1862,I98175,I98320,);
not I_5672 (I98328,I98320);
nor I_5673 (I98345,I178451,I178454);
nor I_5674 (I98362,I98320,I98345);
and I_5675 (I98379,I98320,I98345);
nor I_5676 (I98396,I98379,I98243);
DFFARX1 I_5677 (I98396,I1862,I98175,I98155,);
nand I_5678 (I98427,I178466,I178451);
nor I_5679 (I98444,I98427,I178457);
nand I_5680 (I98461,I98260,I98444);
not I_5681 (I98164,I98461);
nor I_5682 (I98167,I98362,I98461);
nor I_5683 (I98506,I98444,I98226);
nor I_5684 (I98158,I98328,I98506);
nor I_5685 (I98152,I98444,I98345);
not I_5686 (I98551,I98427);
nand I_5687 (I98568,I98345,I98551);
not I_5688 (I98146,I98568);
nor I_5689 (I98149,I98209,I98568);
nor I_5690 (I98161,I98551,I98209);
nand I_5691 (I98627,I98328,I98427);
nor I_5692 (I98143,I98226,I98627);
not I_5693 (I98685,I1869);
or I_5694 (I98702,I213440,I213443);
nand I_5695 (I98719,I213449,I213437);
not I_5696 (I98736,I98719);
nand I_5697 (I98753,I98736,I98702);
not I_5698 (I98770,I98753);
nand I_5699 (I98787,I213455,I213458);
and I_5700 (I98804,I98787,I213452);
DFFARX1 I_5701 (I98804,I1862,I98685,I98830,);
not I_5702 (I98838,I98830);
nor I_5703 (I98855,I213440,I213458);
nor I_5704 (I98872,I98830,I98855);
and I_5705 (I98889,I98830,I98855);
nor I_5706 (I98906,I98889,I98753);
DFFARX1 I_5707 (I98906,I1862,I98685,I98665,);
nand I_5708 (I98937,I213443,I213446);
nor I_5709 (I98954,I98937,I213437);
nand I_5710 (I98971,I98770,I98954);
not I_5711 (I98674,I98971);
nor I_5712 (I98677,I98872,I98971);
nor I_5713 (I99016,I98954,I98736);
nor I_5714 (I98668,I98838,I99016);
nor I_5715 (I98662,I98954,I98855);
not I_5716 (I99061,I98937);
nand I_5717 (I99078,I98855,I99061);
not I_5718 (I98656,I99078);
nor I_5719 (I98659,I98719,I99078);
nor I_5720 (I98671,I99061,I98719);
nand I_5721 (I99137,I98838,I98937);
nor I_5722 (I98653,I98736,I99137);
not I_5723 (I99195,I1869);
or I_5724 (I99212,I166354,I166333);
nand I_5725 (I99229,I166342,I166351);
not I_5726 (I99246,I99229);
nand I_5727 (I99263,I99246,I99212);
not I_5728 (I99280,I99263);
nand I_5729 (I99297,I166348,I166333);
and I_5730 (I99314,I99297,I166339);
DFFARX1 I_5731 (I99314,I1862,I99195,I99340,);
not I_5732 (I99348,I99340);
nor I_5733 (I99365,I166330,I166333);
nor I_5734 (I99382,I99340,I99365);
and I_5735 (I99399,I99340,I99365);
nor I_5736 (I99416,I99399,I99263);
DFFARX1 I_5737 (I99416,I1862,I99195,I99175,);
nand I_5738 (I99447,I166345,I166330);
nor I_5739 (I99464,I99447,I166336);
nand I_5740 (I99481,I99280,I99464);
not I_5741 (I99184,I99481);
nor I_5742 (I99187,I99382,I99481);
nor I_5743 (I99526,I99464,I99246);
nor I_5744 (I99178,I99348,I99526);
nor I_5745 (I99172,I99464,I99365);
not I_5746 (I99571,I99447);
nand I_5747 (I99588,I99365,I99571);
not I_5748 (I99166,I99588);
nor I_5749 (I99169,I99229,I99588);
nor I_5750 (I99181,I99571,I99229);
nand I_5751 (I99647,I99348,I99447);
nor I_5752 (I99163,I99246,I99647);
not I_5753 (I99705,I1869);
or I_5754 (I99722,I170043,I170022);
nand I_5755 (I99739,I170031,I170040);
not I_5756 (I99756,I99739);
nand I_5757 (I99773,I99756,I99722);
not I_5758 (I99790,I99773);
nand I_5759 (I99807,I170037,I170022);
and I_5760 (I99824,I99807,I170028);
DFFARX1 I_5761 (I99824,I1862,I99705,I99850,);
not I_5762 (I99858,I99850);
nor I_5763 (I99875,I170019,I170022);
nor I_5764 (I99892,I99850,I99875);
and I_5765 (I99909,I99850,I99875);
nor I_5766 (I99926,I99909,I99773);
DFFARX1 I_5767 (I99926,I1862,I99705,I99685,);
nand I_5768 (I99957,I170034,I170019);
nor I_5769 (I99974,I99957,I170025);
nand I_5770 (I99991,I99790,I99974);
not I_5771 (I99694,I99991);
nor I_5772 (I99697,I99892,I99991);
nor I_5773 (I100036,I99974,I99756);
nor I_5774 (I99688,I99858,I100036);
nor I_5775 (I99682,I99974,I99875);
not I_5776 (I100081,I99957);
nand I_5777 (I100098,I99875,I100081);
not I_5778 (I99676,I100098);
nor I_5779 (I99679,I99739,I100098);
nor I_5780 (I99691,I100081,I99739);
nand I_5781 (I100157,I99858,I99957);
nor I_5782 (I99673,I99756,I100157);
not I_5783 (I100215,I1869);
or I_5784 (I100232,I205824,I205827);
nand I_5785 (I100249,I205833,I205821);
not I_5786 (I100266,I100249);
nand I_5787 (I100283,I100266,I100232);
not I_5788 (I100300,I100283);
nand I_5789 (I100317,I205839,I205842);
and I_5790 (I100334,I100317,I205836);
DFFARX1 I_5791 (I100334,I1862,I100215,I100360,);
not I_5792 (I100368,I100360);
nor I_5793 (I100385,I205824,I205842);
nor I_5794 (I100402,I100360,I100385);
and I_5795 (I100419,I100360,I100385);
nor I_5796 (I100436,I100419,I100283);
DFFARX1 I_5797 (I100436,I1862,I100215,I100195,);
nand I_5798 (I100467,I205827,I205830);
nor I_5799 (I100484,I100467,I205821);
nand I_5800 (I100501,I100300,I100484);
not I_5801 (I100204,I100501);
nor I_5802 (I100207,I100402,I100501);
nor I_5803 (I100546,I100484,I100266);
nor I_5804 (I100198,I100368,I100546);
nor I_5805 (I100192,I100484,I100385);
not I_5806 (I100591,I100467);
nand I_5807 (I100608,I100385,I100591);
not I_5808 (I100186,I100608);
nor I_5809 (I100189,I100249,I100608);
nor I_5810 (I100201,I100591,I100249);
nand I_5811 (I100667,I100368,I100467);
nor I_5812 (I100183,I100266,I100667);
not I_5813 (I100725,I1869);
or I_5814 (I100742,I380938,I380938);
nand I_5815 (I100759,I380953,I380956);
not I_5816 (I100776,I100759);
nand I_5817 (I100793,I100776,I100742);
not I_5818 (I100810,I100793);
nand I_5819 (I100827,I380944,I380947);
and I_5820 (I100844,I100827,I380941);
DFFARX1 I_5821 (I100844,I1862,I100725,I100870,);
not I_5822 (I100878,I100870);
nor I_5823 (I100895,I380947,I380947);
nor I_5824 (I100912,I100870,I100895);
and I_5825 (I100929,I100870,I100895);
nor I_5826 (I100946,I100929,I100793);
DFFARX1 I_5827 (I100946,I1862,I100725,I100705,);
nand I_5828 (I100977,I380950,I380944);
nor I_5829 (I100994,I100977,I380941);
nand I_5830 (I101011,I100810,I100994);
not I_5831 (I100714,I101011);
nor I_5832 (I100717,I100912,I101011);
nor I_5833 (I101056,I100994,I100776);
nor I_5834 (I100708,I100878,I101056);
nor I_5835 (I100702,I100994,I100895);
not I_5836 (I101101,I100977);
nand I_5837 (I101118,I100895,I101101);
not I_5838 (I100696,I101118);
nor I_5839 (I100699,I100759,I101118);
nor I_5840 (I100711,I101101,I100759);
nand I_5841 (I101177,I100878,I100977);
nor I_5842 (I100693,I100776,I101177);
not I_5843 (I101235,I1869);
or I_5844 (I101252,I270560,I270563);
nand I_5845 (I101269,I270569,I270557);
not I_5846 (I101286,I101269);
nand I_5847 (I101303,I101286,I101252);
not I_5848 (I101320,I101303);
nand I_5849 (I101337,I270575,I270578);
and I_5850 (I101354,I101337,I270572);
DFFARX1 I_5851 (I101354,I1862,I101235,I101380,);
not I_5852 (I101388,I101380);
nor I_5853 (I101405,I270560,I270578);
nor I_5854 (I101422,I101380,I101405);
and I_5855 (I101439,I101380,I101405);
nor I_5856 (I101456,I101439,I101303);
DFFARX1 I_5857 (I101456,I1862,I101235,I101215,);
nand I_5858 (I101487,I270563,I270566);
nor I_5859 (I101504,I101487,I270557);
nand I_5860 (I101521,I101320,I101504);
not I_5861 (I101224,I101521);
nor I_5862 (I101227,I101422,I101521);
nor I_5863 (I101566,I101504,I101286);
nor I_5864 (I101218,I101388,I101566);
nor I_5865 (I101212,I101504,I101405);
not I_5866 (I101611,I101487);
nand I_5867 (I101628,I101405,I101611);
not I_5868 (I101206,I101628);
nor I_5869 (I101209,I101269,I101628);
nor I_5870 (I101221,I101611,I101269);
nand I_5871 (I101687,I101388,I101487);
nor I_5872 (I101203,I101286,I101687);
not I_5873 (I101745,I1869);
or I_5874 (I101762,I315732,I315726);
nand I_5875 (I101779,I315735,I315738);
not I_5876 (I101796,I101779);
nand I_5877 (I101813,I101796,I101762);
not I_5878 (I101830,I101813);
nand I_5879 (I101847,I315729,I315732);
and I_5880 (I101864,I101847,I315726);
DFFARX1 I_5881 (I101864,I1862,I101745,I101890,);
not I_5882 (I101898,I101890);
nor I_5883 (I101915,I315744,I315732);
nor I_5884 (I101932,I101890,I101915);
and I_5885 (I101949,I101890,I101915);
nor I_5886 (I101966,I101949,I101813);
DFFARX1 I_5887 (I101966,I1862,I101745,I101725,);
nand I_5888 (I101997,I315741,I315729);
nor I_5889 (I102014,I101997,I315747);
nand I_5890 (I102031,I101830,I102014);
not I_5891 (I101734,I102031);
nor I_5892 (I101737,I101932,I102031);
nor I_5893 (I102076,I102014,I101796);
nor I_5894 (I101728,I101898,I102076);
nor I_5895 (I101722,I102014,I101915);
not I_5896 (I102121,I101997);
nand I_5897 (I102138,I101915,I102121);
not I_5898 (I101716,I102138);
nor I_5899 (I101719,I101779,I102138);
nor I_5900 (I101731,I102121,I101779);
nand I_5901 (I102197,I101898,I101997);
nor I_5902 (I101713,I101796,I102197);
not I_5903 (I102249,I1869);
and I_5904 (I102266,I180053,I180035);
nor I_5905 (I102283,I102266,I180056);
nand I_5906 (I102300,I180032,I180047);
nor I_5907 (I102317,I102300,I102283);
nor I_5908 (I102223,I102317,I102300);
not I_5909 (I102348,I102317);
not I_5910 (I102365,I102300);
or I_5911 (I102382,I180050,I180032);
nor I_5912 (I102399,I102382,I180038);
nand I_5913 (I102416,I102365,I102399);
not I_5914 (I102238,I102416);
nor I_5915 (I102447,I102317,I180044);
and I_5916 (I102464,I180041,I180035);
nor I_5917 (I102481,I102464,I102317);
nor I_5918 (I102241,I102481,I102416);
nor I_5919 (I102226,I102464,I102399);
nand I_5920 (I102526,I102464,I180044);
not I_5921 (I102543,I102526);
nand I_5922 (I102560,I102399,I102543);
nand I_5923 (I102577,I102348,I102560);
DFFARX1 I_5924 (I102577,I1862,I102249,I102229,);
nand I_5925 (I102235,I102464,I102300);
nand I_5926 (I102232,I102447,I102464);
not I_5927 (I102657,I1869);
and I_5928 (I102674,I240093,I240093);
nor I_5929 (I102691,I102674,I240114);
nand I_5930 (I102708,I240096,I240099);
nor I_5931 (I102725,I102708,I102691);
nor I_5932 (I102631,I102725,I102708);
not I_5933 (I102756,I102725);
not I_5934 (I102773,I102708);
or I_5935 (I102790,I240102,I240111);
nor I_5936 (I102807,I102790,I240108);
nand I_5937 (I102824,I102773,I102807);
not I_5938 (I102646,I102824);
nor I_5939 (I102855,I102725,I240099);
and I_5940 (I102872,I240096,I240105);
nor I_5941 (I102889,I102872,I102725);
nor I_5942 (I102649,I102889,I102824);
nor I_5943 (I102634,I102872,I102807);
nand I_5944 (I102934,I102872,I240099);
not I_5945 (I102951,I102934);
nand I_5946 (I102968,I102807,I102951);
nand I_5947 (I102985,I102756,I102968);
DFFARX1 I_5948 (I102985,I1862,I102657,I102637,);
nand I_5949 (I102643,I102872,I102708);
nand I_5950 (I102640,I102855,I102872);
not I_5951 (I103065,I1869);
and I_5952 (I103082,I269605,I269605);
nor I_5953 (I103099,I103082,I269626);
nand I_5954 (I103116,I269608,I269611);
nor I_5955 (I103133,I103116,I103099);
nor I_5956 (I103039,I103133,I103116);
not I_5957 (I103164,I103133);
not I_5958 (I103181,I103116);
or I_5959 (I103198,I269614,I269623);
nor I_5960 (I103215,I103198,I269620);
nand I_5961 (I103232,I103181,I103215);
not I_5962 (I103054,I103232);
nor I_5963 (I103263,I103133,I269611);
and I_5964 (I103280,I269608,I269617);
nor I_5965 (I103297,I103280,I103133);
nor I_5966 (I103057,I103297,I103232);
nor I_5967 (I103042,I103280,I103215);
nand I_5968 (I103342,I103280,I269611);
not I_5969 (I103359,I103342);
nand I_5970 (I103376,I103215,I103359);
nand I_5971 (I103393,I103164,I103376);
DFFARX1 I_5972 (I103393,I1862,I103065,I103045,);
nand I_5973 (I103051,I103280,I103116);
nand I_5974 (I103048,I103263,I103280);
not I_5975 (I103473,I1869);
and I_5976 (I103490,I223909,I223909);
nor I_5977 (I103507,I103490,I223930);
nand I_5978 (I103524,I223912,I223915);
nor I_5979 (I103541,I103524,I103507);
nor I_5980 (I103447,I103541,I103524);
not I_5981 (I103572,I103541);
not I_5982 (I103589,I103524);
or I_5983 (I103606,I223918,I223927);
nor I_5984 (I103623,I103606,I223924);
nand I_5985 (I103640,I103589,I103623);
not I_5986 (I103462,I103640);
nor I_5987 (I103671,I103541,I223915);
and I_5988 (I103688,I223912,I223921);
nor I_5989 (I103705,I103688,I103541);
nor I_5990 (I103465,I103705,I103640);
nor I_5991 (I103450,I103688,I103623);
nand I_5992 (I103750,I103688,I223915);
not I_5993 (I103767,I103750);
nand I_5994 (I103784,I103623,I103767);
nand I_5995 (I103801,I103572,I103784);
DFFARX1 I_5996 (I103801,I1862,I103473,I103453,);
nand I_5997 (I103459,I103688,I103524);
nand I_5998 (I103456,I103671,I103688);
not I_5999 (I103881,I1869);
and I_6000 (I103898,I178999,I178981);
nor I_6001 (I103915,I103898,I179002);
nand I_6002 (I103932,I178978,I178993);
nor I_6003 (I103949,I103932,I103915);
nor I_6004 (I103855,I103949,I103932);
not I_6005 (I103980,I103949);
not I_6006 (I103997,I103932);
or I_6007 (I104014,I178996,I178978);
nor I_6008 (I104031,I104014,I178984);
nand I_6009 (I104048,I103997,I104031);
not I_6010 (I103870,I104048);
nor I_6011 (I104079,I103949,I178990);
and I_6012 (I104096,I178987,I178981);
nor I_6013 (I104113,I104096,I103949);
nor I_6014 (I103873,I104113,I104048);
nor I_6015 (I103858,I104096,I104031);
nand I_6016 (I104158,I104096,I178990);
not I_6017 (I104175,I104158);
nand I_6018 (I104192,I104031,I104175);
nand I_6019 (I104209,I103980,I104192);
DFFARX1 I_6020 (I104209,I1862,I103881,I103861,);
nand I_6021 (I103867,I104096,I103932);
nand I_6022 (I103864,I104079,I104096);
not I_6023 (I104289,I1869);
and I_6024 (I104306,I1447,I1175);
nor I_6025 (I104323,I104306,I1631);
nand I_6026 (I104340,I903,I1295);
nor I_6027 (I104357,I104340,I104323);
nor I_6028 (I104263,I104357,I104340);
not I_6029 (I104388,I104357);
not I_6030 (I104405,I104340);
or I_6031 (I104422,I1703,I1063);
nor I_6032 (I104439,I104422,I743);
nand I_6033 (I104456,I104405,I104439);
not I_6034 (I104278,I104456);
nor I_6035 (I104487,I104357,I1431);
and I_6036 (I104504,I1183,I1143);
nor I_6037 (I104521,I104504,I104357);
nor I_6038 (I104281,I104521,I104456);
nor I_6039 (I104266,I104504,I104439);
nand I_6040 (I104566,I104504,I1431);
not I_6041 (I104583,I104566);
nand I_6042 (I104600,I104439,I104583);
nand I_6043 (I104617,I104388,I104600);
DFFARX1 I_6044 (I104617,I1862,I104289,I104269,);
nand I_6045 (I104275,I104504,I104340);
nand I_6046 (I104272,I104487,I104504);
not I_6047 (I104697,I1869);
and I_6048 (I104714,I289388,I289397);
nor I_6049 (I104731,I104714,I289379);
nand I_6050 (I104748,I289394,I289382);
nor I_6051 (I104765,I104748,I104731);
nor I_6052 (I104671,I104765,I104748);
not I_6053 (I104796,I104765);
not I_6054 (I104813,I104748);
or I_6055 (I104830,I289376,I289379);
nor I_6056 (I104847,I104830,I289376);
nand I_6057 (I104864,I104813,I104847);
not I_6058 (I104686,I104864);
nor I_6059 (I104895,I104765,I289382);
and I_6060 (I104912,I289385,I289391);
nor I_6061 (I104929,I104912,I104765);
nor I_6062 (I104689,I104929,I104864);
nor I_6063 (I104674,I104912,I104847);
nand I_6064 (I104974,I104912,I289382);
not I_6065 (I104991,I104974);
nand I_6066 (I105008,I104847,I104991);
nand I_6067 (I105025,I104796,I105008);
DFFARX1 I_6068 (I105025,I1862,I104697,I104677,);
nand I_6069 (I104683,I104912,I104748);
nand I_6070 (I104680,I104895,I104912);
not I_6071 (I105105,I1869);
and I_6072 (I105122,I388909,I388903);
nor I_6073 (I105139,I105122,I388906);
nand I_6074 (I105156,I388900,I388900);
nor I_6075 (I105173,I105156,I105139);
nor I_6076 (I105079,I105173,I105156);
not I_6077 (I105204,I105173);
not I_6078 (I105221,I105156);
or I_6079 (I105238,I388897,I388894);
nor I_6080 (I105255,I105238,I388897);
nand I_6081 (I105272,I105221,I105255);
not I_6082 (I105094,I105272);
nor I_6083 (I105303,I105173,I388894);
and I_6084 (I105320,I388903,I388912);
nor I_6085 (I105337,I105320,I105173);
nor I_6086 (I105097,I105337,I105272);
nor I_6087 (I105082,I105320,I105255);
nand I_6088 (I105382,I105320,I388894);
not I_6089 (I105399,I105382);
nand I_6090 (I105416,I105255,I105399);
nand I_6091 (I105433,I105204,I105416);
DFFARX1 I_6092 (I105433,I1862,I105105,I105085,);
nand I_6093 (I105091,I105320,I105156);
nand I_6094 (I105088,I105303,I105320);
not I_6095 (I105513,I1869);
and I_6096 (I105530,I405705,I405699);
nor I_6097 (I105547,I105530,I405702);
nand I_6098 (I105564,I405696,I405696);
nor I_6099 (I105581,I105564,I105547);
nor I_6100 (I105487,I105581,I105564);
not I_6101 (I105612,I105581);
not I_6102 (I105629,I105564);
or I_6103 (I105646,I405693,I405690);
nor I_6104 (I105663,I105646,I405693);
nand I_6105 (I105680,I105629,I105663);
not I_6106 (I105502,I105680);
nor I_6107 (I105711,I105581,I405690);
and I_6108 (I105728,I405699,I405708);
nor I_6109 (I105745,I105728,I105581);
nor I_6110 (I105505,I105745,I105680);
nor I_6111 (I105490,I105728,I105663);
nand I_6112 (I105790,I105728,I405690);
not I_6113 (I105807,I105790);
nand I_6114 (I105824,I105663,I105807);
nand I_6115 (I105841,I105612,I105824);
DFFARX1 I_6116 (I105841,I1862,I105513,I105493,);
nand I_6117 (I105499,I105728,I105564);
nand I_6118 (I105496,I105711,I105728);
not I_6119 (I105921,I1869);
and I_6120 (I105938,I345256,I345241);
nor I_6121 (I105955,I105938,I345244);
nand I_6122 (I105972,I345238,I345253);
nor I_6123 (I105989,I105972,I105955);
nor I_6124 (I105895,I105989,I105972);
not I_6125 (I106020,I105989);
not I_6126 (I106037,I105972);
or I_6127 (I106054,I345241,I345244);
nor I_6128 (I106071,I106054,I345238);
nand I_6129 (I106088,I106037,I106071);
not I_6130 (I105910,I106088);
nor I_6131 (I106119,I105989,I345259);
and I_6132 (I106136,I345250,I345247);
nor I_6133 (I106153,I106136,I105989);
nor I_6134 (I105913,I106153,I106088);
nor I_6135 (I105898,I106136,I106071);
nand I_6136 (I106198,I106136,I345259);
not I_6137 (I106215,I106198);
nand I_6138 (I106232,I106071,I106215);
nand I_6139 (I106249,I106020,I106232);
DFFARX1 I_6140 (I106249,I1862,I105921,I105901,);
nand I_6141 (I105907,I106136,I105972);
nand I_6142 (I105904,I106119,I106136);
not I_6143 (I106329,I1869);
and I_6144 (I106346,I378743,I378737);
nor I_6145 (I106363,I106346,I378740);
nand I_6146 (I106380,I378734,I378734);
nor I_6147 (I106397,I106380,I106363);
nor I_6148 (I106303,I106397,I106380);
not I_6149 (I106428,I106397);
not I_6150 (I106445,I106380);
or I_6151 (I106462,I378731,I378728);
nor I_6152 (I106479,I106462,I378731);
nand I_6153 (I106496,I106445,I106479);
not I_6154 (I106318,I106496);
nor I_6155 (I106527,I106397,I378728);
and I_6156 (I106544,I378737,I378746);
nor I_6157 (I106561,I106544,I106397);
nor I_6158 (I106321,I106561,I106496);
nor I_6159 (I106306,I106544,I106479);
nand I_6160 (I106606,I106544,I378728);
not I_6161 (I106623,I106606);
nand I_6162 (I106640,I106479,I106623);
nand I_6163 (I106657,I106428,I106640);
DFFARX1 I_6164 (I106657,I1862,I106329,I106309,);
nand I_6165 (I106315,I106544,I106380);
nand I_6166 (I106312,I106527,I106544);
not I_6167 (I106737,I1869);
and I_6168 (I106754,I350526,I350511);
nor I_6169 (I106771,I106754,I350514);
nand I_6170 (I106788,I350508,I350523);
nor I_6171 (I106805,I106788,I106771);
nor I_6172 (I106711,I106805,I106788);
not I_6173 (I106836,I106805);
not I_6174 (I106853,I106788);
or I_6175 (I106870,I350511,I350514);
nor I_6176 (I106887,I106870,I350508);
nand I_6177 (I106904,I106853,I106887);
not I_6178 (I106726,I106904);
nor I_6179 (I106935,I106805,I350529);
and I_6180 (I106952,I350520,I350517);
nor I_6181 (I106969,I106952,I106805);
nor I_6182 (I106729,I106969,I106904);
nor I_6183 (I106714,I106952,I106887);
nand I_6184 (I107014,I106952,I350529);
not I_6185 (I107031,I107014);
nand I_6186 (I107048,I106887,I107031);
nand I_6187 (I107065,I106836,I107048);
DFFARX1 I_6188 (I107065,I1862,I106737,I106717,);
nand I_6189 (I106723,I106952,I106788);
nand I_6190 (I106720,I106935,I106952);
not I_6191 (I107145,I1869);
and I_6192 (I107162,I309420,I309405);
nor I_6193 (I107179,I107162,I309408);
nand I_6194 (I107196,I309402,I309417);
nor I_6195 (I107213,I107196,I107179);
nor I_6196 (I107119,I107213,I107196);
not I_6197 (I107244,I107213);
not I_6198 (I107261,I107196);
or I_6199 (I107278,I309405,I309408);
nor I_6200 (I107295,I107278,I309402);
nand I_6201 (I107312,I107261,I107295);
not I_6202 (I107134,I107312);
nor I_6203 (I107343,I107213,I309423);
and I_6204 (I107360,I309414,I309411);
nor I_6205 (I107377,I107360,I107213);
nor I_6206 (I107137,I107377,I107312);
nor I_6207 (I107122,I107360,I107295);
nand I_6208 (I107422,I107360,I309423);
not I_6209 (I107439,I107422);
nand I_6210 (I107456,I107295,I107439);
nand I_6211 (I107473,I107244,I107456);
DFFARX1 I_6212 (I107473,I1862,I107145,I107125,);
nand I_6213 (I107131,I107360,I107196);
nand I_6214 (I107128,I107343,I107360);
not I_6215 (I107553,I1869);
and I_6216 (I107570,I323649,I323634);
nor I_6217 (I107587,I107570,I323637);
nand I_6218 (I107604,I323631,I323646);
nor I_6219 (I107621,I107604,I107587);
nor I_6220 (I107527,I107621,I107604);
not I_6221 (I107652,I107621);
not I_6222 (I107669,I107604);
or I_6223 (I107686,I323634,I323637);
nor I_6224 (I107703,I107686,I323631);
nand I_6225 (I107720,I107669,I107703);
not I_6226 (I107542,I107720);
nor I_6227 (I107751,I107621,I323652);
and I_6228 (I107768,I323643,I323640);
nor I_6229 (I107785,I107768,I107621);
nor I_6230 (I107545,I107785,I107720);
nor I_6231 (I107530,I107768,I107703);
nand I_6232 (I107830,I107768,I323652);
not I_6233 (I107847,I107830);
nand I_6234 (I107864,I107703,I107847);
nand I_6235 (I107881,I107652,I107864);
DFFARX1 I_6236 (I107881,I1862,I107553,I107533,);
nand I_6237 (I107539,I107768,I107604);
nand I_6238 (I107536,I107751,I107768);
not I_6239 (I107961,I1869);
and I_6240 (I107978,I292550,I292559);
nor I_6241 (I107995,I107978,I292541);
nand I_6242 (I108012,I292556,I292544);
nor I_6243 (I108029,I108012,I107995);
nor I_6244 (I107935,I108029,I108012);
not I_6245 (I108060,I108029);
not I_6246 (I108077,I108012);
or I_6247 (I108094,I292538,I292541);
nor I_6248 (I108111,I108094,I292538);
nand I_6249 (I108128,I108077,I108111);
not I_6250 (I107950,I108128);
nor I_6251 (I108159,I108029,I292544);
and I_6252 (I108176,I292547,I292553);
nor I_6253 (I108193,I108176,I108029);
nor I_6254 (I107953,I108193,I108128);
nor I_6255 (I107938,I108176,I108111);
nand I_6256 (I108238,I108176,I292544);
not I_6257 (I108255,I108238);
nand I_6258 (I108272,I108111,I108255);
nand I_6259 (I108289,I108060,I108272);
DFFARX1 I_6260 (I108289,I1862,I107961,I107941,);
nand I_6261 (I107947,I108176,I108012);
nand I_6262 (I107944,I108159,I108176);
not I_6263 (I108369,I1869);
and I_6264 (I108386,I192701,I192683);
nor I_6265 (I108403,I108386,I192704);
nand I_6266 (I108420,I192680,I192695);
nor I_6267 (I108437,I108420,I108403);
nor I_6268 (I108343,I108437,I108420);
not I_6269 (I108468,I108437);
not I_6270 (I108485,I108420);
or I_6271 (I108502,I192698,I192680);
nor I_6272 (I108519,I108502,I192686);
nand I_6273 (I108536,I108485,I108519);
not I_6274 (I108358,I108536);
nor I_6275 (I108567,I108437,I192692);
and I_6276 (I108584,I192689,I192683);
nor I_6277 (I108601,I108584,I108437);
nor I_6278 (I108361,I108601,I108536);
nor I_6279 (I108346,I108584,I108519);
nand I_6280 (I108646,I108584,I192692);
not I_6281 (I108663,I108646);
nand I_6282 (I108680,I108519,I108663);
nand I_6283 (I108697,I108468,I108680);
DFFARX1 I_6284 (I108697,I1862,I108369,I108349,);
nand I_6285 (I108355,I108584,I108420);
nand I_6286 (I108352,I108567,I108584);
not I_6287 (I108777,I1869);
and I_6288 (I108794,I235333,I235333);
nor I_6289 (I108811,I108794,I235354);
nand I_6290 (I108828,I235336,I235339);
nor I_6291 (I108845,I108828,I108811);
nor I_6292 (I108751,I108845,I108828);
not I_6293 (I108876,I108845);
not I_6294 (I108893,I108828);
or I_6295 (I108910,I235342,I235351);
nor I_6296 (I108927,I108910,I235348);
nand I_6297 (I108944,I108893,I108927);
not I_6298 (I108766,I108944);
nor I_6299 (I108975,I108845,I235339);
and I_6300 (I108992,I235336,I235345);
nor I_6301 (I109009,I108992,I108845);
nor I_6302 (I108769,I109009,I108944);
nor I_6303 (I108754,I108992,I108927);
nand I_6304 (I109054,I108992,I235339);
not I_6305 (I109071,I109054);
nand I_6306 (I109088,I108927,I109071);
nand I_6307 (I109105,I108876,I109088);
DFFARX1 I_6308 (I109105,I1862,I108777,I108757,);
nand I_6309 (I108763,I108992,I108828);
nand I_6310 (I108760,I108975,I108992);
not I_6311 (I109185,I1869);
and I_6312 (I109202,I101203,I101206);
nor I_6313 (I109219,I109202,I101224);
nand I_6314 (I109236,I101206,I101209);
nor I_6315 (I109253,I109236,I109219);
nor I_6316 (I109159,I109253,I109236);
not I_6317 (I109284,I109253);
not I_6318 (I109301,I109236);
or I_6319 (I109318,I101227,I101218);
nor I_6320 (I109335,I109318,I101203);
nand I_6321 (I109352,I109301,I109335);
not I_6322 (I109174,I109352);
nor I_6323 (I109383,I109253,I101221);
and I_6324 (I109400,I101215,I101212);
nor I_6325 (I109417,I109400,I109253);
nor I_6326 (I109177,I109417,I109352);
nor I_6327 (I109162,I109400,I109335);
nand I_6328 (I109462,I109400,I101221);
not I_6329 (I109479,I109462);
nand I_6330 (I109496,I109335,I109479);
nand I_6331 (I109513,I109284,I109496);
DFFARX1 I_6332 (I109513,I1862,I109185,I109165,);
nand I_6333 (I109171,I109400,I109236);
nand I_6334 (I109168,I109383,I109400);
not I_6335 (I109593,I1869);
and I_6336 (I109610,I87943,I87946);
nor I_6337 (I109627,I109610,I87964);
nand I_6338 (I109644,I87946,I87949);
nor I_6339 (I109661,I109644,I109627);
nor I_6340 (I109567,I109661,I109644);
not I_6341 (I109692,I109661);
not I_6342 (I109709,I109644);
or I_6343 (I109726,I87967,I87958);
nor I_6344 (I109743,I109726,I87943);
nand I_6345 (I109760,I109709,I109743);
not I_6346 (I109582,I109760);
nor I_6347 (I109791,I109661,I87961);
and I_6348 (I109808,I87955,I87952);
nor I_6349 (I109825,I109808,I109661);
nor I_6350 (I109585,I109825,I109760);
nor I_6351 (I109570,I109808,I109743);
nand I_6352 (I109870,I109808,I87961);
not I_6353 (I109887,I109870);
nand I_6354 (I109904,I109743,I109887);
nand I_6355 (I109921,I109692,I109904);
DFFARX1 I_6356 (I109921,I1862,I109593,I109573,);
nand I_6357 (I109579,I109808,I109644);
nand I_6358 (I109576,I109791,I109808);
not I_6359 (I110001,I1869);
and I_6360 (I110018,I356323,I356308);
nor I_6361 (I110035,I110018,I356311);
nand I_6362 (I110052,I356305,I356320);
nor I_6363 (I110069,I110052,I110035);
nor I_6364 (I109975,I110069,I110052);
not I_6365 (I110100,I110069);
not I_6366 (I110117,I110052);
or I_6367 (I110134,I356308,I356311);
nor I_6368 (I110151,I110134,I356305);
nand I_6369 (I110168,I110117,I110151);
not I_6370 (I109990,I110168);
nor I_6371 (I110199,I110069,I356326);
and I_6372 (I110216,I356317,I356314);
nor I_6373 (I110233,I110216,I110069);
nor I_6374 (I109993,I110233,I110168);
nor I_6375 (I109978,I110216,I110151);
nand I_6376 (I110278,I110216,I356326);
not I_6377 (I110295,I110278);
nand I_6378 (I110312,I110151,I110295);
nand I_6379 (I110329,I110100,I110312);
DFFARX1 I_6380 (I110329,I1862,I110001,I109981,);
nand I_6381 (I109987,I110216,I110052);
nand I_6382 (I109984,I110199,I110216);
not I_6383 (I110409,I1869);
and I_6384 (I110426,I195336,I195318);
nor I_6385 (I110443,I110426,I195339);
nand I_6386 (I110460,I195315,I195330);
nor I_6387 (I110477,I110460,I110443);
nor I_6388 (I110383,I110477,I110460);
not I_6389 (I110508,I110477);
not I_6390 (I110525,I110460);
or I_6391 (I110542,I195333,I195315);
nor I_6392 (I110559,I110542,I195321);
nand I_6393 (I110576,I110525,I110559);
not I_6394 (I110398,I110576);
nor I_6395 (I110607,I110477,I195327);
and I_6396 (I110624,I195324,I195318);
nor I_6397 (I110641,I110624,I110477);
nor I_6398 (I110401,I110641,I110576);
nor I_6399 (I110386,I110624,I110559);
nand I_6400 (I110686,I110624,I195327);
not I_6401 (I110703,I110686);
nand I_6402 (I110720,I110559,I110703);
nand I_6403 (I110737,I110508,I110720);
DFFARX1 I_6404 (I110737,I1862,I110409,I110389,);
nand I_6405 (I110395,I110624,I110460);
nand I_6406 (I110392,I110607,I110624);
not I_6407 (I110817,I1869);
and I_6408 (I110834,I171094,I171076);
nor I_6409 (I110851,I110834,I171097);
nand I_6410 (I110868,I171073,I171088);
nor I_6411 (I110885,I110868,I110851);
nor I_6412 (I110791,I110885,I110868);
not I_6413 (I110916,I110885);
not I_6414 (I110933,I110868);
or I_6415 (I110950,I171091,I171073);
nor I_6416 (I110967,I110950,I171079);
nand I_6417 (I110984,I110933,I110967);
not I_6418 (I110806,I110984);
nor I_6419 (I111015,I110885,I171085);
and I_6420 (I111032,I171082,I171076);
nor I_6421 (I111049,I111032,I110885);
nor I_6422 (I110809,I111049,I110984);
nor I_6423 (I110794,I111032,I110967);
nand I_6424 (I111094,I111032,I171085);
not I_6425 (I111111,I111094);
nand I_6426 (I111128,I110967,I111111);
nand I_6427 (I111145,I110916,I111128);
DFFARX1 I_6428 (I111145,I1862,I110817,I110797,);
nand I_6429 (I110803,I111032,I110868);
nand I_6430 (I110800,I111015,I111032);
not I_6431 (I111225,I1869);
and I_6432 (I111242,I311528,I311513);
nor I_6433 (I111259,I111242,I311516);
nand I_6434 (I111276,I311510,I311525);
nor I_6435 (I111293,I111276,I111259);
nor I_6436 (I111199,I111293,I111276);
not I_6437 (I111324,I111293);
not I_6438 (I111341,I111276);
or I_6439 (I111358,I311513,I311516);
nor I_6440 (I111375,I111358,I311510);
nand I_6441 (I111392,I111341,I111375);
not I_6442 (I111214,I111392);
nor I_6443 (I111423,I111293,I311531);
and I_6444 (I111440,I311522,I311519);
nor I_6445 (I111457,I111440,I111293);
nor I_6446 (I111217,I111457,I111392);
nor I_6447 (I111202,I111440,I111375);
nand I_6448 (I111502,I111440,I311531);
not I_6449 (I111519,I111502);
nand I_6450 (I111536,I111375,I111519);
nand I_6451 (I111553,I111324,I111536);
DFFARX1 I_6452 (I111553,I1862,I111225,I111205,);
nand I_6453 (I111211,I111440,I111276);
nand I_6454 (I111208,I111423,I111440);
not I_6455 (I111633,I1869);
and I_6456 (I111650,I78253,I78256);
nor I_6457 (I111667,I111650,I78274);
nand I_6458 (I111684,I78256,I78259);
nor I_6459 (I111701,I111684,I111667);
nor I_6460 (I111607,I111701,I111684);
not I_6461 (I111732,I111701);
not I_6462 (I111749,I111684);
or I_6463 (I111766,I78277,I78268);
nor I_6464 (I111783,I111766,I78253);
nand I_6465 (I111800,I111749,I111783);
not I_6466 (I111622,I111800);
nor I_6467 (I111831,I111701,I78271);
and I_6468 (I111848,I78265,I78262);
nor I_6469 (I111865,I111848,I111701);
nor I_6470 (I111625,I111865,I111800);
nor I_6471 (I111610,I111848,I111783);
nand I_6472 (I111910,I111848,I78271);
not I_6473 (I111927,I111910);
nand I_6474 (I111944,I111783,I111927);
nand I_6475 (I111961,I111732,I111944);
DFFARX1 I_6476 (I111961,I1862,I111633,I111613,);
nand I_6477 (I111619,I111848,I111684);
nand I_6478 (I111616,I111831,I111848);
not I_6479 (I112041,I1869);
and I_6480 (I112058,I145271,I145253);
nor I_6481 (I112075,I112058,I145274);
nand I_6482 (I112092,I145250,I145265);
nor I_6483 (I112109,I112092,I112075);
nor I_6484 (I112015,I112109,I112092);
not I_6485 (I112140,I112109);
not I_6486 (I112157,I112092);
or I_6487 (I112174,I145268,I145250);
nor I_6488 (I112191,I112174,I145256);
nand I_6489 (I112208,I112157,I112191);
not I_6490 (I112030,I112208);
nor I_6491 (I112239,I112109,I145262);
and I_6492 (I112256,I145259,I145253);
nor I_6493 (I112273,I112256,I112109);
nor I_6494 (I112033,I112273,I112208);
nor I_6495 (I112018,I112256,I112191);
nand I_6496 (I112318,I112256,I145262);
not I_6497 (I112335,I112318);
nand I_6498 (I112352,I112191,I112335);
nand I_6499 (I112369,I112140,I112352);
DFFARX1 I_6500 (I112369,I1862,I112041,I112021,);
nand I_6501 (I112027,I112256,I112092);
nand I_6502 (I112024,I112239,I112256);
not I_6503 (I112449,I1869);
and I_6504 (I112466,I137366,I137348);
nor I_6505 (I112483,I112466,I137369);
nand I_6506 (I112500,I137345,I137360);
nor I_6507 (I112517,I112500,I112483);
nor I_6508 (I112423,I112517,I112500);
not I_6509 (I112548,I112517);
not I_6510 (I112565,I112500);
or I_6511 (I112582,I137363,I137345);
nor I_6512 (I112599,I112582,I137351);
nand I_6513 (I112616,I112565,I112599);
not I_6514 (I112438,I112616);
nor I_6515 (I112647,I112517,I137357);
and I_6516 (I112664,I137354,I137348);
nor I_6517 (I112681,I112664,I112517);
nor I_6518 (I112441,I112681,I112616);
nor I_6519 (I112426,I112664,I112599);
nand I_6520 (I112726,I112664,I137357);
not I_6521 (I112743,I112726);
nand I_6522 (I112760,I112599,I112743);
nand I_6523 (I112777,I112548,I112760);
DFFARX1 I_6524 (I112777,I1862,I112449,I112429,);
nand I_6525 (I112435,I112664,I112500);
nand I_6526 (I112432,I112647,I112664);
not I_6527 (I112857,I1869);
and I_6528 (I112874,I395097,I395091);
nor I_6529 (I112891,I112874,I395094);
nand I_6530 (I112908,I395088,I395088);
nor I_6531 (I112925,I112908,I112891);
nor I_6532 (I112831,I112925,I112908);
not I_6533 (I112956,I112925);
not I_6534 (I112973,I112908);
or I_6535 (I112990,I395085,I395082);
nor I_6536 (I113007,I112990,I395085);
nand I_6537 (I113024,I112973,I113007);
not I_6538 (I112846,I113024);
nor I_6539 (I113055,I112925,I395082);
and I_6540 (I113072,I395091,I395100);
nor I_6541 (I113089,I113072,I112925);
nor I_6542 (I112849,I113089,I113024);
nor I_6543 (I112834,I113072,I113007);
nand I_6544 (I113134,I113072,I395082);
not I_6545 (I113151,I113134);
nand I_6546 (I113168,I113007,I113151);
nand I_6547 (I113185,I112956,I113168);
DFFARX1 I_6548 (I113185,I1862,I112857,I112837,);
nand I_6549 (I112843,I113072,I112908);
nand I_6550 (I112840,I113055,I113072);
not I_6551 (I113265,I1869);
and I_6552 (I113282,I125772,I125754);
nor I_6553 (I113299,I113282,I125775);
nand I_6554 (I113316,I125751,I125766);
nor I_6555 (I113333,I113316,I113299);
nor I_6556 (I113239,I113333,I113316);
not I_6557 (I113364,I113333);
not I_6558 (I113381,I113316);
or I_6559 (I113398,I125769,I125751);
nor I_6560 (I113415,I113398,I125757);
nand I_6561 (I113432,I113381,I113415);
not I_6562 (I113254,I113432);
nor I_6563 (I113463,I113333,I125763);
and I_6564 (I113480,I125760,I125754);
nor I_6565 (I113497,I113480,I113333);
nor I_6566 (I113257,I113497,I113432);
nor I_6567 (I113242,I113480,I113415);
nand I_6568 (I113542,I113480,I125763);
not I_6569 (I113559,I113542);
nand I_6570 (I113576,I113415,I113559);
nand I_6571 (I113593,I113364,I113576);
DFFARX1 I_6572 (I113593,I1862,I113265,I113245,);
nand I_6573 (I113251,I113480,I113316);
nand I_6574 (I113248,I113463,I113480);
not I_6575 (I113673,I1869);
and I_6576 (I113690,I93553,I93556);
nor I_6577 (I113707,I113690,I93574);
nand I_6578 (I113724,I93556,I93559);
nor I_6579 (I113741,I113724,I113707);
nor I_6580 (I113647,I113741,I113724);
not I_6581 (I113772,I113741);
not I_6582 (I113789,I113724);
or I_6583 (I113806,I93577,I93568);
nor I_6584 (I113823,I113806,I93553);
nand I_6585 (I113840,I113789,I113823);
not I_6586 (I113662,I113840);
nor I_6587 (I113871,I113741,I93571);
and I_6588 (I113888,I93565,I93562);
nor I_6589 (I113905,I113888,I113741);
nor I_6590 (I113665,I113905,I113840);
nor I_6591 (I113650,I113888,I113823);
nand I_6592 (I113950,I113888,I93571);
not I_6593 (I113967,I113950);
nand I_6594 (I113984,I113823,I113967);
nand I_6595 (I114001,I113772,I113984);
DFFARX1 I_6596 (I114001,I1862,I113673,I113653,);
nand I_6597 (I113659,I113888,I113724);
nand I_6598 (I113656,I113871,I113888);
not I_6599 (I114081,I1869);
and I_6600 (I114098,I366809,I366803);
nor I_6601 (I114115,I114098,I366806);
nand I_6602 (I114132,I366800,I366800);
nor I_6603 (I114149,I114132,I114115);
nor I_6604 (I114055,I114149,I114132);
not I_6605 (I114180,I114149);
not I_6606 (I114197,I114132);
or I_6607 (I114214,I366797,I366794);
nor I_6608 (I114231,I114214,I366797);
nand I_6609 (I114248,I114197,I114231);
not I_6610 (I114070,I114248);
nor I_6611 (I114279,I114149,I366794);
and I_6612 (I114296,I366803,I366812);
nor I_6613 (I114313,I114296,I114149);
nor I_6614 (I114073,I114313,I114248);
nor I_6615 (I114058,I114296,I114231);
nand I_6616 (I114358,I114296,I366794);
not I_6617 (I114375,I114358);
nand I_6618 (I114392,I114231,I114375);
nand I_6619 (I114409,I114180,I114392);
DFFARX1 I_6620 (I114409,I1862,I114081,I114061,);
nand I_6621 (I114067,I114296,I114132);
nand I_6622 (I114064,I114279,I114296);
not I_6623 (I114489,I1869);
and I_6624 (I114506,I253897,I253897);
nor I_6625 (I114523,I114506,I253918);
nand I_6626 (I114540,I253900,I253903);
nor I_6627 (I114557,I114540,I114523);
nor I_6628 (I114463,I114557,I114540);
not I_6629 (I114588,I114557);
not I_6630 (I114605,I114540);
or I_6631 (I114622,I253906,I253915);
nor I_6632 (I114639,I114622,I253912);
nand I_6633 (I114656,I114605,I114639);
not I_6634 (I114478,I114656);
nor I_6635 (I114687,I114557,I253903);
and I_6636 (I114704,I253900,I253909);
nor I_6637 (I114721,I114704,I114557);
nor I_6638 (I114481,I114721,I114656);
nor I_6639 (I114466,I114704,I114639);
nand I_6640 (I114766,I114704,I253903);
not I_6641 (I114783,I114766);
nand I_6642 (I114800,I114639,I114783);
nand I_6643 (I114817,I114588,I114800);
DFFARX1 I_6644 (I114817,I1862,I114489,I114469,);
nand I_6645 (I114475,I114704,I114540);
nand I_6646 (I114472,I114687,I114704);
not I_6647 (I114897,I1869);
and I_6648 (I114914,I249137,I249137);
nor I_6649 (I114931,I114914,I249158);
nand I_6650 (I114948,I249140,I249143);
nor I_6651 (I114965,I114948,I114931);
nor I_6652 (I114871,I114965,I114948);
not I_6653 (I114996,I114965);
not I_6654 (I115013,I114948);
or I_6655 (I115030,I249146,I249155);
nor I_6656 (I115047,I115030,I249152);
nand I_6657 (I115064,I115013,I115047);
not I_6658 (I114886,I115064);
nor I_6659 (I115095,I114965,I249143);
and I_6660 (I115112,I249140,I249149);
nor I_6661 (I115129,I115112,I114965);
nor I_6662 (I114889,I115129,I115064);
nor I_6663 (I114874,I115112,I115047);
nand I_6664 (I115174,I115112,I249143);
not I_6665 (I115191,I115174);
nand I_6666 (I115208,I115047,I115191);
nand I_6667 (I115225,I114996,I115208);
DFFARX1 I_6668 (I115225,I1862,I114897,I114877,);
nand I_6669 (I114883,I115112,I114948);
nand I_6670 (I114880,I115095,I115112);
not I_6671 (I115305,I1869);
and I_6672 (I115322,I137893,I137875);
nor I_6673 (I115339,I115322,I137896);
nand I_6674 (I115356,I137872,I137887);
nor I_6675 (I115373,I115356,I115339);
nor I_6676 (I115279,I115373,I115356);
not I_6677 (I115404,I115373);
not I_6678 (I115421,I115356);
or I_6679 (I115438,I137890,I137872);
nor I_6680 (I115455,I115438,I137878);
nand I_6681 (I115472,I115421,I115455);
not I_6682 (I115294,I115472);
nor I_6683 (I115503,I115373,I137884);
and I_6684 (I115520,I137881,I137875);
nor I_6685 (I115537,I115520,I115373);
nor I_6686 (I115297,I115537,I115472);
nor I_6687 (I115282,I115520,I115455);
nand I_6688 (I115582,I115520,I137884);
not I_6689 (I115599,I115582);
nand I_6690 (I115616,I115455,I115599);
nand I_6691 (I115633,I115404,I115616);
DFFARX1 I_6692 (I115633,I1862,I115305,I115285,);
nand I_6693 (I115291,I115520,I115356);
nand I_6694 (I115288,I115503,I115520);
not I_6695 (I115713,I1869);
and I_6696 (I115730,I719,I1479);
nor I_6697 (I115747,I115730,I1015);
nand I_6698 (I115764,I1199,I783);
nor I_6699 (I115781,I115764,I115747);
nor I_6700 (I115687,I115781,I115764);
not I_6701 (I115812,I115781);
not I_6702 (I115829,I115764);
or I_6703 (I115846,I1775,I1639);
nor I_6704 (I115863,I115846,I1055);
nand I_6705 (I115880,I115829,I115863);
not I_6706 (I115702,I115880);
nor I_6707 (I115911,I115781,I831);
and I_6708 (I115928,I1663,I1007);
nor I_6709 (I115945,I115928,I115781);
nor I_6710 (I115705,I115945,I115880);
nor I_6711 (I115690,I115928,I115863);
nand I_6712 (I115990,I115928,I831);
not I_6713 (I116007,I115990);
nand I_6714 (I116024,I115863,I116007);
nand I_6715 (I116041,I115812,I116024);
DFFARX1 I_6716 (I116041,I1862,I115713,I115693,);
nand I_6717 (I115699,I115928,I115764);
nand I_6718 (I115696,I115911,I115928);
not I_6719 (I116121,I1869);
and I_6720 (I116138,I274365,I274365);
nor I_6721 (I116155,I116138,I274386);
nand I_6722 (I116172,I274368,I274371);
nor I_6723 (I116189,I116172,I116155);
nor I_6724 (I116095,I116189,I116172);
not I_6725 (I116220,I116189);
not I_6726 (I116237,I116172);
or I_6727 (I116254,I274374,I274383);
nor I_6728 (I116271,I116254,I274380);
nand I_6729 (I116288,I116237,I116271);
not I_6730 (I116110,I116288);
nor I_6731 (I116319,I116189,I274371);
and I_6732 (I116336,I274368,I274377);
nor I_6733 (I116353,I116336,I116189);
nor I_6734 (I116113,I116353,I116288);
nor I_6735 (I116098,I116336,I116271);
nand I_6736 (I116398,I116336,I274371);
not I_6737 (I116415,I116398);
nand I_6738 (I116432,I116271,I116415);
nand I_6739 (I116449,I116220,I116432);
DFFARX1 I_6740 (I116449,I1862,I116121,I116101,);
nand I_6741 (I116107,I116336,I116172);
nand I_6742 (I116104,I116319,I116336);
not I_6743 (I116529,I1869);
and I_6744 (I116546,I26743,I26746);
nor I_6745 (I116563,I116546,I26764);
nand I_6746 (I116580,I26746,I26749);
nor I_6747 (I116597,I116580,I116563);
nor I_6748 (I116503,I116597,I116580);
not I_6749 (I116628,I116597);
not I_6750 (I116645,I116580);
or I_6751 (I116662,I26767,I26758);
nor I_6752 (I116679,I116662,I26743);
nand I_6753 (I116696,I116645,I116679);
not I_6754 (I116518,I116696);
nor I_6755 (I116727,I116597,I26761);
and I_6756 (I116744,I26755,I26752);
nor I_6757 (I116761,I116744,I116597);
nor I_6758 (I116521,I116761,I116696);
nor I_6759 (I116506,I116744,I116679);
nand I_6760 (I116806,I116744,I26761);
not I_6761 (I116823,I116806);
nand I_6762 (I116840,I116679,I116823);
nand I_6763 (I116857,I116628,I116840);
DFFARX1 I_6764 (I116857,I1862,I116529,I116509,);
nand I_6765 (I116515,I116744,I116580);
nand I_6766 (I116512,I116727,I116744);
not I_6767 (I116937,I1869);
and I_6768 (I116954,I144744,I144726);
nor I_6769 (I116971,I116954,I144747);
nand I_6770 (I116988,I144723,I144738);
nor I_6771 (I117005,I116988,I116971);
nor I_6772 (I116911,I117005,I116988);
not I_6773 (I117036,I117005);
not I_6774 (I117053,I116988);
or I_6775 (I117070,I144741,I144723);
nor I_6776 (I117087,I117070,I144729);
nand I_6777 (I117104,I117053,I117087);
not I_6778 (I116926,I117104);
nor I_6779 (I117135,I117005,I144735);
and I_6780 (I117152,I144732,I144726);
nor I_6781 (I117169,I117152,I117005);
nor I_6782 (I116929,I117169,I117104);
nor I_6783 (I116914,I117152,I117087);
nand I_6784 (I117214,I117152,I144735);
not I_6785 (I117231,I117214);
nand I_6786 (I117248,I117087,I117231);
nand I_6787 (I117265,I117036,I117248);
DFFARX1 I_6788 (I117265,I1862,I116937,I116917,);
nand I_6789 (I116923,I117152,I116988);
nand I_6790 (I116920,I117135,I117152);
not I_6791 (I117351,I1869);
or I_6792 (I117368,I322595,I322583);
nand I_6793 (I117385,I322577,I322577);
not I_6794 (I117402,I117385);
nand I_6795 (I117419,I117402,I117368);
not I_6796 (I117436,I117419);
nand I_6797 (I117453,I322580,I322580);
and I_6798 (I117470,I117453,I322586);
DFFARX1 I_6799 (I117470,I1862,I117351,I117496,);
nor I_6800 (I117319,I117496,I117385);
nand I_6801 (I117518,I117436,I117496);
nor I_6802 (I117535,I117496,I117402);
not I_6803 (I117337,I117496);
nor I_6804 (I117566,I322592,I322580);
not I_6805 (I117583,I117566);
nand I_6806 (I117340,I117535,I117566);
not I_6807 (I117614,I322598);
nor I_6808 (I117631,I117496,I322598);
nand I_6809 (I117648,I322583,I322589);
nor I_6810 (I117322,I117648,I117385);
not I_6811 (I117679,I117648);
nor I_6812 (I117696,I117566,I117679);
nor I_6813 (I117343,I117696,I117419);
nand I_6814 (I117727,I117679,I117614);
nand I_6815 (I117328,I117436,I117727);
nand I_6816 (I117758,I117518,I117727);
DFFARX1 I_6817 (I117758,I1862,I117351,I117331,);
nand I_6818 (I117789,I117583,I117648);
nor I_6819 (I117325,I117436,I117789);
nor I_6820 (I117820,I117583,I117648);
nand I_6821 (I117334,I117820,I117631);
not I_6822 (I117878,I1869);
or I_6823 (I117895,I363264,I363261);
nand I_6824 (I117912,I363273,I363276);
not I_6825 (I117929,I117912);
nand I_6826 (I117946,I117929,I117895);
not I_6827 (I117963,I117946);
nand I_6828 (I117980,I363267,I363258);
and I_6829 (I117997,I117980,I363258);
DFFARX1 I_6830 (I117997,I1862,I117878,I118023,);
nor I_6831 (I117846,I118023,I117912);
nand I_6832 (I118045,I117963,I118023);
nor I_6833 (I118062,I118023,I117929);
not I_6834 (I117864,I118023);
nor I_6835 (I118093,I363261,I363258);
not I_6836 (I118110,I118093);
nand I_6837 (I117867,I118062,I118093);
not I_6838 (I118141,I363264);
nor I_6839 (I118158,I118023,I363264);
nand I_6840 (I118175,I363267,I363270);
nor I_6841 (I117849,I118175,I117912);
not I_6842 (I118206,I118175);
nor I_6843 (I118223,I118093,I118206);
nor I_6844 (I117870,I118223,I117946);
nand I_6845 (I118254,I118206,I118141);
nand I_6846 (I117855,I117963,I118254);
nand I_6847 (I118285,I118045,I118254);
DFFARX1 I_6848 (I118285,I1862,I117878,I117858,);
nand I_6849 (I118316,I118110,I118175);
nor I_6850 (I117852,I117963,I118316);
nor I_6851 (I118347,I118110,I118175);
nand I_6852 (I117861,I118347,I118158);
not I_6853 (I118405,I1869);
or I_6854 (I118422,I1831,I1511);
nand I_6855 (I118439,I1375,I663);
not I_6856 (I118456,I118439);
nand I_6857 (I118473,I118456,I118422);
not I_6858 (I118490,I118473);
nand I_6859 (I118507,I1159,I815);
and I_6860 (I118524,I118507,I1215);
DFFARX1 I_6861 (I118524,I1862,I118405,I118550,);
nor I_6862 (I118373,I118550,I118439);
nand I_6863 (I118572,I118490,I118550);
nor I_6864 (I118589,I118550,I118456);
not I_6865 (I118391,I118550);
nor I_6866 (I118620,I1735,I815);
not I_6867 (I118637,I118620);
nand I_6868 (I118394,I118589,I118620);
not I_6869 (I118668,I1127);
nor I_6870 (I118685,I118550,I1127);
nand I_6871 (I118702,I1807,I735);
nor I_6872 (I118376,I118702,I118439);
not I_6873 (I118733,I118702);
nor I_6874 (I118750,I118620,I118733);
nor I_6875 (I118397,I118750,I118473);
nand I_6876 (I118781,I118733,I118668);
nand I_6877 (I118382,I118490,I118781);
nand I_6878 (I118812,I118572,I118781);
DFFARX1 I_6879 (I118812,I1862,I118405,I118385,);
nand I_6880 (I118843,I118637,I118702);
nor I_6881 (I118379,I118490,I118843);
nor I_6882 (I118874,I118637,I118702);
nand I_6883 (I118388,I118874,I118685);
not I_6884 (I118932,I1869);
or I_6885 (I118949,I233429,I233432);
nand I_6886 (I118966,I233435,I233444);
not I_6887 (I118983,I118966);
nand I_6888 (I119000,I118983,I118949);
not I_6889 (I119017,I119000);
nand I_6890 (I119034,I233441,I233447);
and I_6891 (I119051,I119034,I233429);
DFFARX1 I_6892 (I119051,I1862,I118932,I119077,);
nor I_6893 (I118900,I119077,I118966);
nand I_6894 (I119099,I119017,I119077);
nor I_6895 (I119116,I119077,I118983);
not I_6896 (I118918,I119077);
nor I_6897 (I119147,I233432,I233447);
not I_6898 (I119164,I119147);
nand I_6899 (I118921,I119116,I119147);
not I_6900 (I119195,I233450);
nor I_6901 (I119212,I119077,I233450);
nand I_6902 (I119229,I233438,I233435);
nor I_6903 (I118903,I119229,I118966);
not I_6904 (I119260,I119229);
nor I_6905 (I119277,I119147,I119260);
nor I_6906 (I118924,I119277,I119000);
nand I_6907 (I119308,I119260,I119195);
nand I_6908 (I118909,I119017,I119308);
nand I_6909 (I119339,I119099,I119308);
DFFARX1 I_6910 (I119339,I1862,I118932,I118912,);
nand I_6911 (I119370,I119164,I119229);
nor I_6912 (I118906,I119017,I119370);
nor I_6913 (I119401,I119164,I119229);
nand I_6914 (I118915,I119401,I119212);
not I_6915 (I119459,I1869);
or I_6916 (I119476,I244377,I244380);
nand I_6917 (I119493,I244383,I244392);
not I_6918 (I119510,I119493);
nand I_6919 (I119527,I119510,I119476);
not I_6920 (I119544,I119527);
nand I_6921 (I119561,I244389,I244395);
and I_6922 (I119578,I119561,I244377);
DFFARX1 I_6923 (I119578,I1862,I119459,I119604,);
nor I_6924 (I119427,I119604,I119493);
nand I_6925 (I119626,I119544,I119604);
nor I_6926 (I119643,I119604,I119510);
not I_6927 (I119445,I119604);
nor I_6928 (I119674,I244380,I244395);
not I_6929 (I119691,I119674);
nand I_6930 (I119448,I119643,I119674);
not I_6931 (I119722,I244398);
nor I_6932 (I119739,I119604,I244398);
nand I_6933 (I119756,I244386,I244383);
nor I_6934 (I119430,I119756,I119493);
not I_6935 (I119787,I119756);
nor I_6936 (I119804,I119674,I119787);
nor I_6937 (I119451,I119804,I119527);
nand I_6938 (I119835,I119787,I119722);
nand I_6939 (I119436,I119544,I119835);
nand I_6940 (I119866,I119626,I119835);
DFFARX1 I_6941 (I119866,I1862,I119459,I119439,);
nand I_6942 (I119897,I119691,I119756);
nor I_6943 (I119433,I119544,I119897);
nor I_6944 (I119928,I119691,I119756);
nand I_6945 (I119442,I119928,I119739);
not I_6946 (I119986,I1869);
or I_6947 (I120003,I348945,I348933);
nand I_6948 (I120020,I348927,I348927);
not I_6949 (I120037,I120020);
nand I_6950 (I120054,I120037,I120003);
not I_6951 (I120071,I120054);
nand I_6952 (I120088,I348930,I348930);
and I_6953 (I120105,I120088,I348936);
DFFARX1 I_6954 (I120105,I1862,I119986,I120131,);
nor I_6955 (I119954,I120131,I120020);
nand I_6956 (I120153,I120071,I120131);
nor I_6957 (I120170,I120131,I120037);
not I_6958 (I119972,I120131);
nor I_6959 (I120201,I348942,I348930);
not I_6960 (I120218,I120201);
nand I_6961 (I119975,I120170,I120201);
not I_6962 (I120249,I348948);
nor I_6963 (I120266,I120131,I348948);
nand I_6964 (I120283,I348933,I348939);
nor I_6965 (I119957,I120283,I120020);
not I_6966 (I120314,I120283);
nor I_6967 (I120331,I120201,I120314);
nor I_6968 (I119978,I120331,I120054);
nand I_6969 (I120362,I120314,I120249);
nand I_6970 (I119963,I120071,I120362);
nand I_6971 (I120393,I120153,I120362);
DFFARX1 I_6972 (I120393,I1862,I119986,I119966,);
nand I_6973 (I120424,I120218,I120283);
nor I_6974 (I119960,I120071,I120424);
nor I_6975 (I120455,I120218,I120283);
nand I_6976 (I119969,I120455,I120266);
not I_6977 (I120513,I1869);
or I_6978 (I120530,I50206,I50203);
nand I_6979 (I120547,I50209,I50206);
not I_6980 (I120564,I120547);
nand I_6981 (I120581,I120564,I120530);
not I_6982 (I120598,I120581);
nand I_6983 (I120615,I50224,I50227);
and I_6984 (I120632,I120615,I50203);
DFFARX1 I_6985 (I120632,I1862,I120513,I120658,);
nor I_6986 (I120481,I120658,I120547);
nand I_6987 (I120680,I120598,I120658);
nor I_6988 (I120697,I120658,I120564);
not I_6989 (I120499,I120658);
nor I_6990 (I120728,I50221,I50227);
not I_6991 (I120745,I120728);
nand I_6992 (I120502,I120697,I120728);
not I_6993 (I120776,I50212);
nor I_6994 (I120793,I120658,I50212);
nand I_6995 (I120810,I50215,I50218);
nor I_6996 (I120484,I120810,I120547);
not I_6997 (I120841,I120810);
nor I_6998 (I120858,I120728,I120841);
nor I_6999 (I120505,I120858,I120581);
nand I_7000 (I120889,I120841,I120776);
nand I_7001 (I120490,I120598,I120889);
nand I_7002 (I120920,I120680,I120889);
DFFARX1 I_7003 (I120920,I1862,I120513,I120493,);
nand I_7004 (I120951,I120745,I120810);
nor I_7005 (I120487,I120598,I120951);
nor I_7006 (I120982,I120745,I120810);
nand I_7007 (I120496,I120982,I120793);
not I_7008 (I121040,I1869);
or I_7009 (I121057,I116509,I116518);
nand I_7010 (I121074,I116512,I116515);
not I_7011 (I121091,I121074);
nand I_7012 (I121108,I121091,I121057);
not I_7013 (I121125,I121108);
nand I_7014 (I121142,I116506,I116506);
and I_7015 (I121159,I121142,I116503);
DFFARX1 I_7016 (I121159,I1862,I121040,I121185,);
nor I_7017 (I121008,I121185,I121074);
nand I_7018 (I121207,I121125,I121185);
nor I_7019 (I121224,I121185,I121091);
not I_7020 (I121026,I121185);
nor I_7021 (I121255,I116521,I116506);
not I_7022 (I121272,I121255);
nand I_7023 (I121029,I121224,I121255);
not I_7024 (I121303,I116509);
nor I_7025 (I121320,I121185,I116509);
nand I_7026 (I121337,I116512,I116503);
nor I_7027 (I121011,I121337,I121074);
not I_7028 (I121368,I121337);
nor I_7029 (I121385,I121255,I121368);
nor I_7030 (I121032,I121385,I121108);
nand I_7031 (I121416,I121368,I121303);
nand I_7032 (I121017,I121125,I121416);
nand I_7033 (I121447,I121207,I121416);
DFFARX1 I_7034 (I121447,I1862,I121040,I121020,);
nand I_7035 (I121478,I121272,I121337);
nor I_7036 (I121014,I121125,I121478);
nor I_7037 (I121509,I121272,I121337);
nand I_7038 (I121023,I121509,I121320);
not I_7039 (I121567,I1869);
or I_7040 (I121584,I203441,I203444);
nand I_7041 (I121601,I203447,I203456);
not I_7042 (I121618,I121601);
nand I_7043 (I121635,I121618,I121584);
not I_7044 (I121652,I121635);
nand I_7045 (I121669,I203453,I203459);
and I_7046 (I121686,I121669,I203441);
DFFARX1 I_7047 (I121686,I1862,I121567,I121712,);
nor I_7048 (I121535,I121712,I121601);
nand I_7049 (I121734,I121652,I121712);
nor I_7050 (I121751,I121712,I121618);
not I_7051 (I121553,I121712);
nor I_7052 (I121782,I203444,I203459);
not I_7053 (I121799,I121782);
nand I_7054 (I121556,I121751,I121782);
not I_7055 (I121830,I203462);
nor I_7056 (I121847,I121712,I203462);
nand I_7057 (I121864,I203450,I203447);
nor I_7058 (I121538,I121864,I121601);
not I_7059 (I121895,I121864);
nor I_7060 (I121912,I121782,I121895);
nor I_7061 (I121559,I121912,I121635);
nand I_7062 (I121943,I121895,I121830);
nand I_7063 (I121544,I121652,I121943);
nand I_7064 (I121974,I121734,I121943);
DFFARX1 I_7065 (I121974,I1862,I121567,I121547,);
nand I_7066 (I122005,I121799,I121864);
nor I_7067 (I121541,I121652,I122005);
nor I_7068 (I122036,I121799,I121864);
nand I_7069 (I121550,I122036,I121847);
not I_7070 (I122094,I1869);
or I_7071 (I122111,I358958,I358946);
nand I_7072 (I122128,I358940,I358940);
not I_7073 (I122145,I122128);
nand I_7074 (I122162,I122145,I122111);
not I_7075 (I122179,I122162);
nand I_7076 (I122196,I358943,I358943);
and I_7077 (I122213,I122196,I358949);
DFFARX1 I_7078 (I122213,I1862,I122094,I122239,);
nor I_7079 (I122062,I122239,I122128);
nand I_7080 (I122261,I122179,I122239);
nor I_7081 (I122278,I122239,I122145);
not I_7082 (I122080,I122239);
nor I_7083 (I122309,I358955,I358943);
not I_7084 (I122326,I122309);
nand I_7085 (I122083,I122278,I122309);
not I_7086 (I122357,I358961);
nor I_7087 (I122374,I122239,I358961);
nand I_7088 (I122391,I358946,I358952);
nor I_7089 (I122065,I122391,I122128);
not I_7090 (I122422,I122391);
nor I_7091 (I122439,I122309,I122422);
nor I_7092 (I122086,I122439,I122162);
nand I_7093 (I122470,I122422,I122357);
nand I_7094 (I122071,I122179,I122470);
nand I_7095 (I122501,I122261,I122470);
DFFARX1 I_7096 (I122501,I1862,I122094,I122074,);
nand I_7097 (I122532,I122326,I122391);
nor I_7098 (I122068,I122179,I122532);
nor I_7099 (I122563,I122326,I122391);
nand I_7100 (I122077,I122563,I122374);
not I_7101 (I122621,I1869);
or I_7102 (I122638,I238665,I238668);
nand I_7103 (I122655,I238671,I238680);
not I_7104 (I122672,I122655);
nand I_7105 (I122689,I122672,I122638);
not I_7106 (I122706,I122689);
nand I_7107 (I122723,I238677,I238683);
and I_7108 (I122740,I122723,I238665);
DFFARX1 I_7109 (I122740,I1862,I122621,I122766,);
nor I_7110 (I122589,I122766,I122655);
nand I_7111 (I122788,I122706,I122766);
nor I_7112 (I122805,I122766,I122672);
not I_7113 (I122607,I122766);
nor I_7114 (I122836,I238668,I238683);
not I_7115 (I122853,I122836);
nand I_7116 (I122610,I122805,I122836);
not I_7117 (I122884,I238686);
nor I_7118 (I122901,I122766,I238686);
nand I_7119 (I122918,I238674,I238671);
nor I_7120 (I122592,I122918,I122655);
not I_7121 (I122949,I122918);
nor I_7122 (I122966,I122836,I122949);
nor I_7123 (I122613,I122966,I122689);
nand I_7124 (I122997,I122949,I122884);
nand I_7125 (I122598,I122706,I122997);
nand I_7126 (I123028,I122788,I122997);
DFFARX1 I_7127 (I123028,I1862,I122621,I122601,);
nand I_7128 (I123059,I122853,I122918);
nor I_7129 (I122595,I122706,I123059);
nor I_7130 (I123090,I122853,I122918);
nand I_7131 (I122604,I123090,I122901);
not I_7132 (I123148,I1869);
or I_7133 (I123165,I355269,I355257);
nand I_7134 (I123182,I355251,I355251);
not I_7135 (I123199,I123182);
nand I_7136 (I123216,I123199,I123165);
not I_7137 (I123233,I123216);
nand I_7138 (I123250,I355254,I355254);
and I_7139 (I123267,I123250,I355260);
DFFARX1 I_7140 (I123267,I1862,I123148,I123293,);
nor I_7141 (I123116,I123293,I123182);
nand I_7142 (I123315,I123233,I123293);
nor I_7143 (I123332,I123293,I123199);
not I_7144 (I123134,I123293);
nor I_7145 (I123363,I355266,I355254);
not I_7146 (I123380,I123363);
nand I_7147 (I123137,I123332,I123363);
not I_7148 (I123411,I355272);
nor I_7149 (I123428,I123293,I355272);
nand I_7150 (I123445,I355257,I355263);
nor I_7151 (I123119,I123445,I123182);
not I_7152 (I123476,I123445);
nor I_7153 (I123493,I123363,I123476);
nor I_7154 (I123140,I123493,I123216);
nand I_7155 (I123524,I123476,I123411);
nand I_7156 (I123125,I123233,I123524);
nand I_7157 (I123555,I123315,I123524);
DFFARX1 I_7158 (I123555,I1862,I123148,I123128,);
nand I_7159 (I123586,I123380,I123445);
nor I_7160 (I123122,I123233,I123586);
nor I_7161 (I123617,I123380,I123445);
nand I_7162 (I123131,I123617,I123428);
not I_7163 (I123675,I1869);
or I_7164 (I123692,I72646,I72643);
nand I_7165 (I123709,I72649,I72646);
not I_7166 (I123726,I123709);
nand I_7167 (I123743,I123726,I123692);
not I_7168 (I123760,I123743);
nand I_7169 (I123777,I72664,I72667);
and I_7170 (I123794,I123777,I72643);
DFFARX1 I_7171 (I123794,I1862,I123675,I123820,);
nor I_7172 (I123643,I123820,I123709);
nand I_7173 (I123842,I123760,I123820);
nor I_7174 (I123859,I123820,I123726);
not I_7175 (I123661,I123820);
nor I_7176 (I123890,I72661,I72667);
not I_7177 (I123907,I123890);
nand I_7178 (I123664,I123859,I123890);
not I_7179 (I123938,I72652);
nor I_7180 (I123955,I123820,I72652);
nand I_7181 (I123972,I72655,I72658);
nor I_7182 (I123646,I123972,I123709);
not I_7183 (I124003,I123972);
nor I_7184 (I124020,I123890,I124003);
nor I_7185 (I123667,I124020,I123743);
nand I_7186 (I124051,I124003,I123938);
nand I_7187 (I123652,I123760,I124051);
nand I_7188 (I124082,I123842,I124051);
DFFARX1 I_7189 (I124082,I1862,I123675,I123655,);
nand I_7190 (I124113,I123907,I123972);
nor I_7191 (I123649,I123760,I124113);
nor I_7192 (I124144,I123907,I123972);
nand I_7193 (I123658,I124144,I123955);
not I_7194 (I124202,I1869);
or I_7195 (I124219,I227717,I227720);
nand I_7196 (I124236,I227723,I227732);
not I_7197 (I124253,I124236);
nand I_7198 (I124270,I124253,I124219);
not I_7199 (I124287,I124270);
nand I_7200 (I124304,I227729,I227735);
and I_7201 (I124321,I124304,I227717);
DFFARX1 I_7202 (I124321,I1862,I124202,I124347,);
nor I_7203 (I124170,I124347,I124236);
nand I_7204 (I124369,I124287,I124347);
nor I_7205 (I124386,I124347,I124253);
not I_7206 (I124188,I124347);
nor I_7207 (I124417,I227720,I227735);
not I_7208 (I124434,I124417);
nand I_7209 (I124191,I124386,I124417);
not I_7210 (I124465,I227738);
nor I_7211 (I124482,I124347,I227738);
nand I_7212 (I124499,I227726,I227723);
nor I_7213 (I124173,I124499,I124236);
not I_7214 (I124530,I124499);
nor I_7215 (I124547,I124417,I124530);
nor I_7216 (I124194,I124547,I124270);
nand I_7217 (I124578,I124530,I124465);
nand I_7218 (I124179,I124287,I124578);
nand I_7219 (I124609,I124369,I124578);
DFFARX1 I_7220 (I124609,I1862,I124202,I124182,);
nand I_7221 (I124640,I124434,I124499);
nor I_7222 (I124176,I124287,I124640);
nor I_7223 (I124671,I124434,I124499);
nand I_7224 (I124185,I124671,I124482);
not I_7225 (I124729,I1869);
or I_7226 (I124746,I5034,I5034);
nand I_7227 (I124763,I5040,I5043);
not I_7228 (I124780,I124763);
nand I_7229 (I124797,I124780,I124746);
not I_7230 (I124814,I124797);
nand I_7231 (I124831,I5052,I5055);
and I_7232 (I124848,I124831,I5037);
DFFARX1 I_7233 (I124848,I1862,I124729,I124874,);
nor I_7234 (I124697,I124874,I124763);
nand I_7235 (I124896,I124814,I124874);
nor I_7236 (I124913,I124874,I124780);
not I_7237 (I124715,I124874);
nor I_7238 (I124944,I5049,I5055);
not I_7239 (I124961,I124944);
nand I_7240 (I124718,I124913,I124944);
not I_7241 (I124992,I5037);
nor I_7242 (I125009,I124874,I5037);
nand I_7243 (I125026,I5040,I5046);
nor I_7244 (I124700,I125026,I124763);
not I_7245 (I125057,I125026);
nor I_7246 (I125074,I124944,I125057);
nor I_7247 (I124721,I125074,I124797);
nand I_7248 (I125105,I125057,I124992);
nand I_7249 (I124706,I124814,I125105);
nand I_7250 (I125136,I124896,I125105);
DFFARX1 I_7251 (I125136,I1862,I124729,I124709,);
nand I_7252 (I125167,I124961,I125026);
nor I_7253 (I124703,I124814,I125167);
nor I_7254 (I125198,I124961,I125026);
nand I_7255 (I124712,I125198,I125009);
not I_7256 (I125256,I1869);
or I_7257 (I125273,I377408,I377405);
nand I_7258 (I125290,I377417,I377420);
not I_7259 (I125307,I125290);
nand I_7260 (I125324,I125307,I125273);
not I_7261 (I125341,I125324);
nand I_7262 (I125358,I377411,I377402);
and I_7263 (I125375,I125358,I377402);
DFFARX1 I_7264 (I125375,I1862,I125256,I125401,);
nor I_7265 (I125224,I125401,I125290);
nand I_7266 (I125423,I125341,I125401);
nor I_7267 (I125440,I125401,I125307);
not I_7268 (I125242,I125401);
nor I_7269 (I125471,I377405,I377402);
not I_7270 (I125488,I125471);
nand I_7271 (I125245,I125440,I125471);
not I_7272 (I125519,I377408);
nor I_7273 (I125536,I125401,I377408);
nand I_7274 (I125553,I377411,I377414);
nor I_7275 (I125227,I125553,I125290);
not I_7276 (I125584,I125553);
nor I_7277 (I125601,I125471,I125584);
nor I_7278 (I125248,I125601,I125324);
nand I_7279 (I125632,I125584,I125519);
nand I_7280 (I125233,I125341,I125632);
nand I_7281 (I125663,I125423,I125632);
DFFARX1 I_7282 (I125663,I1862,I125256,I125236,);
nand I_7283 (I125694,I125488,I125553);
nor I_7284 (I125230,I125341,I125694);
nor I_7285 (I125725,I125488,I125553);
nand I_7286 (I125239,I125725,I125536);
not I_7287 (I125783,I1869);
or I_7288 (I125800,I244853,I244856);
nand I_7289 (I125817,I244859,I244868);
not I_7290 (I125834,I125817);
nand I_7291 (I125851,I125834,I125800);
not I_7292 (I125868,I125851);
nand I_7293 (I125885,I244865,I244871);
and I_7294 (I125902,I125885,I244853);
DFFARX1 I_7295 (I125902,I1862,I125783,I125928,);
nor I_7296 (I125751,I125928,I125817);
nand I_7297 (I125950,I125868,I125928);
nor I_7298 (I125967,I125928,I125834);
not I_7299 (I125769,I125928);
nor I_7300 (I125998,I244856,I244871);
not I_7301 (I126015,I125998);
nand I_7302 (I125772,I125967,I125998);
not I_7303 (I126046,I244874);
nor I_7304 (I126063,I125928,I244874);
nand I_7305 (I126080,I244862,I244859);
nor I_7306 (I125754,I126080,I125817);
not I_7307 (I126111,I126080);
nor I_7308 (I126128,I125998,I126111);
nor I_7309 (I125775,I126128,I125851);
nand I_7310 (I126159,I126111,I126046);
nand I_7311 (I125760,I125868,I126159);
nand I_7312 (I126190,I125950,I126159);
DFFARX1 I_7313 (I126190,I1862,I125783,I125763,);
nand I_7314 (I126221,I126015,I126080);
nor I_7315 (I125757,I125868,I126221);
nor I_7316 (I126252,I126015,I126080);
nand I_7317 (I125766,I126252,I126063);
not I_7318 (I126310,I1869);
or I_7319 (I126327,I32866,I32863);
nand I_7320 (I126344,I32869,I32866);
not I_7321 (I126361,I126344);
nand I_7322 (I126378,I126361,I126327);
not I_7323 (I126395,I126378);
nand I_7324 (I126412,I32884,I32887);
and I_7325 (I126429,I126412,I32863);
DFFARX1 I_7326 (I126429,I1862,I126310,I126455,);
nor I_7327 (I126278,I126455,I126344);
nand I_7328 (I126477,I126395,I126455);
nor I_7329 (I126494,I126455,I126361);
not I_7330 (I126296,I126455);
nor I_7331 (I126525,I32881,I32887);
not I_7332 (I126542,I126525);
nand I_7333 (I126299,I126494,I126525);
not I_7334 (I126573,I32872);
nor I_7335 (I126590,I126455,I32872);
nand I_7336 (I126607,I32875,I32878);
nor I_7337 (I126281,I126607,I126344);
not I_7338 (I126638,I126607);
nor I_7339 (I126655,I126525,I126638);
nor I_7340 (I126302,I126655,I126378);
nand I_7341 (I126686,I126638,I126573);
nand I_7342 (I126287,I126395,I126686);
nand I_7343 (I126717,I126477,I126686);
DFFARX1 I_7344 (I126717,I1862,I126310,I126290,);
nand I_7345 (I126748,I126542,I126607);
nor I_7346 (I126284,I126395,I126748);
nor I_7347 (I126779,I126542,I126607);
nand I_7348 (I126293,I126779,I126590);
not I_7349 (I126837,I1869);
or I_7350 (I126854,I249613,I249616);
nand I_7351 (I126871,I249619,I249628);
not I_7352 (I126888,I126871);
nand I_7353 (I126905,I126888,I126854);
not I_7354 (I126922,I126905);
nand I_7355 (I126939,I249625,I249631);
and I_7356 (I126956,I126939,I249613);
DFFARX1 I_7357 (I126956,I1862,I126837,I126982,);
nor I_7358 (I126805,I126982,I126871);
nand I_7359 (I127004,I126922,I126982);
nor I_7360 (I127021,I126982,I126888);
not I_7361 (I126823,I126982);
nor I_7362 (I127052,I249616,I249631);
not I_7363 (I127069,I127052);
nand I_7364 (I126826,I127021,I127052);
not I_7365 (I127100,I249634);
nor I_7366 (I127117,I126982,I249634);
nand I_7367 (I127134,I249622,I249619);
nor I_7368 (I126808,I127134,I126871);
not I_7369 (I127165,I127134);
nor I_7370 (I127182,I127052,I127165);
nor I_7371 (I126829,I127182,I126905);
nand I_7372 (I127213,I127165,I127100);
nand I_7373 (I126814,I126922,I127213);
nand I_7374 (I127244,I127004,I127213);
DFFARX1 I_7375 (I127244,I1862,I126837,I126817,);
nand I_7376 (I127275,I127069,I127134);
nor I_7377 (I126811,I126922,I127275);
nor I_7378 (I127306,I127069,I127134);
nand I_7379 (I126820,I127306,I127117);
not I_7380 (I127364,I1869);
or I_7381 (I127381,I80806,I80803);
nand I_7382 (I127398,I80809,I80806);
not I_7383 (I127415,I127398);
nand I_7384 (I127432,I127415,I127381);
not I_7385 (I127449,I127432);
nand I_7386 (I127466,I80824,I80827);
and I_7387 (I127483,I127466,I80803);
DFFARX1 I_7388 (I127483,I1862,I127364,I127509,);
nor I_7389 (I127332,I127509,I127398);
nand I_7390 (I127531,I127449,I127509);
nor I_7391 (I127548,I127509,I127415);
not I_7392 (I127350,I127509);
nor I_7393 (I127579,I80821,I80827);
not I_7394 (I127596,I127579);
nand I_7395 (I127353,I127548,I127579);
not I_7396 (I127627,I80812);
nor I_7397 (I127644,I127509,I80812);
nand I_7398 (I127661,I80815,I80818);
nor I_7399 (I127335,I127661,I127398);
not I_7400 (I127692,I127661);
nor I_7401 (I127709,I127579,I127692);
nor I_7402 (I127356,I127709,I127432);
nand I_7403 (I127740,I127692,I127627);
nand I_7404 (I127341,I127449,I127740);
nand I_7405 (I127771,I127531,I127740);
DFFARX1 I_7406 (I127771,I1862,I127364,I127344,);
nand I_7407 (I127802,I127596,I127661);
nor I_7408 (I127338,I127449,I127802);
nor I_7409 (I127833,I127596,I127661);
nand I_7410 (I127347,I127833,I127644);
not I_7411 (I127891,I1869);
or I_7412 (I127908,I383154,I383151);
nand I_7413 (I127925,I383163,I383166);
not I_7414 (I127942,I127925);
nand I_7415 (I127959,I127942,I127908);
not I_7416 (I127976,I127959);
nand I_7417 (I127993,I383157,I383148);
and I_7418 (I128010,I127993,I383148);
DFFARX1 I_7419 (I128010,I1862,I127891,I128036,);
nor I_7420 (I127859,I128036,I127925);
nand I_7421 (I128058,I127976,I128036);
nor I_7422 (I128075,I128036,I127942);
not I_7423 (I127877,I128036);
nor I_7424 (I128106,I383151,I383148);
not I_7425 (I128123,I128106);
nand I_7426 (I127880,I128075,I128106);
not I_7427 (I128154,I383154);
nor I_7428 (I128171,I128036,I383154);
nand I_7429 (I128188,I383157,I383160);
nor I_7430 (I127862,I128188,I127925);
not I_7431 (I128219,I128188);
nor I_7432 (I128236,I128106,I128219);
nor I_7433 (I127883,I128236,I127959);
nand I_7434 (I128267,I128219,I128154);
nand I_7435 (I127868,I127976,I128267);
nand I_7436 (I128298,I128058,I128267);
DFFARX1 I_7437 (I128298,I1862,I127891,I127871,);
nand I_7438 (I128329,I128123,I128188);
nor I_7439 (I127865,I127976,I128329);
nor I_7440 (I128360,I128123,I128188);
nand I_7441 (I127874,I128360,I128171);
not I_7442 (I128418,I1869);
or I_7443 (I128435,I19606,I19603);
nand I_7444 (I128452,I19609,I19606);
not I_7445 (I128469,I128452);
nand I_7446 (I128486,I128469,I128435);
not I_7447 (I128503,I128486);
nand I_7448 (I128520,I19624,I19627);
and I_7449 (I128537,I128520,I19603);
DFFARX1 I_7450 (I128537,I1862,I128418,I128563,);
nor I_7451 (I128386,I128563,I128452);
nand I_7452 (I128585,I128503,I128563);
nor I_7453 (I128602,I128563,I128469);
not I_7454 (I128404,I128563);
nor I_7455 (I128633,I19621,I19627);
not I_7456 (I128650,I128633);
nand I_7457 (I128407,I128602,I128633);
not I_7458 (I128681,I19612);
nor I_7459 (I128698,I128563,I19612);
nand I_7460 (I128715,I19615,I19618);
nor I_7461 (I128389,I128715,I128452);
not I_7462 (I128746,I128715);
nor I_7463 (I128763,I128633,I128746);
nor I_7464 (I128410,I128763,I128486);
nand I_7465 (I128794,I128746,I128681);
nand I_7466 (I128395,I128503,I128794);
nand I_7467 (I128825,I128585,I128794);
DFFARX1 I_7468 (I128825,I1862,I128418,I128398,);
nand I_7469 (I128856,I128650,I128715);
nor I_7470 (I128392,I128503,I128856);
nor I_7471 (I128887,I128650,I128715);
nand I_7472 (I128401,I128887,I128698);
not I_7473 (I128945,I1869);
or I_7474 (I128962,I823,I1519);
nand I_7475 (I128979,I1191,I983);
not I_7476 (I128996,I128979);
nand I_7477 (I129013,I128996,I128962);
not I_7478 (I129030,I129013);
nand I_7479 (I129047,I1463,I927);
and I_7480 (I129064,I129047,I1711);
DFFARX1 I_7481 (I129064,I1862,I128945,I129090,);
nor I_7482 (I128913,I129090,I128979);
nand I_7483 (I129112,I129030,I129090);
nor I_7484 (I129129,I129090,I128996);
not I_7485 (I128931,I129090);
nor I_7486 (I129160,I703,I927);
not I_7487 (I129177,I129160);
nand I_7488 (I128934,I129129,I129160);
not I_7489 (I129208,I1423);
nor I_7490 (I129225,I129090,I1423);
nand I_7491 (I129242,I1599,I1791);
nor I_7492 (I128916,I129242,I128979);
not I_7493 (I129273,I129242);
nor I_7494 (I129290,I129160,I129273);
nor I_7495 (I128937,I129290,I129013);
nand I_7496 (I129321,I129273,I129208);
nand I_7497 (I128922,I129030,I129321);
nand I_7498 (I129352,I129112,I129321);
DFFARX1 I_7499 (I129352,I1862,I128945,I128925,);
nand I_7500 (I129383,I129177,I129242);
nor I_7501 (I128919,I129030,I129383);
nor I_7502 (I129414,I129177,I129242);
nand I_7503 (I128928,I129414,I129225);
not I_7504 (I129472,I1869);
or I_7505 (I129489,I322068,I322056);
nand I_7506 (I129506,I322050,I322050);
not I_7507 (I129523,I129506);
nand I_7508 (I129540,I129523,I129489);
not I_7509 (I129557,I129540);
nand I_7510 (I129574,I322053,I322053);
and I_7511 (I129591,I129574,I322059);
DFFARX1 I_7512 (I129591,I1862,I129472,I129617,);
nor I_7513 (I129440,I129617,I129506);
nand I_7514 (I129639,I129557,I129617);
nor I_7515 (I129656,I129617,I129523);
not I_7516 (I129458,I129617);
nor I_7517 (I129687,I322065,I322053);
not I_7518 (I129704,I129687);
nand I_7519 (I129461,I129656,I129687);
not I_7520 (I129735,I322071);
nor I_7521 (I129752,I129617,I322071);
nand I_7522 (I129769,I322056,I322062);
nor I_7523 (I129443,I129769,I129506);
not I_7524 (I129800,I129769);
nor I_7525 (I129817,I129687,I129800);
nor I_7526 (I129464,I129817,I129540);
nand I_7527 (I129848,I129800,I129735);
nand I_7528 (I129449,I129557,I129848);
nand I_7529 (I129879,I129639,I129848);
DFFARX1 I_7530 (I129879,I1862,I129472,I129452,);
nand I_7531 (I129910,I129704,I129769);
nor I_7532 (I129446,I129557,I129910);
nor I_7533 (I129941,I129704,I129769);
nand I_7534 (I129455,I129941,I129752);
not I_7535 (I129999,I1869);
or I_7536 (I130016,I9777,I9777);
nand I_7537 (I130033,I9783,I9786);
not I_7538 (I130050,I130033);
nand I_7539 (I130067,I130050,I130016);
not I_7540 (I130084,I130067);
nand I_7541 (I130101,I9795,I9798);
and I_7542 (I130118,I130101,I9780);
DFFARX1 I_7543 (I130118,I1862,I129999,I130144,);
nor I_7544 (I129967,I130144,I130033);
nand I_7545 (I130166,I130084,I130144);
nor I_7546 (I130183,I130144,I130050);
not I_7547 (I129985,I130144);
nor I_7548 (I130214,I9792,I9798);
not I_7549 (I130231,I130214);
nand I_7550 (I129988,I130183,I130214);
not I_7551 (I130262,I9780);
nor I_7552 (I130279,I130144,I9780);
nand I_7553 (I130296,I9783,I9789);
nor I_7554 (I129970,I130296,I130033);
not I_7555 (I130327,I130296);
nor I_7556 (I130344,I130214,I130327);
nor I_7557 (I129991,I130344,I130067);
nand I_7558 (I130375,I130327,I130262);
nand I_7559 (I129976,I130084,I130375);
nand I_7560 (I130406,I130166,I130375);
DFFARX1 I_7561 (I130406,I1862,I129999,I129979,);
nand I_7562 (I130437,I130231,I130296);
nor I_7563 (I129973,I130084,I130437);
nor I_7564 (I130468,I130231,I130296);
nand I_7565 (I129982,I130468,I130279);
not I_7566 (I130526,I1869);
or I_7567 (I130543,I93046,I93043);
nand I_7568 (I130560,I93049,I93046);
not I_7569 (I130577,I130560);
nand I_7570 (I130594,I130577,I130543);
not I_7571 (I130611,I130594);
nand I_7572 (I130628,I93064,I93067);
and I_7573 (I130645,I130628,I93043);
DFFARX1 I_7574 (I130645,I1862,I130526,I130671,);
nor I_7575 (I130494,I130671,I130560);
nand I_7576 (I130693,I130611,I130671);
nor I_7577 (I130710,I130671,I130577);
not I_7578 (I130512,I130671);
nor I_7579 (I130741,I93061,I93067);
not I_7580 (I130758,I130741);
nand I_7581 (I130515,I130710,I130741);
not I_7582 (I130789,I93052);
nor I_7583 (I130806,I130671,I93052);
nand I_7584 (I130823,I93055,I93058);
nor I_7585 (I130497,I130823,I130560);
not I_7586 (I130854,I130823);
nor I_7587 (I130871,I130741,I130854);
nor I_7588 (I130518,I130871,I130594);
nand I_7589 (I130902,I130854,I130789);
nand I_7590 (I130503,I130611,I130902);
nand I_7591 (I130933,I130693,I130902);
DFFARX1 I_7592 (I130933,I1862,I130526,I130506,);
nand I_7593 (I130964,I130758,I130823);
nor I_7594 (I130500,I130611,I130964);
nor I_7595 (I130995,I130758,I130823);
nand I_7596 (I130509,I130995,I130806);
not I_7597 (I131053,I1869);
or I_7598 (I131070,I229145,I229148);
nand I_7599 (I131087,I229151,I229160);
not I_7600 (I131104,I131087);
nand I_7601 (I131121,I131104,I131070);
not I_7602 (I131138,I131121);
nand I_7603 (I131155,I229157,I229163);
and I_7604 (I131172,I131155,I229145);
DFFARX1 I_7605 (I131172,I1862,I131053,I131198,);
nor I_7606 (I131021,I131198,I131087);
nand I_7607 (I131220,I131138,I131198);
nor I_7608 (I131237,I131198,I131104);
not I_7609 (I131039,I131198);
nor I_7610 (I131268,I229148,I229163);
not I_7611 (I131285,I131268);
nand I_7612 (I131042,I131237,I131268);
not I_7613 (I131316,I229166);
nor I_7614 (I131333,I131198,I229166);
nand I_7615 (I131350,I229154,I229151);
nor I_7616 (I131024,I131350,I131087);
not I_7617 (I131381,I131350);
nor I_7618 (I131398,I131268,I131381);
nor I_7619 (I131045,I131398,I131121);
nand I_7620 (I131429,I131381,I131316);
nand I_7621 (I131030,I131138,I131429);
nand I_7622 (I131460,I131220,I131429);
DFFARX1 I_7623 (I131460,I1862,I131053,I131033,);
nand I_7624 (I131491,I131285,I131350);
nor I_7625 (I131027,I131138,I131491);
nor I_7626 (I131522,I131285,I131350);
nand I_7627 (I131036,I131522,I131333);
not I_7628 (I131580,I1869);
or I_7629 (I131597,I385806,I385803);
nand I_7630 (I131614,I385815,I385818);
not I_7631 (I131631,I131614);
nand I_7632 (I131648,I131631,I131597);
not I_7633 (I131665,I131648);
nand I_7634 (I131682,I385809,I385800);
and I_7635 (I131699,I131682,I385800);
DFFARX1 I_7636 (I131699,I1862,I131580,I131725,);
nor I_7637 (I131548,I131725,I131614);
nand I_7638 (I131747,I131665,I131725);
nor I_7639 (I131764,I131725,I131631);
not I_7640 (I131566,I131725);
nor I_7641 (I131795,I385803,I385800);
not I_7642 (I131812,I131795);
nand I_7643 (I131569,I131764,I131795);
not I_7644 (I131843,I385806);
nor I_7645 (I131860,I131725,I385806);
nand I_7646 (I131877,I385809,I385812);
nor I_7647 (I131551,I131877,I131614);
not I_7648 (I131908,I131877);
nor I_7649 (I131925,I131795,I131908);
nor I_7650 (I131572,I131925,I131648);
nand I_7651 (I131956,I131908,I131843);
nand I_7652 (I131557,I131665,I131956);
nand I_7653 (I131987,I131747,I131956);
DFFARX1 I_7654 (I131987,I1862,I131580,I131560,);
nand I_7655 (I132018,I131812,I131877);
nor I_7656 (I131554,I131665,I132018);
nor I_7657 (I132049,I131812,I131877);
nand I_7658 (I131563,I132049,I131860);
not I_7659 (I132107,I1869);
or I_7660 (I132124,I334716,I334704);
nand I_7661 (I132141,I334698,I334698);
not I_7662 (I132158,I132141);
nand I_7663 (I132175,I132158,I132124);
not I_7664 (I132192,I132175);
nand I_7665 (I132209,I334701,I334701);
and I_7666 (I132226,I132209,I334707);
DFFARX1 I_7667 (I132226,I1862,I132107,I132252,);
nor I_7668 (I132075,I132252,I132141);
nand I_7669 (I132274,I132192,I132252);
nor I_7670 (I132291,I132252,I132158);
not I_7671 (I132093,I132252);
nor I_7672 (I132322,I334713,I334701);
not I_7673 (I132339,I132322);
nand I_7674 (I132096,I132291,I132322);
not I_7675 (I132370,I334719);
nor I_7676 (I132387,I132252,I334719);
nand I_7677 (I132404,I334704,I334710);
nor I_7678 (I132078,I132404,I132141);
not I_7679 (I132435,I132404);
nor I_7680 (I132452,I132322,I132435);
nor I_7681 (I132099,I132452,I132175);
nand I_7682 (I132483,I132435,I132370);
nand I_7683 (I132084,I132192,I132483);
nand I_7684 (I132514,I132274,I132483);
DFFARX1 I_7685 (I132514,I1862,I132107,I132087,);
nand I_7686 (I132545,I132339,I132404);
nor I_7687 (I132081,I132192,I132545);
nor I_7688 (I132576,I132339,I132404);
nand I_7689 (I132090,I132576,I132387);
not I_7690 (I132634,I1869);
or I_7691 (I132651,I231525,I231528);
nand I_7692 (I132668,I231531,I231540);
not I_7693 (I132685,I132668);
nand I_7694 (I132702,I132685,I132651);
not I_7695 (I132719,I132702);
nand I_7696 (I132736,I231537,I231543);
and I_7697 (I132753,I132736,I231525);
DFFARX1 I_7698 (I132753,I1862,I132634,I132779,);
nor I_7699 (I132602,I132779,I132668);
nand I_7700 (I132801,I132719,I132779);
nor I_7701 (I132818,I132779,I132685);
not I_7702 (I132620,I132779);
nor I_7703 (I132849,I231528,I231543);
not I_7704 (I132866,I132849);
nand I_7705 (I132623,I132818,I132849);
not I_7706 (I132897,I231546);
nor I_7707 (I132914,I132779,I231546);
nand I_7708 (I132931,I231534,I231531);
nor I_7709 (I132605,I132931,I132668);
not I_7710 (I132962,I132931);
nor I_7711 (I132979,I132849,I132962);
nor I_7712 (I132626,I132979,I132702);
nand I_7713 (I133010,I132962,I132897);
nand I_7714 (I132611,I132719,I133010);
nand I_7715 (I133041,I132801,I133010);
DFFARX1 I_7716 (I133041,I1862,I132634,I132614,);
nand I_7717 (I133072,I132866,I132931);
nor I_7718 (I132608,I132719,I133072);
nor I_7719 (I133103,I132866,I132931);
nand I_7720 (I132617,I133103,I132914);
not I_7721 (I133161,I1869);
or I_7722 (I133178,I218197,I218200);
nand I_7723 (I133195,I218203,I218212);
not I_7724 (I133212,I133195);
nand I_7725 (I133229,I133212,I133178);
not I_7726 (I133246,I133229);
nand I_7727 (I133263,I218209,I218215);
and I_7728 (I133280,I133263,I218197);
DFFARX1 I_7729 (I133280,I1862,I133161,I133306,);
nor I_7730 (I133129,I133306,I133195);
nand I_7731 (I133328,I133246,I133306);
nor I_7732 (I133345,I133306,I133212);
not I_7733 (I133147,I133306);
nor I_7734 (I133376,I218200,I218215);
not I_7735 (I133393,I133376);
nand I_7736 (I133150,I133345,I133376);
not I_7737 (I133424,I218218);
nor I_7738 (I133441,I133306,I218218);
nand I_7739 (I133458,I218206,I218203);
nor I_7740 (I133132,I133458,I133195);
not I_7741 (I133489,I133458);
nor I_7742 (I133506,I133376,I133489);
nor I_7743 (I133153,I133506,I133229);
nand I_7744 (I133537,I133489,I133424);
nand I_7745 (I133138,I133246,I133537);
nand I_7746 (I133568,I133328,I133537);
DFFARX1 I_7747 (I133568,I1862,I133161,I133141,);
nand I_7748 (I133599,I133393,I133458);
nor I_7749 (I133135,I133246,I133599);
nor I_7750 (I133630,I133393,I133458);
nand I_7751 (I133144,I133630,I133441);
not I_7752 (I133688,I1869);
or I_7753 (I133705,I212961,I212964);
nand I_7754 (I133722,I212967,I212976);
not I_7755 (I133739,I133722);
nand I_7756 (I133756,I133739,I133705);
not I_7757 (I133773,I133756);
nand I_7758 (I133790,I212973,I212979);
and I_7759 (I133807,I133790,I212961);
DFFARX1 I_7760 (I133807,I1862,I133688,I133833,);
nor I_7761 (I133656,I133833,I133722);
nand I_7762 (I133855,I133773,I133833);
nor I_7763 (I133872,I133833,I133739);
not I_7764 (I133674,I133833);
nor I_7765 (I133903,I212964,I212979);
not I_7766 (I133920,I133903);
nand I_7767 (I133677,I133872,I133903);
not I_7768 (I133951,I212982);
nor I_7769 (I133968,I133833,I212982);
nand I_7770 (I133985,I212970,I212967);
nor I_7771 (I133659,I133985,I133722);
not I_7772 (I134016,I133985);
nor I_7773 (I134033,I133903,I134016);
nor I_7774 (I133680,I134033,I133756);
nand I_7775 (I134064,I134016,I133951);
nand I_7776 (I133665,I133773,I134064);
nand I_7777 (I134095,I133855,I134064);
DFFARX1 I_7778 (I134095,I1862,I133688,I133668,);
nand I_7779 (I134126,I133920,I133985);
nor I_7780 (I133662,I133773,I134126);
nor I_7781 (I134157,I133920,I133985);
nand I_7782 (I133671,I134157,I133968);
not I_7783 (I134215,I1869);
or I_7784 (I134232,I222957,I222960);
nand I_7785 (I134249,I222963,I222972);
not I_7786 (I134266,I134249);
nand I_7787 (I134283,I134266,I134232);
not I_7788 (I134300,I134283);
nand I_7789 (I134317,I222969,I222975);
and I_7790 (I134334,I134317,I222957);
DFFARX1 I_7791 (I134334,I1862,I134215,I134360,);
nor I_7792 (I134183,I134360,I134249);
nand I_7793 (I134382,I134300,I134360);
nor I_7794 (I134399,I134360,I134266);
not I_7795 (I134201,I134360);
nor I_7796 (I134430,I222960,I222975);
not I_7797 (I134447,I134430);
nand I_7798 (I134204,I134399,I134430);
not I_7799 (I134478,I222978);
nor I_7800 (I134495,I134360,I222978);
nand I_7801 (I134512,I222966,I222963);
nor I_7802 (I134186,I134512,I134249);
not I_7803 (I134543,I134512);
nor I_7804 (I134560,I134430,I134543);
nor I_7805 (I134207,I134560,I134283);
nand I_7806 (I134591,I134543,I134478);
nand I_7807 (I134192,I134300,I134591);
nand I_7808 (I134622,I134382,I134591);
DFFARX1 I_7809 (I134622,I1862,I134215,I134195,);
nand I_7810 (I134653,I134447,I134512);
nor I_7811 (I134189,I134300,I134653);
nor I_7812 (I134684,I134447,I134512);
nand I_7813 (I134198,I134684,I134495);
not I_7814 (I134742,I1869);
or I_7815 (I134759,I304677,I304665);
nand I_7816 (I134776,I304659,I304659);
not I_7817 (I134793,I134776);
nand I_7818 (I134810,I134793,I134759);
not I_7819 (I134827,I134810);
nand I_7820 (I134844,I304662,I304662);
and I_7821 (I134861,I134844,I304668);
DFFARX1 I_7822 (I134861,I1862,I134742,I134887,);
nor I_7823 (I134710,I134887,I134776);
nand I_7824 (I134909,I134827,I134887);
nor I_7825 (I134926,I134887,I134793);
not I_7826 (I134728,I134887);
nor I_7827 (I134957,I304674,I304662);
not I_7828 (I134974,I134957);
nand I_7829 (I134731,I134926,I134957);
not I_7830 (I135005,I304680);
nor I_7831 (I135022,I134887,I304680);
nand I_7832 (I135039,I304665,I304671);
nor I_7833 (I134713,I135039,I134776);
not I_7834 (I135070,I135039);
nor I_7835 (I135087,I134957,I135070);
nor I_7836 (I134734,I135087,I134810);
nand I_7837 (I135118,I135070,I135005);
nand I_7838 (I134719,I134827,I135118);
nand I_7839 (I135149,I134909,I135118);
DFFARX1 I_7840 (I135149,I1862,I134742,I134722,);
nand I_7841 (I135180,I134974,I135039);
nor I_7842 (I134716,I134827,I135180);
nor I_7843 (I135211,I134974,I135039);
nand I_7844 (I134725,I135211,I135022);
not I_7845 (I135269,I1869);
or I_7846 (I135286,I92026,I92023);
nand I_7847 (I135303,I92029,I92026);
not I_7848 (I135320,I135303);
nand I_7849 (I135337,I135320,I135286);
not I_7850 (I135354,I135337);
nand I_7851 (I135371,I92044,I92047);
and I_7852 (I135388,I135371,I92023);
DFFARX1 I_7853 (I135388,I1862,I135269,I135414,);
nor I_7854 (I135237,I135414,I135303);
nand I_7855 (I135436,I135354,I135414);
nor I_7856 (I135453,I135414,I135320);
not I_7857 (I135255,I135414);
nor I_7858 (I135484,I92041,I92047);
not I_7859 (I135501,I135484);
nand I_7860 (I135258,I135453,I135484);
not I_7861 (I135532,I92032);
nor I_7862 (I135549,I135414,I92032);
nand I_7863 (I135566,I92035,I92038);
nor I_7864 (I135240,I135566,I135303);
not I_7865 (I135597,I135566);
nor I_7866 (I135614,I135484,I135597);
nor I_7867 (I135261,I135614,I135337);
nand I_7868 (I135645,I135597,I135532);
nand I_7869 (I135246,I135354,I135645);
nand I_7870 (I135676,I135436,I135645);
DFFARX1 I_7871 (I135676,I1862,I135269,I135249,);
nand I_7872 (I135707,I135501,I135566);
nor I_7873 (I135243,I135354,I135707);
nor I_7874 (I135738,I135501,I135566);
nand I_7875 (I135252,I135738,I135549);
not I_7876 (I135796,I1869);
or I_7877 (I135813,I63976,I63973);
nand I_7878 (I135830,I63979,I63976);
not I_7879 (I135847,I135830);
nand I_7880 (I135864,I135847,I135813);
not I_7881 (I135881,I135864);
nand I_7882 (I135898,I63994,I63997);
and I_7883 (I135915,I135898,I63973);
DFFARX1 I_7884 (I135915,I1862,I135796,I135941,);
nor I_7885 (I135764,I135941,I135830);
nand I_7886 (I135963,I135881,I135941);
nor I_7887 (I135980,I135941,I135847);
not I_7888 (I135782,I135941);
nor I_7889 (I136011,I63991,I63997);
not I_7890 (I136028,I136011);
nand I_7891 (I135785,I135980,I136011);
not I_7892 (I136059,I63982);
nor I_7893 (I136076,I135941,I63982);
nand I_7894 (I136093,I63985,I63988);
nor I_7895 (I135767,I136093,I135830);
not I_7896 (I136124,I136093);
nor I_7897 (I136141,I136011,I136124);
nor I_7898 (I135788,I136141,I135864);
nand I_7899 (I136172,I136124,I136059);
nand I_7900 (I135773,I135881,I136172);
nand I_7901 (I136203,I135963,I136172);
DFFARX1 I_7902 (I136203,I1862,I135796,I135776,);
nand I_7903 (I136234,I136028,I136093);
nor I_7904 (I135770,I135881,I136234);
nor I_7905 (I136265,I136028,I136093);
nand I_7906 (I135779,I136265,I136076);
not I_7907 (I136323,I1869);
or I_7908 (I136340,I362380,I362377);
nand I_7909 (I136357,I362389,I362392);
not I_7910 (I136374,I136357);
nand I_7911 (I136391,I136374,I136340);
not I_7912 (I136408,I136391);
nand I_7913 (I136425,I362383,I362374);
and I_7914 (I136442,I136425,I362374);
DFFARX1 I_7915 (I136442,I1862,I136323,I136468,);
nor I_7916 (I136291,I136468,I136357);
nand I_7917 (I136490,I136408,I136468);
nor I_7918 (I136507,I136468,I136374);
not I_7919 (I136309,I136468);
nor I_7920 (I136538,I362377,I362374);
not I_7921 (I136555,I136538);
nand I_7922 (I136312,I136507,I136538);
not I_7923 (I136586,I362380);
nor I_7924 (I136603,I136468,I362380);
nand I_7925 (I136620,I362383,I362386);
nor I_7926 (I136294,I136620,I136357);
not I_7927 (I136651,I136620);
nor I_7928 (I136668,I136538,I136651);
nor I_7929 (I136315,I136668,I136391);
nand I_7930 (I136699,I136651,I136586);
nand I_7931 (I136300,I136408,I136699);
nand I_7932 (I136730,I136490,I136699);
DFFARX1 I_7933 (I136730,I1862,I136323,I136303,);
nand I_7934 (I136761,I136555,I136620);
nor I_7935 (I136297,I136408,I136761);
nor I_7936 (I136792,I136555,I136620);
nand I_7937 (I136306,I136792,I136603);
not I_7938 (I136850,I1869);
or I_7939 (I136867,I406580,I406577);
nand I_7940 (I136884,I406589,I406592);
not I_7941 (I136901,I136884);
nand I_7942 (I136918,I136901,I136867);
not I_7943 (I136935,I136918);
nand I_7944 (I136952,I406583,I406574);
and I_7945 (I136969,I136952,I406574);
DFFARX1 I_7946 (I136969,I1862,I136850,I136995,);
nor I_7947 (I136818,I136995,I136884);
nand I_7948 (I137017,I136935,I136995);
nor I_7949 (I137034,I136995,I136901);
not I_7950 (I136836,I136995);
nor I_7951 (I137065,I406577,I406574);
not I_7952 (I137082,I137065);
nand I_7953 (I136839,I137034,I137065);
not I_7954 (I137113,I406580);
nor I_7955 (I137130,I136995,I406580);
nand I_7956 (I137147,I406583,I406586);
nor I_7957 (I136821,I137147,I136884);
not I_7958 (I137178,I137147);
nor I_7959 (I137195,I137065,I137178);
nor I_7960 (I136842,I137195,I136918);
nand I_7961 (I137226,I137178,I137113);
nand I_7962 (I136827,I136935,I137226);
nand I_7963 (I137257,I137017,I137226);
DFFARX1 I_7964 (I137257,I1862,I136850,I136830,);
nand I_7965 (I137288,I137082,I137147);
nor I_7966 (I136824,I136935,I137288);
nor I_7967 (I137319,I137082,I137147);
nand I_7968 (I136833,I137319,I137130);
not I_7969 (I137377,I1869);
or I_7970 (I137394,I47146,I47143);
nand I_7971 (I137411,I47149,I47146);
not I_7972 (I137428,I137411);
nand I_7973 (I137445,I137428,I137394);
not I_7974 (I137462,I137445);
nand I_7975 (I137479,I47164,I47167);
and I_7976 (I137496,I137479,I47143);
DFFARX1 I_7977 (I137496,I1862,I137377,I137522,);
nor I_7978 (I137345,I137522,I137411);
nand I_7979 (I137544,I137462,I137522);
nor I_7980 (I137561,I137522,I137428);
not I_7981 (I137363,I137522);
nor I_7982 (I137592,I47161,I47167);
not I_7983 (I137609,I137592);
nand I_7984 (I137366,I137561,I137592);
not I_7985 (I137640,I47152);
nor I_7986 (I137657,I137522,I47152);
nand I_7987 (I137674,I47155,I47158);
nor I_7988 (I137348,I137674,I137411);
not I_7989 (I137705,I137674);
nor I_7990 (I137722,I137592,I137705);
nor I_7991 (I137369,I137722,I137445);
nand I_7992 (I137753,I137705,I137640);
nand I_7993 (I137354,I137462,I137753);
nand I_7994 (I137784,I137544,I137753);
DFFARX1 I_7995 (I137784,I1862,I137377,I137357,);
nand I_7996 (I137815,I137609,I137674);
nor I_7997 (I137351,I137462,I137815);
nor I_7998 (I137846,I137609,I137674);
nand I_7999 (I137360,I137846,I137657);
not I_8000 (I137904,I1869);
or I_8001 (I137921,I110797,I110806);
nand I_8002 (I137938,I110800,I110803);
not I_8003 (I137955,I137938);
nand I_8004 (I137972,I137955,I137921);
not I_8005 (I137989,I137972);
nand I_8006 (I138006,I110794,I110794);
and I_8007 (I138023,I138006,I110791);
DFFARX1 I_8008 (I138023,I1862,I137904,I138049,);
nor I_8009 (I137872,I138049,I137938);
nand I_8010 (I138071,I137989,I138049);
nor I_8011 (I138088,I138049,I137955);
not I_8012 (I137890,I138049);
nor I_8013 (I138119,I110809,I110794);
not I_8014 (I138136,I138119);
nand I_8015 (I137893,I138088,I138119);
not I_8016 (I138167,I110797);
nor I_8017 (I138184,I138049,I110797);
nand I_8018 (I138201,I110800,I110791);
nor I_8019 (I137875,I138201,I137938);
not I_8020 (I138232,I138201);
nor I_8021 (I138249,I138119,I138232);
nor I_8022 (I137896,I138249,I137972);
nand I_8023 (I138280,I138232,I138167);
nand I_8024 (I137881,I137989,I138280);
nand I_8025 (I138311,I138071,I138280);
DFFARX1 I_8026 (I138311,I1862,I137904,I137884,);
nand I_8027 (I138342,I138136,I138201);
nor I_8028 (I137878,I137989,I138342);
nor I_8029 (I138373,I138136,I138201);
nand I_8030 (I137887,I138373,I138184);
not I_8031 (I138431,I1869);
or I_8032 (I138448,I43576,I43573);
nand I_8033 (I138465,I43579,I43576);
not I_8034 (I138482,I138465);
nand I_8035 (I138499,I138482,I138448);
not I_8036 (I138516,I138499);
nand I_8037 (I138533,I43594,I43597);
and I_8038 (I138550,I138533,I43573);
DFFARX1 I_8039 (I138550,I1862,I138431,I138576,);
nor I_8040 (I138399,I138576,I138465);
nand I_8041 (I138598,I138516,I138576);
nor I_8042 (I138615,I138576,I138482);
not I_8043 (I138417,I138576);
nor I_8044 (I138646,I43591,I43597);
not I_8045 (I138663,I138646);
nand I_8046 (I138420,I138615,I138646);
not I_8047 (I138694,I43582);
nor I_8048 (I138711,I138576,I43582);
nand I_8049 (I138728,I43585,I43588);
nor I_8050 (I138402,I138728,I138465);
not I_8051 (I138759,I138728);
nor I_8052 (I138776,I138646,I138759);
nor I_8053 (I138423,I138776,I138499);
nand I_8054 (I138807,I138759,I138694);
nand I_8055 (I138408,I138516,I138807);
nand I_8056 (I138838,I138598,I138807);
DFFARX1 I_8057 (I138838,I1862,I138431,I138411,);
nand I_8058 (I138869,I138663,I138728);
nor I_8059 (I138405,I138516,I138869);
nor I_8060 (I138900,I138663,I138728);
nand I_8061 (I138414,I138900,I138711);
not I_8062 (I138958,I1869);
or I_8063 (I138975,I255325,I255328);
nand I_8064 (I138992,I255331,I255340);
not I_8065 (I139009,I138992);
nand I_8066 (I139026,I139009,I138975);
not I_8067 (I139043,I139026);
nand I_8068 (I139060,I255337,I255343);
and I_8069 (I139077,I139060,I255325);
DFFARX1 I_8070 (I139077,I1862,I138958,I139103,);
nor I_8071 (I138926,I139103,I138992);
nand I_8072 (I139125,I139043,I139103);
nor I_8073 (I139142,I139103,I139009);
not I_8074 (I138944,I139103);
nor I_8075 (I139173,I255328,I255343);
not I_8076 (I139190,I139173);
nand I_8077 (I138947,I139142,I139173);
not I_8078 (I139221,I255346);
nor I_8079 (I139238,I139103,I255346);
nand I_8080 (I139255,I255334,I255331);
nor I_8081 (I138929,I139255,I138992);
not I_8082 (I139286,I139255);
nor I_8083 (I139303,I139173,I139286);
nor I_8084 (I138950,I139303,I139026);
nand I_8085 (I139334,I139286,I139221);
nand I_8086 (I138935,I139043,I139334);
nand I_8087 (I139365,I139125,I139334);
DFFARX1 I_8088 (I139365,I1862,I138958,I138938,);
nand I_8089 (I139396,I139190,I139255);
nor I_8090 (I138932,I139043,I139396);
nor I_8091 (I139427,I139190,I139255);
nand I_8092 (I138941,I139427,I139238);
not I_8093 (I139485,I1869);
or I_8094 (I139502,I205345,I205348);
nand I_8095 (I139519,I205351,I205360);
not I_8096 (I139536,I139519);
nand I_8097 (I139553,I139536,I139502);
not I_8098 (I139570,I139553);
nand I_8099 (I139587,I205357,I205363);
and I_8100 (I139604,I139587,I205345);
DFFARX1 I_8101 (I139604,I1862,I139485,I139630,);
nor I_8102 (I139453,I139630,I139519);
nand I_8103 (I139652,I139570,I139630);
nor I_8104 (I139669,I139630,I139536);
not I_8105 (I139471,I139630);
nor I_8106 (I139700,I205348,I205363);
not I_8107 (I139717,I139700);
nand I_8108 (I139474,I139669,I139700);
not I_8109 (I139748,I205366);
nor I_8110 (I139765,I139630,I205366);
nand I_8111 (I139782,I205354,I205351);
nor I_8112 (I139456,I139782,I139519);
not I_8113 (I139813,I139782);
nor I_8114 (I139830,I139700,I139813);
nor I_8115 (I139477,I139830,I139553);
nand I_8116 (I139861,I139813,I139748);
nand I_8117 (I139462,I139570,I139861);
nand I_8118 (I139892,I139652,I139861);
DFFARX1 I_8119 (I139892,I1862,I139485,I139465,);
nand I_8120 (I139923,I139717,I139782);
nor I_8121 (I139459,I139570,I139923);
nor I_8122 (I139954,I139717,I139782);
nand I_8123 (I139468,I139954,I139765);
not I_8124 (I140012,I1869);
or I_8125 (I140029,I22156,I22153);
nand I_8126 (I140046,I22159,I22156);
not I_8127 (I140063,I140046);
nand I_8128 (I140080,I140063,I140029);
not I_8129 (I140097,I140080);
nand I_8130 (I140114,I22174,I22177);
and I_8131 (I140131,I140114,I22153);
DFFARX1 I_8132 (I140131,I1862,I140012,I140157,);
nor I_8133 (I139980,I140157,I140046);
nand I_8134 (I140179,I140097,I140157);
nor I_8135 (I140196,I140157,I140063);
not I_8136 (I139998,I140157);
nor I_8137 (I140227,I22171,I22177);
not I_8138 (I140244,I140227);
nand I_8139 (I140001,I140196,I140227);
not I_8140 (I140275,I22162);
nor I_8141 (I140292,I140157,I22162);
nand I_8142 (I140309,I22165,I22168);
nor I_8143 (I139983,I140309,I140046);
not I_8144 (I140340,I140309);
nor I_8145 (I140357,I140227,I140340);
nor I_8146 (I140004,I140357,I140080);
nand I_8147 (I140388,I140340,I140275);
nand I_8148 (I139989,I140097,I140388);
nand I_8149 (I140419,I140179,I140388);
DFFARX1 I_8150 (I140419,I1862,I140012,I139992,);
nand I_8151 (I140450,I140244,I140309);
nor I_8152 (I139986,I140097,I140450);
nor I_8153 (I140481,I140244,I140309);
nand I_8154 (I139995,I140481,I140292);
not I_8155 (I140539,I1869);
or I_8156 (I140556,I60406,I60403);
nand I_8157 (I140573,I60409,I60406);
not I_8158 (I140590,I140573);
nand I_8159 (I140607,I140590,I140556);
not I_8160 (I140624,I140607);
nand I_8161 (I140641,I60424,I60427);
and I_8162 (I140658,I140641,I60403);
DFFARX1 I_8163 (I140658,I1862,I140539,I140684,);
nor I_8164 (I140507,I140684,I140573);
nand I_8165 (I140706,I140624,I140684);
nor I_8166 (I140723,I140684,I140590);
not I_8167 (I140525,I140684);
nor I_8168 (I140754,I60421,I60427);
not I_8169 (I140771,I140754);
nand I_8170 (I140528,I140723,I140754);
not I_8171 (I140802,I60412);
nor I_8172 (I140819,I140684,I60412);
nand I_8173 (I140836,I60415,I60418);
nor I_8174 (I140510,I140836,I140573);
not I_8175 (I140867,I140836);
nor I_8176 (I140884,I140754,I140867);
nor I_8177 (I140531,I140884,I140607);
nand I_8178 (I140915,I140867,I140802);
nand I_8179 (I140516,I140624,I140915);
nand I_8180 (I140946,I140706,I140915);
DFFARX1 I_8181 (I140946,I1862,I140539,I140519,);
nand I_8182 (I140977,I140771,I140836);
nor I_8183 (I140513,I140624,I140977);
nor I_8184 (I141008,I140771,I140836);
nand I_8185 (I140522,I141008,I140819);
not I_8186 (I141066,I1869);
or I_8187 (I141083,I294140,I294128);
nand I_8188 (I141100,I294131,I294125);
not I_8189 (I141117,I141100);
nand I_8190 (I141134,I141117,I141083);
not I_8191 (I141151,I141134);
nand I_8192 (I141168,I294122,I294125);
and I_8193 (I141185,I141168,I294119);
DFFARX1 I_8194 (I141185,I1862,I141066,I141211,);
nor I_8195 (I141034,I141211,I141100);
nand I_8196 (I141233,I141151,I141211);
nor I_8197 (I141250,I141211,I141117);
not I_8198 (I141052,I141211);
nor I_8199 (I141281,I294119,I294125);
not I_8200 (I141298,I141281);
nand I_8201 (I141055,I141250,I141281);
not I_8202 (I141329,I294122);
nor I_8203 (I141346,I141211,I294122);
nand I_8204 (I141363,I294137,I294134);
nor I_8205 (I141037,I141363,I141100);
not I_8206 (I141394,I141363);
nor I_8207 (I141411,I141281,I141394);
nor I_8208 (I141058,I141411,I141134);
nand I_8209 (I141442,I141394,I141329);
nand I_8210 (I141043,I141151,I141442);
nand I_8211 (I141473,I141233,I141442);
DFFARX1 I_8212 (I141473,I1862,I141066,I141046,);
nand I_8213 (I141504,I141298,I141363);
nor I_8214 (I141040,I141151,I141504);
nor I_8215 (I141535,I141298,I141363);
nand I_8216 (I141049,I141535,I141346);
not I_8217 (I141593,I1869);
or I_8218 (I141610,I227241,I227244);
nand I_8219 (I141627,I227247,I227256);
not I_8220 (I141644,I141627);
nand I_8221 (I141661,I141644,I141610);
not I_8222 (I141678,I141661);
nand I_8223 (I141695,I227253,I227259);
and I_8224 (I141712,I141695,I227241);
DFFARX1 I_8225 (I141712,I1862,I141593,I141738,);
nor I_8226 (I141561,I141738,I141627);
nand I_8227 (I141760,I141678,I141738);
nor I_8228 (I141777,I141738,I141644);
not I_8229 (I141579,I141738);
nor I_8230 (I141808,I227244,I227259);
not I_8231 (I141825,I141808);
nand I_8232 (I141582,I141777,I141808);
not I_8233 (I141856,I227262);
nor I_8234 (I141873,I141738,I227262);
nand I_8235 (I141890,I227250,I227247);
nor I_8236 (I141564,I141890,I141627);
not I_8237 (I141921,I141890);
nor I_8238 (I141938,I141808,I141921);
nor I_8239 (I141585,I141938,I141661);
nand I_8240 (I141969,I141921,I141856);
nand I_8241 (I141570,I141678,I141969);
nand I_8242 (I142000,I141760,I141969);
DFFARX1 I_8243 (I142000,I1862,I141593,I141573,);
nand I_8244 (I142031,I141825,I141890);
nor I_8245 (I141567,I141678,I142031);
nor I_8246 (I142062,I141825,I141890);
nand I_8247 (I141576,I142062,I141873);
not I_8248 (I142120,I1869);
or I_8249 (I142137,I309947,I309935);
nand I_8250 (I142154,I309929,I309929);
not I_8251 (I142171,I142154);
nand I_8252 (I142188,I142171,I142137);
not I_8253 (I142205,I142188);
nand I_8254 (I142222,I309932,I309932);
and I_8255 (I142239,I142222,I309938);
DFFARX1 I_8256 (I142239,I1862,I142120,I142265,);
nor I_8257 (I142088,I142265,I142154);
nand I_8258 (I142287,I142205,I142265);
nor I_8259 (I142304,I142265,I142171);
not I_8260 (I142106,I142265);
nor I_8261 (I142335,I309944,I309932);
not I_8262 (I142352,I142335);
nand I_8263 (I142109,I142304,I142335);
not I_8264 (I142383,I309950);
nor I_8265 (I142400,I142265,I309950);
nand I_8266 (I142417,I309935,I309941);
nor I_8267 (I142091,I142417,I142154);
not I_8268 (I142448,I142417);
nor I_8269 (I142465,I142335,I142448);
nor I_8270 (I142112,I142465,I142188);
nand I_8271 (I142496,I142448,I142383);
nand I_8272 (I142097,I142205,I142496);
nand I_8273 (I142527,I142287,I142496);
DFFARX1 I_8274 (I142527,I1862,I142120,I142100,);
nand I_8275 (I142558,I142352,I142417);
nor I_8276 (I142094,I142205,I142558);
nor I_8277 (I142589,I142352,I142417);
nand I_8278 (I142103,I142589,I142400);
not I_8279 (I142647,I1869);
or I_8280 (I142664,I56836,I56833);
nand I_8281 (I142681,I56839,I56836);
not I_8282 (I142698,I142681);
nand I_8283 (I142715,I142698,I142664);
not I_8284 (I142732,I142715);
nand I_8285 (I142749,I56854,I56857);
and I_8286 (I142766,I142749,I56833);
DFFARX1 I_8287 (I142766,I1862,I142647,I142792,);
nor I_8288 (I142615,I142792,I142681);
nand I_8289 (I142814,I142732,I142792);
nor I_8290 (I142831,I142792,I142698);
not I_8291 (I142633,I142792);
nor I_8292 (I142862,I56851,I56857);
not I_8293 (I142879,I142862);
nand I_8294 (I142636,I142831,I142862);
not I_8295 (I142910,I56842);
nor I_8296 (I142927,I142792,I56842);
nand I_8297 (I142944,I56845,I56848);
nor I_8298 (I142618,I142944,I142681);
not I_8299 (I142975,I142944);
nor I_8300 (I142992,I142862,I142975);
nor I_8301 (I142639,I142992,I142715);
nand I_8302 (I143023,I142975,I142910);
nand I_8303 (I142624,I142732,I143023);
nand I_8304 (I143054,I142814,I143023);
DFFARX1 I_8305 (I143054,I1862,I142647,I142627,);
nand I_8306 (I143085,I142879,I142944);
nor I_8307 (I142621,I142732,I143085);
nor I_8308 (I143116,I142879,I142944);
nand I_8309 (I142630,I143116,I142927);
not I_8310 (I143174,I1869);
or I_8311 (I143191,I6615,I6615);
nand I_8312 (I143208,I6621,I6624);
not I_8313 (I143225,I143208);
nand I_8314 (I143242,I143225,I143191);
not I_8315 (I143259,I143242);
nand I_8316 (I143276,I6633,I6636);
and I_8317 (I143293,I143276,I6618);
DFFARX1 I_8318 (I143293,I1862,I143174,I143319,);
nor I_8319 (I143142,I143319,I143208);
nand I_8320 (I143341,I143259,I143319);
nor I_8321 (I143358,I143319,I143225);
not I_8322 (I143160,I143319);
nor I_8323 (I143389,I6630,I6636);
not I_8324 (I143406,I143389);
nand I_8325 (I143163,I143358,I143389);
not I_8326 (I143437,I6618);
nor I_8327 (I143454,I143319,I6618);
nand I_8328 (I143471,I6621,I6627);
nor I_8329 (I143145,I143471,I143208);
not I_8330 (I143502,I143471);
nor I_8331 (I143519,I143389,I143502);
nor I_8332 (I143166,I143519,I143242);
nand I_8333 (I143550,I143502,I143437);
nand I_8334 (I143151,I143259,I143550);
nand I_8335 (I143581,I143341,I143550);
DFFARX1 I_8336 (I143581,I1862,I143174,I143154,);
nand I_8337 (I143612,I143406,I143471);
nor I_8338 (I143148,I143259,I143612);
nor I_8339 (I143643,I143406,I143471);
nand I_8340 (I143157,I143643,I143454);
not I_8341 (I143701,I1869);
or I_8342 (I143718,I54796,I54793);
nand I_8343 (I143735,I54799,I54796);
not I_8344 (I143752,I143735);
nand I_8345 (I143769,I143752,I143718);
not I_8346 (I143786,I143769);
nand I_8347 (I143803,I54814,I54817);
and I_8348 (I143820,I143803,I54793);
DFFARX1 I_8349 (I143820,I1862,I143701,I143846,);
nor I_8350 (I143669,I143846,I143735);
nand I_8351 (I143868,I143786,I143846);
nor I_8352 (I143885,I143846,I143752);
not I_8353 (I143687,I143846);
nor I_8354 (I143916,I54811,I54817);
not I_8355 (I143933,I143916);
nand I_8356 (I143690,I143885,I143916);
not I_8357 (I143964,I54802);
nor I_8358 (I143981,I143846,I54802);
nand I_8359 (I143998,I54805,I54808);
nor I_8360 (I143672,I143998,I143735);
not I_8361 (I144029,I143998);
nor I_8362 (I144046,I143916,I144029);
nor I_8363 (I143693,I144046,I143769);
nand I_8364 (I144077,I144029,I143964);
nand I_8365 (I143678,I143786,I144077);
nand I_8366 (I144108,I143868,I144077);
DFFARX1 I_8367 (I144108,I1862,I143701,I143681,);
nand I_8368 (I144139,I143933,I143998);
nor I_8369 (I143675,I143786,I144139);
nor I_8370 (I144170,I143933,I143998);
nand I_8371 (I143684,I144170,I143981);
not I_8372 (I144228,I1869);
or I_8373 (I144245,I353688,I353676);
nand I_8374 (I144262,I353670,I353670);
not I_8375 (I144279,I144262);
nand I_8376 (I144296,I144279,I144245);
not I_8377 (I144313,I144296);
nand I_8378 (I144330,I353673,I353673);
and I_8379 (I144347,I144330,I353679);
DFFARX1 I_8380 (I144347,I1862,I144228,I144373,);
nor I_8381 (I144196,I144373,I144262);
nand I_8382 (I144395,I144313,I144373);
nor I_8383 (I144412,I144373,I144279);
not I_8384 (I144214,I144373);
nor I_8385 (I144443,I353685,I353673);
not I_8386 (I144460,I144443);
nand I_8387 (I144217,I144412,I144443);
not I_8388 (I144491,I353691);
nor I_8389 (I144508,I144373,I353691);
nand I_8390 (I144525,I353676,I353682);
nor I_8391 (I144199,I144525,I144262);
not I_8392 (I144556,I144525);
nor I_8393 (I144573,I144443,I144556);
nor I_8394 (I144220,I144573,I144296);
nand I_8395 (I144604,I144556,I144491);
nand I_8396 (I144205,I144313,I144604);
nand I_8397 (I144635,I144395,I144604);
DFFARX1 I_8398 (I144635,I1862,I144228,I144208,);
nand I_8399 (I144666,I144460,I144525);
nor I_8400 (I144202,I144313,I144666);
nor I_8401 (I144697,I144460,I144525);
nand I_8402 (I144211,I144697,I144508);
not I_8403 (I144755,I1869);
or I_8404 (I144772,I204869,I204872);
nand I_8405 (I144789,I204875,I204884);
not I_8406 (I144806,I144789);
nand I_8407 (I144823,I144806,I144772);
not I_8408 (I144840,I144823);
nand I_8409 (I144857,I204881,I204887);
and I_8410 (I144874,I144857,I204869);
DFFARX1 I_8411 (I144874,I1862,I144755,I144900,);
nor I_8412 (I144723,I144900,I144789);
nand I_8413 (I144922,I144840,I144900);
nor I_8414 (I144939,I144900,I144806);
not I_8415 (I144741,I144900);
nor I_8416 (I144970,I204872,I204887);
not I_8417 (I144987,I144970);
nand I_8418 (I144744,I144939,I144970);
not I_8419 (I145018,I204890);
nor I_8420 (I145035,I144900,I204890);
nand I_8421 (I145052,I204878,I204875);
nor I_8422 (I144726,I145052,I144789);
not I_8423 (I145083,I145052);
nor I_8424 (I145100,I144970,I145083);
nor I_8425 (I144747,I145100,I144823);
nand I_8426 (I145131,I145083,I145018);
nand I_8427 (I144732,I144840,I145131);
nand I_8428 (I145162,I144922,I145131);
DFFARX1 I_8429 (I145162,I1862,I144755,I144735,);
nand I_8430 (I145193,I144987,I145052);
nor I_8431 (I144729,I144840,I145193);
nor I_8432 (I145224,I144987,I145052);
nand I_8433 (I144738,I145224,I145035);
not I_8434 (I145282,I1869);
or I_8435 (I145299,I282933,I282936);
nand I_8436 (I145316,I282939,I282948);
not I_8437 (I145333,I145316);
nand I_8438 (I145350,I145333,I145299);
not I_8439 (I145367,I145350);
nand I_8440 (I145384,I282945,I282951);
and I_8441 (I145401,I145384,I282933);
DFFARX1 I_8442 (I145401,I1862,I145282,I145427,);
nor I_8443 (I145250,I145427,I145316);
nand I_8444 (I145449,I145367,I145427);
nor I_8445 (I145466,I145427,I145333);
not I_8446 (I145268,I145427);
nor I_8447 (I145497,I282936,I282951);
not I_8448 (I145514,I145497);
nand I_8449 (I145271,I145466,I145497);
not I_8450 (I145545,I282954);
nor I_8451 (I145562,I145427,I282954);
nand I_8452 (I145579,I282942,I282939);
nor I_8453 (I145253,I145579,I145316);
not I_8454 (I145610,I145579);
nor I_8455 (I145627,I145497,I145610);
nor I_8456 (I145274,I145627,I145350);
nand I_8457 (I145658,I145610,I145545);
nand I_8458 (I145259,I145367,I145658);
nand I_8459 (I145689,I145449,I145658);
DFFARX1 I_8460 (I145689,I1862,I145282,I145262,);
nand I_8461 (I145720,I145514,I145579);
nor I_8462 (I145256,I145367,I145720);
nor I_8463 (I145751,I145514,I145579);
nand I_8464 (I145265,I145751,I145562);
not I_8465 (I145809,I1869);
or I_8466 (I145826,I299410,I299398);
nand I_8467 (I145843,I299401,I299395);
not I_8468 (I145860,I145843);
nand I_8469 (I145877,I145860,I145826);
not I_8470 (I145894,I145877);
nand I_8471 (I145911,I299392,I299395);
and I_8472 (I145928,I145911,I299389);
DFFARX1 I_8473 (I145928,I1862,I145809,I145954,);
nor I_8474 (I145777,I145954,I145843);
nand I_8475 (I145976,I145894,I145954);
nor I_8476 (I145993,I145954,I145860);
not I_8477 (I145795,I145954);
nor I_8478 (I146024,I299389,I299395);
not I_8479 (I146041,I146024);
nand I_8480 (I145798,I145993,I146024);
not I_8481 (I146072,I299392);
nor I_8482 (I146089,I145954,I299392);
nand I_8483 (I146106,I299407,I299404);
nor I_8484 (I145780,I146106,I145843);
not I_8485 (I146137,I146106);
nor I_8486 (I146154,I146024,I146137);
nor I_8487 (I145801,I146154,I145877);
nand I_8488 (I146185,I146137,I146072);
nand I_8489 (I145786,I145894,I146185);
nand I_8490 (I146216,I145976,I146185);
DFFARX1 I_8491 (I146216,I1862,I145809,I145789,);
nand I_8492 (I146247,I146041,I146106);
nor I_8493 (I145783,I145894,I146247);
nor I_8494 (I146278,I146041,I146106);
nand I_8495 (I145792,I146278,I146089);
not I_8496 (I146336,I1869);
or I_8497 (I146353,I88966,I88963);
nand I_8498 (I146370,I88969,I88966);
not I_8499 (I146387,I146370);
nand I_8500 (I146404,I146387,I146353);
not I_8501 (I146421,I146404);
nand I_8502 (I146438,I88984,I88987);
and I_8503 (I146455,I146438,I88963);
DFFARX1 I_8504 (I146455,I1862,I146336,I146481,);
nor I_8505 (I146304,I146481,I146370);
nand I_8506 (I146503,I146421,I146481);
nor I_8507 (I146520,I146481,I146387);
not I_8508 (I146322,I146481);
nor I_8509 (I146551,I88981,I88987);
not I_8510 (I146568,I146551);
nand I_8511 (I146325,I146520,I146551);
not I_8512 (I146599,I88972);
nor I_8513 (I146616,I146481,I88972);
nand I_8514 (I146633,I88975,I88978);
nor I_8515 (I146307,I146633,I146370);
not I_8516 (I146664,I146633);
nor I_8517 (I146681,I146551,I146664);
nor I_8518 (I146328,I146681,I146404);
nand I_8519 (I146712,I146664,I146599);
nand I_8520 (I146313,I146421,I146712);
nand I_8521 (I146743,I146503,I146712);
DFFARX1 I_8522 (I146743,I1862,I146336,I146316,);
nand I_8523 (I146774,I146568,I146633);
nor I_8524 (I146310,I146421,I146774);
nor I_8525 (I146805,I146568,I146633);
nand I_8526 (I146319,I146805,I146616);
not I_8527 (I146863,I1869);
or I_8528 (I146880,I258657,I258660);
nand I_8529 (I146897,I258663,I258672);
not I_8530 (I146914,I146897);
nand I_8531 (I146931,I146914,I146880);
not I_8532 (I146948,I146931);
nand I_8533 (I146965,I258669,I258675);
and I_8534 (I146982,I146965,I258657);
DFFARX1 I_8535 (I146982,I1862,I146863,I147008,);
nor I_8536 (I146831,I147008,I146897);
nand I_8537 (I147030,I146948,I147008);
nor I_8538 (I147047,I147008,I146914);
not I_8539 (I146849,I147008);
nor I_8540 (I147078,I258660,I258675);
not I_8541 (I147095,I147078);
nand I_8542 (I146852,I147047,I147078);
not I_8543 (I147126,I258678);
nor I_8544 (I147143,I147008,I258678);
nand I_8545 (I147160,I258666,I258663);
nor I_8546 (I146834,I147160,I146897);
not I_8547 (I147191,I147160);
nor I_8548 (I147208,I147078,I147191);
nor I_8549 (I146855,I147208,I146931);
nand I_8550 (I147239,I147191,I147126);
nand I_8551 (I146840,I146948,I147239);
nand I_8552 (I147270,I147030,I147239);
DFFARX1 I_8553 (I147270,I1862,I146863,I146843,);
nand I_8554 (I147301,I147095,I147160);
nor I_8555 (I146837,I146948,I147301);
nor I_8556 (I147332,I147095,I147160);
nand I_8557 (I146846,I147332,I147143);
not I_8558 (I147390,I1869);
or I_8559 (I147407,I87436,I87433);
nand I_8560 (I147424,I87439,I87436);
not I_8561 (I147441,I147424);
nand I_8562 (I147458,I147441,I147407);
not I_8563 (I147475,I147458);
nand I_8564 (I147492,I87454,I87457);
and I_8565 (I147509,I147492,I87433);
DFFARX1 I_8566 (I147509,I1862,I147390,I147535,);
nor I_8567 (I147358,I147535,I147424);
nand I_8568 (I147557,I147475,I147535);
nor I_8569 (I147574,I147535,I147441);
not I_8570 (I147376,I147535);
nor I_8571 (I147605,I87451,I87457);
not I_8572 (I147622,I147605);
nand I_8573 (I147379,I147574,I147605);
not I_8574 (I147653,I87442);
nor I_8575 (I147670,I147535,I87442);
nand I_8576 (I147687,I87445,I87448);
nor I_8577 (I147361,I147687,I147424);
not I_8578 (I147718,I147687);
nor I_8579 (I147735,I147605,I147718);
nor I_8580 (I147382,I147735,I147458);
nand I_8581 (I147766,I147718,I147653);
nand I_8582 (I147367,I147475,I147766);
nand I_8583 (I147797,I147557,I147766);
DFFARX1 I_8584 (I147797,I1862,I147390,I147370,);
nand I_8585 (I147828,I147622,I147687);
nor I_8586 (I147364,I147475,I147828);
nor I_8587 (I147859,I147622,I147687);
nand I_8588 (I147373,I147859,I147670);
not I_8589 (I147917,I1869);
or I_8590 (I147934,I61936,I61933);
nand I_8591 (I147951,I61939,I61936);
not I_8592 (I147968,I147951);
nand I_8593 (I147985,I147968,I147934);
not I_8594 (I148002,I147985);
nand I_8595 (I148019,I61954,I61957);
and I_8596 (I148036,I148019,I61933);
DFFARX1 I_8597 (I148036,I1862,I147917,I148062,);
nor I_8598 (I147885,I148062,I147951);
nand I_8599 (I148084,I148002,I148062);
nor I_8600 (I148101,I148062,I147968);
not I_8601 (I147903,I148062);
nor I_8602 (I148132,I61951,I61957);
not I_8603 (I148149,I148132);
nand I_8604 (I147906,I148101,I148132);
not I_8605 (I148180,I61942);
nor I_8606 (I148197,I148062,I61942);
nand I_8607 (I148214,I61945,I61948);
nor I_8608 (I147888,I148214,I147951);
not I_8609 (I148245,I148214);
nor I_8610 (I148262,I148132,I148245);
nor I_8611 (I147909,I148262,I147985);
nand I_8612 (I148293,I148245,I148180);
nand I_8613 (I147894,I148002,I148293);
nand I_8614 (I148324,I148084,I148293);
DFFARX1 I_8615 (I148324,I1862,I147917,I147897,);
nand I_8616 (I148355,I148149,I148214);
nor I_8617 (I147891,I148002,I148355);
nor I_8618 (I148386,I148149,I148214);
nand I_8619 (I147900,I148386,I148197);
not I_8620 (I148444,I1869);
or I_8621 (I148461,I54286,I54283);
nand I_8622 (I148478,I54289,I54286);
not I_8623 (I148495,I148478);
nand I_8624 (I148512,I148495,I148461);
not I_8625 (I148529,I148512);
nand I_8626 (I148546,I54304,I54307);
and I_8627 (I148563,I148546,I54283);
DFFARX1 I_8628 (I148563,I1862,I148444,I148589,);
nor I_8629 (I148412,I148589,I148478);
nand I_8630 (I148611,I148529,I148589);
nor I_8631 (I148628,I148589,I148495);
not I_8632 (I148430,I148589);
nor I_8633 (I148659,I54301,I54307);
not I_8634 (I148676,I148659);
nand I_8635 (I148433,I148628,I148659);
not I_8636 (I148707,I54292);
nor I_8637 (I148724,I148589,I54292);
nand I_8638 (I148741,I54295,I54298);
nor I_8639 (I148415,I148741,I148478);
not I_8640 (I148772,I148741);
nor I_8641 (I148789,I148659,I148772);
nor I_8642 (I148436,I148789,I148512);
nand I_8643 (I148820,I148772,I148707);
nand I_8644 (I148421,I148529,I148820);
nand I_8645 (I148851,I148611,I148820);
DFFARX1 I_8646 (I148851,I1862,I148444,I148424,);
nand I_8647 (I148882,I148676,I148741);
nor I_8648 (I148418,I148529,I148882);
nor I_8649 (I148913,I148676,I148741);
nand I_8650 (I148427,I148913,I148724);
not I_8651 (I148971,I1869);
or I_8652 (I148988,I200585,I200588);
nand I_8653 (I149005,I200591,I200600);
not I_8654 (I149022,I149005);
nand I_8655 (I149039,I149022,I148988);
not I_8656 (I149056,I149039);
nand I_8657 (I149073,I200597,I200603);
and I_8658 (I149090,I149073,I200585);
DFFARX1 I_8659 (I149090,I1862,I148971,I149116,);
nor I_8660 (I148939,I149116,I149005);
nand I_8661 (I149138,I149056,I149116);
nor I_8662 (I149155,I149116,I149022);
not I_8663 (I148957,I149116);
nor I_8664 (I149186,I200588,I200603);
not I_8665 (I149203,I149186);
nand I_8666 (I148960,I149155,I149186);
not I_8667 (I149234,I200606);
nor I_8668 (I149251,I149116,I200606);
nand I_8669 (I149268,I200594,I200591);
nor I_8670 (I148942,I149268,I149005);
not I_8671 (I149299,I149268);
nor I_8672 (I149316,I149186,I149299);
nor I_8673 (I148963,I149316,I149039);
nand I_8674 (I149347,I149299,I149234);
nand I_8675 (I148948,I149056,I149347);
nand I_8676 (I149378,I149138,I149347);
DFFARX1 I_8677 (I149378,I1862,I148971,I148951,);
nand I_8678 (I149409,I149203,I149268);
nor I_8679 (I148945,I149056,I149409);
nor I_8680 (I149440,I149203,I149268);
nand I_8681 (I148954,I149440,I149251);
not I_8682 (I149498,I1869);
or I_8683 (I149515,I387132,I387129);
nand I_8684 (I149532,I387141,I387144);
not I_8685 (I149549,I149532);
nand I_8686 (I149566,I149549,I149515);
not I_8687 (I149583,I149566);
nand I_8688 (I149600,I387135,I387126);
and I_8689 (I149617,I149600,I387126);
DFFARX1 I_8690 (I149617,I1862,I149498,I149643,);
nor I_8691 (I149466,I149643,I149532);
nand I_8692 (I149665,I149583,I149643);
nor I_8693 (I149682,I149643,I149549);
not I_8694 (I149484,I149643);
nor I_8695 (I149713,I387129,I387126);
not I_8696 (I149730,I149713);
nand I_8697 (I149487,I149682,I149713);
not I_8698 (I149761,I387132);
nor I_8699 (I149778,I149643,I387132);
nand I_8700 (I149795,I387135,I387138);
nor I_8701 (I149469,I149795,I149532);
not I_8702 (I149826,I149795);
nor I_8703 (I149843,I149713,I149826);
nor I_8704 (I149490,I149843,I149566);
nand I_8705 (I149874,I149826,I149761);
nand I_8706 (I149475,I149583,I149874);
nand I_8707 (I149905,I149665,I149874);
DFFARX1 I_8708 (I149905,I1862,I149498,I149478,);
nand I_8709 (I149936,I149730,I149795);
nor I_8710 (I149472,I149583,I149936);
nor I_8711 (I149967,I149730,I149795);
nand I_8712 (I149481,I149967,I149778);
not I_8713 (I150025,I1869);
or I_8714 (I150042,I95086,I95083);
nand I_8715 (I150059,I95089,I95086);
not I_8716 (I150076,I150059);
nand I_8717 (I150093,I150076,I150042);
not I_8718 (I150110,I150093);
nand I_8719 (I150127,I95104,I95107);
and I_8720 (I150144,I150127,I95083);
DFFARX1 I_8721 (I150144,I1862,I150025,I150170,);
nor I_8722 (I149993,I150170,I150059);
nand I_8723 (I150192,I150110,I150170);
nor I_8724 (I150209,I150170,I150076);
not I_8725 (I150011,I150170);
nor I_8726 (I150240,I95101,I95107);
not I_8727 (I150257,I150240);
nand I_8728 (I150014,I150209,I150240);
not I_8729 (I150288,I95092);
nor I_8730 (I150305,I150170,I95092);
nand I_8731 (I150322,I95095,I95098);
nor I_8732 (I149996,I150322,I150059);
not I_8733 (I150353,I150322);
nor I_8734 (I150370,I150240,I150353);
nor I_8735 (I150017,I150370,I150093);
nand I_8736 (I150401,I150353,I150288);
nand I_8737 (I150002,I150110,I150401);
nand I_8738 (I150432,I150192,I150401);
DFFARX1 I_8739 (I150432,I1862,I150025,I150005,);
nand I_8740 (I150463,I150257,I150322);
nor I_8741 (I149999,I150110,I150463);
nor I_8742 (I150494,I150257,I150322);
nand I_8743 (I150008,I150494,I150305);
not I_8744 (I150552,I1869);
or I_8745 (I150569,I382270,I382267);
nand I_8746 (I150586,I382279,I382282);
not I_8747 (I150603,I150586);
nand I_8748 (I150620,I150603,I150569);
not I_8749 (I150637,I150620);
nand I_8750 (I150654,I382273,I382264);
and I_8751 (I150671,I150654,I382264);
DFFARX1 I_8752 (I150671,I1862,I150552,I150697,);
nor I_8753 (I150520,I150697,I150586);
nand I_8754 (I150719,I150637,I150697);
nor I_8755 (I150736,I150697,I150603);
not I_8756 (I150538,I150697);
nor I_8757 (I150767,I382267,I382264);
not I_8758 (I150784,I150767);
nand I_8759 (I150541,I150736,I150767);
not I_8760 (I150815,I382270);
nor I_8761 (I150832,I150697,I382270);
nand I_8762 (I150849,I382273,I382276);
nor I_8763 (I150523,I150849,I150586);
not I_8764 (I150880,I150849);
nor I_8765 (I150897,I150767,I150880);
nor I_8766 (I150544,I150897,I150620);
nand I_8767 (I150928,I150880,I150815);
nand I_8768 (I150529,I150637,I150928);
nand I_8769 (I150959,I150719,I150928);
DFFARX1 I_8770 (I150959,I1862,I150552,I150532,);
nand I_8771 (I150990,I150784,I150849);
nor I_8772 (I150526,I150637,I150990);
nor I_8773 (I151021,I150784,I150849);
nand I_8774 (I150535,I151021,I150832);
not I_8775 (I151079,I1869);
or I_8776 (I151096,I65506,I65503);
nand I_8777 (I151113,I65509,I65506);
not I_8778 (I151130,I151113);
nand I_8779 (I151147,I151130,I151096);
not I_8780 (I151164,I151147);
nand I_8781 (I151181,I65524,I65527);
and I_8782 (I151198,I151181,I65503);
DFFARX1 I_8783 (I151198,I1862,I151079,I151224,);
nor I_8784 (I151047,I151224,I151113);
nand I_8785 (I151246,I151164,I151224);
nor I_8786 (I151263,I151224,I151130);
not I_8787 (I151065,I151224);
nor I_8788 (I151294,I65521,I65527);
not I_8789 (I151311,I151294);
nand I_8790 (I151068,I151263,I151294);
not I_8791 (I151342,I65512);
nor I_8792 (I151359,I151224,I65512);
nand I_8793 (I151376,I65515,I65518);
nor I_8794 (I151050,I151376,I151113);
not I_8795 (I151407,I151376);
nor I_8796 (I151424,I151294,I151407);
nor I_8797 (I151071,I151424,I151147);
nand I_8798 (I151455,I151407,I151342);
nand I_8799 (I151056,I151164,I151455);
nand I_8800 (I151486,I151246,I151455);
DFFARX1 I_8801 (I151486,I1862,I151079,I151059,);
nand I_8802 (I151517,I151311,I151376);
nor I_8803 (I151053,I151164,I151517);
nor I_8804 (I151548,I151311,I151376);
nand I_8805 (I151062,I151548,I151359);
not I_8806 (I151606,I1869);
or I_8807 (I151623,I20116,I20113);
nand I_8808 (I151640,I20119,I20116);
not I_8809 (I151657,I151640);
nand I_8810 (I151674,I151657,I151623);
not I_8811 (I151691,I151674);
nand I_8812 (I151708,I20134,I20137);
and I_8813 (I151725,I151708,I20113);
DFFARX1 I_8814 (I151725,I1862,I151606,I151751,);
nor I_8815 (I151574,I151751,I151640);
nand I_8816 (I151773,I151691,I151751);
nor I_8817 (I151790,I151751,I151657);
not I_8818 (I151592,I151751);
nor I_8819 (I151821,I20131,I20137);
not I_8820 (I151838,I151821);
nand I_8821 (I151595,I151790,I151821);
not I_8822 (I151869,I20122);
nor I_8823 (I151886,I151751,I20122);
nand I_8824 (I151903,I20125,I20128);
nor I_8825 (I151577,I151903,I151640);
not I_8826 (I151934,I151903);
nor I_8827 (I151951,I151821,I151934);
nor I_8828 (I151598,I151951,I151674);
nand I_8829 (I151982,I151934,I151869);
nand I_8830 (I151583,I151691,I151982);
nand I_8831 (I152013,I151773,I151982);
DFFARX1 I_8832 (I152013,I1862,I151606,I151586,);
nand I_8833 (I152044,I151838,I151903);
nor I_8834 (I151580,I151691,I152044);
nor I_8835 (I152075,I151838,I151903);
nand I_8836 (I151589,I152075,I151886);
not I_8837 (I152133,I1869);
or I_8838 (I152150,I403928,I403925);
nand I_8839 (I152167,I403937,I403940);
not I_8840 (I152184,I152167);
nand I_8841 (I152201,I152184,I152150);
not I_8842 (I152218,I152201);
nand I_8843 (I152235,I403931,I403922);
and I_8844 (I152252,I152235,I403922);
DFFARX1 I_8845 (I152252,I1862,I152133,I152278,);
nor I_8846 (I152101,I152278,I152167);
nand I_8847 (I152300,I152218,I152278);
nor I_8848 (I152317,I152278,I152184);
not I_8849 (I152119,I152278);
nor I_8850 (I152348,I403925,I403922);
not I_8851 (I152365,I152348);
nand I_8852 (I152122,I152317,I152348);
not I_8853 (I152396,I403928);
nor I_8854 (I152413,I152278,I403928);
nand I_8855 (I152430,I403931,I403934);
nor I_8856 (I152104,I152430,I152167);
not I_8857 (I152461,I152430);
nor I_8858 (I152478,I152348,I152461);
nor I_8859 (I152125,I152478,I152201);
nand I_8860 (I152509,I152461,I152396);
nand I_8861 (I152110,I152218,I152509);
nand I_8862 (I152540,I152300,I152509);
DFFARX1 I_8863 (I152540,I1862,I152133,I152113,);
nand I_8864 (I152571,I152365,I152430);
nor I_8865 (I152107,I152218,I152571);
nor I_8866 (I152602,I152365,I152430);
nand I_8867 (I152116,I152602,I152413);
not I_8868 (I152660,I1869);
or I_8869 (I152677,I306258,I306246);
nand I_8870 (I152694,I306240,I306240);
not I_8871 (I152711,I152694);
nand I_8872 (I152728,I152711,I152677);
not I_8873 (I152745,I152728);
nand I_8874 (I152762,I306243,I306243);
and I_8875 (I152779,I152762,I306249);
DFFARX1 I_8876 (I152779,I1862,I152660,I152805,);
nor I_8877 (I152628,I152805,I152694);
nand I_8878 (I152827,I152745,I152805);
nor I_8879 (I152844,I152805,I152711);
not I_8880 (I152646,I152805);
nor I_8881 (I152875,I306255,I306243);
not I_8882 (I152892,I152875);
nand I_8883 (I152649,I152844,I152875);
not I_8884 (I152923,I306261);
nor I_8885 (I152940,I152805,I306261);
nand I_8886 (I152957,I306246,I306252);
nor I_8887 (I152631,I152957,I152694);
not I_8888 (I152988,I152957);
nor I_8889 (I153005,I152875,I152988);
nor I_8890 (I152652,I153005,I152728);
nand I_8891 (I153036,I152988,I152923);
nand I_8892 (I152637,I152745,I153036);
nand I_8893 (I153067,I152827,I153036);
DFFARX1 I_8894 (I153067,I1862,I152660,I152640,);
nand I_8895 (I153098,I152892,I152957);
nor I_8896 (I152634,I152745,I153098);
nor I_8897 (I153129,I152892,I152957);
nand I_8898 (I152643,I153129,I152940);
not I_8899 (I153187,I1869);
or I_8900 (I153204,I302045,I302033);
nand I_8901 (I153221,I302036,I302030);
not I_8902 (I153238,I153221);
nand I_8903 (I153255,I153238,I153204);
not I_8904 (I153272,I153255);
nand I_8905 (I153289,I302027,I302030);
and I_8906 (I153306,I153289,I302024);
DFFARX1 I_8907 (I153306,I1862,I153187,I153332,);
nor I_8908 (I153155,I153332,I153221);
nand I_8909 (I153354,I153272,I153332);
nor I_8910 (I153371,I153332,I153238);
not I_8911 (I153173,I153332);
nor I_8912 (I153402,I302024,I302030);
not I_8913 (I153419,I153402);
nand I_8914 (I153176,I153371,I153402);
not I_8915 (I153450,I302027);
nor I_8916 (I153467,I153332,I302027);
nand I_8917 (I153484,I302042,I302039);
nor I_8918 (I153158,I153484,I153221);
not I_8919 (I153515,I153484);
nor I_8920 (I153532,I153402,I153515);
nor I_8921 (I153179,I153532,I153255);
nand I_8922 (I153563,I153515,I153450);
nand I_8923 (I153164,I153272,I153563);
nand I_8924 (I153594,I153354,I153563);
DFFARX1 I_8925 (I153594,I1862,I153187,I153167,);
nand I_8926 (I153625,I153419,I153484);
nor I_8927 (I153161,I153272,I153625);
nor I_8928 (I153656,I153419,I153484);
nand I_8929 (I153170,I153656,I153467);
not I_8930 (I153714,I1869);
or I_8931 (I153731,I104677,I104686);
nand I_8932 (I153748,I104680,I104683);
not I_8933 (I153765,I153748);
nand I_8934 (I153782,I153765,I153731);
not I_8935 (I153799,I153782);
nand I_8936 (I153816,I104674,I104674);
and I_8937 (I153833,I153816,I104671);
DFFARX1 I_8938 (I153833,I1862,I153714,I153859,);
nor I_8939 (I153682,I153859,I153748);
nand I_8940 (I153881,I153799,I153859);
nor I_8941 (I153898,I153859,I153765);
not I_8942 (I153700,I153859);
nor I_8943 (I153929,I104689,I104674);
not I_8944 (I153946,I153929);
nand I_8945 (I153703,I153898,I153929);
not I_8946 (I153977,I104677);
nor I_8947 (I153994,I153859,I104677);
nand I_8948 (I154011,I104680,I104671);
nor I_8949 (I153685,I154011,I153748);
not I_8950 (I154042,I154011);
nor I_8951 (I154059,I153929,I154042);
nor I_8952 (I153706,I154059,I153782);
nand I_8953 (I154090,I154042,I153977);
nand I_8954 (I153691,I153799,I154090);
nand I_8955 (I154121,I153881,I154090);
DFFARX1 I_8956 (I154121,I1862,I153714,I153694,);
nand I_8957 (I154152,I153946,I154011);
nor I_8958 (I153688,I153799,I154152);
nor I_8959 (I154183,I153946,I154011);
nand I_8960 (I153697,I154183,I153994);
not I_8961 (I154241,I1869);
or I_8962 (I154258,I76726,I76723);
nand I_8963 (I154275,I76729,I76726);
not I_8964 (I154292,I154275);
nand I_8965 (I154309,I154292,I154258);
not I_8966 (I154326,I154309);
nand I_8967 (I154343,I76744,I76747);
and I_8968 (I154360,I154343,I76723);
DFFARX1 I_8969 (I154360,I1862,I154241,I154386,);
nor I_8970 (I154209,I154386,I154275);
nand I_8971 (I154408,I154326,I154386);
nor I_8972 (I154425,I154386,I154292);
not I_8973 (I154227,I154386);
nor I_8974 (I154456,I76741,I76747);
not I_8975 (I154473,I154456);
nand I_8976 (I154230,I154425,I154456);
not I_8977 (I154504,I76732);
nor I_8978 (I154521,I154386,I76732);
nand I_8979 (I154538,I76735,I76738);
nor I_8980 (I154212,I154538,I154275);
not I_8981 (I154569,I154538);
nor I_8982 (I154586,I154456,I154569);
nor I_8983 (I154233,I154586,I154309);
nand I_8984 (I154617,I154569,I154504);
nand I_8985 (I154218,I154326,I154617);
nand I_8986 (I154648,I154408,I154617);
DFFARX1 I_8987 (I154648,I1862,I154241,I154221,);
nand I_8988 (I154679,I154473,I154538);
nor I_8989 (I154215,I154326,I154679);
nor I_8990 (I154710,I154473,I154538);
nand I_8991 (I154224,I154710,I154521);
not I_8992 (I154768,I1869);
or I_8993 (I154785,I15016,I15013);
nand I_8994 (I154802,I15019,I15016);
not I_8995 (I154819,I154802);
nand I_8996 (I154836,I154819,I154785);
not I_8997 (I154853,I154836);
nand I_8998 (I154870,I15034,I15037);
and I_8999 (I154887,I154870,I15013);
DFFARX1 I_9000 (I154887,I1862,I154768,I154913,);
nor I_9001 (I154736,I154913,I154802);
nand I_9002 (I154935,I154853,I154913);
nor I_9003 (I154952,I154913,I154819);
not I_9004 (I154754,I154913);
nor I_9005 (I154983,I15031,I15037);
not I_9006 (I155000,I154983);
nand I_9007 (I154757,I154952,I154983);
not I_9008 (I155031,I15022);
nor I_9009 (I155048,I154913,I15022);
nand I_9010 (I155065,I15025,I15028);
nor I_9011 (I154739,I155065,I154802);
not I_9012 (I155096,I155065);
nor I_9013 (I155113,I154983,I155096);
nor I_9014 (I154760,I155113,I154836);
nand I_9015 (I155144,I155096,I155031);
nand I_9016 (I154745,I154853,I155144);
nand I_9017 (I155175,I154935,I155144);
DFFARX1 I_9018 (I155175,I1862,I154768,I154748,);
nand I_9019 (I155206,I155000,I155065);
nor I_9020 (I154742,I154853,I155206);
nor I_9021 (I155237,I155000,I155065);
nand I_9022 (I154751,I155237,I155048);
not I_9023 (I155295,I1869);
or I_9024 (I155312,I27766,I27763);
nand I_9025 (I155329,I27769,I27766);
not I_9026 (I155346,I155329);
nand I_9027 (I155363,I155346,I155312);
not I_9028 (I155380,I155363);
nand I_9029 (I155397,I27784,I27787);
and I_9030 (I155414,I155397,I27763);
DFFARX1 I_9031 (I155414,I1862,I155295,I155440,);
nor I_9032 (I155263,I155440,I155329);
nand I_9033 (I155462,I155380,I155440);
nor I_9034 (I155479,I155440,I155346);
not I_9035 (I155281,I155440);
nor I_9036 (I155510,I27781,I27787);
not I_9037 (I155527,I155510);
nand I_9038 (I155284,I155479,I155510);
not I_9039 (I155558,I27772);
nor I_9040 (I155575,I155440,I27772);
nand I_9041 (I155592,I27775,I27778);
nor I_9042 (I155266,I155592,I155329);
not I_9043 (I155623,I155592);
nor I_9044 (I155640,I155510,I155623);
nor I_9045 (I155287,I155640,I155363);
nand I_9046 (I155671,I155623,I155558);
nand I_9047 (I155272,I155380,I155671);
nand I_9048 (I155702,I155462,I155671);
DFFARX1 I_9049 (I155702,I1862,I155295,I155275,);
nand I_9050 (I155733,I155527,I155592);
nor I_9051 (I155269,I155380,I155733);
nor I_9052 (I155764,I155527,I155592);
nand I_9053 (I155278,I155764,I155575);
not I_9054 (I155822,I1869);
or I_9055 (I155839,I278173,I278176);
nand I_9056 (I155856,I278179,I278188);
not I_9057 (I155873,I155856);
nand I_9058 (I155890,I155873,I155839);
not I_9059 (I155907,I155890);
nand I_9060 (I155924,I278185,I278191);
and I_9061 (I155941,I155924,I278173);
DFFARX1 I_9062 (I155941,I1862,I155822,I155967,);
nor I_9063 (I155790,I155967,I155856);
nand I_9064 (I155989,I155907,I155967);
nor I_9065 (I156006,I155967,I155873);
not I_9066 (I155808,I155967);
nor I_9067 (I156037,I278176,I278191);
not I_9068 (I156054,I156037);
nand I_9069 (I155811,I156006,I156037);
not I_9070 (I156085,I278194);
nor I_9071 (I156102,I155967,I278194);
nand I_9072 (I156119,I278182,I278179);
nor I_9073 (I155793,I156119,I155856);
not I_9074 (I156150,I156119);
nor I_9075 (I156167,I156037,I156150);
nor I_9076 (I155814,I156167,I155890);
nand I_9077 (I156198,I156150,I156085);
nand I_9078 (I155799,I155907,I156198);
nand I_9079 (I156229,I155989,I156198);
DFFARX1 I_9080 (I156229,I1862,I155822,I155802,);
nand I_9081 (I156260,I156054,I156119);
nor I_9082 (I155796,I155907,I156260);
nor I_9083 (I156291,I156054,I156119);
nand I_9084 (I155805,I156291,I156102);
not I_9085 (I156349,I1869);
or I_9086 (I156366,I367684,I367681);
nand I_9087 (I156383,I367693,I367696);
not I_9088 (I156400,I156383);
nand I_9089 (I156417,I156400,I156366);
not I_9090 (I156434,I156417);
nand I_9091 (I156451,I367687,I367678);
and I_9092 (I156468,I156451,I367678);
DFFARX1 I_9093 (I156468,I1862,I156349,I156494,);
nor I_9094 (I156317,I156494,I156383);
nand I_9095 (I156516,I156434,I156494);
nor I_9096 (I156533,I156494,I156400);
not I_9097 (I156335,I156494);
nor I_9098 (I156564,I367681,I367678);
not I_9099 (I156581,I156564);
nand I_9100 (I156338,I156533,I156564);
not I_9101 (I156612,I367684);
nor I_9102 (I156629,I156494,I367684);
nand I_9103 (I156646,I367687,I367690);
nor I_9104 (I156320,I156646,I156383);
not I_9105 (I156677,I156646);
nor I_9106 (I156694,I156564,I156677);
nor I_9107 (I156341,I156694,I156417);
nand I_9108 (I156725,I156677,I156612);
nand I_9109 (I156326,I156434,I156725);
nand I_9110 (I156756,I156516,I156725);
DFFARX1 I_9111 (I156756,I1862,I156349,I156329,);
nand I_9112 (I156787,I156581,I156646);
nor I_9113 (I156323,I156434,I156787);
nor I_9114 (I156818,I156581,I156646);
nand I_9115 (I156332,I156818,I156629);
not I_9116 (I156876,I1869);
or I_9117 (I156893,I254849,I254852);
nand I_9118 (I156910,I254855,I254864);
not I_9119 (I156927,I156910);
nand I_9120 (I156944,I156927,I156893);
not I_9121 (I156961,I156944);
nand I_9122 (I156978,I254861,I254867);
and I_9123 (I156995,I156978,I254849);
DFFARX1 I_9124 (I156995,I1862,I156876,I157021,);
nor I_9125 (I156844,I157021,I156910);
nand I_9126 (I157043,I156961,I157021);
nor I_9127 (I157060,I157021,I156927);
not I_9128 (I156862,I157021);
nor I_9129 (I157091,I254852,I254867);
not I_9130 (I157108,I157091);
nand I_9131 (I156865,I157060,I157091);
not I_9132 (I157139,I254870);
nor I_9133 (I157156,I157021,I254870);
nand I_9134 (I157173,I254858,I254855);
nor I_9135 (I156847,I157173,I156910);
not I_9136 (I157204,I157173);
nor I_9137 (I157221,I157091,I157204);
nor I_9138 (I156868,I157221,I156944);
nand I_9139 (I157252,I157204,I157139);
nand I_9140 (I156853,I156961,I157252);
nand I_9141 (I157283,I157043,I157252);
DFFARX1 I_9142 (I157283,I1862,I156876,I156856,);
nand I_9143 (I157314,I157108,I157173);
nor I_9144 (I156850,I156961,I157314);
nor I_9145 (I157345,I157108,I157173);
nand I_9146 (I156859,I157345,I157156);
not I_9147 (I157403,I1869);
or I_9148 (I157420,I225813,I225816);
nand I_9149 (I157437,I225819,I225828);
not I_9150 (I157454,I157437);
nand I_9151 (I157471,I157454,I157420);
not I_9152 (I157488,I157471);
nand I_9153 (I157505,I225825,I225831);
and I_9154 (I157522,I157505,I225813);
DFFARX1 I_9155 (I157522,I1862,I157403,I157548,);
nor I_9156 (I157371,I157548,I157437);
nand I_9157 (I157570,I157488,I157548);
nor I_9158 (I157587,I157548,I157454);
not I_9159 (I157389,I157548);
nor I_9160 (I157618,I225816,I225831);
not I_9161 (I157635,I157618);
nand I_9162 (I157392,I157587,I157618);
not I_9163 (I157666,I225834);
nor I_9164 (I157683,I157548,I225834);
nand I_9165 (I157700,I225822,I225819);
nor I_9166 (I157374,I157700,I157437);
not I_9167 (I157731,I157700);
nor I_9168 (I157748,I157618,I157731);
nor I_9169 (I157395,I157748,I157471);
nand I_9170 (I157779,I157731,I157666);
nand I_9171 (I157380,I157488,I157779);
nand I_9172 (I157810,I157570,I157779);
DFFARX1 I_9173 (I157810,I1862,I157403,I157383,);
nand I_9174 (I157841,I157635,I157700);
nor I_9175 (I157377,I157488,I157841);
nor I_9176 (I157872,I157635,I157700);
nand I_9177 (I157386,I157872,I157683);
not I_9178 (I157930,I1869);
or I_9179 (I157947,I376082,I376079);
nand I_9180 (I157964,I376091,I376094);
not I_9181 (I157981,I157964);
nand I_9182 (I157998,I157981,I157947);
not I_9183 (I158015,I157998);
nand I_9184 (I158032,I376085,I376076);
and I_9185 (I158049,I158032,I376076);
DFFARX1 I_9186 (I158049,I1862,I157930,I158075,);
nor I_9187 (I157898,I158075,I157964);
nand I_9188 (I158097,I158015,I158075);
nor I_9189 (I158114,I158075,I157981);
not I_9190 (I157916,I158075);
nor I_9191 (I158145,I376079,I376076);
not I_9192 (I158162,I158145);
nand I_9193 (I157919,I158114,I158145);
not I_9194 (I158193,I376082);
nor I_9195 (I158210,I158075,I376082);
nand I_9196 (I158227,I376085,I376088);
nor I_9197 (I157901,I158227,I157964);
not I_9198 (I158258,I158227);
nor I_9199 (I158275,I158145,I158258);
nor I_9200 (I157922,I158275,I157998);
nand I_9201 (I158306,I158258,I158193);
nand I_9202 (I157907,I158015,I158306);
nand I_9203 (I158337,I158097,I158306);
DFFARX1 I_9204 (I158337,I1862,I157930,I157910,);
nand I_9205 (I158368,I158162,I158227);
nor I_9206 (I157904,I158015,I158368);
nor I_9207 (I158399,I158162,I158227);
nand I_9208 (I157913,I158399,I158210);
not I_9209 (I158457,I1869);
or I_9210 (I158474,I99166,I99163);
nand I_9211 (I158491,I99169,I99166);
not I_9212 (I158508,I158491);
nand I_9213 (I158525,I158508,I158474);
not I_9214 (I158542,I158525);
nand I_9215 (I158559,I99184,I99187);
and I_9216 (I158576,I158559,I99163);
DFFARX1 I_9217 (I158576,I1862,I158457,I158602,);
nor I_9218 (I158425,I158602,I158491);
nand I_9219 (I158624,I158542,I158602);
nor I_9220 (I158641,I158602,I158508);
not I_9221 (I158443,I158602);
nor I_9222 (I158672,I99181,I99187);
not I_9223 (I158689,I158672);
nand I_9224 (I158446,I158641,I158672);
not I_9225 (I158720,I99172);
nor I_9226 (I158737,I158602,I99172);
nand I_9227 (I158754,I99175,I99178);
nor I_9228 (I158428,I158754,I158491);
not I_9229 (I158785,I158754);
nor I_9230 (I158802,I158672,I158785);
nor I_9231 (I158449,I158802,I158525);
nand I_9232 (I158833,I158785,I158720);
nand I_9233 (I158434,I158542,I158833);
nand I_9234 (I158864,I158624,I158833);
DFFARX1 I_9235 (I158864,I1862,I158457,I158437,);
nand I_9236 (I158895,I158689,I158754);
nor I_9237 (I158431,I158542,I158895);
nor I_9238 (I158926,I158689,I158754);
nand I_9239 (I158440,I158926,I158737);
not I_9240 (I158984,I1869);
or I_9241 (I159001,I366358,I366355);
nand I_9242 (I159018,I366367,I366370);
not I_9243 (I159035,I159018);
nand I_9244 (I159052,I159035,I159001);
not I_9245 (I159069,I159052);
nand I_9246 (I159086,I366361,I366352);
and I_9247 (I159103,I159086,I366352);
DFFARX1 I_9248 (I159103,I1862,I158984,I159129,);
nor I_9249 (I158952,I159129,I159018);
nand I_9250 (I159151,I159069,I159129);
nor I_9251 (I159168,I159129,I159035);
not I_9252 (I158970,I159129);
nor I_9253 (I159199,I366355,I366352);
not I_9254 (I159216,I159199);
nand I_9255 (I158973,I159168,I159199);
not I_9256 (I159247,I366358);
nor I_9257 (I159264,I159129,I366358);
nand I_9258 (I159281,I366361,I366364);
nor I_9259 (I158955,I159281,I159018);
not I_9260 (I159312,I159281);
nor I_9261 (I159329,I159199,I159312);
nor I_9262 (I158976,I159329,I159052);
nand I_9263 (I159360,I159312,I159247);
nand I_9264 (I158961,I159069,I159360);
nand I_9265 (I159391,I159151,I159360);
DFFARX1 I_9266 (I159391,I1862,I158984,I158964,);
nand I_9267 (I159422,I159216,I159281);
nor I_9268 (I158958,I159069,I159422);
nor I_9269 (I159453,I159216,I159281);
nand I_9270 (I158967,I159453,I159264);
not I_9271 (I159511,I1869);
or I_9272 (I159528,I303623,I303611);
nand I_9273 (I159545,I303605,I303605);
not I_9274 (I159562,I159545);
nand I_9275 (I159579,I159562,I159528);
not I_9276 (I159596,I159579);
nand I_9277 (I159613,I303608,I303608);
and I_9278 (I159630,I159613,I303614);
DFFARX1 I_9279 (I159630,I1862,I159511,I159656,);
nor I_9280 (I159479,I159656,I159545);
nand I_9281 (I159678,I159596,I159656);
nor I_9282 (I159695,I159656,I159562);
not I_9283 (I159497,I159656);
nor I_9284 (I159726,I303620,I303608);
not I_9285 (I159743,I159726);
nand I_9286 (I159500,I159695,I159726);
not I_9287 (I159774,I303626);
nor I_9288 (I159791,I159656,I303626);
nand I_9289 (I159808,I303611,I303617);
nor I_9290 (I159482,I159808,I159545);
not I_9291 (I159839,I159808);
nor I_9292 (I159856,I159726,I159839);
nor I_9293 (I159503,I159856,I159579);
nand I_9294 (I159887,I159839,I159774);
nand I_9295 (I159488,I159596,I159887);
nand I_9296 (I159918,I159678,I159887);
DFFARX1 I_9297 (I159918,I1862,I159511,I159491,);
nand I_9298 (I159949,I159743,I159808);
nor I_9299 (I159485,I159596,I159949);
nor I_9300 (I159980,I159743,I159808);
nand I_9301 (I159494,I159980,I159791);
not I_9302 (I160038,I1869);
or I_9303 (I160055,I241997,I242000);
nand I_9304 (I160072,I242003,I242012);
not I_9305 (I160089,I160072);
nand I_9306 (I160106,I160089,I160055);
not I_9307 (I160123,I160106);
nand I_9308 (I160140,I242009,I242015);
and I_9309 (I160157,I160140,I241997);
DFFARX1 I_9310 (I160157,I1862,I160038,I160183,);
nor I_9311 (I160006,I160183,I160072);
nand I_9312 (I160205,I160123,I160183);
nor I_9313 (I160222,I160183,I160089);
not I_9314 (I160024,I160183);
nor I_9315 (I160253,I242000,I242015);
not I_9316 (I160270,I160253);
nand I_9317 (I160027,I160222,I160253);
not I_9318 (I160301,I242018);
nor I_9319 (I160318,I160183,I242018);
nand I_9320 (I160335,I242006,I242003);
nor I_9321 (I160009,I160335,I160072);
not I_9322 (I160366,I160335);
nor I_9323 (I160383,I160253,I160366);
nor I_9324 (I160030,I160383,I160106);
nand I_9325 (I160414,I160366,I160301);
nand I_9326 (I160015,I160123,I160414);
nand I_9327 (I160445,I160205,I160414);
DFFARX1 I_9328 (I160445,I1862,I160038,I160018,);
nand I_9329 (I160476,I160270,I160335);
nor I_9330 (I160012,I160123,I160476);
nor I_9331 (I160507,I160270,I160335);
nand I_9332 (I160021,I160507,I160318);
not I_9333 (I160565,I1869);
or I_9334 (I160582,I112837,I112846);
nand I_9335 (I160599,I112840,I112843);
not I_9336 (I160616,I160599);
nand I_9337 (I160633,I160616,I160582);
not I_9338 (I160650,I160633);
nand I_9339 (I160667,I112834,I112834);
and I_9340 (I160684,I160667,I112831);
DFFARX1 I_9341 (I160684,I1862,I160565,I160710,);
nor I_9342 (I160533,I160710,I160599);
nand I_9343 (I160732,I160650,I160710);
nor I_9344 (I160749,I160710,I160616);
not I_9345 (I160551,I160710);
nor I_9346 (I160780,I112849,I112834);
not I_9347 (I160797,I160780);
nand I_9348 (I160554,I160749,I160780);
not I_9349 (I160828,I112837);
nor I_9350 (I160845,I160710,I112837);
nand I_9351 (I160862,I112840,I112831);
nor I_9352 (I160536,I160862,I160599);
not I_9353 (I160893,I160862);
nor I_9354 (I160910,I160780,I160893);
nor I_9355 (I160557,I160910,I160633);
nand I_9356 (I160941,I160893,I160828);
nand I_9357 (I160542,I160650,I160941);
nand I_9358 (I160972,I160732,I160941);
DFFARX1 I_9359 (I160972,I1862,I160565,I160545,);
nand I_9360 (I161003,I160797,I160862);
nor I_9361 (I160539,I160650,I161003);
nor I_9362 (I161034,I160797,I160862);
nand I_9363 (I160548,I161034,I160845);
not I_9364 (I161092,I1869);
or I_9365 (I161109,I361054,I361051);
nand I_9366 (I161126,I361063,I361066);
not I_9367 (I161143,I161126);
nand I_9368 (I161160,I161143,I161109);
not I_9369 (I161177,I161160);
nand I_9370 (I161194,I361057,I361048);
and I_9371 (I161211,I161194,I361048);
DFFARX1 I_9372 (I161211,I1862,I161092,I161237,);
nor I_9373 (I161060,I161237,I161126);
nand I_9374 (I161259,I161177,I161237);
nor I_9375 (I161276,I161237,I161143);
not I_9376 (I161078,I161237);
nor I_9377 (I161307,I361051,I361048);
not I_9378 (I161324,I161307);
nand I_9379 (I161081,I161276,I161307);
not I_9380 (I161355,I361054);
nor I_9381 (I161372,I161237,I361054);
nand I_9382 (I161389,I361057,I361060);
nor I_9383 (I161063,I161389,I161126);
not I_9384 (I161420,I161389);
nor I_9385 (I161437,I161307,I161420);
nor I_9386 (I161084,I161437,I161160);
nand I_9387 (I161468,I161420,I161355);
nand I_9388 (I161069,I161177,I161468);
nand I_9389 (I161499,I161259,I161468);
DFFARX1 I_9390 (I161499,I1862,I161092,I161072,);
nand I_9391 (I161530,I161324,I161389);
nor I_9392 (I161066,I161177,I161530);
nor I_9393 (I161561,I161324,I161389);
nand I_9394 (I161075,I161561,I161372);
not I_9395 (I161619,I1869);
or I_9396 (I161636,I40006,I40003);
nand I_9397 (I161653,I40009,I40006);
not I_9398 (I161670,I161653);
nand I_9399 (I161687,I161670,I161636);
not I_9400 (I161704,I161687);
nand I_9401 (I161721,I40024,I40027);
and I_9402 (I161738,I161721,I40003);
DFFARX1 I_9403 (I161738,I1862,I161619,I161764,);
nor I_9404 (I161587,I161764,I161653);
nand I_9405 (I161786,I161704,I161764);
nor I_9406 (I161803,I161764,I161670);
not I_9407 (I161605,I161764);
nor I_9408 (I161834,I40021,I40027);
not I_9409 (I161851,I161834);
nand I_9410 (I161608,I161803,I161834);
not I_9411 (I161882,I40012);
nor I_9412 (I161899,I161764,I40012);
nand I_9413 (I161916,I40015,I40018);
nor I_9414 (I161590,I161916,I161653);
not I_9415 (I161947,I161916);
nor I_9416 (I161964,I161834,I161947);
nor I_9417 (I161611,I161964,I161687);
nand I_9418 (I161995,I161947,I161882);
nand I_9419 (I161596,I161704,I161995);
nand I_9420 (I162026,I161786,I161995);
DFFARX1 I_9421 (I162026,I1862,I161619,I161599,);
nand I_9422 (I162057,I161851,I161916);
nor I_9423 (I161593,I161704,I162057);
nor I_9424 (I162088,I161851,I161916);
nand I_9425 (I161602,I162088,I161899);
not I_9426 (I162146,I1869);
or I_9427 (I162163,I248661,I248664);
nand I_9428 (I162180,I248667,I248676);
not I_9429 (I162197,I162180);
nand I_9430 (I162214,I162197,I162163);
not I_9431 (I162231,I162214);
nand I_9432 (I162248,I248673,I248679);
and I_9433 (I162265,I162248,I248661);
DFFARX1 I_9434 (I162265,I1862,I162146,I162291,);
nor I_9435 (I162114,I162291,I162180);
nand I_9436 (I162313,I162231,I162291);
nor I_9437 (I162330,I162291,I162197);
not I_9438 (I162132,I162291);
nor I_9439 (I162361,I248664,I248679);
not I_9440 (I162378,I162361);
nand I_9441 (I162135,I162330,I162361);
not I_9442 (I162409,I248682);
nor I_9443 (I162426,I162291,I248682);
nand I_9444 (I162443,I248670,I248667);
nor I_9445 (I162117,I162443,I162180);
not I_9446 (I162474,I162443);
nor I_9447 (I162491,I162361,I162474);
nor I_9448 (I162138,I162491,I162214);
nand I_9449 (I162522,I162474,I162409);
nand I_9450 (I162123,I162231,I162522);
nand I_9451 (I162553,I162313,I162522);
DFFARX1 I_9452 (I162553,I1862,I162146,I162126,);
nand I_9453 (I162584,I162378,I162443);
nor I_9454 (I162120,I162231,I162584);
nor I_9455 (I162615,I162378,I162443);
nand I_9456 (I162129,I162615,I162426);
not I_9457 (I162673,I1869);
or I_9458 (I162690,I371220,I371217);
nand I_9459 (I162707,I371229,I371232);
not I_9460 (I162724,I162707);
nand I_9461 (I162741,I162724,I162690);
not I_9462 (I162758,I162741);
nand I_9463 (I162775,I371223,I371214);
and I_9464 (I162792,I162775,I371214);
DFFARX1 I_9465 (I162792,I1862,I162673,I162818,);
nor I_9466 (I162641,I162818,I162707);
nand I_9467 (I162840,I162758,I162818);
nor I_9468 (I162857,I162818,I162724);
not I_9469 (I162659,I162818);
nor I_9470 (I162888,I371217,I371214);
not I_9471 (I162905,I162888);
nand I_9472 (I162662,I162857,I162888);
not I_9473 (I162936,I371220);
nor I_9474 (I162953,I162818,I371220);
nand I_9475 (I162970,I371223,I371226);
nor I_9476 (I162644,I162970,I162707);
not I_9477 (I163001,I162970);
nor I_9478 (I163018,I162888,I163001);
nor I_9479 (I162665,I163018,I162741);
nand I_9480 (I163049,I163001,I162936);
nand I_9481 (I162650,I162758,I163049);
nand I_9482 (I163080,I162840,I163049);
DFFARX1 I_9483 (I163080,I1862,I162673,I162653,);
nand I_9484 (I163111,I162905,I162970);
nor I_9485 (I162647,I162758,I163111);
nor I_9486 (I163142,I162905,I162970);
nand I_9487 (I162656,I163142,I162953);
not I_9488 (I163200,I1869);
or I_9489 (I163217,I369010,I369007);
nand I_9490 (I163234,I369019,I369022);
not I_9491 (I163251,I163234);
nand I_9492 (I163268,I163251,I163217);
not I_9493 (I163285,I163268);
nand I_9494 (I163302,I369013,I369004);
and I_9495 (I163319,I163302,I369004);
DFFARX1 I_9496 (I163319,I1862,I163200,I163345,);
nor I_9497 (I163168,I163345,I163234);
nand I_9498 (I163367,I163285,I163345);
nor I_9499 (I163384,I163345,I163251);
not I_9500 (I163186,I163345);
nor I_9501 (I163415,I369007,I369004);
not I_9502 (I163432,I163415);
nand I_9503 (I163189,I163384,I163415);
not I_9504 (I163463,I369010);
nor I_9505 (I163480,I163345,I369010);
nand I_9506 (I163497,I369013,I369016);
nor I_9507 (I163171,I163497,I163234);
not I_9508 (I163528,I163497);
nor I_9509 (I163545,I163415,I163528);
nor I_9510 (I163192,I163545,I163268);
nand I_9511 (I163576,I163528,I163463);
nand I_9512 (I163177,I163285,I163576);
nand I_9513 (I163607,I163367,I163576);
DFFARX1 I_9514 (I163607,I1862,I163200,I163180,);
nand I_9515 (I163638,I163432,I163497);
nor I_9516 (I163174,I163285,I163638);
nor I_9517 (I163669,I163432,I163497);
nand I_9518 (I163183,I163669,I163480);
not I_9519 (I163727,I1869);
or I_9520 (I163744,I271985,I271988);
nand I_9521 (I163761,I271991,I272000);
not I_9522 (I163778,I163761);
nand I_9523 (I163795,I163778,I163744);
not I_9524 (I163812,I163795);
nand I_9525 (I163829,I271997,I272003);
and I_9526 (I163846,I163829,I271985);
DFFARX1 I_9527 (I163846,I1862,I163727,I163872,);
nor I_9528 (I163695,I163872,I163761);
nand I_9529 (I163894,I163812,I163872);
nor I_9530 (I163911,I163872,I163778);
not I_9531 (I163713,I163872);
nor I_9532 (I163942,I271988,I272003);
not I_9533 (I163959,I163942);
nand I_9534 (I163716,I163911,I163942);
not I_9535 (I163990,I272006);
nor I_9536 (I164007,I163872,I272006);
nand I_9537 (I164024,I271994,I271991);
nor I_9538 (I163698,I164024,I163761);
not I_9539 (I164055,I164024);
nor I_9540 (I164072,I163942,I164055);
nor I_9541 (I163719,I164072,I163795);
nand I_9542 (I164103,I164055,I163990);
nand I_9543 (I163704,I163812,I164103);
nand I_9544 (I164134,I163894,I164103);
DFFARX1 I_9545 (I164134,I1862,I163727,I163707,);
nand I_9546 (I164165,I163959,I164024);
nor I_9547 (I163701,I163812,I164165);
nor I_9548 (I164196,I163959,I164024);
nand I_9549 (I163710,I164196,I164007);
not I_9550 (I164254,I1869);
or I_9551 (I164271,I209629,I209632);
nand I_9552 (I164288,I209635,I209644);
not I_9553 (I164305,I164288);
nand I_9554 (I164322,I164305,I164271);
not I_9555 (I164339,I164322);
nand I_9556 (I164356,I209641,I209647);
and I_9557 (I164373,I164356,I209629);
DFFARX1 I_9558 (I164373,I1862,I164254,I164399,);
nor I_9559 (I164222,I164399,I164288);
nand I_9560 (I164421,I164339,I164399);
nor I_9561 (I164438,I164399,I164305);
not I_9562 (I164240,I164399);
nor I_9563 (I164469,I209632,I209647);
not I_9564 (I164486,I164469);
nand I_9565 (I164243,I164438,I164469);
not I_9566 (I164517,I209650);
nor I_9567 (I164534,I164399,I209650);
nand I_9568 (I164551,I209638,I209635);
nor I_9569 (I164225,I164551,I164288);
not I_9570 (I164582,I164551);
nor I_9571 (I164599,I164469,I164582);
nor I_9572 (I164246,I164599,I164322);
nand I_9573 (I164630,I164582,I164517);
nand I_9574 (I164231,I164339,I164630);
nand I_9575 (I164661,I164421,I164630);
DFFARX1 I_9576 (I164661,I1862,I164254,I164234,);
nand I_9577 (I164692,I164486,I164551);
nor I_9578 (I164228,I164339,I164692);
nor I_9579 (I164723,I164486,I164551);
nand I_9580 (I164237,I164723,I164534);
not I_9581 (I164781,I1869);
or I_9582 (I164798,I42046,I42043);
nand I_9583 (I164815,I42049,I42046);
not I_9584 (I164832,I164815);
nand I_9585 (I164849,I164832,I164798);
not I_9586 (I164866,I164849);
nand I_9587 (I164883,I42064,I42067);
and I_9588 (I164900,I164883,I42043);
DFFARX1 I_9589 (I164900,I1862,I164781,I164926,);
nor I_9590 (I164749,I164926,I164815);
nand I_9591 (I164948,I164866,I164926);
nor I_9592 (I164965,I164926,I164832);
not I_9593 (I164767,I164926);
nor I_9594 (I164996,I42061,I42067);
not I_9595 (I165013,I164996);
nand I_9596 (I164770,I164965,I164996);
not I_9597 (I165044,I42052);
nor I_9598 (I165061,I164926,I42052);
nand I_9599 (I165078,I42055,I42058);
nor I_9600 (I164752,I165078,I164815);
not I_9601 (I165109,I165078);
nor I_9602 (I165126,I164996,I165109);
nor I_9603 (I164773,I165126,I164849);
nand I_9604 (I165157,I165109,I165044);
nand I_9605 (I164758,I164866,I165157);
nand I_9606 (I165188,I164948,I165157);
DFFARX1 I_9607 (I165188,I1862,I164781,I164761,);
nand I_9608 (I165219,I165013,I165078);
nor I_9609 (I164755,I164866,I165219);
nor I_9610 (I165250,I165013,I165078);
nand I_9611 (I164764,I165250,I165061);
not I_9612 (I165308,I1869);
or I_9613 (I165325,I106309,I106318);
nand I_9614 (I165342,I106312,I106315);
not I_9615 (I165359,I165342);
nand I_9616 (I165376,I165359,I165325);
not I_9617 (I165393,I165376);
nand I_9618 (I165410,I106306,I106306);
and I_9619 (I165427,I165410,I106303);
DFFARX1 I_9620 (I165427,I1862,I165308,I165453,);
nor I_9621 (I165276,I165453,I165342);
nand I_9622 (I165475,I165393,I165453);
nor I_9623 (I165492,I165453,I165359);
not I_9624 (I165294,I165453);
nor I_9625 (I165523,I106321,I106306);
not I_9626 (I165540,I165523);
nand I_9627 (I165297,I165492,I165523);
not I_9628 (I165571,I106309);
nor I_9629 (I165588,I165453,I106309);
nand I_9630 (I165605,I106312,I106303);
nor I_9631 (I165279,I165605,I165342);
not I_9632 (I165636,I165605);
nor I_9633 (I165653,I165523,I165636);
nor I_9634 (I165300,I165653,I165376);
nand I_9635 (I165684,I165636,I165571);
nand I_9636 (I165285,I165393,I165684);
nand I_9637 (I165715,I165475,I165684);
DFFARX1 I_9638 (I165715,I1862,I165308,I165288,);
nand I_9639 (I165746,I165540,I165605);
nor I_9640 (I165282,I165393,I165746);
nor I_9641 (I165777,I165540,I165605);
nand I_9642 (I165291,I165777,I165588);
not I_9643 (I165835,I1869);
or I_9644 (I165852,I277697,I277700);
nand I_9645 (I165869,I277703,I277712);
not I_9646 (I165886,I165869);
nand I_9647 (I165903,I165886,I165852);
not I_9648 (I165920,I165903);
nand I_9649 (I165937,I277709,I277715);
and I_9650 (I165954,I165937,I277697);
DFFARX1 I_9651 (I165954,I1862,I165835,I165980,);
nor I_9652 (I165803,I165980,I165869);
nand I_9653 (I166002,I165920,I165980);
nor I_9654 (I166019,I165980,I165886);
not I_9655 (I165821,I165980);
nor I_9656 (I166050,I277700,I277715);
not I_9657 (I166067,I166050);
nand I_9658 (I165824,I166019,I166050);
not I_9659 (I166098,I277718);
nor I_9660 (I166115,I165980,I277718);
nand I_9661 (I166132,I277706,I277703);
nor I_9662 (I165806,I166132,I165869);
not I_9663 (I166163,I166132);
nor I_9664 (I166180,I166050,I166163);
nor I_9665 (I165827,I166180,I165903);
nand I_9666 (I166211,I166163,I166098);
nand I_9667 (I165812,I165920,I166211);
nand I_9668 (I166242,I166002,I166211);
DFFARX1 I_9669 (I166242,I1862,I165835,I165815,);
nand I_9670 (I166273,I166067,I166132);
nor I_9671 (I165809,I165920,I166273);
nor I_9672 (I166304,I166067,I166132);
nand I_9673 (I165818,I166304,I166115);
not I_9674 (I166362,I1869);
or I_9675 (I166379,I357377,I357365);
nand I_9676 (I166396,I357359,I357359);
not I_9677 (I166413,I166396);
nand I_9678 (I166430,I166413,I166379);
not I_9679 (I166447,I166430);
nand I_9680 (I166464,I357362,I357362);
and I_9681 (I166481,I166464,I357368);
DFFARX1 I_9682 (I166481,I1862,I166362,I166507,);
nor I_9683 (I166330,I166507,I166396);
nand I_9684 (I166529,I166447,I166507);
nor I_9685 (I166546,I166507,I166413);
not I_9686 (I166348,I166507);
nor I_9687 (I166577,I357374,I357362);
not I_9688 (I166594,I166577);
nand I_9689 (I166351,I166546,I166577);
not I_9690 (I166625,I357380);
nor I_9691 (I166642,I166507,I357380);
nand I_9692 (I166659,I357365,I357371);
nor I_9693 (I166333,I166659,I166396);
not I_9694 (I166690,I166659);
nor I_9695 (I166707,I166577,I166690);
nor I_9696 (I166354,I166707,I166430);
nand I_9697 (I166738,I166690,I166625);
nand I_9698 (I166339,I166447,I166738);
nand I_9699 (I166769,I166529,I166738);
DFFARX1 I_9700 (I166769,I1862,I166362,I166342,);
nand I_9701 (I166800,I166594,I166659);
nor I_9702 (I166336,I166447,I166800);
nor I_9703 (I166831,I166594,I166659);
nand I_9704 (I166345,I166831,I166642);
not I_9705 (I166889,I1869);
or I_9706 (I166906,I259133,I259136);
nand I_9707 (I166923,I259139,I259148);
not I_9708 (I166940,I166923);
nand I_9709 (I166957,I166940,I166906);
not I_9710 (I166974,I166957);
nand I_9711 (I166991,I259145,I259151);
and I_9712 (I167008,I166991,I259133);
DFFARX1 I_9713 (I167008,I1862,I166889,I167034,);
nor I_9714 (I166857,I167034,I166923);
nand I_9715 (I167056,I166974,I167034);
nor I_9716 (I167073,I167034,I166940);
not I_9717 (I166875,I167034);
nor I_9718 (I167104,I259136,I259151);
not I_9719 (I167121,I167104);
nand I_9720 (I166878,I167073,I167104);
not I_9721 (I167152,I259154);
nor I_9722 (I167169,I167034,I259154);
nand I_9723 (I167186,I259142,I259139);
nor I_9724 (I166860,I167186,I166923);
not I_9725 (I167217,I167186);
nor I_9726 (I167234,I167104,I167217);
nor I_9727 (I166881,I167234,I166957);
nand I_9728 (I167265,I167217,I167152);
nand I_9729 (I166866,I166974,I167265);
nand I_9730 (I167296,I167056,I167265);
DFFARX1 I_9731 (I167296,I1862,I166889,I166869,);
nand I_9732 (I167327,I167121,I167186);
nor I_9733 (I166863,I166974,I167327);
nor I_9734 (I167358,I167121,I167186);
nand I_9735 (I166872,I167358,I167169);
not I_9736 (I167416,I1869);
or I_9737 (I167433,I266273,I266276);
nand I_9738 (I167450,I266279,I266288);
not I_9739 (I167467,I167450);
nand I_9740 (I167484,I167467,I167433);
not I_9741 (I167501,I167484);
nand I_9742 (I167518,I266285,I266291);
and I_9743 (I167535,I167518,I266273);
DFFARX1 I_9744 (I167535,I1862,I167416,I167561,);
nor I_9745 (I167384,I167561,I167450);
nand I_9746 (I167583,I167501,I167561);
nor I_9747 (I167600,I167561,I167467);
not I_9748 (I167402,I167561);
nor I_9749 (I167631,I266276,I266291);
not I_9750 (I167648,I167631);
nand I_9751 (I167405,I167600,I167631);
not I_9752 (I167679,I266294);
nor I_9753 (I167696,I167561,I266294);
nand I_9754 (I167713,I266282,I266279);
nor I_9755 (I167387,I167713,I167450);
not I_9756 (I167744,I167713);
nor I_9757 (I167761,I167631,I167744);
nor I_9758 (I167408,I167761,I167484);
nand I_9759 (I167792,I167744,I167679);
nand I_9760 (I167393,I167501,I167792);
nand I_9761 (I167823,I167583,I167792);
DFFARX1 I_9762 (I167823,I1862,I167416,I167396,);
nand I_9763 (I167854,I167648,I167713);
nor I_9764 (I167390,I167501,I167854);
nor I_9765 (I167885,I167648,I167713);
nand I_9766 (I167399,I167885,I167696);
not I_9767 (I167943,I1869);
or I_9768 (I167960,I378292,I378289);
nand I_9769 (I167977,I378301,I378304);
not I_9770 (I167994,I167977);
nand I_9771 (I168011,I167994,I167960);
not I_9772 (I168028,I168011);
nand I_9773 (I168045,I378295,I378286);
and I_9774 (I168062,I168045,I378286);
DFFARX1 I_9775 (I168062,I1862,I167943,I168088,);
nor I_9776 (I167911,I168088,I167977);
nand I_9777 (I168110,I168028,I168088);
nor I_9778 (I168127,I168088,I167994);
not I_9779 (I167929,I168088);
nor I_9780 (I168158,I378289,I378286);
not I_9781 (I168175,I168158);
nand I_9782 (I167932,I168127,I168158);
not I_9783 (I168206,I378292);
nor I_9784 (I168223,I168088,I378292);
nand I_9785 (I168240,I378295,I378298);
nor I_9786 (I167914,I168240,I167977);
not I_9787 (I168271,I168240);
nor I_9788 (I168288,I168158,I168271);
nor I_9789 (I167935,I168288,I168011);
nand I_9790 (I168319,I168271,I168206);
nand I_9791 (I167920,I168028,I168319);
nand I_9792 (I168350,I168110,I168319);
DFFARX1 I_9793 (I168350,I1862,I167943,I167923,);
nand I_9794 (I168381,I168175,I168240);
nor I_9795 (I167917,I168028,I168381);
nor I_9796 (I168412,I168175,I168240);
nand I_9797 (I167926,I168412,I168223);
not I_9798 (I168470,I1869);
or I_9799 (I168487,I51226,I51223);
nand I_9800 (I168504,I51229,I51226);
not I_9801 (I168521,I168504);
nand I_9802 (I168538,I168521,I168487);
not I_9803 (I168555,I168538);
nand I_9804 (I168572,I51244,I51247);
and I_9805 (I168589,I168572,I51223);
DFFARX1 I_9806 (I168589,I1862,I168470,I168615,);
nor I_9807 (I168438,I168615,I168504);
nand I_9808 (I168637,I168555,I168615);
nor I_9809 (I168654,I168615,I168521);
not I_9810 (I168456,I168615);
nor I_9811 (I168685,I51241,I51247);
not I_9812 (I168702,I168685);
nand I_9813 (I168459,I168654,I168685);
not I_9814 (I168733,I51232);
nor I_9815 (I168750,I168615,I51232);
nand I_9816 (I168767,I51235,I51238);
nor I_9817 (I168441,I168767,I168504);
not I_9818 (I168798,I168767);
nor I_9819 (I168815,I168685,I168798);
nor I_9820 (I168462,I168815,I168538);
nand I_9821 (I168846,I168798,I168733);
nand I_9822 (I168447,I168555,I168846);
nand I_9823 (I168877,I168637,I168846);
DFFARX1 I_9824 (I168877,I1862,I168470,I168450,);
nand I_9825 (I168908,I168702,I168767);
nor I_9826 (I168444,I168555,I168908);
nor I_9827 (I168939,I168702,I168767);
nand I_9828 (I168453,I168939,I168750);
not I_9829 (I168997,I1869);
or I_9830 (I169014,I10831,I10831);
nand I_9831 (I169031,I10837,I10840);
not I_9832 (I169048,I169031);
nand I_9833 (I169065,I169048,I169014);
not I_9834 (I169082,I169065);
nand I_9835 (I169099,I10849,I10852);
and I_9836 (I169116,I169099,I10834);
DFFARX1 I_9837 (I169116,I1862,I168997,I169142,);
nor I_9838 (I168965,I169142,I169031);
nand I_9839 (I169164,I169082,I169142);
nor I_9840 (I169181,I169142,I169048);
not I_9841 (I168983,I169142);
nor I_9842 (I169212,I10846,I10852);
not I_9843 (I169229,I169212);
nand I_9844 (I168986,I169181,I169212);
not I_9845 (I169260,I10834);
nor I_9846 (I169277,I169142,I10834);
nand I_9847 (I169294,I10837,I10843);
nor I_9848 (I168968,I169294,I169031);
not I_9849 (I169325,I169294);
nor I_9850 (I169342,I169212,I169325);
nor I_9851 (I168989,I169342,I169065);
nand I_9852 (I169373,I169325,I169260);
nand I_9853 (I168974,I169082,I169373);
nand I_9854 (I169404,I169164,I169373);
DFFARX1 I_9855 (I169404,I1862,I168997,I168977,);
nand I_9856 (I169435,I169229,I169294);
nor I_9857 (I168971,I169082,I169435);
nor I_9858 (I169466,I169229,I169294);
nand I_9859 (I168980,I169466,I169277);
not I_9860 (I169524,I1869);
or I_9861 (I169541,I298356,I298344);
nand I_9862 (I169558,I298347,I298341);
not I_9863 (I169575,I169558);
nand I_9864 (I169592,I169575,I169541);
not I_9865 (I169609,I169592);
nand I_9866 (I169626,I298338,I298341);
and I_9867 (I169643,I169626,I298335);
DFFARX1 I_9868 (I169643,I1862,I169524,I169669,);
nor I_9869 (I169492,I169669,I169558);
nand I_9870 (I169691,I169609,I169669);
nor I_9871 (I169708,I169669,I169575);
not I_9872 (I169510,I169669);
nor I_9873 (I169739,I298335,I298341);
not I_9874 (I169756,I169739);
nand I_9875 (I169513,I169708,I169739);
not I_9876 (I169787,I298338);
nor I_9877 (I169804,I169669,I298338);
nand I_9878 (I169821,I298353,I298350);
nor I_9879 (I169495,I169821,I169558);
not I_9880 (I169852,I169821);
nor I_9881 (I169869,I169739,I169852);
nor I_9882 (I169516,I169869,I169592);
nand I_9883 (I169900,I169852,I169787);
nand I_9884 (I169501,I169609,I169900);
nand I_9885 (I169931,I169691,I169900);
DFFARX1 I_9886 (I169931,I1862,I169524,I169504,);
nand I_9887 (I169962,I169756,I169821);
nor I_9888 (I169498,I169609,I169962);
nor I_9889 (I169993,I169756,I169821);
nand I_9890 (I169507,I169993,I169804);
not I_9891 (I170051,I1869);
or I_9892 (I170068,I239141,I239144);
nand I_9893 (I170085,I239147,I239156);
not I_9894 (I170102,I170085);
nand I_9895 (I170119,I170102,I170068);
not I_9896 (I170136,I170119);
nand I_9897 (I170153,I239153,I239159);
and I_9898 (I170170,I170153,I239141);
DFFARX1 I_9899 (I170170,I1862,I170051,I170196,);
nor I_9900 (I170019,I170196,I170085);
nand I_9901 (I170218,I170136,I170196);
nor I_9902 (I170235,I170196,I170102);
not I_9903 (I170037,I170196);
nor I_9904 (I170266,I239144,I239159);
not I_9905 (I170283,I170266);
nand I_9906 (I170040,I170235,I170266);
not I_9907 (I170314,I239162);
nor I_9908 (I170331,I170196,I239162);
nand I_9909 (I170348,I239150,I239147);
nor I_9910 (I170022,I170348,I170085);
not I_9911 (I170379,I170348);
nor I_9912 (I170396,I170266,I170379);
nor I_9913 (I170043,I170396,I170119);
nand I_9914 (I170427,I170379,I170314);
nand I_9915 (I170028,I170136,I170427);
nand I_9916 (I170458,I170218,I170427);
DFFARX1 I_9917 (I170458,I1862,I170051,I170031,);
nand I_9918 (I170489,I170283,I170348);
nor I_9919 (I170025,I170136,I170489);
nor I_9920 (I170520,I170283,I170348);
nand I_9921 (I170034,I170520,I170331);
not I_9922 (I170578,I1869);
or I_9923 (I170595,I111205,I111214);
nand I_9924 (I170612,I111208,I111211);
not I_9925 (I170629,I170612);
nand I_9926 (I170646,I170629,I170595);
not I_9927 (I170663,I170646);
nand I_9928 (I170680,I111202,I111202);
and I_9929 (I170697,I170680,I111199);
DFFARX1 I_9930 (I170697,I1862,I170578,I170723,);
nor I_9931 (I170546,I170723,I170612);
nand I_9932 (I170745,I170663,I170723);
nor I_9933 (I170762,I170723,I170629);
not I_9934 (I170564,I170723);
nor I_9935 (I170793,I111217,I111202);
not I_9936 (I170810,I170793);
nand I_9937 (I170567,I170762,I170793);
not I_9938 (I170841,I111205);
nor I_9939 (I170858,I170723,I111205);
nand I_9940 (I170875,I111208,I111199);
nor I_9941 (I170549,I170875,I170612);
not I_9942 (I170906,I170875);
nor I_9943 (I170923,I170793,I170906);
nor I_9944 (I170570,I170923,I170646);
nand I_9945 (I170954,I170906,I170841);
nand I_9946 (I170555,I170663,I170954);
nand I_9947 (I170985,I170745,I170954);
DFFARX1 I_9948 (I170985,I1862,I170578,I170558,);
nand I_9949 (I171016,I170810,I170875);
nor I_9950 (I170552,I170663,I171016);
nor I_9951 (I171047,I170810,I170875);
nand I_9952 (I170561,I171047,I170858);
not I_9953 (I171105,I1869);
or I_9954 (I171122,I241045,I241048);
nand I_9955 (I171139,I241051,I241060);
not I_9956 (I171156,I171139);
nand I_9957 (I171173,I171156,I171122);
not I_9958 (I171190,I171173);
nand I_9959 (I171207,I241057,I241063);
and I_9960 (I171224,I171207,I241045);
DFFARX1 I_9961 (I171224,I1862,I171105,I171250,);
nor I_9962 (I171073,I171250,I171139);
nand I_9963 (I171272,I171190,I171250);
nor I_9964 (I171289,I171250,I171156);
not I_9965 (I171091,I171250);
nor I_9966 (I171320,I241048,I241063);
not I_9967 (I171337,I171320);
nand I_9968 (I171094,I171289,I171320);
not I_9969 (I171368,I241066);
nor I_9970 (I171385,I171250,I241066);
nand I_9971 (I171402,I241054,I241051);
nor I_9972 (I171076,I171402,I171139);
not I_9973 (I171433,I171402);
nor I_9974 (I171450,I171320,I171433);
nor I_9975 (I171097,I171450,I171173);
nand I_9976 (I171481,I171433,I171368);
nand I_9977 (I171082,I171190,I171481);
nand I_9978 (I171512,I171272,I171481);
DFFARX1 I_9979 (I171512,I1862,I171105,I171085,);
nand I_9980 (I171543,I171337,I171402);
nor I_9981 (I171079,I171190,I171543);
nor I_9982 (I171574,I171337,I171402);
nand I_9983 (I171088,I171574,I171385);
not I_9984 (I171632,I1869);
or I_9985 (I171649,I365032,I365029);
nand I_9986 (I171666,I365041,I365044);
not I_9987 (I171683,I171666);
nand I_9988 (I171700,I171683,I171649);
not I_9989 (I171717,I171700);
nand I_9990 (I171734,I365035,I365026);
and I_9991 (I171751,I171734,I365026);
DFFARX1 I_9992 (I171751,I1862,I171632,I171777,);
nor I_9993 (I171600,I171777,I171666);
nand I_9994 (I171799,I171717,I171777);
nor I_9995 (I171816,I171777,I171683);
not I_9996 (I171618,I171777);
nor I_9997 (I171847,I365029,I365026);
not I_9998 (I171864,I171847);
nand I_9999 (I171621,I171816,I171847);
not I_10000 (I171895,I365032);
nor I_10001 (I171912,I171777,I365032);
nand I_10002 (I171929,I365035,I365038);
nor I_10003 (I171603,I171929,I171666);
not I_10004 (I171960,I171929);
nor I_10005 (I171977,I171847,I171960);
nor I_10006 (I171624,I171977,I171700);
nand I_10007 (I172008,I171960,I171895);
nand I_10008 (I171609,I171717,I172008);
nand I_10009 (I172039,I171799,I172008);
DFFARX1 I_10010 (I172039,I1862,I171632,I171612,);
nand I_10011 (I172070,I171864,I171929);
nor I_10012 (I171606,I171717,I172070);
nor I_10013 (I172101,I171864,I171929);
nand I_10014 (I171615,I172101,I171912);
not I_10015 (I172159,I1869);
or I_10016 (I172176,I259609,I259612);
nand I_10017 (I172193,I259615,I259624);
not I_10018 (I172210,I172193);
nand I_10019 (I172227,I172210,I172176);
not I_10020 (I172244,I172227);
nand I_10021 (I172261,I259621,I259627);
and I_10022 (I172278,I172261,I259609);
DFFARX1 I_10023 (I172278,I1862,I172159,I172304,);
nor I_10024 (I172127,I172304,I172193);
nand I_10025 (I172326,I172244,I172304);
nor I_10026 (I172343,I172304,I172210);
not I_10027 (I172145,I172304);
nor I_10028 (I172374,I259612,I259627);
not I_10029 (I172391,I172374);
nand I_10030 (I172148,I172343,I172374);
not I_10031 (I172422,I259630);
nor I_10032 (I172439,I172304,I259630);
nand I_10033 (I172456,I259618,I259615);
nor I_10034 (I172130,I172456,I172193);
not I_10035 (I172487,I172456);
nor I_10036 (I172504,I172374,I172487);
nor I_10037 (I172151,I172504,I172227);
nand I_10038 (I172535,I172487,I172422);
nand I_10039 (I172136,I172244,I172535);
nand I_10040 (I172566,I172326,I172535);
DFFARX1 I_10041 (I172566,I1862,I172159,I172139,);
nand I_10042 (I172597,I172391,I172456);
nor I_10043 (I172133,I172244,I172597);
nor I_10044 (I172628,I172391,I172456);
nand I_10045 (I172142,I172628,I172439);
not I_10046 (I172686,I1869);
or I_10047 (I172703,I326811,I326799);
nand I_10048 (I172720,I326793,I326793);
not I_10049 (I172737,I172720);
nand I_10050 (I172754,I172737,I172703);
not I_10051 (I172771,I172754);
nand I_10052 (I172788,I326796,I326796);
and I_10053 (I172805,I172788,I326802);
DFFARX1 I_10054 (I172805,I1862,I172686,I172831,);
nor I_10055 (I172654,I172831,I172720);
nand I_10056 (I172853,I172771,I172831);
nor I_10057 (I172870,I172831,I172737);
not I_10058 (I172672,I172831);
nor I_10059 (I172901,I326808,I326796);
not I_10060 (I172918,I172901);
nand I_10061 (I172675,I172870,I172901);
not I_10062 (I172949,I326814);
nor I_10063 (I172966,I172831,I326814);
nand I_10064 (I172983,I326799,I326805);
nor I_10065 (I172657,I172983,I172720);
not I_10066 (I173014,I172983);
nor I_10067 (I173031,I172901,I173014);
nor I_10068 (I172678,I173031,I172754);
nand I_10069 (I173062,I173014,I172949);
nand I_10070 (I172663,I172771,I173062);
nand I_10071 (I173093,I172853,I173062);
DFFARX1 I_10072 (I173093,I1862,I172686,I172666,);
nand I_10073 (I173124,I172918,I172983);
nor I_10074 (I172660,I172771,I173124);
nor I_10075 (I173155,I172918,I172983);
nand I_10076 (I172669,I173155,I172966);
not I_10077 (I173213,I1869);
or I_10078 (I173230,I389784,I389781);
nand I_10079 (I173247,I389793,I389796);
not I_10080 (I173264,I173247);
nand I_10081 (I173281,I173264,I173230);
not I_10082 (I173298,I173281);
nand I_10083 (I173315,I389787,I389778);
and I_10084 (I173332,I173315,I389778);
DFFARX1 I_10085 (I173332,I1862,I173213,I173358,);
nor I_10086 (I173181,I173358,I173247);
nand I_10087 (I173380,I173298,I173358);
nor I_10088 (I173397,I173358,I173264);
not I_10089 (I173199,I173358);
nor I_10090 (I173428,I389781,I389778);
not I_10091 (I173445,I173428);
nand I_10092 (I173202,I173397,I173428);
not I_10093 (I173476,I389784);
nor I_10094 (I173493,I173358,I389784);
nand I_10095 (I173510,I389787,I389790);
nor I_10096 (I173184,I173510,I173247);
not I_10097 (I173541,I173510);
nor I_10098 (I173558,I173428,I173541);
nor I_10099 (I173205,I173558,I173281);
nand I_10100 (I173589,I173541,I173476);
nand I_10101 (I173190,I173298,I173589);
nand I_10102 (I173620,I173380,I173589);
DFFARX1 I_10103 (I173620,I1862,I173213,I173193,);
nand I_10104 (I173651,I173445,I173510);
nor I_10105 (I173187,I173298,I173651);
nor I_10106 (I173682,I173445,I173510);
nand I_10107 (I173196,I173682,I173493);
not I_10108 (I173740,I1869);
or I_10109 (I173757,I407464,I407461);
nand I_10110 (I173774,I407473,I407476);
not I_10111 (I173791,I173774);
nand I_10112 (I173808,I173791,I173757);
not I_10113 (I173825,I173808);
nand I_10114 (I173842,I407467,I407458);
and I_10115 (I173859,I173842,I407458);
DFFARX1 I_10116 (I173859,I1862,I173740,I173885,);
nor I_10117 (I173708,I173885,I173774);
nand I_10118 (I173907,I173825,I173885);
nor I_10119 (I173924,I173885,I173791);
not I_10120 (I173726,I173885);
nor I_10121 (I173955,I407461,I407458);
not I_10122 (I173972,I173955);
nand I_10123 (I173729,I173924,I173955);
not I_10124 (I174003,I407464);
nor I_10125 (I174020,I173885,I407464);
nand I_10126 (I174037,I407467,I407470);
nor I_10127 (I173711,I174037,I173774);
not I_10128 (I174068,I174037);
nor I_10129 (I174085,I173955,I174068);
nor I_10130 (I173732,I174085,I173808);
nand I_10131 (I174116,I174068,I174003);
nand I_10132 (I173717,I173825,I174116);
nand I_10133 (I174147,I173907,I174116);
DFFARX1 I_10134 (I174147,I1862,I173740,I173720,);
nand I_10135 (I174178,I173972,I174037);
nor I_10136 (I173714,I173825,I174178);
nor I_10137 (I174209,I173972,I174037);
nand I_10138 (I173723,I174209,I174020);
not I_10139 (I174267,I1869);
or I_10140 (I174284,I338932,I338920);
nand I_10141 (I174301,I338914,I338914);
not I_10142 (I174318,I174301);
nand I_10143 (I174335,I174318,I174284);
not I_10144 (I174352,I174335);
nand I_10145 (I174369,I338917,I338917);
and I_10146 (I174386,I174369,I338923);
DFFARX1 I_10147 (I174386,I1862,I174267,I174412,);
nor I_10148 (I174235,I174412,I174301);
nand I_10149 (I174434,I174352,I174412);
nor I_10150 (I174451,I174412,I174318);
not I_10151 (I174253,I174412);
nor I_10152 (I174482,I338929,I338917);
not I_10153 (I174499,I174482);
nand I_10154 (I174256,I174451,I174482);
not I_10155 (I174530,I338935);
nor I_10156 (I174547,I174412,I338935);
nand I_10157 (I174564,I338920,I338926);
nor I_10158 (I174238,I174564,I174301);
not I_10159 (I174595,I174564);
nor I_10160 (I174612,I174482,I174595);
nor I_10161 (I174259,I174612,I174335);
nand I_10162 (I174643,I174595,I174530);
nand I_10163 (I174244,I174352,I174643);
nand I_10164 (I174674,I174434,I174643);
DFFARX1 I_10165 (I174674,I1862,I174267,I174247,);
nand I_10166 (I174705,I174499,I174564);
nor I_10167 (I174241,I174352,I174705);
nor I_10168 (I174736,I174499,I174564);
nand I_10169 (I174250,I174736,I174547);
not I_10170 (I174794,I1869);
or I_10171 (I174811,I95596,I95593);
nand I_10172 (I174828,I95599,I95596);
not I_10173 (I174845,I174828);
nand I_10174 (I174862,I174845,I174811);
not I_10175 (I174879,I174862);
nand I_10176 (I174896,I95614,I95617);
and I_10177 (I174913,I174896,I95593);
DFFARX1 I_10178 (I174913,I1862,I174794,I174939,);
nor I_10179 (I174762,I174939,I174828);
nand I_10180 (I174961,I174879,I174939);
nor I_10181 (I174978,I174939,I174845);
not I_10182 (I174780,I174939);
nor I_10183 (I175009,I95611,I95617);
not I_10184 (I175026,I175009);
nand I_10185 (I174783,I174978,I175009);
not I_10186 (I175057,I95602);
nor I_10187 (I175074,I174939,I95602);
nand I_10188 (I175091,I95605,I95608);
nor I_10189 (I174765,I175091,I174828);
not I_10190 (I175122,I175091);
nor I_10191 (I175139,I175009,I175122);
nor I_10192 (I174786,I175139,I174862);
nand I_10193 (I175170,I175122,I175057);
nand I_10194 (I174771,I174879,I175170);
nand I_10195 (I175201,I174961,I175170);
DFFARX1 I_10196 (I175201,I1862,I174794,I174774,);
nand I_10197 (I175232,I175026,I175091);
nor I_10198 (I174768,I174879,I175232);
nor I_10199 (I175263,I175026,I175091);
nand I_10200 (I174777,I175263,I175074);
not I_10201 (I175321,I1869);
or I_10202 (I175338,I352634,I352622);
nand I_10203 (I175355,I352616,I352616);
not I_10204 (I175372,I175355);
nand I_10205 (I175389,I175372,I175338);
not I_10206 (I175406,I175389);
nand I_10207 (I175423,I352619,I352619);
and I_10208 (I175440,I175423,I352625);
DFFARX1 I_10209 (I175440,I1862,I175321,I175466,);
nor I_10210 (I175289,I175466,I175355);
nand I_10211 (I175488,I175406,I175466);
nor I_10212 (I175505,I175466,I175372);
not I_10213 (I175307,I175466);
nor I_10214 (I175536,I352631,I352619);
not I_10215 (I175553,I175536);
nand I_10216 (I175310,I175505,I175536);
not I_10217 (I175584,I352637);
nor I_10218 (I175601,I175466,I352637);
nand I_10219 (I175618,I352622,I352628);
nor I_10220 (I175292,I175618,I175355);
not I_10221 (I175649,I175618);
nor I_10222 (I175666,I175536,I175649);
nor I_10223 (I175313,I175666,I175389);
nand I_10224 (I175697,I175649,I175584);
nand I_10225 (I175298,I175406,I175697);
nand I_10226 (I175728,I175488,I175697);
DFFARX1 I_10227 (I175728,I1862,I175321,I175301,);
nand I_10228 (I175759,I175553,I175618);
nor I_10229 (I175295,I175406,I175759);
nor I_10230 (I175790,I175553,I175618);
nand I_10231 (I175304,I175790,I175601);
not I_10232 (I175848,I1869);
or I_10233 (I175865,I262465,I262468);
nand I_10234 (I175882,I262471,I262480);
not I_10235 (I175899,I175882);
nand I_10236 (I175916,I175899,I175865);
not I_10237 (I175933,I175916);
nand I_10238 (I175950,I262477,I262483);
and I_10239 (I175967,I175950,I262465);
DFFARX1 I_10240 (I175967,I1862,I175848,I175993,);
nor I_10241 (I175816,I175993,I175882);
nand I_10242 (I176015,I175933,I175993);
nor I_10243 (I176032,I175993,I175899);
not I_10244 (I175834,I175993);
nor I_10245 (I176063,I262468,I262483);
not I_10246 (I176080,I176063);
nand I_10247 (I175837,I176032,I176063);
not I_10248 (I176111,I262486);
nor I_10249 (I176128,I175993,I262486);
nand I_10250 (I176145,I262474,I262471);
nor I_10251 (I175819,I176145,I175882);
not I_10252 (I176176,I176145);
nor I_10253 (I176193,I176063,I176176);
nor I_10254 (I175840,I176193,I175916);
nand I_10255 (I176224,I176176,I176111);
nand I_10256 (I175825,I175933,I176224);
nand I_10257 (I176255,I176015,I176224);
DFFARX1 I_10258 (I176255,I1862,I175848,I175828,);
nand I_10259 (I176286,I176080,I176145);
nor I_10260 (I175822,I175933,I176286);
nor I_10261 (I176317,I176080,I176145);
nand I_10262 (I175831,I176317,I176128);
not I_10263 (I176375,I1869);
or I_10264 (I176392,I221053,I221056);
nand I_10265 (I176409,I221059,I221068);
not I_10266 (I176426,I176409);
nand I_10267 (I176443,I176426,I176392);
not I_10268 (I176460,I176443);
nand I_10269 (I176477,I221065,I221071);
and I_10270 (I176494,I176477,I221053);
DFFARX1 I_10271 (I176494,I1862,I176375,I176520,);
nor I_10272 (I176343,I176520,I176409);
nand I_10273 (I176542,I176460,I176520);
nor I_10274 (I176559,I176520,I176426);
not I_10275 (I176361,I176520);
nor I_10276 (I176590,I221056,I221071);
not I_10277 (I176607,I176590);
nand I_10278 (I176364,I176559,I176590);
not I_10279 (I176638,I221074);
nor I_10280 (I176655,I176520,I221074);
nand I_10281 (I176672,I221062,I221059);
nor I_10282 (I176346,I176672,I176409);
not I_10283 (I176703,I176672);
nor I_10284 (I176720,I176590,I176703);
nor I_10285 (I176367,I176720,I176443);
nand I_10286 (I176751,I176703,I176638);
nand I_10287 (I176352,I176460,I176751);
nand I_10288 (I176782,I176542,I176751);
DFFARX1 I_10289 (I176782,I1862,I176375,I176355,);
nand I_10290 (I176813,I176607,I176672);
nor I_10291 (I176349,I176460,I176813);
nor I_10292 (I176844,I176607,I176672);
nand I_10293 (I176358,I176844,I176655);
not I_10294 (I176902,I1869);
or I_10295 (I176919,I74686,I74683);
nand I_10296 (I176936,I74689,I74686);
not I_10297 (I176953,I176936);
nand I_10298 (I176970,I176953,I176919);
not I_10299 (I176987,I176970);
nand I_10300 (I177004,I74704,I74707);
and I_10301 (I177021,I177004,I74683);
DFFARX1 I_10302 (I177021,I1862,I176902,I177047,);
nor I_10303 (I176870,I177047,I176936);
nand I_10304 (I177069,I176987,I177047);
nor I_10305 (I177086,I177047,I176953);
not I_10306 (I176888,I177047);
nor I_10307 (I177117,I74701,I74707);
not I_10308 (I177134,I177117);
nand I_10309 (I176891,I177086,I177117);
not I_10310 (I177165,I74692);
nor I_10311 (I177182,I177047,I74692);
nand I_10312 (I177199,I74695,I74698);
nor I_10313 (I176873,I177199,I176936);
not I_10314 (I177230,I177199);
nor I_10315 (I177247,I177117,I177230);
nor I_10316 (I176894,I177247,I176970);
nand I_10317 (I177278,I177230,I177165);
nand I_10318 (I176879,I176987,I177278);
nand I_10319 (I177309,I177069,I177278);
DFFARX1 I_10320 (I177309,I1862,I176902,I176882,);
nand I_10321 (I177340,I177134,I177199);
nor I_10322 (I176876,I176987,I177340);
nor I_10323 (I177371,I177134,I177199);
nand I_10324 (I176885,I177371,I177182);
not I_10325 (I177429,I1869);
or I_10326 (I177446,I23176,I23173);
nand I_10327 (I177463,I23179,I23176);
not I_10328 (I177480,I177463);
nand I_10329 (I177497,I177480,I177446);
not I_10330 (I177514,I177497);
nand I_10331 (I177531,I23194,I23197);
and I_10332 (I177548,I177531,I23173);
DFFARX1 I_10333 (I177548,I1862,I177429,I177574,);
nor I_10334 (I177397,I177574,I177463);
nand I_10335 (I177596,I177514,I177574);
nor I_10336 (I177613,I177574,I177480);
not I_10337 (I177415,I177574);
nor I_10338 (I177644,I23191,I23197);
not I_10339 (I177661,I177644);
nand I_10340 (I177418,I177613,I177644);
not I_10341 (I177692,I23182);
nor I_10342 (I177709,I177574,I23182);
nand I_10343 (I177726,I23185,I23188);
nor I_10344 (I177400,I177726,I177463);
not I_10345 (I177757,I177726);
nor I_10346 (I177774,I177644,I177757);
nor I_10347 (I177421,I177774,I177497);
nand I_10348 (I177805,I177757,I177692);
nand I_10349 (I177406,I177514,I177805);
nand I_10350 (I177836,I177596,I177805);
DFFARX1 I_10351 (I177836,I1862,I177429,I177409,);
nand I_10352 (I177867,I177661,I177726);
nor I_10353 (I177403,I177514,I177867);
nor I_10354 (I177898,I177661,I177726);
nand I_10355 (I177412,I177898,I177709);
not I_10356 (I177956,I1869);
or I_10357 (I177973,I75196,I75193);
nand I_10358 (I177990,I75199,I75196);
not I_10359 (I178007,I177990);
nand I_10360 (I178024,I178007,I177973);
not I_10361 (I178041,I178024);
nand I_10362 (I178058,I75214,I75217);
and I_10363 (I178075,I178058,I75193);
DFFARX1 I_10364 (I178075,I1862,I177956,I178101,);
nor I_10365 (I177924,I178101,I177990);
nand I_10366 (I178123,I178041,I178101);
nor I_10367 (I178140,I178101,I178007);
not I_10368 (I177942,I178101);
nor I_10369 (I178171,I75211,I75217);
not I_10370 (I178188,I178171);
nand I_10371 (I177945,I178140,I178171);
not I_10372 (I178219,I75202);
nor I_10373 (I178236,I178101,I75202);
nand I_10374 (I178253,I75205,I75208);
nor I_10375 (I177927,I178253,I177990);
not I_10376 (I178284,I178253);
nor I_10377 (I178301,I178171,I178284);
nor I_10378 (I177948,I178301,I178024);
nand I_10379 (I178332,I178284,I178219);
nand I_10380 (I177933,I178041,I178332);
nand I_10381 (I178363,I178123,I178332);
DFFARX1 I_10382 (I178363,I1862,I177956,I177936,);
nand I_10383 (I178394,I178188,I178253);
nor I_10384 (I177930,I178041,I178394);
nor I_10385 (I178425,I178188,I178253);
nand I_10386 (I177939,I178425,I178236);
not I_10387 (I178483,I1869);
or I_10388 (I178500,I100696,I100693);
nand I_10389 (I178517,I100699,I100696);
not I_10390 (I178534,I178517);
nand I_10391 (I178551,I178534,I178500);
not I_10392 (I178568,I178551);
nand I_10393 (I178585,I100714,I100717);
and I_10394 (I178602,I178585,I100693);
DFFARX1 I_10395 (I178602,I1862,I178483,I178628,);
nor I_10396 (I178451,I178628,I178517);
nand I_10397 (I178650,I178568,I178628);
nor I_10398 (I178667,I178628,I178534);
not I_10399 (I178469,I178628);
nor I_10400 (I178698,I100711,I100717);
not I_10401 (I178715,I178698);
nand I_10402 (I178472,I178667,I178698);
not I_10403 (I178746,I100702);
nor I_10404 (I178763,I178628,I100702);
nand I_10405 (I178780,I100705,I100708);
nor I_10406 (I178454,I178780,I178517);
not I_10407 (I178811,I178780);
nor I_10408 (I178828,I178698,I178811);
nor I_10409 (I178475,I178828,I178551);
nand I_10410 (I178859,I178811,I178746);
nand I_10411 (I178460,I178568,I178859);
nand I_10412 (I178890,I178650,I178859);
DFFARX1 I_10413 (I178890,I1862,I178483,I178463,);
nand I_10414 (I178921,I178715,I178780);
nor I_10415 (I178457,I178568,I178921);
nor I_10416 (I178952,I178715,I178780);
nand I_10417 (I178466,I178952,I178763);
not I_10418 (I179010,I1869);
or I_10419 (I179027,I254373,I254376);
nand I_10420 (I179044,I254379,I254388);
not I_10421 (I179061,I179044);
nand I_10422 (I179078,I179061,I179027);
not I_10423 (I179095,I179078);
nand I_10424 (I179112,I254385,I254391);
and I_10425 (I179129,I179112,I254373);
DFFARX1 I_10426 (I179129,I1862,I179010,I179155,);
nor I_10427 (I178978,I179155,I179044);
nand I_10428 (I179177,I179095,I179155);
nor I_10429 (I179194,I179155,I179061);
not I_10430 (I178996,I179155);
nor I_10431 (I179225,I254376,I254391);
not I_10432 (I179242,I179225);
nand I_10433 (I178999,I179194,I179225);
not I_10434 (I179273,I254394);
nor I_10435 (I179290,I179155,I254394);
nand I_10436 (I179307,I254382,I254379);
nor I_10437 (I178981,I179307,I179044);
not I_10438 (I179338,I179307);
nor I_10439 (I179355,I179225,I179338);
nor I_10440 (I179002,I179355,I179078);
nand I_10441 (I179386,I179338,I179273);
nand I_10442 (I178987,I179095,I179386);
nand I_10443 (I179417,I179177,I179386);
DFFARX1 I_10444 (I179417,I1862,I179010,I178990,);
nand I_10445 (I179448,I179242,I179307);
nor I_10446 (I178984,I179095,I179448);
nor I_10447 (I179479,I179242,I179307);
nand I_10448 (I178993,I179479,I179290);
not I_10449 (I179537,I1869);
or I_10450 (I179554,I307839,I307827);
nand I_10451 (I179571,I307821,I307821);
not I_10452 (I179588,I179571);
nand I_10453 (I179605,I179588,I179554);
not I_10454 (I179622,I179605);
nand I_10455 (I179639,I307824,I307824);
and I_10456 (I179656,I179639,I307830);
DFFARX1 I_10457 (I179656,I1862,I179537,I179682,);
nor I_10458 (I179505,I179682,I179571);
nand I_10459 (I179704,I179622,I179682);
nor I_10460 (I179721,I179682,I179588);
not I_10461 (I179523,I179682);
nor I_10462 (I179752,I307836,I307824);
not I_10463 (I179769,I179752);
nand I_10464 (I179526,I179721,I179752);
not I_10465 (I179800,I307842);
nor I_10466 (I179817,I179682,I307842);
nand I_10467 (I179834,I307827,I307833);
nor I_10468 (I179508,I179834,I179571);
not I_10469 (I179865,I179834);
nor I_10470 (I179882,I179752,I179865);
nor I_10471 (I179529,I179882,I179605);
nand I_10472 (I179913,I179865,I179800);
nand I_10473 (I179514,I179622,I179913);
nand I_10474 (I179944,I179704,I179913);
DFFARX1 I_10475 (I179944,I1862,I179537,I179517,);
nand I_10476 (I179975,I179769,I179834);
nor I_10477 (I179511,I179622,I179975);
nor I_10478 (I180006,I179769,I179834);
nand I_10479 (I179520,I180006,I179817);
not I_10480 (I180064,I1869);
or I_10481 (I180081,I277221,I277224);
nand I_10482 (I180098,I277227,I277236);
not I_10483 (I180115,I180098);
nand I_10484 (I180132,I180115,I180081);
not I_10485 (I180149,I180132);
nand I_10486 (I180166,I277233,I277239);
and I_10487 (I180183,I180166,I277221);
DFFARX1 I_10488 (I180183,I1862,I180064,I180209,);
nor I_10489 (I180032,I180209,I180098);
nand I_10490 (I180231,I180149,I180209);
nor I_10491 (I180248,I180209,I180115);
not I_10492 (I180050,I180209);
nor I_10493 (I180279,I277224,I277239);
not I_10494 (I180296,I180279);
nand I_10495 (I180053,I180248,I180279);
not I_10496 (I180327,I277242);
nor I_10497 (I180344,I180209,I277242);
nand I_10498 (I180361,I277230,I277227);
nor I_10499 (I180035,I180361,I180098);
not I_10500 (I180392,I180361);
nor I_10501 (I180409,I180279,I180392);
nor I_10502 (I180056,I180409,I180132);
nand I_10503 (I180440,I180392,I180327);
nand I_10504 (I180041,I180149,I180440);
nand I_10505 (I180471,I180231,I180440);
DFFARX1 I_10506 (I180471,I1862,I180064,I180044,);
nand I_10507 (I180502,I180296,I180361);
nor I_10508 (I180038,I180149,I180502);
nor I_10509 (I180533,I180296,I180361);
nand I_10510 (I180047,I180533,I180344);
not I_10511 (I180591,I1869);
or I_10512 (I180608,I77236,I77233);
nand I_10513 (I180625,I77239,I77236);
not I_10514 (I180642,I180625);
nand I_10515 (I180659,I180642,I180608);
not I_10516 (I180676,I180659);
nand I_10517 (I180693,I77254,I77257);
and I_10518 (I180710,I180693,I77233);
DFFARX1 I_10519 (I180710,I1862,I180591,I180736,);
nor I_10520 (I180559,I180736,I180625);
nand I_10521 (I180758,I180676,I180736);
nor I_10522 (I180775,I180736,I180642);
not I_10523 (I180577,I180736);
nor I_10524 (I180806,I77251,I77257);
not I_10525 (I180823,I180806);
nand I_10526 (I180580,I180775,I180806);
not I_10527 (I180854,I77242);
nor I_10528 (I180871,I180736,I77242);
nand I_10529 (I180888,I77245,I77248);
nor I_10530 (I180562,I180888,I180625);
not I_10531 (I180919,I180888);
nor I_10532 (I180936,I180806,I180919);
nor I_10533 (I180583,I180936,I180659);
nand I_10534 (I180967,I180919,I180854);
nand I_10535 (I180568,I180676,I180967);
nand I_10536 (I180998,I180758,I180967);
DFFARX1 I_10537 (I180998,I1862,I180591,I180571,);
nand I_10538 (I181029,I180823,I180888);
nor I_10539 (I180565,I180676,I181029);
nor I_10540 (I181060,I180823,I180888);
nand I_10541 (I180574,I181060,I180871);
not I_10542 (I181118,I1869);
or I_10543 (I181135,I377850,I377847);
nand I_10544 (I181152,I377859,I377862);
not I_10545 (I181169,I181152);
nand I_10546 (I181186,I181169,I181135);
not I_10547 (I181203,I181186);
nand I_10548 (I181220,I377853,I377844);
and I_10549 (I181237,I181220,I377844);
DFFARX1 I_10550 (I181237,I1862,I181118,I181263,);
nor I_10551 (I181086,I181263,I181152);
nand I_10552 (I181285,I181203,I181263);
nor I_10553 (I181302,I181263,I181169);
not I_10554 (I181104,I181263);
nor I_10555 (I181333,I377847,I377844);
not I_10556 (I181350,I181333);
nand I_10557 (I181107,I181302,I181333);
not I_10558 (I181381,I377850);
nor I_10559 (I181398,I181263,I377850);
nand I_10560 (I181415,I377853,I377856);
nor I_10561 (I181089,I181415,I181152);
not I_10562 (I181446,I181415);
nor I_10563 (I181463,I181333,I181446);
nor I_10564 (I181110,I181463,I181186);
nand I_10565 (I181494,I181446,I181381);
nand I_10566 (I181095,I181203,I181494);
nand I_10567 (I181525,I181285,I181494);
DFFARX1 I_10568 (I181525,I1862,I181118,I181098,);
nand I_10569 (I181556,I181350,I181415);
nor I_10570 (I181092,I181203,I181556);
nor I_10571 (I181587,I181350,I181415);
nand I_10572 (I181101,I181587,I181398);
not I_10573 (I181645,I1869);
or I_10574 (I181662,I287289,I287277);
nand I_10575 (I181679,I287280,I287274);
not I_10576 (I181696,I181679);
nand I_10577 (I181713,I181696,I181662);
not I_10578 (I181730,I181713);
nand I_10579 (I181747,I287271,I287274);
and I_10580 (I181764,I181747,I287268);
DFFARX1 I_10581 (I181764,I1862,I181645,I181790,);
nor I_10582 (I181613,I181790,I181679);
nand I_10583 (I181812,I181730,I181790);
nor I_10584 (I181829,I181790,I181696);
not I_10585 (I181631,I181790);
nor I_10586 (I181860,I287268,I287274);
not I_10587 (I181877,I181860);
nand I_10588 (I181634,I181829,I181860);
not I_10589 (I181908,I287271);
nor I_10590 (I181925,I181790,I287271);
nand I_10591 (I181942,I287286,I287283);
nor I_10592 (I181616,I181942,I181679);
not I_10593 (I181973,I181942);
nor I_10594 (I181990,I181860,I181973);
nor I_10595 (I181637,I181990,I181713);
nand I_10596 (I182021,I181973,I181908);
nand I_10597 (I181622,I181730,I182021);
nand I_10598 (I182052,I181812,I182021);
DFFARX1 I_10599 (I182052,I1862,I181645,I181625,);
nand I_10600 (I182083,I181877,I181942);
nor I_10601 (I181619,I181730,I182083);
nor I_10602 (I182114,I181877,I181942);
nand I_10603 (I181628,I182114,I181925);
not I_10604 (I182172,I1869);
or I_10605 (I182189,I346310,I346298);
nand I_10606 (I182206,I346292,I346292);
not I_10607 (I182223,I182206);
nand I_10608 (I182240,I182223,I182189);
not I_10609 (I182257,I182240);
nand I_10610 (I182274,I346295,I346295);
and I_10611 (I182291,I182274,I346301);
DFFARX1 I_10612 (I182291,I1862,I182172,I182317,);
nor I_10613 (I182140,I182317,I182206);
nand I_10614 (I182339,I182257,I182317);
nor I_10615 (I182356,I182317,I182223);
not I_10616 (I182158,I182317);
nor I_10617 (I182387,I346307,I346295);
not I_10618 (I182404,I182387);
nand I_10619 (I182161,I182356,I182387);
not I_10620 (I182435,I346313);
nor I_10621 (I182452,I182317,I346313);
nand I_10622 (I182469,I346298,I346304);
nor I_10623 (I182143,I182469,I182206);
not I_10624 (I182500,I182469);
nor I_10625 (I182517,I182387,I182500);
nor I_10626 (I182164,I182517,I182240);
nand I_10627 (I182548,I182500,I182435);
nand I_10628 (I182149,I182257,I182548);
nand I_10629 (I182579,I182339,I182548);
DFFARX1 I_10630 (I182579,I1862,I182172,I182152,);
nand I_10631 (I182610,I182404,I182469);
nor I_10632 (I182146,I182257,I182610);
nor I_10633 (I182641,I182404,I182469);
nand I_10634 (I182155,I182641,I182452);
not I_10635 (I182699,I1869);
or I_10636 (I182716,I300464,I300452);
nand I_10637 (I182733,I300455,I300449);
not I_10638 (I182750,I182733);
nand I_10639 (I182767,I182750,I182716);
not I_10640 (I182784,I182767);
nand I_10641 (I182801,I300446,I300449);
and I_10642 (I182818,I182801,I300443);
DFFARX1 I_10643 (I182818,I1862,I182699,I182844,);
nor I_10644 (I182667,I182844,I182733);
nand I_10645 (I182866,I182784,I182844);
nor I_10646 (I182883,I182844,I182750);
not I_10647 (I182685,I182844);
nor I_10648 (I182914,I300443,I300449);
not I_10649 (I182931,I182914);
nand I_10650 (I182688,I182883,I182914);
not I_10651 (I182962,I300446);
nor I_10652 (I182979,I182844,I300446);
nand I_10653 (I182996,I300461,I300458);
nor I_10654 (I182670,I182996,I182733);
not I_10655 (I183027,I182996);
nor I_10656 (I183044,I182914,I183027);
nor I_10657 (I182691,I183044,I182767);
nand I_10658 (I183075,I183027,I182962);
nand I_10659 (I182676,I182784,I183075);
nand I_10660 (I183106,I182866,I183075);
DFFARX1 I_10661 (I183106,I1862,I182699,I182679,);
nand I_10662 (I183137,I182931,I182996);
nor I_10663 (I182673,I182784,I183137);
nor I_10664 (I183168,I182931,I182996);
nand I_10665 (I182682,I183168,I182979);
not I_10666 (I183226,I1869);
or I_10667 (I183243,I108757,I108766);
nand I_10668 (I183260,I108760,I108763);
not I_10669 (I183277,I183260);
nand I_10670 (I183294,I183277,I183243);
not I_10671 (I183311,I183294);
nand I_10672 (I183328,I108754,I108754);
and I_10673 (I183345,I183328,I108751);
DFFARX1 I_10674 (I183345,I1862,I183226,I183371,);
nor I_10675 (I183194,I183371,I183260);
nand I_10676 (I183393,I183311,I183371);
nor I_10677 (I183410,I183371,I183277);
not I_10678 (I183212,I183371);
nor I_10679 (I183441,I108769,I108754);
not I_10680 (I183458,I183441);
nand I_10681 (I183215,I183410,I183441);
not I_10682 (I183489,I108757);
nor I_10683 (I183506,I183371,I108757);
nand I_10684 (I183523,I108760,I108751);
nor I_10685 (I183197,I183523,I183260);
not I_10686 (I183554,I183523);
nor I_10687 (I183571,I183441,I183554);
nor I_10688 (I183218,I183571,I183294);
nand I_10689 (I183602,I183554,I183489);
nand I_10690 (I183203,I183311,I183602);
nand I_10691 (I183633,I183393,I183602);
DFFARX1 I_10692 (I183633,I1862,I183226,I183206,);
nand I_10693 (I183664,I183458,I183523);
nor I_10694 (I183200,I183311,I183664);
nor I_10695 (I183695,I183458,I183523);
nand I_10696 (I183209,I183695,I183506);
not I_10697 (I183753,I1869);
or I_10698 (I183770,I79276,I79273);
nand I_10699 (I183787,I79279,I79276);
not I_10700 (I183804,I183787);
nand I_10701 (I183821,I183804,I183770);
not I_10702 (I183838,I183821);
nand I_10703 (I183855,I79294,I79297);
and I_10704 (I183872,I183855,I79273);
DFFARX1 I_10705 (I183872,I1862,I183753,I183898,);
nor I_10706 (I183721,I183898,I183787);
nand I_10707 (I183920,I183838,I183898);
nor I_10708 (I183937,I183898,I183804);
not I_10709 (I183739,I183898);
nor I_10710 (I183968,I79291,I79297);
not I_10711 (I183985,I183968);
nand I_10712 (I183742,I183937,I183968);
not I_10713 (I184016,I79282);
nor I_10714 (I184033,I183898,I79282);
nand I_10715 (I184050,I79285,I79288);
nor I_10716 (I183724,I184050,I183787);
not I_10717 (I184081,I184050);
nor I_10718 (I184098,I183968,I184081);
nor I_10719 (I183745,I184098,I183821);
nand I_10720 (I184129,I184081,I184016);
nand I_10721 (I183730,I183838,I184129);
nand I_10722 (I184160,I183920,I184129);
DFFARX1 I_10723 (I184160,I1862,I183753,I183733,);
nand I_10724 (I184191,I183985,I184050);
nor I_10725 (I183727,I183838,I184191);
nor I_10726 (I184222,I183985,I184050);
nand I_10727 (I183736,I184222,I184033);
not I_10728 (I184280,I1869);
or I_10729 (I184297,I273413,I273416);
nand I_10730 (I184314,I273419,I273428);
not I_10731 (I184331,I184314);
nand I_10732 (I184348,I184331,I184297);
not I_10733 (I184365,I184348);
nand I_10734 (I184382,I273425,I273431);
and I_10735 (I184399,I184382,I273413);
DFFARX1 I_10736 (I184399,I1862,I184280,I184425,);
nor I_10737 (I184248,I184425,I184314);
nand I_10738 (I184447,I184365,I184425);
nor I_10739 (I184464,I184425,I184331);
not I_10740 (I184266,I184425);
nor I_10741 (I184495,I273416,I273431);
not I_10742 (I184512,I184495);
nand I_10743 (I184269,I184464,I184495);
not I_10744 (I184543,I273434);
nor I_10745 (I184560,I184425,I273434);
nand I_10746 (I184577,I273422,I273419);
nor I_10747 (I184251,I184577,I184314);
not I_10748 (I184608,I184577);
nor I_10749 (I184625,I184495,I184608);
nor I_10750 (I184272,I184625,I184348);
nand I_10751 (I184656,I184608,I184543);
nand I_10752 (I184257,I184365,I184656);
nand I_10753 (I184687,I184447,I184656);
DFFARX1 I_10754 (I184687,I1862,I184280,I184260,);
nand I_10755 (I184718,I184512,I184577);
nor I_10756 (I184254,I184365,I184718);
nor I_10757 (I184749,I184512,I184577);
nand I_10758 (I184263,I184749,I184560);
not I_10759 (I184807,I1869);
or I_10760 (I184824,I339459,I339447);
nand I_10761 (I184841,I339441,I339441);
not I_10762 (I184858,I184841);
nand I_10763 (I184875,I184858,I184824);
not I_10764 (I184892,I184875);
nand I_10765 (I184909,I339444,I339444);
and I_10766 (I184926,I184909,I339450);
DFFARX1 I_10767 (I184926,I1862,I184807,I184952,);
nor I_10768 (I184775,I184952,I184841);
nand I_10769 (I184974,I184892,I184952);
nor I_10770 (I184991,I184952,I184858);
not I_10771 (I184793,I184952);
nor I_10772 (I185022,I339456,I339444);
not I_10773 (I185039,I185022);
nand I_10774 (I184796,I184991,I185022);
not I_10775 (I185070,I339462);
nor I_10776 (I185087,I184952,I339462);
nand I_10777 (I185104,I339447,I339453);
nor I_10778 (I184778,I185104,I184841);
not I_10779 (I185135,I185104);
nor I_10780 (I185152,I185022,I185135);
nor I_10781 (I184799,I185152,I184875);
nand I_10782 (I185183,I185135,I185070);
nand I_10783 (I184784,I184892,I185183);
nand I_10784 (I185214,I184974,I185183);
DFFARX1 I_10785 (I185214,I1862,I184807,I184787,);
nand I_10786 (I185245,I185039,I185104);
nor I_10787 (I184781,I184892,I185245);
nor I_10788 (I185276,I185039,I185104);
nand I_10789 (I184790,I185276,I185087);
not I_10790 (I185334,I1869);
or I_10791 (I185351,I305204,I305192);
nand I_10792 (I185368,I305186,I305186);
not I_10793 (I185385,I185368);
nand I_10794 (I185402,I185385,I185351);
not I_10795 (I185419,I185402);
nand I_10796 (I185436,I305189,I305189);
and I_10797 (I185453,I185436,I305195);
DFFARX1 I_10798 (I185453,I1862,I185334,I185479,);
nor I_10799 (I185302,I185479,I185368);
nand I_10800 (I185501,I185419,I185479);
nor I_10801 (I185518,I185479,I185385);
not I_10802 (I185320,I185479);
nor I_10803 (I185549,I305201,I305189);
not I_10804 (I185566,I185549);
nand I_10805 (I185323,I185518,I185549);
not I_10806 (I185597,I305207);
nor I_10807 (I185614,I185479,I305207);
nand I_10808 (I185631,I305192,I305198);
nor I_10809 (I185305,I185631,I185368);
not I_10810 (I185662,I185631);
nor I_10811 (I185679,I185549,I185662);
nor I_10812 (I185326,I185679,I185402);
nand I_10813 (I185710,I185662,I185597);
nand I_10814 (I185311,I185419,I185710);
nand I_10815 (I185741,I185501,I185710);
DFFARX1 I_10816 (I185741,I1862,I185334,I185314,);
nand I_10817 (I185772,I185566,I185631);
nor I_10818 (I185308,I185419,I185772);
nor I_10819 (I185803,I185566,I185631);
nand I_10820 (I185317,I185803,I185614);
not I_10821 (I185861,I1869);
or I_10822 (I185878,I352107,I352095);
nand I_10823 (I185895,I352089,I352089);
not I_10824 (I185912,I185895);
nand I_10825 (I185929,I185912,I185878);
not I_10826 (I185946,I185929);
nand I_10827 (I185963,I352092,I352092);
and I_10828 (I185980,I185963,I352098);
DFFARX1 I_10829 (I185980,I1862,I185861,I186006,);
nor I_10830 (I185829,I186006,I185895);
nand I_10831 (I186028,I185946,I186006);
nor I_10832 (I186045,I186006,I185912);
not I_10833 (I185847,I186006);
nor I_10834 (I186076,I352104,I352092);
not I_10835 (I186093,I186076);
nand I_10836 (I185850,I186045,I186076);
not I_10837 (I186124,I352110);
nor I_10838 (I186141,I186006,I352110);
nand I_10839 (I186158,I352095,I352101);
nor I_10840 (I185832,I186158,I185895);
not I_10841 (I186189,I186158);
nor I_10842 (I186206,I186076,I186189);
nor I_10843 (I185853,I186206,I185929);
nand I_10844 (I186237,I186189,I186124);
nand I_10845 (I185838,I185946,I186237);
nand I_10846 (I186268,I186028,I186237);
DFFARX1 I_10847 (I186268,I1862,I185861,I185841,);
nand I_10848 (I186299,I186093,I186158);
nor I_10849 (I185835,I185946,I186299);
nor I_10850 (I186330,I186093,I186158);
nand I_10851 (I185844,I186330,I186141);
not I_10852 (I186388,I1869);
or I_10853 (I186405,I62446,I62443);
nand I_10854 (I186422,I62449,I62446);
not I_10855 (I186439,I186422);
nand I_10856 (I186456,I186439,I186405);
not I_10857 (I186473,I186456);
nand I_10858 (I186490,I62464,I62467);
and I_10859 (I186507,I186490,I62443);
DFFARX1 I_10860 (I186507,I1862,I186388,I186533,);
nor I_10861 (I186356,I186533,I186422);
nand I_10862 (I186555,I186473,I186533);
nor I_10863 (I186572,I186533,I186439);
not I_10864 (I186374,I186533);
nor I_10865 (I186603,I62461,I62467);
not I_10866 (I186620,I186603);
nand I_10867 (I186377,I186572,I186603);
not I_10868 (I186651,I62452);
nor I_10869 (I186668,I186533,I62452);
nand I_10870 (I186685,I62455,I62458);
nor I_10871 (I186359,I186685,I186422);
not I_10872 (I186716,I186685);
nor I_10873 (I186733,I186603,I186716);
nor I_10874 (I186380,I186733,I186456);
nand I_10875 (I186764,I186716,I186651);
nand I_10876 (I186365,I186473,I186764);
nand I_10877 (I186795,I186555,I186764);
DFFARX1 I_10878 (I186795,I1862,I186388,I186368,);
nand I_10879 (I186826,I186620,I186685);
nor I_10880 (I186362,I186473,I186826);
nor I_10881 (I186857,I186620,I186685);
nand I_10882 (I186371,I186857,I186668);
not I_10883 (I186915,I1869);
or I_10884 (I186932,I357904,I357892);
nand I_10885 (I186949,I357886,I357886);
not I_10886 (I186966,I186949);
nand I_10887 (I186983,I186966,I186932);
not I_10888 (I187000,I186983);
nand I_10889 (I187017,I357889,I357889);
and I_10890 (I187034,I187017,I357895);
DFFARX1 I_10891 (I187034,I1862,I186915,I187060,);
nor I_10892 (I186883,I187060,I186949);
nand I_10893 (I187082,I187000,I187060);
nor I_10894 (I187099,I187060,I186966);
not I_10895 (I186901,I187060);
nor I_10896 (I187130,I357901,I357889);
not I_10897 (I187147,I187130);
nand I_10898 (I186904,I187099,I187130);
not I_10899 (I187178,I357907);
nor I_10900 (I187195,I187060,I357907);
nand I_10901 (I187212,I357892,I357898);
nor I_10902 (I186886,I187212,I186949);
not I_10903 (I187243,I187212);
nor I_10904 (I187260,I187130,I187243);
nor I_10905 (I186907,I187260,I186983);
nand I_10906 (I187291,I187243,I187178);
nand I_10907 (I186892,I187000,I187291);
nand I_10908 (I187322,I187082,I187291);
DFFARX1 I_10909 (I187322,I1862,I186915,I186895,);
nand I_10910 (I187353,I187147,I187212);
nor I_10911 (I186889,I187000,I187353);
nor I_10912 (I187384,I187147,I187212);
nand I_10913 (I186898,I187384,I187195);
not I_10914 (I187442,I1869);
or I_10915 (I187459,I42556,I42553);
nand I_10916 (I187476,I42559,I42556);
not I_10917 (I187493,I187476);
nand I_10918 (I187510,I187493,I187459);
not I_10919 (I187527,I187510);
nand I_10920 (I187544,I42574,I42577);
and I_10921 (I187561,I187544,I42553);
DFFARX1 I_10922 (I187561,I1862,I187442,I187587,);
nor I_10923 (I187410,I187587,I187476);
nand I_10924 (I187609,I187527,I187587);
nor I_10925 (I187626,I187587,I187493);
not I_10926 (I187428,I187587);
nor I_10927 (I187657,I42571,I42577);
not I_10928 (I187674,I187657);
nand I_10929 (I187431,I187626,I187657);
not I_10930 (I187705,I42562);
nor I_10931 (I187722,I187587,I42562);
nand I_10932 (I187739,I42565,I42568);
nor I_10933 (I187413,I187739,I187476);
not I_10934 (I187770,I187739);
nor I_10935 (I187787,I187657,I187770);
nor I_10936 (I187434,I187787,I187510);
nand I_10937 (I187818,I187770,I187705);
nand I_10938 (I187419,I187527,I187818);
nand I_10939 (I187849,I187609,I187818);
DFFARX1 I_10940 (I187849,I1862,I187442,I187422,);
nand I_10941 (I187880,I187674,I187739);
nor I_10942 (I187416,I187527,I187880);
nor I_10943 (I187911,I187674,I187739);
nand I_10944 (I187425,I187911,I187722);
not I_10945 (I187969,I1869);
or I_10946 (I187986,I49186,I49183);
nand I_10947 (I188003,I49189,I49186);
not I_10948 (I188020,I188003);
nand I_10949 (I188037,I188020,I187986);
not I_10950 (I188054,I188037);
nand I_10951 (I188071,I49204,I49207);
and I_10952 (I188088,I188071,I49183);
DFFARX1 I_10953 (I188088,I1862,I187969,I188114,);
nor I_10954 (I187937,I188114,I188003);
nand I_10955 (I188136,I188054,I188114);
nor I_10956 (I188153,I188114,I188020);
not I_10957 (I187955,I188114);
nor I_10958 (I188184,I49201,I49207);
not I_10959 (I188201,I188184);
nand I_10960 (I187958,I188153,I188184);
not I_10961 (I188232,I49192);
nor I_10962 (I188249,I188114,I49192);
nand I_10963 (I188266,I49195,I49198);
nor I_10964 (I187940,I188266,I188003);
not I_10965 (I188297,I188266);
nor I_10966 (I188314,I188184,I188297);
nor I_10967 (I187961,I188314,I188037);
nand I_10968 (I188345,I188297,I188232);
nand I_10969 (I187946,I188054,I188345);
nand I_10970 (I188376,I188136,I188345);
DFFARX1 I_10971 (I188376,I1862,I187969,I187949,);
nand I_10972 (I188407,I188201,I188266);
nor I_10973 (I187943,I188054,I188407);
nor I_10974 (I188438,I188201,I188266);
nand I_10975 (I187952,I188438,I188249);
not I_10976 (I188496,I1869);
or I_10977 (I188513,I14506,I14503);
nand I_10978 (I188530,I14509,I14506);
not I_10979 (I188547,I188530);
nand I_10980 (I188564,I188547,I188513);
not I_10981 (I188581,I188564);
nand I_10982 (I188598,I14524,I14527);
and I_10983 (I188615,I188598,I14503);
DFFARX1 I_10984 (I188615,I1862,I188496,I188641,);
nor I_10985 (I188464,I188641,I188530);
nand I_10986 (I188663,I188581,I188641);
nor I_10987 (I188680,I188641,I188547);
not I_10988 (I188482,I188641);
nor I_10989 (I188711,I14521,I14527);
not I_10990 (I188728,I188711);
nand I_10991 (I188485,I188680,I188711);
not I_10992 (I188759,I14512);
nor I_10993 (I188776,I188641,I14512);
nand I_10994 (I188793,I14515,I14518);
nor I_10995 (I188467,I188793,I188530);
not I_10996 (I188824,I188793);
nor I_10997 (I188841,I188711,I188824);
nor I_10998 (I188488,I188841,I188564);
nand I_10999 (I188872,I188824,I188759);
nand I_11000 (I188473,I188581,I188872);
nand I_11001 (I188903,I188663,I188872);
DFFARX1 I_11002 (I188903,I1862,I188496,I188476,);
nand I_11003 (I188934,I188728,I188793);
nor I_11004 (I188470,I188581,I188934);
nor I_11005 (I188965,I188728,I188793);
nand I_11006 (I188479,I188965,I188776);
not I_11007 (I189023,I1869);
or I_11008 (I189040,I21646,I21643);
nand I_11009 (I189057,I21649,I21646);
not I_11010 (I189074,I189057);
nand I_11011 (I189091,I189074,I189040);
not I_11012 (I189108,I189091);
nand I_11013 (I189125,I21664,I21667);
and I_11014 (I189142,I189125,I21643);
DFFARX1 I_11015 (I189142,I1862,I189023,I189168,);
nor I_11016 (I188991,I189168,I189057);
nand I_11017 (I189190,I189108,I189168);
nor I_11018 (I189207,I189168,I189074);
not I_11019 (I189009,I189168);
nor I_11020 (I189238,I21661,I21667);
not I_11021 (I189255,I189238);
nand I_11022 (I189012,I189207,I189238);
not I_11023 (I189286,I21652);
nor I_11024 (I189303,I189168,I21652);
nand I_11025 (I189320,I21655,I21658);
nor I_11026 (I188994,I189320,I189057);
not I_11027 (I189351,I189320);
nor I_11028 (I189368,I189238,I189351);
nor I_11029 (I189015,I189368,I189091);
nand I_11030 (I189399,I189351,I189286);
nand I_11031 (I189000,I189108,I189399);
nand I_11032 (I189430,I189190,I189399);
DFFARX1 I_11033 (I189430,I1862,I189023,I189003,);
nand I_11034 (I189461,I189255,I189320);
nor I_11035 (I188997,I189108,I189461);
nor I_11036 (I189492,I189255,I189320);
nand I_11037 (I189006,I189492,I189303);
not I_11038 (I189550,I1869);
or I_11039 (I189567,I318379,I318367);
nand I_11040 (I189584,I318361,I318361);
not I_11041 (I189601,I189584);
nand I_11042 (I189618,I189601,I189567);
not I_11043 (I189635,I189618);
nand I_11044 (I189652,I318364,I318364);
and I_11045 (I189669,I189652,I318370);
DFFARX1 I_11046 (I189669,I1862,I189550,I189695,);
nor I_11047 (I189518,I189695,I189584);
nand I_11048 (I189717,I189635,I189695);
nor I_11049 (I189734,I189695,I189601);
not I_11050 (I189536,I189695);
nor I_11051 (I189765,I318376,I318364);
not I_11052 (I189782,I189765);
nand I_11053 (I189539,I189734,I189765);
not I_11054 (I189813,I318382);
nor I_11055 (I189830,I189695,I318382);
nand I_11056 (I189847,I318367,I318373);
nor I_11057 (I189521,I189847,I189584);
not I_11058 (I189878,I189847);
nor I_11059 (I189895,I189765,I189878);
nor I_11060 (I189542,I189895,I189618);
nand I_11061 (I189926,I189878,I189813);
nand I_11062 (I189527,I189635,I189926);
nand I_11063 (I189957,I189717,I189926);
DFFARX1 I_11064 (I189957,I1862,I189550,I189530,);
nand I_11065 (I189988,I189782,I189847);
nor I_11066 (I189524,I189635,I189988);
nor I_11067 (I190019,I189782,I189847);
nand I_11068 (I189533,I190019,I189830);
not I_11069 (I190077,I1869);
or I_11070 (I190094,I400834,I400831);
nand I_11071 (I190111,I400843,I400846);
not I_11072 (I190128,I190111);
nand I_11073 (I190145,I190128,I190094);
not I_11074 (I190162,I190145);
nand I_11075 (I190179,I400837,I400828);
and I_11076 (I190196,I190179,I400828);
DFFARX1 I_11077 (I190196,I1862,I190077,I190222,);
nor I_11078 (I190045,I190222,I190111);
nand I_11079 (I190244,I190162,I190222);
nor I_11080 (I190261,I190222,I190128);
not I_11081 (I190063,I190222);
nor I_11082 (I190292,I400831,I400828);
not I_11083 (I190309,I190292);
nand I_11084 (I190066,I190261,I190292);
not I_11085 (I190340,I400834);
nor I_11086 (I190357,I190222,I400834);
nand I_11087 (I190374,I400837,I400840);
nor I_11088 (I190048,I190374,I190111);
not I_11089 (I190405,I190374);
nor I_11090 (I190422,I190292,I190405);
nor I_11091 (I190069,I190422,I190145);
nand I_11092 (I190453,I190405,I190340);
nand I_11093 (I190054,I190162,I190453);
nand I_11094 (I190484,I190244,I190453);
DFFARX1 I_11095 (I190484,I1862,I190077,I190057,);
nand I_11096 (I190515,I190309,I190374);
nor I_11097 (I190051,I190162,I190515);
nor I_11098 (I190546,I190309,I190374);
nand I_11099 (I190060,I190546,I190357);
not I_11100 (I190604,I1869);
or I_11101 (I190621,I68056,I68053);
nand I_11102 (I190638,I68059,I68056);
not I_11103 (I190655,I190638);
nand I_11104 (I190672,I190655,I190621);
not I_11105 (I190689,I190672);
nand I_11106 (I190706,I68074,I68077);
and I_11107 (I190723,I190706,I68053);
DFFARX1 I_11108 (I190723,I1862,I190604,I190749,);
nor I_11109 (I190572,I190749,I190638);
nand I_11110 (I190771,I190689,I190749);
nor I_11111 (I190788,I190749,I190655);
not I_11112 (I190590,I190749);
nor I_11113 (I190819,I68071,I68077);
not I_11114 (I190836,I190819);
nand I_11115 (I190593,I190788,I190819);
not I_11116 (I190867,I68062);
nor I_11117 (I190884,I190749,I68062);
nand I_11118 (I190901,I68065,I68068);
nor I_11119 (I190575,I190901,I190638);
not I_11120 (I190932,I190901);
nor I_11121 (I190949,I190819,I190932);
nor I_11122 (I190596,I190949,I190672);
nand I_11123 (I190980,I190932,I190867);
nand I_11124 (I190581,I190689,I190980);
nand I_11125 (I191011,I190771,I190980);
DFFARX1 I_11126 (I191011,I1862,I190604,I190584,);
nand I_11127 (I191042,I190836,I190901);
nor I_11128 (I190578,I190689,I191042);
nor I_11129 (I191073,I190836,I190901);
nand I_11130 (I190587,I191073,I190884);
not I_11131 (I191131,I1869);
or I_11132 (I191148,I263893,I263896);
nand I_11133 (I191165,I263899,I263908);
not I_11134 (I191182,I191165);
nand I_11135 (I191199,I191182,I191148);
not I_11136 (I191216,I191199);
nand I_11137 (I191233,I263905,I263911);
and I_11138 (I191250,I191233,I263893);
DFFARX1 I_11139 (I191250,I1862,I191131,I191276,);
nor I_11140 (I191099,I191276,I191165);
nand I_11141 (I191298,I191216,I191276);
nor I_11142 (I191315,I191276,I191182);
not I_11143 (I191117,I191276);
nor I_11144 (I191346,I263896,I263911);
not I_11145 (I191363,I191346);
nand I_11146 (I191120,I191315,I191346);
not I_11147 (I191394,I263914);
nor I_11148 (I191411,I191276,I263914);
nand I_11149 (I191428,I263902,I263899);
nor I_11150 (I191102,I191428,I191165);
not I_11151 (I191459,I191428);
nor I_11152 (I191476,I191346,I191459);
nor I_11153 (I191123,I191476,I191199);
nand I_11154 (I191507,I191459,I191394);
nand I_11155 (I191108,I191216,I191507);
nand I_11156 (I191538,I191298,I191507);
DFFARX1 I_11157 (I191538,I1862,I191131,I191111,);
nand I_11158 (I191569,I191363,I191428);
nor I_11159 (I191105,I191216,I191569);
nor I_11160 (I191600,I191363,I191428);
nand I_11161 (I191114,I191600,I191411);
not I_11162 (I191658,I1869);
or I_11163 (I191675,I204393,I204396);
nand I_11164 (I191692,I204399,I204408);
not I_11165 (I191709,I191692);
nand I_11166 (I191726,I191709,I191675);
not I_11167 (I191743,I191726);
nand I_11168 (I191760,I204405,I204411);
and I_11169 (I191777,I191760,I204393);
DFFARX1 I_11170 (I191777,I1862,I191658,I191803,);
nor I_11171 (I191626,I191803,I191692);
nand I_11172 (I191825,I191743,I191803);
nor I_11173 (I191842,I191803,I191709);
not I_11174 (I191644,I191803);
nor I_11175 (I191873,I204396,I204411);
not I_11176 (I191890,I191873);
nand I_11177 (I191647,I191842,I191873);
not I_11178 (I191921,I204414);
nor I_11179 (I191938,I191803,I204414);
nand I_11180 (I191955,I204402,I204399);
nor I_11181 (I191629,I191955,I191692);
not I_11182 (I191986,I191955);
nor I_11183 (I192003,I191873,I191986);
nor I_11184 (I191650,I192003,I191726);
nand I_11185 (I192034,I191986,I191921);
nand I_11186 (I191635,I191743,I192034);
nand I_11187 (I192065,I191825,I192034);
DFFARX1 I_11188 (I192065,I1862,I191658,I191638,);
nand I_11189 (I192096,I191890,I191955);
nor I_11190 (I191632,I191743,I192096);
nor I_11191 (I192127,I191890,I191955);
nand I_11192 (I191641,I192127,I191938);
not I_11193 (I192185,I1869);
or I_11194 (I192202,I316271,I316259);
nand I_11195 (I192219,I316253,I316253);
not I_11196 (I192236,I192219);
nand I_11197 (I192253,I192236,I192202);
not I_11198 (I192270,I192253);
nand I_11199 (I192287,I316256,I316256);
and I_11200 (I192304,I192287,I316262);
DFFARX1 I_11201 (I192304,I1862,I192185,I192330,);
nor I_11202 (I192153,I192330,I192219);
nand I_11203 (I192352,I192270,I192330);
nor I_11204 (I192369,I192330,I192236);
not I_11205 (I192171,I192330);
nor I_11206 (I192400,I316268,I316256);
not I_11207 (I192417,I192400);
nand I_11208 (I192174,I192369,I192400);
not I_11209 (I192448,I316274);
nor I_11210 (I192465,I192330,I316274);
nand I_11211 (I192482,I316259,I316265);
nor I_11212 (I192156,I192482,I192219);
not I_11213 (I192513,I192482);
nor I_11214 (I192530,I192400,I192513);
nor I_11215 (I192177,I192530,I192253);
nand I_11216 (I192561,I192513,I192448);
nand I_11217 (I192162,I192270,I192561);
nand I_11218 (I192592,I192352,I192561);
DFFARX1 I_11219 (I192592,I1862,I192185,I192165,);
nand I_11220 (I192623,I192417,I192482);
nor I_11221 (I192159,I192270,I192623);
nor I_11222 (I192654,I192417,I192482);
nand I_11223 (I192168,I192654,I192465);
not I_11224 (I192712,I1869);
or I_11225 (I192729,I1647,I1815);
nand I_11226 (I192746,I647,I1743);
not I_11227 (I192763,I192746);
nand I_11228 (I192780,I192763,I192729);
not I_11229 (I192797,I192780);
nand I_11230 (I192814,I751,I839);
and I_11231 (I192831,I192814,I1471);
DFFARX1 I_11232 (I192831,I1862,I192712,I192857,);
nor I_11233 (I192680,I192857,I192746);
nand I_11234 (I192879,I192797,I192857);
nor I_11235 (I192896,I192857,I192763);
not I_11236 (I192698,I192857);
nor I_11237 (I192927,I1351,I839);
not I_11238 (I192944,I192927);
nand I_11239 (I192701,I192896,I192927);
not I_11240 (I192975,I1495);
nor I_11241 (I192992,I192857,I1495);
nand I_11242 (I193009,I1487,I1783);
nor I_11243 (I192683,I193009,I192746);
not I_11244 (I193040,I193009);
nor I_11245 (I193057,I192927,I193040);
nor I_11246 (I192704,I193057,I192780);
nand I_11247 (I193088,I193040,I192975);
nand I_11248 (I192689,I192797,I193088);
nand I_11249 (I193119,I192879,I193088);
DFFARX1 I_11250 (I193119,I1862,I192712,I192692,);
nand I_11251 (I193150,I192944,I193009);
nor I_11252 (I192686,I192797,I193150);
nor I_11253 (I193181,I192944,I193009);
nand I_11254 (I192695,I193181,I192992);
not I_11255 (I193239,I1869);
or I_11256 (I193256,I203917,I203920);
nand I_11257 (I193273,I203923,I203932);
not I_11258 (I193290,I193273);
nand I_11259 (I193307,I193290,I193256);
not I_11260 (I193324,I193307);
nand I_11261 (I193341,I203929,I203935);
and I_11262 (I193358,I193341,I203917);
DFFARX1 I_11263 (I193358,I1862,I193239,I193384,);
nor I_11264 (I193207,I193384,I193273);
nand I_11265 (I193406,I193324,I193384);
nor I_11266 (I193423,I193384,I193290);
not I_11267 (I193225,I193384);
nor I_11268 (I193454,I203920,I203935);
not I_11269 (I193471,I193454);
nand I_11270 (I193228,I193423,I193454);
not I_11271 (I193502,I203938);
nor I_11272 (I193519,I193384,I203938);
nand I_11273 (I193536,I203926,I203923);
nor I_11274 (I193210,I193536,I193273);
not I_11275 (I193567,I193536);
nor I_11276 (I193584,I193454,I193567);
nor I_11277 (I193231,I193584,I193307);
nand I_11278 (I193615,I193567,I193502);
nand I_11279 (I193216,I193324,I193615);
nand I_11280 (I193646,I193406,I193615);
DFFARX1 I_11281 (I193646,I1862,I193239,I193219,);
nand I_11282 (I193677,I193471,I193536);
nor I_11283 (I193213,I193324,I193677);
nor I_11284 (I193708,I193471,I193536);
nand I_11285 (I193222,I193708,I193519);
not I_11286 (I193766,I1869);
or I_11287 (I193783,I275317,I275320);
nand I_11288 (I193800,I275323,I275332);
not I_11289 (I193817,I193800);
nand I_11290 (I193834,I193817,I193783);
not I_11291 (I193851,I193834);
nand I_11292 (I193868,I275329,I275335);
and I_11293 (I193885,I193868,I275317);
DFFARX1 I_11294 (I193885,I1862,I193766,I193911,);
nor I_11295 (I193734,I193911,I193800);
nand I_11296 (I193933,I193851,I193911);
nor I_11297 (I193950,I193911,I193817);
not I_11298 (I193752,I193911);
nor I_11299 (I193981,I275320,I275335);
not I_11300 (I193998,I193981);
nand I_11301 (I193755,I193950,I193981);
not I_11302 (I194029,I275338);
nor I_11303 (I194046,I193911,I275338);
nand I_11304 (I194063,I275326,I275323);
nor I_11305 (I193737,I194063,I193800);
not I_11306 (I194094,I194063);
nor I_11307 (I194111,I193981,I194094);
nor I_11308 (I193758,I194111,I193834);
nand I_11309 (I194142,I194094,I194029);
nand I_11310 (I193743,I193851,I194142);
nand I_11311 (I194173,I193933,I194142);
DFFARX1 I_11312 (I194173,I1862,I193766,I193746,);
nand I_11313 (I194204,I193998,I194063);
nor I_11314 (I193740,I193851,I194204);
nor I_11315 (I194235,I193998,I194063);
nand I_11316 (I193749,I194235,I194046);
not I_11317 (I194293,I1869);
or I_11318 (I194310,I232001,I232004);
nand I_11319 (I194327,I232007,I232016);
not I_11320 (I194344,I194327);
nand I_11321 (I194361,I194344,I194310);
not I_11322 (I194378,I194361);
nand I_11323 (I194395,I232013,I232019);
and I_11324 (I194412,I194395,I232001);
DFFARX1 I_11325 (I194412,I1862,I194293,I194438,);
nor I_11326 (I194261,I194438,I194327);
nand I_11327 (I194460,I194378,I194438);
nor I_11328 (I194477,I194438,I194344);
not I_11329 (I194279,I194438);
nor I_11330 (I194508,I232004,I232019);
not I_11331 (I194525,I194508);
nand I_11332 (I194282,I194477,I194508);
not I_11333 (I194556,I232022);
nor I_11334 (I194573,I194438,I232022);
nand I_11335 (I194590,I232010,I232007);
nor I_11336 (I194264,I194590,I194327);
not I_11337 (I194621,I194590);
nor I_11338 (I194638,I194508,I194621);
nor I_11339 (I194285,I194638,I194361);
nand I_11340 (I194669,I194621,I194556);
nand I_11341 (I194270,I194378,I194669);
nand I_11342 (I194700,I194460,I194669);
DFFARX1 I_11343 (I194700,I1862,I194293,I194273,);
nand I_11344 (I194731,I194525,I194590);
nor I_11345 (I194267,I194378,I194731);
nor I_11346 (I194762,I194525,I194590);
nand I_11347 (I194276,I194762,I194573);
not I_11348 (I194820,I1869);
or I_11349 (I194837,I85906,I85903);
nand I_11350 (I194854,I85909,I85906);
not I_11351 (I194871,I194854);
nand I_11352 (I194888,I194871,I194837);
not I_11353 (I194905,I194888);
nand I_11354 (I194922,I85924,I85927);
and I_11355 (I194939,I194922,I85903);
DFFARX1 I_11356 (I194939,I1862,I194820,I194965,);
nor I_11357 (I194788,I194965,I194854);
nand I_11358 (I194987,I194905,I194965);
nor I_11359 (I195004,I194965,I194871);
not I_11360 (I194806,I194965);
nor I_11361 (I195035,I85921,I85927);
not I_11362 (I195052,I195035);
nand I_11363 (I194809,I195004,I195035);
not I_11364 (I195083,I85912);
nor I_11365 (I195100,I194965,I85912);
nand I_11366 (I195117,I85915,I85918);
nor I_11367 (I194791,I195117,I194854);
not I_11368 (I195148,I195117);
nor I_11369 (I195165,I195035,I195148);
nor I_11370 (I194812,I195165,I194888);
nand I_11371 (I195196,I195148,I195083);
nand I_11372 (I194797,I194905,I195196);
nand I_11373 (I195227,I194987,I195196);
DFFARX1 I_11374 (I195227,I1862,I194820,I194800,);
nand I_11375 (I195258,I195052,I195117);
nor I_11376 (I194794,I194905,I195258);
nor I_11377 (I195289,I195052,I195117);
nand I_11378 (I194803,I195289,I195100);
not I_11379 (I195347,I1869);
or I_11380 (I195364,I71116,I71113);
nand I_11381 (I195381,I71119,I71116);
not I_11382 (I195398,I195381);
nand I_11383 (I195415,I195398,I195364);
not I_11384 (I195432,I195415);
nand I_11385 (I195449,I71134,I71137);
and I_11386 (I195466,I195449,I71113);
DFFARX1 I_11387 (I195466,I1862,I195347,I195492,);
nor I_11388 (I195315,I195492,I195381);
nand I_11389 (I195514,I195432,I195492);
nor I_11390 (I195531,I195492,I195398);
not I_11391 (I195333,I195492);
nor I_11392 (I195562,I71131,I71137);
not I_11393 (I195579,I195562);
nand I_11394 (I195336,I195531,I195562);
not I_11395 (I195610,I71122);
nor I_11396 (I195627,I195492,I71122);
nand I_11397 (I195644,I71125,I71128);
nor I_11398 (I195318,I195644,I195381);
not I_11399 (I195675,I195644);
nor I_11400 (I195692,I195562,I195675);
nor I_11401 (I195339,I195692,I195415);
nand I_11402 (I195723,I195675,I195610);
nand I_11403 (I195324,I195432,I195723);
nand I_11404 (I195754,I195514,I195723);
DFFARX1 I_11405 (I195754,I1862,I195347,I195327,);
nand I_11406 (I195785,I195579,I195644);
nor I_11407 (I195321,I195432,I195785);
nor I_11408 (I195816,I195579,I195644);
nand I_11409 (I195330,I195816,I195627);
not I_11410 (I195874,I1869);
or I_11411 (I195891,I401718,I401715);
nand I_11412 (I195908,I401727,I401730);
not I_11413 (I195925,I195908);
nand I_11414 (I195942,I195925,I195891);
not I_11415 (I195959,I195942);
nand I_11416 (I195976,I401721,I401712);
and I_11417 (I195993,I195976,I401712);
DFFARX1 I_11418 (I195993,I1862,I195874,I196019,);
nor I_11419 (I195842,I196019,I195908);
nand I_11420 (I196041,I195959,I196019);
nor I_11421 (I196058,I196019,I195925);
not I_11422 (I195860,I196019);
nor I_11423 (I196089,I401715,I401712);
not I_11424 (I196106,I196089);
nand I_11425 (I195863,I196058,I196089);
not I_11426 (I196137,I401718);
nor I_11427 (I196154,I196019,I401718);
nand I_11428 (I196171,I401721,I401724);
nor I_11429 (I195845,I196171,I195908);
not I_11430 (I196202,I196171);
nor I_11431 (I196219,I196089,I196202);
nor I_11432 (I195866,I196219,I195942);
nand I_11433 (I196250,I196202,I196137);
nand I_11434 (I195851,I195959,I196250);
nand I_11435 (I196281,I196041,I196250);
DFFARX1 I_11436 (I196281,I1862,I195874,I195854,);
nand I_11437 (I196312,I196106,I196171);
nor I_11438 (I195848,I195959,I196312);
nor I_11439 (I196343,I196106,I196171);
nand I_11440 (I195857,I196343,I196154);
not I_11441 (I196401,I1869);
or I_11442 (I196418,I348418,I348406);
nand I_11443 (I196435,I348400,I348400);
not I_11444 (I196452,I196435);
nand I_11445 (I196469,I196452,I196418);
not I_11446 (I196486,I196469);
nand I_11447 (I196503,I348403,I348403);
and I_11448 (I196520,I196503,I348409);
DFFARX1 I_11449 (I196520,I1862,I196401,I196546,);
nor I_11450 (I196369,I196546,I196435);
nand I_11451 (I196568,I196486,I196546);
nor I_11452 (I196585,I196546,I196452);
not I_11453 (I196387,I196546);
nor I_11454 (I196616,I348415,I348403);
not I_11455 (I196633,I196616);
nand I_11456 (I196390,I196585,I196616);
not I_11457 (I196664,I348421);
nor I_11458 (I196681,I196546,I348421);
nand I_11459 (I196698,I348406,I348412);
nor I_11460 (I196372,I196698,I196435);
not I_11461 (I196729,I196698);
nor I_11462 (I196746,I196616,I196729);
nor I_11463 (I196393,I196746,I196469);
nand I_11464 (I196777,I196729,I196664);
nand I_11465 (I196378,I196486,I196777);
nand I_11466 (I196808,I196568,I196777);
DFFARX1 I_11467 (I196808,I1862,I196401,I196381,);
nand I_11468 (I196839,I196633,I196698);
nor I_11469 (I196375,I196486,I196839);
nor I_11470 (I196870,I196633,I196698);
nand I_11471 (I196384,I196870,I196681);
not I_11472 (I196928,I1869);
or I_11473 (I196945,I98146,I98143);
nand I_11474 (I196962,I98149,I98146);
not I_11475 (I196979,I196962);
nand I_11476 (I196996,I196979,I196945);
not I_11477 (I197013,I196996);
nand I_11478 (I197030,I98164,I98167);
and I_11479 (I197047,I197030,I98143);
DFFARX1 I_11480 (I197047,I1862,I196928,I197073,);
nor I_11481 (I196896,I197073,I196962);
nand I_11482 (I197095,I197013,I197073);
nor I_11483 (I197112,I197073,I196979);
not I_11484 (I196914,I197073);
nor I_11485 (I197143,I98161,I98167);
not I_11486 (I197160,I197143);
nand I_11487 (I196917,I197112,I197143);
not I_11488 (I197191,I98152);
nor I_11489 (I197208,I197073,I98152);
nand I_11490 (I197225,I98155,I98158);
nor I_11491 (I196899,I197225,I196962);
not I_11492 (I197256,I197225);
nor I_11493 (I197273,I197143,I197256);
nor I_11494 (I196920,I197273,I196996);
nand I_11495 (I197304,I197256,I197191);
nand I_11496 (I196905,I197013,I197304);
nand I_11497 (I197335,I197095,I197304);
DFFARX1 I_11498 (I197335,I1862,I196928,I196908,);
nand I_11499 (I197366,I197160,I197225);
nor I_11500 (I196902,I197013,I197366);
nor I_11501 (I197397,I197160,I197225);
nand I_11502 (I196911,I197397,I197208);
not I_11503 (I197455,I1869);
or I_11504 (I197472,I286265,I286268);
nand I_11505 (I197489,I286271,I286280);
not I_11506 (I197506,I197489);
nand I_11507 (I197523,I197506,I197472);
not I_11508 (I197540,I197523);
nand I_11509 (I197557,I286277,I286283);
and I_11510 (I197574,I197557,I286265);
DFFARX1 I_11511 (I197574,I1862,I197455,I197600,);
nor I_11512 (I197423,I197600,I197489);
nand I_11513 (I197622,I197540,I197600);
nor I_11514 (I197639,I197600,I197506);
not I_11515 (I197441,I197600);
nor I_11516 (I197670,I286268,I286283);
not I_11517 (I197687,I197670);
nand I_11518 (I197444,I197639,I197670);
not I_11519 (I197718,I286286);
nor I_11520 (I197735,I197600,I286286);
nand I_11521 (I197752,I286274,I286271);
nor I_11522 (I197426,I197752,I197489);
not I_11523 (I197783,I197752);
nor I_11524 (I197800,I197670,I197783);
nor I_11525 (I197447,I197800,I197523);
nand I_11526 (I197831,I197783,I197718);
nand I_11527 (I197432,I197540,I197831);
nand I_11528 (I197862,I197622,I197831);
DFFARX1 I_11529 (I197862,I1862,I197455,I197435,);
nand I_11530 (I197893,I197687,I197752);
nor I_11531 (I197429,I197540,I197893);
nor I_11532 (I197924,I197687,I197752);
nand I_11533 (I197438,I197924,I197735);
not I_11534 (I197982,I1869);
or I_11535 (I197999,I354215,I354203);
nand I_11536 (I198016,I354197,I354197);
not I_11537 (I198033,I198016);
nand I_11538 (I198050,I198033,I197999);
not I_11539 (I198067,I198050);
nand I_11540 (I198084,I354200,I354200);
and I_11541 (I198101,I198084,I354206);
DFFARX1 I_11542 (I198101,I1862,I197982,I198127,);
nor I_11543 (I197950,I198127,I198016);
nand I_11544 (I198149,I198067,I198127);
nor I_11545 (I198166,I198127,I198033);
not I_11546 (I197968,I198127);
nor I_11547 (I198197,I354212,I354200);
not I_11548 (I198214,I198197);
nand I_11549 (I197971,I198166,I198197);
not I_11550 (I198245,I354218);
nor I_11551 (I198262,I198127,I354218);
nand I_11552 (I198279,I354203,I354209);
nor I_11553 (I197953,I198279,I198016);
not I_11554 (I198310,I198279);
nor I_11555 (I198327,I198197,I198310);
nor I_11556 (I197974,I198327,I198050);
nand I_11557 (I198358,I198310,I198245);
nand I_11558 (I197959,I198067,I198358);
nand I_11559 (I198389,I198149,I198358);
DFFARX1 I_11560 (I198389,I1862,I197982,I197962,);
nand I_11561 (I198420,I198214,I198279);
nor I_11562 (I197956,I198067,I198420);
nor I_11563 (I198451,I198214,I198279);
nand I_11564 (I197965,I198451,I198262);
not I_11565 (I198509,I1869);
or I_11566 (I198526,I329973,I329961);
nand I_11567 (I198543,I329955,I329955);
not I_11568 (I198560,I198543);
nand I_11569 (I198577,I198560,I198526);
not I_11570 (I198594,I198577);
nand I_11571 (I198611,I329958,I329958);
and I_11572 (I198628,I198611,I329964);
DFFARX1 I_11573 (I198628,I1862,I198509,I198654,);
nor I_11574 (I198477,I198654,I198543);
nand I_11575 (I198676,I198594,I198654);
nor I_11576 (I198693,I198654,I198560);
not I_11577 (I198495,I198654);
nor I_11578 (I198724,I329970,I329958);
not I_11579 (I198741,I198724);
nand I_11580 (I198498,I198693,I198724);
not I_11581 (I198772,I329976);
nor I_11582 (I198789,I198654,I329976);
nand I_11583 (I198806,I329961,I329967);
nor I_11584 (I198480,I198806,I198543);
not I_11585 (I198837,I198806);
nor I_11586 (I198854,I198724,I198837);
nor I_11587 (I198501,I198854,I198577);
nand I_11588 (I198885,I198837,I198772);
nand I_11589 (I198486,I198594,I198885);
nand I_11590 (I198916,I198676,I198885);
DFFARX1 I_11591 (I198916,I1862,I198509,I198489,);
nand I_11592 (I198947,I198741,I198806);
nor I_11593 (I198483,I198594,I198947);
nor I_11594 (I198978,I198741,I198806);
nand I_11595 (I198492,I198978,I198789);
not I_11596 (I199036,I1869);
or I_11597 (I199053,I364590,I364587);
nand I_11598 (I199070,I364599,I364602);
not I_11599 (I199087,I199070);
nand I_11600 (I199104,I199087,I199053);
not I_11601 (I199121,I199104);
nand I_11602 (I199138,I364593,I364584);
and I_11603 (I199155,I199138,I364584);
DFFARX1 I_11604 (I199155,I1862,I199036,I199181,);
nor I_11605 (I199004,I199181,I199070);
nand I_11606 (I199203,I199121,I199181);
nor I_11607 (I199220,I199181,I199087);
not I_11608 (I199022,I199181);
nor I_11609 (I199251,I364587,I364584);
not I_11610 (I199268,I199251);
nand I_11611 (I199025,I199220,I199251);
not I_11612 (I199299,I364590);
nor I_11613 (I199316,I199181,I364590);
nand I_11614 (I199333,I364593,I364596);
nor I_11615 (I199007,I199333,I199070);
not I_11616 (I199364,I199333);
nor I_11617 (I199381,I199251,I199364);
nor I_11618 (I199028,I199381,I199104);
nand I_11619 (I199412,I199364,I199299);
nand I_11620 (I199013,I199121,I199412);
nand I_11621 (I199443,I199203,I199412);
DFFARX1 I_11622 (I199443,I1862,I199036,I199016,);
nand I_11623 (I199474,I199268,I199333);
nor I_11624 (I199010,I199121,I199474);
nor I_11625 (I199505,I199268,I199333);
nand I_11626 (I199019,I199505,I199316);
not I_11627 (I199563,I1869);
or I_11628 (I199580,I396856,I396853);
nand I_11629 (I199597,I396865,I396868);
not I_11630 (I199614,I199597);
nand I_11631 (I199631,I199614,I199580);
not I_11632 (I199648,I199631);
nand I_11633 (I199665,I396859,I396850);
and I_11634 (I199682,I199665,I396850);
DFFARX1 I_11635 (I199682,I1862,I199563,I199708,);
nor I_11636 (I199531,I199708,I199597);
nand I_11637 (I199730,I199648,I199708);
nor I_11638 (I199747,I199708,I199614);
not I_11639 (I199549,I199708);
nor I_11640 (I199778,I396853,I396850);
not I_11641 (I199795,I199778);
nand I_11642 (I199552,I199747,I199778);
not I_11643 (I199826,I396856);
nor I_11644 (I199843,I199708,I396856);
nand I_11645 (I199860,I396859,I396862);
nor I_11646 (I199534,I199860,I199597);
not I_11647 (I199891,I199860);
nor I_11648 (I199908,I199778,I199891);
nor I_11649 (I199555,I199908,I199631);
nand I_11650 (I199939,I199891,I199826);
nand I_11651 (I199540,I199648,I199939);
nand I_11652 (I199970,I199730,I199939);
DFFARX1 I_11653 (I199970,I1862,I199563,I199543,);
nand I_11654 (I200001,I199795,I199860);
nor I_11655 (I199537,I199648,I200001);
nor I_11656 (I200032,I199795,I199860);
nand I_11657 (I199546,I200032,I199843);
not I_11658 (I200090,I1869);
or I_11659 (I200107,I364148,I364145);
nand I_11660 (I200124,I364157,I364160);
not I_11661 (I200141,I200124);
nand I_11662 (I200158,I200141,I200107);
not I_11663 (I200175,I200158);
nand I_11664 (I200192,I364151,I364142);
and I_11665 (I200209,I200192,I364142);
DFFARX1 I_11666 (I200209,I1862,I200090,I200235,);
nor I_11667 (I200058,I200235,I200124);
nand I_11668 (I200257,I200175,I200235);
nor I_11669 (I200274,I200235,I200141);
not I_11670 (I200076,I200235);
nor I_11671 (I200305,I364145,I364142);
not I_11672 (I200322,I200305);
nand I_11673 (I200079,I200274,I200305);
not I_11674 (I200353,I364148);
nor I_11675 (I200370,I200235,I364148);
nand I_11676 (I200387,I364151,I364154);
nor I_11677 (I200061,I200387,I200124);
not I_11678 (I200418,I200387);
nor I_11679 (I200435,I200305,I200418);
nor I_11680 (I200082,I200435,I200158);
nand I_11681 (I200466,I200418,I200353);
nand I_11682 (I200067,I200175,I200466);
nand I_11683 (I200497,I200257,I200466);
DFFARX1 I_11684 (I200497,I1862,I200090,I200070,);
nand I_11685 (I200528,I200322,I200387);
nor I_11686 (I200064,I200175,I200528);
nor I_11687 (I200559,I200322,I200387);
nand I_11688 (I200073,I200559,I200370);
not I_11689 (I200614,I1869);
or I_11690 (I200631,I123667,I123652);
nor I_11691 (I200648,I200631,I123646);
nor I_11692 (I200665,I123643,I123664);
or I_11693 (I200682,I200665,I123661);
nor I_11694 (I200699,I123649,I123646);
nand I_11695 (I200716,I200699,I200682);
not I_11696 (I200733,I200716);
nand I_11697 (I200750,I200648,I200733);
nor I_11698 (I200767,I200648,I200733);
nand I_11699 (I200784,I123655,I123658);
nor I_11700 (I200801,I200784,I123643);
nor I_11701 (I200818,I200784,I200801);
not I_11702 (I200835,I200801);
nor I_11703 (I200606,I200835,I200750);
or I_11704 (I200591,I200648,I200835);
nor I_11705 (I200880,I200648,I200801);
nor I_11706 (I200585,I200784,I200880);
nor I_11707 (I200911,I200818,I200880);
nor I_11708 (I200588,I200733,I200911);
nand I_11709 (I200942,I200648,I200801);
nand I_11710 (I200959,I200716,I200942);
DFFARX1 I_11711 (I200959,I1862,I200614,I200594,);
not I_11712 (I200990,I200784);
nor I_11713 (I200603,I200990,I200835);
nand I_11714 (I200600,I200767,I200990);
nor I_11715 (I201035,I200733,I200784);
nand I_11716 (I200597,I201035,I200648);
not I_11717 (I201090,I1869);
or I_11718 (I201107,I103858,I103855);
nor I_11719 (I201124,I201107,I103855);
nor I_11720 (I201141,I103864,I103861);
or I_11721 (I201158,I201141,I103870);
nor I_11722 (I201175,I103873,I103858);
nand I_11723 (I201192,I201175,I201158);
not I_11724 (I201209,I201192);
nand I_11725 (I201226,I201124,I201209);
nor I_11726 (I201243,I201124,I201209);
nand I_11727 (I201260,I103861,I103867);
nor I_11728 (I201277,I201260,I103864);
nor I_11729 (I201294,I201260,I201277);
not I_11730 (I201311,I201277);
nor I_11731 (I201082,I201311,I201226);
or I_11732 (I201067,I201124,I201311);
nor I_11733 (I201356,I201124,I201277);
nor I_11734 (I201061,I201260,I201356);
nor I_11735 (I201387,I201294,I201356);
nor I_11736 (I201064,I201209,I201387);
nand I_11737 (I201418,I201124,I201277);
nand I_11738 (I201435,I201192,I201418);
DFFARX1 I_11739 (I201435,I1862,I201090,I201070,);
not I_11740 (I201466,I201260);
nor I_11741 (I201079,I201466,I201311);
nand I_11742 (I201076,I201243,I201466);
nor I_11743 (I201511,I201209,I201260);
nand I_11744 (I201073,I201511,I201124);
not I_11745 (I201566,I1869);
or I_11746 (I201583,I4001,I3989);
nor I_11747 (I201600,I201583,I3983);
nor I_11748 (I201617,I3986,I3995);
or I_11749 (I201634,I201617,I3998);
nor I_11750 (I201651,I3980,I3983);
nand I_11751 (I201668,I201651,I201634);
not I_11752 (I201685,I201668);
nand I_11753 (I201702,I201600,I201685);
nor I_11754 (I201719,I201600,I201685);
nand I_11755 (I201736,I3986,I3992);
nor I_11756 (I201753,I201736,I3980);
nor I_11757 (I201770,I201736,I201753);
not I_11758 (I201787,I201753);
nor I_11759 (I201558,I201787,I201702);
or I_11760 (I201543,I201600,I201787);
nor I_11761 (I201832,I201600,I201753);
nor I_11762 (I201537,I201736,I201832);
nor I_11763 (I201863,I201770,I201832);
nor I_11764 (I201540,I201685,I201863);
nand I_11765 (I201894,I201600,I201753);
nand I_11766 (I201911,I201668,I201894);
DFFARX1 I_11767 (I201911,I1862,I201566,I201546,);
not I_11768 (I201942,I201736);
nor I_11769 (I201555,I201942,I201787);
nand I_11770 (I201552,I201719,I201942);
nor I_11771 (I201987,I201685,I201736);
nand I_11772 (I201549,I201987,I201600);
not I_11773 (I202042,I1869);
or I_11774 (I202059,I83353,I83362);
nor I_11775 (I202076,I202059,I83377);
nor I_11776 (I202093,I83374,I83356);
or I_11777 (I202110,I202093,I83356);
nor I_11778 (I202127,I83353,I83359);
nand I_11779 (I202144,I202127,I202110);
not I_11780 (I202161,I202144);
nand I_11781 (I202178,I202076,I202161);
nor I_11782 (I202195,I202076,I202161);
nand I_11783 (I202212,I83365,I83368);
nor I_11784 (I202229,I202212,I83371);
nor I_11785 (I202246,I202212,I202229);
not I_11786 (I202263,I202229);
nor I_11787 (I202034,I202263,I202178);
or I_11788 (I202019,I202076,I202263);
nor I_11789 (I202308,I202076,I202229);
nor I_11790 (I202013,I202212,I202308);
nor I_11791 (I202339,I202246,I202308);
nor I_11792 (I202016,I202161,I202339);
nand I_11793 (I202370,I202076,I202229);
nand I_11794 (I202387,I202144,I202370);
DFFARX1 I_11795 (I202387,I1862,I202042,I202022,);
not I_11796 (I202418,I202212);
nor I_11797 (I202031,I202418,I202263);
nand I_11798 (I202028,I202195,I202418);
nor I_11799 (I202463,I202161,I202212);
nand I_11800 (I202025,I202463,I202076);
not I_11801 (I202518,I1869);
or I_11802 (I202535,I67543,I67552);
nor I_11803 (I202552,I202535,I67567);
nor I_11804 (I202569,I67564,I67546);
or I_11805 (I202586,I202569,I67546);
nor I_11806 (I202603,I67543,I67549);
nand I_11807 (I202620,I202603,I202586);
not I_11808 (I202637,I202620);
nand I_11809 (I202654,I202552,I202637);
nor I_11810 (I202671,I202552,I202637);
nand I_11811 (I202688,I67555,I67558);
nor I_11812 (I202705,I202688,I67561);
nor I_11813 (I202722,I202688,I202705);
not I_11814 (I202739,I202705);
nor I_11815 (I202510,I202739,I202654);
or I_11816 (I202495,I202552,I202739);
nor I_11817 (I202784,I202552,I202705);
nor I_11818 (I202489,I202688,I202784);
nor I_11819 (I202815,I202722,I202784);
nor I_11820 (I202492,I202637,I202815);
nand I_11821 (I202846,I202552,I202705);
nand I_11822 (I202863,I202620,I202846);
DFFARX1 I_11823 (I202863,I1862,I202518,I202498,);
not I_11824 (I202894,I202688);
nor I_11825 (I202507,I202894,I202739);
nand I_11826 (I202504,I202671,I202894);
nor I_11827 (I202939,I202637,I202688);
nand I_11828 (I202501,I202939,I202552);
not I_11829 (I202994,I1869);
or I_11830 (I203011,I177421,I177406);
nor I_11831 (I203028,I203011,I177400);
nor I_11832 (I203045,I177397,I177418);
or I_11833 (I203062,I203045,I177415);
nor I_11834 (I203079,I177403,I177400);
nand I_11835 (I203096,I203079,I203062);
not I_11836 (I203113,I203096);
nand I_11837 (I203130,I203028,I203113);
nor I_11838 (I203147,I203028,I203113);
nand I_11839 (I203164,I177409,I177412);
nor I_11840 (I203181,I203164,I177397);
nor I_11841 (I203198,I203164,I203181);
not I_11842 (I203215,I203181);
nor I_11843 (I202986,I203215,I203130);
or I_11844 (I202971,I203028,I203215);
nor I_11845 (I203260,I203028,I203181);
nor I_11846 (I202965,I203164,I203260);
nor I_11847 (I203291,I203198,I203260);
nor I_11848 (I202968,I203113,I203291);
nand I_11849 (I203322,I203028,I203181);
nand I_11850 (I203339,I203096,I203322);
DFFARX1 I_11851 (I203339,I1862,I202994,I202974,);
not I_11852 (I203370,I203164);
nor I_11853 (I202983,I203370,I203215);
nand I_11854 (I202980,I203147,I203370);
nor I_11855 (I203415,I203113,I203164);
nand I_11856 (I202977,I203415,I203028);
not I_11857 (I203470,I1869);
or I_11858 (I203487,I158449,I158434);
nor I_11859 (I203504,I203487,I158428);
nor I_11860 (I203521,I158425,I158446);
or I_11861 (I203538,I203521,I158443);
nor I_11862 (I203555,I158431,I158428);
nand I_11863 (I203572,I203555,I203538);
not I_11864 (I203589,I203572);
nand I_11865 (I203606,I203504,I203589);
nor I_11866 (I203623,I203504,I203589);
nand I_11867 (I203640,I158437,I158440);
nor I_11868 (I203657,I203640,I158425);
nor I_11869 (I203674,I203640,I203657);
not I_11870 (I203691,I203657);
nor I_11871 (I203462,I203691,I203606);
or I_11872 (I203447,I203504,I203691);
nor I_11873 (I203736,I203504,I203657);
nor I_11874 (I203441,I203640,I203736);
nor I_11875 (I203767,I203674,I203736);
nor I_11876 (I203444,I203589,I203767);
nand I_11877 (I203798,I203504,I203657);
nand I_11878 (I203815,I203572,I203798);
DFFARX1 I_11879 (I203815,I1862,I203470,I203450,);
not I_11880 (I203846,I203640);
nor I_11881 (I203459,I203846,I203691);
nand I_11882 (I203456,I203623,I203846);
nor I_11883 (I203891,I203589,I203640);
nand I_11884 (I203453,I203891,I203504);
not I_11885 (I203946,I1869);
or I_11886 (I203963,I399063,I399066);
nor I_11887 (I203980,I203963,I399063);
nor I_11888 (I203997,I399060,I399078);
or I_11889 (I204014,I203997,I399066);
nor I_11890 (I204031,I399069,I399060);
nand I_11891 (I204048,I204031,I204014);
not I_11892 (I204065,I204048);
nand I_11893 (I204082,I203980,I204065);
nor I_11894 (I204099,I203980,I204065);
nand I_11895 (I204116,I399075,I399072);
nor I_11896 (I204133,I204116,I399069);
nor I_11897 (I204150,I204116,I204133);
not I_11898 (I204167,I204133);
nor I_11899 (I203938,I204167,I204082);
or I_11900 (I203923,I203980,I204167);
nor I_11901 (I204212,I203980,I204133);
nor I_11902 (I203917,I204116,I204212);
nor I_11903 (I204243,I204150,I204212);
nor I_11904 (I203920,I204065,I204243);
nand I_11905 (I204274,I203980,I204133);
nand I_11906 (I204291,I204048,I204274);
DFFARX1 I_11907 (I204291,I1862,I203946,I203926,);
not I_11908 (I204322,I204116);
nor I_11909 (I203935,I204322,I204167);
nand I_11910 (I203932,I204099,I204322);
nor I_11911 (I204367,I204065,I204116);
nand I_11912 (I203929,I204367,I203980);
not I_11913 (I204422,I1869);
or I_11914 (I204439,I153706,I153691);
nor I_11915 (I204456,I204439,I153685);
nor I_11916 (I204473,I153682,I153703);
or I_11917 (I204490,I204473,I153700);
nor I_11918 (I204507,I153688,I153685);
nand I_11919 (I204524,I204507,I204490);
not I_11920 (I204541,I204524);
nand I_11921 (I204558,I204456,I204541);
nor I_11922 (I204575,I204456,I204541);
nand I_11923 (I204592,I153694,I153697);
nor I_11924 (I204609,I204592,I153682);
nor I_11925 (I204626,I204592,I204609);
not I_11926 (I204643,I204609);
nor I_11927 (I204414,I204643,I204558);
or I_11928 (I204399,I204456,I204643);
nor I_11929 (I204688,I204456,I204609);
nor I_11930 (I204393,I204592,I204688);
nor I_11931 (I204719,I204626,I204688);
nor I_11932 (I204396,I204541,I204719);
nand I_11933 (I204750,I204456,I204609);
nand I_11934 (I204767,I204524,I204750);
DFFARX1 I_11935 (I204767,I1862,I204422,I204402,);
not I_11936 (I204798,I204592);
nor I_11937 (I204411,I204798,I204643);
nand I_11938 (I204408,I204575,I204798);
nor I_11939 (I204843,I204541,I204592);
nand I_11940 (I204405,I204843,I204456);
not I_11941 (I204898,I1869);
or I_11942 (I204915,I162138,I162123);
nor I_11943 (I204932,I204915,I162117);
nor I_11944 (I204949,I162114,I162135);
or I_11945 (I204966,I204949,I162132);
nor I_11946 (I204983,I162120,I162117);
nand I_11947 (I205000,I204983,I204966);
not I_11948 (I205017,I205000);
nand I_11949 (I205034,I204932,I205017);
nor I_11950 (I205051,I204932,I205017);
nand I_11951 (I205068,I162126,I162129);
nor I_11952 (I205085,I205068,I162114);
nor I_11953 (I205102,I205068,I205085);
not I_11954 (I205119,I205085);
nor I_11955 (I204890,I205119,I205034);
or I_11956 (I204875,I204932,I205119);
nor I_11957 (I205164,I204932,I205085);
nor I_11958 (I204869,I205068,I205164);
nor I_11959 (I205195,I205102,I205164);
nor I_11960 (I204872,I205017,I205195);
nand I_11961 (I205226,I204932,I205085);
nand I_11962 (I205243,I205000,I205226);
DFFARX1 I_11963 (I205243,I1862,I204898,I204878,);
not I_11964 (I205274,I205068);
nor I_11965 (I204887,I205274,I205119);
nand I_11966 (I204884,I205051,I205274);
nor I_11967 (I205319,I205017,I205068);
nand I_11968 (I204881,I205319,I204932);
not I_11969 (I205374,I1869);
or I_11970 (I205391,I384477,I384480);
nor I_11971 (I205408,I205391,I384477);
nor I_11972 (I205425,I384474,I384492);
or I_11973 (I205442,I205425,I384480);
nor I_11974 (I205459,I384483,I384474);
nand I_11975 (I205476,I205459,I205442);
not I_11976 (I205493,I205476);
nand I_11977 (I205510,I205408,I205493);
nor I_11978 (I205527,I205408,I205493);
nand I_11979 (I205544,I384489,I384486);
nor I_11980 (I205561,I205544,I384483);
nor I_11981 (I205578,I205544,I205561);
not I_11982 (I205595,I205561);
nor I_11983 (I205366,I205595,I205510);
or I_11984 (I205351,I205408,I205595);
nor I_11985 (I205640,I205408,I205561);
nor I_11986 (I205345,I205544,I205640);
nor I_11987 (I205671,I205578,I205640);
nor I_11988 (I205348,I205493,I205671);
nand I_11989 (I205702,I205408,I205561);
nand I_11990 (I205719,I205476,I205702);
DFFARX1 I_11991 (I205719,I1862,I205374,I205354,);
not I_11992 (I205750,I205544);
nor I_11993 (I205363,I205750,I205595);
nand I_11994 (I205360,I205527,I205750);
nor I_11995 (I205795,I205493,I205544);
nand I_11996 (I205357,I205795,I205408);
not I_11997 (I205850,I1869);
or I_11998 (I205867,I123140,I123125);
nor I_11999 (I205884,I205867,I123119);
nor I_12000 (I205901,I123116,I123137);
or I_12001 (I205918,I205901,I123134);
nor I_12002 (I205935,I123122,I123119);
nand I_12003 (I205952,I205935,I205918);
not I_12004 (I205969,I205952);
nand I_12005 (I205986,I205884,I205969);
nor I_12006 (I206003,I205884,I205969);
nand I_12007 (I206020,I123128,I123131);
nor I_12008 (I206037,I206020,I123116);
nor I_12009 (I206054,I206020,I206037);
not I_12010 (I206071,I206037);
nor I_12011 (I205842,I206071,I205986);
or I_12012 (I205827,I205884,I206071);
nor I_12013 (I206116,I205884,I206037);
nor I_12014 (I205821,I206020,I206116);
nor I_12015 (I206147,I206054,I206116);
nor I_12016 (I205824,I205969,I206147);
nand I_12017 (I206178,I205884,I206037);
nand I_12018 (I206195,I205952,I206178);
DFFARX1 I_12019 (I206195,I1862,I205850,I205830,);
not I_12020 (I206226,I206020);
nor I_12021 (I205839,I206226,I206071);
nand I_12022 (I205836,I206003,I206226);
nor I_12023 (I206271,I205969,I206020);
nand I_12024 (I205833,I206271,I205884);
not I_12025 (I206326,I1869);
or I_12026 (I206343,I197447,I197432);
nor I_12027 (I206360,I206343,I197426);
nor I_12028 (I206377,I197423,I197444);
or I_12029 (I206394,I206377,I197441);
nor I_12030 (I206411,I197429,I197426);
nand I_12031 (I206428,I206411,I206394);
not I_12032 (I206445,I206428);
nand I_12033 (I206462,I206360,I206445);
nor I_12034 (I206479,I206360,I206445);
nand I_12035 (I206496,I197435,I197438);
nor I_12036 (I206513,I206496,I197423);
nor I_12037 (I206530,I206496,I206513);
not I_12038 (I206547,I206513);
nor I_12039 (I206318,I206547,I206462);
or I_12040 (I206303,I206360,I206547);
nor I_12041 (I206592,I206360,I206513);
nor I_12042 (I206297,I206496,I206592);
nor I_12043 (I206623,I206530,I206592);
nor I_12044 (I206300,I206445,I206623);
nand I_12045 (I206654,I206360,I206513);
nand I_12046 (I206671,I206428,I206654);
DFFARX1 I_12047 (I206671,I1862,I206326,I206306,);
not I_12048 (I206702,I206496);
nor I_12049 (I206315,I206702,I206547);
nand I_12050 (I206312,I206479,I206702);
nor I_12051 (I206747,I206445,I206496);
nand I_12052 (I206309,I206747,I206360);
not I_12053 (I206802,I1869);
or I_12054 (I206819,I47653,I47662);
nor I_12055 (I206836,I206819,I47677);
nor I_12056 (I206853,I47674,I47656);
or I_12057 (I206870,I206853,I47656);
nor I_12058 (I206887,I47653,I47659);
nand I_12059 (I206904,I206887,I206870);
not I_12060 (I206921,I206904);
nand I_12061 (I206938,I206836,I206921);
nor I_12062 (I206955,I206836,I206921);
nand I_12063 (I206972,I47665,I47668);
nor I_12064 (I206989,I206972,I47671);
nor I_12065 (I207006,I206972,I206989);
not I_12066 (I207023,I206989);
nor I_12067 (I206794,I207023,I206938);
or I_12068 (I206779,I206836,I207023);
nor I_12069 (I207068,I206836,I206989);
nor I_12070 (I206773,I206972,I207068);
nor I_12071 (I207099,I207006,I207068);
nor I_12072 (I206776,I206921,I207099);
nand I_12073 (I207130,I206836,I206989);
nand I_12074 (I207147,I206904,I207130);
DFFARX1 I_12075 (I207147,I1862,I206802,I206782,);
not I_12076 (I207178,I206972);
nor I_12077 (I206791,I207178,I207023);
nand I_12078 (I206788,I206955,I207178);
nor I_12079 (I207223,I206921,I206972);
nand I_12080 (I206785,I207223,I206836);
not I_12081 (I207278,I1869);
or I_12082 (I207295,I403483,I403486);
nor I_12083 (I207312,I207295,I403483);
nor I_12084 (I207329,I403480,I403498);
or I_12085 (I207346,I207329,I403486);
nor I_12086 (I207363,I403489,I403480);
nand I_12087 (I207380,I207363,I207346);
not I_12088 (I207397,I207380);
nand I_12089 (I207414,I207312,I207397);
nor I_12090 (I207431,I207312,I207397);
nand I_12091 (I207448,I403495,I403492);
nor I_12092 (I207465,I207448,I403489);
nor I_12093 (I207482,I207448,I207465);
not I_12094 (I207499,I207465);
nor I_12095 (I207270,I207499,I207414);
or I_12096 (I207255,I207312,I207499);
nor I_12097 (I207544,I207312,I207465);
nor I_12098 (I207249,I207448,I207544);
nor I_12099 (I207575,I207482,I207544);
nor I_12100 (I207252,I207397,I207575);
nand I_12101 (I207606,I207312,I207465);
nand I_12102 (I207623,I207380,I207606);
DFFARX1 I_12103 (I207623,I1862,I207278,I207258,);
not I_12104 (I207654,I207448);
nor I_12105 (I207267,I207654,I207499);
nand I_12106 (I207264,I207431,I207654);
nor I_12107 (I207699,I207397,I207448);
nand I_12108 (I207261,I207699,I207312);
not I_12109 (I207754,I1869);
or I_12110 (I207771,I345765,I345786);
nor I_12111 (I207788,I207771,I345771);
nor I_12112 (I207805,I345765,I345783);
or I_12113 (I207822,I207805,I345774);
nor I_12114 (I207839,I345768,I345768);
nand I_12115 (I207856,I207839,I207822);
not I_12116 (I207873,I207856);
nand I_12117 (I207890,I207788,I207873);
nor I_12118 (I207907,I207788,I207873);
nand I_12119 (I207924,I345777,I345780);
nor I_12120 (I207941,I207924,I345771);
nor I_12121 (I207958,I207924,I207941);
not I_12122 (I207975,I207941);
nor I_12123 (I207746,I207975,I207890);
or I_12124 (I207731,I207788,I207975);
nor I_12125 (I208020,I207788,I207941);
nor I_12126 (I207725,I207924,I208020);
nor I_12127 (I208051,I207958,I208020);
nor I_12128 (I207728,I207873,I208051);
nand I_12129 (I208082,I207788,I207941);
nand I_12130 (I208099,I207856,I208082);
DFFARX1 I_12131 (I208099,I1862,I207754,I207734,);
not I_12132 (I208130,I207924);
nor I_12133 (I207743,I208130,I207975);
nand I_12134 (I207740,I207907,I208130);
nor I_12135 (I208175,I207873,I207924);
nand I_12136 (I207737,I208175,I207788);
not I_12137 (I208230,I1869);
or I_12138 (I208247,I338387,I338408);
nor I_12139 (I208264,I208247,I338393);
nor I_12140 (I208281,I338387,I338405);
or I_12141 (I208298,I208281,I338396);
nor I_12142 (I208315,I338390,I338390);
nand I_12143 (I208332,I208315,I208298);
not I_12144 (I208349,I208332);
nand I_12145 (I208366,I208264,I208349);
nor I_12146 (I208383,I208264,I208349);
nand I_12147 (I208400,I338399,I338402);
nor I_12148 (I208417,I208400,I338393);
nor I_12149 (I208434,I208400,I208417);
not I_12150 (I208451,I208417);
nor I_12151 (I208222,I208451,I208366);
or I_12152 (I208207,I208264,I208451);
nor I_12153 (I208496,I208264,I208417);
nor I_12154 (I208201,I208400,I208496);
nor I_12155 (I208527,I208434,I208496);
nor I_12156 (I208204,I208349,I208527);
nand I_12157 (I208558,I208264,I208417);
nand I_12158 (I208575,I208332,I208558);
DFFARX1 I_12159 (I208575,I1862,I208230,I208210,);
not I_12160 (I208606,I208400);
nor I_12161 (I208219,I208606,I208451);
nand I_12162 (I208216,I208383,I208606);
nor I_12163 (I208651,I208349,I208400);
nand I_12164 (I208213,I208651,I208264);
not I_12165 (I208706,I1869);
or I_12166 (I208723,I31333,I31342);
nor I_12167 (I208740,I208723,I31357);
nor I_12168 (I208757,I31354,I31336);
or I_12169 (I208774,I208757,I31336);
nor I_12170 (I208791,I31333,I31339);
nand I_12171 (I208808,I208791,I208774);
not I_12172 (I208825,I208808);
nand I_12173 (I208842,I208740,I208825);
nor I_12174 (I208859,I208740,I208825);
nand I_12175 (I208876,I31345,I31348);
nor I_12176 (I208893,I208876,I31351);
nor I_12177 (I208910,I208876,I208893);
not I_12178 (I208927,I208893);
nor I_12179 (I208698,I208927,I208842);
or I_12180 (I208683,I208740,I208927);
nor I_12181 (I208972,I208740,I208893);
nor I_12182 (I208677,I208876,I208972);
nor I_12183 (I209003,I208910,I208972);
nor I_12184 (I208680,I208825,I209003);
nand I_12185 (I209034,I208740,I208893);
nand I_12186 (I209051,I208808,I209034);
DFFARX1 I_12187 (I209051,I1862,I208706,I208686,);
not I_12188 (I209082,I208876);
nor I_12189 (I208695,I209082,I208927);
nand I_12190 (I208692,I208859,I209082);
nor I_12191 (I209127,I208825,I208876);
nand I_12192 (I208689,I209127,I208740);
not I_12193 (I209182,I1869);
or I_12194 (I209199,I48673,I48682);
nor I_12195 (I209216,I209199,I48697);
nor I_12196 (I209233,I48694,I48676);
or I_12197 (I209250,I209233,I48676);
nor I_12198 (I209267,I48673,I48679);
nand I_12199 (I209284,I209267,I209250);
not I_12200 (I209301,I209284);
nand I_12201 (I209318,I209216,I209301);
nor I_12202 (I209335,I209216,I209301);
nand I_12203 (I209352,I48685,I48688);
nor I_12204 (I209369,I209352,I48691);
nor I_12205 (I209386,I209352,I209369);
not I_12206 (I209403,I209369);
nor I_12207 (I209174,I209403,I209318);
or I_12208 (I209159,I209216,I209403);
nor I_12209 (I209448,I209216,I209369);
nor I_12210 (I209153,I209352,I209448);
nor I_12211 (I209479,I209386,I209448);
nor I_12212 (I209156,I209301,I209479);
nand I_12213 (I209510,I209216,I209369);
nand I_12214 (I209527,I209284,I209510);
DFFARX1 I_12215 (I209527,I1862,I209182,I209162,);
not I_12216 (I209558,I209352);
nor I_12217 (I209171,I209558,I209403);
nand I_12218 (I209168,I209335,I209558);
nor I_12219 (I209603,I209301,I209352);
nand I_12220 (I209165,I209603,I209216);
not I_12221 (I209658,I1869);
or I_12222 (I209675,I86413,I86422);
nor I_12223 (I209692,I209675,I86437);
nor I_12224 (I209709,I86434,I86416);
or I_12225 (I209726,I209709,I86416);
nor I_12226 (I209743,I86413,I86419);
nand I_12227 (I209760,I209743,I209726);
not I_12228 (I209777,I209760);
nand I_12229 (I209794,I209692,I209777);
nor I_12230 (I209811,I209692,I209777);
nand I_12231 (I209828,I86425,I86428);
nor I_12232 (I209845,I209828,I86431);
nor I_12233 (I209862,I209828,I209845);
not I_12234 (I209879,I209845);
nor I_12235 (I209650,I209879,I209794);
or I_12236 (I209635,I209692,I209879);
nor I_12237 (I209924,I209692,I209845);
nor I_12238 (I209629,I209828,I209924);
nor I_12239 (I209955,I209862,I209924);
nor I_12240 (I209632,I209777,I209955);
nand I_12241 (I209986,I209692,I209845);
nand I_12242 (I210003,I209760,I209986);
DFFARX1 I_12243 (I210003,I1862,I209658,I209638,);
not I_12244 (I210034,I209828);
nor I_12245 (I209647,I210034,I209879);
nand I_12246 (I209644,I209811,I210034);
nor I_12247 (I210079,I209777,I209828);
nand I_12248 (I209641,I210079,I209692);
not I_12249 (I210134,I1869);
or I_12250 (I210151,I347873,I347894);
nor I_12251 (I210168,I210151,I347879);
nor I_12252 (I210185,I347873,I347891);
or I_12253 (I210202,I210185,I347882);
nor I_12254 (I210219,I347876,I347876);
nand I_12255 (I210236,I210219,I210202);
not I_12256 (I210253,I210236);
nand I_12257 (I210270,I210168,I210253);
nor I_12258 (I210287,I210168,I210253);
nand I_12259 (I210304,I347885,I347888);
nor I_12260 (I210321,I210304,I347879);
nor I_12261 (I210338,I210304,I210321);
not I_12262 (I210355,I210321);
nor I_12263 (I210126,I210355,I210270);
or I_12264 (I210111,I210168,I210355);
nor I_12265 (I210400,I210168,I210321);
nor I_12266 (I210105,I210304,I210400);
nor I_12267 (I210431,I210338,I210400);
nor I_12268 (I210108,I210253,I210431);
nand I_12269 (I210462,I210168,I210321);
nand I_12270 (I210479,I210236,I210462);
DFFARX1 I_12271 (I210479,I1862,I210134,I210114,);
not I_12272 (I210510,I210304);
nor I_12273 (I210123,I210510,I210355);
nand I_12274 (I210120,I210287,I210510);
nor I_12275 (I210555,I210253,I210304);
nand I_12276 (I210117,I210555,I210168);
not I_12277 (I210610,I1869);
or I_12278 (I210627,I289906,I289903);
nor I_12279 (I210644,I210627,I289912);
nor I_12280 (I210661,I289924,I289909);
or I_12281 (I210678,I210661,I289903);
nor I_12282 (I210695,I289915,I289906);
nand I_12283 (I210712,I210695,I210678);
not I_12284 (I210729,I210712);
nand I_12285 (I210746,I210644,I210729);
nor I_12286 (I210763,I210644,I210729);
nand I_12287 (I210780,I289909,I289921);
nor I_12288 (I210797,I210780,I289918);
nor I_12289 (I210814,I210780,I210797);
not I_12290 (I210831,I210797);
nor I_12291 (I210602,I210831,I210746);
or I_12292 (I210587,I210644,I210831);
nor I_12293 (I210876,I210644,I210797);
nor I_12294 (I210581,I210780,I210876);
nor I_12295 (I210907,I210814,I210876);
nor I_12296 (I210584,I210729,I210907);
nand I_12297 (I210938,I210644,I210797);
nand I_12298 (I210955,I210712,I210938);
DFFARX1 I_12299 (I210955,I1862,I210610,I210590,);
not I_12300 (I210986,I210780);
nor I_12301 (I210599,I210986,I210831);
nand I_12302 (I210596,I210763,I210986);
nor I_12303 (I211031,I210729,I210780);
nand I_12304 (I210593,I211031,I210644);
not I_12305 (I211086,I1869);
or I_12306 (I211103,I41023,I41032);
nor I_12307 (I211120,I211103,I41047);
nor I_12308 (I211137,I41044,I41026);
or I_12309 (I211154,I211137,I41026);
nor I_12310 (I211171,I41023,I41029);
nand I_12311 (I211188,I211171,I211154);
not I_12312 (I211205,I211188);
nand I_12313 (I211222,I211120,I211205);
nor I_12314 (I211239,I211120,I211205);
nand I_12315 (I211256,I41035,I41038);
nor I_12316 (I211273,I211256,I41041);
nor I_12317 (I211290,I211256,I211273);
not I_12318 (I211307,I211273);
nor I_12319 (I211078,I211307,I211222);
or I_12320 (I211063,I211120,I211307);
nor I_12321 (I211352,I211120,I211273);
nor I_12322 (I211057,I211256,I211352);
nor I_12323 (I211383,I211290,I211352);
nor I_12324 (I211060,I211205,I211383);
nand I_12325 (I211414,I211120,I211273);
nand I_12326 (I211431,I211188,I211414);
DFFARX1 I_12327 (I211431,I1862,I211086,I211066,);
not I_12328 (I211462,I211256);
nor I_12329 (I211075,I211462,I211307);
nand I_12330 (I211072,I211239,I211462);
nor I_12331 (I211507,I211205,I211256);
nand I_12332 (I211069,I211507,I211120);
not I_12333 (I211562,I1869);
or I_12334 (I211579,I50713,I50722);
nor I_12335 (I211596,I211579,I50737);
nor I_12336 (I211613,I50734,I50716);
or I_12337 (I211630,I211613,I50716);
nor I_12338 (I211647,I50713,I50719);
nand I_12339 (I211664,I211647,I211630);
not I_12340 (I211681,I211664);
nand I_12341 (I211698,I211596,I211681);
nor I_12342 (I211715,I211596,I211681);
nand I_12343 (I211732,I50725,I50728);
nor I_12344 (I211749,I211732,I50731);
nor I_12345 (I211766,I211732,I211749);
not I_12346 (I211783,I211749);
nor I_12347 (I211554,I211783,I211698);
or I_12348 (I211539,I211596,I211783);
nor I_12349 (I211828,I211596,I211749);
nor I_12350 (I211533,I211732,I211828);
nor I_12351 (I211859,I211766,I211828);
nor I_12352 (I211536,I211681,I211859);
nand I_12353 (I211890,I211596,I211749);
nand I_12354 (I211907,I211664,I211890);
DFFARX1 I_12355 (I211907,I1862,I211562,I211542,);
not I_12356 (I211938,I211732);
nor I_12357 (I211551,I211938,I211783);
nand I_12358 (I211548,I211715,I211938);
nor I_12359 (I211983,I211681,I211732);
nand I_12360 (I211545,I211983,I211596);
not I_12361 (I212038,I1869);
or I_12362 (I212055,I28783,I28792);
nor I_12363 (I212072,I212055,I28807);
nor I_12364 (I212089,I28804,I28786);
or I_12365 (I212106,I212089,I28786);
nor I_12366 (I212123,I28783,I28789);
nand I_12367 (I212140,I212123,I212106);
not I_12368 (I212157,I212140);
nand I_12369 (I212174,I212072,I212157);
nor I_12370 (I212191,I212072,I212157);
nand I_12371 (I212208,I28795,I28798);
nor I_12372 (I212225,I212208,I28801);
nor I_12373 (I212242,I212208,I212225);
not I_12374 (I212259,I212225);
nor I_12375 (I212030,I212259,I212174);
or I_12376 (I212015,I212072,I212259);
nor I_12377 (I212304,I212072,I212225);
nor I_12378 (I212009,I212208,I212304);
nor I_12379 (I212335,I212242,I212304);
nor I_12380 (I212012,I212157,I212335);
nand I_12381 (I212366,I212072,I212225);
nand I_12382 (I212383,I212140,I212366);
DFFARX1 I_12383 (I212383,I1862,I212038,I212018,);
not I_12384 (I212414,I212208);
nor I_12385 (I212027,I212414,I212259);
nand I_12386 (I212024,I212191,I212414);
nor I_12387 (I212459,I212157,I212208);
nand I_12388 (I212021,I212459,I212072);
not I_12389 (I212514,I1869);
or I_12390 (I212531,I319415,I319436);
nor I_12391 (I212548,I212531,I319421);
nor I_12392 (I212565,I319415,I319433);
or I_12393 (I212582,I212565,I319424);
nor I_12394 (I212599,I319418,I319418);
nand I_12395 (I212616,I212599,I212582);
not I_12396 (I212633,I212616);
nand I_12397 (I212650,I212548,I212633);
nor I_12398 (I212667,I212548,I212633);
nand I_12399 (I212684,I319427,I319430);
nor I_12400 (I212701,I212684,I319421);
nor I_12401 (I212718,I212684,I212701);
not I_12402 (I212735,I212701);
nor I_12403 (I212506,I212735,I212650);
or I_12404 (I212491,I212548,I212735);
nor I_12405 (I212780,I212548,I212701);
nor I_12406 (I212485,I212684,I212780);
nor I_12407 (I212811,I212718,I212780);
nor I_12408 (I212488,I212633,I212811);
nand I_12409 (I212842,I212548,I212701);
nand I_12410 (I212859,I212616,I212842);
DFFARX1 I_12411 (I212859,I1862,I212514,I212494,);
not I_12412 (I212890,I212684);
nor I_12413 (I212503,I212890,I212735);
nand I_12414 (I212500,I212667,I212890);
nor I_12415 (I212935,I212633,I212684);
nand I_12416 (I212497,I212935,I212548);
not I_12417 (I212990,I1869);
or I_12418 (I213007,I390665,I390668);
nor I_12419 (I213024,I213007,I390665);
nor I_12420 (I213041,I390662,I390680);
or I_12421 (I213058,I213041,I390668);
nor I_12422 (I213075,I390671,I390662);
nand I_12423 (I213092,I213075,I213058);
not I_12424 (I213109,I213092);
nand I_12425 (I213126,I213024,I213109);
nor I_12426 (I213143,I213024,I213109);
nand I_12427 (I213160,I390677,I390674);
nor I_12428 (I213177,I213160,I390671);
nor I_12429 (I213194,I213160,I213177);
not I_12430 (I213211,I213177);
nor I_12431 (I212982,I213211,I213126);
or I_12432 (I212967,I213024,I213211);
nor I_12433 (I213256,I213024,I213177);
nor I_12434 (I212961,I213160,I213256);
nor I_12435 (I213287,I213194,I213256);
nor I_12436 (I212964,I213109,I213287);
nand I_12437 (I213318,I213024,I213177);
nand I_12438 (I213335,I213092,I213318);
DFFARX1 I_12439 (I213335,I1862,I212990,I212970,);
not I_12440 (I213366,I213160);
nor I_12441 (I212979,I213366,I213211);
nand I_12442 (I212976,I213143,I213366);
nor I_12443 (I213411,I213109,I213160);
nand I_12444 (I212973,I213411,I213024);
not I_12445 (I213466,I1869);
or I_12446 (I213483,I171624,I171609);
nor I_12447 (I213500,I213483,I171603);
nor I_12448 (I213517,I171600,I171621);
or I_12449 (I213534,I213517,I171618);
nor I_12450 (I213551,I171606,I171603);
nand I_12451 (I213568,I213551,I213534);
not I_12452 (I213585,I213568);
nand I_12453 (I213602,I213500,I213585);
nor I_12454 (I213619,I213500,I213585);
nand I_12455 (I213636,I171612,I171615);
nor I_12456 (I213653,I213636,I171600);
nor I_12457 (I213670,I213636,I213653);
not I_12458 (I213687,I213653);
nor I_12459 (I213458,I213687,I213602);
or I_12460 (I213443,I213500,I213687);
nor I_12461 (I213732,I213500,I213653);
nor I_12462 (I213437,I213636,I213732);
nor I_12463 (I213763,I213670,I213732);
nor I_12464 (I213440,I213585,I213763);
nand I_12465 (I213794,I213500,I213653);
nand I_12466 (I213811,I213568,I213794);
DFFARX1 I_12467 (I213811,I1862,I213466,I213446,);
not I_12468 (I213842,I213636);
nor I_12469 (I213455,I213842,I213687);
nand I_12470 (I213452,I213619,I213842);
nor I_12471 (I213887,I213585,I213636);
nand I_12472 (I213449,I213887,I213500);
not I_12473 (I213942,I1869);
or I_12474 (I213959,I186907,I186892);
nor I_12475 (I213976,I213959,I186886);
nor I_12476 (I213993,I186883,I186904);
or I_12477 (I214010,I213993,I186901);
nor I_12478 (I214027,I186889,I186886);
nand I_12479 (I214044,I214027,I214010);
not I_12480 (I214061,I214044);
nand I_12481 (I214078,I213976,I214061);
nor I_12482 (I214095,I213976,I214061);
nand I_12483 (I214112,I186895,I186898);
nor I_12484 (I214129,I214112,I186883);
nor I_12485 (I214146,I214112,I214129);
not I_12486 (I214163,I214129);
nor I_12487 (I213934,I214163,I214078);
or I_12488 (I213919,I213976,I214163);
nor I_12489 (I214208,I213976,I214129);
nor I_12490 (I213913,I214112,I214208);
nor I_12491 (I214239,I214146,I214208);
nor I_12492 (I213916,I214061,I214239);
nand I_12493 (I214270,I213976,I214129);
nand I_12494 (I214287,I214044,I214270);
DFFARX1 I_12495 (I214287,I1862,I213942,I213922,);
not I_12496 (I214318,I214112);
nor I_12497 (I213931,I214318,I214163);
nand I_12498 (I213928,I214095,I214318);
nor I_12499 (I214363,I214061,I214112);
nand I_12500 (I213925,I214363,I213976);
not I_12501 (I214418,I1869);
or I_12502 (I214435,I132099,I132084);
nor I_12503 (I214452,I214435,I132078);
nor I_12504 (I214469,I132075,I132096);
or I_12505 (I214486,I214469,I132093);
nor I_12506 (I214503,I132081,I132078);
nand I_12507 (I214520,I214503,I214486);
not I_12508 (I214537,I214520);
nand I_12509 (I214554,I214452,I214537);
nor I_12510 (I214571,I214452,I214537);
nand I_12511 (I214588,I132087,I132090);
nor I_12512 (I214605,I214588,I132075);
nor I_12513 (I214622,I214588,I214605);
not I_12514 (I214639,I214605);
nor I_12515 (I214410,I214639,I214554);
or I_12516 (I214395,I214452,I214639);
nor I_12517 (I214684,I214452,I214605);
nor I_12518 (I214389,I214588,I214684);
nor I_12519 (I214715,I214622,I214684);
nor I_12520 (I214392,I214537,I214715);
nand I_12521 (I214746,I214452,I214605);
nand I_12522 (I214763,I214520,I214746);
DFFARX1 I_12523 (I214763,I1862,I214418,I214398,);
not I_12524 (I214794,I214588);
nor I_12525 (I214407,I214794,I214639);
nand I_12526 (I214404,I214571,I214794);
nor I_12527 (I214839,I214537,I214588);
nand I_12528 (I214401,I214839,I214452);
not I_12529 (I214894,I1869);
or I_12530 (I214911,I321523,I321544);
nor I_12531 (I214928,I214911,I321529);
nor I_12532 (I214945,I321523,I321541);
or I_12533 (I214962,I214945,I321532);
nor I_12534 (I214979,I321526,I321526);
nand I_12535 (I214996,I214979,I214962);
not I_12536 (I215013,I214996);
nand I_12537 (I215030,I214928,I215013);
nor I_12538 (I215047,I214928,I215013);
nand I_12539 (I215064,I321535,I321538);
nor I_12540 (I215081,I215064,I321529);
nor I_12541 (I215098,I215064,I215081);
not I_12542 (I215115,I215081);
nor I_12543 (I214886,I215115,I215030);
or I_12544 (I214871,I214928,I215115);
nor I_12545 (I215160,I214928,I215081);
nor I_12546 (I214865,I215064,I215160);
nor I_12547 (I215191,I215098,I215160);
nor I_12548 (I214868,I215013,I215191);
nand I_12549 (I215222,I214928,I215081);
nand I_12550 (I215239,I214996,I215222);
DFFARX1 I_12551 (I215239,I1862,I214894,I214874,);
not I_12552 (I215270,I215064);
nor I_12553 (I214883,I215270,I215115);
nand I_12554 (I214880,I215047,I215270);
nor I_12555 (I215315,I215013,I215064);
nand I_12556 (I214877,I215315,I214928);
not I_12557 (I215370,I1869);
or I_12558 (I215387,I72133,I72142);
nor I_12559 (I215404,I215387,I72157);
nor I_12560 (I215421,I72154,I72136);
or I_12561 (I215438,I215421,I72136);
nor I_12562 (I215455,I72133,I72139);
nand I_12563 (I215472,I215455,I215438);
not I_12564 (I215489,I215472);
nand I_12565 (I215506,I215404,I215489);
nor I_12566 (I215523,I215404,I215489);
nand I_12567 (I215540,I72145,I72148);
nor I_12568 (I215557,I215540,I72151);
nor I_12569 (I215574,I215540,I215557);
not I_12570 (I215591,I215557);
nor I_12571 (I215362,I215591,I215506);
or I_12572 (I215347,I215404,I215591);
nor I_12573 (I215636,I215404,I215557);
nor I_12574 (I215341,I215540,I215636);
nor I_12575 (I215667,I215574,I215636);
nor I_12576 (I215344,I215489,I215667);
nand I_12577 (I215698,I215404,I215557);
nand I_12578 (I215715,I215472,I215698);
DFFARX1 I_12579 (I215715,I1862,I215370,I215350,);
not I_12580 (I215746,I215540);
nor I_12581 (I215359,I215746,I215591);
nand I_12582 (I215356,I215523,I215746);
nor I_12583 (I215791,I215489,I215540);
nand I_12584 (I215353,I215791,I215404);
not I_12585 (I215846,I1869);
or I_12586 (I215863,I358413,I358434);
nor I_12587 (I215880,I215863,I358419);
nor I_12588 (I215897,I358413,I358431);
or I_12589 (I215914,I215897,I358422);
nor I_12590 (I215931,I358416,I358416);
nand I_12591 (I215948,I215931,I215914);
not I_12592 (I215965,I215948);
nand I_12593 (I215982,I215880,I215965);
nor I_12594 (I215999,I215880,I215965);
nand I_12595 (I216016,I358425,I358428);
nor I_12596 (I216033,I216016,I358419);
nor I_12597 (I216050,I216016,I216033);
not I_12598 (I216067,I216033);
nor I_12599 (I215838,I216067,I215982);
or I_12600 (I215823,I215880,I216067);
nor I_12601 (I216112,I215880,I216033);
nor I_12602 (I215817,I216016,I216112);
nor I_12603 (I216143,I216050,I216112);
nor I_12604 (I215820,I215965,I216143);
nand I_12605 (I216174,I215880,I216033);
nand I_12606 (I216191,I215948,I216174);
DFFARX1 I_12607 (I216191,I1862,I215846,I215826,);
not I_12608 (I216222,I216016);
nor I_12609 (I215835,I216222,I216067);
nand I_12610 (I215832,I215999,I216222);
nor I_12611 (I216267,I215965,I216016);
nand I_12612 (I215829,I216267,I215880);
not I_12613 (I216322,I1869);
or I_12614 (I216339,I184799,I184784);
nor I_12615 (I216356,I216339,I184778);
nor I_12616 (I216373,I184775,I184796);
or I_12617 (I216390,I216373,I184793);
nor I_12618 (I216407,I184781,I184778);
nand I_12619 (I216424,I216407,I216390);
not I_12620 (I216441,I216424);
nand I_12621 (I216458,I216356,I216441);
nor I_12622 (I216475,I216356,I216441);
nand I_12623 (I216492,I184787,I184790);
nor I_12624 (I216509,I216492,I184775);
nor I_12625 (I216526,I216492,I216509);
not I_12626 (I216543,I216509);
nor I_12627 (I216314,I216543,I216458);
or I_12628 (I216299,I216356,I216543);
nor I_12629 (I216588,I216356,I216509);
nor I_12630 (I216293,I216492,I216588);
nor I_12631 (I216619,I216526,I216588);
nor I_12632 (I216296,I216441,I216619);
nand I_12633 (I216650,I216356,I216509);
nand I_12634 (I216667,I216424,I216650);
DFFARX1 I_12635 (I216667,I1862,I216322,I216302,);
not I_12636 (I216698,I216492);
nor I_12637 (I216311,I216698,I216543);
nand I_12638 (I216308,I216475,I216698);
nor I_12639 (I216743,I216441,I216492);
nand I_12640 (I216305,I216743,I216356);
not I_12641 (I216798,I1869);
or I_12642 (I216815,I369891,I369894);
nor I_12643 (I216832,I216815,I369891);
nor I_12644 (I216849,I369888,I369906);
or I_12645 (I216866,I216849,I369894);
nor I_12646 (I216883,I369897,I369888);
nand I_12647 (I216900,I216883,I216866);
not I_12648 (I216917,I216900);
nand I_12649 (I216934,I216832,I216917);
nor I_12650 (I216951,I216832,I216917);
nand I_12651 (I216968,I369903,I369900);
nor I_12652 (I216985,I216968,I369897);
nor I_12653 (I217002,I216968,I216985);
not I_12654 (I217019,I216985);
nor I_12655 (I216790,I217019,I216934);
or I_12656 (I216775,I216832,I217019);
nor I_12657 (I217064,I216832,I216985);
nor I_12658 (I216769,I216968,I217064);
nor I_12659 (I217095,I217002,I217064);
nor I_12660 (I216772,I216917,I217095);
nand I_12661 (I217126,I216832,I216985);
nand I_12662 (I217143,I216900,I217126);
DFFARX1 I_12663 (I217143,I1862,I216798,I216778,);
not I_12664 (I217174,I216968);
nor I_12665 (I216787,I217174,I217019);
nand I_12666 (I216784,I216951,I217174);
nor I_12667 (I217219,I216917,I216968);
nand I_12668 (I216781,I217219,I216832);
not I_12669 (I217274,I1869);
or I_12670 (I217291,I99673,I99682);
nor I_12671 (I217308,I217291,I99697);
nor I_12672 (I217325,I99694,I99676);
or I_12673 (I217342,I217325,I99676);
nor I_12674 (I217359,I99673,I99679);
nand I_12675 (I217376,I217359,I217342);
not I_12676 (I217393,I217376);
nand I_12677 (I217410,I217308,I217393);
nor I_12678 (I217427,I217308,I217393);
nand I_12679 (I217444,I99685,I99688);
nor I_12680 (I217461,I217444,I99691);
nor I_12681 (I217478,I217444,I217461);
not I_12682 (I217495,I217461);
nor I_12683 (I217266,I217495,I217410);
or I_12684 (I217251,I217308,I217495);
nor I_12685 (I217540,I217308,I217461);
nor I_12686 (I217245,I217444,I217540);
nor I_12687 (I217571,I217478,I217540);
nor I_12688 (I217248,I217393,I217571);
nand I_12689 (I217602,I217308,I217461);
nand I_12690 (I217619,I217376,I217602);
DFFARX1 I_12691 (I217619,I1862,I217274,I217254,);
not I_12692 (I217650,I217444);
nor I_12693 (I217263,I217650,I217495);
nand I_12694 (I217260,I217427,I217650);
nor I_12695 (I217695,I217393,I217444);
nand I_12696 (I217257,I217695,I217308);
not I_12697 (I217750,I1869);
or I_12698 (I217767,I165827,I165812);
nor I_12699 (I217784,I217767,I165806);
nor I_12700 (I217801,I165803,I165824);
or I_12701 (I217818,I217801,I165821);
nor I_12702 (I217835,I165809,I165806);
nand I_12703 (I217852,I217835,I217818);
not I_12704 (I217869,I217852);
nand I_12705 (I217886,I217784,I217869);
nor I_12706 (I217903,I217784,I217869);
nand I_12707 (I217920,I165815,I165818);
nor I_12708 (I217937,I217920,I165803);
nor I_12709 (I217954,I217920,I217937);
not I_12710 (I217971,I217937);
nor I_12711 (I217742,I217971,I217886);
or I_12712 (I217727,I217784,I217971);
nor I_12713 (I218016,I217784,I217937);
nor I_12714 (I217721,I217920,I218016);
nor I_12715 (I218047,I217954,I218016);
nor I_12716 (I217724,I217869,I218047);
nand I_12717 (I218078,I217784,I217937);
nand I_12718 (I218095,I217852,I218078);
DFFARX1 I_12719 (I218095,I1862,I217750,I217730,);
not I_12720 (I218126,I217920);
nor I_12721 (I217739,I218126,I217971);
nand I_12722 (I217736,I217903,I218126);
nor I_12723 (I218171,I217869,I217920);
nand I_12724 (I217733,I218171,I217784);
not I_12725 (I218226,I1869);
or I_12726 (I218243,I160557,I160542);
nor I_12727 (I218260,I218243,I160536);
nor I_12728 (I218277,I160533,I160554);
or I_12729 (I218294,I218277,I160551);
nor I_12730 (I218311,I160539,I160536);
nand I_12731 (I218328,I218311,I218294);
not I_12732 (I218345,I218328);
nand I_12733 (I218362,I218260,I218345);
nor I_12734 (I218379,I218260,I218345);
nand I_12735 (I218396,I160545,I160548);
nor I_12736 (I218413,I218396,I160533);
nor I_12737 (I218430,I218396,I218413);
not I_12738 (I218447,I218413);
nor I_12739 (I218218,I218447,I218362);
or I_12740 (I218203,I218260,I218447);
nor I_12741 (I218492,I218260,I218413);
nor I_12742 (I218197,I218396,I218492);
nor I_12743 (I218523,I218430,I218492);
nor I_12744 (I218200,I218345,I218523);
nand I_12745 (I218554,I218260,I218413);
nand I_12746 (I218571,I218328,I218554);
DFFARX1 I_12747 (I218571,I1862,I218226,I218206,);
not I_12748 (I218602,I218396);
nor I_12749 (I218215,I218602,I218447);
nand I_12750 (I218212,I218379,I218602);
nor I_12751 (I218647,I218345,I218396);
nand I_12752 (I218209,I218647,I218260);
not I_12753 (I218702,I1869);
or I_12754 (I218719,I394201,I394204);
nor I_12755 (I218736,I218719,I394201);
nor I_12756 (I218753,I394198,I394216);
or I_12757 (I218770,I218753,I394204);
nor I_12758 (I218787,I394207,I394198);
nand I_12759 (I218804,I218787,I218770);
not I_12760 (I218821,I218804);
nand I_12761 (I218838,I218736,I218821);
nor I_12762 (I218855,I218736,I218821);
nand I_12763 (I218872,I394213,I394210);
nor I_12764 (I218889,I218872,I394207);
nor I_12765 (I218906,I218872,I218889);
not I_12766 (I218923,I218889);
nor I_12767 (I218694,I218923,I218838);
or I_12768 (I218679,I218736,I218923);
nor I_12769 (I218968,I218736,I218889);
nor I_12770 (I218673,I218872,I218968);
nor I_12771 (I218999,I218906,I218968);
nor I_12772 (I218676,I218821,I218999);
nand I_12773 (I219030,I218736,I218889);
nand I_12774 (I219047,I218804,I219030);
DFFARX1 I_12775 (I219047,I1862,I218702,I218682,);
not I_12776 (I219078,I218872);
nor I_12777 (I218691,I219078,I218923);
nand I_12778 (I218688,I218855,I219078);
nor I_12779 (I219123,I218821,I218872);
nand I_12780 (I218685,I219123,I218736);
not I_12781 (I219178,I1869);
or I_12782 (I219195,I199028,I199013);
nor I_12783 (I219212,I219195,I199007);
nor I_12784 (I219229,I199004,I199025);
or I_12785 (I219246,I219229,I199022);
nor I_12786 (I219263,I199010,I199007);
nand I_12787 (I219280,I219263,I219246);
not I_12788 (I219297,I219280);
nand I_12789 (I219314,I219212,I219297);
nor I_12790 (I219331,I219212,I219297);
nand I_12791 (I219348,I199016,I199019);
nor I_12792 (I219365,I219348,I199004);
nor I_12793 (I219382,I219348,I219365);
not I_12794 (I219399,I219365);
nor I_12795 (I219170,I219399,I219314);
or I_12796 (I219155,I219212,I219399);
nor I_12797 (I219444,I219212,I219365);
nor I_12798 (I219149,I219348,I219444);
nor I_12799 (I219475,I219382,I219444);
nor I_12800 (I219152,I219297,I219475);
nand I_12801 (I219506,I219212,I219365);
nand I_12802 (I219523,I219280,I219506);
DFFARX1 I_12803 (I219523,I1862,I219178,I219158,);
not I_12804 (I219554,I219348);
nor I_12805 (I219167,I219554,I219399);
nand I_12806 (I219164,I219331,I219554);
nor I_12807 (I219599,I219297,I219348);
nand I_12808 (I219161,I219599,I219212);
not I_12809 (I219654,I1869);
or I_12810 (I219671,I127356,I127341);
nor I_12811 (I219688,I219671,I127335);
nor I_12812 (I219705,I127332,I127353);
or I_12813 (I219722,I219705,I127350);
nor I_12814 (I219739,I127338,I127335);
nand I_12815 (I219756,I219739,I219722);
not I_12816 (I219773,I219756);
nand I_12817 (I219790,I219688,I219773);
nor I_12818 (I219807,I219688,I219773);
nand I_12819 (I219824,I127344,I127347);
nor I_12820 (I219841,I219824,I127332);
nor I_12821 (I219858,I219824,I219841);
not I_12822 (I219875,I219841);
nor I_12823 (I219646,I219875,I219790);
or I_12824 (I219631,I219688,I219875);
nor I_12825 (I219920,I219688,I219841);
nor I_12826 (I219625,I219824,I219920);
nor I_12827 (I219951,I219858,I219920);
nor I_12828 (I219628,I219773,I219951);
nand I_12829 (I219982,I219688,I219841);
nand I_12830 (I219999,I219756,I219982);
DFFARX1 I_12831 (I219999,I1862,I219654,I219634,);
not I_12832 (I220030,I219824);
nor I_12833 (I219643,I220030,I219875);
nand I_12834 (I219640,I219807,I220030);
nor I_12835 (I220075,I219773,I219824);
nand I_12836 (I219637,I220075,I219688);
not I_12837 (I220130,I1869);
or I_12838 (I220147,I301500,I301497);
nor I_12839 (I220164,I220147,I301506);
nor I_12840 (I220181,I301518,I301503);
or I_12841 (I220198,I220181,I301497);
nor I_12842 (I220215,I301509,I301500);
nand I_12843 (I220232,I220215,I220198);
not I_12844 (I220249,I220232);
nand I_12845 (I220266,I220164,I220249);
nor I_12846 (I220283,I220164,I220249);
nand I_12847 (I220300,I301503,I301515);
nor I_12848 (I220317,I220300,I301512);
nor I_12849 (I220334,I220300,I220317);
not I_12850 (I220351,I220317);
nor I_12851 (I220122,I220351,I220266);
or I_12852 (I220107,I220164,I220351);
nor I_12853 (I220396,I220164,I220317);
nor I_12854 (I220101,I220300,I220396);
nor I_12855 (I220427,I220334,I220396);
nor I_12856 (I220104,I220249,I220427);
nand I_12857 (I220458,I220164,I220317);
nand I_12858 (I220475,I220232,I220458);
DFFARX1 I_12859 (I220475,I1862,I220130,I220110,);
not I_12860 (I220506,I220300);
nor I_12861 (I220119,I220506,I220351);
nand I_12862 (I220116,I220283,I220506);
nor I_12863 (I220551,I220249,I220300);
nand I_12864 (I220113,I220551,I220164);
not I_12865 (I220606,I1869);
or I_12866 (I220623,I408787,I408790);
nor I_12867 (I220640,I220623,I408787);
nor I_12868 (I220657,I408784,I408802);
or I_12869 (I220674,I220657,I408790);
nor I_12870 (I220691,I408793,I408784);
nand I_12871 (I220708,I220691,I220674);
not I_12872 (I220725,I220708);
nand I_12873 (I220742,I220640,I220725);
nor I_12874 (I220759,I220640,I220725);
nand I_12875 (I220776,I408799,I408796);
nor I_12876 (I220793,I220776,I408793);
nor I_12877 (I220810,I220776,I220793);
not I_12878 (I220827,I220793);
nor I_12879 (I220598,I220827,I220742);
or I_12880 (I220583,I220640,I220827);
nor I_12881 (I220872,I220640,I220793);
nor I_12882 (I220577,I220776,I220872);
nor I_12883 (I220903,I220810,I220872);
nor I_12884 (I220580,I220725,I220903);
nand I_12885 (I220934,I220640,I220793);
nand I_12886 (I220951,I220708,I220934);
DFFARX1 I_12887 (I220951,I1862,I220606,I220586,);
not I_12888 (I220982,I220776);
nor I_12889 (I220595,I220982,I220827);
nand I_12890 (I220592,I220759,I220982);
nor I_12891 (I221027,I220725,I220776);
nand I_12892 (I220589,I221027,I220640);
not I_12893 (I221082,I1869);
or I_12894 (I221099,I290960,I290957);
nor I_12895 (I221116,I221099,I290966);
nor I_12896 (I221133,I290978,I290963);
or I_12897 (I221150,I221133,I290957);
nor I_12898 (I221167,I290969,I290960);
nand I_12899 (I221184,I221167,I221150);
not I_12900 (I221201,I221184);
nand I_12901 (I221218,I221116,I221201);
nor I_12902 (I221235,I221116,I221201);
nand I_12903 (I221252,I290963,I290975);
nor I_12904 (I221269,I221252,I290972);
nor I_12905 (I221286,I221252,I221269);
not I_12906 (I221303,I221269);
nor I_12907 (I221074,I221303,I221218);
or I_12908 (I221059,I221116,I221303);
nor I_12909 (I221348,I221116,I221269);
nor I_12910 (I221053,I221252,I221348);
nor I_12911 (I221379,I221286,I221348);
nor I_12912 (I221056,I221201,I221379);
nand I_12913 (I221410,I221116,I221269);
nand I_12914 (I221427,I221184,I221410);
DFFARX1 I_12915 (I221427,I1862,I221082,I221062,);
not I_12916 (I221458,I221252);
nor I_12917 (I221071,I221458,I221303);
nand I_12918 (I221068,I221235,I221458);
nor I_12919 (I221503,I221201,I221252);
nand I_12920 (I221065,I221503,I221116);
not I_12921 (I221558,I1869);
or I_12922 (I221575,I35413,I35422);
nor I_12923 (I221592,I221575,I35437);
nor I_12924 (I221609,I35434,I35416);
or I_12925 (I221626,I221609,I35416);
nor I_12926 (I221643,I35413,I35419);
nand I_12927 (I221660,I221643,I221626);
not I_12928 (I221677,I221660);
nand I_12929 (I221694,I221592,I221677);
nor I_12930 (I221711,I221592,I221677);
nand I_12931 (I221728,I35425,I35428);
nor I_12932 (I221745,I221728,I35431);
nor I_12933 (I221762,I221728,I221745);
not I_12934 (I221779,I221745);
nor I_12935 (I221550,I221779,I221694);
or I_12936 (I221535,I221592,I221779);
nor I_12937 (I221824,I221592,I221745);
nor I_12938 (I221529,I221728,I221824);
nor I_12939 (I221855,I221762,I221824);
nor I_12940 (I221532,I221677,I221855);
nand I_12941 (I221886,I221592,I221745);
nand I_12942 (I221903,I221660,I221886);
DFFARX1 I_12943 (I221903,I1862,I221558,I221538,);
not I_12944 (I221934,I221728);
nor I_12945 (I221547,I221934,I221779);
nand I_12946 (I221544,I221711,I221934);
nor I_12947 (I221979,I221677,I221728);
nand I_12948 (I221541,I221979,I221592);
not I_12949 (I222034,I1869);
or I_12950 (I222051,I131572,I131557);
nor I_12951 (I222068,I222051,I131551);
nor I_12952 (I222085,I131548,I131569);
or I_12953 (I222102,I222085,I131566);
nor I_12954 (I222119,I131554,I131551);
nand I_12955 (I222136,I222119,I222102);
not I_12956 (I222153,I222136);
nand I_12957 (I222170,I222068,I222153);
nor I_12958 (I222187,I222068,I222153);
nand I_12959 (I222204,I131560,I131563);
nor I_12960 (I222221,I222204,I131548);
nor I_12961 (I222238,I222204,I222221);
not I_12962 (I222255,I222221);
nor I_12963 (I222026,I222255,I222170);
or I_12964 (I222011,I222068,I222255);
nor I_12965 (I222300,I222068,I222221);
nor I_12966 (I222005,I222204,I222300);
nor I_12967 (I222331,I222238,I222300);
nor I_12968 (I222008,I222153,I222331);
nand I_12969 (I222362,I222068,I222221);
nand I_12970 (I222379,I222136,I222362);
DFFARX1 I_12971 (I222379,I1862,I222034,I222014,);
not I_12972 (I222410,I222204);
nor I_12973 (I222023,I222410,I222255);
nand I_12974 (I222020,I222187,I222410);
nor I_12975 (I222455,I222153,I222204);
nand I_12976 (I222017,I222455,I222068);
not I_12977 (I222510,I1869);
or I_12978 (I222527,I327320,I327341);
nor I_12979 (I222544,I222527,I327326);
nor I_12980 (I222561,I327320,I327338);
or I_12981 (I222578,I222561,I327329);
nor I_12982 (I222595,I327323,I327323);
nand I_12983 (I222612,I222595,I222578);
not I_12984 (I222629,I222612);
nand I_12985 (I222646,I222544,I222629);
nor I_12986 (I222663,I222544,I222629);
nand I_12987 (I222680,I327332,I327335);
nor I_12988 (I222697,I222680,I327326);
nor I_12989 (I222714,I222680,I222697);
not I_12990 (I222731,I222697);
nor I_12991 (I222502,I222731,I222646);
or I_12992 (I222487,I222544,I222731);
nor I_12993 (I222776,I222544,I222697);
nor I_12994 (I222481,I222680,I222776);
nor I_12995 (I222807,I222714,I222776);
nor I_12996 (I222484,I222629,I222807);
nand I_12997 (I222838,I222544,I222697);
nand I_12998 (I222855,I222612,I222838);
DFFARX1 I_12999 (I222855,I1862,I222510,I222490,);
not I_13000 (I222886,I222680);
nor I_13001 (I222499,I222886,I222731);
nand I_13002 (I222496,I222663,I222886);
nor I_13003 (I222931,I222629,I222680);
nand I_13004 (I222493,I222931,I222544);
not I_13005 (I222986,I1869);
or I_13006 (I223003,I168462,I168447);
nor I_13007 (I223020,I223003,I168441);
nor I_13008 (I223037,I168438,I168459);
or I_13009 (I223054,I223037,I168456);
nor I_13010 (I223071,I168444,I168441);
nand I_13011 (I223088,I223071,I223054);
not I_13012 (I223105,I223088);
nand I_13013 (I223122,I223020,I223105);
nor I_13014 (I223139,I223020,I223105);
nand I_13015 (I223156,I168450,I168453);
nor I_13016 (I223173,I223156,I168438);
nor I_13017 (I223190,I223156,I223173);
not I_13018 (I223207,I223173);
nor I_13019 (I222978,I223207,I223122);
or I_13020 (I222963,I223020,I223207);
nor I_13021 (I223252,I223020,I223173);
nor I_13022 (I222957,I223156,I223252);
nor I_13023 (I223283,I223190,I223252);
nor I_13024 (I222960,I223105,I223283);
nand I_13025 (I223314,I223020,I223173);
nand I_13026 (I223331,I223088,I223314);
DFFARX1 I_13027 (I223331,I1862,I222986,I222966,);
not I_13028 (I223362,I223156);
nor I_13029 (I222975,I223362,I223207);
nand I_13030 (I222972,I223139,I223362);
nor I_13031 (I223407,I223105,I223156);
nand I_13032 (I222969,I223407,I223020);
not I_13033 (I223462,I1869);
or I_13034 (I223479,I53773,I53782);
nor I_13035 (I223496,I223479,I53797);
nor I_13036 (I223513,I53794,I53776);
or I_13037 (I223530,I223513,I53776);
nor I_13038 (I223547,I53773,I53779);
nand I_13039 (I223564,I223547,I223530);
not I_13040 (I223581,I223564);
nand I_13041 (I223598,I223496,I223581);
nor I_13042 (I223615,I223496,I223581);
nand I_13043 (I223632,I53785,I53788);
nor I_13044 (I223649,I223632,I53791);
nor I_13045 (I223666,I223632,I223649);
not I_13046 (I223683,I223649);
nor I_13047 (I223454,I223683,I223598);
or I_13048 (I223439,I223496,I223683);
nor I_13049 (I223728,I223496,I223649);
nor I_13050 (I223433,I223632,I223728);
nor I_13051 (I223759,I223666,I223728);
nor I_13052 (I223436,I223581,I223759);
nand I_13053 (I223790,I223496,I223649);
nand I_13054 (I223807,I223564,I223790);
DFFARX1 I_13055 (I223807,I1862,I223462,I223442,);
not I_13056 (I223838,I223632);
nor I_13057 (I223451,I223838,I223683);
nand I_13058 (I223448,I223615,I223838);
nor I_13059 (I223883,I223581,I223632);
nand I_13060 (I223445,I223883,I223496);
not I_13061 (I223938,I1869);
or I_13062 (I223955,I325212,I325233);
nor I_13063 (I223972,I223955,I325218);
nor I_13064 (I223989,I325212,I325230);
or I_13065 (I224006,I223989,I325221);
nor I_13066 (I224023,I325215,I325215);
nand I_13067 (I224040,I224023,I224006);
not I_13068 (I224057,I224040);
nand I_13069 (I224074,I223972,I224057);
nor I_13070 (I224091,I223972,I224057);
nand I_13071 (I224108,I325224,I325227);
nor I_13072 (I224125,I224108,I325218);
nor I_13073 (I224142,I224108,I224125);
not I_13074 (I224159,I224125);
nor I_13075 (I223930,I224159,I224074);
or I_13076 (I223915,I223972,I224159);
nor I_13077 (I224204,I223972,I224125);
nor I_13078 (I223909,I224108,I224204);
nor I_13079 (I224235,I224142,I224204);
nor I_13080 (I223912,I224057,I224235);
nand I_13081 (I224266,I223972,I224125);
nand I_13082 (I224283,I224040,I224266);
DFFARX1 I_13083 (I224283,I1862,I223938,I223918,);
not I_13084 (I224314,I224108);
nor I_13085 (I223927,I224314,I224159);
nand I_13086 (I223924,I224091,I224314);
nor I_13087 (I224359,I224057,I224108);
nand I_13088 (I223921,I224359,I223972);
not I_13089 (I224414,I1869);
or I_13090 (I224431,I404809,I404812);
nor I_13091 (I224448,I224431,I404809);
nor I_13092 (I224465,I404806,I404824);
or I_13093 (I224482,I224465,I404812);
nor I_13094 (I224499,I404815,I404806);
nand I_13095 (I224516,I224499,I224482);
not I_13096 (I224533,I224516);
nand I_13097 (I224550,I224448,I224533);
nor I_13098 (I224567,I224448,I224533);
nand I_13099 (I224584,I404821,I404818);
nor I_13100 (I224601,I224584,I404815);
nor I_13101 (I224618,I224584,I224601);
not I_13102 (I224635,I224601);
nor I_13103 (I224406,I224635,I224550);
or I_13104 (I224391,I224448,I224635);
nor I_13105 (I224680,I224448,I224601);
nor I_13106 (I224385,I224584,I224680);
nor I_13107 (I224711,I224618,I224680);
nor I_13108 (I224388,I224533,I224711);
nand I_13109 (I224742,I224448,I224601);
nand I_13110 (I224759,I224516,I224742);
DFFARX1 I_13111 (I224759,I1862,I224414,I224394,);
not I_13112 (I224790,I224584);
nor I_13113 (I224403,I224790,I224635);
nand I_13114 (I224400,I224567,I224790);
nor I_13115 (I224835,I224533,I224584);
nand I_13116 (I224397,I224835,I224448);
not I_13117 (I224890,I1869);
or I_13118 (I224907,I336279,I336300);
nor I_13119 (I224924,I224907,I336285);
nor I_13120 (I224941,I336279,I336297);
or I_13121 (I224958,I224941,I336288);
nor I_13122 (I224975,I336282,I336282);
nand I_13123 (I224992,I224975,I224958);
not I_13124 (I225009,I224992);
nand I_13125 (I225026,I224924,I225009);
nor I_13126 (I225043,I224924,I225009);
nand I_13127 (I225060,I336291,I336294);
nor I_13128 (I225077,I225060,I336285);
nor I_13129 (I225094,I225060,I225077);
not I_13130 (I225111,I225077);
nor I_13131 (I224882,I225111,I225026);
or I_13132 (I224867,I224924,I225111);
nor I_13133 (I225156,I224924,I225077);
nor I_13134 (I224861,I225060,I225156);
nor I_13135 (I225187,I225094,I225156);
nor I_13136 (I224864,I225009,I225187);
nand I_13137 (I225218,I224924,I225077);
nand I_13138 (I225235,I224992,I225218);
DFFARX1 I_13139 (I225235,I1862,I224890,I224870,);
not I_13140 (I225266,I225060);
nor I_13141 (I224879,I225266,I225111);
nand I_13142 (I224876,I225043,I225266);
nor I_13143 (I225311,I225009,I225060);
nand I_13144 (I224873,I225311,I224924);
not I_13145 (I225366,I1869);
or I_13146 (I225383,I380057,I380060);
nor I_13147 (I225400,I225383,I380057);
nor I_13148 (I225417,I380054,I380072);
or I_13149 (I225434,I225417,I380060);
nor I_13150 (I225451,I380063,I380054);
nand I_13151 (I225468,I225451,I225434);
not I_13152 (I225485,I225468);
nand I_13153 (I225502,I225400,I225485);
nor I_13154 (I225519,I225400,I225485);
nand I_13155 (I225536,I380069,I380066);
nor I_13156 (I225553,I225536,I380063);
nor I_13157 (I225570,I225536,I225553);
not I_13158 (I225587,I225553);
nor I_13159 (I225358,I225587,I225502);
or I_13160 (I225343,I225400,I225587);
nor I_13161 (I225632,I225400,I225553);
nor I_13162 (I225337,I225536,I225632);
nor I_13163 (I225663,I225570,I225632);
nor I_13164 (I225340,I225485,I225663);
nand I_13165 (I225694,I225400,I225553);
nand I_13166 (I225711,I225468,I225694);
DFFARX1 I_13167 (I225711,I1862,I225366,I225346,);
not I_13168 (I225742,I225536);
nor I_13169 (I225355,I225742,I225587);
nand I_13170 (I225352,I225519,I225742);
nor I_13171 (I225787,I225485,I225536);
nand I_13172 (I225349,I225787,I225400);
not I_13173 (I225842,I1869);
or I_13174 (I225859,I181110,I181095);
nor I_13175 (I225876,I225859,I181089);
nor I_13176 (I225893,I181086,I181107);
or I_13177 (I225910,I225893,I181104);
nor I_13178 (I225927,I181092,I181089);
nand I_13179 (I225944,I225927,I225910);
not I_13180 (I225961,I225944);
nand I_13181 (I225978,I225876,I225961);
nor I_13182 (I225995,I225876,I225961);
nand I_13183 (I226012,I181098,I181101);
nor I_13184 (I226029,I226012,I181086);
nor I_13185 (I226046,I226012,I226029);
not I_13186 (I226063,I226029);
nor I_13187 (I225834,I226063,I225978);
or I_13188 (I225819,I225876,I226063);
nor I_13189 (I226108,I225876,I226029);
nor I_13190 (I225813,I226012,I226108);
nor I_13191 (I226139,I226046,I226108);
nor I_13192 (I225816,I225961,I226139);
nand I_13193 (I226170,I225876,I226029);
nand I_13194 (I226187,I225944,I226170);
DFFARX1 I_13195 (I226187,I1862,I225842,I225822,);
not I_13196 (I226218,I226012);
nor I_13197 (I225831,I226218,I226063);
nand I_13198 (I225828,I225995,I226218);
nor I_13199 (I226263,I225961,I226012);
nand I_13200 (I225825,I226263,I225876);
not I_13201 (I226318,I1869);
or I_13202 (I226335,I109978,I109975);
nor I_13203 (I226352,I226335,I109975);
nor I_13204 (I226369,I109984,I109981);
or I_13205 (I226386,I226369,I109990);
nor I_13206 (I226403,I109993,I109978);
nand I_13207 (I226420,I226403,I226386);
not I_13208 (I226437,I226420);
nand I_13209 (I226454,I226352,I226437);
nor I_13210 (I226471,I226352,I226437);
nand I_13211 (I226488,I109981,I109987);
nor I_13212 (I226505,I226488,I109984);
nor I_13213 (I226522,I226488,I226505);
not I_13214 (I226539,I226505);
nor I_13215 (I226310,I226539,I226454);
or I_13216 (I226295,I226352,I226539);
nor I_13217 (I226584,I226352,I226505);
nor I_13218 (I226289,I226488,I226584);
nor I_13219 (I226615,I226522,I226584);
nor I_13220 (I226292,I226437,I226615);
nand I_13221 (I226646,I226352,I226505);
nand I_13222 (I226663,I226420,I226646);
DFFARX1 I_13223 (I226663,I1862,I226318,I226298,);
not I_13224 (I226694,I226488);
nor I_13225 (I226307,I226694,I226539);
nand I_13226 (I226304,I226471,I226694);
nor I_13227 (I226739,I226437,I226488);
nand I_13228 (I226301,I226739,I226352);
not I_13229 (I226794,I1869);
or I_13230 (I226811,I398179,I398182);
nor I_13231 (I226828,I226811,I398179);
nor I_13232 (I226845,I398176,I398194);
or I_13233 (I226862,I226845,I398182);
nor I_13234 (I226879,I398185,I398176);
nand I_13235 (I226896,I226879,I226862);
not I_13236 (I226913,I226896);
nand I_13237 (I226930,I226828,I226913);
nor I_13238 (I226947,I226828,I226913);
nand I_13239 (I226964,I398191,I398188);
nor I_13240 (I226981,I226964,I398185);
nor I_13241 (I226998,I226964,I226981);
not I_13242 (I227015,I226981);
nor I_13243 (I226786,I227015,I226930);
or I_13244 (I226771,I226828,I227015);
nor I_13245 (I227060,I226828,I226981);
nor I_13246 (I226765,I226964,I227060);
nor I_13247 (I227091,I226998,I227060);
nor I_13248 (I226768,I226913,I227091);
nand I_13249 (I227122,I226828,I226981);
nand I_13250 (I227139,I226896,I227122);
DFFARX1 I_13251 (I227139,I1862,I226794,I226774,);
not I_13252 (I227170,I226964);
nor I_13253 (I226783,I227170,I227015);
nand I_13254 (I226780,I226947,I227170);
nor I_13255 (I227215,I226913,I226964);
nand I_13256 (I226777,I227215,I226828);
not I_13257 (I227270,I1869);
or I_13258 (I227287,I334171,I334192);
nor I_13259 (I227304,I227287,I334177);
nor I_13260 (I227321,I334171,I334189);
or I_13261 (I227338,I227321,I334180);
nor I_13262 (I227355,I334174,I334174);
nand I_13263 (I227372,I227355,I227338);
not I_13264 (I227389,I227372);
nand I_13265 (I227406,I227304,I227389);
nor I_13266 (I227423,I227304,I227389);
nand I_13267 (I227440,I334183,I334186);
nor I_13268 (I227457,I227440,I334177);
nor I_13269 (I227474,I227440,I227457);
not I_13270 (I227491,I227457);
nor I_13271 (I227262,I227491,I227406);
or I_13272 (I227247,I227304,I227491);
nor I_13273 (I227536,I227304,I227457);
nor I_13274 (I227241,I227440,I227536);
nor I_13275 (I227567,I227474,I227536);
nor I_13276 (I227244,I227389,I227567);
nand I_13277 (I227598,I227304,I227457);
nand I_13278 (I227615,I227372,I227598);
DFFARX1 I_13279 (I227615,I1862,I227270,I227250,);
not I_13280 (I227646,I227440);
nor I_13281 (I227259,I227646,I227491);
nand I_13282 (I227256,I227423,I227646);
nor I_13283 (I227691,I227389,I227440);
nand I_13284 (I227253,I227691,I227304);
not I_13285 (I227746,I1869);
or I_13286 (I227763,I12433,I12421);
nor I_13287 (I227780,I227763,I12415);
nor I_13288 (I227797,I12418,I12427);
or I_13289 (I227814,I227797,I12430);
nor I_13290 (I227831,I12412,I12415);
nand I_13291 (I227848,I227831,I227814);
not I_13292 (I227865,I227848);
nand I_13293 (I227882,I227780,I227865);
nor I_13294 (I227899,I227780,I227865);
nand I_13295 (I227916,I12418,I12424);
nor I_13296 (I227933,I227916,I12412);
nor I_13297 (I227950,I227916,I227933);
not I_13298 (I227967,I227933);
nor I_13299 (I227738,I227967,I227882);
or I_13300 (I227723,I227780,I227967);
nor I_13301 (I228012,I227780,I227933);
nor I_13302 (I227717,I227916,I228012);
nor I_13303 (I228043,I227950,I228012);
nor I_13304 (I227720,I227865,I228043);
nand I_13305 (I228074,I227780,I227933);
nand I_13306 (I228091,I227848,I228074);
DFFARX1 I_13307 (I228091,I1862,I227746,I227726,);
not I_13308 (I228122,I227916);
nor I_13309 (I227735,I228122,I227967);
nand I_13310 (I227732,I227899,I228122);
nor I_13311 (I228167,I227865,I227916);
nand I_13312 (I227729,I228167,I227780);
not I_13313 (I228222,I1869);
or I_13314 (I228239,I351035,I351056);
nor I_13315 (I228256,I228239,I351041);
nor I_13316 (I228273,I351035,I351053);
or I_13317 (I228290,I228273,I351044);
nor I_13318 (I228307,I351038,I351038);
nand I_13319 (I228324,I228307,I228290);
not I_13320 (I228341,I228324);
nand I_13321 (I228358,I228256,I228341);
nor I_13322 (I228375,I228256,I228341);
nand I_13323 (I228392,I351047,I351050);
nor I_13324 (I228409,I228392,I351041);
nor I_13325 (I228426,I228392,I228409);
not I_13326 (I228443,I228409);
nor I_13327 (I228214,I228443,I228358);
or I_13328 (I228199,I228256,I228443);
nor I_13329 (I228488,I228256,I228409);
nor I_13330 (I228193,I228392,I228488);
nor I_13331 (I228519,I228426,I228488);
nor I_13332 (I228196,I228341,I228519);
nand I_13333 (I228550,I228256,I228409);
nand I_13334 (I228567,I228324,I228550);
DFFARX1 I_13335 (I228567,I1862,I228222,I228202,);
not I_13336 (I228598,I228392);
nor I_13337 (I228211,I228598,I228443);
nand I_13338 (I228208,I228375,I228598);
nor I_13339 (I228643,I228341,I228392);
nand I_13340 (I228205,I228643,I228256);
not I_13341 (I228698,I1869);
or I_13342 (I228715,I43063,I43072);
nor I_13343 (I228732,I228715,I43087);
nor I_13344 (I228749,I43084,I43066);
or I_13345 (I228766,I228749,I43066);
nor I_13346 (I228783,I43063,I43069);
nand I_13347 (I228800,I228783,I228766);
not I_13348 (I228817,I228800);
nand I_13349 (I228834,I228732,I228817);
nor I_13350 (I228851,I228732,I228817);
nand I_13351 (I228868,I43075,I43078);
nor I_13352 (I228885,I228868,I43081);
nor I_13353 (I228902,I228868,I228885);
not I_13354 (I228919,I228885);
nor I_13355 (I228690,I228919,I228834);
or I_13356 (I228675,I228732,I228919);
nor I_13357 (I228964,I228732,I228885);
nor I_13358 (I228669,I228868,I228964);
nor I_13359 (I228995,I228902,I228964);
nor I_13360 (I228672,I228817,I228995);
nand I_13361 (I229026,I228732,I228885);
nand I_13362 (I229043,I228800,I229026);
DFFARX1 I_13363 (I229043,I1862,I228698,I228678,);
not I_13364 (I229074,I228868);
nor I_13365 (I228687,I229074,I228919);
nand I_13366 (I228684,I228851,I229074);
nor I_13367 (I229119,I228817,I228868);
nand I_13368 (I228681,I229119,I228732);
not I_13369 (I229174,I1869);
or I_13370 (I229191,I359467,I359488);
nor I_13371 (I229208,I229191,I359473);
nor I_13372 (I229225,I359467,I359485);
or I_13373 (I229242,I229225,I359476);
nor I_13374 (I229259,I359470,I359470);
nand I_13375 (I229276,I229259,I229242);
not I_13376 (I229293,I229276);
nand I_13377 (I229310,I229208,I229293);
nor I_13378 (I229327,I229208,I229293);
nand I_13379 (I229344,I359479,I359482);
nor I_13380 (I229361,I229344,I359473);
nor I_13381 (I229378,I229344,I229361);
not I_13382 (I229395,I229361);
nor I_13383 (I229166,I229395,I229310);
or I_13384 (I229151,I229208,I229395);
nor I_13385 (I229440,I229208,I229361);
nor I_13386 (I229145,I229344,I229440);
nor I_13387 (I229471,I229378,I229440);
nor I_13388 (I229148,I229293,I229471);
nand I_13389 (I229502,I229208,I229361);
nand I_13390 (I229519,I229276,I229502);
DFFARX1 I_13391 (I229519,I1862,I229174,I229154,);
not I_13392 (I229550,I229344);
nor I_13393 (I229163,I229550,I229395);
nand I_13394 (I229160,I229327,I229550);
nor I_13395 (I229595,I229293,I229344);
nand I_13396 (I229157,I229595,I229208);
not I_13397 (I229650,I1869);
or I_13398 (I229667,I70093,I70102);
nor I_13399 (I229684,I229667,I70117);
nor I_13400 (I229701,I70114,I70096);
or I_13401 (I229718,I229701,I70096);
nor I_13402 (I229735,I70093,I70099);
nand I_13403 (I229752,I229735,I229718);
not I_13404 (I229769,I229752);
nand I_13405 (I229786,I229684,I229769);
nor I_13406 (I229803,I229684,I229769);
nand I_13407 (I229820,I70105,I70108);
nor I_13408 (I229837,I229820,I70111);
nor I_13409 (I229854,I229820,I229837);
not I_13410 (I229871,I229837);
nor I_13411 (I229642,I229871,I229786);
or I_13412 (I229627,I229684,I229871);
nor I_13413 (I229916,I229684,I229837);
nor I_13414 (I229621,I229820,I229916);
nor I_13415 (I229947,I229854,I229916);
nor I_13416 (I229624,I229769,I229947);
nand I_13417 (I229978,I229684,I229837);
nand I_13418 (I229995,I229752,I229978);
DFFARX1 I_13419 (I229995,I1862,I229650,I229630,);
not I_13420 (I230026,I229820);
nor I_13421 (I229639,I230026,I229871);
nand I_13422 (I229636,I229803,I230026);
nor I_13423 (I230071,I229769,I229820);
nand I_13424 (I229633,I230071,I229684);
not I_13425 (I230126,I1869);
or I_13426 (I230143,I81313,I81322);
nor I_13427 (I230160,I230143,I81337);
nor I_13428 (I230177,I81334,I81316);
or I_13429 (I230194,I230177,I81316);
nor I_13430 (I230211,I81313,I81319);
nand I_13431 (I230228,I230211,I230194);
not I_13432 (I230245,I230228);
nand I_13433 (I230262,I230160,I230245);
nor I_13434 (I230279,I230160,I230245);
nand I_13435 (I230296,I81325,I81328);
nor I_13436 (I230313,I230296,I81331);
nor I_13437 (I230330,I230296,I230313);
not I_13438 (I230347,I230313);
nor I_13439 (I230118,I230347,I230262);
or I_13440 (I230103,I230160,I230347);
nor I_13441 (I230392,I230160,I230313);
nor I_13442 (I230097,I230296,I230392);
nor I_13443 (I230423,I230330,I230392);
nor I_13444 (I230100,I230245,I230423);
nand I_13445 (I230454,I230160,I230313);
nand I_13446 (I230471,I230228,I230454);
DFFARX1 I_13447 (I230471,I1862,I230126,I230106,);
not I_13448 (I230502,I230296);
nor I_13449 (I230115,I230502,I230347);
nand I_13450 (I230112,I230279,I230502);
nor I_13451 (I230547,I230245,I230296);
nand I_13452 (I230109,I230547,I230160);
not I_13453 (I230602,I1869);
or I_13454 (I230619,I372985,I372988);
nor I_13455 (I230636,I230619,I372985);
nor I_13456 (I230653,I372982,I373000);
or I_13457 (I230670,I230653,I372988);
nor I_13458 (I230687,I372991,I372982);
nand I_13459 (I230704,I230687,I230670);
not I_13460 (I230721,I230704);
nand I_13461 (I230738,I230636,I230721);
nor I_13462 (I230755,I230636,I230721);
nand I_13463 (I230772,I372997,I372994);
nor I_13464 (I230789,I230772,I372991);
nor I_13465 (I230806,I230772,I230789);
not I_13466 (I230823,I230789);
nor I_13467 (I230594,I230823,I230738);
or I_13468 (I230579,I230636,I230823);
nor I_13469 (I230868,I230636,I230789);
nor I_13470 (I230573,I230772,I230868);
nor I_13471 (I230899,I230806,I230868);
nor I_13472 (I230576,I230721,I230899);
nand I_13473 (I230930,I230636,I230789);
nand I_13474 (I230947,I230704,I230930);
DFFARX1 I_13475 (I230947,I1862,I230602,I230582,);
not I_13476 (I230978,I230772);
nor I_13477 (I230591,I230978,I230823);
nand I_13478 (I230588,I230755,I230978);
nor I_13479 (I231023,I230721,I230772);
nand I_13480 (I230585,I231023,I230636);
not I_13481 (I231078,I1869);
or I_13482 (I231095,I114466,I114463);
nor I_13483 (I231112,I231095,I114463);
nor I_13484 (I231129,I114472,I114469);
or I_13485 (I231146,I231129,I114478);
nor I_13486 (I231163,I114481,I114466);
nand I_13487 (I231180,I231163,I231146);
not I_13488 (I231197,I231180);
nand I_13489 (I231214,I231112,I231197);
nor I_13490 (I231231,I231112,I231197);
nand I_13491 (I231248,I114469,I114475);
nor I_13492 (I231265,I231248,I114472);
nor I_13493 (I231282,I231248,I231265);
not I_13494 (I231299,I231265);
nor I_13495 (I231070,I231299,I231214);
or I_13496 (I231055,I231112,I231299);
nor I_13497 (I231344,I231112,I231265);
nor I_13498 (I231049,I231248,I231344);
nor I_13499 (I231375,I231282,I231344);
nor I_13500 (I231052,I231197,I231375);
nand I_13501 (I231406,I231112,I231265);
nand I_13502 (I231423,I231180,I231406);
DFFARX1 I_13503 (I231423,I1862,I231078,I231058,);
not I_13504 (I231454,I231248);
nor I_13505 (I231067,I231454,I231299);
nand I_13506 (I231064,I231231,I231454);
nor I_13507 (I231499,I231197,I231248);
nand I_13508 (I231061,I231499,I231112);
not I_13509 (I231554,I1869);
or I_13510 (I231571,I73153,I73162);
nor I_13511 (I231588,I231571,I73177);
nor I_13512 (I231605,I73174,I73156);
or I_13513 (I231622,I231605,I73156);
nor I_13514 (I231639,I73153,I73159);
nand I_13515 (I231656,I231639,I231622);
not I_13516 (I231673,I231656);
nand I_13517 (I231690,I231588,I231673);
nor I_13518 (I231707,I231588,I231673);
nand I_13519 (I231724,I73165,I73168);
nor I_13520 (I231741,I231724,I73171);
nor I_13521 (I231758,I231724,I231741);
not I_13522 (I231775,I231741);
nor I_13523 (I231546,I231775,I231690);
or I_13524 (I231531,I231588,I231775);
nor I_13525 (I231820,I231588,I231741);
nor I_13526 (I231525,I231724,I231820);
nor I_13527 (I231851,I231758,I231820);
nor I_13528 (I231528,I231673,I231851);
nand I_13529 (I231882,I231588,I231741);
nand I_13530 (I231899,I231656,I231882);
DFFARX1 I_13531 (I231899,I1862,I231554,I231534,);
not I_13532 (I231930,I231724);
nor I_13533 (I231543,I231930,I231775);
nand I_13534 (I231540,I231707,I231930);
nor I_13535 (I231975,I231673,I231724);
nand I_13536 (I231537,I231975,I231588);
not I_13537 (I232030,I1869);
or I_13538 (I232047,I324158,I324179);
nor I_13539 (I232064,I232047,I324164);
nor I_13540 (I232081,I324158,I324176);
or I_13541 (I232098,I232081,I324167);
nor I_13542 (I232115,I324161,I324161);
nand I_13543 (I232132,I232115,I232098);
not I_13544 (I232149,I232132);
nand I_13545 (I232166,I232064,I232149);
nor I_13546 (I232183,I232064,I232149);
nand I_13547 (I232200,I324170,I324173);
nor I_13548 (I232217,I232200,I324164);
nor I_13549 (I232234,I232200,I232217);
not I_13550 (I232251,I232217);
nor I_13551 (I232022,I232251,I232166);
or I_13552 (I232007,I232064,I232251);
nor I_13553 (I232296,I232064,I232217);
nor I_13554 (I232001,I232200,I232296);
nor I_13555 (I232327,I232234,I232296);
nor I_13556 (I232004,I232149,I232327);
nand I_13557 (I232358,I232064,I232217);
nand I_13558 (I232375,I232132,I232358);
DFFARX1 I_13559 (I232375,I1862,I232030,I232010,);
not I_13560 (I232406,I232200);
nor I_13561 (I232019,I232406,I232251);
nand I_13562 (I232016,I232183,I232406);
nor I_13563 (I232451,I232149,I232200);
nand I_13564 (I232013,I232451,I232064);
not I_13565 (I232506,I1869);
or I_13566 (I232523,I79783,I79792);
nor I_13567 (I232540,I232523,I79807);
nor I_13568 (I232557,I79804,I79786);
or I_13569 (I232574,I232557,I79786);
nor I_13570 (I232591,I79783,I79789);
nand I_13571 (I232608,I232591,I232574);
not I_13572 (I232625,I232608);
nand I_13573 (I232642,I232540,I232625);
nor I_13574 (I232659,I232540,I232625);
nand I_13575 (I232676,I79795,I79798);
nor I_13576 (I232693,I232676,I79801);
nor I_13577 (I232710,I232676,I232693);
not I_13578 (I232727,I232693);
nor I_13579 (I232498,I232727,I232642);
or I_13580 (I232483,I232540,I232727);
nor I_13581 (I232772,I232540,I232693);
nor I_13582 (I232477,I232676,I232772);
nor I_13583 (I232803,I232710,I232772);
nor I_13584 (I232480,I232625,I232803);
nand I_13585 (I232834,I232540,I232693);
nand I_13586 (I232851,I232608,I232834);
DFFARX1 I_13587 (I232851,I1862,I232506,I232486,);
not I_13588 (I232882,I232676);
nor I_13589 (I232495,I232882,I232727);
nand I_13590 (I232492,I232659,I232882);
nor I_13591 (I232927,I232625,I232676);
nand I_13592 (I232489,I232927,I232540);
not I_13593 (I232982,I1869);
or I_13594 (I232999,I1759,I1719);
nor I_13595 (I233016,I232999,I1087);
nor I_13596 (I233033,I1383,I1071);
or I_13597 (I233050,I233033,I879);
nor I_13598 (I233067,I887,I727);
nand I_13599 (I233084,I233067,I233050);
not I_13600 (I233101,I233084);
nand I_13601 (I233118,I233016,I233101);
nor I_13602 (I233135,I233016,I233101);
nand I_13603 (I233152,I1135,I895);
nor I_13604 (I233169,I233152,I799);
nor I_13605 (I233186,I233152,I233169);
not I_13606 (I233203,I233169);
nor I_13607 (I232974,I233203,I233118);
or I_13608 (I232959,I233016,I233203);
nor I_13609 (I233248,I233016,I233169);
nor I_13610 (I232953,I233152,I233248);
nor I_13611 (I233279,I233186,I233248);
nor I_13612 (I232956,I233101,I233279);
nand I_13613 (I233310,I233016,I233169);
nand I_13614 (I233327,I233084,I233310);
DFFARX1 I_13615 (I233327,I1862,I232982,I232962,);
not I_13616 (I233358,I233152);
nor I_13617 (I232971,I233358,I233203);
nand I_13618 (I232968,I233135,I233358);
nor I_13619 (I233403,I233101,I233152);
nand I_13620 (I232965,I233403,I233016);
not I_13621 (I233458,I1869);
or I_13622 (I233475,I176367,I176352);
nor I_13623 (I233492,I233475,I176346);
nor I_13624 (I233509,I176343,I176364);
or I_13625 (I233526,I233509,I176361);
nor I_13626 (I233543,I176349,I176346);
nand I_13627 (I233560,I233543,I233526);
not I_13628 (I233577,I233560);
nand I_13629 (I233594,I233492,I233577);
nor I_13630 (I233611,I233492,I233577);
nand I_13631 (I233628,I176355,I176358);
nor I_13632 (I233645,I233628,I176343);
nor I_13633 (I233662,I233628,I233645);
not I_13634 (I233679,I233645);
nor I_13635 (I233450,I233679,I233594);
or I_13636 (I233435,I233492,I233679);
nor I_13637 (I233724,I233492,I233645);
nor I_13638 (I233429,I233628,I233724);
nor I_13639 (I233755,I233662,I233724);
nor I_13640 (I233432,I233577,I233755);
nand I_13641 (I233786,I233492,I233645);
nand I_13642 (I233803,I233560,I233786);
DFFARX1 I_13643 (I233803,I1862,I233458,I233438,);
not I_13644 (I233834,I233628);
nor I_13645 (I233447,I233834,I233679);
nand I_13646 (I233444,I233611,I233834);
nor I_13647 (I233879,I233577,I233628);
nand I_13648 (I233441,I233879,I233492);
not I_13649 (I233934,I1869);
or I_13650 (I233951,I164773,I164758);
nor I_13651 (I233968,I233951,I164752);
nor I_13652 (I233985,I164749,I164770);
or I_13653 (I234002,I233985,I164767);
nor I_13654 (I234019,I164755,I164752);
nand I_13655 (I234036,I234019,I234002);
not I_13656 (I234053,I234036);
nand I_13657 (I234070,I233968,I234053);
nor I_13658 (I234087,I233968,I234053);
nand I_13659 (I234104,I164761,I164764);
nor I_13660 (I234121,I234104,I164749);
nor I_13661 (I234138,I234104,I234121);
not I_13662 (I234155,I234121);
nor I_13663 (I233926,I234155,I234070);
or I_13664 (I233911,I233968,I234155);
nor I_13665 (I234200,I233968,I234121);
nor I_13666 (I233905,I234104,I234200);
nor I_13667 (I234231,I234138,I234200);
nor I_13668 (I233908,I234053,I234231);
nand I_13669 (I234262,I233968,I234121);
nand I_13670 (I234279,I234036,I234262);
DFFARX1 I_13671 (I234279,I1862,I233934,I233914,);
not I_13672 (I234310,I234104);
nor I_13673 (I233923,I234310,I234155);
nand I_13674 (I233920,I234087,I234310);
nor I_13675 (I234355,I234053,I234104);
nand I_13676 (I233917,I234355,I233968);
not I_13677 (I234410,I1869);
or I_13678 (I234427,I191650,I191635);
nor I_13679 (I234444,I234427,I191629);
nor I_13680 (I234461,I191626,I191647);
or I_13681 (I234478,I234461,I191644);
nor I_13682 (I234495,I191632,I191629);
nand I_13683 (I234512,I234495,I234478);
not I_13684 (I234529,I234512);
nand I_13685 (I234546,I234444,I234529);
nor I_13686 (I234563,I234444,I234529);
nand I_13687 (I234580,I191638,I191641);
nor I_13688 (I234597,I234580,I191626);
nor I_13689 (I234614,I234580,I234597);
not I_13690 (I234631,I234597);
nor I_13691 (I234402,I234631,I234546);
or I_13692 (I234387,I234444,I234631);
nor I_13693 (I234676,I234444,I234597);
nor I_13694 (I234381,I234580,I234676);
nor I_13695 (I234707,I234614,I234676);
nor I_13696 (I234384,I234529,I234707);
nand I_13697 (I234738,I234444,I234597);
nand I_13698 (I234755,I234512,I234738);
DFFARX1 I_13699 (I234755,I1862,I234410,I234390,);
not I_13700 (I234786,I234580);
nor I_13701 (I234399,I234786,I234631);
nand I_13702 (I234396,I234563,I234786);
nor I_13703 (I234831,I234529,I234580);
nand I_13704 (I234393,I234831,I234444);
not I_13705 (I234886,I1869);
or I_13706 (I234903,I409229,I409232);
nor I_13707 (I234920,I234903,I409229);
nor I_13708 (I234937,I409226,I409244);
or I_13709 (I234954,I234937,I409232);
nor I_13710 (I234971,I409235,I409226);
nand I_13711 (I234988,I234971,I234954);
not I_13712 (I235005,I234988);
nand I_13713 (I235022,I234920,I235005);
nor I_13714 (I235039,I234920,I235005);
nand I_13715 (I235056,I409241,I409238);
nor I_13716 (I235073,I235056,I409235);
nor I_13717 (I235090,I235056,I235073);
not I_13718 (I235107,I235073);
nor I_13719 (I234878,I235107,I235022);
or I_13720 (I234863,I234920,I235107);
nor I_13721 (I235152,I234920,I235073);
nor I_13722 (I234857,I235056,I235152);
nor I_13723 (I235183,I235090,I235152);
nor I_13724 (I234860,I235005,I235183);
nand I_13725 (I235214,I234920,I235073);
nand I_13726 (I235231,I234988,I235214);
DFFARX1 I_13727 (I235231,I1862,I234886,I234866,);
not I_13728 (I235262,I235056);
nor I_13729 (I234875,I235262,I235107);
nand I_13730 (I234872,I235039,I235262);
nor I_13731 (I235307,I235005,I235056);
nand I_13732 (I234869,I235307,I234920);
not I_13733 (I235362,I1869);
or I_13734 (I235379,I112018,I112015);
nor I_13735 (I235396,I235379,I112015);
nor I_13736 (I235413,I112024,I112021);
or I_13737 (I235430,I235413,I112030);
nor I_13738 (I235447,I112033,I112018);
nand I_13739 (I235464,I235447,I235430);
not I_13740 (I235481,I235464);
nand I_13741 (I235498,I235396,I235481);
nor I_13742 (I235515,I235396,I235481);
nand I_13743 (I235532,I112021,I112027);
nor I_13744 (I235549,I235532,I112024);
nor I_13745 (I235566,I235532,I235549);
not I_13746 (I235583,I235549);
nor I_13747 (I235354,I235583,I235498);
or I_13748 (I235339,I235396,I235583);
nor I_13749 (I235628,I235396,I235549);
nor I_13750 (I235333,I235532,I235628);
nor I_13751 (I235659,I235566,I235628);
nor I_13752 (I235336,I235481,I235659);
nand I_13753 (I235690,I235396,I235549);
nand I_13754 (I235707,I235464,I235690);
DFFARX1 I_13755 (I235707,I1862,I235362,I235342,);
not I_13756 (I235738,I235532);
nor I_13757 (I235351,I235738,I235583);
nand I_13758 (I235348,I235515,I235738);
nor I_13759 (I235783,I235481,I235532);
nand I_13760 (I235345,I235783,I235396);
not I_13761 (I235838,I1869);
or I_13762 (I235855,I144220,I144205);
nor I_13763 (I235872,I235855,I144199);
nor I_13764 (I235889,I144196,I144217);
or I_13765 (I235906,I235889,I144214);
nor I_13766 (I235923,I144202,I144199);
nand I_13767 (I235940,I235923,I235906);
not I_13768 (I235957,I235940);
nand I_13769 (I235974,I235872,I235957);
nor I_13770 (I235991,I235872,I235957);
nand I_13771 (I236008,I144208,I144211);
nor I_13772 (I236025,I236008,I144196);
nor I_13773 (I236042,I236008,I236025);
not I_13774 (I236059,I236025);
nor I_13775 (I235830,I236059,I235974);
or I_13776 (I235815,I235872,I236059);
nor I_13777 (I236104,I235872,I236025);
nor I_13778 (I235809,I236008,I236104);
nor I_13779 (I236135,I236042,I236104);
nor I_13780 (I235812,I235957,I236135);
nand I_13781 (I236166,I235872,I236025);
nand I_13782 (I236183,I235940,I236166);
DFFARX1 I_13783 (I236183,I1862,I235838,I235818,);
not I_13784 (I236214,I236008);
nor I_13785 (I235827,I236214,I236059);
nand I_13786 (I235824,I235991,I236214);
nor I_13787 (I236259,I235957,I236008);
nand I_13788 (I235821,I236259,I235872);
not I_13789 (I236314,I1869);
or I_13790 (I236331,I35923,I35932);
nor I_13791 (I236348,I236331,I35947);
nor I_13792 (I236365,I35944,I35926);
or I_13793 (I236382,I236365,I35926);
nor I_13794 (I236399,I35923,I35929);
nand I_13795 (I236416,I236399,I236382);
not I_13796 (I236433,I236416);
nand I_13797 (I236450,I236348,I236433);
nor I_13798 (I236467,I236348,I236433);
nand I_13799 (I236484,I35935,I35938);
nor I_13800 (I236501,I236484,I35941);
nor I_13801 (I236518,I236484,I236501);
not I_13802 (I236535,I236501);
nor I_13803 (I236306,I236535,I236450);
or I_13804 (I236291,I236348,I236535);
nor I_13805 (I236580,I236348,I236501);
nor I_13806 (I236285,I236484,I236580);
nor I_13807 (I236611,I236518,I236580);
nor I_13808 (I236288,I236433,I236611);
nand I_13809 (I236642,I236348,I236501);
nand I_13810 (I236659,I236416,I236642);
DFFARX1 I_13811 (I236659,I1862,I236314,I236294,);
not I_13812 (I236690,I236484);
nor I_13813 (I236303,I236690,I236535);
nand I_13814 (I236300,I236467,I236690);
nor I_13815 (I236735,I236433,I236484);
nand I_13816 (I236297,I236735,I236348);
not I_13817 (I236790,I1869);
or I_13818 (I236807,I90493,I90502);
nor I_13819 (I236824,I236807,I90517);
nor I_13820 (I236841,I90514,I90496);
or I_13821 (I236858,I236841,I90496);
nor I_13822 (I236875,I90493,I90499);
nand I_13823 (I236892,I236875,I236858);
not I_13824 (I236909,I236892);
nand I_13825 (I236926,I236824,I236909);
nor I_13826 (I236943,I236824,I236909);
nand I_13827 (I236960,I90505,I90508);
nor I_13828 (I236977,I236960,I90511);
nor I_13829 (I236994,I236960,I236977);
not I_13830 (I237011,I236977);
nor I_13831 (I236782,I237011,I236926);
or I_13832 (I236767,I236824,I237011);
nor I_13833 (I237056,I236824,I236977);
nor I_13834 (I236761,I236960,I237056);
nor I_13835 (I237087,I236994,I237056);
nor I_13836 (I236764,I236909,I237087);
nand I_13837 (I237118,I236824,I236977);
nand I_13838 (I237135,I236892,I237118);
DFFARX1 I_13839 (I237135,I1862,I236790,I236770,);
not I_13840 (I237166,I236960);
nor I_13841 (I236779,I237166,I237011);
nand I_13842 (I236776,I236943,I237166);
nor I_13843 (I237211,I236909,I236960);
nand I_13844 (I236773,I237211,I236824);
not I_13845 (I237266,I1869);
or I_13846 (I237283,I4528,I4516);
nor I_13847 (I237300,I237283,I4510);
nor I_13848 (I237317,I4513,I4522);
or I_13849 (I237334,I237317,I4525);
nor I_13850 (I237351,I4507,I4510);
nand I_13851 (I237368,I237351,I237334);
not I_13852 (I237385,I237368);
nand I_13853 (I237402,I237300,I237385);
nor I_13854 (I237419,I237300,I237385);
nand I_13855 (I237436,I4513,I4519);
nor I_13856 (I237453,I237436,I4507);
nor I_13857 (I237470,I237436,I237453);
not I_13858 (I237487,I237453);
nor I_13859 (I237258,I237487,I237402);
or I_13860 (I237243,I237300,I237487);
nor I_13861 (I237532,I237300,I237453);
nor I_13862 (I237237,I237436,I237532);
nor I_13863 (I237563,I237470,I237532);
nor I_13864 (I237240,I237385,I237563);
nand I_13865 (I237594,I237300,I237453);
nand I_13866 (I237611,I237368,I237594);
DFFARX1 I_13867 (I237611,I1862,I237266,I237246,);
not I_13868 (I237642,I237436);
nor I_13869 (I237255,I237642,I237487);
nand I_13870 (I237252,I237419,I237642);
nor I_13871 (I237687,I237385,I237436);
nand I_13872 (I237249,I237687,I237300);
not I_13873 (I237742,I1869);
or I_13874 (I237759,I130518,I130503);
nor I_13875 (I237776,I237759,I130497);
nor I_13876 (I237793,I130494,I130515);
or I_13877 (I237810,I237793,I130512);
nor I_13878 (I237827,I130500,I130497);
nand I_13879 (I237844,I237827,I237810);
not I_13880 (I237861,I237844);
nand I_13881 (I237878,I237776,I237861);
nor I_13882 (I237895,I237776,I237861);
nand I_13883 (I237912,I130506,I130509);
nor I_13884 (I237929,I237912,I130494);
nor I_13885 (I237946,I237912,I237929);
not I_13886 (I237963,I237929);
nor I_13887 (I237734,I237963,I237878);
or I_13888 (I237719,I237776,I237963);
nor I_13889 (I238008,I237776,I237929);
nor I_13890 (I237713,I237912,I238008);
nor I_13891 (I238039,I237946,I238008);
nor I_13892 (I237716,I237861,I238039);
nand I_13893 (I238070,I237776,I237929);
nand I_13894 (I238087,I237844,I238070);
DFFARX1 I_13895 (I238087,I1862,I237742,I237722,);
not I_13896 (I238118,I237912);
nor I_13897 (I237731,I238118,I237963);
nand I_13898 (I237728,I237895,I238118);
nor I_13899 (I238163,I237861,I237912);
nand I_13900 (I237725,I238163,I237776);
not I_13901 (I238218,I1869);
or I_13902 (I238235,I7690,I7678);
nor I_13903 (I238252,I238235,I7672);
nor I_13904 (I238269,I7675,I7684);
or I_13905 (I238286,I238269,I7687);
nor I_13906 (I238303,I7669,I7672);
nand I_13907 (I238320,I238303,I238286);
not I_13908 (I238337,I238320);
nand I_13909 (I238354,I238252,I238337);
nor I_13910 (I238371,I238252,I238337);
nand I_13911 (I238388,I7675,I7681);
nor I_13912 (I238405,I238388,I7669);
nor I_13913 (I238422,I238388,I238405);
not I_13914 (I238439,I238405);
nor I_13915 (I238210,I238439,I238354);
or I_13916 (I238195,I238252,I238439);
nor I_13917 (I238484,I238252,I238405);
nor I_13918 (I238189,I238388,I238484);
nor I_13919 (I238515,I238422,I238484);
nor I_13920 (I238192,I238337,I238515);
nand I_13921 (I238546,I238252,I238405);
nand I_13922 (I238563,I238320,I238546);
DFFARX1 I_13923 (I238563,I1862,I238218,I238198,);
not I_13924 (I238594,I238388);
nor I_13925 (I238207,I238594,I238439);
nand I_13926 (I238204,I238371,I238594);
nor I_13927 (I238639,I238337,I238388);
nand I_13928 (I238201,I238639,I238252);
not I_13929 (I238694,I1869);
or I_13930 (I238711,I63463,I63472);
nor I_13931 (I238728,I238711,I63487);
nor I_13932 (I238745,I63484,I63466);
or I_13933 (I238762,I238745,I63466);
nor I_13934 (I238779,I63463,I63469);
nand I_13935 (I238796,I238779,I238762);
not I_13936 (I238813,I238796);
nand I_13937 (I238830,I238728,I238813);
nor I_13938 (I238847,I238728,I238813);
nand I_13939 (I238864,I63475,I63478);
nor I_13940 (I238881,I238864,I63481);
nor I_13941 (I238898,I238864,I238881);
not I_13942 (I238915,I238881);
nor I_13943 (I238686,I238915,I238830);
or I_13944 (I238671,I238728,I238915);
nor I_13945 (I238960,I238728,I238881);
nor I_13946 (I238665,I238864,I238960);
nor I_13947 (I238991,I238898,I238960);
nor I_13948 (I238668,I238813,I238991);
nand I_13949 (I239022,I238728,I238881);
nand I_13950 (I239039,I238796,I239022);
DFFARX1 I_13951 (I239039,I1862,I238694,I238674,);
not I_13952 (I239070,I238864);
nor I_13953 (I238683,I239070,I238915);
nand I_13954 (I238680,I238847,I239070);
nor I_13955 (I239115,I238813,I238864);
nand I_13956 (I238677,I239115,I238728);
not I_13957 (I239170,I1869);
or I_13958 (I239187,I82843,I82852);
nor I_13959 (I239204,I239187,I82867);
nor I_13960 (I239221,I82864,I82846);
or I_13961 (I239238,I239221,I82846);
nor I_13962 (I239255,I82843,I82849);
nand I_13963 (I239272,I239255,I239238);
not I_13964 (I239289,I239272);
nand I_13965 (I239306,I239204,I239289);
nor I_13966 (I239323,I239204,I239289);
nand I_13967 (I239340,I82855,I82858);
nor I_13968 (I239357,I239340,I82861);
nor I_13969 (I239374,I239340,I239357);
not I_13970 (I239391,I239357);
nor I_13971 (I239162,I239391,I239306);
or I_13972 (I239147,I239204,I239391);
nor I_13973 (I239436,I239204,I239357);
nor I_13974 (I239141,I239340,I239436);
nor I_13975 (I239467,I239374,I239436);
nor I_13976 (I239144,I239289,I239467);
nand I_13977 (I239498,I239204,I239357);
nand I_13978 (I239515,I239272,I239498);
DFFARX1 I_13979 (I239515,I1862,I239170,I239150,);
not I_13980 (I239546,I239340);
nor I_13981 (I239159,I239546,I239391);
nand I_13982 (I239156,I239323,I239546);
nor I_13983 (I239591,I239289,I239340);
nand I_13984 (I239153,I239591,I239204);
not I_13985 (I239646,I1869);
or I_13986 (I239663,I51733,I51742);
nor I_13987 (I239680,I239663,I51757);
nor I_13988 (I239697,I51754,I51736);
or I_13989 (I239714,I239697,I51736);
nor I_13990 (I239731,I51733,I51739);
nand I_13991 (I239748,I239731,I239714);
not I_13992 (I239765,I239748);
nand I_13993 (I239782,I239680,I239765);
nor I_13994 (I239799,I239680,I239765);
nand I_13995 (I239816,I51745,I51748);
nor I_13996 (I239833,I239816,I51751);
nor I_13997 (I239850,I239816,I239833);
not I_13998 (I239867,I239833);
nor I_13999 (I239638,I239867,I239782);
or I_14000 (I239623,I239680,I239867);
nor I_14001 (I239912,I239680,I239833);
nor I_14002 (I239617,I239816,I239912);
nor I_14003 (I239943,I239850,I239912);
nor I_14004 (I239620,I239765,I239943);
nand I_14005 (I239974,I239680,I239833);
nand I_14006 (I239991,I239748,I239974);
DFFARX1 I_14007 (I239991,I1862,I239646,I239626,);
not I_14008 (I240022,I239816);
nor I_14009 (I239635,I240022,I239867);
nand I_14010 (I239632,I239799,I240022);
nor I_14011 (I240067,I239765,I239816);
nand I_14012 (I239629,I240067,I239680);
not I_14013 (I240122,I1869);
or I_14014 (I240139,I173205,I173190);
nor I_14015 (I240156,I240139,I173184);
nor I_14016 (I240173,I173181,I173202);
or I_14017 (I240190,I240173,I173199);
nor I_14018 (I240207,I173187,I173184);
nand I_14019 (I240224,I240207,I240190);
not I_14020 (I240241,I240224);
nand I_14021 (I240258,I240156,I240241);
nor I_14022 (I240275,I240156,I240241);
nand I_14023 (I240292,I173193,I173196);
nor I_14024 (I240309,I240292,I173181);
nor I_14025 (I240326,I240292,I240309);
not I_14026 (I240343,I240309);
nor I_14027 (I240114,I240343,I240258);
or I_14028 (I240099,I240156,I240343);
nor I_14029 (I240388,I240156,I240309);
nor I_14030 (I240093,I240292,I240388);
nor I_14031 (I240419,I240326,I240388);
nor I_14032 (I240096,I240241,I240419);
nand I_14033 (I240450,I240156,I240309);
nand I_14034 (I240467,I240224,I240450);
DFFARX1 I_14035 (I240467,I1862,I240122,I240102,);
not I_14036 (I240498,I240292);
nor I_14037 (I240111,I240498,I240343);
nand I_14038 (I240108,I240275,I240498);
nor I_14039 (I240543,I240241,I240292);
nand I_14040 (I240105,I240543,I240156);
not I_14041 (I240598,I1869);
or I_14042 (I240615,I386245,I386248);
nor I_14043 (I240632,I240615,I386245);
nor I_14044 (I240649,I386242,I386260);
or I_14045 (I240666,I240649,I386248);
nor I_14046 (I240683,I386251,I386242);
nand I_14047 (I240700,I240683,I240666);
not I_14048 (I240717,I240700);
nand I_14049 (I240734,I240632,I240717);
nor I_14050 (I240751,I240632,I240717);
nand I_14051 (I240768,I386257,I386254);
nor I_14052 (I240785,I240768,I386251);
nor I_14053 (I240802,I240768,I240785);
not I_14054 (I240819,I240785);
nor I_14055 (I240590,I240819,I240734);
or I_14056 (I240575,I240632,I240819);
nor I_14057 (I240864,I240632,I240785);
nor I_14058 (I240569,I240768,I240864);
nor I_14059 (I240895,I240802,I240864);
nor I_14060 (I240572,I240717,I240895);
nand I_14061 (I240926,I240632,I240785);
nand I_14062 (I240943,I240700,I240926);
DFFARX1 I_14063 (I240943,I1862,I240598,I240578,);
not I_14064 (I240974,I240768);
nor I_14065 (I240587,I240974,I240819);
nand I_14066 (I240584,I240751,I240974);
nor I_14067 (I241019,I240717,I240768);
nand I_14068 (I240581,I241019,I240632);
not I_14069 (I241074,I1869);
or I_14070 (I241091,I381825,I381828);
nor I_14071 (I241108,I241091,I381825);
nor I_14072 (I241125,I381822,I381840);
or I_14073 (I241142,I241125,I381828);
nor I_14074 (I241159,I381831,I381822);
nand I_14075 (I241176,I241159,I241142);
not I_14076 (I241193,I241176);
nand I_14077 (I241210,I241108,I241193);
nor I_14078 (I241227,I241108,I241193);
nand I_14079 (I241244,I381837,I381834);
nor I_14080 (I241261,I241244,I381831);
nor I_14081 (I241278,I241244,I241261);
not I_14082 (I241295,I241261);
nor I_14083 (I241066,I241295,I241210);
or I_14084 (I241051,I241108,I241295);
nor I_14085 (I241340,I241108,I241261);
nor I_14086 (I241045,I241244,I241340);
nor I_14087 (I241371,I241278,I241340);
nor I_14088 (I241048,I241193,I241371);
nand I_14089 (I241402,I241108,I241261);
nand I_14090 (I241419,I241176,I241402);
DFFARX1 I_14091 (I241419,I1862,I241074,I241054,);
not I_14092 (I241450,I241244);
nor I_14093 (I241063,I241450,I241295);
nand I_14094 (I241060,I241227,I241450);
nor I_14095 (I241495,I241193,I241244);
nand I_14096 (I241057,I241495,I241108);
not I_14097 (I241550,I1869);
or I_14098 (I241567,I391549,I391552);
nor I_14099 (I241584,I241567,I391549);
nor I_14100 (I241601,I391546,I391564);
or I_14101 (I241618,I241601,I391552);
nor I_14102 (I241635,I391555,I391546);
nand I_14103 (I241652,I241635,I241618);
not I_14104 (I241669,I241652);
nand I_14105 (I241686,I241584,I241669);
nor I_14106 (I241703,I241584,I241669);
nand I_14107 (I241720,I391561,I391558);
nor I_14108 (I241737,I241720,I391555);
nor I_14109 (I241754,I241720,I241737);
not I_14110 (I241771,I241737);
nor I_14111 (I241542,I241771,I241686);
or I_14112 (I241527,I241584,I241771);
nor I_14113 (I241816,I241584,I241737);
nor I_14114 (I241521,I241720,I241816);
nor I_14115 (I241847,I241754,I241816);
nor I_14116 (I241524,I241669,I241847);
nand I_14117 (I241878,I241584,I241737);
nand I_14118 (I241895,I241652,I241878);
DFFARX1 I_14119 (I241895,I1862,I241550,I241530,);
not I_14120 (I241926,I241720);
nor I_14121 (I241539,I241926,I241771);
nand I_14122 (I241536,I241703,I241926);
nor I_14123 (I241971,I241669,I241720);
nand I_14124 (I241533,I241971,I241584);
not I_14125 (I242026,I1869);
or I_14126 (I242043,I107938,I107935);
nor I_14127 (I242060,I242043,I107935);
nor I_14128 (I242077,I107944,I107941);
or I_14129 (I242094,I242077,I107950);
nor I_14130 (I242111,I107953,I107938);
nand I_14131 (I242128,I242111,I242094);
not I_14132 (I242145,I242128);
nand I_14133 (I242162,I242060,I242145);
nor I_14134 (I242179,I242060,I242145);
nand I_14135 (I242196,I107941,I107947);
nor I_14136 (I242213,I242196,I107944);
nor I_14137 (I242230,I242196,I242213);
not I_14138 (I242247,I242213);
nor I_14139 (I242018,I242247,I242162);
or I_14140 (I242003,I242060,I242247);
nor I_14141 (I242292,I242060,I242213);
nor I_14142 (I241997,I242196,I242292);
nor I_14143 (I242323,I242230,I242292);
nor I_14144 (I242000,I242145,I242323);
nand I_14145 (I242354,I242060,I242213);
nand I_14146 (I242371,I242128,I242354);
DFFARX1 I_14147 (I242371,I1862,I242026,I242006,);
not I_14148 (I242402,I242196);
nor I_14149 (I242015,I242402,I242247);
nand I_14150 (I242012,I242179,I242402);
nor I_14151 (I242447,I242145,I242196);
nand I_14152 (I242009,I242447,I242060);
not I_14153 (I242502,I1869);
or I_14154 (I242519,I156341,I156326);
nor I_14155 (I242536,I242519,I156320);
nor I_14156 (I242553,I156317,I156338);
or I_14157 (I242570,I242553,I156335);
nor I_14158 (I242587,I156323,I156320);
nand I_14159 (I242604,I242587,I242570);
not I_14160 (I242621,I242604);
nand I_14161 (I242638,I242536,I242621);
nor I_14162 (I242655,I242536,I242621);
nand I_14163 (I242672,I156329,I156332);
nor I_14164 (I242689,I242672,I156317);
nor I_14165 (I242706,I242672,I242689);
not I_14166 (I242723,I242689);
nor I_14167 (I242494,I242723,I242638);
or I_14168 (I242479,I242536,I242723);
nor I_14169 (I242768,I242536,I242689);
nor I_14170 (I242473,I242672,I242768);
nor I_14171 (I242799,I242706,I242768);
nor I_14172 (I242476,I242621,I242799);
nand I_14173 (I242830,I242536,I242689);
nand I_14174 (I242847,I242604,I242830);
DFFARX1 I_14175 (I242847,I1862,I242502,I242482,);
not I_14176 (I242878,I242672);
nor I_14177 (I242491,I242878,I242723);
nand I_14178 (I242488,I242655,I242878);
nor I_14179 (I242923,I242621,I242672);
nand I_14180 (I242485,I242923,I242536);
not I_14181 (I242978,I1869);
or I_14182 (I242995,I292014,I292011);
nor I_14183 (I243012,I242995,I292020);
nor I_14184 (I243029,I292032,I292017);
or I_14185 (I243046,I243029,I292011);
nor I_14186 (I243063,I292023,I292014);
nand I_14187 (I243080,I243063,I243046);
not I_14188 (I243097,I243080);
nand I_14189 (I243114,I243012,I243097);
nor I_14190 (I243131,I243012,I243097);
nand I_14191 (I243148,I292017,I292029);
nor I_14192 (I243165,I243148,I292026);
nor I_14193 (I243182,I243148,I243165);
not I_14194 (I243199,I243165);
nor I_14195 (I242970,I243199,I243114);
or I_14196 (I242955,I243012,I243199);
nor I_14197 (I243244,I243012,I243165);
nor I_14198 (I242949,I243148,I243244);
nor I_14199 (I243275,I243182,I243244);
nor I_14200 (I242952,I243097,I243275);
nand I_14201 (I243306,I243012,I243165);
nand I_14202 (I243323,I243080,I243306);
DFFARX1 I_14203 (I243323,I1862,I242978,I242958,);
not I_14204 (I243354,I243148);
nor I_14205 (I242967,I243354,I243199);
nand I_14206 (I242964,I243131,I243354);
nor I_14207 (I243399,I243097,I243148);
nand I_14208 (I242961,I243399,I243012);
not I_14209 (I243454,I1869);
or I_14210 (I243471,I57343,I57352);
nor I_14211 (I243488,I243471,I57367);
nor I_14212 (I243505,I57364,I57346);
or I_14213 (I243522,I243505,I57346);
nor I_14214 (I243539,I57343,I57349);
nand I_14215 (I243556,I243539,I243522);
not I_14216 (I243573,I243556);
nand I_14217 (I243590,I243488,I243573);
nor I_14218 (I243607,I243488,I243573);
nand I_14219 (I243624,I57355,I57358);
nor I_14220 (I243641,I243624,I57361);
nor I_14221 (I243658,I243624,I243641);
not I_14222 (I243675,I243641);
nor I_14223 (I243446,I243675,I243590);
or I_14224 (I243431,I243488,I243675);
nor I_14225 (I243720,I243488,I243641);
nor I_14226 (I243425,I243624,I243720);
nor I_14227 (I243751,I243658,I243720);
nor I_14228 (I243428,I243573,I243751);
nand I_14229 (I243782,I243488,I243641);
nand I_14230 (I243799,I243556,I243782);
DFFARX1 I_14231 (I243799,I1862,I243454,I243434,);
not I_14232 (I243830,I243624);
nor I_14233 (I243443,I243830,I243675);
nand I_14234 (I243440,I243607,I243830);
nor I_14235 (I243875,I243573,I243624);
nand I_14236 (I243437,I243875,I243488);
not I_14237 (I243930,I1869);
or I_14238 (I243947,I335225,I335246);
nor I_14239 (I243964,I243947,I335231);
nor I_14240 (I243981,I335225,I335243);
or I_14241 (I243998,I243981,I335234);
nor I_14242 (I244015,I335228,I335228);
nand I_14243 (I244032,I244015,I243998);
not I_14244 (I244049,I244032);
nand I_14245 (I244066,I243964,I244049);
nor I_14246 (I244083,I243964,I244049);
nand I_14247 (I244100,I335237,I335240);
nor I_14248 (I244117,I244100,I335231);
nor I_14249 (I244134,I244100,I244117);
not I_14250 (I244151,I244117);
nor I_14251 (I243922,I244151,I244066);
or I_14252 (I243907,I243964,I244151);
nor I_14253 (I244196,I243964,I244117);
nor I_14254 (I243901,I244100,I244196);
nor I_14255 (I244227,I244134,I244196);
nor I_14256 (I243904,I244049,I244227);
nand I_14257 (I244258,I243964,I244117);
nand I_14258 (I244275,I244032,I244258);
DFFARX1 I_14259 (I244275,I1862,I243930,I243910,);
not I_14260 (I244306,I244100);
nor I_14261 (I243919,I244306,I244151);
nand I_14262 (I243916,I244083,I244306);
nor I_14263 (I244351,I244049,I244100);
nand I_14264 (I243913,I244351,I243964);
not I_14265 (I244406,I1869);
or I_14266 (I244423,I108346,I108343);
nor I_14267 (I244440,I244423,I108343);
nor I_14268 (I244457,I108352,I108349);
or I_14269 (I244474,I244457,I108358);
nor I_14270 (I244491,I108361,I108346);
nand I_14271 (I244508,I244491,I244474);
not I_14272 (I244525,I244508);
nand I_14273 (I244542,I244440,I244525);
nor I_14274 (I244559,I244440,I244525);
nand I_14275 (I244576,I108349,I108355);
nor I_14276 (I244593,I244576,I108352);
nor I_14277 (I244610,I244576,I244593);
not I_14278 (I244627,I244593);
nor I_14279 (I244398,I244627,I244542);
or I_14280 (I244383,I244440,I244627);
nor I_14281 (I244672,I244440,I244593);
nor I_14282 (I244377,I244576,I244672);
nor I_14283 (I244703,I244610,I244672);
nor I_14284 (I244380,I244525,I244703);
nand I_14285 (I244734,I244440,I244593);
nand I_14286 (I244751,I244508,I244734);
DFFARX1 I_14287 (I244751,I1862,I244406,I244386,);
not I_14288 (I244782,I244576);
nor I_14289 (I244395,I244782,I244627);
nand I_14290 (I244392,I244559,I244782);
nor I_14291 (I244827,I244525,I244576);
nand I_14292 (I244389,I244827,I244440);
not I_14293 (I244882,I1869);
or I_14294 (I244899,I62953,I62962);
nor I_14295 (I244916,I244899,I62977);
nor I_14296 (I244933,I62974,I62956);
or I_14297 (I244950,I244933,I62956);
nor I_14298 (I244967,I62953,I62959);
nand I_14299 (I244984,I244967,I244950);
not I_14300 (I245001,I244984);
nand I_14301 (I245018,I244916,I245001);
nor I_14302 (I245035,I244916,I245001);
nand I_14303 (I245052,I62965,I62968);
nor I_14304 (I245069,I245052,I62971);
nor I_14305 (I245086,I245052,I245069);
not I_14306 (I245103,I245069);
nor I_14307 (I244874,I245103,I245018);
or I_14308 (I244859,I244916,I245103);
nor I_14309 (I245148,I244916,I245069);
nor I_14310 (I244853,I245052,I245148);
nor I_14311 (I245179,I245086,I245148);
nor I_14312 (I244856,I245001,I245179);
nand I_14313 (I245210,I244916,I245069);
nand I_14314 (I245227,I244984,I245210);
DFFARX1 I_14315 (I245227,I1862,I244882,I244862,);
not I_14316 (I245258,I245052);
nor I_14317 (I244871,I245258,I245103);
nand I_14318 (I244868,I245035,I245258);
nor I_14319 (I245303,I245001,I245052);
nand I_14320 (I244865,I245303,I244916);
not I_14321 (I245358,I1869);
or I_14322 (I245375,I70603,I70612);
nor I_14323 (I245392,I245375,I70627);
nor I_14324 (I245409,I70624,I70606);
or I_14325 (I245426,I245409,I70606);
nor I_14326 (I245443,I70603,I70609);
nand I_14327 (I245460,I245443,I245426);
not I_14328 (I245477,I245460);
nand I_14329 (I245494,I245392,I245477);
nor I_14330 (I245511,I245392,I245477);
nand I_14331 (I245528,I70615,I70618);
nor I_14332 (I245545,I245528,I70621);
nor I_14333 (I245562,I245528,I245545);
not I_14334 (I245579,I245545);
nor I_14335 (I245350,I245579,I245494);
or I_14336 (I245335,I245392,I245579);
nor I_14337 (I245624,I245392,I245545);
nor I_14338 (I245329,I245528,I245624);
nor I_14339 (I245655,I245562,I245624);
nor I_14340 (I245332,I245477,I245655);
nand I_14341 (I245686,I245392,I245545);
nand I_14342 (I245703,I245460,I245686);
DFFARX1 I_14343 (I245703,I1862,I245358,I245338,);
not I_14344 (I245734,I245528);
nor I_14345 (I245347,I245734,I245579);
nand I_14346 (I245344,I245511,I245734);
nor I_14347 (I245779,I245477,I245528);
nand I_14348 (I245341,I245779,I245392);
not I_14349 (I245834,I1869);
or I_14350 (I245851,I8744,I8732);
nor I_14351 (I245868,I245851,I8726);
nor I_14352 (I245885,I8729,I8738);
or I_14353 (I245902,I245885,I8741);
nor I_14354 (I245919,I8723,I8726);
nand I_14355 (I245936,I245919,I245902);
not I_14356 (I245953,I245936);
nand I_14357 (I245970,I245868,I245953);
nor I_14358 (I245987,I245868,I245953);
nand I_14359 (I246004,I8729,I8735);
nor I_14360 (I246021,I246004,I8723);
nor I_14361 (I246038,I246004,I246021);
not I_14362 (I246055,I246021);
nor I_14363 (I245826,I246055,I245970);
or I_14364 (I245811,I245868,I246055);
nor I_14365 (I246100,I245868,I246021);
nor I_14366 (I245805,I246004,I246100);
nor I_14367 (I246131,I246038,I246100);
nor I_14368 (I245808,I245953,I246131);
nand I_14369 (I246162,I245868,I246021);
nand I_14370 (I246179,I245936,I246162);
DFFARX1 I_14371 (I246179,I1862,I245834,I245814,);
not I_14372 (I246210,I246004);
nor I_14373 (I245823,I246210,I246055);
nand I_14374 (I245820,I245987,I246210);
nor I_14375 (I246255,I245953,I246004);
nand I_14376 (I245817,I246255,I245868);
not I_14377 (I246310,I1869);
or I_14378 (I246327,I197974,I197959);
nor I_14379 (I246344,I246327,I197953);
nor I_14380 (I246361,I197950,I197971);
or I_14381 (I246378,I246361,I197968);
nor I_14382 (I246395,I197956,I197953);
nand I_14383 (I246412,I246395,I246378);
not I_14384 (I246429,I246412);
nand I_14385 (I246446,I246344,I246429);
nor I_14386 (I246463,I246344,I246429);
nand I_14387 (I246480,I197962,I197965);
nor I_14388 (I246497,I246480,I197950);
nor I_14389 (I246514,I246480,I246497);
not I_14390 (I246531,I246497);
nor I_14391 (I246302,I246531,I246446);
or I_14392 (I246287,I246344,I246531);
nor I_14393 (I246576,I246344,I246497);
nor I_14394 (I246281,I246480,I246576);
nor I_14395 (I246607,I246514,I246576);
nor I_14396 (I246284,I246429,I246607);
nand I_14397 (I246638,I246344,I246497);
nand I_14398 (I246655,I246412,I246638);
DFFARX1 I_14399 (I246655,I1862,I246310,I246290,);
not I_14400 (I246686,I246480);
nor I_14401 (I246299,I246686,I246531);
nand I_14402 (I246296,I246463,I246686);
nor I_14403 (I246731,I246429,I246480);
nand I_14404 (I246293,I246731,I246344);
not I_14405 (I246786,I1869);
or I_14406 (I246803,I149490,I149475);
nor I_14407 (I246820,I246803,I149469);
nor I_14408 (I246837,I149466,I149487);
or I_14409 (I246854,I246837,I149484);
nor I_14410 (I246871,I149472,I149469);
nand I_14411 (I246888,I246871,I246854);
not I_14412 (I246905,I246888);
nand I_14413 (I246922,I246820,I246905);
nor I_14414 (I246939,I246820,I246905);
nand I_14415 (I246956,I149478,I149481);
nor I_14416 (I246973,I246956,I149466);
nor I_14417 (I246990,I246956,I246973);
not I_14418 (I247007,I246973);
nor I_14419 (I246778,I247007,I246922);
or I_14420 (I246763,I246820,I247007);
nor I_14421 (I247052,I246820,I246973);
nor I_14422 (I246757,I246956,I247052);
nor I_14423 (I247083,I246990,I247052);
nor I_14424 (I246760,I246905,I247083);
nand I_14425 (I247114,I246820,I246973);
nand I_14426 (I247131,I246888,I247114);
DFFARX1 I_14427 (I247131,I1862,I246786,I246766,);
not I_14428 (I247162,I246956);
nor I_14429 (I246775,I247162,I247007);
nand I_14430 (I246772,I246939,I247162);
nor I_14431 (I247207,I246905,I246956);
nand I_14432 (I246769,I247207,I246820);
not I_14433 (I247262,I1869);
or I_14434 (I247279,I8217,I8205);
nor I_14435 (I247296,I247279,I8199);
nor I_14436 (I247313,I8202,I8211);
or I_14437 (I247330,I247313,I8214);
nor I_14438 (I247347,I8196,I8199);
nand I_14439 (I247364,I247347,I247330);
not I_14440 (I247381,I247364);
nand I_14441 (I247398,I247296,I247381);
nor I_14442 (I247415,I247296,I247381);
nand I_14443 (I247432,I8202,I8208);
nor I_14444 (I247449,I247432,I8196);
nor I_14445 (I247466,I247432,I247449);
not I_14446 (I247483,I247449);
nor I_14447 (I247254,I247483,I247398);
or I_14448 (I247239,I247296,I247483);
nor I_14449 (I247528,I247296,I247449);
nor I_14450 (I247233,I247432,I247528);
nor I_14451 (I247559,I247466,I247528);
nor I_14452 (I247236,I247381,I247559);
nand I_14453 (I247590,I247296,I247449);
nand I_14454 (I247607,I247364,I247590);
DFFARX1 I_14455 (I247607,I1862,I247262,I247242,);
not I_14456 (I247638,I247432);
nor I_14457 (I247251,I247638,I247483);
nand I_14458 (I247248,I247415,I247638);
nor I_14459 (I247683,I247381,I247432);
nand I_14460 (I247245,I247683,I247296);
not I_14461 (I247738,I1869);
or I_14462 (I247755,I56323,I56332);
nor I_14463 (I247772,I247755,I56347);
nor I_14464 (I247789,I56344,I56326);
or I_14465 (I247806,I247789,I56326);
nor I_14466 (I247823,I56323,I56329);
nand I_14467 (I247840,I247823,I247806);
not I_14468 (I247857,I247840);
nand I_14469 (I247874,I247772,I247857);
nor I_14470 (I247891,I247772,I247857);
nand I_14471 (I247908,I56335,I56338);
nor I_14472 (I247925,I247908,I56341);
nor I_14473 (I247942,I247908,I247925);
not I_14474 (I247959,I247925);
nor I_14475 (I247730,I247959,I247874);
or I_14476 (I247715,I247772,I247959);
nor I_14477 (I248004,I247772,I247925);
nor I_14478 (I247709,I247908,I248004);
nor I_14479 (I248035,I247942,I248004);
nor I_14480 (I247712,I247857,I248035);
nand I_14481 (I248066,I247772,I247925);
nand I_14482 (I248083,I247840,I248066);
DFFARX1 I_14483 (I248083,I1862,I247738,I247718,);
not I_14484 (I248114,I247908);
nor I_14485 (I247727,I248114,I247959);
nand I_14486 (I247724,I247891,I248114);
nor I_14487 (I248159,I247857,I247908);
nand I_14488 (I247721,I248159,I247772);
not I_14489 (I248214,I1869);
or I_14490 (I248231,I359994,I360015);
nor I_14491 (I248248,I248231,I360000);
nor I_14492 (I248265,I359994,I360012);
or I_14493 (I248282,I248265,I360003);
nor I_14494 (I248299,I359997,I359997);
nand I_14495 (I248316,I248299,I248282);
not I_14496 (I248333,I248316);
nand I_14497 (I248350,I248248,I248333);
nor I_14498 (I248367,I248248,I248333);
nand I_14499 (I248384,I360006,I360009);
nor I_14500 (I248401,I248384,I360000);
nor I_14501 (I248418,I248384,I248401);
not I_14502 (I248435,I248401);
nor I_14503 (I248206,I248435,I248350);
or I_14504 (I248191,I248248,I248435);
nor I_14505 (I248480,I248248,I248401);
nor I_14506 (I248185,I248384,I248480);
nor I_14507 (I248511,I248418,I248480);
nor I_14508 (I248188,I248333,I248511);
nand I_14509 (I248542,I248248,I248401);
nand I_14510 (I248559,I248316,I248542);
DFFARX1 I_14511 (I248559,I1862,I248214,I248194,);
not I_14512 (I248590,I248384);
nor I_14513 (I248203,I248590,I248435);
nand I_14514 (I248200,I248367,I248590);
nor I_14515 (I248635,I248333,I248384);
nand I_14516 (I248197,I248635,I248248);
not I_14517 (I248690,I1869);
or I_14518 (I248707,I410113,I410116);
nor I_14519 (I248724,I248707,I410113);
nor I_14520 (I248741,I410110,I410128);
or I_14521 (I248758,I248741,I410116);
nor I_14522 (I248775,I410119,I410110);
nand I_14523 (I248792,I248775,I248758);
not I_14524 (I248809,I248792);
nand I_14525 (I248826,I248724,I248809);
nor I_14526 (I248843,I248724,I248809);
nand I_14527 (I248860,I410125,I410122);
nor I_14528 (I248877,I248860,I410119);
nor I_14529 (I248894,I248860,I248877);
not I_14530 (I248911,I248877);
nor I_14531 (I248682,I248911,I248826);
or I_14532 (I248667,I248724,I248911);
nor I_14533 (I248956,I248724,I248877);
nor I_14534 (I248661,I248860,I248956);
nor I_14535 (I248987,I248894,I248956);
nor I_14536 (I248664,I248809,I248987);
nand I_14537 (I249018,I248724,I248877);
nand I_14538 (I249035,I248792,I249018);
DFFARX1 I_14539 (I249035,I1862,I248690,I248670,);
not I_14540 (I249066,I248860);
nor I_14541 (I248679,I249066,I248911);
nand I_14542 (I248676,I248843,I249066);
nor I_14543 (I249111,I248809,I248860);
nand I_14544 (I248673,I249111,I248724);
not I_14545 (I249166,I1869);
or I_14546 (I249183,I297811,I297808);
nor I_14547 (I249200,I249183,I297817);
nor I_14548 (I249217,I297829,I297814);
or I_14549 (I249234,I249217,I297808);
nor I_14550 (I249251,I297820,I297811);
nand I_14551 (I249268,I249251,I249234);
not I_14552 (I249285,I249268);
nand I_14553 (I249302,I249200,I249285);
nor I_14554 (I249319,I249200,I249285);
nand I_14555 (I249336,I297814,I297826);
nor I_14556 (I249353,I249336,I297823);
nor I_14557 (I249370,I249336,I249353);
not I_14558 (I249387,I249353);
nor I_14559 (I249158,I249387,I249302);
or I_14560 (I249143,I249200,I249387);
nor I_14561 (I249432,I249200,I249353);
nor I_14562 (I249137,I249336,I249432);
nor I_14563 (I249463,I249370,I249432);
nor I_14564 (I249140,I249285,I249463);
nand I_14565 (I249494,I249200,I249353);
nand I_14566 (I249511,I249268,I249494);
DFFARX1 I_14567 (I249511,I1862,I249166,I249146,);
not I_14568 (I249542,I249336);
nor I_14569 (I249155,I249542,I249387);
nand I_14570 (I249152,I249319,I249542);
nor I_14571 (I249587,I249285,I249336);
nand I_14572 (I249149,I249587,I249200);
not I_14573 (I249642,I1869);
or I_14574 (I249659,I138950,I138935);
nor I_14575 (I249676,I249659,I138929);
nor I_14576 (I249693,I138926,I138947);
or I_14577 (I249710,I249693,I138944);
nor I_14578 (I249727,I138932,I138929);
nand I_14579 (I249744,I249727,I249710);
not I_14580 (I249761,I249744);
nand I_14581 (I249778,I249676,I249761);
nor I_14582 (I249795,I249676,I249761);
nand I_14583 (I249812,I138938,I138941);
nor I_14584 (I249829,I249812,I138926);
nor I_14585 (I249846,I249812,I249829);
not I_14586 (I249863,I249829);
nor I_14587 (I249634,I249863,I249778);
or I_14588 (I249619,I249676,I249863);
nor I_14589 (I249908,I249676,I249829);
nor I_14590 (I249613,I249812,I249908);
nor I_14591 (I249939,I249846,I249908);
nor I_14592 (I249616,I249761,I249939);
nand I_14593 (I249970,I249676,I249829);
nand I_14594 (I249987,I249744,I249970);
DFFARX1 I_14595 (I249987,I1862,I249642,I249622,);
not I_14596 (I250018,I249812);
nor I_14597 (I249631,I250018,I249863);
nand I_14598 (I249628,I249795,I250018);
nor I_14599 (I250063,I249761,I249812);
nand I_14600 (I249625,I250063,I249676);
not I_14601 (I250118,I1869);
or I_14602 (I250135,I370775,I370778);
nor I_14603 (I250152,I250135,I370775);
nor I_14604 (I250169,I370772,I370790);
or I_14605 (I250186,I250169,I370778);
nor I_14606 (I250203,I370781,I370772);
nand I_14607 (I250220,I250203,I250186);
not I_14608 (I250237,I250220);
nand I_14609 (I250254,I250152,I250237);
nor I_14610 (I250271,I250152,I250237);
nand I_14611 (I250288,I370787,I370784);
nor I_14612 (I250305,I250288,I370781);
nor I_14613 (I250322,I250288,I250305);
not I_14614 (I250339,I250305);
nor I_14615 (I250110,I250339,I250254);
or I_14616 (I250095,I250152,I250339);
nor I_14617 (I250384,I250152,I250305);
nor I_14618 (I250089,I250288,I250384);
nor I_14619 (I250415,I250322,I250384);
nor I_14620 (I250092,I250237,I250415);
nand I_14621 (I250446,I250152,I250305);
nand I_14622 (I250463,I250220,I250446);
DFFARX1 I_14623 (I250463,I1862,I250118,I250098,);
not I_14624 (I250494,I250288);
nor I_14625 (I250107,I250494,I250339);
nand I_14626 (I250104,I250271,I250494);
nor I_14627 (I250539,I250237,I250288);
nand I_14628 (I250101,I250539,I250152);
not I_14629 (I250594,I1869);
or I_14630 (I250611,I25213,I25222);
nor I_14631 (I250628,I250611,I25237);
nor I_14632 (I250645,I25234,I25216);
or I_14633 (I250662,I250645,I25216);
nor I_14634 (I250679,I25213,I25219);
nand I_14635 (I250696,I250679,I250662);
not I_14636 (I250713,I250696);
nand I_14637 (I250730,I250628,I250713);
nor I_14638 (I250747,I250628,I250713);
nand I_14639 (I250764,I25225,I25228);
nor I_14640 (I250781,I250764,I25231);
nor I_14641 (I250798,I250764,I250781);
not I_14642 (I250815,I250781);
nor I_14643 (I250586,I250815,I250730);
or I_14644 (I250571,I250628,I250815);
nor I_14645 (I250860,I250628,I250781);
nor I_14646 (I250565,I250764,I250860);
nor I_14647 (I250891,I250798,I250860);
nor I_14648 (I250568,I250713,I250891);
nand I_14649 (I250922,I250628,I250781);
nand I_14650 (I250939,I250696,I250922);
DFFARX1 I_14651 (I250939,I1862,I250594,I250574,);
not I_14652 (I250970,I250764);
nor I_14653 (I250583,I250970,I250815);
nand I_14654 (I250580,I250747,I250970);
nor I_14655 (I251015,I250713,I250764);
nand I_14656 (I250577,I251015,I250628);
not I_14657 (I251070,I1869);
or I_14658 (I251087,I139477,I139462);
nor I_14659 (I251104,I251087,I139456);
nor I_14660 (I251121,I139453,I139474);
or I_14661 (I251138,I251121,I139471);
nor I_14662 (I251155,I139459,I139456);
nand I_14663 (I251172,I251155,I251138);
not I_14664 (I251189,I251172);
nand I_14665 (I251206,I251104,I251189);
nor I_14666 (I251223,I251104,I251189);
nand I_14667 (I251240,I139465,I139468);
nor I_14668 (I251257,I251240,I139453);
nor I_14669 (I251274,I251240,I251257);
not I_14670 (I251291,I251257);
nor I_14671 (I251062,I251291,I251206);
or I_14672 (I251047,I251104,I251291);
nor I_14673 (I251336,I251104,I251257);
nor I_14674 (I251041,I251240,I251336);
nor I_14675 (I251367,I251274,I251336);
nor I_14676 (I251044,I251189,I251367);
nand I_14677 (I251398,I251104,I251257);
nand I_14678 (I251415,I251172,I251398);
DFFARX1 I_14679 (I251415,I1862,I251070,I251050,);
not I_14680 (I251446,I251240);
nor I_14681 (I251059,I251446,I251291);
nand I_14682 (I251056,I251223,I251446);
nor I_14683 (I251491,I251189,I251240);
nand I_14684 (I251053,I251491,I251104);
not I_14685 (I251546,I1869);
or I_14686 (I251563,I308875,I308896);
nor I_14687 (I251580,I251563,I308881);
nor I_14688 (I251597,I308875,I308893);
or I_14689 (I251614,I251597,I308884);
nor I_14690 (I251631,I308878,I308878);
nand I_14691 (I251648,I251631,I251614);
not I_14692 (I251665,I251648);
nand I_14693 (I251682,I251580,I251665);
nor I_14694 (I251699,I251580,I251665);
nand I_14695 (I251716,I308887,I308890);
nor I_14696 (I251733,I251716,I308881);
nor I_14697 (I251750,I251716,I251733);
not I_14698 (I251767,I251733);
nor I_14699 (I251538,I251767,I251682);
or I_14700 (I251523,I251580,I251767);
nor I_14701 (I251812,I251580,I251733);
nor I_14702 (I251517,I251716,I251812);
nor I_14703 (I251843,I251750,I251812);
nor I_14704 (I251520,I251665,I251843);
nand I_14705 (I251874,I251580,I251733);
nand I_14706 (I251891,I251648,I251874);
DFFARX1 I_14707 (I251891,I1862,I251546,I251526,);
not I_14708 (I251922,I251716);
nor I_14709 (I251535,I251922,I251767);
nand I_14710 (I251532,I251699,I251922);
nor I_14711 (I251967,I251665,I251716);
nand I_14712 (I251529,I251967,I251580);
not I_14713 (I252022,I1869);
or I_14714 (I252039,I174259,I174244);
nor I_14715 (I252056,I252039,I174238);
nor I_14716 (I252073,I174235,I174256);
or I_14717 (I252090,I252073,I174253);
nor I_14718 (I252107,I174241,I174238);
nand I_14719 (I252124,I252107,I252090);
not I_14720 (I252141,I252124);
nand I_14721 (I252158,I252056,I252141);
nor I_14722 (I252175,I252056,I252141);
nand I_14723 (I252192,I174247,I174250);
nor I_14724 (I252209,I252192,I174235);
nor I_14725 (I252226,I252192,I252209);
not I_14726 (I252243,I252209);
nor I_14727 (I252014,I252243,I252158);
or I_14728 (I251999,I252056,I252243);
nor I_14729 (I252288,I252056,I252209);
nor I_14730 (I251993,I252192,I252288);
nor I_14731 (I252319,I252226,I252288);
nor I_14732 (I251996,I252141,I252319);
nand I_14733 (I252350,I252056,I252209);
nand I_14734 (I252367,I252124,I252350);
DFFARX1 I_14735 (I252367,I1862,I252022,I252002,);
not I_14736 (I252398,I252192);
nor I_14737 (I252011,I252398,I252243);
nand I_14738 (I252008,I252175,I252398);
nor I_14739 (I252443,I252141,I252192);
nand I_14740 (I252005,I252443,I252056);
not I_14741 (I252498,I1869);
or I_14742 (I252515,I404367,I404370);
nor I_14743 (I252532,I252515,I404367);
nor I_14744 (I252549,I404364,I404382);
or I_14745 (I252566,I252549,I404370);
nor I_14746 (I252583,I404373,I404364);
nand I_14747 (I252600,I252583,I252566);
not I_14748 (I252617,I252600);
nand I_14749 (I252634,I252532,I252617);
nor I_14750 (I252651,I252532,I252617);
nand I_14751 (I252668,I404379,I404376);
nor I_14752 (I252685,I252668,I404373);
nor I_14753 (I252702,I252668,I252685);
not I_14754 (I252719,I252685);
nor I_14755 (I252490,I252719,I252634);
or I_14756 (I252475,I252532,I252719);
nor I_14757 (I252764,I252532,I252685);
nor I_14758 (I252469,I252668,I252764);
nor I_14759 (I252795,I252702,I252764);
nor I_14760 (I252472,I252617,I252795);
nand I_14761 (I252826,I252532,I252685);
nand I_14762 (I252843,I252600,I252826);
DFFARX1 I_14763 (I252843,I1862,I252498,I252478,);
not I_14764 (I252874,I252668);
nor I_14765 (I252487,I252874,I252719);
nand I_14766 (I252484,I252651,I252874);
nor I_14767 (I252919,I252617,I252668);
nand I_14768 (I252481,I252919,I252532);
not I_14769 (I252974,I1869);
or I_14770 (I252991,I69583,I69592);
nor I_14771 (I253008,I252991,I69607);
nor I_14772 (I253025,I69604,I69586);
or I_14773 (I253042,I253025,I69586);
nor I_14774 (I253059,I69583,I69589);
nand I_14775 (I253076,I253059,I253042);
not I_14776 (I253093,I253076);
nand I_14777 (I253110,I253008,I253093);
nor I_14778 (I253127,I253008,I253093);
nand I_14779 (I253144,I69595,I69598);
nor I_14780 (I253161,I253144,I69601);
nor I_14781 (I253178,I253144,I253161);
not I_14782 (I253195,I253161);
nor I_14783 (I252966,I253195,I253110);
or I_14784 (I252951,I253008,I253195);
nor I_14785 (I253240,I253008,I253161);
nor I_14786 (I252945,I253144,I253240);
nor I_14787 (I253271,I253178,I253240);
nor I_14788 (I252948,I253093,I253271);
nand I_14789 (I253302,I253008,I253161);
nand I_14790 (I253319,I253076,I253302);
DFFARX1 I_14791 (I253319,I1862,I252974,I252954,);
not I_14792 (I253350,I253144);
nor I_14793 (I252963,I253350,I253195);
nand I_14794 (I252960,I253127,I253350);
nor I_14795 (I253395,I253093,I253144);
nand I_14796 (I252957,I253395,I253008);
not I_14797 (I253450,I1869);
or I_14798 (I253467,I128937,I128922);
nor I_14799 (I253484,I253467,I128916);
nor I_14800 (I253501,I128913,I128934);
or I_14801 (I253518,I253501,I128931);
nor I_14802 (I253535,I128919,I128916);
nand I_14803 (I253552,I253535,I253518);
not I_14804 (I253569,I253552);
nand I_14805 (I253586,I253484,I253569);
nor I_14806 (I253603,I253484,I253569);
nand I_14807 (I253620,I128925,I128928);
nor I_14808 (I253637,I253620,I128913);
nor I_14809 (I253654,I253620,I253637);
not I_14810 (I253671,I253637);
nor I_14811 (I253442,I253671,I253586);
or I_14812 (I253427,I253484,I253671);
nor I_14813 (I253716,I253484,I253637);
nor I_14814 (I253421,I253620,I253716);
nor I_14815 (I253747,I253654,I253716);
nor I_14816 (I253424,I253569,I253747);
nand I_14817 (I253778,I253484,I253637);
nand I_14818 (I253795,I253552,I253778);
DFFARX1 I_14819 (I253795,I1862,I253450,I253430,);
not I_14820 (I253826,I253620);
nor I_14821 (I253439,I253826,I253671);
nand I_14822 (I253436,I253603,I253826);
nor I_14823 (I253871,I253569,I253620);
nand I_14824 (I253433,I253871,I253484);
not I_14825 (I253926,I1869);
or I_14826 (I253943,I306767,I306788);
nor I_14827 (I253960,I253943,I306773);
nor I_14828 (I253977,I306767,I306785);
or I_14829 (I253994,I253977,I306776);
nor I_14830 (I254011,I306770,I306770);
nand I_14831 (I254028,I254011,I253994);
not I_14832 (I254045,I254028);
nand I_14833 (I254062,I253960,I254045);
nor I_14834 (I254079,I253960,I254045);
nand I_14835 (I254096,I306779,I306782);
nor I_14836 (I254113,I254096,I306773);
nor I_14837 (I254130,I254096,I254113);
not I_14838 (I254147,I254113);
nor I_14839 (I253918,I254147,I254062);
or I_14840 (I253903,I253960,I254147);
nor I_14841 (I254192,I253960,I254113);
nor I_14842 (I253897,I254096,I254192);
nor I_14843 (I254223,I254130,I254192);
nor I_14844 (I253900,I254045,I254223);
nand I_14845 (I254254,I253960,I254113);
nand I_14846 (I254271,I254028,I254254);
DFFARX1 I_14847 (I254271,I1862,I253926,I253906,);
not I_14848 (I254302,I254096);
nor I_14849 (I253915,I254302,I254147);
nand I_14850 (I253912,I254079,I254302);
nor I_14851 (I254347,I254045,I254096);
nand I_14852 (I253909,I254347,I253960);
not I_14853 (I254402,I1869);
or I_14854 (I254419,I390223,I390226);
nor I_14855 (I254436,I254419,I390223);
nor I_14856 (I254453,I390220,I390238);
or I_14857 (I254470,I254453,I390226);
nor I_14858 (I254487,I390229,I390220);
nand I_14859 (I254504,I254487,I254470);
not I_14860 (I254521,I254504);
nand I_14861 (I254538,I254436,I254521);
nor I_14862 (I254555,I254436,I254521);
nand I_14863 (I254572,I390235,I390232);
nor I_14864 (I254589,I254572,I390229);
nor I_14865 (I254606,I254572,I254589);
not I_14866 (I254623,I254589);
nor I_14867 (I254394,I254623,I254538);
or I_14868 (I254379,I254436,I254623);
nor I_14869 (I254668,I254436,I254589);
nor I_14870 (I254373,I254572,I254668);
nor I_14871 (I254699,I254606,I254668);
nor I_14872 (I254376,I254521,I254699);
nand I_14873 (I254730,I254436,I254589);
nand I_14874 (I254747,I254504,I254730);
DFFARX1 I_14875 (I254747,I1862,I254402,I254382,);
not I_14876 (I254778,I254572);
nor I_14877 (I254391,I254778,I254623);
nand I_14878 (I254388,I254555,I254778);
nor I_14879 (I254823,I254521,I254572);
nand I_14880 (I254385,I254823,I254436);
not I_14881 (I254878,I1869);
or I_14882 (I254895,I406135,I406138);
nor I_14883 (I254912,I254895,I406135);
nor I_14884 (I254929,I406132,I406150);
or I_14885 (I254946,I254929,I406138);
nor I_14886 (I254963,I406141,I406132);
nand I_14887 (I254980,I254963,I254946);
not I_14888 (I254997,I254980);
nand I_14889 (I255014,I254912,I254997);
nor I_14890 (I255031,I254912,I254997);
nand I_14891 (I255048,I406147,I406144);
nor I_14892 (I255065,I255048,I406141);
nor I_14893 (I255082,I255048,I255065);
not I_14894 (I255099,I255065);
nor I_14895 (I254870,I255099,I255014);
or I_14896 (I254855,I254912,I255099);
nor I_14897 (I255144,I254912,I255065);
nor I_14898 (I254849,I255048,I255144);
nor I_14899 (I255175,I255082,I255144);
nor I_14900 (I254852,I254997,I255175);
nand I_14901 (I255206,I254912,I255065);
nand I_14902 (I255223,I254980,I255206);
DFFARX1 I_14903 (I255223,I1862,I254878,I254858,);
not I_14904 (I255254,I255048);
nor I_14905 (I254867,I255254,I255099);
nand I_14906 (I254864,I255031,I255254);
nor I_14907 (I255299,I254997,I255048);
nand I_14908 (I254861,I255299,I254912);
not I_14909 (I255354,I1869);
or I_14910 (I255371,I320469,I320490);
nor I_14911 (I255388,I255371,I320475);
nor I_14912 (I255405,I320469,I320487);
or I_14913 (I255422,I255405,I320478);
nor I_14914 (I255439,I320472,I320472);
nand I_14915 (I255456,I255439,I255422);
not I_14916 (I255473,I255456);
nand I_14917 (I255490,I255388,I255473);
nor I_14918 (I255507,I255388,I255473);
nand I_14919 (I255524,I320481,I320484);
nor I_14920 (I255541,I255524,I320475);
nor I_14921 (I255558,I255524,I255541);
not I_14922 (I255575,I255541);
nor I_14923 (I255346,I255575,I255490);
or I_14924 (I255331,I255388,I255575);
nor I_14925 (I255620,I255388,I255541);
nor I_14926 (I255325,I255524,I255620);
nor I_14927 (I255651,I255558,I255620);
nor I_14928 (I255328,I255473,I255651);
nand I_14929 (I255682,I255388,I255541);
nand I_14930 (I255699,I255456,I255682);
DFFARX1 I_14931 (I255699,I1862,I255354,I255334,);
not I_14932 (I255730,I255524);
nor I_14933 (I255343,I255730,I255575);
nand I_14934 (I255340,I255507,I255730);
nor I_14935 (I255775,I255473,I255524);
nand I_14936 (I255337,I255775,I255388);
not I_14937 (I255830,I1869);
or I_14938 (I255847,I141058,I141043);
nor I_14939 (I255864,I255847,I141037);
nor I_14940 (I255881,I141034,I141055);
or I_14941 (I255898,I255881,I141052);
nor I_14942 (I255915,I141040,I141037);
nand I_14943 (I255932,I255915,I255898);
not I_14944 (I255949,I255932);
nand I_14945 (I255966,I255864,I255949);
nor I_14946 (I255983,I255864,I255949);
nand I_14947 (I256000,I141046,I141049);
nor I_14948 (I256017,I256000,I141034);
nor I_14949 (I256034,I256000,I256017);
not I_14950 (I256051,I256017);
nor I_14951 (I255822,I256051,I255966);
or I_14952 (I255807,I255864,I256051);
nor I_14953 (I256096,I255864,I256017);
nor I_14954 (I255801,I256000,I256096);
nor I_14955 (I256127,I256034,I256096);
nor I_14956 (I255804,I255949,I256127);
nand I_14957 (I256158,I255864,I256017);
nand I_14958 (I256175,I255932,I256158);
DFFARX1 I_14959 (I256175,I1862,I255830,I255810,);
not I_14960 (I256206,I256000);
nor I_14961 (I255819,I256206,I256051);
nand I_14962 (I255816,I255983,I256206);
nor I_14963 (I256251,I255949,I256000);
nand I_14964 (I255813,I256251,I255864);
not I_14965 (I256306,I1869);
or I_14966 (I256323,I286744,I286741);
nor I_14967 (I256340,I256323,I286750);
nor I_14968 (I256357,I286762,I286747);
or I_14969 (I256374,I256357,I286741);
nor I_14970 (I256391,I286753,I286744);
nand I_14971 (I256408,I256391,I256374);
not I_14972 (I256425,I256408);
nand I_14973 (I256442,I256340,I256425);
nor I_14974 (I256459,I256340,I256425);
nand I_14975 (I256476,I286747,I286759);
nor I_14976 (I256493,I256476,I286756);
nor I_14977 (I256510,I256476,I256493);
not I_14978 (I256527,I256493);
nor I_14979 (I256298,I256527,I256442);
or I_14980 (I256283,I256340,I256527);
nor I_14981 (I256572,I256340,I256493);
nor I_14982 (I256277,I256476,I256572);
nor I_14983 (I256603,I256510,I256572);
nor I_14984 (I256280,I256425,I256603);
nand I_14985 (I256634,I256340,I256493);
nand I_14986 (I256651,I256408,I256634);
DFFARX1 I_14987 (I256651,I1862,I256306,I256286,);
not I_14988 (I256682,I256476);
nor I_14989 (I256295,I256682,I256527);
nand I_14990 (I256292,I256459,I256682);
nor I_14991 (I256727,I256425,I256476);
nand I_14992 (I256289,I256727,I256340);
not I_14993 (I256782,I1869);
or I_14994 (I256799,I314672,I314693);
nor I_14995 (I256816,I256799,I314678);
nor I_14996 (I256833,I314672,I314690);
or I_14997 (I256850,I256833,I314681);
nor I_14998 (I256867,I314675,I314675);
nand I_14999 (I256884,I256867,I256850);
not I_15000 (I256901,I256884);
nand I_15001 (I256918,I256816,I256901);
nor I_15002 (I256935,I256816,I256901);
nand I_15003 (I256952,I314684,I314687);
nor I_15004 (I256969,I256952,I314678);
nor I_15005 (I256986,I256952,I256969);
not I_15006 (I257003,I256969);
nor I_15007 (I256774,I257003,I256918);
or I_15008 (I256759,I256816,I257003);
nor I_15009 (I257048,I256816,I256969);
nor I_15010 (I256753,I256952,I257048);
nor I_15011 (I257079,I256986,I257048);
nor I_15012 (I256756,I256901,I257079);
nand I_15013 (I257110,I256816,I256969);
nand I_15014 (I257127,I256884,I257110);
DFFARX1 I_15015 (I257127,I1862,I256782,I256762,);
not I_15016 (I257158,I256952);
nor I_15017 (I256771,I257158,I257003);
nand I_15018 (I256768,I256935,I257158);
nor I_15019 (I257203,I256901,I256952);
nand I_15020 (I256765,I257203,I256816);
not I_15021 (I257258,I1869);
or I_15022 (I257275,I48163,I48172);
nor I_15023 (I257292,I257275,I48187);
nor I_15024 (I257309,I48184,I48166);
or I_15025 (I257326,I257309,I48166);
nor I_15026 (I257343,I48163,I48169);
nand I_15027 (I257360,I257343,I257326);
not I_15028 (I257377,I257360);
nand I_15029 (I257394,I257292,I257377);
nor I_15030 (I257411,I257292,I257377);
nand I_15031 (I257428,I48175,I48178);
nor I_15032 (I257445,I257428,I48181);
nor I_15033 (I257462,I257428,I257445);
not I_15034 (I257479,I257445);
nor I_15035 (I257250,I257479,I257394);
or I_15036 (I257235,I257292,I257479);
nor I_15037 (I257524,I257292,I257445);
nor I_15038 (I257229,I257428,I257524);
nor I_15039 (I257555,I257462,I257524);
nor I_15040 (I257232,I257377,I257555);
nand I_15041 (I257586,I257292,I257445);
nand I_15042 (I257603,I257360,I257586);
DFFARX1 I_15043 (I257603,I1862,I257258,I257238,);
not I_15044 (I257634,I257428);
nor I_15045 (I257247,I257634,I257479);
nand I_15046 (I257244,I257411,I257634);
nor I_15047 (I257679,I257377,I257428);
nand I_15048 (I257241,I257679,I257292);
not I_15049 (I257734,I1869);
or I_15050 (I257751,I373427,I373430);
nor I_15051 (I257768,I257751,I373427);
nor I_15052 (I257785,I373424,I373442);
or I_15053 (I257802,I257785,I373430);
nor I_15054 (I257819,I373433,I373424);
nand I_15055 (I257836,I257819,I257802);
not I_15056 (I257853,I257836);
nand I_15057 (I257870,I257768,I257853);
nor I_15058 (I257887,I257768,I257853);
nand I_15059 (I257904,I373439,I373436);
nor I_15060 (I257921,I257904,I373433);
nor I_15061 (I257938,I257904,I257921);
not I_15062 (I257955,I257921);
nor I_15063 (I257726,I257955,I257870);
or I_15064 (I257711,I257768,I257955);
nor I_15065 (I258000,I257768,I257921);
nor I_15066 (I257705,I257904,I258000);
nor I_15067 (I258031,I257938,I258000);
nor I_15068 (I257708,I257853,I258031);
nand I_15069 (I258062,I257768,I257921);
nand I_15070 (I258079,I257836,I258062);
DFFARX1 I_15071 (I258079,I1862,I257734,I257714,);
not I_15072 (I258110,I257904);
nor I_15073 (I257723,I258110,I257955);
nand I_15074 (I257720,I257887,I258110);
nor I_15075 (I258155,I257853,I257904);
nand I_15076 (I257717,I258155,I257768);
not I_15077 (I258210,I1869);
or I_15078 (I258227,I18073,I18082);
nor I_15079 (I258244,I258227,I18097);
nor I_15080 (I258261,I18094,I18076);
or I_15081 (I258278,I258261,I18076);
nor I_15082 (I258295,I18073,I18079);
nand I_15083 (I258312,I258295,I258278);
not I_15084 (I258329,I258312);
nand I_15085 (I258346,I258244,I258329);
nor I_15086 (I258363,I258244,I258329);
nand I_15087 (I258380,I18085,I18088);
nor I_15088 (I258397,I258380,I18091);
nor I_15089 (I258414,I258380,I258397);
not I_15090 (I258431,I258397);
nor I_15091 (I258202,I258431,I258346);
or I_15092 (I258187,I258244,I258431);
nor I_15093 (I258476,I258244,I258397);
nor I_15094 (I258181,I258380,I258476);
nor I_15095 (I258507,I258414,I258476);
nor I_15096 (I258184,I258329,I258507);
nand I_15097 (I258538,I258244,I258397);
nand I_15098 (I258555,I258312,I258538);
DFFARX1 I_15099 (I258555,I1862,I258210,I258190,);
not I_15100 (I258586,I258380);
nor I_15101 (I258199,I258586,I258431);
nand I_15102 (I258196,I258363,I258586);
nor I_15103 (I258631,I258329,I258380);
nand I_15104 (I258193,I258631,I258244);
not I_15105 (I258686,I1869);
or I_15106 (I258703,I147382,I147367);
nor I_15107 (I258720,I258703,I147361);
nor I_15108 (I258737,I147358,I147379);
or I_15109 (I258754,I258737,I147376);
nor I_15110 (I258771,I147364,I147361);
nand I_15111 (I258788,I258771,I258754);
not I_15112 (I258805,I258788);
nand I_15113 (I258822,I258720,I258805);
nor I_15114 (I258839,I258720,I258805);
nand I_15115 (I258856,I147370,I147373);
nor I_15116 (I258873,I258856,I147358);
nor I_15117 (I258890,I258856,I258873);
not I_15118 (I258907,I258873);
nor I_15119 (I258678,I258907,I258822);
or I_15120 (I258663,I258720,I258907);
nor I_15121 (I258952,I258720,I258873);
nor I_15122 (I258657,I258856,I258952);
nor I_15123 (I258983,I258890,I258952);
nor I_15124 (I258660,I258805,I258983);
nand I_15125 (I259014,I258720,I258873);
nand I_15126 (I259031,I258788,I259014);
DFFARX1 I_15127 (I259031,I1862,I258686,I258666,);
not I_15128 (I259062,I258856);
nor I_15129 (I258675,I259062,I258907);
nand I_15130 (I258672,I258839,I259062);
nor I_15131 (I259107,I258805,I258856);
nand I_15132 (I258669,I259107,I258720);
not I_15133 (I259162,I1869);
or I_15134 (I259179,I317307,I317328);
nor I_15135 (I259196,I259179,I317313);
nor I_15136 (I259213,I317307,I317325);
or I_15137 (I259230,I259213,I317316);
nor I_15138 (I259247,I317310,I317310);
nand I_15139 (I259264,I259247,I259230);
not I_15140 (I259281,I259264);
nand I_15141 (I259298,I259196,I259281);
nor I_15142 (I259315,I259196,I259281);
nand I_15143 (I259332,I317319,I317322);
nor I_15144 (I259349,I259332,I317313);
nor I_15145 (I259366,I259332,I259349);
not I_15146 (I259383,I259349);
nor I_15147 (I259154,I259383,I259298);
or I_15148 (I259139,I259196,I259383);
nor I_15149 (I259428,I259196,I259349);
nor I_15150 (I259133,I259332,I259428);
nor I_15151 (I259459,I259366,I259428);
nor I_15152 (I259136,I259281,I259459);
nand I_15153 (I259490,I259196,I259349);
nand I_15154 (I259507,I259264,I259490);
DFFARX1 I_15155 (I259507,I1862,I259162,I259142,);
not I_15156 (I259538,I259332);
nor I_15157 (I259151,I259538,I259383);
nand I_15158 (I259148,I259315,I259538);
nor I_15159 (I259583,I259281,I259332);
nand I_15160 (I259145,I259583,I259196);
not I_15161 (I259638,I1869);
or I_15162 (I259655,I181637,I181622);
nor I_15163 (I259672,I259655,I181616);
nor I_15164 (I259689,I181613,I181634);
or I_15165 (I259706,I259689,I181631);
nor I_15166 (I259723,I181619,I181616);
nand I_15167 (I259740,I259723,I259706);
not I_15168 (I259757,I259740);
nand I_15169 (I259774,I259672,I259757);
nor I_15170 (I259791,I259672,I259757);
nand I_15171 (I259808,I181625,I181628);
nor I_15172 (I259825,I259808,I181613);
nor I_15173 (I259842,I259808,I259825);
not I_15174 (I259859,I259825);
nor I_15175 (I259630,I259859,I259774);
or I_15176 (I259615,I259672,I259859);
nor I_15177 (I259904,I259672,I259825);
nor I_15178 (I259609,I259808,I259904);
nor I_15179 (I259935,I259842,I259904);
nor I_15180 (I259612,I259757,I259935);
nand I_15181 (I259966,I259672,I259825);
nand I_15182 (I259983,I259740,I259966);
DFFARX1 I_15183 (I259983,I1862,I259638,I259618,);
not I_15184 (I260014,I259808);
nor I_15185 (I259627,I260014,I259859);
nand I_15186 (I259624,I259791,I260014);
nor I_15187 (I260059,I259757,I259808);
nand I_15188 (I259621,I260059,I259672);
not I_15189 (I260114,I1869);
or I_15190 (I260131,I374311,I374314);
nor I_15191 (I260148,I260131,I374311);
nor I_15192 (I260165,I374308,I374326);
or I_15193 (I260182,I260165,I374314);
nor I_15194 (I260199,I374317,I374308);
nand I_15195 (I260216,I260199,I260182);
not I_15196 (I260233,I260216);
nand I_15197 (I260250,I260148,I260233);
nor I_15198 (I260267,I260148,I260233);
nand I_15199 (I260284,I374323,I374320);
nor I_15200 (I260301,I260284,I374317);
nor I_15201 (I260318,I260284,I260301);
not I_15202 (I260335,I260301);
nor I_15203 (I260106,I260335,I260250);
or I_15204 (I260091,I260148,I260335);
nor I_15205 (I260380,I260148,I260301);
nor I_15206 (I260085,I260284,I260380);
nor I_15207 (I260411,I260318,I260380);
nor I_15208 (I260088,I260233,I260411);
nand I_15209 (I260442,I260148,I260301);
nand I_15210 (I260459,I260216,I260442);
DFFARX1 I_15211 (I260459,I1862,I260114,I260094,);
not I_15212 (I260490,I260284);
nor I_15213 (I260103,I260490,I260335);
nand I_15214 (I260100,I260267,I260490);
nor I_15215 (I260535,I260233,I260284);
nand I_15216 (I260097,I260535,I260148);
not I_15217 (I260590,I1869);
or I_15218 (I260607,I106714,I106711);
nor I_15219 (I260624,I260607,I106711);
nor I_15220 (I260641,I106720,I106717);
or I_15221 (I260658,I260641,I106726);
nor I_15222 (I260675,I106729,I106714);
nand I_15223 (I260692,I260675,I260658);
not I_15224 (I260709,I260692);
nand I_15225 (I260726,I260624,I260709);
nor I_15226 (I260743,I260624,I260709);
nand I_15227 (I260760,I106717,I106723);
nor I_15228 (I260777,I260760,I106720);
nor I_15229 (I260794,I260760,I260777);
not I_15230 (I260811,I260777);
nor I_15231 (I260582,I260811,I260726);
or I_15232 (I260567,I260624,I260811);
nor I_15233 (I260856,I260624,I260777);
nor I_15234 (I260561,I260760,I260856);
nor I_15235 (I260887,I260794,I260856);
nor I_15236 (I260564,I260709,I260887);
nand I_15237 (I260918,I260624,I260777);
nand I_15238 (I260935,I260692,I260918);
DFFARX1 I_15239 (I260935,I1862,I260590,I260570,);
not I_15240 (I260966,I260760);
nor I_15241 (I260579,I260966,I260811);
nand I_15242 (I260576,I260743,I260966);
nor I_15243 (I261011,I260709,I260760);
nand I_15244 (I260573,I261011,I260624);
not I_15245 (I261066,I1869);
or I_15246 (I261083,I376521,I376524);
nor I_15247 (I261100,I261083,I376521);
nor I_15248 (I261117,I376518,I376536);
or I_15249 (I261134,I261117,I376524);
nor I_15250 (I261151,I376527,I376518);
nand I_15251 (I261168,I261151,I261134);
not I_15252 (I261185,I261168);
nand I_15253 (I261202,I261100,I261185);
nor I_15254 (I261219,I261100,I261185);
nand I_15255 (I261236,I376533,I376530);
nor I_15256 (I261253,I261236,I376527);
nor I_15257 (I261270,I261236,I261253);
not I_15258 (I261287,I261253);
nor I_15259 (I261058,I261287,I261202);
or I_15260 (I261043,I261100,I261287);
nor I_15261 (I261332,I261100,I261253);
nor I_15262 (I261037,I261236,I261332);
nor I_15263 (I261363,I261270,I261332);
nor I_15264 (I261040,I261185,I261363);
nand I_15265 (I261394,I261100,I261253);
nand I_15266 (I261411,I261168,I261394);
DFFARX1 I_15267 (I261411,I1862,I261066,I261046,);
not I_15268 (I261442,I261236);
nor I_15269 (I261055,I261442,I261287);
nand I_15270 (I261052,I261219,I261442);
nor I_15271 (I261487,I261185,I261236);
nand I_15272 (I261049,I261487,I261100);
not I_15273 (I261542,I1869);
or I_15274 (I261559,I21133,I21142);
nor I_15275 (I261576,I261559,I21157);
nor I_15276 (I261593,I21154,I21136);
or I_15277 (I261610,I261593,I21136);
nor I_15278 (I261627,I21133,I21139);
nand I_15279 (I261644,I261627,I261610);
not I_15280 (I261661,I261644);
nand I_15281 (I261678,I261576,I261661);
nor I_15282 (I261695,I261576,I261661);
nand I_15283 (I261712,I21145,I21148);
nor I_15284 (I261729,I261712,I21151);
nor I_15285 (I261746,I261712,I261729);
not I_15286 (I261763,I261729);
nor I_15287 (I261534,I261763,I261678);
or I_15288 (I261519,I261576,I261763);
nor I_15289 (I261808,I261576,I261729);
nor I_15290 (I261513,I261712,I261808);
nor I_15291 (I261839,I261746,I261808);
nor I_15292 (I261516,I261661,I261839);
nand I_15293 (I261870,I261576,I261729);
nand I_15294 (I261887,I261644,I261870);
DFFARX1 I_15295 (I261887,I1862,I261542,I261522,);
not I_15296 (I261918,I261712);
nor I_15297 (I261531,I261918,I261763);
nand I_15298 (I261528,I261695,I261918);
nor I_15299 (I261963,I261661,I261712);
nand I_15300 (I261525,I261963,I261576);
not I_15301 (I262018,I1869);
or I_15302 (I262035,I27253,I27262);
nor I_15303 (I262052,I262035,I27277);
nor I_15304 (I262069,I27274,I27256);
or I_15305 (I262086,I262069,I27256);
nor I_15306 (I262103,I27253,I27259);
nand I_15307 (I262120,I262103,I262086);
not I_15308 (I262137,I262120);
nand I_15309 (I262154,I262052,I262137);
nor I_15310 (I262171,I262052,I262137);
nand I_15311 (I262188,I27265,I27268);
nor I_15312 (I262205,I262188,I27271);
nor I_15313 (I262222,I262188,I262205);
not I_15314 (I262239,I262205);
nor I_15315 (I262010,I262239,I262154);
or I_15316 (I261995,I262052,I262239);
nor I_15317 (I262284,I262052,I262205);
nor I_15318 (I261989,I262188,I262284);
nor I_15319 (I262315,I262222,I262284);
nor I_15320 (I261992,I262137,I262315);
nand I_15321 (I262346,I262052,I262205);
nand I_15322 (I262363,I262120,I262346);
DFFARX1 I_15323 (I262363,I1862,I262018,I261998,);
not I_15324 (I262394,I262188);
nor I_15325 (I262007,I262394,I262239);
nand I_15326 (I262004,I262171,I262394);
nor I_15327 (I262439,I262137,I262188);
nand I_15328 (I262001,I262439,I262052);
not I_15329 (I262494,I1869);
or I_15330 (I262511,I78763,I78772);
nor I_15331 (I262528,I262511,I78787);
nor I_15332 (I262545,I78784,I78766);
or I_15333 (I262562,I262545,I78766);
nor I_15334 (I262579,I78763,I78769);
nand I_15335 (I262596,I262579,I262562);
not I_15336 (I262613,I262596);
nand I_15337 (I262630,I262528,I262613);
nor I_15338 (I262647,I262528,I262613);
nand I_15339 (I262664,I78775,I78778);
nor I_15340 (I262681,I262664,I78781);
nor I_15341 (I262698,I262664,I262681);
not I_15342 (I262715,I262681);
nor I_15343 (I262486,I262715,I262630);
or I_15344 (I262471,I262528,I262715);
nor I_15345 (I262760,I262528,I262681);
nor I_15346 (I262465,I262664,I262760);
nor I_15347 (I262791,I262698,I262760);
nor I_15348 (I262468,I262613,I262791);
nand I_15349 (I262822,I262528,I262681);
nand I_15350 (I262839,I262596,I262822);
DFFARX1 I_15351 (I262839,I1862,I262494,I262474,);
not I_15352 (I262870,I262664);
nor I_15353 (I262483,I262870,I262715);
nand I_15354 (I262480,I262647,I262870);
nor I_15355 (I262915,I262613,I262664);
nand I_15356 (I262477,I262915,I262528);
not I_15357 (I262970,I1869);
or I_15358 (I262987,I40513,I40522);
nor I_15359 (I263004,I262987,I40537);
nor I_15360 (I263021,I40534,I40516);
or I_15361 (I263038,I263021,I40516);
nor I_15362 (I263055,I40513,I40519);
nand I_15363 (I263072,I263055,I263038);
not I_15364 (I263089,I263072);
nand I_15365 (I263106,I263004,I263089);
nor I_15366 (I263123,I263004,I263089);
nand I_15367 (I263140,I40525,I40528);
nor I_15368 (I263157,I263140,I40531);
nor I_15369 (I263174,I263140,I263157);
not I_15370 (I263191,I263157);
nor I_15371 (I262962,I263191,I263106);
or I_15372 (I262947,I263004,I263191);
nor I_15373 (I263236,I263004,I263157);
nor I_15374 (I262941,I263140,I263236);
nor I_15375 (I263267,I263174,I263236);
nor I_15376 (I262944,I263089,I263267);
nand I_15377 (I263298,I263004,I263157);
nand I_15378 (I263315,I263072,I263298);
DFFARX1 I_15379 (I263315,I1862,I262970,I262950,);
not I_15380 (I263346,I263140);
nor I_15381 (I262959,I263346,I263191);
nand I_15382 (I262956,I263123,I263346);
nor I_15383 (I263391,I263089,I263140);
nand I_15384 (I262953,I263391,I263004);
not I_15385 (I263446,I1869);
or I_15386 (I263463,I64993,I65002);
nor I_15387 (I263480,I263463,I65017);
nor I_15388 (I263497,I65014,I64996);
or I_15389 (I263514,I263497,I64996);
nor I_15390 (I263531,I64993,I64999);
nand I_15391 (I263548,I263531,I263514);
not I_15392 (I263565,I263548);
nand I_15393 (I263582,I263480,I263565);
nor I_15394 (I263599,I263480,I263565);
nand I_15395 (I263616,I65005,I65008);
nor I_15396 (I263633,I263616,I65011);
nor I_15397 (I263650,I263616,I263633);
not I_15398 (I263667,I263633);
nor I_15399 (I263438,I263667,I263582);
or I_15400 (I263423,I263480,I263667);
nor I_15401 (I263712,I263480,I263633);
nor I_15402 (I263417,I263616,I263712);
nor I_15403 (I263743,I263650,I263712);
nor I_15404 (I263420,I263565,I263743);
nand I_15405 (I263774,I263480,I263633);
nand I_15406 (I263791,I263548,I263774);
DFFARX1 I_15407 (I263791,I1862,I263446,I263426,);
not I_15408 (I263822,I263616);
nor I_15409 (I263435,I263822,I263667);
nand I_15410 (I263432,I263599,I263822);
nor I_15411 (I263867,I263565,I263616);
nand I_15412 (I263429,I263867,I263480);
not I_15413 (I263922,I1869);
or I_15414 (I263939,I66013,I66022);
nor I_15415 (I263956,I263939,I66037);
nor I_15416 (I263973,I66034,I66016);
or I_15417 (I263990,I263973,I66016);
nor I_15418 (I264007,I66013,I66019);
nand I_15419 (I264024,I264007,I263990);
not I_15420 (I264041,I264024);
nand I_15421 (I264058,I263956,I264041);
nor I_15422 (I264075,I263956,I264041);
nand I_15423 (I264092,I66025,I66028);
nor I_15424 (I264109,I264092,I66031);
nor I_15425 (I264126,I264092,I264109);
not I_15426 (I264143,I264109);
nor I_15427 (I263914,I264143,I264058);
or I_15428 (I263899,I263956,I264143);
nor I_15429 (I264188,I263956,I264109);
nor I_15430 (I263893,I264092,I264188);
nor I_15431 (I264219,I264126,I264188);
nor I_15432 (I263896,I264041,I264219);
nand I_15433 (I264250,I263956,I264109);
nand I_15434 (I264267,I264024,I264250);
DFFARX1 I_15435 (I264267,I1862,I263922,I263902,);
not I_15436 (I264298,I264092);
nor I_15437 (I263911,I264298,I264143);
nand I_15438 (I263908,I264075,I264298);
nor I_15439 (I264343,I264041,I264092);
nand I_15440 (I263905,I264343,I263956);
not I_15441 (I264398,I1869);
or I_15442 (I264415,I45103,I45112);
nor I_15443 (I264432,I264415,I45127);
nor I_15444 (I264449,I45124,I45106);
or I_15445 (I264466,I264449,I45106);
nor I_15446 (I264483,I45103,I45109);
nand I_15447 (I264500,I264483,I264466);
not I_15448 (I264517,I264500);
nand I_15449 (I264534,I264432,I264517);
nor I_15450 (I264551,I264432,I264517);
nand I_15451 (I264568,I45115,I45118);
nor I_15452 (I264585,I264568,I45121);
nor I_15453 (I264602,I264568,I264585);
not I_15454 (I264619,I264585);
nor I_15455 (I264390,I264619,I264534);
or I_15456 (I264375,I264432,I264619);
nor I_15457 (I264664,I264432,I264585);
nor I_15458 (I264369,I264568,I264664);
nor I_15459 (I264695,I264602,I264664);
nor I_15460 (I264372,I264517,I264695);
nand I_15461 (I264726,I264432,I264585);
nand I_15462 (I264743,I264500,I264726);
DFFARX1 I_15463 (I264743,I1862,I264398,I264378,);
not I_15464 (I264774,I264568);
nor I_15465 (I264387,I264774,I264619);
nand I_15466 (I264384,I264551,I264774);
nor I_15467 (I264819,I264517,I264568);
nand I_15468 (I264381,I264819,I264432);
not I_15469 (I264874,I1869);
or I_15470 (I264891,I68563,I68572);
nor I_15471 (I264908,I264891,I68587);
nor I_15472 (I264925,I68584,I68566);
or I_15473 (I264942,I264925,I68566);
nor I_15474 (I264959,I68563,I68569);
nand I_15475 (I264976,I264959,I264942);
not I_15476 (I264993,I264976);
nand I_15477 (I265010,I264908,I264993);
nor I_15478 (I265027,I264908,I264993);
nand I_15479 (I265044,I68575,I68578);
nor I_15480 (I265061,I265044,I68581);
nor I_15481 (I265078,I265044,I265061);
not I_15482 (I265095,I265061);
nor I_15483 (I264866,I265095,I265010);
or I_15484 (I264851,I264908,I265095);
nor I_15485 (I265140,I264908,I265061);
nor I_15486 (I264845,I265044,I265140);
nor I_15487 (I265171,I265078,I265140);
nor I_15488 (I264848,I264993,I265171);
nand I_15489 (I265202,I264908,I265061);
nand I_15490 (I265219,I264976,I265202);
DFFARX1 I_15491 (I265219,I1862,I264874,I264854,);
not I_15492 (I265250,I265044);
nor I_15493 (I264863,I265250,I265095);
nand I_15494 (I264860,I265027,I265250);
nor I_15495 (I265295,I264993,I265044);
nand I_15496 (I264857,I265295,I264908);
not I_15497 (I265350,I1869);
or I_15498 (I265367,I140004,I139989);
nor I_15499 (I265384,I265367,I139983);
nor I_15500 (I265401,I139980,I140001);
or I_15501 (I265418,I265401,I139998);
nor I_15502 (I265435,I139986,I139983);
nand I_15503 (I265452,I265435,I265418);
not I_15504 (I265469,I265452);
nand I_15505 (I265486,I265384,I265469);
nor I_15506 (I265503,I265384,I265469);
nand I_15507 (I265520,I139992,I139995);
nor I_15508 (I265537,I265520,I139980);
nor I_15509 (I265554,I265520,I265537);
not I_15510 (I265571,I265537);
nor I_15511 (I265342,I265571,I265486);
or I_15512 (I265327,I265384,I265571);
nor I_15513 (I265616,I265384,I265537);
nor I_15514 (I265321,I265520,I265616);
nor I_15515 (I265647,I265554,I265616);
nor I_15516 (I265324,I265469,I265647);
nand I_15517 (I265678,I265384,I265537);
nand I_15518 (I265695,I265452,I265678);
DFFARX1 I_15519 (I265695,I1862,I265350,I265330,);
not I_15520 (I265726,I265520);
nor I_15521 (I265339,I265726,I265571);
nand I_15522 (I265336,I265503,I265726);
nor I_15523 (I265771,I265469,I265520);
nand I_15524 (I265333,I265771,I265384);
not I_15525 (I265826,I1869);
or I_15526 (I265843,I96103,I96112);
nor I_15527 (I265860,I265843,I96127);
nor I_15528 (I265877,I96124,I96106);
or I_15529 (I265894,I265877,I96106);
nor I_15530 (I265911,I96103,I96109);
nand I_15531 (I265928,I265911,I265894);
not I_15532 (I265945,I265928);
nand I_15533 (I265962,I265860,I265945);
nor I_15534 (I265979,I265860,I265945);
nand I_15535 (I265996,I96115,I96118);
nor I_15536 (I266013,I265996,I96121);
nor I_15537 (I266030,I265996,I266013);
not I_15538 (I266047,I266013);
nor I_15539 (I265818,I266047,I265962);
or I_15540 (I265803,I265860,I266047);
nor I_15541 (I266092,I265860,I266013);
nor I_15542 (I265797,I265996,I266092);
nor I_15543 (I266123,I266030,I266092);
nor I_15544 (I265800,I265945,I266123);
nand I_15545 (I266154,I265860,I266013);
nand I_15546 (I266171,I265928,I266154);
DFFARX1 I_15547 (I266171,I1862,I265826,I265806,);
not I_15548 (I266202,I265996);
nor I_15549 (I265815,I266202,I266047);
nand I_15550 (I265812,I265979,I266202);
nor I_15551 (I266247,I265945,I265996);
nand I_15552 (I265809,I266247,I265860);
not I_15553 (I266302,I1869);
or I_15554 (I266319,I84883,I84892);
nor I_15555 (I266336,I266319,I84907);
nor I_15556 (I266353,I84904,I84886);
or I_15557 (I266370,I266353,I84886);
nor I_15558 (I266387,I84883,I84889);
nand I_15559 (I266404,I266387,I266370);
not I_15560 (I266421,I266404);
nand I_15561 (I266438,I266336,I266421);
nor I_15562 (I266455,I266336,I266421);
nand I_15563 (I266472,I84895,I84898);
nor I_15564 (I266489,I266472,I84901);
nor I_15565 (I266506,I266472,I266489);
not I_15566 (I266523,I266489);
nor I_15567 (I266294,I266523,I266438);
or I_15568 (I266279,I266336,I266523);
nor I_15569 (I266568,I266336,I266489);
nor I_15570 (I266273,I266472,I266568);
nor I_15571 (I266599,I266506,I266568);
nor I_15572 (I266276,I266421,I266599);
nand I_15573 (I266630,I266336,I266489);
nand I_15574 (I266647,I266404,I266630);
DFFARX1 I_15575 (I266647,I1862,I266302,I266282,);
not I_15576 (I266678,I266472);
nor I_15577 (I266291,I266678,I266523);
nand I_15578 (I266288,I266455,I266678);
nor I_15579 (I266723,I266421,I266472);
nand I_15580 (I266285,I266723,I266336);
not I_15581 (I266778,I1869);
or I_15582 (I266795,I17053,I17062);
nor I_15583 (I266812,I266795,I17077);
nor I_15584 (I266829,I17074,I17056);
or I_15585 (I266846,I266829,I17056);
nor I_15586 (I266863,I17053,I17059);
nand I_15587 (I266880,I266863,I266846);
not I_15588 (I266897,I266880);
nand I_15589 (I266914,I266812,I266897);
nor I_15590 (I266931,I266812,I266897);
nand I_15591 (I266948,I17065,I17068);
nor I_15592 (I266965,I266948,I17071);
nor I_15593 (I266982,I266948,I266965);
not I_15594 (I266999,I266965);
nor I_15595 (I266770,I266999,I266914);
or I_15596 (I266755,I266812,I266999);
nor I_15597 (I267044,I266812,I266965);
nor I_15598 (I266749,I266948,I267044);
nor I_15599 (I267075,I266982,I267044);
nor I_15600 (I266752,I266897,I267075);
nand I_15601 (I267106,I266812,I266965);
nand I_15602 (I267123,I266880,I267106);
DFFARX1 I_15603 (I267123,I1862,I266778,I266758,);
not I_15604 (I267154,I266948);
nor I_15605 (I266767,I267154,I266999);
nand I_15606 (I266764,I266931,I267154);
nor I_15607 (I267199,I266897,I266948);
nand I_15608 (I266761,I267199,I266812);
not I_15609 (I267254,I1869);
or I_15610 (I267271,I15523,I15532);
nor I_15611 (I267288,I267271,I15547);
nor I_15612 (I267305,I15544,I15526);
or I_15613 (I267322,I267305,I15526);
nor I_15614 (I267339,I15523,I15529);
nand I_15615 (I267356,I267339,I267322);
not I_15616 (I267373,I267356);
nand I_15617 (I267390,I267288,I267373);
nor I_15618 (I267407,I267288,I267373);
nand I_15619 (I267424,I15535,I15538);
nor I_15620 (I267441,I267424,I15541);
nor I_15621 (I267458,I267424,I267441);
not I_15622 (I267475,I267441);
nor I_15623 (I267246,I267475,I267390);
or I_15624 (I267231,I267288,I267475);
nor I_15625 (I267520,I267288,I267441);
nor I_15626 (I267225,I267424,I267520);
nor I_15627 (I267551,I267458,I267520);
nor I_15628 (I267228,I267373,I267551);
nand I_15629 (I267582,I267288,I267441);
nand I_15630 (I267599,I267356,I267582);
DFFARX1 I_15631 (I267599,I1862,I267254,I267234,);
not I_15632 (I267630,I267424);
nor I_15633 (I267243,I267630,I267475);
nand I_15634 (I267240,I267407,I267630);
nor I_15635 (I267675,I267373,I267424);
nand I_15636 (I267237,I267675,I267288);
not I_15637 (I267730,I1869);
or I_15638 (I267747,I293068,I293065);
nor I_15639 (I267764,I267747,I293074);
nor I_15640 (I267781,I293086,I293071);
or I_15641 (I267798,I267781,I293065);
nor I_15642 (I267815,I293077,I293068);
nand I_15643 (I267832,I267815,I267798);
not I_15644 (I267849,I267832);
nand I_15645 (I267866,I267764,I267849);
nor I_15646 (I267883,I267764,I267849);
nand I_15647 (I267900,I293071,I293083);
nor I_15648 (I267917,I267900,I293080);
nor I_15649 (I267934,I267900,I267917);
not I_15650 (I267951,I267917);
nor I_15651 (I267722,I267951,I267866);
or I_15652 (I267707,I267764,I267951);
nor I_15653 (I267996,I267764,I267917);
nor I_15654 (I267701,I267900,I267996);
nor I_15655 (I268027,I267934,I267996);
nor I_15656 (I267704,I267849,I268027);
nand I_15657 (I268058,I267764,I267917);
nand I_15658 (I268075,I267832,I268058);
DFFARX1 I_15659 (I268075,I1862,I267730,I267710,);
not I_15660 (I268106,I267900);
nor I_15661 (I267719,I268106,I267951);
nand I_15662 (I267716,I267883,I268106);
nor I_15663 (I268151,I267849,I267900);
nand I_15664 (I267713,I268151,I267764);
not I_15665 (I268206,I1869);
or I_15666 (I268223,I59893,I59902);
nor I_15667 (I268240,I268223,I59917);
nor I_15668 (I268257,I59914,I59896);
or I_15669 (I268274,I268257,I59896);
nor I_15670 (I268291,I59893,I59899);
nand I_15671 (I268308,I268291,I268274);
not I_15672 (I268325,I268308);
nand I_15673 (I268342,I268240,I268325);
nor I_15674 (I268359,I268240,I268325);
nand I_15675 (I268376,I59905,I59908);
nor I_15676 (I268393,I268376,I59911);
nor I_15677 (I268410,I268376,I268393);
not I_15678 (I268427,I268393);
nor I_15679 (I268198,I268427,I268342);
or I_15680 (I268183,I268240,I268427);
nor I_15681 (I268472,I268240,I268393);
nor I_15682 (I268177,I268376,I268472);
nor I_15683 (I268503,I268410,I268472);
nor I_15684 (I268180,I268325,I268503);
nand I_15685 (I268534,I268240,I268393);
nand I_15686 (I268551,I268308,I268534);
DFFARX1 I_15687 (I268551,I1862,I268206,I268186,);
not I_15688 (I268582,I268376);
nor I_15689 (I268195,I268582,I268427);
nand I_15690 (I268192,I268359,I268582);
nor I_15691 (I268627,I268325,I268376);
nand I_15692 (I268189,I268627,I268240);
not I_15693 (I268682,I1869);
or I_15694 (I268699,I343657,I343678);
nor I_15695 (I268716,I268699,I343663);
nor I_15696 (I268733,I343657,I343675);
or I_15697 (I268750,I268733,I343666);
nor I_15698 (I268767,I343660,I343660);
nand I_15699 (I268784,I268767,I268750);
not I_15700 (I268801,I268784);
nand I_15701 (I268818,I268716,I268801);
nor I_15702 (I268835,I268716,I268801);
nand I_15703 (I268852,I343669,I343672);
nor I_15704 (I268869,I268852,I343663);
nor I_15705 (I268886,I268852,I268869);
not I_15706 (I268903,I268869);
nor I_15707 (I268674,I268903,I268818);
or I_15708 (I268659,I268716,I268903);
nor I_15709 (I268948,I268716,I268869);
nor I_15710 (I268653,I268852,I268948);
nor I_15711 (I268979,I268886,I268948);
nor I_15712 (I268656,I268801,I268979);
nand I_15713 (I269010,I268716,I268869);
nand I_15714 (I269027,I268784,I269010);
DFFARX1 I_15715 (I269027,I1862,I268682,I268662,);
not I_15716 (I269058,I268852);
nor I_15717 (I268671,I269058,I268903);
nand I_15718 (I268668,I268835,I269058);
nor I_15719 (I269103,I268801,I268852);
nand I_15720 (I268665,I269103,I268716);
not I_15721 (I269158,I1869);
or I_15722 (I269175,I30823,I30832);
nor I_15723 (I269192,I269175,I30847);
nor I_15724 (I269209,I30844,I30826);
or I_15725 (I269226,I269209,I30826);
nor I_15726 (I269243,I30823,I30829);
nand I_15727 (I269260,I269243,I269226);
not I_15728 (I269277,I269260);
nand I_15729 (I269294,I269192,I269277);
nor I_15730 (I269311,I269192,I269277);
nand I_15731 (I269328,I30835,I30838);
nor I_15732 (I269345,I269328,I30841);
nor I_15733 (I269362,I269328,I269345);
not I_15734 (I269379,I269345);
nor I_15735 (I269150,I269379,I269294);
or I_15736 (I269135,I269192,I269379);
nor I_15737 (I269424,I269192,I269345);
nor I_15738 (I269129,I269328,I269424);
nor I_15739 (I269455,I269362,I269424);
nor I_15740 (I269132,I269277,I269455);
nand I_15741 (I269486,I269192,I269345);
nand I_15742 (I269503,I269260,I269486);
DFFARX1 I_15743 (I269503,I1862,I269158,I269138,);
not I_15744 (I269534,I269328);
nor I_15745 (I269147,I269534,I269379);
nand I_15746 (I269144,I269311,I269534);
nor I_15747 (I269579,I269277,I269328);
nand I_15748 (I269141,I269579,I269192);
not I_15749 (I269634,I1869);
or I_15750 (I269651,I86923,I86932);
nor I_15751 (I269668,I269651,I86947);
nor I_15752 (I269685,I86944,I86926);
or I_15753 (I269702,I269685,I86926);
nor I_15754 (I269719,I86923,I86929);
nand I_15755 (I269736,I269719,I269702);
not I_15756 (I269753,I269736);
nand I_15757 (I269770,I269668,I269753);
nor I_15758 (I269787,I269668,I269753);
nand I_15759 (I269804,I86935,I86938);
nor I_15760 (I269821,I269804,I86941);
nor I_15761 (I269838,I269804,I269821);
not I_15762 (I269855,I269821);
nor I_15763 (I269626,I269855,I269770);
or I_15764 (I269611,I269668,I269855);
nor I_15765 (I269900,I269668,I269821);
nor I_15766 (I269605,I269804,I269900);
nor I_15767 (I269931,I269838,I269900);
nor I_15768 (I269608,I269753,I269931);
nand I_15769 (I269962,I269668,I269821);
nand I_15770 (I269979,I269736,I269962);
DFFARX1 I_15771 (I269979,I1862,I269634,I269614,);
not I_15772 (I270010,I269804);
nor I_15773 (I269623,I270010,I269855);
nand I_15774 (I269620,I269787,I270010);
nor I_15775 (I270055,I269753,I269804);
nand I_15776 (I269617,I270055,I269668);
not I_15777 (I270110,I1869);
or I_15778 (I270127,I365471,I365474);
nor I_15779 (I270144,I270127,I365471);
nor I_15780 (I270161,I365468,I365486);
or I_15781 (I270178,I270161,I365474);
nor I_15782 (I270195,I365477,I365468);
nand I_15783 (I270212,I270195,I270178);
not I_15784 (I270229,I270212);
nand I_15785 (I270246,I270144,I270229);
nor I_15786 (I270263,I270144,I270229);
nand I_15787 (I270280,I365483,I365480);
nor I_15788 (I270297,I270280,I365477);
nor I_15789 (I270314,I270280,I270297);
not I_15790 (I270331,I270297);
nor I_15791 (I270102,I270331,I270246);
or I_15792 (I270087,I270144,I270331);
nor I_15793 (I270376,I270144,I270297);
nor I_15794 (I270081,I270280,I270376);
nor I_15795 (I270407,I270314,I270376);
nor I_15796 (I270084,I270229,I270407);
nand I_15797 (I270438,I270144,I270297);
nand I_15798 (I270455,I270212,I270438);
DFFARX1 I_15799 (I270455,I1862,I270110,I270090,);
not I_15800 (I270486,I270280);
nor I_15801 (I270099,I270486,I270331);
nand I_15802 (I270096,I270263,I270486);
nor I_15803 (I270531,I270229,I270280);
nand I_15804 (I270093,I270531,I270144);
not I_15805 (I270586,I1869);
or I_15806 (I270603,I44593,I44602);
nor I_15807 (I270620,I270603,I44617);
nor I_15808 (I270637,I44614,I44596);
or I_15809 (I270654,I270637,I44596);
nor I_15810 (I270671,I44593,I44599);
nand I_15811 (I270688,I270671,I270654);
not I_15812 (I270705,I270688);
nand I_15813 (I270722,I270620,I270705);
nor I_15814 (I270739,I270620,I270705);
nand I_15815 (I270756,I44605,I44608);
nor I_15816 (I270773,I270756,I44611);
nor I_15817 (I270790,I270756,I270773);
not I_15818 (I270807,I270773);
nor I_15819 (I270578,I270807,I270722);
or I_15820 (I270563,I270620,I270807);
nor I_15821 (I270852,I270620,I270773);
nor I_15822 (I270557,I270756,I270852);
nor I_15823 (I270883,I270790,I270852);
nor I_15824 (I270560,I270705,I270883);
nand I_15825 (I270914,I270620,I270773);
nand I_15826 (I270931,I270688,I270914);
DFFARX1 I_15827 (I270931,I1862,I270586,I270566,);
not I_15828 (I270962,I270756);
nor I_15829 (I270575,I270962,I270807);
nand I_15830 (I270572,I270739,I270962);
nor I_15831 (I271007,I270705,I270756);
nand I_15832 (I270569,I271007,I270620);
not I_15833 (I271062,I1869);
or I_15834 (I271079,I385361,I385364);
nor I_15835 (I271096,I271079,I385361);
nor I_15836 (I271113,I385358,I385376);
or I_15837 (I271130,I271113,I385364);
nor I_15838 (I271147,I385367,I385358);
nand I_15839 (I271164,I271147,I271130);
not I_15840 (I271181,I271164);
nand I_15841 (I271198,I271096,I271181);
nor I_15842 (I271215,I271096,I271181);
nand I_15843 (I271232,I385373,I385370);
nor I_15844 (I271249,I271232,I385367);
nor I_15845 (I271266,I271232,I271249);
not I_15846 (I271283,I271249);
nor I_15847 (I271054,I271283,I271198);
or I_15848 (I271039,I271096,I271283);
nor I_15849 (I271328,I271096,I271249);
nor I_15850 (I271033,I271232,I271328);
nor I_15851 (I271359,I271266,I271328);
nor I_15852 (I271036,I271181,I271359);
nand I_15853 (I271390,I271096,I271249);
nand I_15854 (I271407,I271164,I271390);
DFFARX1 I_15855 (I271407,I1862,I271062,I271042,);
not I_15856 (I271438,I271232);
nor I_15857 (I271051,I271438,I271283);
nand I_15858 (I271048,I271215,I271438);
nor I_15859 (I271483,I271181,I271232);
nand I_15860 (I271045,I271483,I271096);
not I_15861 (I271538,I1869);
or I_15862 (I271555,I112426,I112423);
nor I_15863 (I271572,I271555,I112423);
nor I_15864 (I271589,I112432,I112429);
or I_15865 (I271606,I271589,I112438);
nor I_15866 (I271623,I112441,I112426);
nand I_15867 (I271640,I271623,I271606);
not I_15868 (I271657,I271640);
nand I_15869 (I271674,I271572,I271657);
nor I_15870 (I271691,I271572,I271657);
nand I_15871 (I271708,I112429,I112435);
nor I_15872 (I271725,I271708,I112432);
nor I_15873 (I271742,I271708,I271725);
not I_15874 (I271759,I271725);
nor I_15875 (I271530,I271759,I271674);
or I_15876 (I271515,I271572,I271759);
nor I_15877 (I271804,I271572,I271725);
nor I_15878 (I271509,I271708,I271804);
nor I_15879 (I271835,I271742,I271804);
nor I_15880 (I271512,I271657,I271835);
nand I_15881 (I271866,I271572,I271725);
nand I_15882 (I271883,I271640,I271866);
DFFARX1 I_15883 (I271883,I1862,I271538,I271518,);
not I_15884 (I271914,I271708);
nor I_15885 (I271527,I271914,I271759);
nand I_15886 (I271524,I271691,I271914);
nor I_15887 (I271959,I271657,I271708);
nand I_15888 (I271521,I271959,I271572);
not I_15889 (I272014,I1869);
or I_15890 (I272031,I188488,I188473);
nor I_15891 (I272048,I272031,I188467);
nor I_15892 (I272065,I188464,I188485);
or I_15893 (I272082,I272065,I188482);
nor I_15894 (I272099,I188470,I188467);
nand I_15895 (I272116,I272099,I272082);
not I_15896 (I272133,I272116);
nand I_15897 (I272150,I272048,I272133);
nor I_15898 (I272167,I272048,I272133);
nand I_15899 (I272184,I188476,I188479);
nor I_15900 (I272201,I272184,I188464);
nor I_15901 (I272218,I272184,I272201);
not I_15902 (I272235,I272201);
nor I_15903 (I272006,I272235,I272150);
or I_15904 (I271991,I272048,I272235);
nor I_15905 (I272280,I272048,I272201);
nor I_15906 (I271985,I272184,I272280);
nor I_15907 (I272311,I272218,I272280);
nor I_15908 (I271988,I272133,I272311);
nand I_15909 (I272342,I272048,I272201);
nand I_15910 (I272359,I272116,I272342);
DFFARX1 I_15911 (I272359,I1862,I272014,I271994,);
not I_15912 (I272390,I272184);
nor I_15913 (I272003,I272390,I272235);
nand I_15914 (I272000,I272167,I272390);
nor I_15915 (I272435,I272133,I272184);
nand I_15916 (I271997,I272435,I272048);
not I_15917 (I272490,I1869);
or I_15918 (I272507,I132626,I132611);
nor I_15919 (I272524,I272507,I132605);
nor I_15920 (I272541,I132602,I132623);
or I_15921 (I272558,I272541,I132620);
nor I_15922 (I272575,I132608,I132605);
nand I_15923 (I272592,I272575,I272558);
not I_15924 (I272609,I272592);
nand I_15925 (I272626,I272524,I272609);
nor I_15926 (I272643,I272524,I272609);
nand I_15927 (I272660,I132614,I132617);
nor I_15928 (I272677,I272660,I132602);
nor I_15929 (I272694,I272660,I272677);
not I_15930 (I272711,I272677);
nor I_15931 (I272482,I272711,I272626);
or I_15932 (I272467,I272524,I272711);
nor I_15933 (I272756,I272524,I272677);
nor I_15934 (I272461,I272660,I272756);
nor I_15935 (I272787,I272694,I272756);
nor I_15936 (I272464,I272609,I272787);
nand I_15937 (I272818,I272524,I272677);
nand I_15938 (I272835,I272592,I272818);
DFFARX1 I_15939 (I272835,I1862,I272490,I272470,);
not I_15940 (I272866,I272660);
nor I_15941 (I272479,I272866,I272711);
nand I_15942 (I272476,I272643,I272866);
nor I_15943 (I272911,I272609,I272660);
nand I_15944 (I272473,I272911,I272524);
not I_15945 (I272966,I1869);
or I_15946 (I272983,I194285,I194270);
nor I_15947 (I273000,I272983,I194264);
nor I_15948 (I273017,I194261,I194282);
or I_15949 (I273034,I273017,I194279);
nor I_15950 (I273051,I194267,I194264);
nand I_15951 (I273068,I273051,I273034);
not I_15952 (I273085,I273068);
nand I_15953 (I273102,I273000,I273085);
nor I_15954 (I273119,I273000,I273085);
nand I_15955 (I273136,I194273,I194276);
nor I_15956 (I273153,I273136,I194261);
nor I_15957 (I273170,I273136,I273153);
not I_15958 (I273187,I273153);
nor I_15959 (I272958,I273187,I273102);
or I_15960 (I272943,I273000,I273187);
nor I_15961 (I273232,I273000,I273153);
nor I_15962 (I272937,I273136,I273232);
nor I_15963 (I273263,I273170,I273232);
nor I_15964 (I272940,I273085,I273263);
nand I_15965 (I273294,I273000,I273153);
nand I_15966 (I273311,I273068,I273294);
DFFARX1 I_15967 (I273311,I1862,I272966,I272946,);
not I_15968 (I273342,I273136);
nor I_15969 (I272955,I273342,I273187);
nand I_15970 (I272952,I273119,I273342);
nor I_15971 (I273387,I273085,I273136);
nand I_15972 (I272949,I273387,I273000);
not I_15973 (I273442,I1869);
or I_15974 (I273459,I310983,I311004);
nor I_15975 (I273476,I273459,I310989);
nor I_15976 (I273493,I310983,I311001);
or I_15977 (I273510,I273493,I310992);
nor I_15978 (I273527,I310986,I310986);
nand I_15979 (I273544,I273527,I273510);
not I_15980 (I273561,I273544);
nand I_15981 (I273578,I273476,I273561);
nor I_15982 (I273595,I273476,I273561);
nand I_15983 (I273612,I310995,I310998);
nor I_15984 (I273629,I273612,I310989);
nor I_15985 (I273646,I273612,I273629);
not I_15986 (I273663,I273629);
nor I_15987 (I273434,I273663,I273578);
or I_15988 (I273419,I273476,I273663);
nor I_15989 (I273708,I273476,I273629);
nor I_15990 (I273413,I273612,I273708);
nor I_15991 (I273739,I273646,I273708);
nor I_15992 (I273416,I273561,I273739);
nand I_15993 (I273770,I273476,I273629);
nand I_15994 (I273787,I273544,I273770);
DFFARX1 I_15995 (I273787,I1862,I273442,I273422,);
not I_15996 (I273818,I273612);
nor I_15997 (I273431,I273818,I273663);
nand I_15998 (I273428,I273595,I273818);
nor I_15999 (I273863,I273561,I273612);
nand I_16000 (I273425,I273863,I273476);
not I_16001 (I273918,I1869);
or I_16002 (I273935,I401273,I401276);
nor I_16003 (I273952,I273935,I401273);
nor I_16004 (I273969,I401270,I401288);
or I_16005 (I273986,I273969,I401276);
nor I_16006 (I274003,I401279,I401270);
nand I_16007 (I274020,I274003,I273986);
not I_16008 (I274037,I274020);
nand I_16009 (I274054,I273952,I274037);
nor I_16010 (I274071,I273952,I274037);
nand I_16011 (I274088,I401285,I401282);
nor I_16012 (I274105,I274088,I401279);
nor I_16013 (I274122,I274088,I274105);
not I_16014 (I274139,I274105);
nor I_16015 (I273910,I274139,I274054);
or I_16016 (I273895,I273952,I274139);
nor I_16017 (I274184,I273952,I274105);
nor I_16018 (I273889,I274088,I274184);
nor I_16019 (I274215,I274122,I274184);
nor I_16020 (I273892,I274037,I274215);
nand I_16021 (I274246,I273952,I274105);
nand I_16022 (I274263,I274020,I274246);
DFFARX1 I_16023 (I274263,I1862,I273918,I273898,);
not I_16024 (I274294,I274088);
nor I_16025 (I273907,I274294,I274139);
nand I_16026 (I273904,I274071,I274294);
nor I_16027 (I274339,I274037,I274088);
nand I_16028 (I273901,I274339,I273952);
not I_16029 (I274394,I1869);
or I_16030 (I274411,I146855,I146840);
nor I_16031 (I274428,I274411,I146834);
nor I_16032 (I274445,I146831,I146852);
or I_16033 (I274462,I274445,I146849);
nor I_16034 (I274479,I146837,I146834);
nand I_16035 (I274496,I274479,I274462);
not I_16036 (I274513,I274496);
nand I_16037 (I274530,I274428,I274513);
nor I_16038 (I274547,I274428,I274513);
nand I_16039 (I274564,I146843,I146846);
nor I_16040 (I274581,I274564,I146831);
nor I_16041 (I274598,I274564,I274581);
not I_16042 (I274615,I274581);
nor I_16043 (I274386,I274615,I274530);
or I_16044 (I274371,I274428,I274615);
nor I_16045 (I274660,I274428,I274581);
nor I_16046 (I274365,I274564,I274660);
nor I_16047 (I274691,I274598,I274660);
nor I_16048 (I274368,I274513,I274691);
nand I_16049 (I274722,I274428,I274581);
nand I_16050 (I274739,I274496,I274722);
DFFARX1 I_16051 (I274739,I1862,I274394,I274374,);
not I_16052 (I274770,I274564);
nor I_16053 (I274383,I274770,I274615);
nand I_16054 (I274380,I274547,I274770);
nor I_16055 (I274815,I274513,I274564);
nand I_16056 (I274377,I274815,I274428);
not I_16057 (I274870,I1869);
or I_16058 (I274887,I187961,I187946);
nor I_16059 (I274904,I274887,I187940);
nor I_16060 (I274921,I187937,I187958);
or I_16061 (I274938,I274921,I187955);
nor I_16062 (I274955,I187943,I187940);
nand I_16063 (I274972,I274955,I274938);
not I_16064 (I274989,I274972);
nand I_16065 (I275006,I274904,I274989);
nor I_16066 (I275023,I274904,I274989);
nand I_16067 (I275040,I187949,I187952);
nor I_16068 (I275057,I275040,I187937);
nor I_16069 (I275074,I275040,I275057);
not I_16070 (I275091,I275057);
nor I_16071 (I274862,I275091,I275006);
or I_16072 (I274847,I274904,I275091);
nor I_16073 (I275136,I274904,I275057);
nor I_16074 (I274841,I275040,I275136);
nor I_16075 (I275167,I275074,I275136);
nor I_16076 (I274844,I274989,I275167);
nand I_16077 (I275198,I274904,I275057);
nand I_16078 (I275215,I274972,I275198);
DFFARX1 I_16079 (I275215,I1862,I274870,I274850,);
not I_16080 (I275246,I275040);
nor I_16081 (I274859,I275246,I275091);
nand I_16082 (I274856,I275023,I275246);
nor I_16083 (I275291,I274989,I275040);
nand I_16084 (I274853,I275291,I274904);
not I_16085 (I275346,I1869);
or I_16086 (I275363,I5582,I5570);
nor I_16087 (I275380,I275363,I5564);
nor I_16088 (I275397,I5567,I5576);
or I_16089 (I275414,I275397,I5579);
nor I_16090 (I275431,I5561,I5564);
nand I_16091 (I275448,I275431,I275414);
not I_16092 (I275465,I275448);
nand I_16093 (I275482,I275380,I275465);
nor I_16094 (I275499,I275380,I275465);
nand I_16095 (I275516,I5567,I5573);
nor I_16096 (I275533,I275516,I5561);
nor I_16097 (I275550,I275516,I275533);
not I_16098 (I275567,I275533);
nor I_16099 (I275338,I275567,I275482);
or I_16100 (I275323,I275380,I275567);
nor I_16101 (I275612,I275380,I275533);
nor I_16102 (I275317,I275516,I275612);
nor I_16103 (I275643,I275550,I275612);
nor I_16104 (I275320,I275465,I275643);
nand I_16105 (I275674,I275380,I275533);
nand I_16106 (I275691,I275448,I275674);
DFFARX1 I_16107 (I275691,I1862,I275346,I275326,);
not I_16108 (I275722,I275516);
nor I_16109 (I275335,I275722,I275567);
nand I_16110 (I275332,I275499,I275722);
nor I_16111 (I275767,I275465,I275516);
nand I_16112 (I275329,I275767,I275380);
not I_16113 (I275822,I1869);
or I_16114 (I275839,I32353,I32362);
nor I_16115 (I275856,I275839,I32377);
nor I_16116 (I275873,I32374,I32356);
or I_16117 (I275890,I275873,I32356);
nor I_16118 (I275907,I32353,I32359);
nand I_16119 (I275924,I275907,I275890);
not I_16120 (I275941,I275924);
nand I_16121 (I275958,I275856,I275941);
nor I_16122 (I275975,I275856,I275941);
nand I_16123 (I275992,I32365,I32368);
nor I_16124 (I276009,I275992,I32371);
nor I_16125 (I276026,I275992,I276009);
not I_16126 (I276043,I276009);
nor I_16127 (I275814,I276043,I275958);
or I_16128 (I275799,I275856,I276043);
nor I_16129 (I276088,I275856,I276009);
nor I_16130 (I275793,I275992,I276088);
nor I_16131 (I276119,I276026,I276088);
nor I_16132 (I275796,I275941,I276119);
nand I_16133 (I276150,I275856,I276009);
nand I_16134 (I276167,I275924,I276150);
DFFARX1 I_16135 (I276167,I1862,I275822,I275802,);
not I_16136 (I276198,I275992);
nor I_16137 (I275811,I276198,I276043);
nand I_16138 (I275808,I275975,I276198);
nor I_16139 (I276243,I275941,I275992);
nand I_16140 (I275805,I276243,I275856);
not I_16141 (I276298,I1869);
or I_16142 (I276315,I190069,I190054);
nor I_16143 (I276332,I276315,I190048);
nor I_16144 (I276349,I190045,I190066);
or I_16145 (I276366,I276349,I190063);
nor I_16146 (I276383,I190051,I190048);
nand I_16147 (I276400,I276383,I276366);
not I_16148 (I276417,I276400);
nand I_16149 (I276434,I276332,I276417);
nor I_16150 (I276451,I276332,I276417);
nand I_16151 (I276468,I190057,I190060);
nor I_16152 (I276485,I276468,I190045);
nor I_16153 (I276502,I276468,I276485);
not I_16154 (I276519,I276485);
nor I_16155 (I276290,I276519,I276434);
or I_16156 (I276275,I276332,I276519);
nor I_16157 (I276564,I276332,I276485);
nor I_16158 (I276269,I276468,I276564);
nor I_16159 (I276595,I276502,I276564);
nor I_16160 (I276272,I276417,I276595);
nand I_16161 (I276626,I276332,I276485);
nand I_16162 (I276643,I276400,I276626);
DFFARX1 I_16163 (I276643,I1862,I276298,I276278,);
not I_16164 (I276674,I276468);
nor I_16165 (I276287,I276674,I276519);
nand I_16166 (I276284,I276451,I276674);
nor I_16167 (I276719,I276417,I276468);
nand I_16168 (I276281,I276719,I276332);
not I_16169 (I276774,I1869);
or I_16170 (I276791,I98653,I98662);
nor I_16171 (I276808,I276791,I98677);
nor I_16172 (I276825,I98674,I98656);
or I_16173 (I276842,I276825,I98656);
nor I_16174 (I276859,I98653,I98659);
nand I_16175 (I276876,I276859,I276842);
not I_16176 (I276893,I276876);
nand I_16177 (I276910,I276808,I276893);
nor I_16178 (I276927,I276808,I276893);
nand I_16179 (I276944,I98665,I98668);
nor I_16180 (I276961,I276944,I98671);
nor I_16181 (I276978,I276944,I276961);
not I_16182 (I276995,I276961);
nor I_16183 (I276766,I276995,I276910);
or I_16184 (I276751,I276808,I276995);
nor I_16185 (I277040,I276808,I276961);
nor I_16186 (I276745,I276944,I277040);
nor I_16187 (I277071,I276978,I277040);
nor I_16188 (I276748,I276893,I277071);
nand I_16189 (I277102,I276808,I276961);
nand I_16190 (I277119,I276876,I277102);
DFFARX1 I_16191 (I277119,I1862,I276774,I276754,);
not I_16192 (I277150,I276944);
nor I_16193 (I276763,I277150,I276995);
nand I_16194 (I276760,I276927,I277150);
nor I_16195 (I277195,I276893,I276944);
nand I_16196 (I276757,I277195,I276808);
not I_16197 (I277250,I1869);
or I_16198 (I277267,I53263,I53272);
nor I_16199 (I277284,I277267,I53287);
nor I_16200 (I277301,I53284,I53266);
or I_16201 (I277318,I277301,I53266);
nor I_16202 (I277335,I53263,I53269);
nand I_16203 (I277352,I277335,I277318);
not I_16204 (I277369,I277352);
nand I_16205 (I277386,I277284,I277369);
nor I_16206 (I277403,I277284,I277369);
nand I_16207 (I277420,I53275,I53278);
nor I_16208 (I277437,I277420,I53281);
nor I_16209 (I277454,I277420,I277437);
not I_16210 (I277471,I277437);
nor I_16211 (I277242,I277471,I277386);
or I_16212 (I277227,I277284,I277471);
nor I_16213 (I277516,I277284,I277437);
nor I_16214 (I277221,I277420,I277516);
nor I_16215 (I277547,I277454,I277516);
nor I_16216 (I277224,I277369,I277547);
nand I_16217 (I277578,I277284,I277437);
nand I_16218 (I277595,I277352,I277578);
DFFARX1 I_16219 (I277595,I1862,I277250,I277230,);
not I_16220 (I277626,I277420);
nor I_16221 (I277239,I277626,I277471);
nand I_16222 (I277236,I277403,I277626);
nor I_16223 (I277671,I277369,I277420);
nand I_16224 (I277233,I277671,I277284);
not I_16225 (I277726,I1869);
or I_16226 (I277743,I310456,I310477);
nor I_16227 (I277760,I277743,I310462);
nor I_16228 (I277777,I310456,I310474);
or I_16229 (I277794,I277777,I310465);
nor I_16230 (I277811,I310459,I310459);
nand I_16231 (I277828,I277811,I277794);
not I_16232 (I277845,I277828);
nand I_16233 (I277862,I277760,I277845);
nor I_16234 (I277879,I277760,I277845);
nand I_16235 (I277896,I310468,I310471);
nor I_16236 (I277913,I277896,I310462);
nor I_16237 (I277930,I277896,I277913);
not I_16238 (I277947,I277913);
nor I_16239 (I277718,I277947,I277862);
or I_16240 (I277703,I277760,I277947);
nor I_16241 (I277992,I277760,I277913);
nor I_16242 (I277697,I277896,I277992);
nor I_16243 (I278023,I277930,I277992);
nor I_16244 (I277700,I277845,I278023);
nand I_16245 (I278054,I277760,I277913);
nand I_16246 (I278071,I277828,I278054);
DFFARX1 I_16247 (I278071,I1862,I277726,I277706,);
not I_16248 (I278102,I277896);
nor I_16249 (I277715,I278102,I277947);
nand I_16250 (I277712,I277879,I278102);
nor I_16251 (I278147,I277845,I277896);
nand I_16252 (I277709,I278147,I277760);
not I_16253 (I278202,I1869);
or I_16254 (I278219,I314145,I314166);
nor I_16255 (I278236,I278219,I314151);
nor I_16256 (I278253,I314145,I314163);
or I_16257 (I278270,I278253,I314154);
nor I_16258 (I278287,I314148,I314148);
nand I_16259 (I278304,I278287,I278270);
not I_16260 (I278321,I278304);
nand I_16261 (I278338,I278236,I278321);
nor I_16262 (I278355,I278236,I278321);
nand I_16263 (I278372,I314157,I314160);
nor I_16264 (I278389,I278372,I314151);
nor I_16265 (I278406,I278372,I278389);
not I_16266 (I278423,I278389);
nor I_16267 (I278194,I278423,I278338);
or I_16268 (I278179,I278236,I278423);
nor I_16269 (I278468,I278236,I278389);
nor I_16270 (I278173,I278372,I278468);
nor I_16271 (I278499,I278406,I278468);
nor I_16272 (I278176,I278321,I278499);
nand I_16273 (I278530,I278236,I278389);
nand I_16274 (I278547,I278304,I278530);
DFFARX1 I_16275 (I278547,I1862,I278202,I278182,);
not I_16276 (I278578,I278372);
nor I_16277 (I278191,I278578,I278423);
nand I_16278 (I278188,I278355,I278578);
nor I_16279 (I278623,I278321,I278372);
nand I_16280 (I278185,I278623,I278236);
not I_16281 (I278678,I1869);
or I_16282 (I278695,I403041,I403044);
nor I_16283 (I278712,I278695,I403041);
nor I_16284 (I278729,I403038,I403056);
or I_16285 (I278746,I278729,I403044);
nor I_16286 (I278763,I403047,I403038);
nand I_16287 (I278780,I278763,I278746);
not I_16288 (I278797,I278780);
nand I_16289 (I278814,I278712,I278797);
nor I_16290 (I278831,I278712,I278797);
nand I_16291 (I278848,I403053,I403050);
nor I_16292 (I278865,I278848,I403047);
nor I_16293 (I278882,I278848,I278865);
not I_16294 (I278899,I278865);
nor I_16295 (I278670,I278899,I278814);
or I_16296 (I278655,I278712,I278899);
nor I_16297 (I278944,I278712,I278865);
nor I_16298 (I278649,I278848,I278944);
nor I_16299 (I278975,I278882,I278944);
nor I_16300 (I278652,I278797,I278975);
nand I_16301 (I279006,I278712,I278865);
nand I_16302 (I279023,I278780,I279006);
DFFARX1 I_16303 (I279023,I1862,I278678,I278658,);
not I_16304 (I279054,I278848);
nor I_16305 (I278667,I279054,I278899);
nand I_16306 (I278664,I278831,I279054);
nor I_16307 (I279099,I278797,I278848);
nand I_16308 (I278661,I279099,I278712);
not I_16309 (I279154,I1869);
or I_16310 (I279171,I399505,I399508);
nor I_16311 (I279188,I279171,I399505);
nor I_16312 (I279205,I399502,I399520);
or I_16313 (I279222,I279205,I399508);
nor I_16314 (I279239,I399511,I399502);
nand I_16315 (I279256,I279239,I279222);
not I_16316 (I279273,I279256);
nand I_16317 (I279290,I279188,I279273);
nor I_16318 (I279307,I279188,I279273);
nand I_16319 (I279324,I399517,I399514);
nor I_16320 (I279341,I279324,I399511);
nor I_16321 (I279358,I279324,I279341);
not I_16322 (I279375,I279341);
nor I_16323 (I279146,I279375,I279290);
or I_16324 (I279131,I279188,I279375);
nor I_16325 (I279420,I279188,I279341);
nor I_16326 (I279125,I279324,I279420);
nor I_16327 (I279451,I279358,I279420);
nor I_16328 (I279128,I279273,I279451);
nand I_16329 (I279482,I279188,I279341);
nand I_16330 (I279499,I279256,I279482);
DFFARX1 I_16331 (I279499,I1862,I279154,I279134,);
not I_16332 (I279530,I279324);
nor I_16333 (I279143,I279530,I279375);
nand I_16334 (I279140,I279307,I279530);
nor I_16335 (I279575,I279273,I279324);
nand I_16336 (I279137,I279575,I279188);
not I_16337 (I279630,I1869);
or I_16338 (I279647,I327847,I327868);
nor I_16339 (I279664,I279647,I327853);
nor I_16340 (I279681,I327847,I327865);
or I_16341 (I279698,I279681,I327856);
nor I_16342 (I279715,I327850,I327850);
nand I_16343 (I279732,I279715,I279698);
not I_16344 (I279749,I279732);
nand I_16345 (I279766,I279664,I279749);
nor I_16346 (I279783,I279664,I279749);
nand I_16347 (I279800,I327859,I327862);
nor I_16348 (I279817,I279800,I327853);
nor I_16349 (I279834,I279800,I279817);
not I_16350 (I279851,I279817);
nor I_16351 (I279622,I279851,I279766);
or I_16352 (I279607,I279664,I279851);
nor I_16353 (I279896,I279664,I279817);
nor I_16354 (I279601,I279800,I279896);
nor I_16355 (I279927,I279834,I279896);
nor I_16356 (I279604,I279749,I279927);
nand I_16357 (I279958,I279664,I279817);
nand I_16358 (I279975,I279732,I279958);
DFFARX1 I_16359 (I279975,I1862,I279630,I279610,);
not I_16360 (I280006,I279800);
nor I_16361 (I279619,I280006,I279851);
nand I_16362 (I279616,I279783,I280006);
nor I_16363 (I280051,I279749,I279800);
nand I_16364 (I279613,I280051,I279664);
not I_16365 (I280106,I1869);
or I_16366 (I280123,I387571,I387574);
nor I_16367 (I280140,I280123,I387571);
nor I_16368 (I280157,I387568,I387586);
or I_16369 (I280174,I280157,I387574);
nor I_16370 (I280191,I387577,I387568);
nand I_16371 (I280208,I280191,I280174);
not I_16372 (I280225,I280208);
nand I_16373 (I280242,I280140,I280225);
nor I_16374 (I280259,I280140,I280225);
nand I_16375 (I280276,I387583,I387580);
nor I_16376 (I280293,I280276,I387577);
nor I_16377 (I280310,I280276,I280293);
not I_16378 (I280327,I280293);
nor I_16379 (I280098,I280327,I280242);
or I_16380 (I280083,I280140,I280327);
nor I_16381 (I280372,I280140,I280293);
nor I_16382 (I280077,I280276,I280372);
nor I_16383 (I280403,I280310,I280372);
nor I_16384 (I280080,I280225,I280403);
nand I_16385 (I280434,I280140,I280293);
nand I_16386 (I280451,I280208,I280434);
DFFARX1 I_16387 (I280451,I1862,I280106,I280086,);
not I_16388 (I280482,I280276);
nor I_16389 (I280095,I280482,I280327);
nand I_16390 (I280092,I280259,I280482);
nor I_16391 (I280527,I280225,I280276);
nand I_16392 (I280089,I280527,I280140);
not I_16393 (I280582,I1869);
or I_16394 (I280599,I9271,I9259);
nor I_16395 (I280616,I280599,I9253);
nor I_16396 (I280633,I9256,I9265);
or I_16397 (I280650,I280633,I9268);
nor I_16398 (I280667,I9250,I9253);
nand I_16399 (I280684,I280667,I280650);
not I_16400 (I280701,I280684);
nand I_16401 (I280718,I280616,I280701);
nor I_16402 (I280735,I280616,I280701);
nand I_16403 (I280752,I9256,I9262);
nor I_16404 (I280769,I280752,I9250);
nor I_16405 (I280786,I280752,I280769);
not I_16406 (I280803,I280769);
nor I_16407 (I280574,I280803,I280718);
or I_16408 (I280559,I280616,I280803);
nor I_16409 (I280848,I280616,I280769);
nor I_16410 (I280553,I280752,I280848);
nor I_16411 (I280879,I280786,I280848);
nor I_16412 (I280556,I280701,I280879);
nand I_16413 (I280910,I280616,I280769);
nand I_16414 (I280927,I280684,I280910);
DFFARX1 I_16415 (I280927,I1862,I280582,I280562,);
not I_16416 (I280958,I280752);
nor I_16417 (I280571,I280958,I280803);
nand I_16418 (I280568,I280735,I280958);
nor I_16419 (I281003,I280701,I280752);
nand I_16420 (I280565,I281003,I280616);
not I_16421 (I281058,I1869);
or I_16422 (I281075,I407903,I407906);
nor I_16423 (I281092,I281075,I407903);
nor I_16424 (I281109,I407900,I407918);
or I_16425 (I281126,I281109,I407906);
nor I_16426 (I281143,I407909,I407900);
nand I_16427 (I281160,I281143,I281126);
not I_16428 (I281177,I281160);
nand I_16429 (I281194,I281092,I281177);
nor I_16430 (I281211,I281092,I281177);
nand I_16431 (I281228,I407915,I407912);
nor I_16432 (I281245,I281228,I407909);
nor I_16433 (I281262,I281228,I281245);
not I_16434 (I281279,I281245);
nor I_16435 (I281050,I281279,I281194);
or I_16436 (I281035,I281092,I281279);
nor I_16437 (I281324,I281092,I281245);
nor I_16438 (I281029,I281228,I281324);
nor I_16439 (I281355,I281262,I281324);
nor I_16440 (I281032,I281177,I281355);
nand I_16441 (I281386,I281092,I281245);
nand I_16442 (I281403,I281160,I281386);
DFFARX1 I_16443 (I281403,I1862,I281058,I281038,);
not I_16444 (I281434,I281228);
nor I_16445 (I281047,I281434,I281279);
nand I_16446 (I281044,I281211,I281434);
nor I_16447 (I281479,I281177,I281228);
nand I_16448 (I281041,I281479,I281092);
not I_16449 (I281534,I1869);
or I_16450 (I281551,I101713,I101722);
nor I_16451 (I281568,I281551,I101737);
nor I_16452 (I281585,I101734,I101716);
or I_16453 (I281602,I281585,I101716);
nor I_16454 (I281619,I101713,I101719);
nand I_16455 (I281636,I281619,I281602);
not I_16456 (I281653,I281636);
nand I_16457 (I281670,I281568,I281653);
nor I_16458 (I281687,I281568,I281653);
nand I_16459 (I281704,I101725,I101728);
nor I_16460 (I281721,I281704,I101731);
nor I_16461 (I281738,I281704,I281721);
not I_16462 (I281755,I281721);
nor I_16463 (I281526,I281755,I281670);
or I_16464 (I281511,I281568,I281755);
nor I_16465 (I281800,I281568,I281721);
nor I_16466 (I281505,I281704,I281800);
nor I_16467 (I281831,I281738,I281800);
nor I_16468 (I281508,I281653,I281831);
nand I_16469 (I281862,I281568,I281721);
nand I_16470 (I281879,I281636,I281862);
DFFARX1 I_16471 (I281879,I1862,I281534,I281514,);
not I_16472 (I281910,I281704);
nor I_16473 (I281523,I281910,I281755);
nand I_16474 (I281520,I281687,I281910);
nor I_16475 (I281955,I281653,I281704);
nand I_16476 (I281517,I281955,I281568);
not I_16477 (I282010,I1869);
or I_16478 (I282027,I388455,I388458);
nor I_16479 (I282044,I282027,I388455);
nor I_16480 (I282061,I388452,I388470);
or I_16481 (I282078,I282061,I388458);
nor I_16482 (I282095,I388461,I388452);
nand I_16483 (I282112,I282095,I282078);
not I_16484 (I282129,I282112);
nand I_16485 (I282146,I282044,I282129);
nor I_16486 (I282163,I282044,I282129);
nand I_16487 (I282180,I388467,I388464);
nor I_16488 (I282197,I282180,I388461);
nor I_16489 (I282214,I282180,I282197);
not I_16490 (I282231,I282197);
nor I_16491 (I282002,I282231,I282146);
or I_16492 (I281987,I282044,I282231);
nor I_16493 (I282276,I282044,I282197);
nor I_16494 (I281981,I282180,I282276);
nor I_16495 (I282307,I282214,I282276);
nor I_16496 (I281984,I282129,I282307);
nand I_16497 (I282338,I282044,I282197);
nand I_16498 (I282355,I282112,I282338);
DFFARX1 I_16499 (I282355,I1862,I282010,I281990,);
not I_16500 (I282386,I282180);
nor I_16501 (I281999,I282386,I282231);
nand I_16502 (I281996,I282163,I282386);
nor I_16503 (I282431,I282129,I282180);
nand I_16504 (I281993,I282431,I282044);
not I_16505 (I282486,I1869);
or I_16506 (I282503,I382709,I382712);
nor I_16507 (I282520,I282503,I382709);
nor I_16508 (I282537,I382706,I382724);
or I_16509 (I282554,I282537,I382712);
nor I_16510 (I282571,I382715,I382706);
nand I_16511 (I282588,I282571,I282554);
not I_16512 (I282605,I282588);
nand I_16513 (I282622,I282520,I282605);
nor I_16514 (I282639,I282520,I282605);
nand I_16515 (I282656,I382721,I382718);
nor I_16516 (I282673,I282656,I382715);
nor I_16517 (I282690,I282656,I282673);
not I_16518 (I282707,I282673);
nor I_16519 (I282478,I282707,I282622);
or I_16520 (I282463,I282520,I282707);
nor I_16521 (I282752,I282520,I282673);
nor I_16522 (I282457,I282656,I282752);
nor I_16523 (I282783,I282690,I282752);
nor I_16524 (I282460,I282605,I282783);
nand I_16525 (I282814,I282520,I282673);
nand I_16526 (I282831,I282588,I282814);
DFFARX1 I_16527 (I282831,I1862,I282486,I282466,);
not I_16528 (I282862,I282656);
nor I_16529 (I282475,I282862,I282707);
nand I_16530 (I282472,I282639,I282862);
nor I_16531 (I282907,I282605,I282656);
nand I_16532 (I282469,I282907,I282520);
not I_16533 (I282962,I1869);
or I_16534 (I282979,I297284,I297281);
nor I_16535 (I282996,I282979,I297290);
nor I_16536 (I283013,I297302,I297287);
or I_16537 (I283030,I283013,I297281);
nor I_16538 (I283047,I297293,I297284);
nand I_16539 (I283064,I283047,I283030);
not I_16540 (I283081,I283064);
nand I_16541 (I283098,I282996,I283081);
nor I_16542 (I283115,I282996,I283081);
nand I_16543 (I283132,I297287,I297299);
nor I_16544 (I283149,I283132,I297296);
nor I_16545 (I283166,I283132,I283149);
not I_16546 (I283183,I283149);
nor I_16547 (I282954,I283183,I283098);
or I_16548 (I282939,I282996,I283183);
nor I_16549 (I283228,I282996,I283149);
nor I_16550 (I282933,I283132,I283228);
nor I_16551 (I283259,I283166,I283228);
nor I_16552 (I282936,I283081,I283259);
nand I_16553 (I283290,I282996,I283149);
nand I_16554 (I283307,I283064,I283290);
DFFARX1 I_16555 (I283307,I1862,I282962,I282942,);
not I_16556 (I283338,I283132);
nor I_16557 (I282951,I283338,I283183);
nand I_16558 (I282948,I283115,I283338);
nor I_16559 (I283383,I283081,I283132);
nand I_16560 (I282945,I283383,I282996);
not I_16561 (I283438,I1869);
or I_16562 (I283455,I29293,I29302);
nor I_16563 (I283472,I283455,I29317);
nor I_16564 (I283489,I29314,I29296);
or I_16565 (I283506,I283489,I29296);
nor I_16566 (I283523,I29293,I29299);
nand I_16567 (I283540,I283523,I283506);
not I_16568 (I283557,I283540);
nand I_16569 (I283574,I283472,I283557);
nor I_16570 (I283591,I283472,I283557);
nand I_16571 (I283608,I29305,I29308);
nor I_16572 (I283625,I283608,I29311);
nor I_16573 (I283642,I283608,I283625);
not I_16574 (I283659,I283625);
nor I_16575 (I283430,I283659,I283574);
or I_16576 (I283415,I283472,I283659);
nor I_16577 (I283704,I283472,I283625);
nor I_16578 (I283409,I283608,I283704);
nor I_16579 (I283735,I283642,I283704);
nor I_16580 (I283412,I283557,I283735);
nand I_16581 (I283766,I283472,I283625);
nand I_16582 (I283783,I283540,I283766);
DFFARX1 I_16583 (I283783,I1862,I283438,I283418,);
not I_16584 (I283814,I283608);
nor I_16585 (I283427,I283814,I283659);
nand I_16586 (I283424,I283591,I283814);
nor I_16587 (I283859,I283557,I283608);
nand I_16588 (I283421,I283859,I283472);
not I_16589 (I283914,I1869);
or I_16590 (I283931,I31843,I31852);
nor I_16591 (I283948,I283931,I31867);
nor I_16592 (I283965,I31864,I31846);
or I_16593 (I283982,I283965,I31846);
nor I_16594 (I283999,I31843,I31849);
nand I_16595 (I284016,I283999,I283982);
not I_16596 (I284033,I284016);
nand I_16597 (I284050,I283948,I284033);
nor I_16598 (I284067,I283948,I284033);
nand I_16599 (I284084,I31855,I31858);
nor I_16600 (I284101,I284084,I31861);
nor I_16601 (I284118,I284084,I284101);
not I_16602 (I284135,I284101);
nor I_16603 (I283906,I284135,I284050);
or I_16604 (I283891,I283948,I284135);
nor I_16605 (I284180,I283948,I284101);
nor I_16606 (I283885,I284084,I284180);
nor I_16607 (I284211,I284118,I284180);
nor I_16608 (I283888,I284033,I284211);
nand I_16609 (I284242,I283948,I284101);
nand I_16610 (I284259,I284016,I284242);
DFFARX1 I_16611 (I284259,I1862,I283914,I283894,);
not I_16612 (I284290,I284084);
nor I_16613 (I283903,I284290,I284135);
nand I_16614 (I283900,I284067,I284290);
nor I_16615 (I284335,I284033,I284084);
nand I_16616 (I283897,I284335,I283948);
not I_16617 (I284390,I1869);
or I_16618 (I284407,I1327,I943);
nor I_16619 (I284424,I284407,I759);
nor I_16620 (I284441,I791,I1855);
or I_16621 (I284458,I284441,I967);
nor I_16622 (I284475,I1823,I767);
nand I_16623 (I284492,I284475,I284458);
not I_16624 (I284509,I284492);
nand I_16625 (I284526,I284424,I284509);
nor I_16626 (I284543,I284424,I284509);
nand I_16627 (I284560,I1567,I1543);
nor I_16628 (I284577,I284560,I1207);
nor I_16629 (I284594,I284560,I284577);
not I_16630 (I284611,I284577);
nor I_16631 (I284382,I284611,I284526);
or I_16632 (I284367,I284424,I284611);
nor I_16633 (I284656,I284424,I284577);
nor I_16634 (I284361,I284560,I284656);
nor I_16635 (I284687,I284594,I284656);
nor I_16636 (I284364,I284509,I284687);
nand I_16637 (I284718,I284424,I284577);
nand I_16638 (I284735,I284492,I284718);
DFFARX1 I_16639 (I284735,I1862,I284390,I284370,);
not I_16640 (I284766,I284560);
nor I_16641 (I284379,I284766,I284611);
nand I_16642 (I284376,I284543,I284766);
nor I_16643 (I284811,I284509,I284560);
nand I_16644 (I284373,I284811,I284424);
not I_16645 (I284866,I1869);
or I_16646 (I284883,I391991,I391994);
nor I_16647 (I284900,I284883,I391991);
nor I_16648 (I284917,I391988,I392006);
or I_16649 (I284934,I284917,I391994);
nor I_16650 (I284951,I391997,I391988);
nand I_16651 (I284968,I284951,I284934);
not I_16652 (I284985,I284968);
nand I_16653 (I285002,I284900,I284985);
nor I_16654 (I285019,I284900,I284985);
nand I_16655 (I285036,I392003,I392000);
nor I_16656 (I285053,I285036,I391997);
nor I_16657 (I285070,I285036,I285053);
not I_16658 (I285087,I285053);
nor I_16659 (I284858,I285087,I285002);
or I_16660 (I284843,I284900,I285087);
nor I_16661 (I285132,I284900,I285053);
nor I_16662 (I284837,I285036,I285132);
nor I_16663 (I285163,I285070,I285132);
nor I_16664 (I284840,I284985,I285163);
nand I_16665 (I285194,I284900,I285053);
nand I_16666 (I285211,I284968,I285194);
DFFARX1 I_16667 (I285211,I1862,I284866,I284846,);
not I_16668 (I285242,I285036);
nor I_16669 (I284855,I285242,I285087);
nand I_16670 (I284852,I285019,I285242);
nor I_16671 (I285287,I284985,I285036);
nand I_16672 (I284849,I285287,I284900);
not I_16673 (I285342,I1869);
or I_16674 (I285359,I174786,I174771);
nor I_16675 (I285376,I285359,I174765);
nor I_16676 (I285393,I174762,I174783);
or I_16677 (I285410,I285393,I174780);
nor I_16678 (I285427,I174768,I174765);
nand I_16679 (I285444,I285427,I285410);
not I_16680 (I285461,I285444);
nand I_16681 (I285478,I285376,I285461);
nor I_16682 (I285495,I285376,I285461);
nand I_16683 (I285512,I174774,I174777);
nor I_16684 (I285529,I285512,I174762);
nor I_16685 (I285546,I285512,I285529);
not I_16686 (I285563,I285529);
nor I_16687 (I285334,I285563,I285478);
or I_16688 (I285319,I285376,I285563);
nor I_16689 (I285608,I285376,I285529);
nor I_16690 (I285313,I285512,I285608);
nor I_16691 (I285639,I285546,I285608);
nor I_16692 (I285316,I285461,I285639);
nand I_16693 (I285670,I285376,I285529);
nand I_16694 (I285687,I285444,I285670);
DFFARX1 I_16695 (I285687,I1862,I285342,I285322,);
not I_16696 (I285718,I285512);
nor I_16697 (I285331,I285718,I285563);
nand I_16698 (I285328,I285495,I285718);
nor I_16699 (I285763,I285461,I285512);
nand I_16700 (I285325,I285763,I285376);
not I_16701 (I285818,I1869);
or I_16702 (I285835,I23683,I23692);
nor I_16703 (I285852,I285835,I23707);
nor I_16704 (I285869,I23704,I23686);
or I_16705 (I285886,I285869,I23686);
nor I_16706 (I285903,I23683,I23689);
nand I_16707 (I285920,I285903,I285886);
not I_16708 (I285937,I285920);
nand I_16709 (I285954,I285852,I285937);
nor I_16710 (I285971,I285852,I285937);
nand I_16711 (I285988,I23695,I23698);
nor I_16712 (I286005,I285988,I23701);
nor I_16713 (I286022,I285988,I286005);
not I_16714 (I286039,I286005);
nor I_16715 (I285810,I286039,I285954);
or I_16716 (I285795,I285852,I286039);
nor I_16717 (I286084,I285852,I286005);
nor I_16718 (I285789,I285988,I286084);
nor I_16719 (I286115,I286022,I286084);
nor I_16720 (I285792,I285937,I286115);
nand I_16721 (I286146,I285852,I286005);
nand I_16722 (I286163,I285920,I286146);
DFFARX1 I_16723 (I286163,I1862,I285818,I285798,);
not I_16724 (I286194,I285988);
nor I_16725 (I285807,I286194,I286039);
nand I_16726 (I285804,I285971,I286194);
nor I_16727 (I286239,I285937,I285988);
nand I_16728 (I285801,I286239,I285852);
not I_16729 (I286294,I1869);
or I_16730 (I286311,I36943,I36952);
nor I_16731 (I286328,I286311,I36967);
nor I_16732 (I286345,I36964,I36946);
or I_16733 (I286362,I286345,I36946);
nor I_16734 (I286379,I36943,I36949);
nand I_16735 (I286396,I286379,I286362);
not I_16736 (I286413,I286396);
nand I_16737 (I286430,I286328,I286413);
nor I_16738 (I286447,I286328,I286413);
nand I_16739 (I286464,I36955,I36958);
nor I_16740 (I286481,I286464,I36961);
nor I_16741 (I286498,I286464,I286481);
not I_16742 (I286515,I286481);
nor I_16743 (I286286,I286515,I286430);
or I_16744 (I286271,I286328,I286515);
nor I_16745 (I286560,I286328,I286481);
nor I_16746 (I286265,I286464,I286560);
nor I_16747 (I286591,I286498,I286560);
nor I_16748 (I286268,I286413,I286591);
nand I_16749 (I286622,I286328,I286481);
nand I_16750 (I286639,I286396,I286622);
DFFARX1 I_16751 (I286639,I1862,I286294,I286274,);
not I_16752 (I286670,I286464);
nor I_16753 (I286283,I286670,I286515);
nand I_16754 (I286280,I286447,I286670);
nor I_16755 (I286715,I286413,I286464);
nand I_16756 (I286277,I286715,I286328);
not I_16757 (I286770,I1869);
or I_16758 (I286787,I29803,I29824);
nand I_16759 (I286804,I29818,I29806);
not I_16760 (I286821,I286804);
nand I_16761 (I286838,I286821,I286787);
not I_16762 (I286855,I286838);
nand I_16763 (I286872,I29809,I29815);
nor I_16764 (I286889,I286872,I29821);
nor I_16765 (I286906,I286838,I286889);
or I_16766 (I286923,I286889,I286855);
nand I_16767 (I286747,I286838,I286889);
nand I_16768 (I286954,I286889,I286855);
and I_16769 (I286971,I286804,I286872);
nor I_16770 (I286988,I286906,I286971);
nor I_16771 (I287005,I29806,I29812);
not I_16772 (I287022,I29827);
nor I_16773 (I287039,I287022,I287005);
nor I_16774 (I286741,I287039,I286804);
nand I_16775 (I287070,I287039,I286923);
nor I_16776 (I286762,I286804,I287070);
nor I_16777 (I286744,I287039,I286988);
not I_16778 (I286756,I287039);
nor I_16779 (I287129,I287039,I29803);
or I_16780 (I287146,I287022,I29803);
nand I_16781 (I287163,I287146,I286954);
DFFARX1 I_16782 (I287163,I1862,I286770,I286750,);
nor I_16783 (I287194,I287022,I29803);
nor I_16784 (I287211,I287039,I287194);
nand I_16785 (I286759,I287211,I286889);
nor I_16786 (I287242,I287022,I286838);
nand I_16787 (I286753,I287242,I287129);
not I_16788 (I287297,I1869);
or I_16789 (I287314,I207270,I207252);
nand I_16790 (I287331,I207264,I207255);
not I_16791 (I287348,I287331);
nand I_16792 (I287365,I287348,I287314);
not I_16793 (I287382,I287365);
nand I_16794 (I287399,I207261,I207252);
nor I_16795 (I287416,I287399,I207249);
nor I_16796 (I287433,I287365,I287416);
or I_16797 (I287450,I287416,I287382);
nand I_16798 (I287274,I287365,I287416);
nand I_16799 (I287481,I287416,I287382);
and I_16800 (I287498,I287331,I287399);
nor I_16801 (I287515,I287433,I287498);
nor I_16802 (I287532,I207267,I207258);
not I_16803 (I287549,I207249);
nor I_16804 (I287566,I287549,I287532);
nor I_16805 (I287268,I287566,I287331);
nand I_16806 (I287597,I287566,I287450);
nor I_16807 (I287289,I287331,I287597);
nor I_16808 (I287271,I287566,I287515);
not I_16809 (I287283,I287566);
nor I_16810 (I287656,I287566,I207255);
or I_16811 (I287673,I287549,I207255);
nand I_16812 (I287690,I287673,I287481);
DFFARX1 I_16813 (I287690,I1862,I287297,I287277,);
nor I_16814 (I287721,I287549,I207255);
nor I_16815 (I287738,I287566,I287721);
nand I_16816 (I287286,I287738,I287416);
nor I_16817 (I287769,I287549,I287365);
nand I_16818 (I287280,I287769,I287656);
not I_16819 (I287824,I1869);
or I_16820 (I287841,I250110,I250092);
nand I_16821 (I287858,I250104,I250095);
not I_16822 (I287875,I287858);
nand I_16823 (I287892,I287875,I287841);
not I_16824 (I287909,I287892);
nand I_16825 (I287926,I250101,I250092);
nor I_16826 (I287943,I287926,I250089);
nor I_16827 (I287960,I287892,I287943);
or I_16828 (I287977,I287943,I287909);
nand I_16829 (I287801,I287892,I287943);
nand I_16830 (I288008,I287943,I287909);
and I_16831 (I288025,I287858,I287926);
nor I_16832 (I288042,I287960,I288025);
nor I_16833 (I288059,I250107,I250098);
not I_16834 (I288076,I250089);
nor I_16835 (I288093,I288076,I288059);
nor I_16836 (I287795,I288093,I287858);
nand I_16837 (I288124,I288093,I287977);
nor I_16838 (I287816,I287858,I288124);
nor I_16839 (I287798,I288093,I288042);
not I_16840 (I287810,I288093);
nor I_16841 (I288183,I288093,I250095);
or I_16842 (I288200,I288076,I250095);
nand I_16843 (I288217,I288200,I288008);
DFFARX1 I_16844 (I288217,I1862,I287824,I287804,);
nor I_16845 (I288248,I288076,I250095);
nor I_16846 (I288265,I288093,I288248);
nand I_16847 (I287813,I288265,I287943);
nor I_16848 (I288296,I288076,I287892);
nand I_16849 (I287807,I288296,I288183);
not I_16850 (I288351,I1869);
or I_16851 (I288368,I337333,I337345);
nand I_16852 (I288385,I337348,I337351);
not I_16853 (I288402,I288385);
nand I_16854 (I288419,I288402,I288368);
not I_16855 (I288436,I288419);
nand I_16856 (I288453,I337333,I337336);
nor I_16857 (I288470,I288453,I337339);
nor I_16858 (I288487,I288419,I288470);
or I_16859 (I288504,I288470,I288436);
nand I_16860 (I288328,I288419,I288470);
nand I_16861 (I288535,I288470,I288436);
and I_16862 (I288552,I288385,I288453);
nor I_16863 (I288569,I288487,I288552);
nor I_16864 (I288586,I337342,I337339);
not I_16865 (I288603,I337354);
nor I_16866 (I288620,I288603,I288586);
nor I_16867 (I288322,I288620,I288385);
nand I_16868 (I288651,I288620,I288504);
nor I_16869 (I288343,I288385,I288651);
nor I_16870 (I288325,I288620,I288569);
not I_16871 (I288337,I288620);
nor I_16872 (I288710,I288620,I337336);
or I_16873 (I288727,I288603,I337336);
nand I_16874 (I288744,I288727,I288535);
DFFARX1 I_16875 (I288744,I1862,I288351,I288331,);
nor I_16876 (I288775,I288603,I337336);
nor I_16877 (I288792,I288620,I288775);
nand I_16878 (I288340,I288792,I288470);
nor I_16879 (I288823,I288603,I288419);
nand I_16880 (I288334,I288823,I288710);
not I_16881 (I288878,I1869);
or I_16882 (I288895,I349981,I349993);
nand I_16883 (I288912,I349996,I349999);
not I_16884 (I288929,I288912);
nand I_16885 (I288946,I288929,I288895);
not I_16886 (I288963,I288946);
nand I_16887 (I288980,I349981,I349984);
nor I_16888 (I288997,I288980,I349987);
nor I_16889 (I289014,I288946,I288997);
or I_16890 (I289031,I288997,I288963);
nand I_16891 (I288855,I288946,I288997);
nand I_16892 (I289062,I288997,I288963);
and I_16893 (I289079,I288912,I288980);
nor I_16894 (I289096,I289014,I289079);
nor I_16895 (I289113,I349990,I349987);
not I_16896 (I289130,I350002);
nor I_16897 (I289147,I289130,I289113);
nor I_16898 (I288849,I289147,I288912);
nand I_16899 (I289178,I289147,I289031);
nor I_16900 (I288870,I288912,I289178);
nor I_16901 (I288852,I289147,I289096);
not I_16902 (I288864,I289147);
nor I_16903 (I289237,I289147,I349984);
or I_16904 (I289254,I289130,I349984);
nand I_16905 (I289271,I289254,I289062);
DFFARX1 I_16906 (I289271,I1862,I288878,I288858,);
nor I_16907 (I289302,I289130,I349984);
nor I_16908 (I289319,I289147,I289302);
nand I_16909 (I288867,I289319,I288997);
nor I_16910 (I289350,I289130,I288946);
nand I_16911 (I288861,I289350,I289237);
not I_16912 (I289405,I1869);
or I_16913 (I289422,I103042,I103054);
nand I_16914 (I289439,I103048,I103048);
not I_16915 (I289456,I289439);
nand I_16916 (I289473,I289456,I289422);
not I_16917 (I289490,I289473);
nand I_16918 (I289507,I103057,I103039);
nor I_16919 (I289524,I289507,I103045);
nor I_16920 (I289541,I289473,I289524);
or I_16921 (I289558,I289524,I289490);
nand I_16922 (I289382,I289473,I289524);
nand I_16923 (I289589,I289524,I289490);
and I_16924 (I289606,I289439,I289507);
nor I_16925 (I289623,I289541,I289606);
nor I_16926 (I289640,I103042,I103045);
not I_16927 (I289657,I103051);
nor I_16928 (I289674,I289657,I289640);
nor I_16929 (I289376,I289674,I289439);
nand I_16930 (I289705,I289674,I289558);
nor I_16931 (I289397,I289439,I289705);
nor I_16932 (I289379,I289674,I289623);
not I_16933 (I289391,I289674);
nor I_16934 (I289764,I289674,I103039);
or I_16935 (I289781,I289657,I103039);
nand I_16936 (I289798,I289781,I289589);
DFFARX1 I_16937 (I289798,I1862,I289405,I289385,);
nor I_16938 (I289829,I289657,I103039);
nor I_16939 (I289846,I289674,I289829);
nand I_16940 (I289394,I289846,I289524);
nor I_16941 (I289877,I289657,I289473);
nand I_16942 (I289388,I289877,I289764);
not I_16943 (I289932,I1869);
or I_16944 (I289949,I389336,I389339);
nand I_16945 (I289966,I389345,I389342);
not I_16946 (I289983,I289966);
nand I_16947 (I290000,I289983,I289949);
not I_16948 (I290017,I290000);
nand I_16949 (I290034,I389345,I389351);
nor I_16950 (I290051,I290034,I389336);
nor I_16951 (I290068,I290000,I290051);
or I_16952 (I290085,I290051,I290017);
nand I_16953 (I289909,I290000,I290051);
nand I_16954 (I290116,I290051,I290017);
and I_16955 (I290133,I289966,I290034);
nor I_16956 (I290150,I290068,I290133);
nor I_16957 (I290167,I389339,I389342);
not I_16958 (I290184,I389348);
nor I_16959 (I290201,I290184,I290167);
nor I_16960 (I289903,I290201,I289966);
nand I_16961 (I290232,I290201,I290085);
nor I_16962 (I289924,I289966,I290232);
nor I_16963 (I289906,I290201,I290150);
not I_16964 (I289918,I290201);
nor I_16965 (I290291,I290201,I389354);
or I_16966 (I290308,I290184,I389354);
nand I_16967 (I290325,I290308,I290116);
DFFARX1 I_16968 (I290325,I1862,I289932,I289912,);
nor I_16969 (I290356,I290184,I389354);
nor I_16970 (I290373,I290201,I290356);
nand I_16971 (I289921,I290373,I290051);
nor I_16972 (I290404,I290184,I290000);
nand I_16973 (I289915,I290404,I290291);
not I_16974 (I290459,I1869);
or I_16975 (I290476,I135767,I135785);
nand I_16976 (I290493,I135782,I135776);
not I_16977 (I290510,I290493);
nand I_16978 (I290527,I290510,I290476);
not I_16979 (I290544,I290527);
nand I_16980 (I290561,I135773,I135764);
nor I_16981 (I290578,I290561,I135788);
nor I_16982 (I290595,I290527,I290578);
or I_16983 (I290612,I290578,I290544);
nand I_16984 (I290436,I290527,I290578);
nand I_16985 (I290643,I290578,I290544);
and I_16986 (I290660,I290493,I290561);
nor I_16987 (I290677,I290595,I290660);
nor I_16988 (I290694,I135770,I135764);
not I_16989 (I290711,I135779);
nor I_16990 (I290728,I290711,I290694);
nor I_16991 (I290430,I290728,I290493);
nand I_16992 (I290759,I290728,I290612);
nor I_16993 (I290451,I290493,I290759);
nor I_16994 (I290433,I290728,I290677);
not I_16995 (I290445,I290728);
nor I_16996 (I290818,I290728,I135767);
or I_16997 (I290835,I290711,I135767);
nand I_16998 (I290852,I290835,I290643);
DFFARX1 I_16999 (I290852,I1862,I290459,I290439,);
nor I_17000 (I290883,I290711,I135767);
nor I_17001 (I290900,I290728,I290883);
nand I_17002 (I290448,I290900,I290578);
nor I_17003 (I290931,I290711,I290527);
nand I_17004 (I290442,I290931,I290818);
not I_17005 (I290986,I1869);
or I_17006 (I291003,I155266,I155284);
nand I_17007 (I291020,I155281,I155275);
not I_17008 (I291037,I291020);
nand I_17009 (I291054,I291037,I291003);
not I_17010 (I291071,I291054);
nand I_17011 (I291088,I155272,I155263);
nor I_17012 (I291105,I291088,I155287);
nor I_17013 (I291122,I291054,I291105);
or I_17014 (I291139,I291105,I291071);
nand I_17015 (I290963,I291054,I291105);
nand I_17016 (I291170,I291105,I291071);
and I_17017 (I291187,I291020,I291088);
nor I_17018 (I291204,I291122,I291187);
nor I_17019 (I291221,I155269,I155263);
not I_17020 (I291238,I155278);
nor I_17021 (I291255,I291238,I291221);
nor I_17022 (I290957,I291255,I291020);
nand I_17023 (I291286,I291255,I291139);
nor I_17024 (I290978,I291020,I291286);
nor I_17025 (I290960,I291255,I291204);
not I_17026 (I290972,I291255);
nor I_17027 (I291345,I291255,I155266);
or I_17028 (I291362,I291238,I155266);
nand I_17029 (I291379,I291362,I291170);
DFFARX1 I_17030 (I291379,I1862,I290986,I290966,);
nor I_17031 (I291410,I291238,I155266);
nor I_17032 (I291427,I291255,I291410);
nand I_17033 (I290975,I291427,I291105);
nor I_17034 (I291458,I291238,I291054);
nand I_17035 (I290969,I291458,I291345);
not I_17036 (I291513,I1869);
or I_17037 (I291530,I211078,I211060);
nand I_17038 (I291547,I211072,I211063);
not I_17039 (I291564,I291547);
nand I_17040 (I291581,I291564,I291530);
not I_17041 (I291598,I291581);
nand I_17042 (I291615,I211069,I211060);
nor I_17043 (I291632,I291615,I211057);
nor I_17044 (I291649,I291581,I291632);
or I_17045 (I291666,I291632,I291598);
nand I_17046 (I291490,I291581,I291632);
nand I_17047 (I291697,I291632,I291598);
and I_17048 (I291714,I291547,I291615);
nor I_17049 (I291731,I291649,I291714);
nor I_17050 (I291748,I211075,I211066);
not I_17051 (I291765,I211057);
nor I_17052 (I291782,I291765,I291748);
nor I_17053 (I291484,I291782,I291547);
nand I_17054 (I291813,I291782,I291666);
nor I_17055 (I291505,I291547,I291813);
nor I_17056 (I291487,I291782,I291731);
not I_17057 (I291499,I291782);
nor I_17058 (I291872,I291782,I211063);
or I_17059 (I291889,I291765,I211063);
nand I_17060 (I291906,I291889,I291697);
DFFARX1 I_17061 (I291906,I1862,I291513,I291493,);
nor I_17062 (I291937,I291765,I211063);
nor I_17063 (I291954,I291782,I291937);
nand I_17064 (I291502,I291954,I291632);
nor I_17065 (I291985,I291765,I291581);
nand I_17066 (I291496,I291985,I291872);
not I_17067 (I292040,I1869);
or I_17068 (I292057,I138402,I138420);
nand I_17069 (I292074,I138417,I138411);
not I_17070 (I292091,I292074);
nand I_17071 (I292108,I292091,I292057);
not I_17072 (I292125,I292108);
nand I_17073 (I292142,I138408,I138399);
nor I_17074 (I292159,I292142,I138423);
nor I_17075 (I292176,I292108,I292159);
or I_17076 (I292193,I292159,I292125);
nand I_17077 (I292017,I292108,I292159);
nand I_17078 (I292224,I292159,I292125);
and I_17079 (I292241,I292074,I292142);
nor I_17080 (I292258,I292176,I292241);
nor I_17081 (I292275,I138405,I138399);
not I_17082 (I292292,I138414);
nor I_17083 (I292309,I292292,I292275);
nor I_17084 (I292011,I292309,I292074);
nand I_17085 (I292340,I292309,I292193);
nor I_17086 (I292032,I292074,I292340);
nor I_17087 (I292014,I292309,I292258);
not I_17088 (I292026,I292309);
nor I_17089 (I292399,I292309,I138402);
or I_17090 (I292416,I292292,I138402);
nand I_17091 (I292433,I292416,I292224);
DFFARX1 I_17092 (I292433,I1862,I292040,I292020,);
nor I_17093 (I292464,I292292,I138402);
nor I_17094 (I292481,I292309,I292464);
nand I_17095 (I292029,I292481,I292159);
nor I_17096 (I292512,I292292,I292108);
nand I_17097 (I292023,I292512,I292399);
not I_17098 (I292567,I1869);
or I_17099 (I292584,I49693,I49714);
nand I_17100 (I292601,I49708,I49696);
not I_17101 (I292618,I292601);
nand I_17102 (I292635,I292618,I292584);
not I_17103 (I292652,I292635);
nand I_17104 (I292669,I49699,I49705);
nor I_17105 (I292686,I292669,I49711);
nor I_17106 (I292703,I292635,I292686);
or I_17107 (I292720,I292686,I292652);
nand I_17108 (I292544,I292635,I292686);
nand I_17109 (I292751,I292686,I292652);
and I_17110 (I292768,I292601,I292669);
nor I_17111 (I292785,I292703,I292768);
nor I_17112 (I292802,I49696,I49702);
not I_17113 (I292819,I49717);
nor I_17114 (I292836,I292819,I292802);
nor I_17115 (I292538,I292836,I292601);
nand I_17116 (I292867,I292836,I292720);
nor I_17117 (I292559,I292601,I292867);
nor I_17118 (I292541,I292836,I292785);
not I_17119 (I292553,I292836);
nor I_17120 (I292926,I292836,I49693);
or I_17121 (I292943,I292819,I49693);
nand I_17122 (I292960,I292943,I292751);
DFFARX1 I_17123 (I292960,I1862,I292567,I292547,);
nor I_17124 (I292991,I292819,I49693);
nor I_17125 (I293008,I292836,I292991);
nand I_17126 (I292556,I293008,I292686);
nor I_17127 (I293039,I292819,I292635);
nand I_17128 (I292550,I293039,I292926);
not I_17129 (I293094,I1869);
or I_17130 (I293111,I1535,I711);
nand I_17131 (I293128,I631,I1671);
not I_17132 (I293145,I293128);
nand I_17133 (I293162,I293145,I293111);
not I_17134 (I293179,I293162);
nand I_17135 (I293196,I1111,I655);
nor I_17136 (I293213,I293196,I1583);
nor I_17137 (I293230,I293162,I293213);
or I_17138 (I293247,I293213,I293179);
nand I_17139 (I293071,I293162,I293213);
nand I_17140 (I293278,I293213,I293179);
and I_17141 (I293295,I293128,I293196);
nor I_17142 (I293312,I293230,I293295);
nor I_17143 (I293329,I1439,I687);
not I_17144 (I293346,I1391);
nor I_17145 (I293363,I293346,I293329);
nor I_17146 (I293065,I293363,I293128);
nand I_17147 (I293394,I293363,I293247);
nor I_17148 (I293086,I293128,I293394);
nor I_17149 (I293068,I293363,I293312);
not I_17150 (I293080,I293363);
nor I_17151 (I293453,I293363,I1079);
or I_17152 (I293470,I293346,I1079);
nand I_17153 (I293487,I293470,I293278);
DFFARX1 I_17154 (I293487,I1862,I293094,I293074,);
nor I_17155 (I293518,I293346,I1079);
nor I_17156 (I293535,I293363,I293518);
nand I_17157 (I293083,I293535,I293213);
nor I_17158 (I293566,I293346,I293162);
nand I_17159 (I293077,I293566,I293453);
not I_17160 (I293621,I1869);
or I_17161 (I293638,I207746,I207728);
nand I_17162 (I293655,I207740,I207731);
not I_17163 (I293672,I293655);
nand I_17164 (I293689,I293672,I293638);
not I_17165 (I293706,I293689);
nand I_17166 (I293723,I207737,I207728);
nor I_17167 (I293740,I293723,I207725);
nor I_17168 (I293757,I293689,I293740);
or I_17169 (I293774,I293740,I293706);
nand I_17170 (I293598,I293689,I293740);
nand I_17171 (I293805,I293740,I293706);
and I_17172 (I293822,I293655,I293723);
nor I_17173 (I293839,I293757,I293822);
nor I_17174 (I293856,I207743,I207734);
not I_17175 (I293873,I207725);
nor I_17176 (I293890,I293873,I293856);
nor I_17177 (I293592,I293890,I293655);
nand I_17178 (I293921,I293890,I293774);
nor I_17179 (I293613,I293655,I293921);
nor I_17180 (I293595,I293890,I293839);
not I_17181 (I293607,I293890);
nor I_17182 (I293980,I293890,I207731);
or I_17183 (I293997,I293873,I207731);
nand I_17184 (I294014,I293997,I293805);
DFFARX1 I_17185 (I294014,I1862,I293621,I293601,);
nor I_17186 (I294045,I293873,I207731);
nor I_17187 (I294062,I293890,I294045);
nand I_17188 (I293610,I294062,I293740);
nor I_17189 (I294093,I293873,I293689);
nand I_17190 (I293604,I294093,I293980);
not I_17191 (I294148,I1869);
or I_17192 (I294165,I278670,I278652);
nand I_17193 (I294182,I278664,I278655);
not I_17194 (I294199,I294182);
nand I_17195 (I294216,I294199,I294165);
not I_17196 (I294233,I294216);
nand I_17197 (I294250,I278661,I278652);
nor I_17198 (I294267,I294250,I278649);
nor I_17199 (I294284,I294216,I294267);
or I_17200 (I294301,I294267,I294233);
nand I_17201 (I294125,I294216,I294267);
nand I_17202 (I294332,I294267,I294233);
and I_17203 (I294349,I294182,I294250);
nor I_17204 (I294366,I294284,I294349);
nor I_17205 (I294383,I278667,I278658);
not I_17206 (I294400,I278649);
nor I_17207 (I294417,I294400,I294383);
nor I_17208 (I294119,I294417,I294182);
nand I_17209 (I294448,I294417,I294301);
nor I_17210 (I294140,I294182,I294448);
nor I_17211 (I294122,I294417,I294366);
not I_17212 (I294134,I294417);
nor I_17213 (I294507,I294417,I278655);
or I_17214 (I294524,I294400,I278655);
nand I_17215 (I294541,I294524,I294332);
DFFARX1 I_17216 (I294541,I1862,I294148,I294128,);
nor I_17217 (I294572,I294400,I278655);
nor I_17218 (I294589,I294417,I294572);
nand I_17219 (I294137,I294589,I294267);
nor I_17220 (I294620,I294400,I294216);
nand I_17221 (I294131,I294620,I294507);
not I_17222 (I294675,I1869);
or I_17223 (I294692,I267246,I267228);
nand I_17224 (I294709,I267240,I267231);
not I_17225 (I294726,I294709);
nand I_17226 (I294743,I294726,I294692);
not I_17227 (I294760,I294743);
nand I_17228 (I294777,I267237,I267228);
nor I_17229 (I294794,I294777,I267225);
nor I_17230 (I294811,I294743,I294794);
or I_17231 (I294828,I294794,I294760);
nand I_17232 (I294652,I294743,I294794);
nand I_17233 (I294859,I294794,I294760);
and I_17234 (I294876,I294709,I294777);
nor I_17235 (I294893,I294811,I294876);
nor I_17236 (I294910,I267243,I267234);
not I_17237 (I294927,I267225);
nor I_17238 (I294944,I294927,I294910);
nor I_17239 (I294646,I294944,I294709);
nand I_17240 (I294975,I294944,I294828);
nor I_17241 (I294667,I294709,I294975);
nor I_17242 (I294649,I294944,I294893);
not I_17243 (I294661,I294944);
nor I_17244 (I295034,I294944,I267231);
or I_17245 (I295051,I294927,I267231);
nand I_17246 (I295068,I295051,I294859);
DFFARX1 I_17247 (I295068,I1862,I294675,I294655,);
nor I_17248 (I295099,I294927,I267231);
nor I_17249 (I295116,I294944,I295099);
nand I_17250 (I294664,I295116,I294794);
nor I_17251 (I295147,I294927,I294743);
nand I_17252 (I294658,I295147,I295034);
not I_17253 (I295202,I1869);
or I_17254 (I295219,I118903,I118921);
nand I_17255 (I295236,I118918,I118912);
not I_17256 (I295253,I295236);
nand I_17257 (I295270,I295253,I295219);
not I_17258 (I295287,I295270);
nand I_17259 (I295304,I118909,I118900);
nor I_17260 (I295321,I295304,I118924);
nor I_17261 (I295338,I295270,I295321);
or I_17262 (I295355,I295321,I295287);
nand I_17263 (I295179,I295270,I295321);
nand I_17264 (I295386,I295321,I295287);
and I_17265 (I295403,I295236,I295304);
nor I_17266 (I295420,I295338,I295403);
nor I_17267 (I295437,I118906,I118900);
not I_17268 (I295454,I118915);
nor I_17269 (I295471,I295454,I295437);
nor I_17270 (I295173,I295471,I295236);
nand I_17271 (I295502,I295471,I295355);
nor I_17272 (I295194,I295236,I295502);
nor I_17273 (I295176,I295471,I295420);
not I_17274 (I295188,I295471);
nor I_17275 (I295561,I295471,I118903);
or I_17276 (I295578,I295454,I118903);
nand I_17277 (I295595,I295578,I295386);
DFFARX1 I_17278 (I295595,I1862,I295202,I295182,);
nor I_17279 (I295626,I295454,I118903);
nor I_17280 (I295643,I295471,I295626);
nand I_17281 (I295191,I295643,I295321);
nor I_17282 (I295674,I295454,I295270);
nand I_17283 (I295185,I295674,I295561);
not I_17284 (I295729,I1869);
or I_17285 (I295746,I222502,I222484);
nand I_17286 (I295763,I222496,I222487);
not I_17287 (I295780,I295763);
nand I_17288 (I295797,I295780,I295746);
not I_17289 (I295814,I295797);
nand I_17290 (I295831,I222493,I222484);
nor I_17291 (I295848,I295831,I222481);
nor I_17292 (I295865,I295797,I295848);
or I_17293 (I295882,I295848,I295814);
nand I_17294 (I295706,I295797,I295848);
nand I_17295 (I295913,I295848,I295814);
and I_17296 (I295930,I295763,I295831);
nor I_17297 (I295947,I295865,I295930);
nor I_17298 (I295964,I222499,I222490);
not I_17299 (I295981,I222481);
nor I_17300 (I295998,I295981,I295964);
nor I_17301 (I295700,I295998,I295763);
nand I_17302 (I296029,I295998,I295882);
nor I_17303 (I295721,I295763,I296029);
nor I_17304 (I295703,I295998,I295947);
not I_17305 (I295715,I295998);
nor I_17306 (I296088,I295998,I222487);
or I_17307 (I296105,I295981,I222487);
nand I_17308 (I296122,I296105,I295913);
DFFARX1 I_17309 (I296122,I1862,I295729,I295709,);
nor I_17310 (I296153,I295981,I222487);
nor I_17311 (I296170,I295998,I296153);
nand I_17312 (I295718,I296170,I295848);
nor I_17313 (I296201,I295981,I295797);
nand I_17314 (I295712,I296201,I296088);
not I_17315 (I296256,I1869);
or I_17316 (I296273,I365910,I365913);
nand I_17317 (I296290,I365919,I365916);
not I_17318 (I296307,I296290);
nand I_17319 (I296324,I296307,I296273);
not I_17320 (I296341,I296324);
nand I_17321 (I296358,I365919,I365925);
nor I_17322 (I296375,I296358,I365910);
nor I_17323 (I296392,I296324,I296375);
or I_17324 (I296409,I296375,I296341);
nand I_17325 (I296233,I296324,I296375);
nand I_17326 (I296440,I296375,I296341);
and I_17327 (I296457,I296290,I296358);
nor I_17328 (I296474,I296392,I296457);
nor I_17329 (I296491,I365913,I365916);
not I_17330 (I296508,I365922);
nor I_17331 (I296525,I296508,I296491);
nor I_17332 (I296227,I296525,I296290);
nand I_17333 (I296556,I296525,I296409);
nor I_17334 (I296248,I296290,I296556);
nor I_17335 (I296230,I296525,I296474);
not I_17336 (I296242,I296525);
nor I_17337 (I296615,I296525,I365928);
or I_17338 (I296632,I296508,I365928);
nand I_17339 (I296649,I296632,I296440);
DFFARX1 I_17340 (I296649,I1862,I296256,I296236,);
nor I_17341 (I296680,I296508,I365928);
nor I_17342 (I296697,I296525,I296680);
nand I_17343 (I296245,I296697,I296375);
nor I_17344 (I296728,I296508,I296324);
nand I_17345 (I296239,I296728,I296615);
not I_17346 (I296783,I1869);
or I_17347 (I296800,I409668,I409671);
nand I_17348 (I296817,I409677,I409674);
not I_17349 (I296834,I296817);
nand I_17350 (I296851,I296834,I296800);
not I_17351 (I296868,I296851);
nand I_17352 (I296885,I409677,I409683);
nor I_17353 (I296902,I296885,I409668);
nor I_17354 (I296919,I296851,I296902);
or I_17355 (I296936,I296902,I296868);
nand I_17356 (I296760,I296851,I296902);
nand I_17357 (I296967,I296902,I296868);
and I_17358 (I296984,I296817,I296885);
nor I_17359 (I297001,I296919,I296984);
nor I_17360 (I297018,I409671,I409674);
not I_17361 (I297035,I409680);
nor I_17362 (I297052,I297035,I297018);
nor I_17363 (I296754,I297052,I296817);
nand I_17364 (I297083,I297052,I296936);
nor I_17365 (I296775,I296817,I297083);
nor I_17366 (I296757,I297052,I297001);
not I_17367 (I296769,I297052);
nor I_17368 (I297142,I297052,I409686);
or I_17369 (I297159,I297035,I409686);
nand I_17370 (I297176,I297159,I296967);
DFFARX1 I_17371 (I297176,I1862,I296783,I296763,);
nor I_17372 (I297207,I297035,I409686);
nor I_17373 (I297224,I297052,I297207);
nand I_17374 (I296772,I297224,I296902);
nor I_17375 (I297255,I297035,I296851);
nand I_17376 (I296766,I297255,I297142);
not I_17377 (I297310,I1869);
or I_17378 (I297327,I153158,I153176);
nand I_17379 (I297344,I153173,I153167);
not I_17380 (I297361,I297344);
nand I_17381 (I297378,I297361,I297327);
not I_17382 (I297395,I297378);
nand I_17383 (I297412,I153164,I153155);
nor I_17384 (I297429,I297412,I153179);
nor I_17385 (I297446,I297378,I297429);
or I_17386 (I297463,I297429,I297395);
nand I_17387 (I297287,I297378,I297429);
nand I_17388 (I297494,I297429,I297395);
and I_17389 (I297511,I297344,I297412);
nor I_17390 (I297528,I297446,I297511);
nor I_17391 (I297545,I153161,I153155);
not I_17392 (I297562,I153170);
nor I_17393 (I297579,I297562,I297545);
nor I_17394 (I297281,I297579,I297344);
nand I_17395 (I297610,I297579,I297463);
nor I_17396 (I297302,I297344,I297610);
nor I_17397 (I297284,I297579,I297528);
not I_17398 (I297296,I297579);
nor I_17399 (I297669,I297579,I153158);
or I_17400 (I297686,I297562,I153158);
nand I_17401 (I297703,I297686,I297494);
DFFARX1 I_17402 (I297703,I1862,I297310,I297290,);
nor I_17403 (I297734,I297562,I153158);
nor I_17404 (I297751,I297579,I297734);
nand I_17405 (I297299,I297751,I297429);
nor I_17406 (I297782,I297562,I297378);
nand I_17407 (I297293,I297782,I297669);
not I_17408 (I297837,I1869);
or I_17409 (I297854,I59383,I59404);
nand I_17410 (I297871,I59398,I59386);
not I_17411 (I297888,I297871);
nand I_17412 (I297905,I297888,I297854);
not I_17413 (I297922,I297905);
nand I_17414 (I297939,I59389,I59395);
nor I_17415 (I297956,I297939,I59401);
nor I_17416 (I297973,I297905,I297956);
or I_17417 (I297990,I297956,I297922);
nand I_17418 (I297814,I297905,I297956);
nand I_17419 (I298021,I297956,I297922);
and I_17420 (I298038,I297871,I297939);
nor I_17421 (I298055,I297973,I298038);
nor I_17422 (I298072,I59386,I59392);
not I_17423 (I298089,I59407);
nor I_17424 (I298106,I298089,I298072);
nor I_17425 (I297808,I298106,I297871);
nand I_17426 (I298137,I298106,I297990);
nor I_17427 (I297829,I297871,I298137);
nor I_17428 (I297811,I298106,I298055);
not I_17429 (I297823,I298106);
nor I_17430 (I298196,I298106,I59383);
or I_17431 (I298213,I298089,I59383);
nand I_17432 (I298230,I298213,I298021);
DFFARX1 I_17433 (I298230,I1862,I297837,I297817,);
nor I_17434 (I298261,I298089,I59383);
nor I_17435 (I298278,I298106,I298261);
nand I_17436 (I297826,I298278,I297956);
nor I_17437 (I298309,I298089,I297905);
nand I_17438 (I297820,I298309,I298196);
not I_17439 (I298364,I1869);
or I_17440 (I298381,I340495,I340507);
nand I_17441 (I298398,I340510,I340513);
not I_17442 (I298415,I298398);
nand I_17443 (I298432,I298415,I298381);
not I_17444 (I298449,I298432);
nand I_17445 (I298466,I340495,I340498);
nor I_17446 (I298483,I298466,I340501);
nor I_17447 (I298500,I298432,I298483);
or I_17448 (I298517,I298483,I298449);
nand I_17449 (I298341,I298432,I298483);
nand I_17450 (I298548,I298483,I298449);
and I_17451 (I298565,I298398,I298466);
nor I_17452 (I298582,I298500,I298565);
nor I_17453 (I298599,I340504,I340501);
not I_17454 (I298616,I340516);
nor I_17455 (I298633,I298616,I298599);
nor I_17456 (I298335,I298633,I298398);
nand I_17457 (I298664,I298633,I298517);
nor I_17458 (I298356,I298398,I298664);
nor I_17459 (I298338,I298633,I298582);
not I_17460 (I298350,I298633);
nor I_17461 (I298723,I298633,I340498);
or I_17462 (I298740,I298616,I340498);
nand I_17463 (I298757,I298740,I298548);
DFFARX1 I_17464 (I298757,I1862,I298364,I298344,);
nor I_17465 (I298788,I298616,I340498);
nor I_17466 (I298805,I298633,I298788);
nand I_17467 (I298353,I298805,I298483);
nor I_17468 (I298836,I298616,I298432);
nand I_17469 (I298347,I298836,I298723);
not I_17470 (I298891,I1869);
or I_17471 (I298908,I16033,I16054);
nand I_17472 (I298925,I16048,I16036);
not I_17473 (I298942,I298925);
nand I_17474 (I298959,I298942,I298908);
not I_17475 (I298976,I298959);
nand I_17476 (I298993,I16039,I16045);
nor I_17477 (I299010,I298993,I16051);
nor I_17478 (I299027,I298959,I299010);
or I_17479 (I299044,I299010,I298976);
nand I_17480 (I298868,I298959,I299010);
nand I_17481 (I299075,I299010,I298976);
and I_17482 (I299092,I298925,I298993);
nor I_17483 (I299109,I299027,I299092);
nor I_17484 (I299126,I16036,I16042);
not I_17485 (I299143,I16057);
nor I_17486 (I299160,I299143,I299126);
nor I_17487 (I298862,I299160,I298925);
nand I_17488 (I299191,I299160,I299044);
nor I_17489 (I298883,I298925,I299191);
nor I_17490 (I298865,I299160,I299109);
not I_17491 (I298877,I299160);
nor I_17492 (I299250,I299160,I16033);
or I_17493 (I299267,I299143,I16033);
nand I_17494 (I299284,I299267,I299075);
DFFARX1 I_17495 (I299284,I1862,I298891,I298871,);
nor I_17496 (I299315,I299143,I16033);
nor I_17497 (I299332,I299160,I299315);
nand I_17498 (I298880,I299332,I299010);
nor I_17499 (I299363,I299143,I298959);
nand I_17500 (I298874,I299363,I299250);
not I_17501 (I299418,I1869);
or I_17502 (I299435,I375634,I375637);
nand I_17503 (I299452,I375643,I375640);
not I_17504 (I299469,I299452);
nand I_17505 (I299486,I299469,I299435);
not I_17506 (I299503,I299486);
nand I_17507 (I299520,I375643,I375649);
nor I_17508 (I299537,I299520,I375634);
nor I_17509 (I299554,I299486,I299537);
or I_17510 (I299571,I299537,I299503);
nand I_17511 (I299395,I299486,I299537);
nand I_17512 (I299602,I299537,I299503);
and I_17513 (I299619,I299452,I299520);
nor I_17514 (I299636,I299554,I299619);
nor I_17515 (I299653,I375637,I375640);
not I_17516 (I299670,I375646);
nor I_17517 (I299687,I299670,I299653);
nor I_17518 (I299389,I299687,I299452);
nand I_17519 (I299718,I299687,I299571);
nor I_17520 (I299410,I299452,I299718);
nor I_17521 (I299392,I299687,I299636);
not I_17522 (I299404,I299687);
nor I_17523 (I299777,I299687,I375652);
or I_17524 (I299794,I299670,I375652);
nand I_17525 (I299811,I299794,I299602);
DFFARX1 I_17526 (I299811,I1862,I299418,I299398,);
nor I_17527 (I299842,I299670,I375652);
nor I_17528 (I299859,I299687,I299842);
nand I_17529 (I299407,I299859,I299537);
nor I_17530 (I299890,I299670,I299486);
nand I_17531 (I299401,I299890,I299777);
not I_17532 (I299945,I1869);
or I_17533 (I299962,I94573,I94594);
nand I_17534 (I299979,I94588,I94576);
not I_17535 (I299996,I299979);
nand I_17536 (I300013,I299996,I299962);
not I_17537 (I300030,I300013);
nand I_17538 (I300047,I94579,I94585);
nor I_17539 (I300064,I300047,I94591);
nor I_17540 (I300081,I300013,I300064);
or I_17541 (I300098,I300064,I300030);
nand I_17542 (I299922,I300013,I300064);
nand I_17543 (I300129,I300064,I300030);
and I_17544 (I300146,I299979,I300047);
nor I_17545 (I300163,I300081,I300146);
nor I_17546 (I300180,I94576,I94582);
not I_17547 (I300197,I94597);
nor I_17548 (I300214,I300197,I300180);
nor I_17549 (I299916,I300214,I299979);
nand I_17550 (I300245,I300214,I300098);
nor I_17551 (I299937,I299979,I300245);
nor I_17552 (I299919,I300214,I300163);
not I_17553 (I299931,I300214);
nor I_17554 (I300304,I300214,I94573);
or I_17555 (I300321,I300197,I94573);
nand I_17556 (I300338,I300321,I300129);
DFFARX1 I_17557 (I300338,I1862,I299945,I299925,);
nor I_17558 (I300369,I300197,I94573);
nor I_17559 (I300386,I300214,I300369);
nand I_17560 (I299934,I300386,I300064);
nor I_17561 (I300417,I300197,I300013);
nand I_17562 (I299928,I300417,I300304);
not I_17563 (I300472,I1869);
or I_17564 (I300489,I11888,I11903);
nand I_17565 (I300506,I11891,I11891);
not I_17566 (I300523,I300506);
nand I_17567 (I300540,I300523,I300489);
not I_17568 (I300557,I300540);
nand I_17569 (I300574,I11894,I11897);
nor I_17570 (I300591,I300574,I11906);
nor I_17571 (I300608,I300540,I300591);
or I_17572 (I300625,I300591,I300557);
nand I_17573 (I300449,I300540,I300591);
nand I_17574 (I300656,I300591,I300557);
and I_17575 (I300673,I300506,I300574);
nor I_17576 (I300690,I300608,I300673);
nor I_17577 (I300707,I11888,I11885);
not I_17578 (I300724,I11900);
nor I_17579 (I300741,I300724,I300707);
nor I_17580 (I300443,I300741,I300506);
nand I_17581 (I300772,I300741,I300625);
nor I_17582 (I300464,I300506,I300772);
nor I_17583 (I300446,I300741,I300690);
not I_17584 (I300458,I300741);
nor I_17585 (I300831,I300741,I11885);
or I_17586 (I300848,I300724,I11885);
nand I_17587 (I300865,I300848,I300656);
DFFARX1 I_17588 (I300865,I1862,I300472,I300452,);
nor I_17589 (I300896,I300724,I11885);
nor I_17590 (I300913,I300741,I300896);
nand I_17591 (I300461,I300913,I300591);
nor I_17592 (I300944,I300724,I300540);
nand I_17593 (I300455,I300944,I300831);
not I_17594 (I300999,I1869);
or I_17595 (I301016,I392872,I392875);
nand I_17596 (I301033,I392881,I392878);
not I_17597 (I301050,I301033);
nand I_17598 (I301067,I301050,I301016);
not I_17599 (I301084,I301067);
nand I_17600 (I301101,I392881,I392887);
nor I_17601 (I301118,I301101,I392872);
nor I_17602 (I301135,I301067,I301118);
or I_17603 (I301152,I301118,I301084);
nand I_17604 (I300976,I301067,I301118);
nand I_17605 (I301183,I301118,I301084);
and I_17606 (I301200,I301033,I301101);
nor I_17607 (I301217,I301135,I301200);
nor I_17608 (I301234,I392875,I392878);
not I_17609 (I301251,I392884);
nor I_17610 (I301268,I301251,I301234);
nor I_17611 (I300970,I301268,I301033);
nand I_17612 (I301299,I301268,I301152);
nor I_17613 (I300991,I301033,I301299);
nor I_17614 (I300973,I301268,I301217);
not I_17615 (I300985,I301268);
nor I_17616 (I301358,I301268,I392890);
or I_17617 (I301375,I301251,I392890);
nand I_17618 (I301392,I301375,I301183);
DFFARX1 I_17619 (I301392,I1862,I300999,I300979,);
nor I_17620 (I301423,I301251,I392890);
nor I_17621 (I301440,I301268,I301423);
nand I_17622 (I300988,I301440,I301118);
nor I_17623 (I301471,I301251,I301067);
nand I_17624 (I300982,I301471,I301358);
not I_17625 (I301526,I1869);
or I_17626 (I301543,I6091,I6106);
nand I_17627 (I301560,I6094,I6094);
not I_17628 (I301577,I301560);
nand I_17629 (I301594,I301577,I301543);
not I_17630 (I301611,I301594);
nand I_17631 (I301628,I6097,I6100);
nor I_17632 (I301645,I301628,I6109);
nor I_17633 (I301662,I301594,I301645);
or I_17634 (I301679,I301645,I301611);
nand I_17635 (I301503,I301594,I301645);
nand I_17636 (I301710,I301645,I301611);
and I_17637 (I301727,I301560,I301628);
nor I_17638 (I301744,I301662,I301727);
nor I_17639 (I301761,I6091,I6088);
not I_17640 (I301778,I6103);
nor I_17641 (I301795,I301778,I301761);
nor I_17642 (I301497,I301795,I301560);
nand I_17643 (I301826,I301795,I301679);
nor I_17644 (I301518,I301560,I301826);
nor I_17645 (I301500,I301795,I301744);
not I_17646 (I301512,I301795);
nor I_17647 (I301885,I301795,I6088);
or I_17648 (I301902,I301778,I6088);
nand I_17649 (I301919,I301902,I301710);
DFFARX1 I_17650 (I301919,I1862,I301526,I301506,);
nor I_17651 (I301950,I301778,I6088);
nor I_17652 (I301967,I301795,I301950);
nand I_17653 (I301515,I301967,I301645);
nor I_17654 (I301998,I301778,I301594);
nand I_17655 (I301509,I301998,I301885);
not I_17656 (I302053,I1869);
or I_17657 (I302070,I164225,I164243);
nand I_17658 (I302087,I164240,I164234);
not I_17659 (I302104,I302087);
nand I_17660 (I302121,I302104,I302070);
not I_17661 (I302138,I302121);
nand I_17662 (I302155,I164231,I164222);
nor I_17663 (I302172,I302155,I164246);
nor I_17664 (I302189,I302121,I302172);
or I_17665 (I302206,I302172,I302138);
nand I_17666 (I302030,I302121,I302172);
nand I_17667 (I302237,I302172,I302138);
and I_17668 (I302254,I302087,I302155);
nor I_17669 (I302271,I302189,I302254);
nor I_17670 (I302288,I164228,I164222);
not I_17671 (I302305,I164237);
nor I_17672 (I302322,I302305,I302288);
nor I_17673 (I302024,I302322,I302087);
nand I_17674 (I302353,I302322,I302206);
nor I_17675 (I302045,I302087,I302353);
nor I_17676 (I302027,I302322,I302271);
not I_17677 (I302039,I302322);
nor I_17678 (I302412,I302322,I164225);
or I_17679 (I302429,I302305,I164225);
nand I_17680 (I302446,I302429,I302237);
DFFARX1 I_17681 (I302446,I1862,I302053,I302033,);
nor I_17682 (I302477,I302305,I164225);
nor I_17683 (I302494,I302322,I302477);
nand I_17684 (I302042,I302494,I302172);
nor I_17685 (I302525,I302305,I302121);
nand I_17686 (I302036,I302525,I302412);
not I_17687 (I302580,I1869);
or I_17688 (I302597,I216790,I216772);
nand I_17689 (I302614,I216784,I216775);
not I_17690 (I302631,I302614);
nand I_17691 (I302648,I302631,I302597);
not I_17692 (I302665,I302648);
nand I_17693 (I302682,I216781,I216772);
nor I_17694 (I302699,I302682,I216769);
nor I_17695 (I302716,I302648,I302699);
or I_17696 (I302733,I302699,I302665);
nand I_17697 (I302557,I302648,I302699);
nand I_17698 (I302764,I302699,I302665);
and I_17699 (I302781,I302614,I302682);
nor I_17700 (I302798,I302716,I302781);
nor I_17701 (I302815,I216787,I216778);
not I_17702 (I302832,I216769);
nor I_17703 (I302849,I302832,I302815);
nor I_17704 (I302551,I302849,I302614);
nand I_17705 (I302880,I302849,I302733);
nor I_17706 (I302572,I302614,I302880);
nor I_17707 (I302554,I302849,I302798);
not I_17708 (I302566,I302849);
nor I_17709 (I302939,I302849,I216775);
or I_17710 (I302956,I302832,I216775);
nand I_17711 (I302973,I302956,I302764);
DFFARX1 I_17712 (I302973,I1862,I302580,I302560,);
nor I_17713 (I303004,I302832,I216775);
nor I_17714 (I303021,I302849,I303004);
nand I_17715 (I302569,I303021,I302699);
nor I_17716 (I303052,I302832,I302648);
nand I_17717 (I302563,I303052,I302939);
not I_17718 (I303107,I1869);
nor I_17719 (I303124,I239635,I239623);
not I_17720 (I303141,I239620);
not I_17721 (I303158,I239617);
nor I_17722 (I303175,I303158,I303124);
nand I_17723 (I303192,I303175,I239620);
not I_17724 (I303081,I303192);
nor I_17725 (I303223,I303158,I303141);
and I_17726 (I303240,I303192,I239620);
nor I_17727 (I303257,I303223,I239620);
nand I_17728 (I303274,I239623,I239629);
not I_17729 (I303291,I303274);
nand I_17730 (I303308,I303291,I303257);
nor I_17731 (I303325,I239638,I239632);
not I_17732 (I303342,I239626);
nor I_17733 (I303359,I303342,I239617);
nor I_17734 (I303078,I303359,I303192);
not I_17735 (I303390,I303359);
or I_17736 (I303093,I303308,I303359);
nor I_17737 (I303421,I303359,I303274);
nand I_17738 (I303090,I303223,I303421);
nor I_17739 (I303452,I303325,I303342);
nand I_17740 (I303469,I303291,I303452);
not I_17741 (I303096,I303469);
nor I_17742 (I303099,I303240,I303469);
or I_17743 (I303514,I303359,I303452);
nor I_17744 (I303084,I303291,I303514);
nor I_17745 (I303545,I303452,I239620);
nand I_17746 (I303562,I303545,I303291);
nand I_17747 (I303579,I303390,I303562);
DFFARX1 I_17748 (I303579,I1862,I303107,I303087,);
not I_17749 (I303634,I1869);
nor I_17750 (I303651,I226307,I226295);
not I_17751 (I303668,I226292);
not I_17752 (I303685,I226289);
nor I_17753 (I303702,I303685,I303651);
nand I_17754 (I303719,I303702,I226292);
not I_17755 (I303608,I303719);
nor I_17756 (I303750,I303685,I303668);
and I_17757 (I303767,I303719,I226292);
nor I_17758 (I303784,I303750,I226292);
nand I_17759 (I303801,I226295,I226301);
not I_17760 (I303818,I303801);
nand I_17761 (I303835,I303818,I303784);
nor I_17762 (I303852,I226310,I226304);
not I_17763 (I303869,I226298);
nor I_17764 (I303886,I303869,I226289);
nor I_17765 (I303605,I303886,I303719);
not I_17766 (I303917,I303886);
or I_17767 (I303620,I303835,I303886);
nor I_17768 (I303948,I303886,I303801);
nand I_17769 (I303617,I303750,I303948);
nor I_17770 (I303979,I303852,I303869);
nand I_17771 (I303996,I303818,I303979);
not I_17772 (I303623,I303996);
nor I_17773 (I303626,I303767,I303996);
or I_17774 (I304041,I303886,I303979);
nor I_17775 (I303611,I303818,I304041);
nor I_17776 (I304072,I303979,I226292);
nand I_17777 (I304089,I304072,I303818);
nand I_17778 (I304106,I303917,I304089);
DFFARX1 I_17779 (I304106,I1862,I303634,I303614,);
not I_17780 (I304161,I1869);
nor I_17781 (I304178,I235827,I235815);
not I_17782 (I304195,I235812);
not I_17783 (I304212,I235809);
nor I_17784 (I304229,I304212,I304178);
nand I_17785 (I304246,I304229,I235812);
not I_17786 (I304135,I304246);
nor I_17787 (I304277,I304212,I304195);
and I_17788 (I304294,I304246,I235812);
nor I_17789 (I304311,I304277,I235812);
nand I_17790 (I304328,I235815,I235821);
not I_17791 (I304345,I304328);
nand I_17792 (I304362,I304345,I304311);
nor I_17793 (I304379,I235830,I235824);
not I_17794 (I304396,I235818);
nor I_17795 (I304413,I304396,I235809);
nor I_17796 (I304132,I304413,I304246);
not I_17797 (I304444,I304413);
or I_17798 (I304147,I304362,I304413);
nor I_17799 (I304475,I304413,I304328);
nand I_17800 (I304144,I304277,I304475);
nor I_17801 (I304506,I304379,I304396);
nand I_17802 (I304523,I304345,I304506);
not I_17803 (I304150,I304523);
nor I_17804 (I304153,I304294,I304523);
or I_17805 (I304568,I304413,I304506);
nor I_17806 (I304138,I304345,I304568);
nor I_17807 (I304599,I304506,I235812);
nand I_17808 (I304616,I304599,I304345);
nand I_17809 (I304633,I304444,I304616);
DFFARX1 I_17810 (I304633,I1862,I304161,I304141,);
not I_17811 (I304688,I1869);
nor I_17812 (I304705,I397734,I397737);
not I_17813 (I304722,I397749);
not I_17814 (I304739,I397740);
nor I_17815 (I304756,I304739,I304705);
nand I_17816 (I304773,I304756,I397749);
not I_17817 (I304662,I304773);
nor I_17818 (I304804,I304739,I304722);
and I_17819 (I304821,I304773,I397743);
nor I_17820 (I304838,I304804,I397743);
nand I_17821 (I304855,I397740,I397746);
not I_17822 (I304872,I304855);
nand I_17823 (I304889,I304872,I304838);
nor I_17824 (I304906,I397737,I397752);
not I_17825 (I304923,I397743);
nor I_17826 (I304940,I304923,I397734);
nor I_17827 (I304659,I304940,I304773);
not I_17828 (I304971,I304940);
or I_17829 (I304674,I304889,I304940);
nor I_17830 (I305002,I304940,I304855);
nand I_17831 (I304671,I304804,I305002);
nor I_17832 (I305033,I304906,I304923);
nand I_17833 (I305050,I304872,I305033);
not I_17834 (I304677,I305050);
nor I_17835 (I304680,I304821,I305050);
or I_17836 (I305095,I304940,I305033);
nor I_17837 (I304665,I304872,I305095);
nor I_17838 (I305126,I305033,I397743);
nand I_17839 (I305143,I305126,I304872);
nand I_17840 (I305160,I304971,I305143);
DFFARX1 I_17841 (I305160,I1862,I304688,I304668,);
not I_17842 (I305215,I1869);
nor I_17843 (I305232,I91516,I91513);
not I_17844 (I305249,I91531);
not I_17845 (I305266,I91522);
nor I_17846 (I305283,I305266,I305232);
nand I_17847 (I305300,I305283,I91531);
not I_17848 (I305189,I305300);
nor I_17849 (I305331,I305266,I305249);
and I_17850 (I305348,I305300,I91537);
nor I_17851 (I305365,I305331,I91537);
nand I_17852 (I305382,I91534,I91525);
not I_17853 (I305399,I305382);
nand I_17854 (I305416,I305399,I305365);
nor I_17855 (I305433,I91513,I91516);
not I_17856 (I305450,I91528);
nor I_17857 (I305467,I305450,I91519);
nor I_17858 (I305186,I305467,I305300);
not I_17859 (I305498,I305467);
or I_17860 (I305201,I305416,I305467);
nor I_17861 (I305529,I305467,I305382);
nand I_17862 (I305198,I305331,I305529);
nor I_17863 (I305560,I305433,I305450);
nand I_17864 (I305577,I305399,I305560);
not I_17865 (I305204,I305577);
nor I_17866 (I305207,I305348,I305577);
or I_17867 (I305622,I305467,I305560);
nor I_17868 (I305192,I305399,I305622);
nor I_17869 (I305653,I305560,I91537);
nand I_17870 (I305670,I305653,I305399);
nand I_17871 (I305687,I305498,I305670);
DFFARX1 I_17872 (I305687,I1862,I305215,I305195,);
not I_17873 (I305742,I1869);
nor I_17874 (I305759,I11358,I11361);
not I_17875 (I305776,I11373);
not I_17876 (I305793,I11364);
nor I_17877 (I305810,I305793,I305759);
nand I_17878 (I305827,I305810,I11373);
not I_17879 (I305716,I305827);
nor I_17880 (I305858,I305793,I305776);
and I_17881 (I305875,I305827,I11361);
nor I_17882 (I305892,I305858,I11361);
nand I_17883 (I305909,I11367,I11364);
not I_17884 (I305926,I305909);
nand I_17885 (I305943,I305926,I305892);
nor I_17886 (I305960,I11379,I11376);
not I_17887 (I305977,I11370);
nor I_17888 (I305994,I305977,I11358);
nor I_17889 (I305713,I305994,I305827);
not I_17890 (I306025,I305994);
or I_17891 (I305728,I305943,I305994);
nor I_17892 (I306056,I305994,I305909);
nand I_17893 (I305725,I305858,I306056);
nor I_17894 (I306087,I305960,I305977);
nand I_17895 (I306104,I305926,I306087);
not I_17896 (I305731,I306104);
nor I_17897 (I305734,I305875,I306104);
or I_17898 (I306149,I305994,I306087);
nor I_17899 (I305719,I305926,I306149);
nor I_17900 (I306180,I306087,I11361);
nand I_17901 (I306197,I306180,I305926);
nand I_17902 (I306214,I306025,I306197);
DFFARX1 I_17903 (I306214,I1862,I305742,I305722,);
not I_17904 (I306269,I1869);
nor I_17905 (I306286,I362816,I362819);
not I_17906 (I306303,I362831);
not I_17907 (I306320,I362822);
nor I_17908 (I306337,I306320,I306286);
nand I_17909 (I306354,I306337,I362831);
not I_17910 (I306243,I306354);
nor I_17911 (I306385,I306320,I306303);
and I_17912 (I306402,I306354,I362825);
nor I_17913 (I306419,I306385,I362825);
nand I_17914 (I306436,I362822,I362828);
not I_17915 (I306453,I306436);
nand I_17916 (I306470,I306453,I306419);
nor I_17917 (I306487,I362819,I362834);
not I_17918 (I306504,I362825);
nor I_17919 (I306521,I306504,I362816);
nor I_17920 (I306240,I306521,I306354);
not I_17921 (I306552,I306521);
or I_17922 (I306255,I306470,I306521);
nor I_17923 (I306583,I306521,I306436);
nand I_17924 (I306252,I306385,I306583);
nor I_17925 (I306614,I306487,I306504);
nand I_17926 (I306631,I306453,I306614);
not I_17927 (I306258,I306631);
nor I_17928 (I306261,I306402,I306631);
or I_17929 (I306676,I306521,I306614);
nor I_17930 (I306246,I306453,I306676);
nor I_17931 (I306707,I306614,I362825);
nand I_17932 (I306724,I306707,I306453);
nand I_17933 (I306741,I306552,I306724);
DFFARX1 I_17934 (I306741,I1862,I306269,I306249,);
not I_17935 (I306796,I1869);
nor I_17936 (I306813,I281999,I281987);
not I_17937 (I306830,I281984);
not I_17938 (I306847,I281981);
nor I_17939 (I306864,I306847,I306813);
nand I_17940 (I306881,I306864,I281984);
not I_17941 (I306770,I306881);
nor I_17942 (I306912,I306847,I306830);
and I_17943 (I306929,I306881,I281984);
nor I_17944 (I306946,I306912,I281984);
nand I_17945 (I306963,I281987,I281993);
not I_17946 (I306980,I306963);
nand I_17947 (I306997,I306980,I306946);
nor I_17948 (I307014,I282002,I281996);
not I_17949 (I307031,I281990);
nor I_17950 (I307048,I307031,I281981);
nor I_17951 (I306767,I307048,I306881);
not I_17952 (I307079,I307048);
or I_17953 (I306782,I306997,I307048);
nor I_17954 (I307110,I307048,I306963);
nand I_17955 (I306779,I306912,I307110);
nor I_17956 (I307141,I307014,I307031);
nand I_17957 (I307158,I306980,I307141);
not I_17958 (I306785,I307158);
nor I_17959 (I306788,I306929,I307158);
or I_17960 (I307203,I307048,I307141);
nor I_17961 (I306773,I306980,I307203);
nor I_17962 (I307234,I307141,I281984);
nand I_17963 (I307251,I307234,I306980);
nand I_17964 (I307268,I307079,I307251);
DFFARX1 I_17965 (I307268,I1862,I306796,I306776,);
not I_17966 (I307323,I1869);
nor I_17967 (I307340,I46126,I46123);
not I_17968 (I307357,I46141);
not I_17969 (I307374,I46132);
nor I_17970 (I307391,I307374,I307340);
nand I_17971 (I307408,I307391,I46141);
not I_17972 (I307297,I307408);
nor I_17973 (I307439,I307374,I307357);
and I_17974 (I307456,I307408,I46147);
nor I_17975 (I307473,I307439,I46147);
nand I_17976 (I307490,I46144,I46135);
not I_17977 (I307507,I307490);
nand I_17978 (I307524,I307507,I307473);
nor I_17979 (I307541,I46123,I46126);
not I_17980 (I307558,I46138);
nor I_17981 (I307575,I307558,I46129);
nor I_17982 (I307294,I307575,I307408);
not I_17983 (I307606,I307575);
or I_17984 (I307309,I307524,I307575);
nor I_17985 (I307637,I307575,I307490);
nand I_17986 (I307306,I307439,I307637);
nor I_17987 (I307668,I307541,I307558);
nand I_17988 (I307685,I307507,I307668);
not I_17989 (I307312,I307685);
nor I_17990 (I307315,I307456,I307685);
or I_17991 (I307730,I307575,I307668);
nor I_17992 (I307300,I307507,I307730);
nor I_17993 (I307761,I307668,I46147);
nand I_17994 (I307778,I307761,I307507);
nand I_17995 (I307795,I307606,I307778);
DFFARX1 I_17996 (I307795,I1862,I307323,I307303,);
not I_17997 (I307850,I1869);
nor I_17998 (I307867,I20626,I20623);
not I_17999 (I307884,I20641);
not I_18000 (I307901,I20632);
nor I_18001 (I307918,I307901,I307867);
nand I_18002 (I307935,I307918,I20641);
not I_18003 (I307824,I307935);
nor I_18004 (I307966,I307901,I307884);
and I_18005 (I307983,I307935,I20647);
nor I_18006 (I308000,I307966,I20647);
nand I_18007 (I308017,I20644,I20635);
not I_18008 (I308034,I308017);
nand I_18009 (I308051,I308034,I308000);
nor I_18010 (I308068,I20623,I20626);
not I_18011 (I308085,I20638);
nor I_18012 (I308102,I308085,I20629);
nor I_18013 (I307821,I308102,I307935);
not I_18014 (I308133,I308102);
or I_18015 (I307836,I308051,I308102);
nor I_18016 (I308164,I308102,I308017);
nand I_18017 (I307833,I307966,I308164);
nor I_18018 (I308195,I308068,I308085);
nand I_18019 (I308212,I308034,I308195);
not I_18020 (I307839,I308212);
nor I_18021 (I307842,I307983,I308212);
or I_18022 (I308257,I308102,I308195);
nor I_18023 (I307827,I308034,I308257);
nor I_18024 (I308288,I308195,I20647);
nand I_18025 (I308305,I308288,I308034);
nand I_18026 (I308322,I308133,I308305);
DFFARX1 I_18027 (I308322,I1862,I307850,I307830,);
not I_18028 (I308377,I1869);
nor I_18029 (I308394,I57856,I57853);
not I_18030 (I308411,I57871);
not I_18031 (I308428,I57862);
nor I_18032 (I308445,I308428,I308394);
nand I_18033 (I308462,I308445,I57871);
not I_18034 (I308351,I308462);
nor I_18035 (I308493,I308428,I308411);
and I_18036 (I308510,I308462,I57877);
nor I_18037 (I308527,I308493,I57877);
nand I_18038 (I308544,I57874,I57865);
not I_18039 (I308561,I308544);
nand I_18040 (I308578,I308561,I308527);
nor I_18041 (I308595,I57853,I57856);
not I_18042 (I308612,I57868);
nor I_18043 (I308629,I308612,I57859);
nor I_18044 (I308348,I308629,I308462);
not I_18045 (I308660,I308629);
or I_18046 (I308363,I308578,I308629);
nor I_18047 (I308691,I308629,I308544);
nand I_18048 (I308360,I308493,I308691);
nor I_18049 (I308722,I308595,I308612);
nand I_18050 (I308739,I308561,I308722);
not I_18051 (I308366,I308739);
nor I_18052 (I308369,I308510,I308739);
or I_18053 (I308784,I308629,I308722);
nor I_18054 (I308354,I308561,I308784);
nor I_18055 (I308815,I308722,I57877);
nand I_18056 (I308832,I308815,I308561);
nand I_18057 (I308849,I308660,I308832);
DFFARX1 I_18058 (I308849,I1862,I308377,I308357,);
not I_18059 (I308904,I1869);
nor I_18060 (I308921,I146304,I146328);
not I_18061 (I308938,I146313);
not I_18062 (I308955,I146307);
nor I_18063 (I308972,I308955,I308921);
nand I_18064 (I308989,I308972,I146313);
not I_18065 (I308878,I308989);
nor I_18066 (I309020,I308955,I308938);
and I_18067 (I309037,I308989,I146310);
nor I_18068 (I309054,I309020,I146310);
nand I_18069 (I309071,I146304,I146319);
not I_18070 (I309088,I309071);
nand I_18071 (I309105,I309088,I309054);
nor I_18072 (I309122,I146316,I146307);
not I_18073 (I309139,I146325);
nor I_18074 (I309156,I309139,I146322);
nor I_18075 (I308875,I309156,I308989);
not I_18076 (I309187,I309156);
or I_18077 (I308890,I309105,I309156);
nor I_18078 (I309218,I309156,I309071);
nand I_18079 (I308887,I309020,I309218);
nor I_18080 (I309249,I309122,I309139);
nand I_18081 (I309266,I309088,I309249);
not I_18082 (I308893,I309266);
nor I_18083 (I308896,I309037,I309266);
or I_18084 (I309311,I309156,I309249);
nor I_18085 (I308881,I309088,I309311);
nor I_18086 (I309342,I309249,I146310);
nand I_18087 (I309359,I309342,I309088);
nand I_18088 (I309376,I309187,I309359);
DFFARX1 I_18089 (I309376,I1862,I308904,I308884,);
not I_18090 (I309431,I1869);
nor I_18091 (I309448,I25726,I25723);
not I_18092 (I309465,I25741);
not I_18093 (I309482,I25732);
nor I_18094 (I309499,I309482,I309448);
nand I_18095 (I309516,I309499,I25741);
not I_18096 (I309405,I309516);
nor I_18097 (I309547,I309482,I309465);
and I_18098 (I309564,I309516,I25747);
nor I_18099 (I309581,I309547,I25747);
nand I_18100 (I309598,I25744,I25735);
not I_18101 (I309615,I309598);
nand I_18102 (I309632,I309615,I309581);
nor I_18103 (I309649,I25723,I25726);
not I_18104 (I309666,I25738);
nor I_18105 (I309683,I309666,I25729);
nor I_18106 (I309402,I309683,I309516);
not I_18107 (I309714,I309683);
or I_18108 (I309417,I309632,I309683);
nor I_18109 (I309745,I309683,I309598);
nand I_18110 (I309414,I309547,I309745);
nor I_18111 (I309776,I309649,I309666);
nand I_18112 (I309793,I309615,I309776);
not I_18113 (I309420,I309793);
nor I_18114 (I309423,I309564,I309793);
or I_18115 (I309838,I309683,I309776);
nor I_18116 (I309408,I309615,I309838);
nor I_18117 (I309869,I309776,I25747);
nand I_18118 (I309886,I309869,I309615);
nand I_18119 (I309903,I309714,I309886);
DFFARX1 I_18120 (I309903,I1862,I309431,I309411,);
not I_18121 (I309958,I1869);
nor I_18122 (I309975,I266767,I266755);
not I_18123 (I309992,I266752);
not I_18124 (I310009,I266749);
nor I_18125 (I310026,I310009,I309975);
nand I_18126 (I310043,I310026,I266752);
not I_18127 (I309932,I310043);
nor I_18128 (I310074,I310009,I309992);
and I_18129 (I310091,I310043,I266752);
nor I_18130 (I310108,I310074,I266752);
nand I_18131 (I310125,I266755,I266761);
not I_18132 (I310142,I310125);
nand I_18133 (I310159,I310142,I310108);
nor I_18134 (I310176,I266770,I266764);
not I_18135 (I310193,I266758);
nor I_18136 (I310210,I310193,I266749);
nor I_18137 (I309929,I310210,I310043);
not I_18138 (I310241,I310210);
or I_18139 (I309944,I310159,I310210);
nor I_18140 (I310272,I310210,I310125);
nand I_18141 (I309941,I310074,I310272);
nor I_18142 (I310303,I310176,I310193);
nand I_18143 (I310320,I310142,I310303);
not I_18144 (I309947,I310320);
nor I_18145 (I309950,I310091,I310320);
or I_18146 (I310365,I310210,I310303);
nor I_18147 (I309935,I310142,I310365);
nor I_18148 (I310396,I310303,I266752);
nand I_18149 (I310413,I310396,I310142);
nand I_18150 (I310430,I310241,I310413);
DFFARX1 I_18151 (I310430,I1862,I309958,I309938,);
not I_18152 (I310485,I1869);
nor I_18153 (I310502,I371656,I371659);
not I_18154 (I310519,I371671);
not I_18155 (I310536,I371662);
nor I_18156 (I310553,I310536,I310502);
nand I_18157 (I310570,I310553,I371671);
not I_18158 (I310459,I310570);
nor I_18159 (I310601,I310536,I310519);
and I_18160 (I310618,I310570,I371665);
nor I_18161 (I310635,I310601,I371665);
nand I_18162 (I310652,I371662,I371668);
not I_18163 (I310669,I310652);
nand I_18164 (I310686,I310669,I310635);
nor I_18165 (I310703,I371659,I371674);
not I_18166 (I310720,I371665);
nor I_18167 (I310737,I310720,I371656);
nor I_18168 (I310456,I310737,I310570);
not I_18169 (I310768,I310737);
or I_18170 (I310471,I310686,I310737);
nor I_18171 (I310799,I310737,I310652);
nand I_18172 (I310468,I310601,I310799);
nor I_18173 (I310830,I310703,I310720);
nand I_18174 (I310847,I310669,I310830);
not I_18175 (I310474,I310847);
nor I_18176 (I310477,I310618,I310847);
or I_18177 (I310892,I310737,I310830);
nor I_18178 (I310462,I310669,I310892);
nor I_18179 (I310923,I310830,I371665);
nand I_18180 (I310940,I310923,I310669);
nand I_18181 (I310957,I310768,I310940);
DFFARX1 I_18182 (I310957,I1862,I310485,I310465,);
not I_18183 (I311012,I1869);
nor I_18184 (I311029,I94066,I94063);
not I_18185 (I311046,I94081);
not I_18186 (I311063,I94072);
nor I_18187 (I311080,I311063,I311029);
nand I_18188 (I311097,I311080,I94081);
not I_18189 (I310986,I311097);
nor I_18190 (I311128,I311063,I311046);
and I_18191 (I311145,I311097,I94087);
nor I_18192 (I311162,I311128,I94087);
nand I_18193 (I311179,I94084,I94075);
not I_18194 (I311196,I311179);
nand I_18195 (I311213,I311196,I311162);
nor I_18196 (I311230,I94063,I94066);
not I_18197 (I311247,I94078);
nor I_18198 (I311264,I311247,I94069);
nor I_18199 (I310983,I311264,I311097);
not I_18200 (I311295,I311264);
or I_18201 (I310998,I311213,I311264);
nor I_18202 (I311326,I311264,I311179);
nand I_18203 (I310995,I311128,I311326);
nor I_18204 (I311357,I311230,I311247);
nand I_18205 (I311374,I311196,I311357);
not I_18206 (I311001,I311374);
nor I_18207 (I311004,I311145,I311374);
or I_18208 (I311419,I311264,I311357);
nor I_18209 (I310989,I311196,I311419);
nor I_18210 (I311450,I311357,I94087);
nand I_18211 (I311467,I311450,I311196);
nand I_18212 (I311484,I311295,I311467);
DFFARX1 I_18213 (I311484,I1862,I311012,I310992,);
not I_18214 (I311539,I1869);
nor I_18215 (I311556,I122062,I122086);
not I_18216 (I311573,I122071);
not I_18217 (I311590,I122065);
nor I_18218 (I311607,I311590,I311556);
nand I_18219 (I311624,I311607,I122071);
not I_18220 (I311513,I311624);
nor I_18221 (I311655,I311590,I311573);
and I_18222 (I311672,I311624,I122068);
nor I_18223 (I311689,I311655,I122068);
nand I_18224 (I311706,I122062,I122077);
not I_18225 (I311723,I311706);
nand I_18226 (I311740,I311723,I311689);
nor I_18227 (I311757,I122074,I122065);
not I_18228 (I311774,I122083);
nor I_18229 (I311791,I311774,I122080);
nor I_18230 (I311510,I311791,I311624);
not I_18231 (I311822,I311791);
or I_18232 (I311525,I311740,I311791);
nor I_18233 (I311853,I311791,I311706);
nand I_18234 (I311522,I311655,I311853);
nor I_18235 (I311884,I311757,I311774);
nand I_18236 (I311901,I311723,I311884);
not I_18237 (I311528,I311901);
nor I_18238 (I311531,I311672,I311901);
or I_18239 (I311946,I311791,I311884);
nor I_18240 (I311516,I311723,I311946);
nor I_18241 (I311977,I311884,I122068);
nand I_18242 (I311994,I311977,I311723);
nand I_18243 (I312011,I311822,I311994);
DFFARX1 I_18244 (I312011,I1862,I311539,I311519,);
not I_18245 (I312066,I1869);
nor I_18246 (I312083,I280095,I280083);
not I_18247 (I312100,I280080);
not I_18248 (I312117,I280077);
nor I_18249 (I312134,I312117,I312083);
nand I_18250 (I312151,I312134,I280080);
not I_18251 (I312040,I312151);
nor I_18252 (I312182,I312117,I312100);
and I_18253 (I312199,I312151,I280080);
nor I_18254 (I312216,I312182,I280080);
nand I_18255 (I312233,I280083,I280089);
not I_18256 (I312250,I312233);
nand I_18257 (I312267,I312250,I312216);
nor I_18258 (I312284,I280098,I280092);
not I_18259 (I312301,I280086);
nor I_18260 (I312318,I312301,I280077);
nor I_18261 (I312037,I312318,I312151);
not I_18262 (I312349,I312318);
or I_18263 (I312052,I312267,I312318);
nor I_18264 (I312380,I312318,I312233);
nand I_18265 (I312049,I312182,I312380);
nor I_18266 (I312411,I312284,I312301);
nand I_18267 (I312428,I312250,I312411);
not I_18268 (I312055,I312428);
nor I_18269 (I312058,I312199,I312428);
or I_18270 (I312473,I312318,I312411);
nor I_18271 (I312043,I312250,I312473);
nor I_18272 (I312504,I312411,I280080);
nand I_18273 (I312521,I312504,I312250);
nand I_18274 (I312538,I312349,I312521);
DFFARX1 I_18275 (I312538,I1862,I312066,I312046,);
not I_18276 (I312593,I1869);
nor I_18277 (I312610,I37456,I37453);
not I_18278 (I312627,I37471);
not I_18279 (I312644,I37462);
nor I_18280 (I312661,I312644,I312610);
nand I_18281 (I312678,I312661,I37471);
not I_18282 (I312567,I312678);
nor I_18283 (I312709,I312644,I312627);
and I_18284 (I312726,I312678,I37477);
nor I_18285 (I312743,I312709,I37477);
nand I_18286 (I312760,I37474,I37465);
not I_18287 (I312777,I312760);
nand I_18288 (I312794,I312777,I312743);
nor I_18289 (I312811,I37453,I37456);
not I_18290 (I312828,I37468);
nor I_18291 (I312845,I312828,I37459);
nor I_18292 (I312564,I312845,I312678);
not I_18293 (I312876,I312845);
or I_18294 (I312579,I312794,I312845);
nor I_18295 (I312907,I312845,I312760);
nand I_18296 (I312576,I312709,I312907);
nor I_18297 (I312938,I312811,I312828);
nand I_18298 (I312955,I312777,I312938);
not I_18299 (I312582,I312955);
nor I_18300 (I312585,I312726,I312955);
or I_18301 (I313000,I312845,I312938);
nor I_18302 (I312570,I312777,I313000);
nor I_18303 (I313031,I312938,I37477);
nand I_18304 (I313048,I313031,I312777);
nand I_18305 (I313065,I312876,I313048);
DFFARX1 I_18306 (I313065,I1862,I312593,I312573,);
not I_18307 (I313120,I1869);
nor I_18308 (I313137,I247251,I247239);
not I_18309 (I313154,I247236);
not I_18310 (I313171,I247233);
nor I_18311 (I313188,I313171,I313137);
nand I_18312 (I313205,I313188,I247236);
not I_18313 (I313094,I313205);
nor I_18314 (I313236,I313171,I313154);
and I_18315 (I313253,I313205,I247236);
nor I_18316 (I313270,I313236,I247236);
nand I_18317 (I313287,I247239,I247245);
not I_18318 (I313304,I313287);
nand I_18319 (I313321,I313304,I313270);
nor I_18320 (I313338,I247254,I247248);
not I_18321 (I313355,I247242);
nor I_18322 (I313372,I313355,I247233);
nor I_18323 (I313091,I313372,I313205);
not I_18324 (I313403,I313372);
or I_18325 (I313106,I313321,I313372);
nor I_18326 (I313434,I313372,I313287);
nand I_18327 (I313103,I313236,I313434);
nor I_18328 (I313465,I313338,I313355);
nand I_18329 (I313482,I313304,I313465);
not I_18330 (I313109,I313482);
nor I_18331 (I313112,I313253,I313482);
or I_18332 (I313527,I313372,I313465);
nor I_18333 (I313097,I313304,I313527);
nor I_18334 (I313558,I313465,I247236);
nand I_18335 (I313575,I313558,I313304);
nand I_18336 (I313592,I313403,I313575);
DFFARX1 I_18337 (I313592,I1862,I313120,I313100,);
not I_18338 (I313647,I1869);
nor I_18339 (I313664,I41536,I41533);
not I_18340 (I313681,I41551);
not I_18341 (I313698,I41542);
nor I_18342 (I313715,I313698,I313664);
nand I_18343 (I313732,I313715,I41551);
not I_18344 (I313621,I313732);
nor I_18345 (I313763,I313698,I313681);
and I_18346 (I313780,I313732,I41557);
nor I_18347 (I313797,I313763,I41557);
nand I_18348 (I313814,I41554,I41545);
not I_18349 (I313831,I313814);
nand I_18350 (I313848,I313831,I313797);
nor I_18351 (I313865,I41533,I41536);
not I_18352 (I313882,I41548);
nor I_18353 (I313899,I313882,I41539);
nor I_18354 (I313618,I313899,I313732);
not I_18355 (I313930,I313899);
or I_18356 (I313633,I313848,I313899);
nor I_18357 (I313961,I313899,I313814);
nand I_18358 (I313630,I313763,I313961);
nor I_18359 (I313992,I313865,I313882);
nand I_18360 (I314009,I313831,I313992);
not I_18361 (I313636,I314009);
nor I_18362 (I313639,I313780,I314009);
or I_18363 (I314054,I313899,I313992);
nor I_18364 (I313624,I313831,I314054);
nor I_18365 (I314085,I313992,I41557);
nand I_18366 (I314102,I314085,I313831);
nand I_18367 (I314119,I313930,I314102);
DFFARX1 I_18368 (I314119,I1862,I313647,I313627,);
not I_18369 (I314174,I1869);
nor I_18370 (I314191,I89476,I89473);
not I_18371 (I314208,I89491);
not I_18372 (I314225,I89482);
nor I_18373 (I314242,I314225,I314191);
nand I_18374 (I314259,I314242,I89491);
not I_18375 (I314148,I314259);
nor I_18376 (I314290,I314225,I314208);
and I_18377 (I314307,I314259,I89497);
nor I_18378 (I314324,I314290,I89497);
nand I_18379 (I314341,I89494,I89485);
not I_18380 (I314358,I314341);
nand I_18381 (I314375,I314358,I314324);
nor I_18382 (I314392,I89473,I89476);
not I_18383 (I314409,I89488);
nor I_18384 (I314426,I314409,I89479);
nor I_18385 (I314145,I314426,I314259);
not I_18386 (I314457,I314426);
or I_18387 (I314160,I314375,I314426);
nor I_18388 (I314488,I314426,I314341);
nand I_18389 (I314157,I314290,I314488);
nor I_18390 (I314519,I314392,I314409);
nand I_18391 (I314536,I314358,I314519);
not I_18392 (I314163,I314536);
nor I_18393 (I314166,I314307,I314536);
or I_18394 (I314581,I314426,I314519);
nor I_18395 (I314151,I314358,I314581);
nor I_18396 (I314612,I314519,I89497);
nand I_18397 (I314629,I314612,I314358);
nand I_18398 (I314646,I314457,I314629);
DFFARX1 I_18399 (I314646,I1862,I314174,I314154,);
not I_18400 (I314701,I1869);
nor I_18401 (I314718,I58366,I58363);
not I_18402 (I314735,I58381);
not I_18403 (I314752,I58372);
nor I_18404 (I314769,I314752,I314718);
nand I_18405 (I314786,I314769,I58381);
not I_18406 (I314675,I314786);
nor I_18407 (I314817,I314752,I314735);
and I_18408 (I314834,I314786,I58387);
nor I_18409 (I314851,I314817,I58387);
nand I_18410 (I314868,I58384,I58375);
not I_18411 (I314885,I314868);
nand I_18412 (I314902,I314885,I314851);
nor I_18413 (I314919,I58363,I58366);
not I_18414 (I314936,I58378);
nor I_18415 (I314953,I314936,I58369);
nor I_18416 (I314672,I314953,I314786);
not I_18417 (I314984,I314953);
or I_18418 (I314687,I314902,I314953);
nor I_18419 (I315015,I314953,I314868);
nand I_18420 (I314684,I314817,I315015);
nor I_18421 (I315046,I314919,I314936);
nand I_18422 (I315063,I314885,I315046);
not I_18423 (I314690,I315063);
nor I_18424 (I314693,I314834,I315063);
or I_18425 (I315108,I314953,I315046);
nor I_18426 (I314678,I314885,I315108);
nor I_18427 (I315139,I315046,I58387);
nand I_18428 (I315156,I315139,I314885);
nand I_18429 (I315173,I314984,I315156);
DFFARX1 I_18430 (I315173,I1862,I314701,I314681,);
not I_18431 (I315228,I1869);
nor I_18432 (I315245,I379612,I379615);
not I_18433 (I315262,I379627);
not I_18434 (I315279,I379618);
nor I_18435 (I315296,I315279,I315245);
nand I_18436 (I315313,I315296,I379627);
not I_18437 (I315202,I315313);
nor I_18438 (I315344,I315279,I315262);
and I_18439 (I315361,I315313,I379621);
nor I_18440 (I315378,I315344,I379621);
nand I_18441 (I315395,I379618,I379624);
not I_18442 (I315412,I315395);
nand I_18443 (I315429,I315412,I315378);
nor I_18444 (I315446,I379615,I379630);
not I_18445 (I315463,I379621);
nor I_18446 (I315480,I315463,I379612);
nor I_18447 (I315199,I315480,I315313);
not I_18448 (I315511,I315480);
or I_18449 (I315214,I315429,I315480);
nor I_18450 (I315542,I315480,I315395);
nand I_18451 (I315211,I315344,I315542);
nor I_18452 (I315573,I315446,I315463);
nand I_18453 (I315590,I315412,I315573);
not I_18454 (I315217,I315590);
nor I_18455 (I315220,I315361,I315590);
or I_18456 (I315635,I315480,I315573);
nor I_18457 (I315205,I315412,I315635);
nor I_18458 (I315666,I315573,I379621);
nand I_18459 (I315683,I315666,I315412);
nand I_18460 (I315700,I315511,I315683);
DFFARX1 I_18461 (I315700,I1862,I315228,I315208,);
not I_18462 (I315755,I1869);
nor I_18463 (I315772,I83866,I83863);
not I_18464 (I315789,I83881);
not I_18465 (I315806,I83872);
nor I_18466 (I315823,I315806,I315772);
nand I_18467 (I315840,I315823,I83881);
not I_18468 (I315729,I315840);
nor I_18469 (I315871,I315806,I315789);
and I_18470 (I315888,I315840,I83887);
nor I_18471 (I315905,I315871,I83887);
nand I_18472 (I315922,I83884,I83875);
not I_18473 (I315939,I315922);
nand I_18474 (I315956,I315939,I315905);
nor I_18475 (I315973,I83863,I83866);
not I_18476 (I315990,I83878);
nor I_18477 (I316007,I315990,I83869);
nor I_18478 (I315726,I316007,I315840);
not I_18479 (I316038,I316007);
or I_18480 (I315741,I315956,I316007);
nor I_18481 (I316069,I316007,I315922);
nand I_18482 (I315738,I315871,I316069);
nor I_18483 (I316100,I315973,I315990);
nand I_18484 (I316117,I315939,I316100);
not I_18485 (I315744,I316117);
nor I_18486 (I315747,I315888,I316117);
or I_18487 (I316162,I316007,I316100);
nor I_18488 (I315732,I315939,I316162);
nor I_18489 (I316193,I316100,I83887);
nand I_18490 (I316210,I316193,I315939);
nand I_18491 (I316227,I316038,I316210);
DFFARX1 I_18492 (I316227,I1862,I315755,I315735,);
not I_18493 (I316282,I1869);
nor I_18494 (I316299,I300973,I300970);
not I_18495 (I316316,I300979);
not I_18496 (I316333,I300976);
nor I_18497 (I316350,I316333,I316299);
nand I_18498 (I316367,I316350,I300979);
not I_18499 (I316256,I316367);
nor I_18500 (I316398,I316333,I316316);
and I_18501 (I316415,I316367,I300982);
nor I_18502 (I316432,I316398,I300982);
nand I_18503 (I316449,I300985,I300976);
not I_18504 (I316466,I316449);
nand I_18505 (I316483,I316466,I316432);
nor I_18506 (I316500,I300991,I300988);
not I_18507 (I316517,I300970);
nor I_18508 (I316534,I316517,I300973);
nor I_18509 (I316253,I316534,I316367);
not I_18510 (I316565,I316534);
or I_18511 (I316268,I316483,I316534);
nor I_18512 (I316596,I316534,I316449);
nand I_18513 (I316265,I316398,I316596);
nor I_18514 (I316627,I316500,I316517);
nand I_18515 (I316644,I316466,I316627);
not I_18516 (I316271,I316644);
nor I_18517 (I316274,I316415,I316644);
or I_18518 (I316689,I316534,I316627);
nor I_18519 (I316259,I316466,I316689);
nor I_18520 (I316720,I316627,I300982);
nand I_18521 (I316737,I316720,I316466);
nand I_18522 (I316754,I316565,I316737);
DFFARX1 I_18523 (I316754,I1862,I316282,I316262,);
not I_18524 (I316809,I1869);
nor I_18525 (I316826,I24196,I24193);
not I_18526 (I316843,I24211);
not I_18527 (I316860,I24202);
nor I_18528 (I316877,I316860,I316826);
nand I_18529 (I316894,I316877,I24211);
not I_18530 (I316783,I316894);
nor I_18531 (I316925,I316860,I316843);
and I_18532 (I316942,I316894,I24217);
nor I_18533 (I316959,I316925,I24217);
nand I_18534 (I316976,I24214,I24205);
not I_18535 (I316993,I316976);
nand I_18536 (I317010,I316993,I316959);
nor I_18537 (I317027,I24193,I24196);
not I_18538 (I317044,I24208);
nor I_18539 (I317061,I317044,I24199);
nor I_18540 (I316780,I317061,I316894);
not I_18541 (I317092,I317061);
or I_18542 (I316795,I317010,I317061);
nor I_18543 (I317123,I317061,I316976);
nand I_18544 (I316792,I316925,I317123);
nor I_18545 (I317154,I317027,I317044);
nand I_18546 (I317171,I316993,I317154);
not I_18547 (I316798,I317171);
nor I_18548 (I316801,I316942,I317171);
or I_18549 (I317216,I317061,I317154);
nor I_18550 (I316786,I316993,I317216);
nor I_18551 (I317247,I317154,I24217);
nand I_18552 (I317264,I317247,I316993);
nand I_18553 (I317281,I317092,I317264);
DFFARX1 I_18554 (I317281,I1862,I316809,I316789,);
not I_18555 (I317336,I1869);
nor I_18556 (I317353,I34396,I34393);
not I_18557 (I317370,I34411);
not I_18558 (I317387,I34402);
nor I_18559 (I317404,I317387,I317353);
nand I_18560 (I317421,I317404,I34411);
not I_18561 (I317310,I317421);
nor I_18562 (I317452,I317387,I317370);
and I_18563 (I317469,I317421,I34417);
nor I_18564 (I317486,I317452,I34417);
nand I_18565 (I317503,I34414,I34405);
not I_18566 (I317520,I317503);
nand I_18567 (I317537,I317520,I317486);
nor I_18568 (I317554,I34393,I34396);
not I_18569 (I317571,I34408);
nor I_18570 (I317588,I317571,I34399);
nor I_18571 (I317307,I317588,I317421);
not I_18572 (I317619,I317588);
or I_18573 (I317322,I317537,I317588);
nor I_18574 (I317650,I317588,I317503);
nand I_18575 (I317319,I317452,I317650);
nor I_18576 (I317681,I317554,I317571);
nand I_18577 (I317698,I317520,I317681);
not I_18578 (I317325,I317698);
nor I_18579 (I317328,I317469,I317698);
or I_18580 (I317743,I317588,I317681);
nor I_18581 (I317313,I317520,I317743);
nor I_18582 (I317774,I317681,I34417);
nand I_18583 (I317791,I317774,I317520);
nand I_18584 (I317808,I317619,I317791);
DFFARX1 I_18585 (I317808,I1862,I317336,I317316,);
not I_18586 (I317863,I1869);
nor I_18587 (I317880,I157371,I157395);
not I_18588 (I317897,I157380);
not I_18589 (I317914,I157374);
nor I_18590 (I317931,I317914,I317880);
nand I_18591 (I317948,I317931,I157380);
not I_18592 (I317837,I317948);
nor I_18593 (I317979,I317914,I317897);
and I_18594 (I317996,I317948,I157377);
nor I_18595 (I318013,I317979,I157377);
nand I_18596 (I318030,I157371,I157386);
not I_18597 (I318047,I318030);
nand I_18598 (I318064,I318047,I318013);
nor I_18599 (I318081,I157383,I157374);
not I_18600 (I318098,I157392);
nor I_18601 (I318115,I318098,I157389);
nor I_18602 (I317834,I318115,I317948);
not I_18603 (I318146,I318115);
or I_18604 (I317849,I318064,I318115);
nor I_18605 (I318177,I318115,I318030);
nand I_18606 (I317846,I317979,I318177);
nor I_18607 (I318208,I318081,I318098);
nand I_18608 (I318225,I318047,I318208);
not I_18609 (I317852,I318225);
nor I_18610 (I317855,I317996,I318225);
or I_18611 (I318270,I318115,I318208);
nor I_18612 (I317840,I318047,I318270);
nor I_18613 (I318301,I318208,I157377);
nand I_18614 (I318318,I318301,I318047);
nand I_18615 (I318335,I318146,I318318);
DFFARX1 I_18616 (I318335,I1862,I317863,I317843,);
not I_18617 (I318390,I1869);
nor I_18618 (I318407,I270099,I270087);
not I_18619 (I318424,I270084);
not I_18620 (I318441,I270081);
nor I_18621 (I318458,I318441,I318407);
nand I_18622 (I318475,I318458,I270084);
not I_18623 (I318364,I318475);
nor I_18624 (I318506,I318441,I318424);
and I_18625 (I318523,I318475,I270084);
nor I_18626 (I318540,I318506,I270084);
nand I_18627 (I318557,I270087,I270093);
not I_18628 (I318574,I318557);
nand I_18629 (I318591,I318574,I318540);
nor I_18630 (I318608,I270102,I270096);
not I_18631 (I318625,I270090);
nor I_18632 (I318642,I318625,I270081);
nor I_18633 (I318361,I318642,I318475);
not I_18634 (I318673,I318642);
or I_18635 (I318376,I318591,I318642);
nor I_18636 (I318704,I318642,I318557);
nand I_18637 (I318373,I318506,I318704);
nor I_18638 (I318735,I318608,I318625);
nand I_18639 (I318752,I318574,I318735);
not I_18640 (I318379,I318752);
nor I_18641 (I318382,I318523,I318752);
or I_18642 (I318797,I318642,I318735);
nor I_18643 (I318367,I318574,I318797);
nor I_18644 (I318828,I318735,I270084);
nand I_18645 (I318845,I318828,I318574);
nand I_18646 (I318862,I318673,I318845);
DFFARX1 I_18647 (I318862,I1862,I318390,I318370,);
not I_18648 (I318917,I1869);
nor I_18649 (I318934,I52756,I52753);
not I_18650 (I318951,I52771);
not I_18651 (I318968,I52762);
nor I_18652 (I318985,I318968,I318934);
nand I_18653 (I319002,I318985,I52771);
not I_18654 (I318891,I319002);
nor I_18655 (I319033,I318968,I318951);
and I_18656 (I319050,I319002,I52777);
nor I_18657 (I319067,I319033,I52777);
nand I_18658 (I319084,I52774,I52765);
not I_18659 (I319101,I319084);
nand I_18660 (I319118,I319101,I319067);
nor I_18661 (I319135,I52753,I52756);
not I_18662 (I319152,I52768);
nor I_18663 (I319169,I319152,I52759);
nor I_18664 (I318888,I319169,I319002);
not I_18665 (I319200,I319169);
or I_18666 (I318903,I319118,I319169);
nor I_18667 (I319231,I319169,I319084);
nand I_18668 (I318900,I319033,I319231);
nor I_18669 (I319262,I319135,I319152);
nand I_18670 (I319279,I319101,I319262);
not I_18671 (I318906,I319279);
nor I_18672 (I318909,I319050,I319279);
or I_18673 (I319324,I319169,I319262);
nor I_18674 (I318894,I319101,I319324);
nor I_18675 (I319355,I319262,I52777);
nand I_18676 (I319372,I319355,I319101);
nand I_18677 (I319389,I319200,I319372);
DFFARX1 I_18678 (I319389,I1862,I318917,I318897,);
not I_18679 (I319444,I1869);
nor I_18680 (I319461,I102226,I102241);
not I_18681 (I319478,I102229);
not I_18682 (I319495,I102223);
nor I_18683 (I319512,I319495,I319461);
nand I_18684 (I319529,I319512,I102229);
not I_18685 (I319418,I319529);
nor I_18686 (I319560,I319495,I319478);
and I_18687 (I319577,I319529,I102238);
nor I_18688 (I319594,I319560,I102238);
nand I_18689 (I319611,I102223,I102232);
not I_18690 (I319628,I319611);
nand I_18691 (I319645,I319628,I319594);
nor I_18692 (I319662,I102235,I102226);
not I_18693 (I319679,I102229);
nor I_18694 (I319696,I319679,I102232);
nor I_18695 (I319415,I319696,I319529);
not I_18696 (I319727,I319696);
or I_18697 (I319430,I319645,I319696);
nor I_18698 (I319758,I319696,I319611);
nand I_18699 (I319427,I319560,I319758);
nor I_18700 (I319789,I319662,I319679);
nand I_18701 (I319806,I319628,I319789);
not I_18702 (I319433,I319806);
nor I_18703 (I319436,I319577,I319806);
or I_18704 (I319851,I319696,I319789);
nor I_18705 (I319421,I319628,I319851);
nor I_18706 (I319882,I319789,I102238);
nand I_18707 (I319899,I319882,I319628);
nand I_18708 (I319916,I319727,I319899);
DFFARX1 I_18709 (I319916,I1862,I319444,I319424,);
not I_18710 (I319971,I1869);
nor I_18711 (I319988,I236779,I236767);
not I_18712 (I320005,I236764);
not I_18713 (I320022,I236761);
nor I_18714 (I320039,I320022,I319988);
nand I_18715 (I320056,I320039,I236764);
not I_18716 (I319945,I320056);
nor I_18717 (I320087,I320022,I320005);
and I_18718 (I320104,I320056,I236764);
nor I_18719 (I320121,I320087,I236764);
nand I_18720 (I320138,I236767,I236773);
not I_18721 (I320155,I320138);
nand I_18722 (I320172,I320155,I320121);
nor I_18723 (I320189,I236782,I236776);
not I_18724 (I320206,I236770);
nor I_18725 (I320223,I320206,I236761);
nor I_18726 (I319942,I320223,I320056);
not I_18727 (I320254,I320223);
or I_18728 (I319957,I320172,I320223);
nor I_18729 (I320285,I320223,I320138);
nand I_18730 (I319954,I320087,I320285);
nor I_18731 (I320316,I320189,I320206);
nand I_18732 (I320333,I320155,I320316);
not I_18733 (I319960,I320333);
nor I_18734 (I319963,I320104,I320333);
or I_18735 (I320378,I320223,I320316);
nor I_18736 (I319948,I320155,I320378);
nor I_18737 (I320409,I320316,I236764);
nand I_18738 (I320426,I320409,I320155);
nand I_18739 (I320443,I320254,I320426);
DFFARX1 I_18740 (I320443,I1862,I319971,I319951,);
not I_18741 (I320498,I1869);
nor I_18742 (I320515,I150520,I150544);
not I_18743 (I320532,I150529);
not I_18744 (I320549,I150523);
nor I_18745 (I320566,I320549,I320515);
nand I_18746 (I320583,I320566,I150529);
not I_18747 (I320472,I320583);
nor I_18748 (I320614,I320549,I320532);
and I_18749 (I320631,I320583,I150526);
nor I_18750 (I320648,I320614,I150526);
nand I_18751 (I320665,I150520,I150535);
not I_18752 (I320682,I320665);
nand I_18753 (I320699,I320682,I320648);
nor I_18754 (I320716,I150532,I150523);
not I_18755 (I320733,I150541);
nor I_18756 (I320750,I320733,I150538);
nor I_18757 (I320469,I320750,I320583);
not I_18758 (I320781,I320750);
or I_18759 (I320484,I320699,I320750);
nor I_18760 (I320812,I320750,I320665);
nand I_18761 (I320481,I320614,I320812);
nor I_18762 (I320843,I320716,I320733);
nand I_18763 (I320860,I320682,I320843);
not I_18764 (I320487,I320860);
nor I_18765 (I320490,I320631,I320860);
or I_18766 (I320905,I320750,I320843);
nor I_18767 (I320475,I320682,I320905);
nor I_18768 (I320936,I320843,I150526);
nand I_18769 (I320953,I320936,I320682);
nand I_18770 (I320970,I320781,I320953);
DFFARX1 I_18771 (I320970,I1862,I320498,I320478,);
not I_18772 (I321025,I1869);
nor I_18773 (I321042,I96616,I96613);
not I_18774 (I321059,I96631);
not I_18775 (I321076,I96622);
nor I_18776 (I321093,I321076,I321042);
nand I_18777 (I321110,I321093,I96631);
not I_18778 (I320999,I321110);
nor I_18779 (I321141,I321076,I321059);
and I_18780 (I321158,I321110,I96637);
nor I_18781 (I321175,I321141,I96637);
nand I_18782 (I321192,I96634,I96625);
not I_18783 (I321209,I321192);
nand I_18784 (I321226,I321209,I321175);
nor I_18785 (I321243,I96613,I96616);
not I_18786 (I321260,I96628);
nor I_18787 (I321277,I321260,I96619);
nor I_18788 (I320996,I321277,I321110);
not I_18789 (I321308,I321277);
or I_18790 (I321011,I321226,I321277);
nor I_18791 (I321339,I321277,I321192);
nand I_18792 (I321008,I321141,I321339);
nor I_18793 (I321370,I321243,I321260);
nand I_18794 (I321387,I321209,I321370);
not I_18795 (I321014,I321387);
nor I_18796 (I321017,I321158,I321387);
or I_18797 (I321432,I321277,I321370);
nor I_18798 (I321002,I321209,I321432);
nor I_18799 (I321463,I321370,I96637);
nand I_18800 (I321480,I321463,I321209);
nand I_18801 (I321497,I321308,I321480);
DFFARX1 I_18802 (I321497,I1862,I321025,I321005,);
not I_18803 (I321552,I1869);
nor I_18804 (I321569,I136291,I136315);
not I_18805 (I321586,I136300);
not I_18806 (I321603,I136294);
nor I_18807 (I321620,I321603,I321569);
nand I_18808 (I321637,I321620,I136300);
not I_18809 (I321526,I321637);
nor I_18810 (I321668,I321603,I321586);
and I_18811 (I321685,I321637,I136297);
nor I_18812 (I321702,I321668,I136297);
nand I_18813 (I321719,I136291,I136306);
not I_18814 (I321736,I321719);
nand I_18815 (I321753,I321736,I321702);
nor I_18816 (I321770,I136303,I136294);
not I_18817 (I321787,I136312);
nor I_18818 (I321804,I321787,I136309);
nor I_18819 (I321523,I321804,I321637);
not I_18820 (I321835,I321804);
or I_18821 (I321538,I321753,I321804);
nor I_18822 (I321866,I321804,I321719);
nand I_18823 (I321535,I321668,I321866);
nor I_18824 (I321897,I321770,I321787);
nand I_18825 (I321914,I321736,I321897);
not I_18826 (I321541,I321914);
nor I_18827 (I321544,I321685,I321914);
or I_18828 (I321959,I321804,I321897);
nor I_18829 (I321529,I321736,I321959);
nor I_18830 (I321990,I321897,I136297);
nand I_18831 (I322007,I321990,I321736);
nand I_18832 (I322024,I321835,I322007);
DFFARX1 I_18833 (I322024,I1862,I321552,I321532,);
not I_18834 (I322079,I1869);
nor I_18835 (I322096,I237731,I237719);
not I_18836 (I322113,I237716);
not I_18837 (I322130,I237713);
nor I_18838 (I322147,I322130,I322096);
nand I_18839 (I322164,I322147,I237716);
not I_18840 (I322053,I322164);
nor I_18841 (I322195,I322130,I322113);
and I_18842 (I322212,I322164,I237716);
nor I_18843 (I322229,I322195,I237716);
nand I_18844 (I322246,I237719,I237725);
not I_18845 (I322263,I322246);
nand I_18846 (I322280,I322263,I322229);
nor I_18847 (I322297,I237734,I237728);
not I_18848 (I322314,I237722);
nor I_18849 (I322331,I322314,I237713);
nor I_18850 (I322050,I322331,I322164);
not I_18851 (I322362,I322331);
or I_18852 (I322065,I322280,I322331);
nor I_18853 (I322393,I322331,I322246);
nand I_18854 (I322062,I322195,I322393);
nor I_18855 (I322424,I322297,I322314);
nand I_18856 (I322441,I322263,I322424);
not I_18857 (I322068,I322441);
nor I_18858 (I322071,I322212,I322441);
or I_18859 (I322486,I322331,I322424);
nor I_18860 (I322056,I322263,I322486);
nor I_18861 (I322517,I322424,I237716);
nand I_18862 (I322534,I322517,I322263);
nand I_18863 (I322551,I322362,I322534);
DFFARX1 I_18864 (I322551,I1862,I322079,I322059,);
not I_18865 (I322606,I1869);
nor I_18866 (I322623,I224403,I224391);
not I_18867 (I322640,I224388);
not I_18868 (I322657,I224385);
nor I_18869 (I322674,I322657,I322623);
nand I_18870 (I322691,I322674,I224388);
not I_18871 (I322580,I322691);
nor I_18872 (I322722,I322657,I322640);
and I_18873 (I322739,I322691,I224388);
nor I_18874 (I322756,I322722,I224388);
nand I_18875 (I322773,I224391,I224397);
not I_18876 (I322790,I322773);
nand I_18877 (I322807,I322790,I322756);
nor I_18878 (I322824,I224406,I224400);
not I_18879 (I322841,I224394);
nor I_18880 (I322858,I322841,I224385);
nor I_18881 (I322577,I322858,I322691);
not I_18882 (I322889,I322858);
or I_18883 (I322592,I322807,I322858);
nor I_18884 (I322920,I322858,I322773);
nand I_18885 (I322589,I322722,I322920);
nor I_18886 (I322951,I322824,I322841);
nand I_18887 (I322968,I322790,I322951);
not I_18888 (I322595,I322968);
nor I_18889 (I322598,I322739,I322968);
or I_18890 (I323013,I322858,I322951);
nor I_18891 (I322583,I322790,I323013);
nor I_18892 (I323044,I322951,I224388);
nand I_18893 (I323061,I323044,I322790);
nand I_18894 (I323078,I322889,I323061);
DFFARX1 I_18895 (I323078,I1862,I322606,I322586,);
not I_18896 (I323133,I1869);
nor I_18897 (I323150,I392430,I392433);
not I_18898 (I323167,I392445);
not I_18899 (I323184,I392436);
nor I_18900 (I323201,I323184,I323150);
nand I_18901 (I323218,I323201,I392445);
not I_18902 (I323107,I323218);
nor I_18903 (I323249,I323184,I323167);
and I_18904 (I323266,I323218,I392439);
nor I_18905 (I323283,I323249,I392439);
nand I_18906 (I323300,I392436,I392442);
not I_18907 (I323317,I323300);
nand I_18908 (I323334,I323317,I323283);
nor I_18909 (I323351,I392433,I392448);
not I_18910 (I323368,I392439);
nor I_18911 (I323385,I323368,I392430);
nor I_18912 (I323104,I323385,I323218);
not I_18913 (I323416,I323385);
or I_18914 (I323119,I323334,I323385);
nor I_18915 (I323447,I323385,I323300);
nand I_18916 (I323116,I323249,I323447);
nor I_18917 (I323478,I323351,I323368);
nand I_18918 (I323495,I323317,I323478);
not I_18919 (I323122,I323495);
nor I_18920 (I323125,I323266,I323495);
or I_18921 (I323540,I323385,I323478);
nor I_18922 (I323110,I323317,I323540);
nor I_18923 (I323571,I323478,I392439);
nand I_18924 (I323588,I323571,I323317);
nand I_18925 (I323605,I323416,I323588);
DFFARX1 I_18926 (I323605,I1862,I323133,I323113,);
not I_18927 (I323660,I1869);
nor I_18928 (I323677,I287798,I287795);
not I_18929 (I323694,I287804);
not I_18930 (I323711,I287801);
nor I_18931 (I323728,I323711,I323677);
nand I_18932 (I323745,I323728,I287804);
not I_18933 (I323634,I323745);
nor I_18934 (I323776,I323711,I323694);
and I_18935 (I323793,I323745,I287807);
nor I_18936 (I323810,I323776,I287807);
nand I_18937 (I323827,I287810,I287801);
not I_18938 (I323844,I323827);
nand I_18939 (I323861,I323844,I323810);
nor I_18940 (I323878,I287816,I287813);
not I_18941 (I323895,I287795);
nor I_18942 (I323912,I323895,I287798);
nor I_18943 (I323631,I323912,I323745);
not I_18944 (I323943,I323912);
or I_18945 (I323646,I323861,I323912);
nor I_18946 (I323974,I323912,I323827);
nand I_18947 (I323643,I323776,I323974);
nor I_18948 (I324005,I323878,I323895);
nand I_18949 (I324022,I323844,I324005);
not I_18950 (I323649,I324022);
nor I_18951 (I323652,I323793,I324022);
or I_18952 (I324067,I323912,I324005);
nor I_18953 (I323637,I323844,I324067);
nor I_18954 (I324098,I324005,I287807);
nand I_18955 (I324115,I324098,I323844);
nand I_18956 (I324132,I323943,I324115);
DFFARX1 I_18957 (I324132,I1862,I323660,I323640,);
not I_18958 (I324187,I1869);
nor I_18959 (I324204,I391104,I391107);
not I_18960 (I324221,I391119);
not I_18961 (I324238,I391110);
nor I_18962 (I324255,I324238,I324204);
nand I_18963 (I324272,I324255,I391119);
not I_18964 (I324161,I324272);
nor I_18965 (I324303,I324238,I324221);
and I_18966 (I324320,I324272,I391113);
nor I_18967 (I324337,I324303,I391113);
nand I_18968 (I324354,I391110,I391116);
not I_18969 (I324371,I324354);
nand I_18970 (I324388,I324371,I324337);
nor I_18971 (I324405,I391107,I391122);
not I_18972 (I324422,I391113);
nor I_18973 (I324439,I324422,I391104);
nor I_18974 (I324158,I324439,I324272);
not I_18975 (I324470,I324439);
or I_18976 (I324173,I324388,I324439);
nor I_18977 (I324501,I324439,I324354);
nand I_18978 (I324170,I324303,I324501);
nor I_18979 (I324532,I324405,I324422);
nand I_18980 (I324549,I324371,I324532);
not I_18981 (I324176,I324549);
nor I_18982 (I324179,I324320,I324549);
or I_18983 (I324594,I324439,I324532);
nor I_18984 (I324164,I324371,I324594);
nor I_18985 (I324625,I324532,I391113);
nand I_18986 (I324642,I324625,I324371);
nand I_18987 (I324659,I324470,I324642);
DFFARX1 I_18988 (I324659,I1862,I324187,I324167,);
not I_18989 (I324714,I1869);
nor I_18990 (I324731,I104266,I104281);
not I_18991 (I324748,I104269);
not I_18992 (I324765,I104263);
nor I_18993 (I324782,I324765,I324731);
nand I_18994 (I324799,I324782,I104269);
not I_18995 (I324688,I324799);
nor I_18996 (I324830,I324765,I324748);
and I_18997 (I324847,I324799,I104278);
nor I_18998 (I324864,I324830,I104278);
nand I_18999 (I324881,I104263,I104272);
not I_19000 (I324898,I324881);
nand I_19001 (I324915,I324898,I324864);
nor I_19002 (I324932,I104275,I104266);
not I_19003 (I324949,I104269);
nor I_19004 (I324966,I324949,I104272);
nor I_19005 (I324685,I324966,I324799);
not I_19006 (I324997,I324966);
or I_19007 (I324700,I324915,I324966);
nor I_19008 (I325028,I324966,I324881);
nand I_19009 (I324697,I324830,I325028);
nor I_19010 (I325059,I324932,I324949);
nand I_19011 (I325076,I324898,I325059);
not I_19012 (I324703,I325076);
nor I_19013 (I324706,I324847,I325076);
or I_19014 (I325121,I324966,I325059);
nor I_19015 (I324691,I324898,I325121);
nor I_19016 (I325152,I325059,I104278);
nand I_19017 (I325169,I325152,I324898);
nand I_19018 (I325186,I324997,I325169);
DFFARX1 I_19019 (I325186,I1862,I324714,I324694,);
not I_19020 (I325241,I1869);
nor I_19021 (I325258,I236303,I236291);
not I_19022 (I325275,I236288);
not I_19023 (I325292,I236285);
nor I_19024 (I325309,I325292,I325258);
nand I_19025 (I325326,I325309,I236288);
not I_19026 (I325215,I325326);
nor I_19027 (I325357,I325292,I325275);
and I_19028 (I325374,I325326,I236288);
nor I_19029 (I325391,I325357,I236288);
nand I_19030 (I325408,I236291,I236297);
not I_19031 (I325425,I325408);
nand I_19032 (I325442,I325425,I325391);
nor I_19033 (I325459,I236306,I236300);
not I_19034 (I325476,I236294);
nor I_19035 (I325493,I325476,I236285);
nor I_19036 (I325212,I325493,I325326);
not I_19037 (I325524,I325493);
or I_19038 (I325227,I325442,I325493);
nor I_19039 (I325555,I325493,I325408);
nand I_19040 (I325224,I325357,I325555);
nor I_19041 (I325586,I325459,I325476);
nand I_19042 (I325603,I325425,I325586);
not I_19043 (I325230,I325603);
nor I_19044 (I325233,I325374,I325603);
or I_19045 (I325648,I325493,I325586);
nor I_19046 (I325218,I325425,I325648);
nor I_19047 (I325679,I325586,I236288);
nand I_19048 (I325696,I325679,I325425);
nand I_19049 (I325713,I325524,I325696);
DFFARX1 I_19050 (I325713,I1862,I325241,I325221,);
not I_19051 (I325768,I1869);
nor I_19052 (I325785,I252963,I252951);
not I_19053 (I325802,I252948);
not I_19054 (I325819,I252945);
nor I_19055 (I325836,I325819,I325785);
nand I_19056 (I325853,I325836,I252948);
not I_19057 (I325742,I325853);
nor I_19058 (I325884,I325819,I325802);
and I_19059 (I325901,I325853,I252948);
nor I_19060 (I325918,I325884,I252948);
nand I_19061 (I325935,I252951,I252957);
not I_19062 (I325952,I325935);
nand I_19063 (I325969,I325952,I325918);
nor I_19064 (I325986,I252966,I252960);
not I_19065 (I326003,I252954);
nor I_19066 (I326020,I326003,I252945);
nor I_19067 (I325739,I326020,I325853);
not I_19068 (I326051,I326020);
or I_19069 (I325754,I325969,I326020);
nor I_19070 (I326082,I326020,I325935);
nand I_19071 (I325751,I325884,I326082);
nor I_19072 (I326113,I325986,I326003);
nand I_19073 (I326130,I325952,I326113);
not I_19074 (I325757,I326130);
nor I_19075 (I325760,I325901,I326130);
or I_19076 (I326175,I326020,I326113);
nor I_19077 (I325745,I325952,I326175);
nor I_19078 (I326206,I326113,I252948);
nand I_19079 (I326223,I326206,I325952);
nand I_19080 (I326240,I326051,I326223);
DFFARX1 I_19081 (I326240,I1862,I325768,I325748,);
not I_19082 (I326295,I1869);
nor I_19083 (I326312,I367236,I367239);
not I_19084 (I326329,I367251);
not I_19085 (I326346,I367242);
nor I_19086 (I326363,I326346,I326312);
nand I_19087 (I326380,I326363,I367251);
not I_19088 (I326269,I326380);
nor I_19089 (I326411,I326346,I326329);
and I_19090 (I326428,I326380,I367245);
nor I_19091 (I326445,I326411,I367245);
nand I_19092 (I326462,I367242,I367248);
not I_19093 (I326479,I326462);
nand I_19094 (I326496,I326479,I326445);
nor I_19095 (I326513,I367239,I367254);
not I_19096 (I326530,I367245);
nor I_19097 (I326547,I326530,I367236);
nor I_19098 (I326266,I326547,I326380);
not I_19099 (I326578,I326547);
or I_19100 (I326281,I326496,I326547);
nor I_19101 (I326609,I326547,I326462);
nand I_19102 (I326278,I326411,I326609);
nor I_19103 (I326640,I326513,I326530);
nand I_19104 (I326657,I326479,I326640);
not I_19105 (I326284,I326657);
nor I_19106 (I326287,I326428,I326657);
or I_19107 (I326702,I326547,I326640);
nor I_19108 (I326272,I326479,I326702);
nor I_19109 (I326733,I326640,I367245);
nand I_19110 (I326750,I326733,I326479);
nand I_19111 (I326767,I326578,I326750);
DFFARX1 I_19112 (I326767,I1862,I326295,I326275,);
not I_19113 (I326822,I1869);
nor I_19114 (I326839,I279143,I279131);
not I_19115 (I326856,I279128);
not I_19116 (I326873,I279125);
nor I_19117 (I326890,I326873,I326839);
nand I_19118 (I326907,I326890,I279128);
not I_19119 (I326796,I326907);
nor I_19120 (I326938,I326873,I326856);
and I_19121 (I326955,I326907,I279128);
nor I_19122 (I326972,I326938,I279128);
nand I_19123 (I326989,I279131,I279137);
not I_19124 (I327006,I326989);
nand I_19125 (I327023,I327006,I326972);
nor I_19126 (I327040,I279146,I279140);
not I_19127 (I327057,I279134);
nor I_19128 (I327074,I327057,I279125);
nor I_19129 (I326793,I327074,I326907);
not I_19130 (I327105,I327074);
or I_19131 (I326808,I327023,I327074);
nor I_19132 (I327136,I327074,I326989);
nand I_19133 (I326805,I326938,I327136);
nor I_19134 (I327167,I327040,I327057);
nand I_19135 (I327184,I327006,I327167);
not I_19136 (I326811,I327184);
nor I_19137 (I326814,I326955,I327184);
or I_19138 (I327229,I327074,I327167);
nor I_19139 (I326799,I327006,I327229);
nor I_19140 (I327260,I327167,I279128);
nand I_19141 (I327277,I327260,I327006);
nand I_19142 (I327294,I327105,I327277);
DFFARX1 I_19143 (I327294,I1862,I326822,I326802,);
not I_19144 (I327349,I1869);
nor I_19145 (I327366,I55816,I55813);
not I_19146 (I327383,I55831);
not I_19147 (I327400,I55822);
nor I_19148 (I327417,I327400,I327366);
nand I_19149 (I327434,I327417,I55831);
not I_19150 (I327323,I327434);
nor I_19151 (I327465,I327400,I327383);
and I_19152 (I327482,I327434,I55837);
nor I_19153 (I327499,I327465,I55837);
nand I_19154 (I327516,I55834,I55825);
not I_19155 (I327533,I327516);
nand I_19156 (I327550,I327533,I327499);
nor I_19157 (I327567,I55813,I55816);
not I_19158 (I327584,I55828);
nor I_19159 (I327601,I327584,I55819);
nor I_19160 (I327320,I327601,I327434);
not I_19161 (I327632,I327601);
or I_19162 (I327335,I327550,I327601);
nor I_19163 (I327663,I327601,I327516);
nand I_19164 (I327332,I327465,I327663);
nor I_19165 (I327694,I327567,I327584);
nand I_19166 (I327711,I327533,I327694);
not I_19167 (I327338,I327711);
nor I_19168 (I327341,I327482,I327711);
or I_19169 (I327756,I327601,I327694);
nor I_19170 (I327326,I327533,I327756);
nor I_19171 (I327787,I327694,I55837);
nand I_19172 (I327804,I327787,I327533);
nand I_19173 (I327821,I327632,I327804);
DFFARX1 I_19174 (I327821,I1862,I327349,I327329,);
not I_19175 (I327876,I1869);
nor I_19176 (I327893,I28276,I28273);
not I_19177 (I327910,I28291);
not I_19178 (I327927,I28282);
nor I_19179 (I327944,I327927,I327893);
nand I_19180 (I327961,I327944,I28291);
not I_19181 (I327850,I327961);
nor I_19182 (I327992,I327927,I327910);
and I_19183 (I328009,I327961,I28297);
nor I_19184 (I328026,I327992,I28297);
nand I_19185 (I328043,I28294,I28285);
not I_19186 (I328060,I328043);
nand I_19187 (I328077,I328060,I328026);
nor I_19188 (I328094,I28273,I28276);
not I_19189 (I328111,I28288);
nor I_19190 (I328128,I328111,I28279);
nor I_19191 (I327847,I328128,I327961);
not I_19192 (I328159,I328128);
or I_19193 (I327862,I328077,I328128);
nor I_19194 (I328190,I328128,I328043);
nand I_19195 (I327859,I327992,I328190);
nor I_19196 (I328221,I328094,I328111);
nand I_19197 (I328238,I328060,I328221);
not I_19198 (I327865,I328238);
nor I_19199 (I327868,I328009,I328238);
or I_19200 (I328283,I328128,I328221);
nor I_19201 (I327853,I328060,I328283);
nor I_19202 (I328314,I328221,I28297);
nand I_19203 (I328331,I328314,I328060);
nand I_19204 (I328348,I328159,I328331);
DFFARX1 I_19205 (I328348,I1862,I327876,I327856,);
not I_19206 (I328403,I1869);
nor I_19207 (I328420,I180559,I180583);
not I_19208 (I328437,I180568);
not I_19209 (I328454,I180562);
nor I_19210 (I328471,I328454,I328420);
nand I_19211 (I328488,I328471,I180568);
not I_19212 (I328377,I328488);
nor I_19213 (I328519,I328454,I328437);
and I_19214 (I328536,I328488,I180565);
nor I_19215 (I328553,I328519,I180565);
nand I_19216 (I328570,I180559,I180574);
not I_19217 (I328587,I328570);
nand I_19218 (I328604,I328587,I328553);
nor I_19219 (I328621,I180571,I180562);
not I_19220 (I328638,I180580);
nor I_19221 (I328655,I328638,I180577);
nor I_19222 (I328374,I328655,I328488);
not I_19223 (I328686,I328655);
or I_19224 (I328389,I328604,I328655);
nor I_19225 (I328717,I328655,I328570);
nand I_19226 (I328386,I328519,I328717);
nor I_19227 (I328748,I328621,I328638);
nand I_19228 (I328765,I328587,I328748);
not I_19229 (I328392,I328765);
nor I_19230 (I328395,I328536,I328765);
or I_19231 (I328810,I328655,I328748);
nor I_19232 (I328380,I328587,I328810);
nor I_19233 (I328841,I328748,I180565);
nand I_19234 (I328858,I328841,I328587);
nand I_19235 (I328875,I328686,I328858);
DFFARX1 I_19236 (I328875,I1862,I328403,I328383,);
not I_19237 (I328930,I1869);
nor I_19238 (I328947,I386684,I386687);
not I_19239 (I328964,I386699);
not I_19240 (I328981,I386690);
nor I_19241 (I328998,I328981,I328947);
nand I_19242 (I329015,I328998,I386699);
not I_19243 (I328904,I329015);
nor I_19244 (I329046,I328981,I328964);
and I_19245 (I329063,I329015,I386693);
nor I_19246 (I329080,I329046,I386693);
nand I_19247 (I329097,I386690,I386696);
not I_19248 (I329114,I329097);
nand I_19249 (I329131,I329114,I329080);
nor I_19250 (I329148,I386687,I386702);
not I_19251 (I329165,I386693);
nor I_19252 (I329182,I329165,I386684);
nor I_19253 (I328901,I329182,I329015);
not I_19254 (I329213,I329182);
or I_19255 (I328916,I329131,I329182);
nor I_19256 (I329244,I329182,I329097);
nand I_19257 (I328913,I329046,I329244);
nor I_19258 (I329275,I329148,I329165);
nand I_19259 (I329292,I329114,I329275);
not I_19260 (I328919,I329292);
nor I_19261 (I328922,I329063,I329292);
or I_19262 (I329337,I329182,I329275);
nor I_19263 (I328907,I329114,I329337);
nor I_19264 (I329368,I329275,I386693);
nand I_19265 (I329385,I329368,I329114);
nand I_19266 (I329402,I329213,I329385);
DFFARX1 I_19267 (I329402,I1862,I328930,I328910,);
not I_19268 (I329457,I1869);
nor I_19269 (I329474,I115282,I115297);
not I_19270 (I329491,I115285);
not I_19271 (I329508,I115279);
nor I_19272 (I329525,I329508,I329474);
nand I_19273 (I329542,I329525,I115285);
not I_19274 (I329431,I329542);
nor I_19275 (I329573,I329508,I329491);
and I_19276 (I329590,I329542,I115294);
nor I_19277 (I329607,I329573,I115294);
nand I_19278 (I329624,I115279,I115288);
not I_19279 (I329641,I329624);
nand I_19280 (I329658,I329641,I329607);
nor I_19281 (I329675,I115291,I115282);
not I_19282 (I329692,I115285);
nor I_19283 (I329709,I329692,I115288);
nor I_19284 (I329428,I329709,I329542);
not I_19285 (I329740,I329709);
or I_19286 (I329443,I329658,I329709);
nor I_19287 (I329771,I329709,I329624);
nand I_19288 (I329440,I329573,I329771);
nor I_19289 (I329802,I329675,I329692);
nand I_19290 (I329819,I329641,I329802);
not I_19291 (I329446,I329819);
nor I_19292 (I329449,I329590,I329819);
or I_19293 (I329864,I329709,I329802);
nor I_19294 (I329434,I329641,I329864);
nor I_19295 (I329895,I329802,I115294);
nand I_19296 (I329912,I329895,I329641);
nand I_19297 (I329929,I329740,I329912);
DFFARX1 I_19298 (I329929,I1862,I329457,I329437,);
not I_19299 (I329984,I1869);
nor I_19300 (I330001,I284855,I284843);
not I_19301 (I330018,I284840);
not I_19302 (I330035,I284837);
nor I_19303 (I330052,I330035,I330001);
nand I_19304 (I330069,I330052,I284840);
not I_19305 (I329958,I330069);
nor I_19306 (I330100,I330035,I330018);
and I_19307 (I330117,I330069,I284840);
nor I_19308 (I330134,I330100,I284840);
nand I_19309 (I330151,I284843,I284849);
not I_19310 (I330168,I330151);
nand I_19311 (I330185,I330168,I330134);
nor I_19312 (I330202,I284858,I284852);
not I_19313 (I330219,I284846);
nor I_19314 (I330236,I330219,I284837);
nor I_19315 (I329955,I330236,I330069);
not I_19316 (I330267,I330236);
or I_19317 (I329970,I330185,I330236);
nor I_19318 (I330298,I330236,I330151);
nand I_19319 (I329967,I330100,I330298);
nor I_19320 (I330329,I330202,I330219);
nand I_19321 (I330346,I330168,I330329);
not I_19322 (I329973,I330346);
nor I_19323 (I329976,I330117,I330346);
or I_19324 (I330391,I330236,I330329);
nor I_19325 (I329961,I330168,I330391);
nor I_19326 (I330422,I330329,I284840);
nand I_19327 (I330439,I330422,I330168);
nand I_19328 (I330456,I330267,I330439);
DFFARX1 I_19329 (I330456,I1862,I329984,I329964,);
not I_19330 (I330511,I1869);
nor I_19331 (I330528,I13996,I13993);
not I_19332 (I330545,I14011);
not I_19333 (I330562,I14002);
nor I_19334 (I330579,I330562,I330528);
nand I_19335 (I330596,I330579,I14011);
not I_19336 (I330485,I330596);
nor I_19337 (I330627,I330562,I330545);
and I_19338 (I330644,I330596,I14017);
nor I_19339 (I330661,I330627,I14017);
nand I_19340 (I330678,I14014,I14005);
not I_19341 (I330695,I330678);
nand I_19342 (I330712,I330695,I330661);
nor I_19343 (I330729,I13993,I13996);
not I_19344 (I330746,I14008);
nor I_19345 (I330763,I330746,I13999);
nor I_19346 (I330482,I330763,I330596);
not I_19347 (I330794,I330763);
or I_19348 (I330497,I330712,I330763);
nor I_19349 (I330825,I330763,I330678);
nand I_19350 (I330494,I330627,I330825);
nor I_19351 (I330856,I330729,I330746);
nand I_19352 (I330873,I330695,I330856);
not I_19353 (I330500,I330873);
nor I_19354 (I330503,I330644,I330873);
or I_19355 (I330918,I330763,I330856);
nor I_19356 (I330488,I330695,I330918);
nor I_19357 (I330949,I330856,I14017);
nand I_19358 (I330966,I330949,I330695);
nand I_19359 (I330983,I330794,I330966);
DFFARX1 I_19360 (I330983,I1862,I330511,I330491,);
not I_19361 (I331038,I1869);
nor I_19362 (I331055,I91006,I91003);
not I_19363 (I331072,I91021);
not I_19364 (I331089,I91012);
nor I_19365 (I331106,I331089,I331055);
nand I_19366 (I331123,I331106,I91021);
not I_19367 (I331012,I331123);
nor I_19368 (I331154,I331089,I331072);
and I_19369 (I331171,I331123,I91027);
nor I_19370 (I331188,I331154,I91027);
nand I_19371 (I331205,I91024,I91015);
not I_19372 (I331222,I331205);
nand I_19373 (I331239,I331222,I331188);
nor I_19374 (I331256,I91003,I91006);
not I_19375 (I331273,I91018);
nor I_19376 (I331290,I331273,I91009);
nor I_19377 (I331009,I331290,I331123);
not I_19378 (I331321,I331290);
or I_19379 (I331024,I331239,I331290);
nor I_19380 (I331352,I331290,I331205);
nand I_19381 (I331021,I331154,I331352);
nor I_19382 (I331383,I331256,I331273);
nand I_19383 (I331400,I331222,I331383);
not I_19384 (I331027,I331400);
nor I_19385 (I331030,I331171,I331400);
or I_19386 (I331445,I331290,I331383);
nor I_19387 (I331015,I331222,I331445);
nor I_19388 (I331476,I331383,I91027);
nand I_19389 (I331493,I331476,I331222);
nand I_19390 (I331510,I331321,I331493);
DFFARX1 I_19391 (I331510,I1862,I331038,I331018,);
not I_19392 (I331565,I1869);
nor I_19393 (I331582,I273907,I273895);
not I_19394 (I331599,I273892);
not I_19395 (I331616,I273889);
nor I_19396 (I331633,I331616,I331582);
nand I_19397 (I331650,I331633,I273892);
not I_19398 (I331539,I331650);
nor I_19399 (I331681,I331616,I331599);
and I_19400 (I331698,I331650,I273892);
nor I_19401 (I331715,I331681,I273892);
nand I_19402 (I331732,I273895,I273901);
not I_19403 (I331749,I331732);
nand I_19404 (I331766,I331749,I331715);
nor I_19405 (I331783,I273910,I273904);
not I_19406 (I331800,I273898);
nor I_19407 (I331817,I331800,I273889);
nor I_19408 (I331536,I331817,I331650);
not I_19409 (I331848,I331817);
or I_19410 (I331551,I331766,I331817);
nor I_19411 (I331879,I331817,I331732);
nand I_19412 (I331548,I331681,I331879);
nor I_19413 (I331910,I331783,I331800);
nand I_19414 (I331927,I331749,I331910);
not I_19415 (I331554,I331927);
nor I_19416 (I331557,I331698,I331927);
or I_19417 (I331972,I331817,I331910);
nor I_19418 (I331542,I331749,I331972);
nor I_19419 (I332003,I331910,I273892);
nand I_19420 (I332020,I332003,I331749);
nand I_19421 (I332037,I331848,I332020);
DFFARX1 I_19422 (I332037,I1862,I331565,I331545,);
not I_19423 (I332092,I1869);
nor I_19424 (I332109,I218691,I218679);
not I_19425 (I332126,I218676);
not I_19426 (I332143,I218673);
nor I_19427 (I332160,I332143,I332109);
nand I_19428 (I332177,I332160,I218676);
not I_19429 (I332066,I332177);
nor I_19430 (I332208,I332143,I332126);
and I_19431 (I332225,I332177,I218676);
nor I_19432 (I332242,I332208,I218676);
nand I_19433 (I332259,I218679,I218685);
not I_19434 (I332276,I332259);
nand I_19435 (I332293,I332276,I332242);
nor I_19436 (I332310,I218694,I218688);
not I_19437 (I332327,I218682);
nor I_19438 (I332344,I332327,I218673);
nor I_19439 (I332063,I332344,I332177);
not I_19440 (I332375,I332344);
or I_19441 (I332078,I332293,I332344);
nor I_19442 (I332406,I332344,I332259);
nand I_19443 (I332075,I332208,I332406);
nor I_19444 (I332437,I332310,I332327);
nand I_19445 (I332454,I332276,I332437);
not I_19446 (I332081,I332454);
nor I_19447 (I332084,I332225,I332454);
or I_19448 (I332499,I332344,I332437);
nor I_19449 (I332069,I332276,I332499);
nor I_19450 (I332530,I332437,I218676);
nand I_19451 (I332547,I332530,I332276);
nand I_19452 (I332564,I332375,I332547);
DFFARX1 I_19453 (I332564,I1862,I332092,I332072,);
not I_19454 (I332619,I1869);
nor I_19455 (I332636,I75706,I75703);
not I_19456 (I332653,I75721);
not I_19457 (I332670,I75712);
nor I_19458 (I332687,I332670,I332636);
nand I_19459 (I332704,I332687,I75721);
not I_19460 (I332593,I332704);
nor I_19461 (I332735,I332670,I332653);
and I_19462 (I332752,I332704,I75727);
nor I_19463 (I332769,I332735,I75727);
nand I_19464 (I332786,I75724,I75715);
not I_19465 (I332803,I332786);
nand I_19466 (I332820,I332803,I332769);
nor I_19467 (I332837,I75703,I75706);
not I_19468 (I332854,I75718);
nor I_19469 (I332871,I332854,I75709);
nor I_19470 (I332590,I332871,I332704);
not I_19471 (I332902,I332871);
or I_19472 (I332605,I332820,I332871);
nor I_19473 (I332933,I332871,I332786);
nand I_19474 (I332602,I332735,I332933);
nor I_19475 (I332964,I332837,I332854);
nand I_19476 (I332981,I332803,I332964);
not I_19477 (I332608,I332981);
nor I_19478 (I332611,I332752,I332981);
or I_19479 (I333026,I332871,I332964);
nor I_19480 (I332596,I332803,I333026);
nor I_19481 (I333057,I332964,I75727);
nand I_19482 (I333074,I333057,I332803);
nand I_19483 (I333091,I332902,I333074);
DFFARX1 I_19484 (I333091,I1862,I332619,I332599,);
not I_19485 (I333146,I1869);
nor I_19486 (I333163,I55306,I55303);
not I_19487 (I333180,I55321);
not I_19488 (I333197,I55312);
nor I_19489 (I333214,I333197,I333163);
nand I_19490 (I333231,I333214,I55321);
not I_19491 (I333120,I333231);
nor I_19492 (I333262,I333197,I333180);
and I_19493 (I333279,I333231,I55327);
nor I_19494 (I333296,I333262,I55327);
nand I_19495 (I333313,I55324,I55315);
not I_19496 (I333330,I333313);
nand I_19497 (I333347,I333330,I333296);
nor I_19498 (I333364,I55303,I55306);
not I_19499 (I333381,I55318);
nor I_19500 (I333398,I333381,I55309);
nor I_19501 (I333117,I333398,I333231);
not I_19502 (I333429,I333398);
or I_19503 (I333132,I333347,I333398);
nor I_19504 (I333460,I333398,I333313);
nand I_19505 (I333129,I333262,I333460);
nor I_19506 (I333491,I333364,I333381);
nand I_19507 (I333508,I333330,I333491);
not I_19508 (I333135,I333508);
nor I_19509 (I333138,I333279,I333508);
or I_19510 (I333553,I333398,I333491);
nor I_19511 (I333123,I333330,I333553);
nor I_19512 (I333584,I333491,I55327);
nand I_19513 (I333601,I333584,I333330);
nand I_19514 (I333618,I333429,I333601);
DFFARX1 I_19515 (I333618,I1862,I333146,I333126,);
not I_19516 (I333673,I1869);
nor I_19517 (I333690,I163695,I163719);
not I_19518 (I333707,I163704);
not I_19519 (I333724,I163698);
nor I_19520 (I333741,I333724,I333690);
nand I_19521 (I333758,I333741,I163704);
not I_19522 (I333647,I333758);
nor I_19523 (I333789,I333724,I333707);
and I_19524 (I333806,I333758,I163701);
nor I_19525 (I333823,I333789,I163701);
nand I_19526 (I333840,I163695,I163710);
not I_19527 (I333857,I333840);
nand I_19528 (I333874,I333857,I333823);
nor I_19529 (I333891,I163707,I163698);
not I_19530 (I333908,I163716);
nor I_19531 (I333925,I333908,I163713);
nor I_19532 (I333644,I333925,I333758);
not I_19533 (I333956,I333925);
or I_19534 (I333659,I333874,I333925);
nor I_19535 (I333987,I333925,I333840);
nand I_19536 (I333656,I333789,I333987);
nor I_19537 (I334018,I333891,I333908);
nand I_19538 (I334035,I333857,I334018);
not I_19539 (I333662,I334035);
nor I_19540 (I333665,I333806,I334035);
or I_19541 (I334080,I333925,I334018);
nor I_19542 (I333650,I333857,I334080);
nor I_19543 (I334111,I334018,I163701);
nand I_19544 (I334128,I334111,I333857);
nand I_19545 (I334145,I333956,I334128);
DFFARX1 I_19546 (I334145,I1862,I333673,I333653,);
not I_19547 (I334200,I1869);
nor I_19548 (I334217,I33376,I33373);
not I_19549 (I334234,I33391);
not I_19550 (I334251,I33382);
nor I_19551 (I334268,I334251,I334217);
nand I_19552 (I334285,I334268,I33391);
not I_19553 (I334174,I334285);
nor I_19554 (I334316,I334251,I334234);
and I_19555 (I334333,I334285,I33397);
nor I_19556 (I334350,I334316,I33397);
nand I_19557 (I334367,I33394,I33385);
not I_19558 (I334384,I334367);
nand I_19559 (I334401,I334384,I334350);
nor I_19560 (I334418,I33373,I33376);
not I_19561 (I334435,I33388);
nor I_19562 (I334452,I334435,I33379);
nor I_19563 (I334171,I334452,I334285);
not I_19564 (I334483,I334452);
or I_19565 (I334186,I334401,I334452);
nor I_19566 (I334514,I334452,I334367);
nand I_19567 (I334183,I334316,I334514);
nor I_19568 (I334545,I334418,I334435);
nand I_19569 (I334562,I334384,I334545);
not I_19570 (I334189,I334562);
nor I_19571 (I334192,I334333,I334562);
or I_19572 (I334607,I334452,I334545);
nor I_19573 (I334177,I334384,I334607);
nor I_19574 (I334638,I334545,I33397);
nand I_19575 (I334655,I334638,I334384);
nand I_19576 (I334672,I334483,I334655);
DFFARX1 I_19577 (I334672,I1862,I334200,I334180,);
not I_19578 (I334727,I1869);
nor I_19579 (I334744,I69076,I69073);
not I_19580 (I334761,I69091);
not I_19581 (I334778,I69082);
nor I_19582 (I334795,I334778,I334744);
nand I_19583 (I334812,I334795,I69091);
not I_19584 (I334701,I334812);
nor I_19585 (I334843,I334778,I334761);
and I_19586 (I334860,I334812,I69097);
nor I_19587 (I334877,I334843,I69097);
nand I_19588 (I334894,I69094,I69085);
not I_19589 (I334911,I334894);
nand I_19590 (I334928,I334911,I334877);
nor I_19591 (I334945,I69073,I69076);
not I_19592 (I334962,I69088);
nor I_19593 (I334979,I334962,I69079);
nor I_19594 (I334698,I334979,I334812);
not I_19595 (I335010,I334979);
or I_19596 (I334713,I334928,I334979);
nor I_19597 (I335041,I334979,I334894);
nand I_19598 (I334710,I334843,I335041);
nor I_19599 (I335072,I334945,I334962);
nand I_19600 (I335089,I334911,I335072);
not I_19601 (I334716,I335089);
nor I_19602 (I334719,I334860,I335089);
or I_19603 (I335134,I334979,I335072);
nor I_19604 (I334704,I334911,I335134);
nor I_19605 (I335165,I335072,I69097);
nand I_19606 (I335182,I335165,I334911);
nand I_19607 (I335199,I335010,I335182);
DFFARX1 I_19608 (I335199,I1862,I334727,I334707,);
not I_19609 (I335254,I1869);
nor I_19610 (I335271,I73666,I73663);
not I_19611 (I335288,I73681);
not I_19612 (I335305,I73672);
nor I_19613 (I335322,I335305,I335271);
nand I_19614 (I335339,I335322,I73681);
not I_19615 (I335228,I335339);
nor I_19616 (I335370,I335305,I335288);
and I_19617 (I335387,I335339,I73687);
nor I_19618 (I335404,I335370,I73687);
nand I_19619 (I335421,I73684,I73675);
not I_19620 (I335438,I335421);
nand I_19621 (I335455,I335438,I335404);
nor I_19622 (I335472,I73663,I73666);
not I_19623 (I335489,I73678);
nor I_19624 (I335506,I335489,I73669);
nor I_19625 (I335225,I335506,I335339);
not I_19626 (I335537,I335506);
or I_19627 (I335240,I335455,I335506);
nor I_19628 (I335568,I335506,I335421);
nand I_19629 (I335237,I335370,I335568);
nor I_19630 (I335599,I335472,I335489);
nand I_19631 (I335616,I335438,I335599);
not I_19632 (I335243,I335616);
nor I_19633 (I335246,I335387,I335616);
or I_19634 (I335661,I335506,I335599);
nor I_19635 (I335231,I335438,I335661);
nor I_19636 (I335692,I335599,I73687);
nand I_19637 (I335709,I335692,I335438);
nand I_19638 (I335726,I335537,I335709);
DFFARX1 I_19639 (I335726,I1862,I335254,I335234,);
not I_19640 (I335781,I1869);
nor I_19641 (I335798,I229639,I229627);
not I_19642 (I335815,I229624);
not I_19643 (I335832,I229621);
nor I_19644 (I335849,I335832,I335798);
nand I_19645 (I335866,I335849,I229624);
not I_19646 (I335755,I335866);
nor I_19647 (I335897,I335832,I335815);
and I_19648 (I335914,I335866,I229624);
nor I_19649 (I335931,I335897,I229624);
nand I_19650 (I335948,I229627,I229633);
not I_19651 (I335965,I335948);
nand I_19652 (I335982,I335965,I335931);
nor I_19653 (I335999,I229642,I229636);
not I_19654 (I336016,I229630);
nor I_19655 (I336033,I336016,I229621);
nor I_19656 (I335752,I336033,I335866);
not I_19657 (I336064,I336033);
or I_19658 (I335767,I335982,I336033);
nor I_19659 (I336095,I336033,I335948);
nand I_19660 (I335764,I335897,I336095);
nor I_19661 (I336126,I335999,I336016);
nand I_19662 (I336143,I335965,I336126);
not I_19663 (I335770,I336143);
nor I_19664 (I335773,I335914,I336143);
or I_19665 (I336188,I336033,I336126);
nor I_19666 (I335758,I335965,I336188);
nor I_19667 (I336219,I336126,I229624);
nand I_19668 (I336236,I336219,I335965);
nand I_19669 (I336253,I336064,I336236);
DFFARX1 I_19670 (I336253,I1862,I335781,I335761,);
not I_19671 (I336308,I1869);
nor I_19672 (I336325,I33886,I33883);
not I_19673 (I336342,I33901);
not I_19674 (I336359,I33892);
nor I_19675 (I336376,I336359,I336325);
nand I_19676 (I336393,I336376,I33901);
not I_19677 (I336282,I336393);
nor I_19678 (I336424,I336359,I336342);
and I_19679 (I336441,I336393,I33907);
nor I_19680 (I336458,I336424,I33907);
nand I_19681 (I336475,I33904,I33895);
not I_19682 (I336492,I336475);
nand I_19683 (I336509,I336492,I336458);
nor I_19684 (I336526,I33883,I33886);
not I_19685 (I336543,I33898);
nor I_19686 (I336560,I336543,I33889);
nor I_19687 (I336279,I336560,I336393);
not I_19688 (I336591,I336560);
or I_19689 (I336294,I336509,I336560);
nor I_19690 (I336622,I336560,I336475);
nand I_19691 (I336291,I336424,I336622);
nor I_19692 (I336653,I336526,I336543);
nand I_19693 (I336670,I336492,I336653);
not I_19694 (I336297,I336670);
nor I_19695 (I336300,I336441,I336670);
or I_19696 (I336715,I336560,I336653);
nor I_19697 (I336285,I336492,I336715);
nor I_19698 (I336746,I336653,I33907);
nand I_19699 (I336763,I336746,I336492);
nand I_19700 (I336780,I336591,I336763);
DFFARX1 I_19701 (I336780,I1862,I336308,I336288,);
not I_19702 (I336835,I1869);
nor I_19703 (I336852,I66526,I66523);
not I_19704 (I336869,I66541);
not I_19705 (I336886,I66532);
nor I_19706 (I336903,I336886,I336852);
nand I_19707 (I336920,I336903,I66541);
not I_19708 (I336809,I336920);
nor I_19709 (I336951,I336886,I336869);
and I_19710 (I336968,I336920,I66547);
nor I_19711 (I336985,I336951,I66547);
nand I_19712 (I337002,I66544,I66535);
not I_19713 (I337019,I337002);
nand I_19714 (I337036,I337019,I336985);
nor I_19715 (I337053,I66523,I66526);
not I_19716 (I337070,I66538);
nor I_19717 (I337087,I337070,I66529);
nor I_19718 (I336806,I337087,I336920);
not I_19719 (I337118,I337087);
or I_19720 (I336821,I337036,I337087);
nor I_19721 (I337149,I337087,I337002);
nand I_19722 (I336818,I336951,I337149);
nor I_19723 (I337180,I337053,I337070);
nand I_19724 (I337197,I337019,I337180);
not I_19725 (I336824,I337197);
nor I_19726 (I336827,I336968,I337197);
or I_19727 (I337242,I337087,I337180);
nor I_19728 (I336812,I337019,I337242);
nor I_19729 (I337273,I337180,I66547);
nand I_19730 (I337290,I337273,I337019);
nand I_19731 (I337307,I337118,I337290);
DFFARX1 I_19732 (I337307,I1862,I336835,I336815,);
not I_19733 (I337362,I1869);
nor I_19734 (I337379,I189518,I189542);
not I_19735 (I337396,I189527);
not I_19736 (I337413,I189521);
nor I_19737 (I337430,I337413,I337379);
nand I_19738 (I337447,I337430,I189527);
not I_19739 (I337336,I337447);
nor I_19740 (I337478,I337413,I337396);
and I_19741 (I337495,I337447,I189524);
nor I_19742 (I337512,I337478,I189524);
nand I_19743 (I337529,I189518,I189533);
not I_19744 (I337546,I337529);
nand I_19745 (I337563,I337546,I337512);
nor I_19746 (I337580,I189530,I189521);
not I_19747 (I337597,I189539);
nor I_19748 (I337614,I337597,I189536);
nor I_19749 (I337333,I337614,I337447);
not I_19750 (I337645,I337614);
or I_19751 (I337348,I337563,I337614);
nor I_19752 (I337676,I337614,I337529);
nand I_19753 (I337345,I337478,I337676);
nor I_19754 (I337707,I337580,I337597);
nand I_19755 (I337724,I337546,I337707);
not I_19756 (I337351,I337724);
nor I_19757 (I337354,I337495,I337724);
or I_19758 (I337769,I337614,I337707);
nor I_19759 (I337339,I337546,I337769);
nor I_19760 (I337800,I337707,I189524);
nand I_19761 (I337817,I337800,I337546);
nand I_19762 (I337834,I337645,I337817);
DFFARX1 I_19763 (I337834,I1862,I337362,I337342,);
not I_19764 (I337889,I1869);
nor I_19765 (I337906,I200058,I200082);
not I_19766 (I337923,I200067);
not I_19767 (I337940,I200061);
nor I_19768 (I337957,I337940,I337906);
nand I_19769 (I337974,I337957,I200067);
not I_19770 (I337863,I337974);
nor I_19771 (I338005,I337940,I337923);
and I_19772 (I338022,I337974,I200064);
nor I_19773 (I338039,I338005,I200064);
nand I_19774 (I338056,I200058,I200073);
not I_19775 (I338073,I338056);
nand I_19776 (I338090,I338073,I338039);
nor I_19777 (I338107,I200070,I200061);
not I_19778 (I338124,I200079);
nor I_19779 (I338141,I338124,I200076);
nor I_19780 (I337860,I338141,I337974);
not I_19781 (I338172,I338141);
or I_19782 (I337875,I338090,I338141);
nor I_19783 (I338203,I338141,I338056);
nand I_19784 (I337872,I338005,I338203);
nor I_19785 (I338234,I338107,I338124);
nand I_19786 (I338251,I338073,I338234);
not I_19787 (I337878,I338251);
nor I_19788 (I337881,I338022,I338251);
or I_19789 (I338296,I338141,I338234);
nor I_19790 (I337866,I338073,I338296);
nor I_19791 (I338327,I338234,I200064);
nand I_19792 (I338344,I338327,I338073);
nand I_19793 (I338361,I338172,I338344);
DFFARX1 I_19794 (I338361,I1862,I337889,I337869,);
not I_19795 (I338416,I1869);
nor I_19796 (I338433,I149993,I150017);
not I_19797 (I338450,I150002);
not I_19798 (I338467,I149996);
nor I_19799 (I338484,I338467,I338433);
nand I_19800 (I338501,I338484,I150002);
not I_19801 (I338390,I338501);
nor I_19802 (I338532,I338467,I338450);
and I_19803 (I338549,I338501,I149999);
nor I_19804 (I338566,I338532,I149999);
nand I_19805 (I338583,I149993,I150008);
not I_19806 (I338600,I338583);
nand I_19807 (I338617,I338600,I338566);
nor I_19808 (I338634,I150005,I149996);
not I_19809 (I338651,I150014);
nor I_19810 (I338668,I338651,I150011);
nor I_19811 (I338387,I338668,I338501);
not I_19812 (I338699,I338668);
or I_19813 (I338402,I338617,I338668);
nor I_19814 (I338730,I338668,I338583);
nand I_19815 (I338399,I338532,I338730);
nor I_19816 (I338761,I338634,I338651);
nand I_19817 (I338778,I338600,I338761);
not I_19818 (I338405,I338778);
nor I_19819 (I338408,I338549,I338778);
or I_19820 (I338823,I338668,I338761);
nor I_19821 (I338393,I338600,I338823);
nor I_19822 (I338854,I338761,I149999);
nand I_19823 (I338871,I338854,I338600);
nand I_19824 (I338888,I338699,I338871);
DFFARX1 I_19825 (I338888,I1862,I338416,I338396,);
not I_19826 (I338943,I1869);
nor I_19827 (I338960,I264387,I264375);
not I_19828 (I338977,I264372);
not I_19829 (I338994,I264369);
nor I_19830 (I339011,I338994,I338960);
nand I_19831 (I339028,I339011,I264372);
not I_19832 (I338917,I339028);
nor I_19833 (I339059,I338994,I338977);
and I_19834 (I339076,I339028,I264372);
nor I_19835 (I339093,I339059,I264372);
nand I_19836 (I339110,I264375,I264381);
not I_19837 (I339127,I339110);
nand I_19838 (I339144,I339127,I339093);
nor I_19839 (I339161,I264390,I264384);
not I_19840 (I339178,I264378);
nor I_19841 (I339195,I339178,I264369);
nor I_19842 (I338914,I339195,I339028);
not I_19843 (I339226,I339195);
or I_19844 (I338929,I339144,I339195);
nor I_19845 (I339257,I339195,I339110);
nand I_19846 (I338926,I339059,I339257);
nor I_19847 (I339288,I339161,I339178);
nand I_19848 (I339305,I339127,I339288);
not I_19849 (I338932,I339305);
nor I_19850 (I338935,I339076,I339305);
or I_19851 (I339350,I339195,I339288);
nor I_19852 (I338920,I339127,I339350);
nor I_19853 (I339381,I339288,I264372);
nand I_19854 (I339398,I339381,I339127);
nand I_19855 (I339415,I339226,I339398);
DFFARX1 I_19856 (I339415,I1862,I338943,I338923,);
not I_19857 (I339470,I1869);
nor I_19858 (I339487,I395524,I395527);
not I_19859 (I339504,I395539);
not I_19860 (I339521,I395530);
nor I_19861 (I339538,I339521,I339487);
nand I_19862 (I339555,I339538,I395539);
not I_19863 (I339444,I339555);
nor I_19864 (I339586,I339521,I339504);
and I_19865 (I339603,I339555,I395533);
nor I_19866 (I339620,I339586,I395533);
nand I_19867 (I339637,I395530,I395536);
not I_19868 (I339654,I339637);
nand I_19869 (I339671,I339654,I339620);
nor I_19870 (I339688,I395527,I395542);
not I_19871 (I339705,I395533);
nor I_19872 (I339722,I339705,I395524);
nor I_19873 (I339441,I339722,I339555);
not I_19874 (I339753,I339722);
or I_19875 (I339456,I339671,I339722);
nor I_19876 (I339784,I339722,I339637);
nand I_19877 (I339453,I339586,I339784);
nor I_19878 (I339815,I339688,I339705);
nand I_19879 (I339832,I339654,I339815);
not I_19880 (I339459,I339832);
nor I_19881 (I339462,I339603,I339832);
or I_19882 (I339877,I339722,I339815);
nor I_19883 (I339447,I339654,I339877);
nor I_19884 (I339908,I339815,I395533);
nand I_19885 (I339925,I339908,I339654);
nand I_19886 (I339942,I339753,I339925);
DFFARX1 I_19887 (I339942,I1862,I339470,I339450,);
not I_19888 (I339997,I1869);
nor I_19889 (I340014,I158952,I158976);
not I_19890 (I340031,I158961);
not I_19891 (I340048,I158955);
nor I_19892 (I340065,I340048,I340014);
nand I_19893 (I340082,I340065,I158961);
not I_19894 (I339971,I340082);
nor I_19895 (I340113,I340048,I340031);
and I_19896 (I340130,I340082,I158958);
nor I_19897 (I340147,I340113,I158958);
nand I_19898 (I340164,I158952,I158967);
not I_19899 (I340181,I340164);
nand I_19900 (I340198,I340181,I340147);
nor I_19901 (I340215,I158964,I158955);
not I_19902 (I340232,I158973);
nor I_19903 (I340249,I340232,I158970);
nor I_19904 (I339968,I340249,I340082);
not I_19905 (I340280,I340249);
or I_19906 (I339983,I340198,I340249);
nor I_19907 (I340311,I340249,I340164);
nand I_19908 (I339980,I340113,I340311);
nor I_19909 (I340342,I340215,I340232);
nand I_19910 (I340359,I340181,I340342);
not I_19911 (I339986,I340359);
nor I_19912 (I339989,I340130,I340359);
or I_19913 (I340404,I340249,I340342);
nor I_19914 (I339974,I340181,I340404);
nor I_19915 (I340435,I340342,I158958);
nand I_19916 (I340452,I340435,I340181);
nand I_19917 (I340469,I340280,I340452);
DFFARX1 I_19918 (I340469,I1862,I339997,I339977,);
not I_19919 (I340524,I1869);
nor I_19920 (I340541,I295703,I295700);
not I_19921 (I340558,I295709);
not I_19922 (I340575,I295706);
nor I_19923 (I340592,I340575,I340541);
nand I_19924 (I340609,I340592,I295709);
not I_19925 (I340498,I340609);
nor I_19926 (I340640,I340575,I340558);
and I_19927 (I340657,I340609,I295712);
nor I_19928 (I340674,I340640,I295712);
nand I_19929 (I340691,I295715,I295706);
not I_19930 (I340708,I340691);
nand I_19931 (I340725,I340708,I340674);
nor I_19932 (I340742,I295721,I295718);
not I_19933 (I340759,I295700);
nor I_19934 (I340776,I340759,I295703);
nor I_19935 (I340495,I340776,I340609);
not I_19936 (I340807,I340776);
or I_19937 (I340510,I340725,I340776);
nor I_19938 (I340838,I340776,I340691);
nand I_19939 (I340507,I340640,I340838);
nor I_19940 (I340869,I340742,I340759);
nand I_19941 (I340886,I340708,I340869);
not I_19942 (I340513,I340886);
nor I_19943 (I340516,I340657,I340886);
or I_19944 (I340931,I340776,I340869);
nor I_19945 (I340501,I340708,I340931);
nor I_19946 (I340962,I340869,I295712);
nand I_19947 (I340979,I340962,I340708);
nand I_19948 (I340996,I340807,I340979);
DFFARX1 I_19949 (I340996,I1862,I340524,I340504,);
not I_19950 (I341051,I1869);
nor I_19951 (I341068,I405248,I405251);
not I_19952 (I341085,I405263);
not I_19953 (I341102,I405254);
nor I_19954 (I341119,I341102,I341068);
nand I_19955 (I341136,I341119,I405263);
not I_19956 (I341025,I341136);
nor I_19957 (I341167,I341102,I341085);
and I_19958 (I341184,I341136,I405257);
nor I_19959 (I341201,I341167,I405257);
nand I_19960 (I341218,I405254,I405260);
not I_19961 (I341235,I341218);
nand I_19962 (I341252,I341235,I341201);
nor I_19963 (I341269,I405251,I405266);
not I_19964 (I341286,I405257);
nor I_19965 (I341303,I341286,I405248);
nor I_19966 (I341022,I341303,I341136);
not I_19967 (I341334,I341303);
or I_19968 (I341037,I341252,I341303);
nor I_19969 (I341365,I341303,I341218);
nand I_19970 (I341034,I341167,I341365);
nor I_19971 (I341396,I341269,I341286);
nand I_19972 (I341413,I341235,I341396);
not I_19973 (I341040,I341413);
nor I_19974 (I341043,I341184,I341413);
or I_19975 (I341458,I341303,I341396);
nor I_19976 (I341028,I341235,I341458);
nor I_19977 (I341489,I341396,I405257);
nand I_19978 (I341506,I341489,I341235);
nand I_19979 (I341523,I341334,I341506);
DFFARX1 I_19980 (I341523,I1862,I341051,I341031,);
not I_19981 (I341578,I1869);
nor I_19982 (I341595,I172654,I172678);
not I_19983 (I341612,I172663);
not I_19984 (I341629,I172657);
nor I_19985 (I341646,I341629,I341595);
nand I_19986 (I341663,I341646,I172663);
not I_19987 (I341552,I341663);
nor I_19988 (I341694,I341629,I341612);
and I_19989 (I341711,I341663,I172660);
nor I_19990 (I341728,I341694,I172660);
nand I_19991 (I341745,I172654,I172669);
not I_19992 (I341762,I341745);
nand I_19993 (I341779,I341762,I341728);
nor I_19994 (I341796,I172666,I172657);
not I_19995 (I341813,I172675);
nor I_19996 (I341830,I341813,I172672);
nor I_19997 (I341549,I341830,I341663);
not I_19998 (I341861,I341830);
or I_19999 (I341564,I341779,I341830);
nor I_20000 (I341892,I341830,I341745);
nand I_20001 (I341561,I341694,I341892);
nor I_20002 (I341923,I341796,I341813);
nand I_20003 (I341940,I341762,I341923);
not I_20004 (I341567,I341940);
nor I_20005 (I341570,I341711,I341940);
or I_20006 (I341985,I341830,I341923);
nor I_20007 (I341555,I341762,I341985);
nor I_20008 (I342016,I341923,I172660);
nand I_20009 (I342033,I342016,I341762);
nand I_20010 (I342050,I341861,I342033);
DFFARX1 I_20011 (I342050,I1862,I341578,I341558,);
not I_20012 (I342105,I1869);
nor I_20013 (I342122,I206315,I206303);
not I_20014 (I342139,I206300);
not I_20015 (I342156,I206297);
nor I_20016 (I342173,I342156,I342122);
nand I_20017 (I342190,I342173,I206300);
not I_20018 (I342079,I342190);
nor I_20019 (I342221,I342156,I342139);
and I_20020 (I342238,I342190,I206300);
nor I_20021 (I342255,I342221,I206300);
nand I_20022 (I342272,I206303,I206309);
not I_20023 (I342289,I342272);
nand I_20024 (I342306,I342289,I342255);
nor I_20025 (I342323,I206318,I206312);
not I_20026 (I342340,I206306);
nor I_20027 (I342357,I342340,I206297);
nor I_20028 (I342076,I342357,I342190);
not I_20029 (I342388,I342357);
or I_20030 (I342091,I342306,I342357);
nor I_20031 (I342419,I342357,I342272);
nand I_20032 (I342088,I342221,I342419);
nor I_20033 (I342450,I342323,I342340);
nand I_20034 (I342467,I342289,I342450);
not I_20035 (I342094,I342467);
nor I_20036 (I342097,I342238,I342467);
or I_20037 (I342512,I342357,I342450);
nor I_20038 (I342082,I342289,I342512);
nor I_20039 (I342543,I342450,I206300);
nand I_20040 (I342560,I342543,I342289);
nand I_20041 (I342577,I342388,I342560);
DFFARX1 I_20042 (I342577,I1862,I342105,I342085,);
not I_20043 (I342632,I1869);
nor I_20044 (I342649,I202031,I202019);
not I_20045 (I342666,I202016);
not I_20046 (I342683,I202013);
nor I_20047 (I342700,I342683,I342649);
nand I_20048 (I342717,I342700,I202016);
not I_20049 (I342606,I342717);
nor I_20050 (I342748,I342683,I342666);
and I_20051 (I342765,I342717,I202016);
nor I_20052 (I342782,I342748,I202016);
nand I_20053 (I342799,I202019,I202025);
not I_20054 (I342816,I342799);
nand I_20055 (I342833,I342816,I342782);
nor I_20056 (I342850,I202034,I202028);
not I_20057 (I342867,I202022);
nor I_20058 (I342884,I342867,I202013);
nor I_20059 (I342603,I342884,I342717);
not I_20060 (I342915,I342884);
or I_20061 (I342618,I342833,I342884);
nor I_20062 (I342946,I342884,I342799);
nand I_20063 (I342615,I342748,I342946);
nor I_20064 (I342977,I342850,I342867);
nand I_20065 (I342994,I342816,I342977);
not I_20066 (I342621,I342994);
nor I_20067 (I342624,I342765,I342994);
or I_20068 (I343039,I342884,I342977);
nor I_20069 (I342609,I342816,I343039);
nor I_20070 (I343070,I342977,I202016);
nand I_20071 (I343087,I343070,I342816);
nand I_20072 (I343104,I342915,I343087);
DFFARX1 I_20073 (I343104,I1862,I342632,I342612,);
not I_20074 (I343159,I1869);
nor I_20075 (I343176,I115690,I115705);
not I_20076 (I343193,I115693);
not I_20077 (I343210,I115687);
nor I_20078 (I343227,I343210,I343176);
nand I_20079 (I343244,I343227,I115693);
not I_20080 (I343133,I343244);
nor I_20081 (I343275,I343210,I343193);
and I_20082 (I343292,I343244,I115702);
nor I_20083 (I343309,I343275,I115702);
nand I_20084 (I343326,I115687,I115696);
not I_20085 (I343343,I343326);
nand I_20086 (I343360,I343343,I343309);
nor I_20087 (I343377,I115699,I115690);
not I_20088 (I343394,I115693);
nor I_20089 (I343411,I343394,I115696);
nor I_20090 (I343130,I343411,I343244);
not I_20091 (I343442,I343411);
or I_20092 (I343145,I343360,I343411);
nor I_20093 (I343473,I343411,I343326);
nand I_20094 (I343142,I343275,I343473);
nor I_20095 (I343504,I343377,I343394);
nand I_20096 (I343521,I343343,I343504);
not I_20097 (I343148,I343521);
nor I_20098 (I343151,I343292,I343521);
or I_20099 (I343566,I343411,I343504);
nor I_20100 (I343136,I343343,I343566);
nor I_20101 (I343597,I343504,I115702);
nand I_20102 (I343614,I343597,I343343);
nand I_20103 (I343631,I343442,I343614);
DFFARX1 I_20104 (I343631,I1862,I343159,I343139,);
not I_20105 (I343686,I1869);
nor I_20106 (I343703,I122589,I122613);
not I_20107 (I343720,I122598);
not I_20108 (I343737,I122592);
nor I_20109 (I343754,I343737,I343703);
nand I_20110 (I343771,I343754,I122598);
not I_20111 (I343660,I343771);
nor I_20112 (I343802,I343737,I343720);
and I_20113 (I343819,I343771,I122595);
nor I_20114 (I343836,I343802,I122595);
nand I_20115 (I343853,I122589,I122604);
not I_20116 (I343870,I343853);
nand I_20117 (I343887,I343870,I343836);
nor I_20118 (I343904,I122601,I122592);
not I_20119 (I343921,I122610);
nor I_20120 (I343938,I343921,I122607);
nor I_20121 (I343657,I343938,I343771);
not I_20122 (I343969,I343938);
or I_20123 (I343672,I343887,I343938);
nor I_20124 (I344000,I343938,I343853);
nand I_20125 (I343669,I343802,I344000);
nor I_20126 (I344031,I343904,I343921);
nand I_20127 (I344048,I343870,I344031);
not I_20128 (I343675,I344048);
nor I_20129 (I343678,I343819,I344048);
or I_20130 (I344093,I343938,I344031);
nor I_20131 (I343663,I343870,I344093);
nor I_20132 (I344124,I344031,I122595);
nand I_20133 (I344141,I344124,I343870);
nand I_20134 (I344158,I343969,I344141);
DFFARX1 I_20135 (I344158,I1862,I343686,I343666,);
not I_20136 (I344213,I1869);
nor I_20137 (I344230,I187410,I187434);
not I_20138 (I344247,I187419);
not I_20139 (I344264,I187413);
nor I_20140 (I344281,I344264,I344230);
nand I_20141 (I344298,I344281,I187419);
not I_20142 (I344187,I344298);
nor I_20143 (I344329,I344264,I344247);
and I_20144 (I344346,I344298,I187416);
nor I_20145 (I344363,I344329,I187416);
nand I_20146 (I344380,I187410,I187425);
not I_20147 (I344397,I344380);
nand I_20148 (I344414,I344397,I344363);
nor I_20149 (I344431,I187422,I187413);
not I_20150 (I344448,I187431);
nor I_20151 (I344465,I344448,I187428);
nor I_20152 (I344184,I344465,I344298);
not I_20153 (I344496,I344465);
or I_20154 (I344199,I344414,I344465);
nor I_20155 (I344527,I344465,I344380);
nand I_20156 (I344196,I344329,I344527);
nor I_20157 (I344558,I344431,I344448);
nand I_20158 (I344575,I344397,I344558);
not I_20159 (I344202,I344575);
nor I_20160 (I344205,I344346,I344575);
or I_20161 (I344620,I344465,I344558);
nor I_20162 (I344190,I344397,I344620);
nor I_20163 (I344651,I344558,I187416);
nand I_20164 (I344668,I344651,I344397);
nand I_20165 (I344685,I344496,I344668);
DFFARX1 I_20166 (I344685,I1862,I344213,I344193,);
not I_20167 (I344740,I1869);
nor I_20168 (I344757,I198477,I198501);
not I_20169 (I344774,I198486);
not I_20170 (I344791,I198480);
nor I_20171 (I344808,I344791,I344757);
nand I_20172 (I344825,I344808,I198486);
not I_20173 (I344714,I344825);
nor I_20174 (I344856,I344791,I344774);
and I_20175 (I344873,I344825,I198483);
nor I_20176 (I344890,I344856,I198483);
nand I_20177 (I344907,I198477,I198492);
not I_20178 (I344924,I344907);
nand I_20179 (I344941,I344924,I344890);
nor I_20180 (I344958,I198489,I198480);
not I_20181 (I344975,I198498);
nor I_20182 (I344992,I344975,I198495);
nor I_20183 (I344711,I344992,I344825);
not I_20184 (I345023,I344992);
or I_20185 (I344726,I344941,I344992);
nor I_20186 (I345054,I344992,I344907);
nand I_20187 (I344723,I344856,I345054);
nor I_20188 (I345085,I344958,I344975);
nand I_20189 (I345102,I344924,I345085);
not I_20190 (I344729,I345102);
nor I_20191 (I344732,I344873,I345102);
or I_20192 (I345147,I344992,I345085);
nor I_20193 (I344717,I344924,I345147);
nor I_20194 (I345178,I345085,I198483);
nand I_20195 (I345195,I345178,I344924);
nand I_20196 (I345212,I345023,I345195);
DFFARX1 I_20197 (I345212,I1862,I344740,I344720,);
not I_20198 (I345267,I1869);
nor I_20199 (I345284,I217739,I217727);
not I_20200 (I345301,I217724);
not I_20201 (I345318,I217721);
nor I_20202 (I345335,I345318,I345284);
nand I_20203 (I345352,I345335,I217724);
not I_20204 (I345241,I345352);
nor I_20205 (I345383,I345318,I345301);
and I_20206 (I345400,I345352,I217724);
nor I_20207 (I345417,I345383,I217724);
nand I_20208 (I345434,I217727,I217733);
not I_20209 (I345451,I345434);
nand I_20210 (I345468,I345451,I345417);
nor I_20211 (I345485,I217742,I217736);
not I_20212 (I345502,I217730);
nor I_20213 (I345519,I345502,I217721);
nor I_20214 (I345238,I345519,I345352);
not I_20215 (I345550,I345519);
or I_20216 (I345253,I345468,I345519);
nor I_20217 (I345581,I345519,I345434);
nand I_20218 (I345250,I345383,I345581);
nor I_20219 (I345612,I345485,I345502);
nand I_20220 (I345629,I345451,I345612);
not I_20221 (I345256,I345629);
nor I_20222 (I345259,I345400,I345629);
or I_20223 (I345674,I345519,I345612);
nor I_20224 (I345244,I345451,I345674);
nor I_20225 (I345705,I345612,I217724);
nand I_20226 (I345722,I345705,I345451);
nand I_20227 (I345739,I345550,I345722);
DFFARX1 I_20228 (I345739,I1862,I345267,I345247,);
not I_20229 (I345794,I1869);
nor I_20230 (I345811,I84376,I84373);
not I_20231 (I345828,I84391);
not I_20232 (I345845,I84382);
nor I_20233 (I345862,I345845,I345811);
nand I_20234 (I345879,I345862,I84391);
not I_20235 (I345768,I345879);
nor I_20236 (I345910,I345845,I345828);
and I_20237 (I345927,I345879,I84397);
nor I_20238 (I345944,I345910,I84397);
nand I_20239 (I345961,I84394,I84385);
not I_20240 (I345978,I345961);
nand I_20241 (I345995,I345978,I345944);
nor I_20242 (I346012,I84373,I84376);
not I_20243 (I346029,I84388);
nor I_20244 (I346046,I346029,I84379);
nor I_20245 (I345765,I346046,I345879);
not I_20246 (I346077,I346046);
or I_20247 (I345780,I345995,I346046);
nor I_20248 (I346108,I346046,I345961);
nand I_20249 (I345777,I345910,I346108);
nor I_20250 (I346139,I346012,I346029);
nand I_20251 (I346156,I345978,I346139);
not I_20252 (I345783,I346156);
nor I_20253 (I345786,I345927,I346156);
or I_20254 (I346201,I346046,I346139);
nor I_20255 (I345771,I345978,I346201);
nor I_20256 (I346232,I346139,I84397);
nand I_20257 (I346249,I346232,I345978);
nand I_20258 (I346266,I346077,I346249);
DFFARX1 I_20259 (I346266,I1862,I345794,I345774,);
not I_20260 (I346321,I1869);
nor I_20261 (I346338,I398618,I398621);
not I_20262 (I346355,I398633);
not I_20263 (I346372,I398624);
nor I_20264 (I346389,I346372,I346338);
nand I_20265 (I346406,I346389,I398633);
not I_20266 (I346295,I346406);
nor I_20267 (I346437,I346372,I346355);
and I_20268 (I346454,I346406,I398627);
nor I_20269 (I346471,I346437,I398627);
nand I_20270 (I346488,I398624,I398630);
not I_20271 (I346505,I346488);
nand I_20272 (I346522,I346505,I346471);
nor I_20273 (I346539,I398621,I398636);
not I_20274 (I346556,I398627);
nor I_20275 (I346573,I346556,I398618);
nor I_20276 (I346292,I346573,I346406);
not I_20277 (I346604,I346573);
or I_20278 (I346307,I346522,I346573);
nor I_20279 (I346635,I346573,I346488);
nand I_20280 (I346304,I346437,I346635);
nor I_20281 (I346666,I346539,I346556);
nand I_20282 (I346683,I346505,I346666);
not I_20283 (I346310,I346683);
nor I_20284 (I346313,I346454,I346683);
or I_20285 (I346728,I346573,I346666);
nor I_20286 (I346298,I346505,I346728);
nor I_20287 (I346759,I346666,I398627);
nand I_20288 (I346776,I346759,I346505);
nand I_20289 (I346793,I346604,I346776);
DFFARX1 I_20290 (I346793,I1862,I346321,I346301,);
not I_20291 (I346848,I1869);
nor I_20292 (I346865,I302554,I302551);
not I_20293 (I346882,I302560);
not I_20294 (I346899,I302557);
nor I_20295 (I346916,I346899,I346865);
nand I_20296 (I346933,I346916,I302560);
not I_20297 (I346822,I346933);
nor I_20298 (I346964,I346899,I346882);
and I_20299 (I346981,I346933,I302563);
nor I_20300 (I346998,I346964,I302563);
nand I_20301 (I347015,I302566,I302557);
not I_20302 (I347032,I347015);
nand I_20303 (I347049,I347032,I346998);
nor I_20304 (I347066,I302572,I302569);
not I_20305 (I347083,I302551);
nor I_20306 (I347100,I347083,I302554);
nor I_20307 (I346819,I347100,I346933);
not I_20308 (I347131,I347100);
or I_20309 (I346834,I347049,I347100);
nor I_20310 (I347162,I347100,I347015);
nand I_20311 (I346831,I346964,I347162);
nor I_20312 (I347193,I347066,I347083);
nand I_20313 (I347210,I347032,I347193);
not I_20314 (I346837,I347210);
nor I_20315 (I346840,I346981,I347210);
or I_20316 (I347255,I347100,I347193);
nor I_20317 (I346825,I347032,I347255);
nor I_20318 (I347286,I347193,I302563);
nand I_20319 (I347303,I347286,I347032);
nand I_20320 (I347320,I347131,I347303);
DFFARX1 I_20321 (I347320,I1862,I346848,I346828,);
not I_20322 (I347375,I1869);
nor I_20323 (I347392,I124170,I124194);
not I_20324 (I347409,I124179);
not I_20325 (I347426,I124173);
nor I_20326 (I347443,I347426,I347392);
nand I_20327 (I347460,I347443,I124179);
not I_20328 (I347349,I347460);
nor I_20329 (I347491,I347426,I347409);
and I_20330 (I347508,I347460,I124176);
nor I_20331 (I347525,I347491,I124176);
nand I_20332 (I347542,I124170,I124185);
not I_20333 (I347559,I347542);
nand I_20334 (I347576,I347559,I347525);
nor I_20335 (I347593,I124182,I124173);
not I_20336 (I347610,I124191);
nor I_20337 (I347627,I347610,I124188);
nor I_20338 (I347346,I347627,I347460);
not I_20339 (I347658,I347627);
or I_20340 (I347361,I347576,I347627);
nor I_20341 (I347689,I347627,I347542);
nand I_20342 (I347358,I347491,I347689);
nor I_20343 (I347720,I347593,I347610);
nand I_20344 (I347737,I347559,I347720);
not I_20345 (I347364,I347737);
nor I_20346 (I347367,I347508,I347737);
or I_20347 (I347782,I347627,I347720);
nor I_20348 (I347352,I347559,I347782);
nor I_20349 (I347813,I347720,I124176);
nand I_20350 (I347830,I347813,I347559);
nand I_20351 (I347847,I347658,I347830);
DFFARX1 I_20352 (I347847,I1862,I347375,I347355,);
not I_20353 (I347902,I1869);
nor I_20354 (I347919,I279619,I279607);
not I_20355 (I347936,I279604);
not I_20356 (I347953,I279601);
nor I_20357 (I347970,I347953,I347919);
nand I_20358 (I347987,I347970,I279604);
not I_20359 (I347876,I347987);
nor I_20360 (I348018,I347953,I347936);
and I_20361 (I348035,I347987,I279604);
nor I_20362 (I348052,I348018,I279604);
nand I_20363 (I348069,I279607,I279613);
not I_20364 (I348086,I348069);
nand I_20365 (I348103,I348086,I348052);
nor I_20366 (I348120,I279622,I279616);
not I_20367 (I348137,I279610);
nor I_20368 (I348154,I348137,I279601);
nor I_20369 (I347873,I348154,I347987);
not I_20370 (I348185,I348154);
or I_20371 (I347888,I348103,I348154);
nor I_20372 (I348216,I348154,I348069);
nand I_20373 (I347885,I348018,I348216);
nor I_20374 (I348247,I348120,I348137);
nand I_20375 (I348264,I348086,I348247);
not I_20376 (I347891,I348264);
nor I_20377 (I347894,I348035,I348264);
or I_20378 (I348309,I348154,I348247);
nor I_20379 (I347879,I348086,I348309);
nor I_20380 (I348340,I348247,I279604);
nand I_20381 (I348357,I348340,I348086);
nand I_20382 (I348374,I348185,I348357);
DFFARX1 I_20383 (I348374,I1862,I347902,I347882,);
not I_20384 (I348429,I1869);
nor I_20385 (I348446,I255819,I255807);
not I_20386 (I348463,I255804);
not I_20387 (I348480,I255801);
nor I_20388 (I348497,I348480,I348446);
nand I_20389 (I348514,I348497,I255804);
not I_20390 (I348403,I348514);
nor I_20391 (I348545,I348480,I348463);
and I_20392 (I348562,I348514,I255804);
nor I_20393 (I348579,I348545,I255804);
nand I_20394 (I348596,I255807,I255813);
not I_20395 (I348613,I348596);
nand I_20396 (I348630,I348613,I348579);
nor I_20397 (I348647,I255822,I255816);
not I_20398 (I348664,I255810);
nor I_20399 (I348681,I348664,I255801);
nor I_20400 (I348400,I348681,I348514);
not I_20401 (I348712,I348681);
or I_20402 (I348415,I348630,I348681);
nor I_20403 (I348743,I348681,I348596);
nand I_20404 (I348412,I348545,I348743);
nor I_20405 (I348774,I348647,I348664);
nand I_20406 (I348791,I348613,I348774);
not I_20407 (I348418,I348791);
nor I_20408 (I348421,I348562,I348791);
or I_20409 (I348836,I348681,I348774);
nor I_20410 (I348406,I348613,I348836);
nor I_20411 (I348867,I348774,I255804);
nand I_20412 (I348884,I348867,I348613);
nand I_20413 (I348901,I348712,I348884);
DFFARX1 I_20414 (I348901,I1862,I348429,I348409,);
not I_20415 (I348956,I1869);
nor I_20416 (I348973,I361490,I361493);
not I_20417 (I348990,I361505);
not I_20418 (I349007,I361496);
nor I_20419 (I349024,I349007,I348973);
nand I_20420 (I349041,I349024,I361505);
not I_20421 (I348930,I349041);
nor I_20422 (I349072,I349007,I348990);
and I_20423 (I349089,I349041,I361499);
nor I_20424 (I349106,I349072,I361499);
nand I_20425 (I349123,I361496,I361502);
not I_20426 (I349140,I349123);
nand I_20427 (I349157,I349140,I349106);
nor I_20428 (I349174,I361493,I361508);
not I_20429 (I349191,I361499);
nor I_20430 (I349208,I349191,I361490);
nor I_20431 (I348927,I349208,I349041);
not I_20432 (I349239,I349208);
or I_20433 (I348942,I349157,I349208);
nor I_20434 (I349270,I349208,I349123);
nand I_20435 (I348939,I349072,I349270);
nor I_20436 (I349301,I349174,I349191);
nand I_20437 (I349318,I349140,I349301);
not I_20438 (I348945,I349318);
nor I_20439 (I348948,I349089,I349318);
or I_20440 (I349363,I349208,I349301);
nor I_20441 (I348933,I349140,I349363);
nor I_20442 (I349394,I349301,I361499);
nand I_20443 (I349411,I349394,I349140);
nand I_20444 (I349428,I349239,I349411);
DFFARX1 I_20445 (I349428,I1862,I348956,I348936,);
not I_20446 (I349483,I1869);
nor I_20447 (I349500,I26236,I26233);
not I_20448 (I349517,I26251);
not I_20449 (I349534,I26242);
nor I_20450 (I349551,I349534,I349500);
nand I_20451 (I349568,I349551,I26251);
not I_20452 (I349457,I349568);
nor I_20453 (I349599,I349534,I349517);
and I_20454 (I349616,I349568,I26257);
nor I_20455 (I349633,I349599,I26257);
nand I_20456 (I349650,I26254,I26245);
not I_20457 (I349667,I349650);
nand I_20458 (I349684,I349667,I349633);
nor I_20459 (I349701,I26233,I26236);
not I_20460 (I349718,I26248);
nor I_20461 (I349735,I349718,I26239);
nor I_20462 (I349454,I349735,I349568);
not I_20463 (I349766,I349735);
or I_20464 (I349469,I349684,I349735);
nor I_20465 (I349797,I349735,I349650);
nand I_20466 (I349466,I349599,I349797);
nor I_20467 (I349828,I349701,I349718);
nand I_20468 (I349845,I349667,I349828);
not I_20469 (I349472,I349845);
nor I_20470 (I349475,I349616,I349845);
or I_20471 (I349890,I349735,I349828);
nor I_20472 (I349460,I349667,I349890);
nor I_20473 (I349921,I349828,I26257);
nand I_20474 (I349938,I349921,I349667);
nand I_20475 (I349955,I349766,I349938);
DFFARX1 I_20476 (I349955,I1862,I349483,I349463,);
not I_20477 (I350010,I1869);
nor I_20478 (I350027,I237255,I237243);
not I_20479 (I350044,I237240);
not I_20480 (I350061,I237237);
nor I_20481 (I350078,I350061,I350027);
nand I_20482 (I350095,I350078,I237240);
not I_20483 (I349984,I350095);
nor I_20484 (I350126,I350061,I350044);
and I_20485 (I350143,I350095,I237240);
nor I_20486 (I350160,I350126,I237240);
nand I_20487 (I350177,I237243,I237249);
not I_20488 (I350194,I350177);
nand I_20489 (I350211,I350194,I350160);
nor I_20490 (I350228,I237258,I237252);
not I_20491 (I350245,I237246);
nor I_20492 (I350262,I350245,I237237);
nor I_20493 (I349981,I350262,I350095);
not I_20494 (I350293,I350262);
or I_20495 (I349996,I350211,I350262);
nor I_20496 (I350324,I350262,I350177);
nand I_20497 (I349993,I350126,I350324);
nor I_20498 (I350355,I350228,I350245);
nand I_20499 (I350372,I350194,I350355);
not I_20500 (I349999,I350372);
nor I_20501 (I350002,I350143,I350372);
or I_20502 (I350417,I350262,I350355);
nor I_20503 (I349987,I350194,I350417);
nor I_20504 (I350448,I350355,I237240);
nand I_20505 (I350465,I350448,I350194);
nand I_20506 (I350482,I350293,I350465);
DFFARX1 I_20507 (I350482,I1862,I350010,I349990,);
not I_20508 (I350537,I1869);
nor I_20509 (I350554,I211551,I211539);
not I_20510 (I350571,I211536);
not I_20511 (I350588,I211533);
nor I_20512 (I350605,I350588,I350554);
nand I_20513 (I350622,I350605,I211536);
not I_20514 (I350511,I350622);
nor I_20515 (I350653,I350588,I350571);
and I_20516 (I350670,I350622,I211536);
nor I_20517 (I350687,I350653,I211536);
nand I_20518 (I350704,I211539,I211545);
not I_20519 (I350721,I350704);
nand I_20520 (I350738,I350721,I350687);
nor I_20521 (I350755,I211554,I211548);
not I_20522 (I350772,I211542);
nor I_20523 (I350789,I350772,I211533);
nor I_20524 (I350508,I350789,I350622);
not I_20525 (I350820,I350789);
or I_20526 (I350523,I350738,I350789);
nor I_20527 (I350851,I350789,I350704);
nand I_20528 (I350520,I350653,I350851);
nor I_20529 (I350882,I350755,I350772);
nand I_20530 (I350899,I350721,I350882);
not I_20531 (I350526,I350899);
nor I_20532 (I350529,I350670,I350899);
or I_20533 (I350944,I350789,I350882);
nor I_20534 (I350514,I350721,I350944);
nor I_20535 (I350975,I350882,I211536);
nand I_20536 (I350992,I350975,I350721);
nand I_20537 (I351009,I350820,I350992);
DFFARX1 I_20538 (I351009,I1862,I350537,I350517,);
not I_20539 (I351064,I1869);
nor I_20540 (I351081,I219167,I219155);
not I_20541 (I351098,I219152);
not I_20542 (I351115,I219149);
nor I_20543 (I351132,I351115,I351081);
nand I_20544 (I351149,I351132,I219152);
not I_20545 (I351038,I351149);
nor I_20546 (I351180,I351115,I351098);
and I_20547 (I351197,I351149,I219152);
nor I_20548 (I351214,I351180,I219152);
nand I_20549 (I351231,I219155,I219161);
not I_20550 (I351248,I351231);
nand I_20551 (I351265,I351248,I351214);
nor I_20552 (I351282,I219170,I219164);
not I_20553 (I351299,I219158);
nor I_20554 (I351316,I351299,I219149);
nor I_20555 (I351035,I351316,I351149);
not I_20556 (I351347,I351316);
or I_20557 (I351050,I351265,I351316);
nor I_20558 (I351378,I351316,I351231);
nand I_20559 (I351047,I351180,I351378);
nor I_20560 (I351409,I351282,I351299);
nand I_20561 (I351426,I351248,I351409);
not I_20562 (I351053,I351426);
nor I_20563 (I351056,I351197,I351426);
or I_20564 (I351471,I351316,I351409);
nor I_20565 (I351041,I351248,I351471);
nor I_20566 (I351502,I351409,I219152);
nand I_20567 (I351519,I351502,I351248);
nand I_20568 (I351536,I351347,I351519);
DFFARX1 I_20569 (I351536,I1862,I351064,I351044,);
not I_20570 (I351591,I1869);
nor I_20571 (I351608,I142088,I142112);
not I_20572 (I351625,I142097);
not I_20573 (I351642,I142091);
nor I_20574 (I351659,I351642,I351608);
nand I_20575 (I351676,I351659,I142097);
not I_20576 (I351565,I351676);
nor I_20577 (I351707,I351642,I351625);
and I_20578 (I351724,I351676,I142094);
nor I_20579 (I351741,I351707,I142094);
nand I_20580 (I351758,I142088,I142103);
not I_20581 (I351775,I351758);
nand I_20582 (I351792,I351775,I351741);
nor I_20583 (I351809,I142100,I142091);
not I_20584 (I351826,I142109);
nor I_20585 (I351843,I351826,I142106);
nor I_20586 (I351562,I351843,I351676);
not I_20587 (I351874,I351843);
or I_20588 (I351577,I351792,I351843);
nor I_20589 (I351905,I351843,I351758);
nand I_20590 (I351574,I351707,I351905);
nor I_20591 (I351936,I351809,I351826);
nand I_20592 (I351953,I351775,I351936);
not I_20593 (I351580,I351953);
nor I_20594 (I351583,I351724,I351953);
or I_20595 (I351998,I351843,I351936);
nor I_20596 (I351568,I351775,I351998);
nor I_20597 (I352029,I351936,I142094);
nand I_20598 (I352046,I352029,I351775);
nand I_20599 (I352063,I351874,I352046);
DFFARX1 I_20600 (I352063,I1862,I351591,I351571,);
not I_20601 (I352118,I1869);
nor I_20602 (I352135,I295176,I295173);
not I_20603 (I352152,I295182);
not I_20604 (I352169,I295179);
nor I_20605 (I352186,I352169,I352135);
nand I_20606 (I352203,I352186,I295182);
not I_20607 (I352092,I352203);
nor I_20608 (I352234,I352169,I352152);
and I_20609 (I352251,I352203,I295185);
nor I_20610 (I352268,I352234,I295185);
nand I_20611 (I352285,I295188,I295179);
not I_20612 (I352302,I352285);
nand I_20613 (I352319,I352302,I352268);
nor I_20614 (I352336,I295194,I295191);
not I_20615 (I352353,I295173);
nor I_20616 (I352370,I352353,I295176);
nor I_20617 (I352089,I352370,I352203);
not I_20618 (I352401,I352370);
or I_20619 (I352104,I352319,I352370);
nor I_20620 (I352432,I352370,I352285);
nand I_20621 (I352101,I352234,I352432);
nor I_20622 (I352463,I352336,I352353);
nand I_20623 (I352480,I352302,I352463);
not I_20624 (I352107,I352480);
nor I_20625 (I352110,I352251,I352480);
or I_20626 (I352525,I352370,I352463);
nor I_20627 (I352095,I352302,I352525);
nor I_20628 (I352556,I352463,I295185);
nand I_20629 (I352573,I352556,I352302);
nand I_20630 (I352590,I352401,I352573);
DFFARX1 I_20631 (I352590,I1862,I352118,I352098,);
not I_20632 (I352645,I1869);
nor I_20633 (I352662,I1239,I1311);
not I_20634 (I352679,I1167);
not I_20635 (I352696,I1615);
nor I_20636 (I352713,I352696,I352662);
nand I_20637 (I352730,I352713,I1167);
not I_20638 (I352619,I352730);
nor I_20639 (I352761,I352696,I352679);
and I_20640 (I352778,I352730,I1335);
nor I_20641 (I352795,I352761,I1335);
nand I_20642 (I352812,I671,I1655);
not I_20643 (I352829,I352812);
nand I_20644 (I352846,I352829,I352795);
nor I_20645 (I352863,I1319,I863);
not I_20646 (I352880,I855);
nor I_20647 (I352897,I352880,I1551);
nor I_20648 (I352616,I352897,I352730);
not I_20649 (I352928,I352897);
or I_20650 (I352631,I352846,I352897);
nor I_20651 (I352959,I352897,I352812);
nand I_20652 (I352628,I352761,I352959);
nor I_20653 (I352990,I352863,I352880);
nand I_20654 (I353007,I352829,I352990);
not I_20655 (I352634,I353007);
nor I_20656 (I352637,I352778,I353007);
or I_20657 (I353052,I352897,I352990);
nor I_20658 (I352622,I352829,I353052);
nor I_20659 (I353083,I352990,I1335);
nand I_20660 (I353100,I353083,I352829);
nand I_20661 (I353117,I352928,I353100);
DFFARX1 I_20662 (I353117,I1862,I352645,I352625,);
not I_20663 (I353172,I1869);
nor I_20664 (I353189,I119427,I119451);
not I_20665 (I353206,I119436);
not I_20666 (I353223,I119430);
nor I_20667 (I353240,I353223,I353189);
nand I_20668 (I353257,I353240,I119436);
not I_20669 (I353146,I353257);
nor I_20670 (I353288,I353223,I353206);
and I_20671 (I353305,I353257,I119433);
nor I_20672 (I353322,I353288,I119433);
nand I_20673 (I353339,I119427,I119442);
not I_20674 (I353356,I353339);
nand I_20675 (I353373,I353356,I353322);
nor I_20676 (I353390,I119439,I119430);
not I_20677 (I353407,I119448);
nor I_20678 (I353424,I353407,I119445);
nor I_20679 (I353143,I353424,I353257);
not I_20680 (I353455,I353424);
or I_20681 (I353158,I353373,I353424);
nor I_20682 (I353486,I353424,I353339);
nand I_20683 (I353155,I353288,I353486);
nor I_20684 (I353517,I353390,I353407);
nand I_20685 (I353534,I353356,I353517);
not I_20686 (I353161,I353534);
nor I_20687 (I353164,I353305,I353534);
or I_20688 (I353579,I353424,I353517);
nor I_20689 (I353149,I353356,I353579);
nor I_20690 (I353610,I353517,I119433);
nand I_20691 (I353627,I353610,I353356);
nand I_20692 (I353644,I353455,I353627);
DFFARX1 I_20693 (I353644,I1862,I353172,I353152,);
not I_20694 (I353699,I1869);
nor I_20695 (I353716,I113650,I113665);
not I_20696 (I353733,I113653);
not I_20697 (I353750,I113647);
nor I_20698 (I353767,I353750,I353716);
nand I_20699 (I353784,I353767,I113653);
not I_20700 (I353673,I353784);
nor I_20701 (I353815,I353750,I353733);
and I_20702 (I353832,I353784,I113662);
nor I_20703 (I353849,I353815,I113662);
nand I_20704 (I353866,I113647,I113656);
not I_20705 (I353883,I353866);
nand I_20706 (I353900,I353883,I353849);
nor I_20707 (I353917,I113659,I113650);
not I_20708 (I353934,I113653);
nor I_20709 (I353951,I353934,I113656);
nor I_20710 (I353670,I353951,I353784);
not I_20711 (I353982,I353951);
or I_20712 (I353685,I353900,I353951);
nor I_20713 (I354013,I353951,I353866);
nand I_20714 (I353682,I353815,I354013);
nor I_20715 (I354044,I353917,I353934);
nand I_20716 (I354061,I353883,I354044);
not I_20717 (I353688,I354061);
nor I_20718 (I353691,I353832,I354061);
or I_20719 (I354106,I353951,I354044);
nor I_20720 (I353676,I353883,I354106);
nor I_20721 (I354137,I354044,I113662);
nand I_20722 (I354154,I354137,I353883);
nand I_20723 (I354171,I353982,I354154);
DFFARX1 I_20724 (I354171,I1862,I353699,I353679,);
not I_20725 (I354226,I1869);
nor I_20726 (I354243,I148939,I148963);
not I_20727 (I354260,I148948);
not I_20728 (I354277,I148942);
nor I_20729 (I354294,I354277,I354243);
nand I_20730 (I354311,I354294,I148948);
not I_20731 (I354200,I354311);
nor I_20732 (I354342,I354277,I354260);
and I_20733 (I354359,I354311,I148945);
nor I_20734 (I354376,I354342,I148945);
nand I_20735 (I354393,I148939,I148954);
not I_20736 (I354410,I354393);
nand I_20737 (I354427,I354410,I354376);
nor I_20738 (I354444,I148951,I148942);
not I_20739 (I354461,I148960);
nor I_20740 (I354478,I354461,I148957);
nor I_20741 (I354197,I354478,I354311);
not I_20742 (I354509,I354478);
or I_20743 (I354212,I354427,I354478);
nor I_20744 (I354540,I354478,I354393);
nand I_20745 (I354209,I354342,I354540);
nor I_20746 (I354571,I354444,I354461);
nand I_20747 (I354588,I354410,I354571);
not I_20748 (I354215,I354588);
nor I_20749 (I354218,I354359,I354588);
or I_20750 (I354633,I354478,I354571);
nor I_20751 (I354203,I354410,I354633);
nor I_20752 (I354664,I354571,I148945);
nand I_20753 (I354681,I354664,I354410);
nand I_20754 (I354698,I354509,I354681);
DFFARX1 I_20755 (I354698,I1862,I354226,I354206,);
not I_20756 (I354753,I1869);
nor I_20757 (I354770,I376960,I376963);
not I_20758 (I354787,I376975);
not I_20759 (I354804,I376966);
nor I_20760 (I354821,I354804,I354770);
nand I_20761 (I354838,I354821,I376975);
not I_20762 (I354727,I354838);
nor I_20763 (I354869,I354804,I354787);
and I_20764 (I354886,I354838,I376969);
nor I_20765 (I354903,I354869,I376969);
nand I_20766 (I354920,I376966,I376972);
not I_20767 (I354937,I354920);
nand I_20768 (I354954,I354937,I354903);
nor I_20769 (I354971,I376963,I376978);
not I_20770 (I354988,I376969);
nor I_20771 (I355005,I354988,I376960);
nor I_20772 (I354724,I355005,I354838);
not I_20773 (I355036,I355005);
or I_20774 (I354739,I354954,I355005);
nor I_20775 (I355067,I355005,I354920);
nand I_20776 (I354736,I354869,I355067);
nor I_20777 (I355098,I354971,I354988);
nand I_20778 (I355115,I354937,I355098);
not I_20779 (I354742,I355115);
nor I_20780 (I354745,I354886,I355115);
or I_20781 (I355160,I355005,I355098);
nor I_20782 (I354730,I354937,I355160);
nor I_20783 (I355191,I355098,I376969);
nand I_20784 (I355208,I355191,I354937);
nand I_20785 (I355225,I355036,I355208);
DFFARX1 I_20786 (I355225,I1862,I354753,I354733,);
not I_20787 (I355280,I1869);
nor I_20788 (I355297,I141561,I141585);
not I_20789 (I355314,I141570);
not I_20790 (I355331,I141564);
nor I_20791 (I355348,I355331,I355297);
nand I_20792 (I355365,I355348,I141570);
not I_20793 (I355254,I355365);
nor I_20794 (I355396,I355331,I355314);
and I_20795 (I355413,I355365,I141567);
nor I_20796 (I355430,I355396,I141567);
nand I_20797 (I355447,I141561,I141576);
not I_20798 (I355464,I355447);
nand I_20799 (I355481,I355464,I355430);
nor I_20800 (I355498,I141573,I141564);
not I_20801 (I355515,I141582);
nor I_20802 (I355532,I355515,I141579);
nor I_20803 (I355251,I355532,I355365);
not I_20804 (I355563,I355532);
or I_20805 (I355266,I355481,I355532);
nor I_20806 (I355594,I355532,I355447);
nand I_20807 (I355263,I355396,I355594);
nor I_20808 (I355625,I355498,I355515);
nand I_20809 (I355642,I355464,I355625);
not I_20810 (I355269,I355642);
nor I_20811 (I355272,I355413,I355642);
or I_20812 (I355687,I355532,I355625);
nor I_20813 (I355257,I355464,I355687);
nor I_20814 (I355718,I355625,I141567);
nand I_20815 (I355735,I355718,I355464);
nand I_20816 (I355752,I355563,I355735);
DFFARX1 I_20817 (I355752,I1862,I355280,I355260,);
not I_20818 (I355807,I1869);
nor I_20819 (I355824,I151047,I151071);
not I_20820 (I355841,I151056);
not I_20821 (I355858,I151050);
nor I_20822 (I355875,I355858,I355824);
nand I_20823 (I355892,I355875,I151056);
not I_20824 (I355781,I355892);
nor I_20825 (I355923,I355858,I355841);
and I_20826 (I355940,I355892,I151053);
nor I_20827 (I355957,I355923,I151053);
nand I_20828 (I355974,I151047,I151062);
not I_20829 (I355991,I355974);
nand I_20830 (I356008,I355991,I355957);
nor I_20831 (I356025,I151059,I151050);
not I_20832 (I356042,I151068);
nor I_20833 (I356059,I356042,I151065);
nor I_20834 (I355778,I356059,I355892);
not I_20835 (I356090,I356059);
or I_20836 (I355793,I356008,I356059);
nor I_20837 (I356121,I356059,I355974);
nand I_20838 (I355790,I355923,I356121);
nor I_20839 (I356152,I356025,I356042);
nand I_20840 (I356169,I355991,I356152);
not I_20841 (I355796,I356169);
nor I_20842 (I355799,I355940,I356169);
or I_20843 (I356214,I356059,I356152);
nor I_20844 (I355784,I355991,I356214);
nor I_20845 (I356245,I356152,I151053);
nand I_20846 (I356262,I356245,I355991);
nand I_20847 (I356279,I356090,I356262);
DFFARX1 I_20848 (I356279,I1862,I355807,I355787,);
not I_20849 (I356334,I1869);
nor I_20850 (I356351,I399944,I399947);
not I_20851 (I356368,I399959);
not I_20852 (I356385,I399950);
nor I_20853 (I356402,I356385,I356351);
nand I_20854 (I356419,I356402,I399959);
not I_20855 (I356308,I356419);
nor I_20856 (I356450,I356385,I356368);
and I_20857 (I356467,I356419,I399953);
nor I_20858 (I356484,I356450,I399953);
nand I_20859 (I356501,I399950,I399956);
not I_20860 (I356518,I356501);
nand I_20861 (I356535,I356518,I356484);
nor I_20862 (I356552,I399947,I399962);
not I_20863 (I356569,I399953);
nor I_20864 (I356586,I356569,I399944);
nor I_20865 (I356305,I356586,I356419);
not I_20866 (I356617,I356586);
or I_20867 (I356320,I356535,I356586);
nor I_20868 (I356648,I356586,I356501);
nand I_20869 (I356317,I356450,I356648);
nor I_20870 (I356679,I356552,I356569);
nand I_20871 (I356696,I356518,I356679);
not I_20872 (I356323,I356696);
nor I_20873 (I356326,I356467,I356696);
or I_20874 (I356741,I356586,I356679);
nor I_20875 (I356311,I356518,I356741);
nor I_20876 (I356772,I356679,I399953);
nand I_20877 (I356789,I356772,I356518);
nand I_20878 (I356806,I356617,I356789);
DFFARX1 I_20879 (I356806,I1862,I356334,I356314,);
not I_20880 (I356861,I1869);
nor I_20881 (I356878,I400386,I400389);
not I_20882 (I356895,I400401);
not I_20883 (I356912,I400392);
nor I_20884 (I356929,I356912,I356878);
nand I_20885 (I356946,I356929,I400401);
not I_20886 (I356835,I356946);
nor I_20887 (I356977,I356912,I356895);
and I_20888 (I356994,I356946,I400395);
nor I_20889 (I357011,I356977,I400395);
nand I_20890 (I357028,I400392,I400398);
not I_20891 (I357045,I357028);
nand I_20892 (I357062,I357045,I357011);
nor I_20893 (I357079,I400389,I400404);
not I_20894 (I357096,I400395);
nor I_20895 (I357113,I357096,I400386);
nor I_20896 (I356832,I357113,I356946);
not I_20897 (I357144,I357113);
or I_20898 (I356847,I357062,I357113);
nor I_20899 (I357175,I357113,I357028);
nand I_20900 (I356844,I356977,I357175);
nor I_20901 (I357206,I357079,I357096);
nand I_20902 (I357223,I357045,I357206);
not I_20903 (I356850,I357223);
nor I_20904 (I356853,I356994,I357223);
or I_20905 (I357268,I357113,I357206);
nor I_20906 (I356838,I357045,I357268);
nor I_20907 (I357299,I357206,I400395);
nand I_20908 (I357316,I357299,I357045);
nand I_20909 (I357333,I357144,I357316);
DFFARX1 I_20910 (I357333,I1862,I356861,I356841,);
not I_20911 (I357388,I1869);
nor I_20912 (I357405,I242967,I242955);
not I_20913 (I357422,I242952);
not I_20914 (I357439,I242949);
nor I_20915 (I357456,I357439,I357405);
nand I_20916 (I357473,I357456,I242952);
not I_20917 (I357362,I357473);
nor I_20918 (I357504,I357439,I357422);
and I_20919 (I357521,I357473,I242952);
nor I_20920 (I357538,I357504,I242952);
nand I_20921 (I357555,I242955,I242961);
not I_20922 (I357572,I357555);
nand I_20923 (I357589,I357572,I357538);
nor I_20924 (I357606,I242970,I242964);
not I_20925 (I357623,I242958);
nor I_20926 (I357640,I357623,I242949);
nor I_20927 (I357359,I357640,I357473);
not I_20928 (I357671,I357640);
or I_20929 (I357374,I357589,I357640);
nor I_20930 (I357702,I357640,I357555);
nand I_20931 (I357371,I357504,I357702);
nor I_20932 (I357733,I357606,I357623);
nand I_20933 (I357750,I357572,I357733);
not I_20934 (I357377,I357750);
nor I_20935 (I357380,I357521,I357750);
or I_20936 (I357795,I357640,I357733);
nor I_20937 (I357365,I357572,I357795);
nor I_20938 (I357826,I357733,I242952);
nand I_20939 (I357843,I357826,I357572);
nand I_20940 (I357860,I357671,I357843);
DFFARX1 I_20941 (I357860,I1862,I357388,I357368,);
not I_20942 (I357915,I1869);
nor I_20943 (I357932,I242491,I242479);
not I_20944 (I357949,I242476);
not I_20945 (I357966,I242473);
nor I_20946 (I357983,I357966,I357932);
nand I_20947 (I358000,I357983,I242476);
not I_20948 (I357889,I358000);
nor I_20949 (I358031,I357966,I357949);
and I_20950 (I358048,I358000,I242476);
nor I_20951 (I358065,I358031,I242476);
nand I_20952 (I358082,I242479,I242485);
not I_20953 (I358099,I358082);
nand I_20954 (I358116,I358099,I358065);
nor I_20955 (I358133,I242494,I242488);
not I_20956 (I358150,I242482);
nor I_20957 (I358167,I358150,I242473);
nor I_20958 (I357886,I358167,I358000);
not I_20959 (I358198,I358167);
or I_20960 (I357901,I358116,I358167);
nor I_20961 (I358229,I358167,I358082);
nand I_20962 (I357898,I358031,I358229);
nor I_20963 (I358260,I358133,I358150);
nand I_20964 (I358277,I358099,I358260);
not I_20965 (I357904,I358277);
nor I_20966 (I357907,I358048,I358277);
or I_20967 (I358322,I358167,I358260);
nor I_20968 (I357892,I358099,I358322);
nor I_20969 (I358353,I358260,I242476);
nand I_20970 (I358370,I358353,I358099);
nand I_20971 (I358387,I358198,I358370);
DFFARX1 I_20972 (I358387,I1862,I357915,I357895,);
not I_20973 (I358442,I1869);
nor I_20974 (I358459,I140507,I140531);
not I_20975 (I358476,I140516);
not I_20976 (I358493,I140510);
nor I_20977 (I358510,I358493,I358459);
nand I_20978 (I358527,I358510,I140516);
not I_20979 (I358416,I358527);
nor I_20980 (I358558,I358493,I358476);
and I_20981 (I358575,I358527,I140513);
nor I_20982 (I358592,I358558,I140513);
nand I_20983 (I358609,I140507,I140522);
not I_20984 (I358626,I358609);
nand I_20985 (I358643,I358626,I358592);
nor I_20986 (I358660,I140519,I140510);
not I_20987 (I358677,I140528);
nor I_20988 (I358694,I358677,I140525);
nor I_20989 (I358413,I358694,I358527);
not I_20990 (I358725,I358694);
or I_20991 (I358428,I358643,I358694);
nor I_20992 (I358756,I358694,I358609);
nand I_20993 (I358425,I358558,I358756);
nor I_20994 (I358787,I358660,I358677);
nand I_20995 (I358804,I358626,I358787);
not I_20996 (I358431,I358804);
nor I_20997 (I358434,I358575,I358804);
or I_20998 (I358849,I358694,I358787);
nor I_20999 (I358419,I358626,I358849);
nor I_21000 (I358880,I358787,I140513);
nand I_21001 (I358897,I358880,I358626);
nand I_21002 (I358914,I358725,I358897);
DFFARX1 I_21003 (I358914,I1862,I358442,I358422,);
not I_21004 (I358969,I1869);
nor I_21005 (I358986,I373866,I373869);
not I_21006 (I359003,I373881);
not I_21007 (I359020,I373872);
nor I_21008 (I359037,I359020,I358986);
nand I_21009 (I359054,I359037,I373881);
not I_21010 (I358943,I359054);
nor I_21011 (I359085,I359020,I359003);
and I_21012 (I359102,I359054,I373875);
nor I_21013 (I359119,I359085,I373875);
nand I_21014 (I359136,I373872,I373878);
not I_21015 (I359153,I359136);
nand I_21016 (I359170,I359153,I359119);
nor I_21017 (I359187,I373869,I373884);
not I_21018 (I359204,I373875);
nor I_21019 (I359221,I359204,I373866);
nor I_21020 (I358940,I359221,I359054);
not I_21021 (I359252,I359221);
or I_21022 (I358955,I359170,I359221);
nor I_21023 (I359283,I359221,I359136);
nand I_21024 (I358952,I359085,I359283);
nor I_21025 (I359314,I359187,I359204);
nand I_21026 (I359331,I359153,I359314);
not I_21027 (I358958,I359331);
nor I_21028 (I358961,I359102,I359331);
or I_21029 (I359376,I359221,I359314);
nor I_21030 (I358946,I359153,I359376);
nor I_21031 (I359407,I359314,I373875);
nand I_21032 (I359424,I359407,I359153);
nand I_21033 (I359441,I359252,I359424);
DFFARX1 I_21034 (I359441,I1862,I358969,I358949,);
not I_21035 (I359496,I1869);
nor I_21036 (I359513,I77746,I77743);
not I_21037 (I359530,I77761);
not I_21038 (I359547,I77752);
nor I_21039 (I359564,I359547,I359513);
nand I_21040 (I359581,I359564,I77761);
not I_21041 (I359470,I359581);
nor I_21042 (I359612,I359547,I359530);
and I_21043 (I359629,I359581,I77767);
nor I_21044 (I359646,I359612,I77767);
nand I_21045 (I359663,I77764,I77755);
not I_21046 (I359680,I359663);
nand I_21047 (I359697,I359680,I359646);
nor I_21048 (I359714,I77743,I77746);
not I_21049 (I359731,I77758);
nor I_21050 (I359748,I359731,I77749);
nor I_21051 (I359467,I359748,I359581);
not I_21052 (I359779,I359748);
or I_21053 (I359482,I359697,I359748);
nor I_21054 (I359810,I359748,I359663);
nand I_21055 (I359479,I359612,I359810);
nor I_21056 (I359841,I359714,I359731);
nand I_21057 (I359858,I359680,I359841);
not I_21058 (I359485,I359858);
nor I_21059 (I359488,I359629,I359858);
or I_21060 (I359903,I359748,I359841);
nor I_21061 (I359473,I359680,I359903);
nor I_21062 (I359934,I359841,I77767);
nand I_21063 (I359951,I359934,I359680);
nand I_21064 (I359968,I359779,I359951);
DFFARX1 I_21065 (I359968,I1862,I359496,I359476,);
not I_21066 (I360023,I1869);
nor I_21067 (I360040,I60916,I60913);
not I_21068 (I360057,I60931);
not I_21069 (I360074,I60922);
nor I_21070 (I360091,I360074,I360040);
nand I_21071 (I360108,I360091,I60931);
not I_21072 (I359997,I360108);
nor I_21073 (I360139,I360074,I360057);
and I_21074 (I360156,I360108,I60937);
nor I_21075 (I360173,I360139,I60937);
nand I_21076 (I360190,I60934,I60925);
not I_21077 (I360207,I360190);
nand I_21078 (I360224,I360207,I360173);
nor I_21079 (I360241,I60913,I60916);
not I_21080 (I360258,I60928);
nor I_21081 (I360275,I360258,I60919);
nor I_21082 (I359994,I360275,I360108);
not I_21083 (I360306,I360275);
or I_21084 (I360009,I360224,I360275);
nor I_21085 (I360337,I360275,I360190);
nand I_21086 (I360006,I360139,I360337);
nor I_21087 (I360368,I360241,I360258);
nand I_21088 (I360385,I360207,I360368);
not I_21089 (I360012,I360385);
nor I_21090 (I360015,I360156,I360385);
or I_21091 (I360430,I360275,I360368);
nor I_21092 (I360000,I360207,I360430);
nor I_21093 (I360461,I360368,I60937);
nand I_21094 (I360478,I360461,I360207);
nand I_21095 (I360495,I360306,I360478);
DFFARX1 I_21096 (I360495,I1862,I360023,I360003,);
not I_21097 (I360550,I1869);
nor I_21098 (I360567,I262007,I261995);
not I_21099 (I360584,I261992);
not I_21100 (I360601,I261989);
nor I_21101 (I360618,I360601,I360567);
nand I_21102 (I360635,I360618,I261992);
not I_21103 (I360524,I360635);
nor I_21104 (I360666,I360601,I360584);
and I_21105 (I360683,I360635,I261992);
nor I_21106 (I360700,I360666,I261992);
nand I_21107 (I360717,I261995,I262001);
not I_21108 (I360734,I360717);
nand I_21109 (I360751,I360734,I360700);
nor I_21110 (I360768,I262010,I262004);
not I_21111 (I360785,I261998);
nor I_21112 (I360802,I360785,I261989);
nor I_21113 (I360521,I360802,I360635);
not I_21114 (I360833,I360802);
or I_21115 (I360536,I360751,I360802);
nor I_21116 (I360864,I360802,I360717);
nand I_21117 (I360533,I360666,I360864);
nor I_21118 (I360895,I360768,I360785);
nand I_21119 (I360912,I360734,I360895);
not I_21120 (I360539,I360912);
nor I_21121 (I360542,I360683,I360912);
or I_21122 (I360957,I360802,I360895);
nor I_21123 (I360527,I360734,I360957);
nor I_21124 (I360988,I360895,I261992);
nand I_21125 (I361005,I360988,I360734);
nand I_21126 (I361022,I360833,I361005);
DFFARX1 I_21127 (I361022,I1862,I360550,I360530,);
not I_21128 (I361074,I1869);
and I_21129 (I361091,I243913,I243919);
nor I_21130 (I361108,I361091,I243907);
nand I_21131 (I361125,I243904,I243901);
nor I_21132 (I361142,I361125,I361108);
not I_21133 (I361063,I361142);
not I_21134 (I361173,I361125);
or I_21135 (I361190,I243910,I243922);
nor I_21136 (I361207,I361190,I243904);
nor I_21137 (I361224,I361207,I361173);
nand I_21138 (I361241,I243901,I243916);
nor I_21139 (I361258,I361241,I243907);
not I_21140 (I361275,I361258);
nor I_21141 (I361292,I361142,I361275);
nand I_21142 (I361060,I361292,I361207);
nor I_21143 (I361048,I361275,I361224);
nand I_21144 (I361054,I361207,I361275);
nor I_21145 (I361351,I361142,I361241);
nand I_21146 (I361368,I361351,I361207);
nand I_21147 (I361385,I361275,I361368);
DFFARX1 I_21148 (I361385,I1862,I361074,I361057,);
not I_21149 (I361416,I361241);
or I_21150 (I361433,I361207,I361416);
nor I_21151 (I361051,I361173,I361433);
nor I_21152 (I361464,I361142,I361416);
nand I_21153 (I361066,I361464,I361173);
not I_21154 (I361516,I1869);
and I_21155 (I361533,I328919,I328904);
nor I_21156 (I361550,I361533,I328907);
nand I_21157 (I361567,I328901,I328901);
nor I_21158 (I361584,I361567,I361550);
not I_21159 (I361505,I361584);
not I_21160 (I361615,I361567);
or I_21161 (I361632,I328904,I328922);
nor I_21162 (I361649,I361632,I328913);
nor I_21163 (I361666,I361649,I361615);
nand I_21164 (I361683,I328916,I328910);
nor I_21165 (I361700,I361683,I328907);
not I_21166 (I361717,I361700);
nor I_21167 (I361734,I361584,I361717);
nand I_21168 (I361502,I361734,I361649);
nor I_21169 (I361490,I361717,I361666);
nand I_21170 (I361496,I361649,I361717);
nor I_21171 (I361793,I361584,I361683);
nand I_21172 (I361810,I361793,I361649);
nand I_21173 (I361827,I361717,I361810);
DFFARX1 I_21174 (I361827,I1862,I361516,I361499,);
not I_21175 (I361858,I361683);
or I_21176 (I361875,I361649,I361858);
nor I_21177 (I361493,I361615,I361875);
nor I_21178 (I361906,I361584,I361858);
nand I_21179 (I361508,I361906,I361615);
not I_21180 (I361958,I1869);
and I_21181 (I361975,I37987,I37963);
nor I_21182 (I361992,I361975,I37969);
nand I_21183 (I362009,I37984,I37966);
nor I_21184 (I362026,I362009,I361992);
not I_21185 (I361947,I362026);
not I_21186 (I362057,I362009);
or I_21187 (I362074,I37963,I37966);
nor I_21188 (I362091,I362074,I37978);
nor I_21189 (I362108,I362091,I362057);
nand I_21190 (I362125,I37972,I37975);
nor I_21191 (I362142,I362125,I37981);
not I_21192 (I362159,I362142);
nor I_21193 (I362176,I362026,I362159);
nand I_21194 (I361944,I362176,I362091);
nor I_21195 (I361932,I362159,I362108);
nand I_21196 (I361938,I362091,I362159);
nor I_21197 (I362235,I362026,I362125);
nand I_21198 (I362252,I362235,I362091);
nand I_21199 (I362269,I362159,I362252);
DFFARX1 I_21200 (I362269,I1862,I361958,I361941,);
not I_21201 (I362300,I362125);
or I_21202 (I362317,I362091,I362300);
nor I_21203 (I361935,I362057,I362317);
nor I_21204 (I362348,I362026,I362300);
nand I_21205 (I361950,I362348,I362057);
not I_21206 (I362400,I1869);
and I_21207 (I362417,I260097,I260103);
nor I_21208 (I362434,I362417,I260091);
nand I_21209 (I362451,I260088,I260085);
nor I_21210 (I362468,I362451,I362434);
not I_21211 (I362389,I362468);
not I_21212 (I362499,I362451);
or I_21213 (I362516,I260094,I260106);
nor I_21214 (I362533,I362516,I260088);
nor I_21215 (I362550,I362533,I362499);
nand I_21216 (I362567,I260085,I260100);
nor I_21217 (I362584,I362567,I260091);
not I_21218 (I362601,I362584);
nor I_21219 (I362618,I362468,I362601);
nand I_21220 (I362386,I362618,I362533);
nor I_21221 (I362374,I362601,I362550);
nand I_21222 (I362380,I362533,I362601);
nor I_21223 (I362677,I362468,I362567);
nand I_21224 (I362694,I362677,I362533);
nand I_21225 (I362711,I362601,I362694);
DFFARX1 I_21226 (I362711,I1862,I362400,I362383,);
not I_21227 (I362742,I362567);
or I_21228 (I362759,I362533,I362742);
nor I_21229 (I362377,I362499,I362759);
nor I_21230 (I362790,I362468,I362742);
nand I_21231 (I362392,I362790,I362499);
not I_21232 (I362842,I1869);
and I_21233 (I362859,I1887,I1875);
nor I_21234 (I362876,I362859,I1893);
nand I_21235 (I362893,I1881,I1878);
nor I_21236 (I362910,I362893,I362876);
not I_21237 (I362831,I362910);
not I_21238 (I362941,I362893);
or I_21239 (I362958,I1875,I1872);
nor I_21240 (I362975,I362958,I1872);
nor I_21241 (I362992,I362975,I362941);
nand I_21242 (I363009,I1884,I1878);
nor I_21243 (I363026,I363009,I1890);
not I_21244 (I363043,I363026);
nor I_21245 (I363060,I362910,I363043);
nand I_21246 (I362828,I363060,I362975);
nor I_21247 (I362816,I363043,I362992);
nand I_21248 (I362822,I362975,I363043);
nor I_21249 (I363119,I362910,I363009);
nand I_21250 (I363136,I363119,I362975);
nand I_21251 (I363153,I363043,I363136);
DFFARX1 I_21252 (I363153,I1862,I362842,I362825,);
not I_21253 (I363184,I363009);
or I_21254 (I363201,I362975,I363184);
nor I_21255 (I362819,I362941,I363201);
nor I_21256 (I363232,I362910,I363184);
nand I_21257 (I362834,I363232,I362941);
not I_21258 (I363284,I1869);
and I_21259 (I363301,I194788,I194788);
nor I_21260 (I363318,I363301,I194812);
nand I_21261 (I363335,I194809,I194797);
nor I_21262 (I363352,I363335,I363318);
not I_21263 (I363273,I363352);
not I_21264 (I363383,I363335);
or I_21265 (I363400,I194791,I194791);
nor I_21266 (I363417,I363400,I194794);
nor I_21267 (I363434,I363417,I363383);
nand I_21268 (I363451,I194803,I194806);
nor I_21269 (I363468,I363451,I194800);
not I_21270 (I363485,I363468);
nor I_21271 (I363502,I363352,I363485);
nand I_21272 (I363270,I363502,I363417);
nor I_21273 (I363258,I363485,I363434);
nand I_21274 (I363264,I363417,I363485);
nor I_21275 (I363561,I363352,I363451);
nand I_21276 (I363578,I363561,I363417);
nand I_21277 (I363595,I363485,I363578);
DFFARX1 I_21278 (I363595,I1862,I363284,I363267,);
not I_21279 (I363626,I363451);
or I_21280 (I363643,I363417,I363626);
nor I_21281 (I363261,I363383,I363643);
nor I_21282 (I363674,I363352,I363626);
nand I_21283 (I363276,I363674,I363383);
not I_21284 (I363726,I1869);
and I_21285 (I363743,I347364,I347349);
nor I_21286 (I363760,I363743,I347352);
nand I_21287 (I363777,I347346,I347346);
nor I_21288 (I363794,I363777,I363760);
not I_21289 (I363715,I363794);
not I_21290 (I363825,I363777);
or I_21291 (I363842,I347349,I347367);
nor I_21292 (I363859,I363842,I347358);
nor I_21293 (I363876,I363859,I363825);
nand I_21294 (I363893,I347361,I347355);
nor I_21295 (I363910,I363893,I347352);
not I_21296 (I363927,I363910);
nor I_21297 (I363944,I363794,I363927);
nand I_21298 (I363712,I363944,I363859);
nor I_21299 (I363700,I363927,I363876);
nand I_21300 (I363706,I363859,I363927);
nor I_21301 (I364003,I363794,I363893);
nand I_21302 (I364020,I364003,I363859);
nand I_21303 (I364037,I363927,I364020);
DFFARX1 I_21304 (I364037,I1862,I363726,I363709,);
not I_21305 (I364068,I363893);
or I_21306 (I364085,I363859,I364068);
nor I_21307 (I363703,I363825,I364085);
nor I_21308 (I364116,I363794,I364068);
nand I_21309 (I363718,I364116,I363825);
not I_21310 (I364168,I1869);
and I_21311 (I364185,I16567,I16543);
nor I_21312 (I364202,I364185,I16549);
nand I_21313 (I364219,I16564,I16546);
nor I_21314 (I364236,I364219,I364202);
not I_21315 (I364157,I364236);
not I_21316 (I364267,I364219);
or I_21317 (I364284,I16543,I16546);
nor I_21318 (I364301,I364284,I16558);
nor I_21319 (I364318,I364301,I364267);
nand I_21320 (I364335,I16552,I16555);
nor I_21321 (I364352,I364335,I16561);
not I_21322 (I364369,I364352);
nor I_21323 (I364386,I364236,I364369);
nand I_21324 (I364154,I364386,I364301);
nor I_21325 (I364142,I364369,I364318);
nand I_21326 (I364148,I364301,I364369);
nor I_21327 (I364445,I364236,I364335);
nand I_21328 (I364462,I364445,I364301);
nand I_21329 (I364479,I364369,I364462);
DFFARX1 I_21330 (I364479,I1862,I364168,I364151,);
not I_21331 (I364510,I364335);
or I_21332 (I364527,I364301,I364510);
nor I_21333 (I364145,I364267,I364527);
nor I_21334 (I364558,I364236,I364510);
nand I_21335 (I364160,I364558,I364267);
not I_21336 (I364610,I1869);
and I_21337 (I364627,I288343,I288325);
nor I_21338 (I364644,I364627,I288340);
nand I_21339 (I364661,I288337,I288328);
nor I_21340 (I364678,I364661,I364644);
not I_21341 (I364599,I364678);
not I_21342 (I364709,I364661);
or I_21343 (I364726,I288322,I288328);
nor I_21344 (I364743,I364726,I288322);
nor I_21345 (I364760,I364743,I364709);
nand I_21346 (I364777,I288331,I288334);
nor I_21347 (I364794,I364777,I288325);
not I_21348 (I364811,I364794);
nor I_21349 (I364828,I364678,I364811);
nand I_21350 (I364596,I364828,I364743);
nor I_21351 (I364584,I364811,I364760);
nand I_21352 (I364590,I364743,I364811);
nor I_21353 (I364887,I364678,I364777);
nand I_21354 (I364904,I364887,I364743);
nand I_21355 (I364921,I364811,I364904);
DFFARX1 I_21356 (I364921,I1862,I364610,I364593,);
not I_21357 (I364952,I364777);
or I_21358 (I364969,I364743,I364952);
nor I_21359 (I364587,I364709,I364969);
nor I_21360 (I365000,I364678,I364952);
nand I_21361 (I364602,I365000,I364709);
not I_21362 (I365052,I1869);
and I_21363 (I365069,I245817,I245823);
nor I_21364 (I365086,I365069,I245811);
nand I_21365 (I365103,I245808,I245805);
nor I_21366 (I365120,I365103,I365086);
not I_21367 (I365041,I365120);
not I_21368 (I365151,I365103);
or I_21369 (I365168,I245814,I245826);
nor I_21370 (I365185,I365168,I245808);
nor I_21371 (I365202,I365185,I365151);
nand I_21372 (I365219,I245805,I245820);
nor I_21373 (I365236,I365219,I245811);
not I_21374 (I365253,I365236);
nor I_21375 (I365270,I365120,I365253);
nand I_21376 (I365038,I365270,I365185);
nor I_21377 (I365026,I365253,I365202);
nand I_21378 (I365032,I365185,I365253);
nor I_21379 (I365329,I365120,I365219);
nand I_21380 (I365346,I365329,I365185);
nand I_21381 (I365363,I365253,I365346);
DFFARX1 I_21382 (I365363,I1862,I365052,I365035,);
not I_21383 (I365394,I365219);
or I_21384 (I365411,I365185,I365394);
nor I_21385 (I365029,I365151,I365411);
nor I_21386 (I365442,I365120,I365394);
nand I_21387 (I365044,I365442,I365151);
not I_21388 (I365494,I1869);
and I_21389 (I365511,I283421,I283427);
nor I_21390 (I365528,I365511,I283415);
nand I_21391 (I365545,I283412,I283409);
nor I_21392 (I365562,I365545,I365528);
not I_21393 (I365483,I365562);
not I_21394 (I365593,I365545);
or I_21395 (I365610,I283418,I283430);
nor I_21396 (I365627,I365610,I283412);
nor I_21397 (I365644,I365627,I365593);
nand I_21398 (I365661,I283409,I283424);
nor I_21399 (I365678,I365661,I283415);
not I_21400 (I365695,I365678);
nor I_21401 (I365712,I365562,I365695);
nand I_21402 (I365480,I365712,I365627);
nor I_21403 (I365468,I365695,I365644);
nand I_21404 (I365474,I365627,I365695);
nor I_21405 (I365771,I365562,I365661);
nand I_21406 (I365788,I365771,I365627);
nand I_21407 (I365805,I365695,I365788);
DFFARX1 I_21408 (I365805,I1862,I365494,I365477,);
not I_21409 (I365836,I365661);
or I_21410 (I365853,I365627,I365836);
nor I_21411 (I365471,I365593,I365853);
nor I_21412 (I365884,I365562,I365836);
nand I_21413 (I365486,I365884,I365593);
not I_21414 (I365936,I1869);
and I_21415 (I365953,I136818,I136818);
nor I_21416 (I365970,I365953,I136842);
nand I_21417 (I365987,I136839,I136827);
nor I_21418 (I366004,I365987,I365970);
not I_21419 (I365925,I366004);
not I_21420 (I366035,I365987);
or I_21421 (I366052,I136821,I136821);
nor I_21422 (I366069,I366052,I136824);
nor I_21423 (I366086,I366069,I366035);
nand I_21424 (I366103,I136833,I136836);
nor I_21425 (I366120,I366103,I136830);
not I_21426 (I366137,I366120);
nor I_21427 (I366154,I366004,I366137);
nand I_21428 (I365922,I366154,I366069);
nor I_21429 (I365910,I366137,I366086);
nand I_21430 (I365916,I366069,I366137);
nor I_21431 (I366213,I366004,I366103);
nand I_21432 (I366230,I366213,I366069);
nand I_21433 (I366247,I366137,I366230);
DFFARX1 I_21434 (I366247,I1862,I365936,I365919,);
not I_21435 (I366278,I366103);
or I_21436 (I366295,I366069,I366278);
nor I_21437 (I365913,I366035,I366295);
nor I_21438 (I366326,I366004,I366278);
nand I_21439 (I365928,I366326,I366035);
not I_21440 (I366378,I1869);
and I_21441 (I366395,I133656,I133656);
nor I_21442 (I366412,I366395,I133680);
nand I_21443 (I366429,I133677,I133665);
nor I_21444 (I366446,I366429,I366412);
not I_21445 (I366367,I366446);
not I_21446 (I366477,I366429);
or I_21447 (I366494,I133659,I133659);
nor I_21448 (I366511,I366494,I133662);
nor I_21449 (I366528,I366511,I366477);
nand I_21450 (I366545,I133671,I133674);
nor I_21451 (I366562,I366545,I133668);
not I_21452 (I366579,I366562);
nor I_21453 (I366596,I366446,I366579);
nand I_21454 (I366364,I366596,I366511);
nor I_21455 (I366352,I366579,I366528);
nand I_21456 (I366358,I366511,I366579);
nor I_21457 (I366655,I366446,I366545);
nand I_21458 (I366672,I366655,I366511);
nand I_21459 (I366689,I366579,I366672);
DFFARX1 I_21460 (I366689,I1862,I366378,I366361,);
not I_21461 (I366720,I366545);
or I_21462 (I366737,I366511,I366720);
nor I_21463 (I366355,I366477,I366737);
nor I_21464 (I366768,I366446,I366720);
nand I_21465 (I366370,I366768,I366477);
not I_21466 (I366820,I1869);
and I_21467 (I366837,I17587,I17563);
nor I_21468 (I366854,I366837,I17569);
nand I_21469 (I366871,I17584,I17566);
nor I_21470 (I366888,I366871,I366854);
not I_21471 (I366809,I366888);
not I_21472 (I366919,I366871);
or I_21473 (I366936,I17563,I17566);
nor I_21474 (I366953,I366936,I17578);
nor I_21475 (I366970,I366953,I366919);
nand I_21476 (I366987,I17572,I17575);
nor I_21477 (I367004,I366987,I17581);
not I_21478 (I367021,I367004);
nor I_21479 (I367038,I366888,I367021);
nand I_21480 (I366806,I367038,I366953);
nor I_21481 (I366794,I367021,I366970);
nand I_21482 (I366800,I366953,I367021);
nor I_21483 (I367097,I366888,I366987);
nand I_21484 (I367114,I367097,I366953);
nand I_21485 (I367131,I367021,I367114);
DFFARX1 I_21486 (I367131,I1862,I366820,I366803,);
not I_21487 (I367162,I366987);
or I_21488 (I367179,I366953,I367162);
nor I_21489 (I366797,I366919,I367179);
nor I_21490 (I367210,I366888,I367162);
nand I_21491 (I366812,I367210,I366919);
not I_21492 (I367262,I1869);
and I_21493 (I367279,I154736,I154736);
nor I_21494 (I367296,I367279,I154760);
nand I_21495 (I367313,I154757,I154745);
nor I_21496 (I367330,I367313,I367296);
not I_21497 (I367251,I367330);
not I_21498 (I367361,I367313);
or I_21499 (I367378,I154739,I154739);
nor I_21500 (I367395,I367378,I154742);
nor I_21501 (I367412,I367395,I367361);
nand I_21502 (I367429,I154751,I154754);
nor I_21503 (I367446,I367429,I154748);
not I_21504 (I367463,I367446);
nor I_21505 (I367480,I367330,I367463);
nand I_21506 (I367248,I367480,I367395);
nor I_21507 (I367236,I367463,I367412);
nand I_21508 (I367242,I367395,I367463);
nor I_21509 (I367539,I367330,I367429);
nand I_21510 (I367556,I367539,I367395);
nand I_21511 (I367573,I367463,I367556);
DFFARX1 I_21512 (I367573,I1862,I367262,I367245,);
not I_21513 (I367604,I367429);
or I_21514 (I367621,I367395,I367604);
nor I_21515 (I367239,I367361,I367621);
nor I_21516 (I367652,I367330,I367604);
nand I_21517 (I367254,I367652,I367361);
not I_21518 (I367704,I1869);
and I_21519 (I367721,I110383,I110389);
nor I_21520 (I367738,I367721,I110389);
nand I_21521 (I367755,I110392,I110398);
nor I_21522 (I367772,I367755,I367738);
not I_21523 (I367693,I367772);
not I_21524 (I367803,I367755);
or I_21525 (I367820,I110386,I110386);
nor I_21526 (I367837,I367820,I110401);
nor I_21527 (I367854,I367837,I367803);
nand I_21528 (I367871,I110395,I110383);
nor I_21529 (I367888,I367871,I110392);
not I_21530 (I367905,I367888);
nor I_21531 (I367922,I367772,I367905);
nand I_21532 (I367690,I367922,I367837);
nor I_21533 (I367678,I367905,I367854);
nand I_21534 (I367684,I367837,I367905);
nor I_21535 (I367981,I367772,I367871);
nand I_21536 (I367998,I367981,I367837);
nand I_21537 (I368015,I367905,I367998);
DFFARX1 I_21538 (I368015,I1862,I367704,I367687,);
not I_21539 (I368046,I367871);
or I_21540 (I368063,I367837,I368046);
nor I_21541 (I367681,I367803,I368063);
nor I_21542 (I368094,I367772,I368046);
nand I_21543 (I367696,I368094,I367803);
not I_21544 (I368146,I1869);
and I_21545 (I368163,I262953,I262959);
nor I_21546 (I368180,I368163,I262947);
nand I_21547 (I368197,I262944,I262941);
nor I_21548 (I368214,I368197,I368180);
not I_21549 (I368135,I368214);
not I_21550 (I368245,I368197);
or I_21551 (I368262,I262950,I262962);
nor I_21552 (I368279,I368262,I262944);
nor I_21553 (I368296,I368279,I368245);
nand I_21554 (I368313,I262941,I262956);
nor I_21555 (I368330,I368313,I262947);
not I_21556 (I368347,I368330);
nor I_21557 (I368364,I368214,I368347);
nand I_21558 (I368132,I368364,I368279);
nor I_21559 (I368120,I368347,I368296);
nand I_21560 (I368126,I368279,I368347);
nor I_21561 (I368423,I368214,I368313);
nand I_21562 (I368440,I368423,I368279);
nand I_21563 (I368457,I368347,I368440);
DFFARX1 I_21564 (I368457,I1862,I368146,I368129,);
not I_21565 (I368488,I368313);
or I_21566 (I368505,I368279,I368488);
nor I_21567 (I368123,I368245,I368505);
nor I_21568 (I368536,I368214,I368488);
nand I_21569 (I368138,I368536,I368245);
not I_21570 (I368588,I1869);
and I_21571 (I368605,I58897,I58873);
nor I_21572 (I368622,I368605,I58879);
nand I_21573 (I368639,I58894,I58876);
nor I_21574 (I368656,I368639,I368622);
not I_21575 (I368577,I368656);
not I_21576 (I368687,I368639);
or I_21577 (I368704,I58873,I58876);
nor I_21578 (I368721,I368704,I58888);
nor I_21579 (I368738,I368721,I368687);
nand I_21580 (I368755,I58882,I58885);
nor I_21581 (I368772,I368755,I58891);
not I_21582 (I368789,I368772);
nor I_21583 (I368806,I368656,I368789);
nand I_21584 (I368574,I368806,I368721);
nor I_21585 (I368562,I368789,I368738);
nand I_21586 (I368568,I368721,I368789);
nor I_21587 (I368865,I368656,I368755);
nand I_21588 (I368882,I368865,I368721);
nand I_21589 (I368899,I368789,I368882);
DFFARX1 I_21590 (I368899,I1862,I368588,I368571,);
not I_21591 (I368930,I368755);
or I_21592 (I368947,I368721,I368930);
nor I_21593 (I368565,I368687,I368947);
nor I_21594 (I368978,I368656,I368930);
nand I_21595 (I368580,I368978,I368687);
not I_21596 (I369030,I1869);
and I_21597 (I369047,I330500,I330485);
nor I_21598 (I369064,I369047,I330488);
nand I_21599 (I369081,I330482,I330482);
nor I_21600 (I369098,I369081,I369064);
not I_21601 (I369019,I369098);
not I_21602 (I369129,I369081);
or I_21603 (I369146,I330485,I330503);
nor I_21604 (I369163,I369146,I330494);
nor I_21605 (I369180,I369163,I369129);
nand I_21606 (I369197,I330497,I330491);
nor I_21607 (I369214,I369197,I330488);
not I_21608 (I369231,I369214);
nor I_21609 (I369248,I369098,I369231);
nand I_21610 (I369016,I369248,I369163);
nor I_21611 (I369004,I369231,I369180);
nand I_21612 (I369010,I369163,I369231);
nor I_21613 (I369307,I369098,I369197);
nand I_21614 (I369324,I369307,I369163);
nand I_21615 (I369341,I369231,I369324);
DFFARX1 I_21616 (I369341,I1862,I369030,I369013,);
not I_21617 (I369372,I369197);
or I_21618 (I369389,I369163,I369372);
nor I_21619 (I369007,I369129,I369389);
nor I_21620 (I369420,I369098,I369372);
nand I_21621 (I369022,I369420,I369129);
not I_21622 (I369472,I1869);
and I_21623 (I369489,I312582,I312567);
nor I_21624 (I369506,I369489,I312570);
nand I_21625 (I369523,I312564,I312564);
nor I_21626 (I369540,I369523,I369506);
not I_21627 (I369461,I369540);
not I_21628 (I369571,I369523);
or I_21629 (I369588,I312567,I312585);
nor I_21630 (I369605,I369588,I312576);
nor I_21631 (I369622,I369605,I369571);
nand I_21632 (I369639,I312579,I312573);
nor I_21633 (I369656,I369639,I312570);
not I_21634 (I369673,I369656);
nor I_21635 (I369690,I369540,I369673);
nand I_21636 (I369458,I369690,I369605);
nor I_21637 (I369446,I369673,I369622);
nand I_21638 (I369452,I369605,I369673);
nor I_21639 (I369749,I369540,I369639);
nand I_21640 (I369766,I369749,I369605);
nand I_21641 (I369783,I369673,I369766);
DFFARX1 I_21642 (I369783,I1862,I369472,I369455,);
not I_21643 (I369814,I369639);
or I_21644 (I369831,I369605,I369814);
nor I_21645 (I369449,I369571,I369831);
nor I_21646 (I369862,I369540,I369814);
nand I_21647 (I369464,I369862,I369571);
not I_21648 (I369914,I1869);
and I_21649 (I369931,I152101,I152101);
nor I_21650 (I369948,I369931,I152125);
nand I_21651 (I369965,I152122,I152110);
nor I_21652 (I369982,I369965,I369948);
not I_21653 (I369903,I369982);
not I_21654 (I370013,I369965);
or I_21655 (I370030,I152104,I152104);
nor I_21656 (I370047,I370030,I152107);
nor I_21657 (I370064,I370047,I370013);
nand I_21658 (I370081,I152116,I152119);
nor I_21659 (I370098,I370081,I152113);
not I_21660 (I370115,I370098);
nor I_21661 (I370132,I369982,I370115);
nand I_21662 (I369900,I370132,I370047);
nor I_21663 (I369888,I370115,I370064);
nand I_21664 (I369894,I370047,I370115);
nor I_21665 (I370191,I369982,I370081);
nand I_21666 (I370208,I370191,I370047);
nand I_21667 (I370225,I370115,I370208);
DFFARX1 I_21668 (I370225,I1862,I369914,I369897,);
not I_21669 (I370256,I370081);
or I_21670 (I370273,I370047,I370256);
nor I_21671 (I369891,I370013,I370273);
nor I_21672 (I370304,I369982,I370256);
nand I_21673 (I369906,I370304,I370013);
not I_21674 (I370356,I1869);
and I_21675 (I370373,I172127,I172127);
nor I_21676 (I370390,I370373,I172151);
nand I_21677 (I370407,I172148,I172136);
nor I_21678 (I370424,I370407,I370390);
not I_21679 (I370345,I370424);
not I_21680 (I370455,I370407);
or I_21681 (I370472,I172130,I172130);
nor I_21682 (I370489,I370472,I172133);
nor I_21683 (I370506,I370489,I370455);
nand I_21684 (I370523,I172142,I172145);
nor I_21685 (I370540,I370523,I172139);
not I_21686 (I370557,I370540);
nor I_21687 (I370574,I370424,I370557);
nand I_21688 (I370342,I370574,I370489);
nor I_21689 (I370330,I370557,I370506);
nand I_21690 (I370336,I370489,I370557);
nor I_21691 (I370633,I370424,I370523);
nand I_21692 (I370650,I370633,I370489);
nand I_21693 (I370667,I370557,I370650);
DFFARX1 I_21694 (I370667,I1862,I370356,I370339,);
not I_21695 (I370698,I370523);
or I_21696 (I370715,I370489,I370698);
nor I_21697 (I370333,I370455,I370715);
nor I_21698 (I370746,I370424,I370698);
nand I_21699 (I370348,I370746,I370455);
not I_21700 (I370798,I1869);
and I_21701 (I370815,I253433,I253439);
nor I_21702 (I370832,I370815,I253427);
nand I_21703 (I370849,I253424,I253421);
nor I_21704 (I370866,I370849,I370832);
not I_21705 (I370787,I370866);
not I_21706 (I370897,I370849);
or I_21707 (I370914,I253430,I253442);
nor I_21708 (I370931,I370914,I253424);
nor I_21709 (I370948,I370931,I370897);
nand I_21710 (I370965,I253421,I253436);
nor I_21711 (I370982,I370965,I253427);
not I_21712 (I370999,I370982);
nor I_21713 (I371016,I370866,I370999);
nand I_21714 (I370784,I371016,I370931);
nor I_21715 (I370772,I370999,I370948);
nand I_21716 (I370778,I370931,I370999);
nor I_21717 (I371075,I370866,I370965);
nand I_21718 (I371092,I371075,I370931);
nand I_21719 (I371109,I370999,I371092);
DFFARX1 I_21720 (I371109,I1862,I370798,I370781,);
not I_21721 (I371140,I370965);
or I_21722 (I371157,I370931,I371140);
nor I_21723 (I370775,I370897,I371157);
nor I_21724 (I371188,I370866,I371140);
nand I_21725 (I370790,I371188,I370897);
not I_21726 (I371240,I1869);
and I_21727 (I371257,I341567,I341552);
nor I_21728 (I371274,I371257,I341555);
nand I_21729 (I371291,I341549,I341549);
nor I_21730 (I371308,I371291,I371274);
not I_21731 (I371229,I371308);
not I_21732 (I371339,I371291);
or I_21733 (I371356,I341552,I341570);
nor I_21734 (I371373,I371356,I341561);
nor I_21735 (I371390,I371373,I371339);
nand I_21736 (I371407,I341564,I341558);
nor I_21737 (I371424,I371407,I341555);
not I_21738 (I371441,I371424);
nor I_21739 (I371458,I371308,I371441);
nand I_21740 (I371226,I371458,I371373);
nor I_21741 (I371214,I371441,I371390);
nand I_21742 (I371220,I371373,I371441);
nor I_21743 (I371517,I371308,I371407);
nand I_21744 (I371534,I371517,I371373);
nand I_21745 (I371551,I371441,I371534);
DFFARX1 I_21746 (I371551,I1862,I371240,I371223,);
not I_21747 (I371582,I371407);
or I_21748 (I371599,I371373,I371582);
nor I_21749 (I371217,I371339,I371599);
nor I_21750 (I371630,I371308,I371582);
nand I_21751 (I371232,I371630,I371339);
not I_21752 (I371682,I1869);
and I_21753 (I371699,I154209,I154209);
nor I_21754 (I371716,I371699,I154233);
nand I_21755 (I371733,I154230,I154218);
nor I_21756 (I371750,I371733,I371716);
not I_21757 (I371671,I371750);
not I_21758 (I371781,I371733);
or I_21759 (I371798,I154212,I154212);
nor I_21760 (I371815,I371798,I154215);
nor I_21761 (I371832,I371815,I371781);
nand I_21762 (I371849,I154224,I154227);
nor I_21763 (I371866,I371849,I154221);
not I_21764 (I371883,I371866);
nor I_21765 (I371900,I371750,I371883);
nand I_21766 (I371668,I371900,I371815);
nor I_21767 (I371656,I371883,I371832);
nand I_21768 (I371662,I371815,I371883);
nor I_21769 (I371959,I371750,I371849);
nand I_21770 (I371976,I371959,I371815);
nand I_21771 (I371993,I371883,I371976);
DFFARX1 I_21772 (I371993,I1862,I371682,I371665,);
not I_21773 (I372024,I371849);
or I_21774 (I372041,I371815,I372024);
nor I_21775 (I371659,I371781,I372041);
nor I_21776 (I372072,I371750,I372024);
nand I_21777 (I371674,I372072,I371781);
not I_21778 (I372124,I1869);
and I_21779 (I372141,I323122,I323107);
nor I_21780 (I372158,I372141,I323110);
nand I_21781 (I372175,I323104,I323104);
nor I_21782 (I372192,I372175,I372158);
not I_21783 (I372113,I372192);
not I_21784 (I372223,I372175);
or I_21785 (I372240,I323107,I323125);
nor I_21786 (I372257,I372240,I323116);
nor I_21787 (I372274,I372257,I372223);
nand I_21788 (I372291,I323119,I323113);
nor I_21789 (I372308,I372291,I323110);
not I_21790 (I372325,I372308);
nor I_21791 (I372342,I372192,I372325);
nand I_21792 (I372110,I372342,I372257);
nor I_21793 (I372098,I372325,I372274);
nand I_21794 (I372104,I372257,I372325);
nor I_21795 (I372401,I372192,I372291);
nand I_21796 (I372418,I372401,I372257);
nand I_21797 (I372435,I372325,I372418);
DFFARX1 I_21798 (I372435,I1862,I372124,I372107,);
not I_21799 (I372466,I372291);
or I_21800 (I372483,I372257,I372466);
nor I_21801 (I372101,I372223,I372483);
nor I_21802 (I372514,I372192,I372466);
nand I_21803 (I372116,I372514,I372223);
not I_21804 (I372566,I1869);
and I_21805 (I372583,I226777,I226783);
nor I_21806 (I372600,I372583,I226771);
nand I_21807 (I372617,I226768,I226765);
nor I_21808 (I372634,I372617,I372600);
not I_21809 (I372555,I372634);
not I_21810 (I372665,I372617);
or I_21811 (I372682,I226774,I226786);
nor I_21812 (I372699,I372682,I226768);
nor I_21813 (I372716,I372699,I372665);
nand I_21814 (I372733,I226765,I226780);
nor I_21815 (I372750,I372733,I226771);
not I_21816 (I372767,I372750);
nor I_21817 (I372784,I372634,I372767);
nand I_21818 (I372552,I372784,I372699);
nor I_21819 (I372540,I372767,I372716);
nand I_21820 (I372546,I372699,I372767);
nor I_21821 (I372843,I372634,I372733);
nand I_21822 (I372860,I372843,I372699);
nand I_21823 (I372877,I372767,I372860);
DFFARX1 I_21824 (I372877,I1862,I372566,I372549,);
not I_21825 (I372908,I372733);
or I_21826 (I372925,I372699,I372908);
nor I_21827 (I372543,I372665,I372925);
nor I_21828 (I372956,I372634,I372908);
nand I_21829 (I372558,I372956,I372665);
not I_21830 (I373008,I1869);
and I_21831 (I373025,I975,I1751);
nor I_21832 (I373042,I373025,I1039);
nand I_21833 (I373059,I1103,I1399);
nor I_21834 (I373076,I373059,I373042);
not I_21835 (I372997,I373076);
not I_21836 (I373107,I373059);
or I_21837 (I373124,I911,I1695);
nor I_21838 (I373141,I373124,I847);
nor I_21839 (I373158,I373141,I373107);
nand I_21840 (I373175,I1023,I951);
nor I_21841 (I373192,I373175,I1367);
not I_21842 (I373209,I373192);
nor I_21843 (I373226,I373076,I373209);
nand I_21844 (I372994,I373226,I373141);
nor I_21845 (I372982,I373209,I373158);
nand I_21846 (I372988,I373141,I373209);
nor I_21847 (I373285,I373076,I373175);
nand I_21848 (I373302,I373285,I373141);
nand I_21849 (I373319,I373209,I373302);
DFFARX1 I_21850 (I373319,I1862,I373008,I372991,);
not I_21851 (I373350,I373175);
or I_21852 (I373367,I373141,I373350);
nor I_21853 (I372985,I373107,I373367);
nor I_21854 (I373398,I373076,I373350);
nand I_21855 (I373000,I373398,I373107);
not I_21856 (I373450,I1869);
and I_21857 (I373467,I92557,I92533);
nor I_21858 (I373484,I373467,I92539);
nand I_21859 (I373501,I92554,I92536);
nor I_21860 (I373518,I373501,I373484);
not I_21861 (I373439,I373518);
not I_21862 (I373549,I373501);
or I_21863 (I373566,I92533,I92536);
nor I_21864 (I373583,I373566,I92548);
nor I_21865 (I373600,I373583,I373549);
nand I_21866 (I373617,I92542,I92545);
nor I_21867 (I373634,I373617,I92551);
not I_21868 (I373651,I373634);
nor I_21869 (I373668,I373518,I373651);
nand I_21870 (I373436,I373668,I373583);
nor I_21871 (I373424,I373651,I373600);
nand I_21872 (I373430,I373583,I373651);
nor I_21873 (I373727,I373518,I373617);
nand I_21874 (I373744,I373727,I373583);
nand I_21875 (I373761,I373651,I373744);
DFFARX1 I_21876 (I373761,I1862,I373450,I373433,);
not I_21877 (I373792,I373617);
or I_21878 (I373809,I373583,I373792);
nor I_21879 (I373427,I373549,I373809);
nor I_21880 (I373840,I373518,I373792);
nand I_21881 (I373442,I373840,I373549);
not I_21882 (I373892,I1869);
and I_21883 (I373909,I193734,I193734);
nor I_21884 (I373926,I373909,I193758);
nand I_21885 (I373943,I193755,I193743);
nor I_21886 (I373960,I373943,I373926);
not I_21887 (I373881,I373960);
not I_21888 (I373991,I373943);
or I_21889 (I374008,I193737,I193737);
nor I_21890 (I374025,I374008,I193740);
nor I_21891 (I374042,I374025,I373991);
nand I_21892 (I374059,I193749,I193752);
nor I_21893 (I374076,I374059,I193746);
not I_21894 (I374093,I374076);
nor I_21895 (I374110,I373960,I374093);
nand I_21896 (I373878,I374110,I374025);
nor I_21897 (I373866,I374093,I374042);
nand I_21898 (I373872,I374025,I374093);
nor I_21899 (I374169,I373960,I374059);
nand I_21900 (I374186,I374169,I374025);
nand I_21901 (I374203,I374093,I374186);
DFFARX1 I_21902 (I374203,I1862,I373892,I373875,);
not I_21903 (I374234,I374059);
or I_21904 (I374251,I374025,I374234);
nor I_21905 (I373869,I373991,I374251);
nor I_21906 (I374282,I373960,I374234);
nand I_21907 (I373884,I374282,I373991);
not I_21908 (I374334,I1869);
and I_21909 (I374351,I296248,I296230);
nor I_21910 (I374368,I374351,I296245);
nand I_21911 (I374385,I296242,I296233);
nor I_21912 (I374402,I374385,I374368);
not I_21913 (I374323,I374402);
not I_21914 (I374433,I374385);
or I_21915 (I374450,I296227,I296233);
nor I_21916 (I374467,I374450,I296227);
nor I_21917 (I374484,I374467,I374433);
nand I_21918 (I374501,I296236,I296239);
nor I_21919 (I374518,I374501,I296230);
not I_21920 (I374535,I374518);
nor I_21921 (I374552,I374402,I374535);
nand I_21922 (I374320,I374552,I374467);
nor I_21923 (I374308,I374535,I374484);
nand I_21924 (I374314,I374467,I374535);
nor I_21925 (I374611,I374402,I374501);
nand I_21926 (I374628,I374611,I374467);
nand I_21927 (I374645,I374535,I374628);
DFFARX1 I_21928 (I374645,I1862,I374334,I374317,);
not I_21929 (I374676,I374501);
or I_21930 (I374693,I374467,I374676);
nor I_21931 (I374311,I374433,I374693);
nor I_21932 (I374724,I374402,I374676);
nand I_21933 (I374326,I374724,I374433);
not I_21934 (I374776,I1869);
and I_21935 (I374793,I167911,I167911);
nor I_21936 (I374810,I374793,I167935);
nand I_21937 (I374827,I167932,I167920);
nor I_21938 (I374844,I374827,I374810);
not I_21939 (I374765,I374844);
not I_21940 (I374875,I374827);
or I_21941 (I374892,I167914,I167914);
nor I_21942 (I374909,I374892,I167917);
nor I_21943 (I374926,I374909,I374875);
nand I_21944 (I374943,I167926,I167929);
nor I_21945 (I374960,I374943,I167923);
not I_21946 (I374977,I374960);
nor I_21947 (I374994,I374844,I374977);
nand I_21948 (I374762,I374994,I374909);
nor I_21949 (I374750,I374977,I374926);
nand I_21950 (I374756,I374909,I374977);
nor I_21951 (I375053,I374844,I374943);
nand I_21952 (I375070,I375053,I374909);
nand I_21953 (I375087,I374977,I375070);
DFFARX1 I_21954 (I375087,I1862,I374776,I374759,);
not I_21955 (I375118,I374943);
or I_21956 (I375135,I374909,I375118);
nor I_21957 (I374753,I374875,I375135);
nor I_21958 (I375166,I374844,I375118);
nand I_21959 (I374768,I375166,I374875);
not I_21960 (I375218,I1869);
and I_21961 (I375235,I234393,I234399);
nor I_21962 (I375252,I375235,I234387);
nand I_21963 (I375269,I234384,I234381);
nor I_21964 (I375286,I375269,I375252);
not I_21965 (I375207,I375286);
not I_21966 (I375317,I375269);
or I_21967 (I375334,I234390,I234402);
nor I_21968 (I375351,I375334,I234384);
nor I_21969 (I375368,I375351,I375317);
nand I_21970 (I375385,I234381,I234396);
nor I_21971 (I375402,I375385,I234387);
not I_21972 (I375419,I375402);
nor I_21973 (I375436,I375286,I375419);
nand I_21974 (I375204,I375436,I375351);
nor I_21975 (I375192,I375419,I375368);
nand I_21976 (I375198,I375351,I375419);
nor I_21977 (I375495,I375286,I375385);
nand I_21978 (I375512,I375495,I375351);
nand I_21979 (I375529,I375419,I375512);
DFFARX1 I_21980 (I375529,I1862,I375218,I375201,);
not I_21981 (I375560,I375385);
or I_21982 (I375577,I375351,I375560);
nor I_21983 (I375195,I375317,I375577);
nor I_21984 (I375608,I375286,I375560);
nand I_21985 (I375210,I375608,I375317);
not I_21986 (I375660,I1869);
and I_21987 (I375677,I213925,I213931);
nor I_21988 (I375694,I375677,I213919);
nand I_21989 (I375711,I213916,I213913);
nor I_21990 (I375728,I375711,I375694);
not I_21991 (I375649,I375728);
not I_21992 (I375759,I375711);
or I_21993 (I375776,I213922,I213934);
nor I_21994 (I375793,I375776,I213916);
nor I_21995 (I375810,I375793,I375759);
nand I_21996 (I375827,I213913,I213928);
nor I_21997 (I375844,I375827,I213919);
not I_21998 (I375861,I375844);
nor I_21999 (I375878,I375728,I375861);
nand I_22000 (I375646,I375878,I375793);
nor I_22001 (I375634,I375861,I375810);
nand I_22002 (I375640,I375793,I375861);
nor I_22003 (I375937,I375728,I375827);
nand I_22004 (I375954,I375937,I375793);
nand I_22005 (I375971,I375861,I375954);
DFFARX1 I_22006 (I375971,I1862,I375660,I375643,);
not I_22007 (I376002,I375827);
or I_22008 (I376019,I375793,I376002);
nor I_22009 (I375637,I375759,I376019);
nor I_22010 (I376050,I375728,I376002);
nand I_22011 (I375652,I376050,I375759);
not I_22012 (I376102,I1869);
and I_22013 (I376119,I74197,I74173);
nor I_22014 (I376136,I376119,I74179);
nand I_22015 (I376153,I74194,I74176);
nor I_22016 (I376170,I376153,I376136);
not I_22017 (I376091,I376170);
not I_22018 (I376201,I376153);
or I_22019 (I376218,I74173,I74176);
nor I_22020 (I376235,I376218,I74188);
nor I_22021 (I376252,I376235,I376201);
nand I_22022 (I376269,I74182,I74185);
nor I_22023 (I376286,I376269,I74191);
not I_22024 (I376303,I376286);
nor I_22025 (I376320,I376170,I376303);
nand I_22026 (I376088,I376320,I376235);
nor I_22027 (I376076,I376303,I376252);
nand I_22028 (I376082,I376235,I376303);
nor I_22029 (I376379,I376170,I376269);
nand I_22030 (I376396,I376379,I376235);
nand I_22031 (I376413,I376303,I376396);
DFFARX1 I_22032 (I376413,I1862,I376102,I376085,);
not I_22033 (I376444,I376269);
or I_22034 (I376461,I376235,I376444);
nor I_22035 (I376079,I376201,I376461);
nor I_22036 (I376492,I376170,I376444);
nand I_22037 (I376094,I376492,I376201);
not I_22038 (I376544,I1869);
and I_22039 (I376561,I210117,I210123);
nor I_22040 (I376578,I376561,I210111);
nand I_22041 (I376595,I210108,I210105);
nor I_22042 (I376612,I376595,I376578);
not I_22043 (I376533,I376612);
not I_22044 (I376643,I376595);
or I_22045 (I376660,I210114,I210126);
nor I_22046 (I376677,I376660,I210108);
nor I_22047 (I376694,I376677,I376643);
nand I_22048 (I376711,I210105,I210120);
nor I_22049 (I376728,I376711,I210111);
not I_22050 (I376745,I376728);
nor I_22051 (I376762,I376612,I376745);
nand I_22052 (I376530,I376762,I376677);
nor I_22053 (I376518,I376745,I376694);
nand I_22054 (I376524,I376677,I376745);
nor I_22055 (I376821,I376612,I376711);
nand I_22056 (I376838,I376821,I376677);
nand I_22057 (I376855,I376745,I376838);
DFFARX1 I_22058 (I376855,I1862,I376544,I376527,);
not I_22059 (I376886,I376711);
or I_22060 (I376903,I376677,I376886);
nor I_22061 (I376521,I376643,I376903);
nor I_22062 (I376934,I376612,I376886);
nand I_22063 (I376536,I376934,I376643);
not I_22064 (I376986,I1869);
and I_22065 (I377003,I151574,I151574);
nor I_22066 (I377020,I377003,I151598);
nand I_22067 (I377037,I151595,I151583);
nor I_22068 (I377054,I377037,I377020);
not I_22069 (I376975,I377054);
not I_22070 (I377085,I377037);
or I_22071 (I377102,I151577,I151577);
nor I_22072 (I377119,I377102,I151580);
nor I_22073 (I377136,I377119,I377085);
nand I_22074 (I377153,I151589,I151592);
nor I_22075 (I377170,I377153,I151586);
not I_22076 (I377187,I377170);
nor I_22077 (I377204,I377054,I377187);
nand I_22078 (I376972,I377204,I377119);
nor I_22079 (I376960,I377187,I377136);
nand I_22080 (I376966,I377119,I377187);
nor I_22081 (I377263,I377054,I377153);
nand I_22082 (I377280,I377263,I377119);
nand I_22083 (I377297,I377187,I377280);
DFFARX1 I_22084 (I377297,I1862,I376986,I376969,);
not I_22085 (I377328,I377153);
or I_22086 (I377345,I377119,I377328);
nor I_22087 (I376963,I377085,I377345);
nor I_22088 (I377376,I377054,I377328);
nand I_22089 (I376978,I377376,I377085);
not I_22090 (I377428,I1869);
and I_22091 (I377445,I342094,I342079);
nor I_22092 (I377462,I377445,I342082);
nand I_22093 (I377479,I342076,I342076);
nor I_22094 (I377496,I377479,I377462);
not I_22095 (I377417,I377496);
not I_22096 (I377527,I377479);
or I_22097 (I377544,I342079,I342097);
nor I_22098 (I377561,I377544,I342088);
nor I_22099 (I377578,I377561,I377527);
nand I_22100 (I377595,I342091,I342085);
nor I_22101 (I377612,I377595,I342082);
not I_22102 (I377629,I377612);
nor I_22103 (I377646,I377496,I377629);
nand I_22104 (I377414,I377646,I377561);
nor I_22105 (I377402,I377629,I377578);
nand I_22106 (I377408,I377561,I377629);
nor I_22107 (I377705,I377496,I377595);
nand I_22108 (I377722,I377705,I377561);
nand I_22109 (I377739,I377629,I377722);
DFFARX1 I_22110 (I377739,I1862,I377428,I377411,);
not I_22111 (I377770,I377595);
or I_22112 (I377787,I377561,I377770);
nor I_22113 (I377405,I377527,I377787);
nor I_22114 (I377818,I377496,I377770);
nand I_22115 (I377420,I377818,I377527);
not I_22116 (I377870,I1869);
and I_22117 (I377887,I61447,I61423);
nor I_22118 (I377904,I377887,I61429);
nand I_22119 (I377921,I61444,I61426);
nor I_22120 (I377938,I377921,I377904);
not I_22121 (I377859,I377938);
not I_22122 (I377969,I377921);
or I_22123 (I377986,I61423,I61426);
nor I_22124 (I378003,I377986,I61438);
nor I_22125 (I378020,I378003,I377969);
nand I_22126 (I378037,I61432,I61435);
nor I_22127 (I378054,I378037,I61441);
not I_22128 (I378071,I378054);
nor I_22129 (I378088,I377938,I378071);
nand I_22130 (I377856,I378088,I378003);
nor I_22131 (I377844,I378071,I378020);
nand I_22132 (I377850,I378003,I378071);
nor I_22133 (I378147,I377938,I378037);
nand I_22134 (I378164,I378147,I378003);
nand I_22135 (I378181,I378071,I378164);
DFFARX1 I_22136 (I378181,I1862,I377870,I377853,);
not I_22137 (I378212,I378037);
or I_22138 (I378229,I378003,I378212);
nor I_22139 (I377847,I377969,I378229);
nor I_22140 (I378260,I377938,I378212);
nand I_22141 (I377862,I378260,I377969);
not I_22142 (I378312,I1869);
and I_22143 (I378329,I116911,I116917);
nor I_22144 (I378346,I378329,I116917);
nand I_22145 (I378363,I116920,I116926);
nor I_22146 (I378380,I378363,I378346);
not I_22147 (I378301,I378380);
not I_22148 (I378411,I378363);
or I_22149 (I378428,I116914,I116914);
nor I_22150 (I378445,I378428,I116929);
nor I_22151 (I378462,I378445,I378411);
nand I_22152 (I378479,I116923,I116911);
nor I_22153 (I378496,I378479,I116920);
not I_22154 (I378513,I378496);
nor I_22155 (I378530,I378380,I378513);
nand I_22156 (I378298,I378530,I378445);
nor I_22157 (I378286,I378513,I378462);
nand I_22158 (I378292,I378445,I378513);
nor I_22159 (I378589,I378380,I378479);
nand I_22160 (I378606,I378589,I378445);
nand I_22161 (I378623,I378513,I378606);
DFFARX1 I_22162 (I378623,I1862,I378312,I378295,);
not I_22163 (I378654,I378479);
or I_22164 (I378671,I378445,I378654);
nor I_22165 (I378289,I378411,I378671);
nor I_22166 (I378702,I378380,I378654);
nand I_22167 (I378304,I378702,I378411);
not I_22168 (I378754,I1869);
and I_22169 (I378771,I109567,I109573);
nor I_22170 (I378788,I378771,I109573);
nand I_22171 (I378805,I109576,I109582);
nor I_22172 (I378822,I378805,I378788);
not I_22173 (I378743,I378822);
not I_22174 (I378853,I378805);
or I_22175 (I378870,I109570,I109570);
nor I_22176 (I378887,I378870,I109585);
nor I_22177 (I378904,I378887,I378853);
nand I_22178 (I378921,I109579,I109567);
nor I_22179 (I378938,I378921,I109576);
not I_22180 (I378955,I378938);
nor I_22181 (I378972,I378822,I378955);
nand I_22182 (I378740,I378972,I378887);
nor I_22183 (I378728,I378955,I378904);
nand I_22184 (I378734,I378887,I378955);
nor I_22185 (I379031,I378822,I378921);
nand I_22186 (I379048,I379031,I378887);
nand I_22187 (I379065,I378955,I379048);
DFFARX1 I_22188 (I379065,I1862,I378754,I378737,);
not I_22189 (I379096,I378921);
or I_22190 (I379113,I378887,I379096);
nor I_22191 (I378731,I378853,I379113);
nor I_22192 (I379144,I378822,I379096);
nand I_22193 (I378746,I379144,I378853);
not I_22194 (I379196,I1869);
and I_22195 (I379213,I269141,I269147);
nor I_22196 (I379230,I379213,I269135);
nand I_22197 (I379247,I269132,I269129);
nor I_22198 (I379264,I379247,I379230);
not I_22199 (I379185,I379264);
not I_22200 (I379295,I379247);
or I_22201 (I379312,I269138,I269150);
nor I_22202 (I379329,I379312,I269132);
nor I_22203 (I379346,I379329,I379295);
nand I_22204 (I379363,I269129,I269144);
nor I_22205 (I379380,I379363,I269135);
not I_22206 (I379397,I379380);
nor I_22207 (I379414,I379264,I379397);
nand I_22208 (I379182,I379414,I379329);
nor I_22209 (I379170,I379397,I379346);
nand I_22210 (I379176,I379329,I379397);
nor I_22211 (I379473,I379264,I379363);
nand I_22212 (I379490,I379473,I379329);
nand I_22213 (I379507,I379397,I379490);
DFFARX1 I_22214 (I379507,I1862,I379196,I379179,);
not I_22215 (I379538,I379363);
or I_22216 (I379555,I379329,I379538);
nor I_22217 (I379173,I379295,I379555);
nor I_22218 (I379586,I379264,I379538);
nand I_22219 (I379188,I379586,I379295);
not I_22220 (I379638,I1869);
and I_22221 (I379655,I157898,I157898);
nor I_22222 (I379672,I379655,I157922);
nand I_22223 (I379689,I157919,I157907);
nor I_22224 (I379706,I379689,I379672);
not I_22225 (I379627,I379706);
not I_22226 (I379737,I379689);
or I_22227 (I379754,I157901,I157901);
nor I_22228 (I379771,I379754,I157904);
nor I_22229 (I379788,I379771,I379737);
nand I_22230 (I379805,I157913,I157916);
nor I_22231 (I379822,I379805,I157910);
not I_22232 (I379839,I379822);
nor I_22233 (I379856,I379706,I379839);
nand I_22234 (I379624,I379856,I379771);
nor I_22235 (I379612,I379839,I379788);
nand I_22236 (I379618,I379771,I379839);
nor I_22237 (I379915,I379706,I379805);
nand I_22238 (I379932,I379915,I379771);
nand I_22239 (I379949,I379839,I379932);
DFFARX1 I_22240 (I379949,I1862,I379638,I379621,);
not I_22241 (I379980,I379805);
or I_22242 (I379997,I379771,I379980);
nor I_22243 (I379615,I379737,I379997);
nor I_22244 (I380028,I379706,I379980);
nand I_22245 (I379630,I380028,I379737);
not I_22246 (I380080,I1869);
and I_22247 (I380097,I67057,I67033);
nor I_22248 (I380114,I380097,I67039);
nand I_22249 (I380131,I67054,I67036);
nor I_22250 (I380148,I380131,I380114);
not I_22251 (I380069,I380148);
not I_22252 (I380179,I380131);
or I_22253 (I380196,I67033,I67036);
nor I_22254 (I380213,I380196,I67048);
nor I_22255 (I380230,I380213,I380179);
nand I_22256 (I380247,I67042,I67045);
nor I_22257 (I380264,I380247,I67051);
not I_22258 (I380281,I380264);
nor I_22259 (I380298,I380148,I380281);
nand I_22260 (I380066,I380298,I380213);
nor I_22261 (I380054,I380281,I380230);
nand I_22262 (I380060,I380213,I380281);
nor I_22263 (I380357,I380148,I380247);
nand I_22264 (I380374,I380357,I380213);
nand I_22265 (I380391,I380281,I380374);
DFFARX1 I_22266 (I380391,I1862,I380080,I380063,);
not I_22267 (I380422,I380247);
or I_22268 (I380439,I380213,I380422);
nor I_22269 (I380057,I380179,I380439);
nor I_22270 (I380470,I380148,I380422);
nand I_22271 (I380072,I380470,I380179);
not I_22272 (I380522,I1869);
and I_22273 (I380539,I30337,I30313);
nor I_22274 (I380556,I380539,I30319);
nand I_22275 (I380573,I30334,I30316);
nor I_22276 (I380590,I380573,I380556);
not I_22277 (I380511,I380590);
not I_22278 (I380621,I380573);
or I_22279 (I380638,I30313,I30316);
nor I_22280 (I380655,I380638,I30328);
nor I_22281 (I380672,I380655,I380621);
nand I_22282 (I380689,I30322,I30325);
nor I_22283 (I380706,I380689,I30331);
not I_22284 (I380723,I380706);
nor I_22285 (I380740,I380590,I380723);
nand I_22286 (I380508,I380740,I380655);
nor I_22287 (I380496,I380723,I380672);
nand I_22288 (I380502,I380655,I380723);
nor I_22289 (I380799,I380590,I380689);
nand I_22290 (I380816,I380799,I380655);
nand I_22291 (I380833,I380723,I380816);
DFFARX1 I_22292 (I380833,I1862,I380522,I380505,);
not I_22293 (I380864,I380689);
or I_22294 (I380881,I380655,I380864);
nor I_22295 (I380499,I380621,I380881);
nor I_22296 (I380912,I380590,I380864);
nand I_22297 (I380514,I380912,I380621);
not I_22298 (I380964,I1869);
and I_22299 (I380981,I125224,I125224);
nor I_22300 (I380998,I380981,I125248);
nand I_22301 (I381015,I125245,I125233);
nor I_22302 (I381032,I381015,I380998);
not I_22303 (I380953,I381032);
not I_22304 (I381063,I381015);
or I_22305 (I381080,I125227,I125227);
nor I_22306 (I381097,I381080,I125230);
nor I_22307 (I381114,I381097,I381063);
nand I_22308 (I381131,I125239,I125242);
nor I_22309 (I381148,I381131,I125236);
not I_22310 (I381165,I381148);
nor I_22311 (I381182,I381032,I381165);
nand I_22312 (I380950,I381182,I381097);
nor I_22313 (I380938,I381165,I381114);
nand I_22314 (I380944,I381097,I381165);
nor I_22315 (I381241,I381032,I381131);
nand I_22316 (I381258,I381241,I381097);
nand I_22317 (I381275,I381165,I381258);
DFFARX1 I_22318 (I381275,I1862,I380964,I380947,);
not I_22319 (I381306,I381131);
or I_22320 (I381323,I381097,I381306);
nor I_22321 (I380941,I381063,I381323);
nor I_22322 (I381354,I381032,I381306);
nand I_22323 (I380956,I381354,I381063);
not I_22324 (I381406,I1869);
and I_22325 (I381423,I22687,I22663);
nor I_22326 (I381440,I381423,I22669);
nand I_22327 (I381457,I22684,I22666);
nor I_22328 (I381474,I381457,I381440);
not I_22329 (I381395,I381474);
not I_22330 (I381505,I381457);
or I_22331 (I381522,I22663,I22666);
nor I_22332 (I381539,I381522,I22678);
nor I_22333 (I381556,I381539,I381505);
nand I_22334 (I381573,I22672,I22675);
nor I_22335 (I381590,I381573,I22681);
not I_22336 (I381607,I381590);
nor I_22337 (I381624,I381474,I381607);
nand I_22338 (I381392,I381624,I381539);
nor I_22339 (I381380,I381607,I381556);
nand I_22340 (I381386,I381539,I381607);
nor I_22341 (I381683,I381474,I381573);
nand I_22342 (I381700,I381683,I381539);
nand I_22343 (I381717,I381607,I381700);
DFFARX1 I_22344 (I381717,I1862,I381406,I381389,);
not I_22345 (I381748,I381573);
or I_22346 (I381765,I381539,I381748);
nor I_22347 (I381383,I381505,I381765);
nor I_22348 (I381796,I381474,I381748);
nand I_22349 (I381398,I381796,I381505);
not I_22350 (I381848,I1869);
and I_22351 (I381865,I220113,I220119);
nor I_22352 (I381882,I381865,I220107);
nand I_22353 (I381899,I220104,I220101);
nor I_22354 (I381916,I381899,I381882);
not I_22355 (I381837,I381916);
not I_22356 (I381947,I381899);
or I_22357 (I381964,I220110,I220122);
nor I_22358 (I381981,I381964,I220104);
nor I_22359 (I381998,I381981,I381947);
nand I_22360 (I382015,I220101,I220116);
nor I_22361 (I382032,I382015,I220107);
not I_22362 (I382049,I382032);
nor I_22363 (I382066,I381916,I382049);
nand I_22364 (I381834,I382066,I381981);
nor I_22365 (I381822,I382049,I381998);
nand I_22366 (I381828,I381981,I382049);
nor I_22367 (I382125,I381916,I382015);
nand I_22368 (I382142,I382125,I381981);
nand I_22369 (I382159,I382049,I382142);
DFFARX1 I_22370 (I382159,I1862,I381848,I381831,);
not I_22371 (I382190,I382015);
or I_22372 (I382207,I381981,I382190);
nor I_22373 (I381825,I381947,I382207);
nor I_22374 (I382238,I381916,I382190);
nand I_22375 (I381840,I382238,I381947);
not I_22376 (I382290,I1869);
and I_22377 (I382307,I349472,I349457);
nor I_22378 (I382324,I382307,I349460);
nand I_22379 (I382341,I349454,I349454);
nor I_22380 (I382358,I382341,I382324);
not I_22381 (I382279,I382358);
not I_22382 (I382389,I382341);
or I_22383 (I382406,I349457,I349475);
nor I_22384 (I382423,I382406,I349466);
nor I_22385 (I382440,I382423,I382389);
nand I_22386 (I382457,I349469,I349463);
nor I_22387 (I382474,I382457,I349460);
not I_22388 (I382491,I382474);
nor I_22389 (I382508,I382358,I382491);
nand I_22390 (I382276,I382508,I382423);
nor I_22391 (I382264,I382491,I382440);
nand I_22392 (I382270,I382423,I382491);
nor I_22393 (I382567,I382358,I382457);
nand I_22394 (I382584,I382567,I382423);
nand I_22395 (I382601,I382491,I382584);
DFFARX1 I_22396 (I382601,I1862,I382290,I382273,);
not I_22397 (I382632,I382457);
or I_22398 (I382649,I382423,I382632);
nor I_22399 (I382267,I382389,I382649);
nor I_22400 (I382680,I382358,I382632);
nand I_22401 (I382282,I382680,I382389);
not I_22402 (I382732,I1869);
and I_22403 (I382749,I288870,I288852);
nor I_22404 (I382766,I382749,I288867);
nand I_22405 (I382783,I288864,I288855);
nor I_22406 (I382800,I382783,I382766);
not I_22407 (I382721,I382800);
not I_22408 (I382831,I382783);
or I_22409 (I382848,I288849,I288855);
nor I_22410 (I382865,I382848,I288849);
nor I_22411 (I382882,I382865,I382831);
nand I_22412 (I382899,I288858,I288861);
nor I_22413 (I382916,I382899,I288852);
not I_22414 (I382933,I382916);
nor I_22415 (I382950,I382800,I382933);
nand I_22416 (I382718,I382950,I382865);
nor I_22417 (I382706,I382933,I382882);
nand I_22418 (I382712,I382865,I382933);
nor I_22419 (I383009,I382800,I382899);
nand I_22420 (I383026,I383009,I382865);
nand I_22421 (I383043,I382933,I383026);
DFFARX1 I_22422 (I383043,I1862,I382732,I382715,);
not I_22423 (I383074,I382899);
or I_22424 (I383091,I382865,I383074);
nor I_22425 (I382709,I382831,I383091);
nor I_22426 (I383122,I382800,I383074);
nand I_22427 (I382724,I383122,I382831);
not I_22428 (I383174,I1869);
and I_22429 (I383191,I272949,I272955);
nor I_22430 (I383208,I383191,I272943);
nand I_22431 (I383225,I272940,I272937);
nor I_22432 (I383242,I383225,I383208);
not I_22433 (I383163,I383242);
not I_22434 (I383273,I383225);
or I_22435 (I383290,I272946,I272958);
nor I_22436 (I383307,I383290,I272940);
nor I_22437 (I383324,I383307,I383273);
nand I_22438 (I383341,I272937,I272952);
nor I_22439 (I383358,I383341,I272943);
not I_22440 (I383375,I383358);
nor I_22441 (I383392,I383242,I383375);
nand I_22442 (I383160,I383392,I383307);
nor I_22443 (I383148,I383375,I383324);
nand I_22444 (I383154,I383307,I383375);
nor I_22445 (I383451,I383242,I383341);
nand I_22446 (I383468,I383451,I383307);
nand I_22447 (I383485,I383375,I383468);
DFFARX1 I_22448 (I383485,I1862,I383174,I383157,);
not I_22449 (I383516,I383341);
or I_22450 (I383533,I383307,I383516);
nor I_22451 (I383151,I383273,I383533);
nor I_22452 (I383564,I383242,I383516);
nand I_22453 (I383166,I383564,I383273);
not I_22454 (I383616,I1869);
and I_22455 (I383633,I183721,I183721);
nor I_22456 (I383650,I383633,I183745);
nand I_22457 (I383667,I183742,I183730);
nor I_22458 (I383684,I383667,I383650);
not I_22459 (I383605,I383684);
not I_22460 (I383715,I383667);
or I_22461 (I383732,I183724,I183724);
nor I_22462 (I383749,I383732,I183727);
nor I_22463 (I383766,I383749,I383715);
nand I_22464 (I383783,I183736,I183739);
nor I_22465 (I383800,I383783,I183733);
not I_22466 (I383817,I383800);
nor I_22467 (I383834,I383684,I383817);
nand I_22468 (I383602,I383834,I383749);
nor I_22469 (I383590,I383817,I383766);
nand I_22470 (I383596,I383749,I383817);
nor I_22471 (I383893,I383684,I383783);
nand I_22472 (I383910,I383893,I383749);
nand I_22473 (I383927,I383817,I383910);
DFFARX1 I_22474 (I383927,I1862,I383616,I383599,);
not I_22475 (I383958,I383783);
or I_22476 (I383975,I383749,I383958);
nor I_22477 (I383593,I383715,I383975);
nor I_22478 (I384006,I383684,I383958);
nand I_22479 (I383608,I384006,I383715);
not I_22480 (I384058,I1869);
and I_22481 (I384075,I102631,I102637);
nor I_22482 (I384092,I384075,I102637);
nand I_22483 (I384109,I102640,I102646);
nor I_22484 (I384126,I384109,I384092);
not I_22485 (I384047,I384126);
not I_22486 (I384157,I384109);
or I_22487 (I384174,I102634,I102634);
nor I_22488 (I384191,I384174,I102649);
nor I_22489 (I384208,I384191,I384157);
nand I_22490 (I384225,I102643,I102631);
nor I_22491 (I384242,I384225,I102640);
not I_22492 (I384259,I384242);
nor I_22493 (I384276,I384126,I384259);
nand I_22494 (I384044,I384276,I384191);
nor I_22495 (I384032,I384259,I384208);
nand I_22496 (I384038,I384191,I384259);
nor I_22497 (I384335,I384126,I384225);
nand I_22498 (I384352,I384335,I384191);
nand I_22499 (I384369,I384259,I384352);
DFFARX1 I_22500 (I384369,I1862,I384058,I384041,);
not I_22501 (I384400,I384225);
or I_22502 (I384417,I384191,I384400);
nor I_22503 (I384035,I384157,I384417);
nor I_22504 (I384448,I384126,I384400);
nand I_22505 (I384050,I384448,I384157);
not I_22506 (I384500,I1869);
and I_22507 (I384517,I326284,I326269);
nor I_22508 (I384534,I384517,I326272);
nand I_22509 (I384551,I326266,I326266);
nor I_22510 (I384568,I384551,I384534);
not I_22511 (I384489,I384568);
not I_22512 (I384599,I384551);
or I_22513 (I384616,I326269,I326287);
nor I_22514 (I384633,I384616,I326278);
nor I_22515 (I384650,I384633,I384599);
nand I_22516 (I384667,I326281,I326275);
nor I_22517 (I384684,I384667,I326272);
not I_22518 (I384701,I384684);
nor I_22519 (I384718,I384568,I384701);
nand I_22520 (I384486,I384718,I384633);
nor I_22521 (I384474,I384701,I384650);
nand I_22522 (I384480,I384633,I384701);
nor I_22523 (I384777,I384568,I384667);
nand I_22524 (I384794,I384777,I384633);
nand I_22525 (I384811,I384701,I384794);
DFFARX1 I_22526 (I384811,I1862,I384500,I384483,);
not I_22527 (I384842,I384667);
or I_22528 (I384859,I384633,I384842);
nor I_22529 (I384477,I384599,I384859);
nor I_22530 (I384890,I384568,I384842);
nand I_22531 (I384492,I384890,I384599);
not I_22532 (I384942,I1869);
and I_22533 (I384959,I119954,I119954);
nor I_22534 (I384976,I384959,I119978);
nand I_22535 (I384993,I119975,I119963);
nor I_22536 (I385010,I384993,I384976);
not I_22537 (I384931,I385010);
not I_22538 (I385041,I384993);
or I_22539 (I385058,I119957,I119957);
nor I_22540 (I385075,I385058,I119960);
nor I_22541 (I385092,I385075,I385041);
nand I_22542 (I385109,I119969,I119972);
nor I_22543 (I385126,I385109,I119966);
not I_22544 (I385143,I385126);
nor I_22545 (I385160,I385010,I385143);
nand I_22546 (I384928,I385160,I385075);
nor I_22547 (I384916,I385143,I385092);
nand I_22548 (I384922,I385075,I385143);
nor I_22549 (I385219,I385010,I385109);
nand I_22550 (I385236,I385219,I385075);
nand I_22551 (I385253,I385143,I385236);
DFFARX1 I_22552 (I385253,I1862,I384942,I384925,);
not I_22553 (I385284,I385109);
or I_22554 (I385301,I385075,I385284);
nor I_22555 (I384919,I385041,I385301);
nor I_22556 (I385332,I385010,I385284);
nand I_22557 (I384934,I385332,I385041);
not I_22558 (I385384,I1869);
and I_22559 (I385401,I274853,I274859);
nor I_22560 (I385418,I385401,I274847);
nand I_22561 (I385435,I274844,I274841);
nor I_22562 (I385452,I385435,I385418);
not I_22563 (I385373,I385452);
not I_22564 (I385483,I385435);
or I_22565 (I385500,I274850,I274862);
nor I_22566 (I385517,I385500,I274844);
nor I_22567 (I385534,I385517,I385483);
nand I_22568 (I385551,I274841,I274856);
nor I_22569 (I385568,I385551,I274847);
not I_22570 (I385585,I385568);
nor I_22571 (I385602,I385452,I385585);
nand I_22572 (I385370,I385602,I385517);
nor I_22573 (I385358,I385585,I385534);
nand I_22574 (I385364,I385517,I385585);
nor I_22575 (I385661,I385452,I385551);
nand I_22576 (I385678,I385661,I385517);
nand I_22577 (I385695,I385585,I385678);
DFFARX1 I_22578 (I385695,I1862,I385384,I385367,);
not I_22579 (I385726,I385551);
or I_22580 (I385743,I385517,I385726);
nor I_22581 (I385361,I385483,I385743);
nor I_22582 (I385774,I385452,I385726);
nand I_22583 (I385376,I385774,I385483);
not I_22584 (I385826,I1869);
and I_22585 (I385843,I88477,I88453);
nor I_22586 (I385860,I385843,I88459);
nand I_22587 (I385877,I88474,I88456);
nor I_22588 (I385894,I385877,I385860);
not I_22589 (I385815,I385894);
not I_22590 (I385925,I385877);
or I_22591 (I385942,I88453,I88456);
nor I_22592 (I385959,I385942,I88468);
nor I_22593 (I385976,I385959,I385925);
nand I_22594 (I385993,I88462,I88465);
nor I_22595 (I386010,I385993,I88471);
not I_22596 (I386027,I386010);
nor I_22597 (I386044,I385894,I386027);
nand I_22598 (I385812,I386044,I385959);
nor I_22599 (I385800,I386027,I385976);
nand I_22600 (I385806,I385959,I386027);
nor I_22601 (I386103,I385894,I385993);
nand I_22602 (I386120,I386103,I385959);
nand I_22603 (I386137,I386027,I386120);
DFFARX1 I_22604 (I386137,I1862,I385826,I385809,);
not I_22605 (I386168,I385993);
or I_22606 (I386185,I385959,I386168);
nor I_22607 (I385803,I385925,I386185);
nor I_22608 (I386216,I385894,I386168);
nand I_22609 (I385818,I386216,I385925);
not I_22610 (I386268,I1869);
and I_22611 (I386285,I105895,I105901);
nor I_22612 (I386302,I386285,I105901);
nand I_22613 (I386319,I105904,I105910);
nor I_22614 (I386336,I386319,I386302);
not I_22615 (I386257,I386336);
not I_22616 (I386367,I386319);
or I_22617 (I386384,I105898,I105898);
nor I_22618 (I386401,I386384,I105913);
nor I_22619 (I386418,I386401,I386367);
nand I_22620 (I386435,I105907,I105895);
nor I_22621 (I386452,I386435,I105904);
not I_22622 (I386469,I386452);
nor I_22623 (I386486,I386336,I386469);
nand I_22624 (I386254,I386486,I386401);
nor I_22625 (I386242,I386469,I386418);
nand I_22626 (I386248,I386401,I386469);
nor I_22627 (I386545,I386336,I386435);
nand I_22628 (I386562,I386545,I386401);
nand I_22629 (I386579,I386469,I386562);
DFFARX1 I_22630 (I386579,I1862,I386268,I386251,);
not I_22631 (I386610,I386435);
or I_22632 (I386627,I386401,I386610);
nor I_22633 (I386245,I386367,I386627);
nor I_22634 (I386658,I386336,I386610);
nand I_22635 (I386260,I386658,I386367);
not I_22636 (I386710,I1869);
and I_22637 (I386727,I190572,I190572);
nor I_22638 (I386744,I386727,I190596);
nand I_22639 (I386761,I190593,I190581);
nor I_22640 (I386778,I386761,I386744);
not I_22641 (I386699,I386778);
not I_22642 (I386809,I386761);
or I_22643 (I386826,I190575,I190575);
nor I_22644 (I386843,I386826,I190578);
nor I_22645 (I386860,I386843,I386809);
nand I_22646 (I386877,I190587,I190590);
nor I_22647 (I386894,I386877,I190584);
not I_22648 (I386911,I386894);
nor I_22649 (I386928,I386778,I386911);
nand I_22650 (I386696,I386928,I386843);
nor I_22651 (I386684,I386911,I386860);
nand I_22652 (I386690,I386843,I386911);
nor I_22653 (I386987,I386778,I386877);
nand I_22654 (I387004,I386987,I386843);
nand I_22655 (I387021,I386911,I387004);
DFFARX1 I_22656 (I387021,I1862,I386710,I386693,);
not I_22657 (I387052,I386877);
or I_22658 (I387069,I386843,I387052);
nor I_22659 (I386687,I386809,I387069);
nor I_22660 (I387100,I386778,I387052);
nand I_22661 (I386702,I387100,I386809);
not I_22662 (I387152,I1869);
and I_22663 (I387169,I52267,I52243);
nor I_22664 (I387186,I387169,I52249);
nand I_22665 (I387203,I52264,I52246);
nor I_22666 (I387220,I387203,I387186);
not I_22667 (I387141,I387220);
not I_22668 (I387251,I387203);
or I_22669 (I387268,I52243,I52246);
nor I_22670 (I387285,I387268,I52258);
nor I_22671 (I387302,I387285,I387251);
nand I_22672 (I387319,I52252,I52255);
nor I_22673 (I387336,I387319,I52261);
not I_22674 (I387353,I387336);
nor I_22675 (I387370,I387220,I387353);
nand I_22676 (I387138,I387370,I387285);
nor I_22677 (I387126,I387353,I387302);
nand I_22678 (I387132,I387285,I387353);
nor I_22679 (I387429,I387220,I387319);
nand I_22680 (I387446,I387429,I387285);
nand I_22681 (I387463,I387353,I387446);
DFFARX1 I_22682 (I387463,I1862,I387152,I387135,);
not I_22683 (I387494,I387319);
or I_22684 (I387511,I387285,I387494);
nor I_22685 (I387129,I387251,I387511);
nor I_22686 (I387542,I387220,I387494);
nand I_22687 (I387144,I387542,I387251);
not I_22688 (I387594,I1869);
and I_22689 (I387611,I127859,I127859);
nor I_22690 (I387628,I387611,I127883);
nand I_22691 (I387645,I127880,I127868);
nor I_22692 (I387662,I387645,I387628);
not I_22693 (I387583,I387662);
not I_22694 (I387693,I387645);
or I_22695 (I387710,I127862,I127862);
nor I_22696 (I387727,I387710,I127865);
nor I_22697 (I387744,I387727,I387693);
nand I_22698 (I387761,I127874,I127877);
nor I_22699 (I387778,I387761,I127871);
not I_22700 (I387795,I387778);
nor I_22701 (I387812,I387662,I387795);
nand I_22702 (I387580,I387812,I387727);
nor I_22703 (I387568,I387795,I387744);
nand I_22704 (I387574,I387727,I387795);
nor I_22705 (I387871,I387662,I387761);
nand I_22706 (I387888,I387871,I387727);
nand I_22707 (I387905,I387795,I387888);
DFFARX1 I_22708 (I387905,I1862,I387594,I387577,);
not I_22709 (I387936,I387761);
or I_22710 (I387953,I387727,I387936);
nor I_22711 (I387571,I387693,I387953);
nor I_22712 (I387984,I387662,I387936);
nand I_22713 (I387586,I387984,I387693);
not I_22714 (I388036,I1869);
and I_22715 (I388053,I284373,I284379);
nor I_22716 (I388070,I388053,I284367);
nand I_22717 (I388087,I284364,I284361);
nor I_22718 (I388104,I388087,I388070);
not I_22719 (I388025,I388104);
not I_22720 (I388135,I388087);
or I_22721 (I388152,I284370,I284382);
nor I_22722 (I388169,I388152,I284364);
nor I_22723 (I388186,I388169,I388135);
nand I_22724 (I388203,I284361,I284376);
nor I_22725 (I388220,I388203,I284367);
not I_22726 (I388237,I388220);
nor I_22727 (I388254,I388104,I388237);
nand I_22728 (I388022,I388254,I388169);
nor I_22729 (I388010,I388237,I388186);
nand I_22730 (I388016,I388169,I388237);
nor I_22731 (I388313,I388104,I388203);
nand I_22732 (I388330,I388313,I388169);
nand I_22733 (I388347,I388237,I388330);
DFFARX1 I_22734 (I388347,I1862,I388036,I388019,);
not I_22735 (I388378,I388203);
or I_22736 (I388395,I388169,I388378);
nor I_22737 (I388013,I388135,I388395);
nor I_22738 (I388426,I388104,I388378);
nand I_22739 (I388028,I388426,I388135);
not I_22740 (I388478,I1869);
and I_22741 (I388495,I76237,I76213);
nor I_22742 (I388512,I388495,I76219);
nand I_22743 (I388529,I76234,I76216);
nor I_22744 (I388546,I388529,I388512);
not I_22745 (I388467,I388546);
not I_22746 (I388577,I388529);
or I_22747 (I388594,I76213,I76216);
nor I_22748 (I388611,I388594,I76228);
nor I_22749 (I388628,I388611,I388577);
nand I_22750 (I388645,I76222,I76225);
nor I_22751 (I388662,I388645,I76231);
not I_22752 (I388679,I388662);
nor I_22753 (I388696,I388546,I388679);
nand I_22754 (I388464,I388696,I388611);
nor I_22755 (I388452,I388679,I388628);
nand I_22756 (I388458,I388611,I388679);
nor I_22757 (I388755,I388546,I388645);
nand I_22758 (I388772,I388755,I388611);
nand I_22759 (I388789,I388679,I388772);
DFFARX1 I_22760 (I388789,I1862,I388478,I388461,);
not I_22761 (I388820,I388645);
or I_22762 (I388837,I388611,I388820);
nor I_22763 (I388455,I388577,I388837);
nor I_22764 (I388868,I388546,I388820);
nand I_22765 (I388470,I388868,I388577);
not I_22766 (I388920,I1869);
and I_22767 (I388937,I111607,I111613);
nor I_22768 (I388954,I388937,I111613);
nand I_22769 (I388971,I111616,I111622);
nor I_22770 (I388988,I388971,I388954);
not I_22771 (I388909,I388988);
not I_22772 (I389019,I388971);
or I_22773 (I389036,I111610,I111610);
nor I_22774 (I389053,I389036,I111625);
nor I_22775 (I389070,I389053,I389019);
nand I_22776 (I389087,I111619,I111607);
nor I_22777 (I389104,I389087,I111616);
not I_22778 (I389121,I389104);
nor I_22779 (I389138,I388988,I389121);
nand I_22780 (I388906,I389138,I389053);
nor I_22781 (I388894,I389121,I389070);
nand I_22782 (I388900,I389053,I389121);
nor I_22783 (I389197,I388988,I389087);
nand I_22784 (I389214,I389197,I389053);
nand I_22785 (I389231,I389121,I389214);
DFFARX1 I_22786 (I389231,I1862,I388920,I388903,);
not I_22787 (I389262,I389087);
or I_22788 (I389279,I389053,I389262);
nor I_22789 (I388897,I389019,I389279);
nor I_22790 (I389310,I388988,I389262);
nand I_22791 (I388912,I389310,I389019);
not I_22792 (I389362,I1869);
and I_22793 (I389379,I24727,I24703);
nor I_22794 (I389396,I389379,I24709);
nand I_22795 (I389413,I24724,I24706);
nor I_22796 (I389430,I389413,I389396);
not I_22797 (I389351,I389430);
not I_22798 (I389461,I389413);
or I_22799 (I389478,I24703,I24706);
nor I_22800 (I389495,I389478,I24718);
nor I_22801 (I389512,I389495,I389461);
nand I_22802 (I389529,I24712,I24715);
nor I_22803 (I389546,I389529,I24721);
not I_22804 (I389563,I389546);
nor I_22805 (I389580,I389430,I389563);
nand I_22806 (I389348,I389580,I389495);
nor I_22807 (I389336,I389563,I389512);
nand I_22808 (I389342,I389495,I389563);
nor I_22809 (I389639,I389430,I389529);
nand I_22810 (I389656,I389639,I389495);
nand I_22811 (I389673,I389563,I389656);
DFFARX1 I_22812 (I389673,I1862,I389362,I389345,);
not I_22813 (I389704,I389529);
or I_22814 (I389721,I389495,I389704);
nor I_22815 (I389339,I389461,I389721);
nor I_22816 (I389752,I389430,I389704);
nand I_22817 (I389354,I389752,I389461);
not I_22818 (I389804,I1869);
and I_22819 (I389821,I228205,I228211);
nor I_22820 (I389838,I389821,I228199);
nand I_22821 (I389855,I228196,I228193);
nor I_22822 (I389872,I389855,I389838);
not I_22823 (I389793,I389872);
not I_22824 (I389903,I389855);
or I_22825 (I389920,I228202,I228214);
nor I_22826 (I389937,I389920,I228196);
nor I_22827 (I389954,I389937,I389903);
nand I_22828 (I389971,I228193,I228208);
nor I_22829 (I389988,I389971,I228199);
not I_22830 (I390005,I389988);
nor I_22831 (I390022,I389872,I390005);
nand I_22832 (I389790,I390022,I389937);
nor I_22833 (I389778,I390005,I389954);
nand I_22834 (I389784,I389937,I390005);
nor I_22835 (I390081,I389872,I389971);
nand I_22836 (I390098,I390081,I389937);
nand I_22837 (I390115,I390005,I390098);
DFFARX1 I_22838 (I390115,I1862,I389804,I389787,);
not I_22839 (I390146,I389971);
or I_22840 (I390163,I389937,I390146);
nor I_22841 (I389781,I389903,I390163);
nor I_22842 (I390194,I389872,I390146);
nand I_22843 (I389796,I390194,I389903);
not I_22844 (I390246,I1869);
and I_22845 (I390263,I81847,I81823);
nor I_22846 (I390280,I390263,I81829);
nand I_22847 (I390297,I81844,I81826);
nor I_22848 (I390314,I390297,I390280);
not I_22849 (I390235,I390314);
not I_22850 (I390345,I390297);
or I_22851 (I390362,I81823,I81826);
nor I_22852 (I390379,I390362,I81838);
nor I_22853 (I390396,I390379,I390345);
nand I_22854 (I390413,I81832,I81835);
nor I_22855 (I390430,I390413,I81841);
not I_22856 (I390447,I390430);
nor I_22857 (I390464,I390314,I390447);
nand I_22858 (I390232,I390464,I390379);
nor I_22859 (I390220,I390447,I390396);
nand I_22860 (I390226,I390379,I390447);
nor I_22861 (I390523,I390314,I390413);
nand I_22862 (I390540,I390523,I390379);
nand I_22863 (I390557,I390447,I390540);
DFFARX1 I_22864 (I390557,I1862,I390246,I390229,);
not I_22865 (I390588,I390413);
or I_22866 (I390605,I390379,I390588);
nor I_22867 (I390223,I390345,I390605);
nor I_22868 (I390636,I390314,I390588);
nand I_22869 (I390238,I390636,I390345);
not I_22870 (I390688,I1869);
and I_22871 (I390705,I85417,I85393);
nor I_22872 (I390722,I390705,I85399);
nand I_22873 (I390739,I85414,I85396);
nor I_22874 (I390756,I390739,I390722);
not I_22875 (I390677,I390756);
not I_22876 (I390787,I390739);
or I_22877 (I390804,I85393,I85396);
nor I_22878 (I390821,I390804,I85408);
nor I_22879 (I390838,I390821,I390787);
nand I_22880 (I390855,I85402,I85405);
nor I_22881 (I390872,I390855,I85411);
not I_22882 (I390889,I390872);
nor I_22883 (I390906,I390756,I390889);
nand I_22884 (I390674,I390906,I390821);
nor I_22885 (I390662,I390889,I390838);
nand I_22886 (I390668,I390821,I390889);
nor I_22887 (I390965,I390756,I390855);
nand I_22888 (I390982,I390965,I390821);
nand I_22889 (I390999,I390889,I390982);
DFFARX1 I_22890 (I390999,I1862,I390688,I390671,);
not I_22891 (I391030,I390855);
or I_22892 (I391047,I390821,I391030);
nor I_22893 (I390665,I390787,I391047);
nor I_22894 (I391078,I390756,I391030);
nand I_22895 (I390680,I391078,I390787);
not I_22896 (I391130,I1869);
and I_22897 (I391147,I271045,I271051);
nor I_22898 (I391164,I391147,I271039);
nand I_22899 (I391181,I271036,I271033);
nor I_22900 (I391198,I391181,I391164);
not I_22901 (I391119,I391198);
not I_22902 (I391229,I391181);
or I_22903 (I391246,I271042,I271054);
nor I_22904 (I391263,I391246,I271036);
nor I_22905 (I391280,I391263,I391229);
nand I_22906 (I391297,I271033,I271048);
nor I_22907 (I391314,I391297,I271039);
not I_22908 (I391331,I391314);
nor I_22909 (I391348,I391198,I391331);
nand I_22910 (I391116,I391348,I391263);
nor I_22911 (I391104,I391331,I391280);
nand I_22912 (I391110,I391263,I391331);
nor I_22913 (I391407,I391198,I391297);
nand I_22914 (I391424,I391407,I391263);
nand I_22915 (I391441,I391331,I391424);
DFFARX1 I_22916 (I391441,I1862,I391130,I391113,);
not I_22917 (I391472,I391297);
or I_22918 (I391489,I391263,I391472);
nor I_22919 (I391107,I391229,I391489);
nor I_22920 (I391520,I391198,I391472);
nand I_22921 (I391122,I391520,I391229);
not I_22922 (I391572,I1869);
and I_22923 (I391589,I222017,I222023);
nor I_22924 (I391606,I391589,I222011);
nand I_22925 (I391623,I222008,I222005);
nor I_22926 (I391640,I391623,I391606);
not I_22927 (I391561,I391640);
not I_22928 (I391671,I391623);
or I_22929 (I391688,I222014,I222026);
nor I_22930 (I391705,I391688,I222008);
nor I_22931 (I391722,I391705,I391671);
nand I_22932 (I391739,I222005,I222020);
nor I_22933 (I391756,I391739,I222011);
not I_22934 (I391773,I391756);
nor I_22935 (I391790,I391640,I391773);
nand I_22936 (I391558,I391790,I391705);
nor I_22937 (I391546,I391773,I391722);
nand I_22938 (I391552,I391705,I391773);
nor I_22939 (I391849,I391640,I391739);
nand I_22940 (I391866,I391849,I391705);
nand I_22941 (I391883,I391773,I391866);
DFFARX1 I_22942 (I391883,I1862,I391572,I391555,);
not I_22943 (I391914,I391739);
or I_22944 (I391931,I391705,I391914);
nor I_22945 (I391549,I391671,I391931);
nor I_22946 (I391962,I391640,I391914);
nand I_22947 (I391564,I391962,I391671);
not I_22948 (I392014,I1869);
and I_22949 (I392031,I318906,I318891);
nor I_22950 (I392048,I392031,I318894);
nand I_22951 (I392065,I318888,I318888);
nor I_22952 (I392082,I392065,I392048);
not I_22953 (I392003,I392082);
not I_22954 (I392113,I392065);
or I_22955 (I392130,I318891,I318909);
nor I_22956 (I392147,I392130,I318900);
nor I_22957 (I392164,I392147,I392113);
nand I_22958 (I392181,I318903,I318897);
nor I_22959 (I392198,I392181,I318894);
not I_22960 (I392215,I392198);
nor I_22961 (I392232,I392082,I392215);
nand I_22962 (I392000,I392232,I392147);
nor I_22963 (I391988,I392215,I392164);
nand I_22964 (I391994,I392147,I392215);
nor I_22965 (I392291,I392082,I392181);
nand I_22966 (I392308,I392291,I392147);
nand I_22967 (I392325,I392215,I392308);
DFFARX1 I_22968 (I392325,I1862,I392014,I391997,);
not I_22969 (I392356,I392181);
or I_22970 (I392373,I392147,I392356);
nor I_22971 (I391991,I392113,I392373);
nor I_22972 (I392404,I392082,I392356);
nand I_22973 (I392006,I392404,I392113);
not I_22974 (I392456,I1869);
and I_22975 (I392473,I182667,I182667);
nor I_22976 (I392490,I392473,I182691);
nand I_22977 (I392507,I182688,I182676);
nor I_22978 (I392524,I392507,I392490);
not I_22979 (I392445,I392524);
not I_22980 (I392555,I392507);
or I_22981 (I392572,I182670,I182670);
nor I_22982 (I392589,I392572,I182673);
nor I_22983 (I392606,I392589,I392555);
nand I_22984 (I392623,I182682,I182685);
nor I_22985 (I392640,I392623,I182679);
not I_22986 (I392657,I392640);
nor I_22987 (I392674,I392524,I392657);
nand I_22988 (I392442,I392674,I392589);
nor I_22989 (I392430,I392657,I392606);
nand I_22990 (I392436,I392589,I392657);
nor I_22991 (I392733,I392524,I392623);
nand I_22992 (I392750,I392733,I392589);
nand I_22993 (I392767,I392657,I392750);
DFFARX1 I_22994 (I392767,I1862,I392456,I392439,);
not I_22995 (I392798,I392623);
or I_22996 (I392815,I392589,I392798);
nor I_22997 (I392433,I392555,I392815);
nor I_22998 (I392846,I392524,I392798);
nand I_22999 (I392448,I392846,I392555);
not I_23000 (I392898,I1869);
and I_23001 (I392915,I223445,I223451);
nor I_23002 (I392932,I392915,I223439);
nand I_23003 (I392949,I223436,I223433);
nor I_23004 (I392966,I392949,I392932);
not I_23005 (I392887,I392966);
not I_23006 (I392997,I392949);
or I_23007 (I393014,I223442,I223454);
nor I_23008 (I393031,I393014,I223436);
nor I_23009 (I393048,I393031,I392997);
nand I_23010 (I393065,I223433,I223448);
nor I_23011 (I393082,I393065,I223439);
not I_23012 (I393099,I393082);
nor I_23013 (I393116,I392966,I393099);
nand I_23014 (I392884,I393116,I393031);
nor I_23015 (I392872,I393099,I393048);
nand I_23016 (I392878,I393031,I393099);
nor I_23017 (I393175,I392966,I393065);
nand I_23018 (I393192,I393175,I393031);
nand I_23019 (I393209,I393099,I393192);
DFFARX1 I_23020 (I393209,I1862,I392898,I392881,);
not I_23021 (I393240,I393065);
or I_23022 (I393257,I393031,I393240);
nor I_23023 (I392875,I392997,I393257);
nor I_23024 (I393288,I392966,I393240);
nand I_23025 (I392890,I393288,I392997);
not I_23026 (I393340,I1869);
and I_23027 (I393357,I103447,I103453);
nor I_23028 (I393374,I393357,I103453);
nand I_23029 (I393391,I103456,I103462);
nor I_23030 (I393408,I393391,I393374);
not I_23031 (I393329,I393408);
not I_23032 (I393439,I393391);
or I_23033 (I393456,I103450,I103450);
nor I_23034 (I393473,I393456,I103465);
nor I_23035 (I393490,I393473,I393439);
nand I_23036 (I393507,I103459,I103447);
nor I_23037 (I393524,I393507,I103456);
not I_23038 (I393541,I393524);
nor I_23039 (I393558,I393408,I393541);
nand I_23040 (I393326,I393558,I393473);
nor I_23041 (I393314,I393541,I393490);
nand I_23042 (I393320,I393473,I393541);
nor I_23043 (I393617,I393408,I393507);
nand I_23044 (I393634,I393617,I393473);
nand I_23045 (I393651,I393541,I393634);
DFFARX1 I_23046 (I393651,I1862,I393340,I393323,);
not I_23047 (I393682,I393507);
or I_23048 (I393699,I393473,I393682);
nor I_23049 (I393317,I393439,I393699);
nor I_23050 (I393730,I393408,I393682);
nand I_23051 (I393332,I393730,I393439);
not I_23052 (I393782,I1869);
and I_23053 (I393799,I12954,I12942);
nor I_23054 (I393816,I393799,I12960);
nand I_23055 (I393833,I12948,I12945);
nor I_23056 (I393850,I393833,I393816);
not I_23057 (I393771,I393850);
not I_23058 (I393881,I393833);
or I_23059 (I393898,I12942,I12939);
nor I_23060 (I393915,I393898,I12939);
nor I_23061 (I393932,I393915,I393881);
nand I_23062 (I393949,I12951,I12945);
nor I_23063 (I393966,I393949,I12957);
not I_23064 (I393983,I393966);
nor I_23065 (I394000,I393850,I393983);
nand I_23066 (I393768,I394000,I393915);
nor I_23067 (I393756,I393983,I393932);
nand I_23068 (I393762,I393915,I393983);
nor I_23069 (I394059,I393850,I393949);
nand I_23070 (I394076,I394059,I393915);
nand I_23071 (I394093,I393983,I394076);
DFFARX1 I_23072 (I394093,I1862,I393782,I393765,);
not I_23073 (I394124,I393949);
or I_23074 (I394141,I393915,I394124);
nor I_23075 (I393759,I393881,I394141);
nor I_23076 (I394172,I393850,I394124);
nand I_23077 (I393774,I394172,I393881);
not I_23078 (I394224,I1869);
and I_23079 (I394241,I173708,I173708);
nor I_23080 (I394258,I394241,I173732);
nand I_23081 (I394275,I173729,I173717);
nor I_23082 (I394292,I394275,I394258);
not I_23083 (I394213,I394292);
not I_23084 (I394323,I394275);
or I_23085 (I394340,I173711,I173711);
nor I_23086 (I394357,I394340,I173714);
nor I_23087 (I394374,I394357,I394323);
nand I_23088 (I394391,I173723,I173726);
nor I_23089 (I394408,I394391,I173720);
not I_23090 (I394425,I394408);
nor I_23091 (I394442,I394292,I394425);
nand I_23092 (I394210,I394442,I394357);
nor I_23093 (I394198,I394425,I394374);
nand I_23094 (I394204,I394357,I394425);
nor I_23095 (I394501,I394292,I394391);
nand I_23096 (I394518,I394501,I394357);
nand I_23097 (I394535,I394425,I394518);
DFFARX1 I_23098 (I394535,I1862,I394224,I394207,);
not I_23099 (I394566,I394391);
or I_23100 (I394583,I394357,I394566);
nor I_23101 (I394201,I394323,I394583);
nor I_23102 (I394614,I394292,I394566);
nand I_23103 (I394216,I394614,I394323);
not I_23104 (I394666,I1869);
and I_23105 (I394683,I232965,I232971);
nor I_23106 (I394700,I394683,I232959);
nand I_23107 (I394717,I232956,I232953);
nor I_23108 (I394734,I394717,I394700);
not I_23109 (I394655,I394734);
not I_23110 (I394765,I394717);
or I_23111 (I394782,I232962,I232974);
nor I_23112 (I394799,I394782,I232956);
nor I_23113 (I394816,I394799,I394765);
nand I_23114 (I394833,I232953,I232968);
nor I_23115 (I394850,I394833,I232959);
not I_23116 (I394867,I394850);
nor I_23117 (I394884,I394734,I394867);
nand I_23118 (I394652,I394884,I394799);
nor I_23119 (I394640,I394867,I394816);
nand I_23120 (I394646,I394799,I394867);
nor I_23121 (I394943,I394734,I394833);
nand I_23122 (I394960,I394943,I394799);
nand I_23123 (I394977,I394867,I394960);
DFFARX1 I_23124 (I394977,I1862,I394666,I394649,);
not I_23125 (I395008,I394833);
or I_23126 (I395025,I394799,I395008);
nor I_23127 (I394643,I394765,I395025);
nor I_23128 (I395056,I394734,I395008);
nand I_23129 (I394658,I395056,I394765);
not I_23130 (I395108,I1869);
and I_23131 (I395125,I3468,I3456);
nor I_23132 (I395142,I395125,I3474);
nand I_23133 (I395159,I3462,I3459);
nor I_23134 (I395176,I395159,I395142);
not I_23135 (I395097,I395176);
not I_23136 (I395207,I395159);
or I_23137 (I395224,I3456,I3453);
nor I_23138 (I395241,I395224,I3453);
nor I_23139 (I395258,I395241,I395207);
nand I_23140 (I395275,I3465,I3459);
nor I_23141 (I395292,I395275,I3471);
not I_23142 (I395309,I395292);
nor I_23143 (I395326,I395176,I395309);
nand I_23144 (I395094,I395326,I395241);
nor I_23145 (I395082,I395309,I395258);
nand I_23146 (I395088,I395241,I395309);
nor I_23147 (I395385,I395176,I395275);
nand I_23148 (I395402,I395385,I395241);
nand I_23149 (I395419,I395309,I395402);
DFFARX1 I_23150 (I395419,I1862,I395108,I395091,);
not I_23151 (I395450,I395275);
or I_23152 (I395467,I395241,I395450);
nor I_23153 (I395085,I395207,I395467);
nor I_23154 (I395498,I395176,I395450);
nand I_23155 (I395100,I395498,I395207);
not I_23156 (I395550,I1869);
and I_23157 (I395567,I258193,I258199);
nor I_23158 (I395584,I395567,I258187);
nand I_23159 (I395601,I258184,I258181);
nor I_23160 (I395618,I395601,I395584);
not I_23161 (I395539,I395618);
not I_23162 (I395649,I395601);
or I_23163 (I395666,I258190,I258202);
nor I_23164 (I395683,I395666,I258184);
nor I_23165 (I395700,I395683,I395649);
nand I_23166 (I395717,I258181,I258196);
nor I_23167 (I395734,I395717,I258187);
not I_23168 (I395751,I395734);
nor I_23169 (I395768,I395618,I395751);
nand I_23170 (I395536,I395768,I395683);
nor I_23171 (I395524,I395751,I395700);
nand I_23172 (I395530,I395683,I395751);
nor I_23173 (I395827,I395618,I395717);
nand I_23174 (I395844,I395827,I395683);
nand I_23175 (I395861,I395751,I395844);
DFFARX1 I_23176 (I395861,I1862,I395550,I395533,);
not I_23177 (I395892,I395717);
or I_23178 (I395909,I395683,I395892);
nor I_23179 (I395527,I395649,I395909);
nor I_23180 (I395940,I395618,I395892);
nand I_23181 (I395542,I395940,I395649);
not I_23182 (I395992,I1869);
and I_23183 (I396009,I339986,I339971);
nor I_23184 (I396026,I396009,I339974);
nand I_23185 (I396043,I339968,I339968);
nor I_23186 (I396060,I396043,I396026);
not I_23187 (I395981,I396060);
not I_23188 (I396091,I396043);
or I_23189 (I396108,I339971,I339989);
nor I_23190 (I396125,I396108,I339980);
nor I_23191 (I396142,I396125,I396091);
nand I_23192 (I396159,I339983,I339977);
nor I_23193 (I396176,I396159,I339974);
not I_23194 (I396193,I396176);
nor I_23195 (I396210,I396060,I396193);
nand I_23196 (I395978,I396210,I396125);
nor I_23197 (I395966,I396193,I396142);
nand I_23198 (I395972,I396125,I396193);
nor I_23199 (I396269,I396060,I396159);
nand I_23200 (I396286,I396269,I396125);
nand I_23201 (I396303,I396193,I396286);
DFFARX1 I_23202 (I396303,I1862,I395992,I395975,);
not I_23203 (I396334,I396159);
or I_23204 (I396351,I396125,I396334);
nor I_23205 (I395969,I396091,I396351);
nor I_23206 (I396382,I396060,I396334);
nand I_23207 (I395984,I396382,I396091);
not I_23208 (I396434,I1869);
and I_23209 (I396451,I220589,I220595);
nor I_23210 (I396468,I396451,I220583);
nand I_23211 (I396485,I220580,I220577);
nor I_23212 (I396502,I396485,I396468);
not I_23213 (I396423,I396502);
not I_23214 (I396533,I396485);
or I_23215 (I396550,I220586,I220598);
nor I_23216 (I396567,I396550,I220580);
nor I_23217 (I396584,I396567,I396533);
nand I_23218 (I396601,I220577,I220592);
nor I_23219 (I396618,I396601,I220583);
not I_23220 (I396635,I396618);
nor I_23221 (I396652,I396502,I396635);
nand I_23222 (I396420,I396652,I396567);
nor I_23223 (I396408,I396635,I396584);
nand I_23224 (I396414,I396567,I396635);
nor I_23225 (I396711,I396502,I396601);
nand I_23226 (I396728,I396711,I396567);
nand I_23227 (I396745,I396635,I396728);
DFFARX1 I_23228 (I396745,I1862,I396434,I396417,);
not I_23229 (I396776,I396601);
or I_23230 (I396793,I396567,I396776);
nor I_23231 (I396411,I396533,I396793);
nor I_23232 (I396824,I396502,I396776);
nand I_23233 (I396426,I396824,I396533);
not I_23234 (I396876,I1869);
and I_23235 (I396893,I256765,I256771);
nor I_23236 (I396910,I396893,I256759);
nand I_23237 (I396927,I256756,I256753);
nor I_23238 (I396944,I396927,I396910);
not I_23239 (I396865,I396944);
not I_23240 (I396975,I396927);
or I_23241 (I396992,I256762,I256774);
nor I_23242 (I397009,I396992,I256756);
nor I_23243 (I397026,I397009,I396975);
nand I_23244 (I397043,I256753,I256768);
nor I_23245 (I397060,I397043,I256759);
not I_23246 (I397077,I397060);
nor I_23247 (I397094,I396944,I397077);
nand I_23248 (I396862,I397094,I397009);
nor I_23249 (I396850,I397077,I397026);
nand I_23250 (I396856,I397009,I397077);
nor I_23251 (I397153,I396944,I397043);
nand I_23252 (I397170,I397153,I397009);
nand I_23253 (I397187,I397077,I397170);
DFFARX1 I_23254 (I397187,I1862,I396876,I396859,);
not I_23255 (I397218,I397043);
or I_23256 (I397235,I397009,I397218);
nor I_23257 (I396853,I396975,I397235);
nor I_23258 (I397266,I396944,I397218);
nand I_23259 (I396868,I397266,I396975);
not I_23260 (I397318,I1869);
and I_23261 (I397335,I263429,I263435);
nor I_23262 (I397352,I397335,I263423);
nand I_23263 (I397369,I263420,I263417);
nor I_23264 (I397386,I397369,I397352);
not I_23265 (I397307,I397386);
not I_23266 (I397417,I397369);
or I_23267 (I397434,I263426,I263438);
nor I_23268 (I397451,I397434,I263420);
nor I_23269 (I397468,I397451,I397417);
nand I_23270 (I397485,I263417,I263432);
nor I_23271 (I397502,I397485,I263423);
not I_23272 (I397519,I397502);
nor I_23273 (I397536,I397386,I397519);
nand I_23274 (I397304,I397536,I397451);
nor I_23275 (I397292,I397519,I397468);
nand I_23276 (I397298,I397451,I397519);
nor I_23277 (I397595,I397386,I397485);
nand I_23278 (I397612,I397595,I397451);
nand I_23279 (I397629,I397519,I397612);
DFFARX1 I_23280 (I397629,I1862,I397318,I397301,);
not I_23281 (I397660,I397485);
or I_23282 (I397677,I397451,I397660);
nor I_23283 (I397295,I397417,I397677);
nor I_23284 (I397708,I397386,I397660);
nand I_23285 (I397310,I397708,I397417);
not I_23286 (I397760,I1869);
and I_23287 (I397777,I39007,I38983);
nor I_23288 (I397794,I397777,I38989);
nand I_23289 (I397811,I39004,I38986);
nor I_23290 (I397828,I397811,I397794);
not I_23291 (I397749,I397828);
not I_23292 (I397859,I397811);
or I_23293 (I397876,I38983,I38986);
nor I_23294 (I397893,I397876,I38998);
nor I_23295 (I397910,I397893,I397859);
nand I_23296 (I397927,I38992,I38995);
nor I_23297 (I397944,I397927,I39001);
not I_23298 (I397961,I397944);
nor I_23299 (I397978,I397828,I397961);
nand I_23300 (I397746,I397978,I397893);
nor I_23301 (I397734,I397961,I397910);
nand I_23302 (I397740,I397893,I397961);
nor I_23303 (I398037,I397828,I397927);
nand I_23304 (I398054,I398037,I397893);
nand I_23305 (I398071,I397961,I398054);
DFFARX1 I_23306 (I398071,I1862,I397760,I397743,);
not I_23307 (I398102,I397927);
or I_23308 (I398119,I397893,I398102);
nor I_23309 (I397737,I397859,I398119);
nor I_23310 (I398150,I397828,I398102);
nand I_23311 (I397752,I398150,I397859);
not I_23312 (I398202,I1869);
and I_23313 (I398219,I46657,I46633);
nor I_23314 (I398236,I398219,I46639);
nand I_23315 (I398253,I46654,I46636);
nor I_23316 (I398270,I398253,I398236);
not I_23317 (I398191,I398270);
not I_23318 (I398301,I398253);
or I_23319 (I398318,I46633,I46636);
nor I_23320 (I398335,I398318,I46648);
nor I_23321 (I398352,I398335,I398301);
nand I_23322 (I398369,I46642,I46645);
nor I_23323 (I398386,I398369,I46651);
not I_23324 (I398403,I398386);
nor I_23325 (I398420,I398270,I398403);
nand I_23326 (I398188,I398420,I398335);
nor I_23327 (I398176,I398403,I398352);
nand I_23328 (I398182,I398335,I398403);
nor I_23329 (I398479,I398270,I398369);
nand I_23330 (I398496,I398479,I398335);
nand I_23331 (I398513,I398403,I398496);
DFFARX1 I_23332 (I398513,I1862,I398202,I398185,);
not I_23333 (I398544,I398369);
or I_23334 (I398561,I398335,I398544);
nor I_23335 (I398179,I398301,I398561);
nor I_23336 (I398592,I398270,I398544);
nand I_23337 (I398194,I398592,I398301);
not I_23338 (I398644,I1869);
and I_23339 (I398661,I252481,I252487);
nor I_23340 (I398678,I398661,I252475);
nand I_23341 (I398695,I252472,I252469);
nor I_23342 (I398712,I398695,I398678);
not I_23343 (I398633,I398712);
not I_23344 (I398743,I398695);
or I_23345 (I398760,I252478,I252490);
nor I_23346 (I398777,I398760,I252472);
nor I_23347 (I398794,I398777,I398743);
nand I_23348 (I398811,I252469,I252484);
nor I_23349 (I398828,I398811,I252475);
not I_23350 (I398845,I398828);
nor I_23351 (I398862,I398712,I398845);
nand I_23352 (I398630,I398862,I398777);
nor I_23353 (I398618,I398845,I398794);
nand I_23354 (I398624,I398777,I398845);
nor I_23355 (I398921,I398712,I398811);
nand I_23356 (I398938,I398921,I398777);
nand I_23357 (I398955,I398845,I398938);
DFFARX1 I_23358 (I398955,I1862,I398644,I398627,);
not I_23359 (I398986,I398811);
or I_23360 (I399003,I398777,I398986);
nor I_23361 (I398621,I398743,I399003);
nor I_23362 (I399034,I398712,I398986);
nand I_23363 (I398636,I399034,I398743);
not I_23364 (I399086,I1869);
and I_23365 (I399103,I100207,I100183);
nor I_23366 (I399120,I399103,I100189);
nand I_23367 (I399137,I100204,I100186);
nor I_23368 (I399154,I399137,I399120);
not I_23369 (I399075,I399154);
not I_23370 (I399185,I399137);
or I_23371 (I399202,I100183,I100186);
nor I_23372 (I399219,I399202,I100198);
nor I_23373 (I399236,I399219,I399185);
nand I_23374 (I399253,I100192,I100195);
nor I_23375 (I399270,I399253,I100201);
not I_23376 (I399287,I399270);
nor I_23377 (I399304,I399154,I399287);
nand I_23378 (I399072,I399304,I399219);
nor I_23379 (I399060,I399287,I399236);
nand I_23380 (I399066,I399219,I399287);
nor I_23381 (I399363,I399154,I399253);
nand I_23382 (I399380,I399363,I399219);
nand I_23383 (I399397,I399287,I399380);
DFFARX1 I_23384 (I399397,I1862,I399086,I399069,);
not I_23385 (I399428,I399253);
or I_23386 (I399445,I399219,I399428);
nor I_23387 (I399063,I399185,I399445);
nor I_23388 (I399476,I399154,I399428);
nand I_23389 (I399078,I399476,I399185);
not I_23390 (I399528,I1869);
and I_23391 (I399545,I354742,I354727);
nor I_23392 (I399562,I399545,I354730);
nand I_23393 (I399579,I354724,I354724);
nor I_23394 (I399596,I399579,I399562);
not I_23395 (I399517,I399596);
not I_23396 (I399627,I399579);
or I_23397 (I399644,I354727,I354745);
nor I_23398 (I399661,I399644,I354736);
nor I_23399 (I399678,I399661,I399627);
nand I_23400 (I399695,I354739,I354733);
nor I_23401 (I399712,I399695,I354730);
not I_23402 (I399729,I399712);
nor I_23403 (I399746,I399596,I399729);
nand I_23404 (I399514,I399746,I399661);
nor I_23405 (I399502,I399729,I399678);
nand I_23406 (I399508,I399661,I399729);
nor I_23407 (I399805,I399596,I399695);
nand I_23408 (I399822,I399805,I399661);
nand I_23409 (I399839,I399729,I399822);
DFFARX1 I_23410 (I399839,I1862,I399528,I399511,);
not I_23411 (I399870,I399695);
or I_23412 (I399887,I399661,I399870);
nor I_23413 (I399505,I399627,I399887);
nor I_23414 (I399918,I399596,I399870);
nand I_23415 (I399520,I399918,I399627);
not I_23416 (I399970,I1869);
and I_23417 (I399987,I285325,I285331);
nor I_23418 (I400004,I399987,I285319);
nand I_23419 (I400021,I285316,I285313);
nor I_23420 (I400038,I400021,I400004);
not I_23421 (I399959,I400038);
not I_23422 (I400069,I400021);
or I_23423 (I400086,I285322,I285334);
nor I_23424 (I400103,I400086,I285316);
nor I_23425 (I400120,I400103,I400069);
nand I_23426 (I400137,I285313,I285328);
nor I_23427 (I400154,I400137,I285319);
not I_23428 (I400171,I400154);
nor I_23429 (I400188,I400038,I400171);
nand I_23430 (I399956,I400188,I400103);
nor I_23431 (I399944,I400171,I400120);
nand I_23432 (I399950,I400103,I400171);
nor I_23433 (I400247,I400038,I400137);
nand I_23434 (I400264,I400247,I400103);
nand I_23435 (I400281,I400171,I400264);
DFFARX1 I_23436 (I400281,I1862,I399970,I399953,);
not I_23437 (I400312,I400137);
or I_23438 (I400329,I400103,I400312);
nor I_23439 (I399947,I400069,I400329);
nor I_23440 (I400360,I400038,I400312);
nand I_23441 (I399962,I400360,I400069);
not I_23442 (I400412,I1869);
and I_23443 (I400429,I212497,I212503);
nor I_23444 (I400446,I400429,I212491);
nand I_23445 (I400463,I212488,I212485);
nor I_23446 (I400480,I400463,I400446);
not I_23447 (I400401,I400480);
not I_23448 (I400511,I400463);
or I_23449 (I400528,I212494,I212506);
nor I_23450 (I400545,I400528,I212488);
nor I_23451 (I400562,I400545,I400511);
nand I_23452 (I400579,I212485,I212500);
nor I_23453 (I400596,I400579,I212491);
not I_23454 (I400613,I400596);
nor I_23455 (I400630,I400480,I400613);
nand I_23456 (I400398,I400630,I400545);
nor I_23457 (I400386,I400613,I400562);
nand I_23458 (I400392,I400545,I400613);
nor I_23459 (I400689,I400480,I400579);
nand I_23460 (I400706,I400689,I400545);
nand I_23461 (I400723,I400613,I400706);
DFFARX1 I_23462 (I400723,I1862,I400412,I400395,);
not I_23463 (I400754,I400579);
or I_23464 (I400771,I400545,I400754);
nor I_23465 (I400389,I400511,I400771);
nor I_23466 (I400802,I400480,I400754);
nand I_23467 (I400404,I400802,I400511);
not I_23468 (I400854,I1869);
and I_23469 (I400871,I97657,I97633);
nor I_23470 (I400888,I400871,I97639);
nand I_23471 (I400905,I97654,I97636);
nor I_23472 (I400922,I400905,I400888);
not I_23473 (I400843,I400922);
not I_23474 (I400953,I400905);
or I_23475 (I400970,I97633,I97636);
nor I_23476 (I400987,I400970,I97648);
nor I_23477 (I401004,I400987,I400953);
nand I_23478 (I401021,I97642,I97645);
nor I_23479 (I401038,I401021,I97651);
not I_23480 (I401055,I401038);
nor I_23481 (I401072,I400922,I401055);
nand I_23482 (I400840,I401072,I400987);
nor I_23483 (I400828,I401055,I401004);
nand I_23484 (I400834,I400987,I401055);
nor I_23485 (I401131,I400922,I401021);
nand I_23486 (I401148,I401131,I400987);
nand I_23487 (I401165,I401055,I401148);
DFFARX1 I_23488 (I401165,I1862,I400854,I400837,);
not I_23489 (I401196,I401021);
or I_23490 (I401213,I400987,I401196);
nor I_23491 (I400831,I400953,I401213);
nor I_23492 (I401244,I400922,I401196);
nand I_23493 (I400846,I401244,I400953);
not I_23494 (I401296,I1869);
and I_23495 (I401313,I293613,I293595);
nor I_23496 (I401330,I401313,I293610);
nand I_23497 (I401347,I293607,I293598);
nor I_23498 (I401364,I401347,I401330);
not I_23499 (I401285,I401364);
not I_23500 (I401395,I401347);
or I_23501 (I401412,I293592,I293598);
nor I_23502 (I401429,I401412,I293592);
nor I_23503 (I401446,I401429,I401395);
nand I_23504 (I401463,I293601,I293604);
nor I_23505 (I401480,I401463,I293595);
not I_23506 (I401497,I401480);
nor I_23507 (I401514,I401364,I401497);
nand I_23508 (I401282,I401514,I401429);
nor I_23509 (I401270,I401497,I401446);
nand I_23510 (I401276,I401429,I401497);
nor I_23511 (I401573,I401364,I401463);
nand I_23512 (I401590,I401573,I401429);
nand I_23513 (I401607,I401497,I401590);
DFFARX1 I_23514 (I401607,I1862,I401296,I401279,);
not I_23515 (I401638,I401463);
or I_23516 (I401655,I401429,I401638);
nor I_23517 (I401273,I401395,I401655);
nor I_23518 (I401686,I401364,I401638);
nand I_23519 (I401288,I401686,I401395);
not I_23520 (I401738,I1869);
and I_23521 (I401755,I240581,I240587);
nor I_23522 (I401772,I401755,I240575);
nand I_23523 (I401789,I240572,I240569);
nor I_23524 (I401806,I401789,I401772);
not I_23525 (I401727,I401806);
not I_23526 (I401837,I401789);
or I_23527 (I401854,I240578,I240590);
nor I_23528 (I401871,I401854,I240572);
nor I_23529 (I401888,I401871,I401837);
nand I_23530 (I401905,I240569,I240584);
nor I_23531 (I401922,I401905,I240575);
not I_23532 (I401939,I401922);
nor I_23533 (I401956,I401806,I401939);
nand I_23534 (I401724,I401956,I401871);
nor I_23535 (I401712,I401939,I401888);
nand I_23536 (I401718,I401871,I401939);
nor I_23537 (I402015,I401806,I401905);
nand I_23538 (I402032,I402015,I401871);
nand I_23539 (I402049,I401939,I402032);
DFFARX1 I_23540 (I402049,I1862,I401738,I401721,);
not I_23541 (I402080,I401905);
or I_23542 (I402097,I401871,I402080);
nor I_23543 (I401715,I401837,I402097);
nor I_23544 (I402128,I401806,I402080);
nand I_23545 (I401730,I402128,I401837);
not I_23546 (I402180,I1869);
and I_23547 (I402197,I19117,I19093);
nor I_23548 (I402214,I402197,I19099);
nand I_23549 (I402231,I19114,I19096);
nor I_23550 (I402248,I402231,I402214);
not I_23551 (I402169,I402248);
not I_23552 (I402279,I402231);
or I_23553 (I402296,I19093,I19096);
nor I_23554 (I402313,I402296,I19108);
nor I_23555 (I402330,I402313,I402279);
nand I_23556 (I402347,I19102,I19105);
nor I_23557 (I402364,I402347,I19111);
not I_23558 (I402381,I402364);
nor I_23559 (I402398,I402248,I402381);
nand I_23560 (I402166,I402398,I402313);
nor I_23561 (I402154,I402381,I402330);
nand I_23562 (I402160,I402313,I402381);
nor I_23563 (I402457,I402248,I402347);
nand I_23564 (I402474,I402457,I402313);
nand I_23565 (I402491,I402381,I402474);
DFFARX1 I_23566 (I402491,I1862,I402180,I402163,);
not I_23567 (I402522,I402347);
or I_23568 (I402539,I402313,I402522);
nor I_23569 (I402157,I402279,I402539);
nor I_23570 (I402570,I402248,I402522);
nand I_23571 (I402172,I402570,I402279);
not I_23572 (I402622,I1869);
and I_23573 (I402639,I196896,I196896);
nor I_23574 (I402656,I402639,I196920);
nand I_23575 (I402673,I196917,I196905);
nor I_23576 (I402690,I402673,I402656);
not I_23577 (I402611,I402690);
not I_23578 (I402721,I402673);
or I_23579 (I402738,I196899,I196899);
nor I_23580 (I402755,I402738,I196902);
nor I_23581 (I402772,I402755,I402721);
nand I_23582 (I402789,I196911,I196914);
nor I_23583 (I402806,I402789,I196908);
not I_23584 (I402823,I402806);
nor I_23585 (I402840,I402690,I402823);
nand I_23586 (I402608,I402840,I402755);
nor I_23587 (I402596,I402823,I402772);
nand I_23588 (I402602,I402755,I402823);
nor I_23589 (I402899,I402690,I402789);
nand I_23590 (I402916,I402899,I402755);
nand I_23591 (I402933,I402823,I402916);
DFFARX1 I_23592 (I402933,I1862,I402622,I402605,);
not I_23593 (I402964,I402789);
or I_23594 (I402981,I402755,I402964);
nor I_23595 (I402599,I402721,I402981);
nor I_23596 (I403012,I402690,I402964);
nand I_23597 (I402614,I403012,I402721);
not I_23598 (I403064,I1869);
and I_23599 (I403081,I271521,I271527);
nor I_23600 (I403098,I403081,I271515);
nand I_23601 (I403115,I271512,I271509);
nor I_23602 (I403132,I403115,I403098);
not I_23603 (I403053,I403132);
not I_23604 (I403163,I403115);
or I_23605 (I403180,I271518,I271530);
nor I_23606 (I403197,I403180,I271512);
nor I_23607 (I403214,I403197,I403163);
nand I_23608 (I403231,I271509,I271524);
nor I_23609 (I403248,I403231,I271515);
not I_23610 (I403265,I403248);
nor I_23611 (I403282,I403132,I403265);
nand I_23612 (I403050,I403282,I403197);
nor I_23613 (I403038,I403265,I403214);
nand I_23614 (I403044,I403197,I403265);
nor I_23615 (I403341,I403132,I403231);
nand I_23616 (I403358,I403341,I403197);
nand I_23617 (I403375,I403265,I403358);
DFFARX1 I_23618 (I403375,I1862,I403064,I403047,);
not I_23619 (I403406,I403231);
or I_23620 (I403423,I403197,I403406);
nor I_23621 (I403041,I403163,I403423);
nor I_23622 (I403454,I403132,I403406);
nand I_23623 (I403056,I403454,I403163);
not I_23624 (I403506,I1869);
and I_23625 (I403523,I265333,I265339);
nor I_23626 (I403540,I403523,I265327);
nand I_23627 (I403557,I265324,I265321);
nor I_23628 (I403574,I403557,I403540);
not I_23629 (I403495,I403574);
not I_23630 (I403605,I403557);
or I_23631 (I403622,I265330,I265342);
nor I_23632 (I403639,I403622,I265324);
nor I_23633 (I403656,I403639,I403605);
nand I_23634 (I403673,I265321,I265336);
nor I_23635 (I403690,I403673,I265327);
not I_23636 (I403707,I403690);
nor I_23637 (I403724,I403574,I403707);
nand I_23638 (I403492,I403724,I403639);
nor I_23639 (I403480,I403707,I403656);
nand I_23640 (I403486,I403639,I403707);
nor I_23641 (I403783,I403574,I403673);
nand I_23642 (I403800,I403783,I403639);
nand I_23643 (I403817,I403707,I403800);
DFFARX1 I_23644 (I403817,I1862,I403506,I403489,);
not I_23645 (I403848,I403673);
or I_23646 (I403865,I403639,I403848);
nor I_23647 (I403483,I403605,I403865);
nor I_23648 (I403896,I403574,I403848);
nand I_23649 (I403498,I403896,I403605);
not I_23650 (I403948,I1869);
and I_23651 (I403965,I2414,I2402);
nor I_23652 (I403982,I403965,I2420);
nand I_23653 (I403999,I2408,I2405);
nor I_23654 (I404016,I403999,I403982);
not I_23655 (I403937,I404016);
not I_23656 (I404047,I403999);
or I_23657 (I404064,I2402,I2399);
nor I_23658 (I404081,I404064,I2399);
nor I_23659 (I404098,I404081,I404047);
nand I_23660 (I404115,I2411,I2405);
nor I_23661 (I404132,I404115,I2417);
not I_23662 (I404149,I404132);
nor I_23663 (I404166,I404016,I404149);
nand I_23664 (I403934,I404166,I404081);
nor I_23665 (I403922,I404149,I404098);
nand I_23666 (I403928,I404081,I404149);
nor I_23667 (I404225,I404016,I404115);
nand I_23668 (I404242,I404225,I404081);
nand I_23669 (I404259,I404149,I404242);
DFFARX1 I_23670 (I404259,I1862,I403948,I403931,);
not I_23671 (I404290,I404115);
or I_23672 (I404307,I404081,I404290);
nor I_23673 (I403925,I404047,I404307);
nor I_23674 (I404338,I404016,I404290);
nand I_23675 (I403940,I404338,I404047);
not I_23676 (I404390,I1869);
and I_23677 (I404407,I344729,I344714);
nor I_23678 (I404424,I404407,I344717);
nand I_23679 (I404441,I344711,I344711);
nor I_23680 (I404458,I404441,I404424);
not I_23681 (I404379,I404458);
not I_23682 (I404489,I404441);
or I_23683 (I404506,I344714,I344732);
nor I_23684 (I404523,I404506,I344723);
nor I_23685 (I404540,I404523,I404489);
nand I_23686 (I404557,I344726,I344720);
nor I_23687 (I404574,I404557,I344717);
not I_23688 (I404591,I404574);
nor I_23689 (I404608,I404458,I404591);
nand I_23690 (I404376,I404608,I404523);
nor I_23691 (I404364,I404591,I404540);
nand I_23692 (I404370,I404523,I404591);
nor I_23693 (I404667,I404458,I404557);
nand I_23694 (I404684,I404667,I404523);
nand I_23695 (I404701,I404591,I404684);
DFFARX1 I_23696 (I404701,I1862,I404390,I404373,);
not I_23697 (I404732,I404557);
or I_23698 (I404749,I404523,I404732);
nor I_23699 (I404367,I404489,I404749);
nor I_23700 (I404780,I404458,I404732);
nand I_23701 (I404382,I404780,I404489);
not I_23702 (I404832,I1869);
and I_23703 (I404849,I316798,I316783);
nor I_23704 (I404866,I404849,I316786);
nand I_23705 (I404883,I316780,I316780);
nor I_23706 (I404900,I404883,I404866);
not I_23707 (I404821,I404900);
not I_23708 (I404931,I404883);
or I_23709 (I404948,I316783,I316801);
nor I_23710 (I404965,I404948,I316792);
nor I_23711 (I404982,I404965,I404931);
nand I_23712 (I404999,I316795,I316789);
nor I_23713 (I405016,I404999,I316786);
not I_23714 (I405033,I405016);
nor I_23715 (I405050,I404900,I405033);
nand I_23716 (I404818,I405050,I404965);
nor I_23717 (I404806,I405033,I404982);
nand I_23718 (I404812,I404965,I405033);
nor I_23719 (I405109,I404900,I404999);
nand I_23720 (I405126,I405109,I404965);
nand I_23721 (I405143,I405033,I405126);
DFFARX1 I_23722 (I405143,I1862,I404832,I404815,);
not I_23723 (I405174,I404999);
or I_23724 (I405191,I404965,I405174);
nor I_23725 (I404809,I404931,I405191);
nor I_23726 (I405222,I404900,I405174);
nand I_23727 (I404824,I405222,I404931);
not I_23728 (I405274,I1869);
and I_23729 (I405291,I328392,I328377);
nor I_23730 (I405308,I405291,I328380);
nand I_23731 (I405325,I328374,I328374);
nor I_23732 (I405342,I405325,I405308);
not I_23733 (I405263,I405342);
not I_23734 (I405373,I405325);
or I_23735 (I405390,I328377,I328395);
nor I_23736 (I405407,I405390,I328386);
nor I_23737 (I405424,I405407,I405373);
nand I_23738 (I405441,I328389,I328383);
nor I_23739 (I405458,I405441,I328380);
not I_23740 (I405475,I405458);
nor I_23741 (I405492,I405342,I405475);
nand I_23742 (I405260,I405492,I405407);
nor I_23743 (I405248,I405475,I405424);
nand I_23744 (I405254,I405407,I405475);
nor I_23745 (I405551,I405342,I405441);
nand I_23746 (I405568,I405551,I405407);
nand I_23747 (I405585,I405475,I405568);
DFFARX1 I_23748 (I405585,I1862,I405274,I405257,);
not I_23749 (I405616,I405441);
or I_23750 (I405633,I405407,I405616);
nor I_23751 (I405251,I405373,I405633);
nor I_23752 (I405664,I405342,I405616);
nand I_23753 (I405266,I405664,I405373);
not I_23754 (I405716,I1869);
and I_23755 (I405733,I97147,I97123);
nor I_23756 (I405750,I405733,I97129);
nand I_23757 (I405767,I97144,I97126);
nor I_23758 (I405784,I405767,I405750);
not I_23759 (I405705,I405784);
not I_23760 (I405815,I405767);
or I_23761 (I405832,I97123,I97126);
nor I_23762 (I405849,I405832,I97138);
nor I_23763 (I405866,I405849,I405815);
nand I_23764 (I405883,I97132,I97135);
nor I_23765 (I405900,I405883,I97141);
not I_23766 (I405917,I405900);
nor I_23767 (I405934,I405784,I405917);
nand I_23768 (I405702,I405934,I405849);
nor I_23769 (I405690,I405917,I405866);
nand I_23770 (I405696,I405849,I405917);
nor I_23771 (I405993,I405784,I405883);
nand I_23772 (I406010,I405993,I405849);
nand I_23773 (I406027,I405917,I406010);
DFFARX1 I_23774 (I406027,I1862,I405716,I405699,);
not I_23775 (I406058,I405883);
or I_23776 (I406075,I405849,I406058);
nor I_23777 (I405693,I405815,I406075);
nor I_23778 (I406106,I405784,I406058);
nand I_23779 (I405708,I406106,I405815);
not I_23780 (I406158,I1869);
and I_23781 (I406175,I332081,I332066);
nor I_23782 (I406192,I406175,I332069);
nand I_23783 (I406209,I332063,I332063);
nor I_23784 (I406226,I406209,I406192);
not I_23785 (I406147,I406226);
not I_23786 (I406257,I406209);
or I_23787 (I406274,I332066,I332084);
nor I_23788 (I406291,I406274,I332075);
nor I_23789 (I406308,I406291,I406257);
nand I_23790 (I406325,I332078,I332072);
nor I_23791 (I406342,I406325,I332069);
not I_23792 (I406359,I406342);
nor I_23793 (I406376,I406226,I406359);
nand I_23794 (I406144,I406376,I406291);
nor I_23795 (I406132,I406359,I406308);
nand I_23796 (I406138,I406291,I406359);
nor I_23797 (I406435,I406226,I406325);
nand I_23798 (I406452,I406435,I406291);
nand I_23799 (I406469,I406359,I406452);
DFFARX1 I_23800 (I406469,I1862,I406158,I406141,);
not I_23801 (I406500,I406325);
or I_23802 (I406517,I406291,I406500);
nor I_23803 (I406135,I406257,I406517);
nor I_23804 (I406548,I406226,I406500);
nand I_23805 (I406150,I406548,I406257);
not I_23806 (I406600,I1869);
and I_23807 (I406617,I343148,I343133);
nor I_23808 (I406634,I406617,I343136);
nand I_23809 (I406651,I343130,I343130);
nor I_23810 (I406668,I406651,I406634);
not I_23811 (I406589,I406668);
not I_23812 (I406699,I406651);
or I_23813 (I406716,I343133,I343151);
nor I_23814 (I406733,I406716,I343142);
nor I_23815 (I406750,I406733,I406699);
nand I_23816 (I406767,I343145,I343139);
nor I_23817 (I406784,I406767,I343136);
not I_23818 (I406801,I406784);
nor I_23819 (I406818,I406668,I406801);
nand I_23820 (I406586,I406818,I406733);
nor I_23821 (I406574,I406801,I406750);
nand I_23822 (I406580,I406733,I406801);
nor I_23823 (I406877,I406668,I406767);
nand I_23824 (I406894,I406877,I406733);
nand I_23825 (I406911,I406801,I406894);
DFFARX1 I_23826 (I406911,I1862,I406600,I406583,);
not I_23827 (I406942,I406767);
or I_23828 (I406959,I406733,I406942);
nor I_23829 (I406577,I406699,I406959);
nor I_23830 (I406990,I406668,I406942);
nand I_23831 (I406592,I406990,I406699);
not I_23832 (I407042,I1869);
and I_23833 (I407059,I321014,I320999);
nor I_23834 (I407076,I407059,I321002);
nand I_23835 (I407093,I320996,I320996);
nor I_23836 (I407110,I407093,I407076);
not I_23837 (I407031,I407110);
not I_23838 (I407141,I407093);
or I_23839 (I407158,I320999,I321017);
nor I_23840 (I407175,I407158,I321008);
nor I_23841 (I407192,I407175,I407141);
nand I_23842 (I407209,I321011,I321005);
nor I_23843 (I407226,I407209,I321002);
not I_23844 (I407243,I407226);
nor I_23845 (I407260,I407110,I407243);
nand I_23846 (I407028,I407260,I407175);
nor I_23847 (I407016,I407243,I407192);
nand I_23848 (I407022,I407175,I407243);
nor I_23849 (I407319,I407110,I407209);
nand I_23850 (I407336,I407319,I407175);
nand I_23851 (I407353,I407243,I407336);
DFFARX1 I_23852 (I407353,I1862,I407042,I407025,);
not I_23853 (I407384,I407209);
or I_23854 (I407401,I407175,I407384);
nor I_23855 (I407019,I407141,I407401);
nor I_23856 (I407432,I407110,I407384);
nand I_23857 (I407034,I407432,I407141);
not I_23858 (I407484,I1869);
and I_23859 (I407501,I165276,I165276);
nor I_23860 (I407518,I407501,I165300);
nand I_23861 (I407535,I165297,I165285);
nor I_23862 (I407552,I407535,I407518);
not I_23863 (I407473,I407552);
not I_23864 (I407583,I407535);
or I_23865 (I407600,I165279,I165279);
nor I_23866 (I407617,I407600,I165282);
nor I_23867 (I407634,I407617,I407583);
nand I_23868 (I407651,I165291,I165294);
nor I_23869 (I407668,I407651,I165288);
not I_23870 (I407685,I407668);
nor I_23871 (I407702,I407552,I407685);
nand I_23872 (I407470,I407702,I407617);
nor I_23873 (I407458,I407685,I407634);
nand I_23874 (I407464,I407617,I407685);
nor I_23875 (I407761,I407552,I407651);
nand I_23876 (I407778,I407761,I407617);
nand I_23877 (I407795,I407685,I407778);
DFFARX1 I_23878 (I407795,I1862,I407484,I407467,);
not I_23879 (I407826,I407651);
or I_23880 (I407843,I407617,I407826);
nor I_23881 (I407461,I407583,I407843);
nor I_23882 (I407874,I407552,I407826);
nand I_23883 (I407476,I407874,I407583);
not I_23884 (I407926,I1869);
and I_23885 (I407943,I344202,I344187);
nor I_23886 (I407960,I407943,I344190);
nand I_23887 (I407977,I344184,I344184);
nor I_23888 (I407994,I407977,I407960);
not I_23889 (I407915,I407994);
not I_23890 (I408025,I407977);
or I_23891 (I408042,I344187,I344205);
nor I_23892 (I408059,I408042,I344196);
nor I_23893 (I408076,I408059,I408025);
nand I_23894 (I408093,I344199,I344193);
nor I_23895 (I408110,I408093,I344190);
not I_23896 (I408127,I408110);
nor I_23897 (I408144,I407994,I408127);
nand I_23898 (I407912,I408144,I408059);
nor I_23899 (I407900,I408127,I408076);
nand I_23900 (I407906,I408059,I408127);
nor I_23901 (I408203,I407994,I408093);
nand I_23902 (I408220,I408203,I408059);
nand I_23903 (I408237,I408127,I408220);
DFFARX1 I_23904 (I408237,I1862,I407926,I407909,);
not I_23905 (I408268,I408093);
or I_23906 (I408285,I408059,I408268);
nor I_23907 (I407903,I408025,I408285);
nor I_23908 (I408316,I407994,I408268);
nand I_23909 (I407918,I408316,I408025);
not I_23910 (I408368,I1869);
and I_23911 (I408385,I143669,I143669);
nor I_23912 (I408402,I408385,I143693);
nand I_23913 (I408419,I143690,I143678);
nor I_23914 (I408436,I408419,I408402);
not I_23915 (I408357,I408436);
not I_23916 (I408467,I408419);
or I_23917 (I408484,I143672,I143672);
nor I_23918 (I408501,I408484,I143675);
nor I_23919 (I408518,I408501,I408467);
nand I_23920 (I408535,I143684,I143687);
nor I_23921 (I408552,I408535,I143681);
not I_23922 (I408569,I408552);
nor I_23923 (I408586,I408436,I408569);
nand I_23924 (I408354,I408586,I408501);
nor I_23925 (I408342,I408569,I408518);
nand I_23926 (I408348,I408501,I408569);
nor I_23927 (I408645,I408436,I408535);
nand I_23928 (I408662,I408645,I408501);
nand I_23929 (I408679,I408569,I408662);
DFFARX1 I_23930 (I408679,I1862,I408368,I408351,);
not I_23931 (I408710,I408535);
or I_23932 (I408727,I408501,I408710);
nor I_23933 (I408345,I408467,I408727);
nor I_23934 (I408758,I408436,I408710);
nand I_23935 (I408360,I408758,I408467);
not I_23936 (I408810,I1869);
and I_23937 (I408827,I351580,I351565);
nor I_23938 (I408844,I408827,I351568);
nand I_23939 (I408861,I351562,I351562);
nor I_23940 (I408878,I408861,I408844);
not I_23941 (I408799,I408878);
not I_23942 (I408909,I408861);
or I_23943 (I408926,I351565,I351583);
nor I_23944 (I408943,I408926,I351574);
nor I_23945 (I408960,I408943,I408909);
nand I_23946 (I408977,I351577,I351571);
nor I_23947 (I408994,I408977,I351568);
not I_23948 (I409011,I408994);
nor I_23949 (I409028,I408878,I409011);
nand I_23950 (I408796,I409028,I408943);
nor I_23951 (I408784,I409011,I408960);
nand I_23952 (I408790,I408943,I409011);
nor I_23953 (I409087,I408878,I408977);
nand I_23954 (I409104,I409087,I408943);
nand I_23955 (I409121,I409011,I409104);
DFFARX1 I_23956 (I409121,I1862,I408810,I408793,);
not I_23957 (I409152,I408977);
or I_23958 (I409169,I408943,I409152);
nor I_23959 (I408787,I408909,I409169);
nor I_23960 (I409200,I408878,I409152);
nand I_23961 (I408802,I409200,I408909);
not I_23962 (I409252,I1869);
and I_23963 (I409269,I356850,I356835);
nor I_23964 (I409286,I409269,I356838);
nand I_23965 (I409303,I356832,I356832);
nor I_23966 (I409320,I409303,I409286);
not I_23967 (I409241,I409320);
not I_23968 (I409351,I409303);
or I_23969 (I409368,I356835,I356853);
nor I_23970 (I409385,I409368,I356844);
nor I_23971 (I409402,I409385,I409351);
nand I_23972 (I409419,I356847,I356841);
nor I_23973 (I409436,I409419,I356838);
not I_23974 (I409453,I409436);
nor I_23975 (I409470,I409320,I409453);
nand I_23976 (I409238,I409470,I409385);
nor I_23977 (I409226,I409453,I409402);
nand I_23978 (I409232,I409385,I409453);
nor I_23979 (I409529,I409320,I409419);
nand I_23980 (I409546,I409529,I409385);
nand I_23981 (I409563,I409453,I409546);
DFFARX1 I_23982 (I409563,I1862,I409252,I409235,);
not I_23983 (I409594,I409419);
or I_23984 (I409611,I409385,I409594);
nor I_23985 (I409229,I409351,I409611);
nor I_23986 (I409642,I409320,I409594);
nand I_23987 (I409244,I409642,I409351);
not I_23988 (I409694,I1869);
and I_23989 (I409711,I113239,I113245);
nor I_23990 (I409728,I409711,I113245);
nand I_23991 (I409745,I113248,I113254);
nor I_23992 (I409762,I409745,I409728);
not I_23993 (I409683,I409762);
not I_23994 (I409793,I409745);
or I_23995 (I409810,I113242,I113242);
nor I_23996 (I409827,I409810,I113257);
nor I_23997 (I409844,I409827,I409793);
nand I_23998 (I409861,I113251,I113239);
nor I_23999 (I409878,I409861,I113248);
not I_24000 (I409895,I409878);
nor I_24001 (I409912,I409762,I409895);
nand I_24002 (I409680,I409912,I409827);
nor I_24003 (I409668,I409895,I409844);
nand I_24004 (I409674,I409827,I409895);
nor I_24005 (I409971,I409762,I409861);
nand I_24006 (I409988,I409971,I409827);
nand I_24007 (I410005,I409895,I409988);
DFFARX1 I_24008 (I410005,I1862,I409694,I409677,);
not I_24009 (I410036,I409861);
or I_24010 (I410053,I409827,I410036);
nor I_24011 (I409671,I409793,I410053);
nor I_24012 (I410084,I409762,I410036);
nand I_24013 (I409686,I410084,I409793);
not I_24014 (I410136,I1869);
and I_24015 (I410153,I80317,I80293);
nor I_24016 (I410170,I410153,I80299);
nand I_24017 (I410187,I80314,I80296);
nor I_24018 (I410204,I410187,I410170);
not I_24019 (I410125,I410204);
not I_24020 (I410235,I410187);
or I_24021 (I410252,I80293,I80296);
nor I_24022 (I410269,I410252,I80308);
nor I_24023 (I410286,I410269,I410235);
nand I_24024 (I410303,I80302,I80305);
nor I_24025 (I410320,I410303,I80311);
not I_24026 (I410337,I410320);
nor I_24027 (I410354,I410204,I410337);
nand I_24028 (I410122,I410354,I410269);
nor I_24029 (I410110,I410337,I410286);
nand I_24030 (I410116,I410269,I410337);
nor I_24031 (I410413,I410204,I410303);
nand I_24032 (I410430,I410413,I410269);
nand I_24033 (I410447,I410337,I410430);
DFFARX1 I_24034 (I410447,I1862,I410136,I410119,);
not I_24035 (I410478,I410303);
or I_24036 (I410495,I410269,I410478);
nor I_24037 (I410113,I410235,I410495);
nor I_24038 (I410526,I410204,I410478);
nand I_24039 (I410128,I410526,I410235);
not I_24040 (I410578,I1869);
and I_24041 (I410595,I34927,I34903);
nor I_24042 (I410612,I410595,I34909);
nand I_24043 (I410629,I34924,I34906);
nor I_24044 (I410646,I410629,I410612);
not I_24045 (I410567,I410646);
not I_24046 (I410677,I410629);
or I_24047 (I410694,I34903,I34906);
nor I_24048 (I410711,I410694,I34918);
nor I_24049 (I410728,I410711,I410677);
nand I_24050 (I410745,I34912,I34915);
nor I_24051 (I410762,I410745,I34921);
not I_24052 (I410779,I410762);
nor I_24053 (I410796,I410646,I410779);
nand I_24054 (I410564,I410796,I410711);
nor I_24055 (I410552,I410779,I410728);
nand I_24056 (I410558,I410711,I410779);
nor I_24057 (I410855,I410646,I410745);
nand I_24058 (I410872,I410855,I410711);
nand I_24059 (I410889,I410779,I410872);
DFFARX1 I_24060 (I410889,I1862,I410578,I410561,);
not I_24061 (I410920,I410745);
or I_24062 (I410937,I410711,I410920);
nor I_24063 (I410555,I410677,I410937);
nor I_24064 (I410968,I410646,I410920);
nand I_24065 (I410570,I410968,I410677);
endmodule


