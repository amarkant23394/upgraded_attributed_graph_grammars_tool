module test_I16818_rst(I1477_rst,I16818_rst);
,I16818_rst);
input I1477_rst;
output I16818_rst;
wire ;
not I_0(I16818_rst,I1477_rst);
endmodule


