module test_I6294(I1477,I1470,I4068,I3969,I6294);
input I1477,I1470,I4068,I3969;
output I6294;
wire I3963,I3966,I3954,I6346,I6363,I6380,I6329,I6493,I4181,I4034,I6541;
nor I_0(I3963,I4181,I4034);
or I_1(I3966,I4068,I4034);
not I_2(I3954,I4068);
nand I_3(I6346,I3969,I3954);
and I_4(I6363,I6346,I3963);
DFFARX1 I_5(I6363,I1470,I6329,,,I6380,);
not I_6(I6329,I1477);
DFFARX1 I_7(I3966,I1470,I6329,,,I6493,);
DFFARX1 I_8(I1470,,,I4181,);
DFFARX1 I_9(I1470,,,I4034,);
and I_10(I6294,I6380,I6541);
DFFARX1 I_11(I6493,I1470,I6329,,,I6541,);
endmodule


