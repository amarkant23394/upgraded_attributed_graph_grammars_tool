module test_I4629(I2441,I1303,I1477,I2294,I1247,I1470,I1239,I2215,I4629);
input I2441,I1303,I1477,I2294,I1247,I1470,I1239,I2215;
output I4629;
wire I2167,I2540,I2173,I2181,I2328,I2509,I2557,I2232,I2458,I2311,I2633;
nand I_0(I2167,I2633,I2328);
nor I_1(I4629,I2167,I2173);
DFFARX1 I_2(I1247,I1470,I2181,,,I2540,);
nand I_3(I2173,I2557,I2509);
not I_4(I2181,I1477);
nor I_5(I2328,I2232,I2311);
nor I_6(I2509,I2458,I2232);
and I_7(I2557,I2540,I1303);
DFFARX1 I_8(I2215,I1470,I2181,,,I2232,);
DFFARX1 I_9(I2441,I1470,I2181,,,I2458,);
not I_10(I2311,I2294);
DFFARX1 I_11(I1239,I1470,I2181,,,I2633,);
endmodule


