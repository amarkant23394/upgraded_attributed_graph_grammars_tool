module test_I16257(I14438,I1477,I13542,I14520,I1470,I13296,I16257);
input I14438,I1477,I13542,I14520,I1470,I13296;
output I16257;
wire I14338,I13177,I14341,I14472,I14455,I14537,I14605,I14370;
DFFARX1 I_0(I14605,I1470,I14370,,,I14338,);
nand I_1(I13177,I13296,I13542);
nand I_2(I16257,I14341,I14338);
DFFARX1 I_3(I14455,I1470,I14370,,,I14341,);
nand I_4(I14472,I14455,I14438);
DFFARX1 I_5(I13177,I1470,I14370,,,I14455,);
DFFARX1 I_6(I14520,I1470,I14370,,,I14537,);
and I_7(I14605,I14537,I14472);
not I_8(I14370,I1477);
endmodule


