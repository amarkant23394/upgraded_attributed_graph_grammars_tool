module test_final(IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_7_r_2,blif_reset_net_7_r_2,N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2);
input IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_7_r_2,blif_reset_net_7_r_2;
output N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2;
wire N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_573_7_r_12,n_549_7_r_12,n_569_7_r_12,n_452_7_r_12,N6147_9_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12,n4_7_l_2,n10_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2;
nor I_0(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_1(N1508_0_r_12,n30_12,n37_12);
nor I_2(N1507_6_r_12,n25_12,n39_12);
nor I_3(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_4(n1_12,blif_clk_net_7_r_2,n10_2,G42_7_r_12,);
nor I_5(n_572_7_r_12,n23_12,n24_12);
nand I_6(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_7(n_549_7_r_12,n27_12,n28_12);
nand I_8(n_569_7_r_12,n25_12,n26_12);
nand I_9(n_452_7_r_12,IN_1_1_l_12,IN_2_1_l_12);
nand I_10(N6147_9_r_12,n30_12,n31_12);
nor I_11(N6134_9_r_12,n35_12,n36_12);
not I_12(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_13(n1_12,n_573_7_r_12);
not I_14(n23_12,n36_12);
nor I_15(n24_12,IN_3_1_l_12,n_452_7_r_12);
nand I_16(n25_12,n23_12,n40_12);
not I_17(n26_12,n35_12);
not I_18(n27_12,N6134_9_r_12);
nand I_19(n28_12,n26_12,n29_12);
not I_20(n29_12,n24_12);
nand I_21(n30_12,n33_12,n41_12);
nand I_22(n31_12,n32_12,n33_12);
nor I_23(n32_12,n26_12,n34_12);
nor I_24(n33_12,IN_1_2_l_12,IN_2_2_l_12);
nor I_25(n34_12,IN_5_2_l_12,n42_12);
nor I_26(n35_12,IN_1_3_l_12,n38_12);
nand I_27(n36_12,IN_1_10_l_12,IN_2_10_l_12);
nand I_28(n37_12,n23_12,n35_12);
or I_29(n38_12,IN_2_3_l_12,IN_3_3_l_12);
not I_30(n39_12,n30_12);
or I_31(n40_12,IN_3_10_l_12,IN_4_10_l_12);
nor I_32(n41_12,n34_12,n36_12);
nor I_33(n42_12,IN_3_2_l_12,IN_4_2_l_12);
nor I_34(N1371_0_r_2,n32_2,n35_2);
nor I_35(N1508_0_r_2,n32_2,n55_2);
not I_36(N1372_1_r_2,n54_2);
nor I_37(N1508_1_r_2,n59_2,n54_2);
nor I_38(N6147_2_r_2,n42_2,n43_2);
nor I_39(N1507_6_r_2,n40_2,n53_2);
nor I_40(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_41(n4_7_r_2,blif_clk_net_7_r_2,n10_2,G42_7_r_2,);
nor I_42(n_572_7_r_2,n36_2,n37_2);
or I_43(n_573_7_r_2,n34_2,n35_2);
nor I_44(n_549_7_r_2,n40_2,n41_2);
nand I_45(n_569_7_r_2,n38_2,n39_2);
nor I_46(n_452_7_r_2,n59_2,n35_2);
nor I_47(n4_7_l_2,n_549_7_r_12,G42_7_r_12);
not I_48(n10_2,blif_reset_net_7_r_2);
DFFARX1 I_49(n4_7_l_2,blif_clk_net_7_r_2,n10_2,n59_2,);
not I_50(n33_2,n59_2);
and I_51(N3_8_l_2,n49_2,n_572_7_r_12);
DFFARX1 I_52(N3_8_l_2,blif_clk_net_7_r_2,n10_2,n32_internal_2,);
not I_53(n32_2,n32_internal_2);
nor I_54(n4_7_r_2,n59_2,n36_2);
not I_55(n34_2,n39_2);
nor I_56(n35_2,N1507_6_r_12,N1508_6_r_12);
nor I_57(n36_2,n_572_7_r_12,n_549_7_r_12);
or I_58(n37_2,N1507_6_r_12,N1371_0_r_12);
not I_59(n38_2,n40_2);
nand I_60(n39_2,n45_2,n57_2);
nor I_61(n40_2,n47_2,N1371_0_r_12);
nor I_62(n41_2,n32_2,n36_2);
not I_63(n42_2,n53_2);
nand I_64(n43_2,n44_2,n45_2);
nand I_65(n44_2,n38_2,n46_2);
not I_66(n45_2,N1371_0_r_12);
nand I_67(n46_2,n47_2,n48_2);
nand I_68(n47_2,n_569_7_r_12,N1508_0_r_12);
or I_69(n48_2,N1508_6_r_12,N6147_9_r_12);
nand I_70(n49_2,N1508_0_r_12,N1507_6_r_12);
nand I_71(n50_2,n51_2,n52_2);
not I_72(n51_2,n47_2);
nand I_73(n52_2,n38_2,n53_2);
nor I_74(n53_2,N1507_6_r_12,n_572_7_r_12);
nand I_75(n54_2,n42_2,n56_2);
nor I_76(n55_2,n34_2,n56_2);
nor I_77(n56_2,N1508_6_r_12,N6147_9_r_12);
nand I_78(n57_2,n58_2,G42_7_r_12);
not I_79(n58_2,N1508_6_r_12);
endmodule


