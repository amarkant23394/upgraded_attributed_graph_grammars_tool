module test_I2173(I1303,I1247,I1477,I1327,I1470,I2198,I2424,I1271,I2173);
input I1303,I1247,I1477,I1327,I1470,I2198,I2424,I1271;
output I2173;
wire I2540,I2441,I2181,I2509,I2557,I2232,I2458,I2215;
DFFARX1 I_0(I1247,I1470,I2181,,,I2540,);
and I_1(I2441,I2424,I1327);
nand I_2(I2173,I2557,I2509);
not I_3(I2181,I1477);
nor I_4(I2509,I2458,I2232);
and I_5(I2557,I2540,I1303);
DFFARX1 I_6(I2215,I1470,I2181,,,I2232,);
DFFARX1 I_7(I2441,I1470,I2181,,,I2458,);
and I_8(I2215,I2198,I1271);
endmodule


