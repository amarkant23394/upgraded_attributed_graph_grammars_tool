module test_I17375(I15594,I16162,I1477,I15832,I1470,I15585,I17375);
input I15594,I16162,I1477,I15832,I1470,I15585;
output I17375;
wire I17413,I15597,I17775,I17532,I17854,I17871,I17447,I17464;
not I_0(I17413,I1477);
nor I_1(I15597,I15832,I16162);
DFFARX1 I_2(I15585,I1470,I17413,,,I17775,);
not I_3(I17532,I15597);
nand I_4(I17854,I17775,I17464);
and I_5(I17871,I17532,I17854);
nor I_6(I17447,I15597);
nand I_7(I17464,I17447,I15594);
DFFARX1 I_8(I17871,I1470,I17413,,,I17375,);
endmodule


