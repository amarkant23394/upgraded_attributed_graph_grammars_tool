module test_I5416(I1477,I3504,I1470,I1498,I5416);
input I1477,I3504,I1470,I1498;
output I5416;
wire I3388,I3350,I3668,I3521,I5122,I3555,I3589,I1495,I3405,I3685,I3356,I3572;
nand I_0(I5416,I5122,I3356);
not I_1(I3388,I1477);
DFFARX1 I_2(I3685,I1470,I3388,,,I3350,);
DFFARX1 I_3(I1470,I3388,,,I3668,);
nor I_4(I3521,I3504,I1495);
not I_5(I5122,I3350);
DFFARX1 I_6(I1470,I3388,,,I3555,);
and I_7(I3589,I3521,I3572);
DFFARX1 I_8(I1470,,,I1495,);
or I_9(I3405,I1495);
and I_10(I3685,I3668,I1498);
DFFARX1 I_11(I3589,I1470,I3388,,,I3356,);
nand I_12(I3572,I3555,I3405);
endmodule


