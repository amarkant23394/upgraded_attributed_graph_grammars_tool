module test_I7714(I6442,I3966,I3957,I1470_clk,I1477_rst,I7714);
input I6442,I3966,I3957,I1470_clk,I1477_rst;
output I7714;
wire I6843,I6826,I6493,I6781,I6329_rst,I6297;
and I_0(I6843,I6493,I6826);
nand I_1(I6826,I6781,I6442);
DFFARX1 I_2 (I3966,I1470_clk,I6329_rst,I6493);
DFFARX1 I_3 (I3957,I1470_clk,I6329_rst,I6781);
not I_4(I6329_rst,I1477_rst);
DFFARX1 I_5 (I6843,I1470_clk,I6329_rst,I6297);
not I_6(I7714,I6297);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule