module test_I2575(I1911,I2344,I2022,I1294,I1301,I2575);
input I1911,I2344,I2022,I1294,I1301;
output I2575;
wire I2668,I3120,I2897,I3137,I2600,I3103,I2583,I2651,I1914,I1923,I3086;
nand I_0(I2668,I2651,I1914);
nand I_1(I3120,I3103,I2668);
nand I_2(I2897,I2600,I1923);
and I_3(I3137,I2897,I3120);
not I_4(I2600,I1911);
not I_5(I3103,I3086);
DFFARX1 I_6(I3137,I1294,I2583,,,I2575,);
not I_7(I2583,I1301);
nor I_8(I2651,I2600);
DFFARX1 I_9(I1294,,,I1914,);
nand I_10(I1923,I2022,I2344);
DFFARX1 I_11(I1294,I2583,,,I3086,);
endmodule


