module test_final(G18_1_l_3,G15_1_l_3,IN_1_1_l_3,IN_4_1_l_3,IN_5_1_l_3,IN_7_1_l_3,IN_9_1_l_3,IN_10_1_l_3,IN_1_3_l_3,IN_2_3_l_3,IN_4_3_l_3,blif_clk_net_1_r_17,blif_reset_net_1_r_17,G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17);
input G18_1_l_3,G15_1_l_3,IN_1_1_l_3,IN_4_1_l_3,IN_5_1_l_3,IN_7_1_l_3,IN_9_1_l_3,IN_10_1_l_3,IN_1_3_l_3,IN_2_3_l_3,IN_4_3_l_3,blif_clk_net_1_r_17,blif_reset_net_1_r_17;
output G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17;
wire G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3,n4_1_l_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n_431_0_l_17,n6_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17;
DFFARX1 I_0(n4_1_r_3,blif_clk_net_1_r_17,n6_17,G42_1_r_3,);
nor I_1(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_2(n_573_1_r_3,n26_3,n27_3);
nor I_3(n_549_1_r_3,n40_3,n32_3);
nand I_4(n_569_1_r_3,n27_3,n31_3);
and I_5(n_452_1_r_3,G18_1_l_3,n26_3);
nor I_6(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_7(N3_2_r_3,blif_clk_net_1_r_17,n6_17,G199_2_r_3,);
DFFARX1 I_8(n_572_1_l_3,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_3,);
nor I_9(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_10(n4_1_l_3,G18_1_l_3,IN_1_1_l_3);
DFFARX1 I_11(n4_1_l_3,blif_clk_net_1_r_17,n6_17,G42_1_l_3,);
not I_12(n22_3,G42_1_l_3);
DFFARX1 I_13(IN_1_3_l_3,blif_clk_net_1_r_17,n6_17,n40_3,);
DFFARX1 I_14(IN_2_3_l_3,blif_clk_net_1_r_17,n6_17,n25_internal_3,);
not I_15(n25_3,n25_internal_3);
nor I_16(n4_1_r_3,n40_3,n36_3);
nor I_17(N3_2_r_3,n26_3,n37_3);
nor I_18(n_572_1_l_3,G15_1_l_3,IN_7_1_l_3);
DFFARX1 I_19(G42_1_l_3,blif_clk_net_1_r_17,n6_17,ACVQN1_3_r_3,);
nor I_20(n26_3,IN_5_1_l_3,IN_9_1_l_3);
not I_21(n27_3,IN_10_1_l_3);
nor I_22(n28_3,IN_10_1_l_3,n29_3);
nor I_23(n29_3,G15_1_l_3,n30_3);
not I_24(n30_3,IN_4_1_l_3);
nor I_25(n31_3,IN_9_1_l_3,n40_3);
nor I_26(n32_3,n25_3,n33_3);
nand I_27(n33_3,IN_4_3_l_3,n22_3);
or I_28(n34_3,IN_9_1_l_3,IN_10_1_l_3);
nand I_29(n35_3,IN_4_3_l_3,ACVQN1_3_r_3);
nor I_30(n36_3,G18_1_l_3,IN_5_1_l_3);
nor I_31(n37_3,n38_3,n39_3);
not I_32(n38_3,n_572_1_l_3);
nand I_33(n39_3,n27_3,n30_3);
DFFARX1 I_34(n4_1_r_17,blif_clk_net_1_r_17,n6_17,G42_1_r_17,);
nor I_35(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_36(n_573_1_r_17,n20_17,n21_17);
nand I_37(n_549_1_r_17,n23_17,n24_17);
nand I_38(n_569_1_r_17,n21_17,n22_17);
not I_39(n_452_1_r_17,n23_17);
DFFARX1 I_40(n19_17,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_17,);
nor I_41(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_42(N1_4_r_17,blif_clk_net_1_r_17,n6_17,G199_4_r_17,);
DFFARX1 I_43(n5_17,blif_clk_net_1_r_17,n6_17,G214_4_r_17,);
or I_44(n_431_0_l_17,n26_17,G42_1_r_3);
not I_45(n6_17,blif_reset_net_1_r_17);
DFFARX1 I_46(n_431_0_l_17,blif_clk_net_1_r_17,n6_17,n20_internal_17,);
not I_47(n20_17,n20_internal_17);
DFFARX1 I_48(ACVQN2_3_r_3,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_17,);
DFFARX1 I_49(G42_1_r_3,blif_clk_net_1_r_17,n6_17,n19_internal_17,);
not I_50(n19_17,n19_internal_17);
nor I_51(n4_1_r_17,n5_17,n25_17);
not I_52(n2_17,n29_17);
DFFARX1 I_53(n2_17,blif_clk_net_1_r_17,n6_17,n17_internal_17,);
not I_54(n17_17,n17_internal_17);
nor I_55(N1_4_r_17,n29_17,n31_17);
not I_56(n5_17,n_266_and_0_3_r_3);
and I_57(n21_17,n32_17,G199_2_r_3);
not I_58(n22_17,n25_17);
nand I_59(n23_17,n20_17,n22_17);
nand I_60(n24_17,n19_17,n22_17);
nand I_61(n25_17,n30_17,n_42_2_r_3);
and I_62(n26_17,n27_17,n_573_1_r_3);
nor I_63(n27_17,n28_17,n_452_1_r_3);
not I_64(n28_17,n_569_1_r_3);
nor I_65(n29_17,n28_17,n_572_1_r_3);
and I_66(n30_17,n5_17,n_572_1_r_3);
nor I_67(n31_17,n21_17,n_266_and_0_3_r_3);
nor I_68(n32_17,n_549_1_r_3,n_266_and_0_3_r_3);
endmodule


