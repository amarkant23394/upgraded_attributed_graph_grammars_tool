module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_6,blif_reset_net_1_r_6,G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_6,blif_reset_net_1_r_6;
output G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6;
wire G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_452_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10,N3_2_l_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10,N3_2_l_6,n4_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6;
DFFARX1 I_0(n4_1_r_10,blif_clk_net_1_r_6,n4_6,G42_1_r_10,);
nor I_1(n_572_1_r_10,n26_10,n3_10);
nand I_2(n_573_1_r_10,n16_10,n18_10);
nand I_3(n_549_1_r_10,n19_10,n20_10);
nor I_4(n_452_1_r_10,n25_10,n21_10);
nor I_5(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_6(N3_2_r_10,blif_clk_net_1_r_6,n4_6,G199_2_r_10,);
DFFARX1 I_7(G199_4_l_10,blif_clk_net_1_r_6,n4_6,ACVQN2_3_r_10,);
nor I_8(n_266_and_0_3_r_10,n17_10,n13_10);
and I_9(N3_2_l_10,IN_6_2_l_10,n23_10);
DFFARX1 I_10(N3_2_l_10,blif_clk_net_1_r_6,n4_6,n25_10,);
not I_11(n16_10,n25_10);
DFFARX1 I_12(IN_1_3_l_10,blif_clk_net_1_r_6,n4_6,n26_10,);
DFFARX1 I_13(IN_2_3_l_10,blif_clk_net_1_r_6,n4_6,ACVQN1_3_l_10,);
and I_14(N1_4_l_10,IN_6_4_l_10,n24_10);
DFFARX1 I_15(N1_4_l_10,blif_clk_net_1_r_6,n4_6,G199_4_l_10,);
DFFARX1 I_16(IN_3_4_l_10,blif_clk_net_1_r_6,n4_6,n27_10,);
not I_17(n17_10,n27_10);
nor I_18(n4_1_r_10,n27_10,n21_10);
nor I_19(N3_2_r_10,n16_10,n22_10);
not I_20(n3_10,n18_10);
DFFARX1 I_21(n3_10,blif_clk_net_1_r_6,n4_6,n13_internal_10,);
not I_22(n13_10,n13_internal_10);
nand I_23(n18_10,IN_4_3_l_10,ACVQN1_3_l_10);
not I_24(n19_10,n_452_1_r_10);
nand I_25(n20_10,n16_10,n26_10);
nor I_26(n21_10,IN_1_2_l_10,IN_3_2_l_10);
and I_27(n22_10,n26_10,n21_10);
nand I_28(n23_10,IN_2_2_l_10,IN_3_2_l_10);
nand I_29(n24_10,IN_1_4_l_10,IN_2_4_l_10);
DFFARX1 I_30(n4_1_r_6,blif_clk_net_1_r_6,n4_6,G42_1_r_6,);
nor I_31(n_572_1_r_6,n27_6,n28_6);
nand I_32(n_573_1_r_6,n18_6,n19_6);
nor I_33(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_34(n_569_1_r_6,n19_6,n20_6);
nor I_35(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_36(N1_4_r_6,blif_clk_net_1_r_6,n4_6,G199_4_r_6,);
DFFARX1 I_37(n_42_2_l_6,blif_clk_net_1_r_6,n4_6,G214_4_r_6,);
DFFARX1 I_38(n_42_2_l_6,blif_clk_net_1_r_6,n4_6,ACVQN1_5_r_6,);
not I_39(P6_5_r_6,P6_5_r_internal_6);
and I_40(N3_2_l_6,n23_6,G199_2_r_10);
not I_41(n4_6,blif_reset_net_1_r_6);
DFFARX1 I_42(N3_2_l_6,blif_clk_net_1_r_6,n4_6,n27_6,);
not I_43(n17_6,n27_6);
DFFARX1 I_44(n_266_and_0_3_r_10,blif_clk_net_1_r_6,n4_6,n28_6,);
DFFARX1 I_45(n_549_1_r_10,blif_clk_net_1_r_6,n4_6,n26_6,);
and I_46(N1_4_l_6,n25_6,n_573_1_r_10);
DFFARX1 I_47(N1_4_l_6,blif_clk_net_1_r_6,n4_6,n29_6,);
not I_48(n18_6,n29_6);
DFFARX1 I_49(n_549_1_r_10,blif_clk_net_1_r_6,n4_6,G214_4_l_6,);
not I_50(n12_6,G214_4_l_6);
nor I_51(n4_1_r_6,n28_6,n22_6);
nor I_52(N1_4_r_6,n12_6,n24_6);
nor I_53(n_42_2_l_6,G42_1_r_10,ACVQN2_3_r_10);
DFFARX1 I_54(G214_4_l_6,blif_clk_net_1_r_6,n4_6,P6_5_r_internal_6,);
nand I_55(n19_6,n26_6,n_572_1_r_10);
not I_56(n20_6,n_42_2_l_6);
nor I_57(n21_6,n17_6,n28_6);
and I_58(n22_6,n26_6,n_572_1_r_10);
nand I_59(n23_6,G42_1_r_10,n_572_1_r_10);
nor I_60(n24_6,n17_6,n18_6);
nand I_61(n25_6,n_573_1_r_10,n_42_2_r_10);
endmodule


