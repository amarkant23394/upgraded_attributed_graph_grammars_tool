module test_I3226(I2668,I2702,I1294,I1301,I3226);
input I2668,I2702,I1294,I1301;
output I3226;
wire I3622,I2554,I2866,I3814,I3246,I3797,I3715,I3698,I2572;
DFFARX1 I_0(I2572,I1294,I3246,,,I3622,);
not I_1(I2554,I2866);
DFFARX1 I_2(I1294,,,I2866,);
nand I_3(I3226,I3715,I3814);
nor I_4(I3814,I3622,I3797);
not I_5(I3246,I1301);
not I_6(I3797,I3715);
not I_7(I3715,I3698);
DFFARX1 I_8(I2554,I1294,I3246,,,I3698,);
nor I_9(I2572,I2668,I2702);
endmodule


