module test_I4518(I1477,I2328,I2557,I1470,I2509,I4518);
input I1477,I2328,I2557,I1470,I2509;
output I4518;
wire I2167,I4629,I2173,I4544,I2181,I4869,I2149,I4674,I2155,I2678,I2345,I4691,I2633,I2695;
nand I_0(I2167,I2633,I2328);
nor I_1(I4629,I2167,I2173);
nand I_2(I2173,I2557,I2509);
nand I_3(I4518,I4869,I4691);
not I_4(I4544,I1477);
not I_5(I2181,I1477);
DFFARX1 I_6(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_7(I2695,I1470,I2181,,,I2149,);
DFFARX1 I_8(I2155,I1470,I4544,,,I4674,);
DFFARX1 I_9(I2633,I1470,I2181,,,I2155,);
nand I_10(I2678,I2633);
DFFARX1 I_11(I1470,I2181,,,I2345,);
nor I_12(I4691,I4674,I4629);
DFFARX1 I_13(I1470,I2181,,,I2633,);
and I_14(I2695,I2345,I2678);
endmodule


