module test_I17447(I13908,I15645,I1477,I13758,I13764,I1470,I17447);
input I13908,I15645,I1477,I13758,I13764,I1470;
output I17447;
wire I15662,I13749,I13743,I15832,I16052,I15611,I15679,I15597,I15588,I16145,I16162,I16069,I16086,I15696,I14162,I15628;
nand I_0(I15662,I15645,I13764);
nand I_1(I13749,I14162,I13908);
DFFARX1 I_2(I1470,,,I13743,);
nand I_3(I15832,I15628,I13749);
DFFARX1 I_4(I1470,I15611,,,I16052,);
not I_5(I15611,I1477);
nor I_6(I15679,I15628);
nor I_7(I15597,I15832,I16162);
DFFARX1 I_8(I16086,I1470,I15611,,,I15588,);
not I_9(I16145,I16069);
and I_10(I16162,I15696,I16145);
not I_11(I16069,I16052);
nor I_12(I16086,I16069,I15662);
nand I_13(I15696,I15679,I13758);
DFFARX1 I_14(I1470,,,I14162,);
not I_15(I15628,I13743);
nor I_16(I17447,I15597,I15588);
endmodule


