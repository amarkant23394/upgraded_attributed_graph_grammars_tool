module test_I8998(I5368,I5070,I5642,I6924,I8998);
input I5368,I5070,I5642,I6924;
output I8998;
wire I6992,I6975,I7026,I7057,I6881,I5097;
not I_0(I8998,I6881);
nand I_1(I6992,I6975,I5097);
nor I_2(I6975,I6924,I5070);
not I_3(I7026,I5070);
not I_4(I7057,I7026);
nand I_5(I6881,I6992,I7057);
nand I_6(I5097,I5642,I5368);
endmodule


