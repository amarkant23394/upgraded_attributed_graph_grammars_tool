module test_I9032(I6992,I1477,I7057,I1470,I7221,I5642,I9032);
input I6992,I1477,I7057,I1470,I7221,I5642;
output I9032;
wire I8998,I5105,I7461,I5067,I9015,I6881,I6907,I7269,I6890,I6899,I7444;
not I_0(I8998,I6881);
not I_1(I5105,I1477);
and I_2(I9032,I9015,I6890);
and I_3(I7461,I7221,I7444);
DFFARX1 I_4(I5642,I1470,I5105,,,I5067,);
nor I_5(I9015,I8998,I6899);
nand I_6(I6881,I6992,I7057);
not I_7(I6907,I1477);
DFFARX1 I_8(I5067,I1470,I6907,,,I7269,);
not I_9(I6890,I7269);
DFFARX1 I_10(I7461,I1470,I6907,,,I6899,);
nand I_11(I7444,I6992);
endmodule


