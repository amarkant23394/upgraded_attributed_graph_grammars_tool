module test_I15594(I1477,I15764,I14066,I1470,I13755,I14196,I15594);
input I1477,I15764,I14066,I1470,I13755,I14196;
output I15594;
wire I14083,I13767,I13746,I15815,I13775,I15611,I15798,I15781,I15928;
DFFARX1 I_0(I14066,I1470,I13775,,,I14083,);
DFFARX1 I_1(I14196,I1470,I13775,,,I13767,);
not I_2(I13746,I14083);
DFFARX1 I_3(I15798,I1470,I15611,,,I15815,);
not I_4(I13775,I1477);
not I_5(I15611,I1477);
or I_6(I15594,I15928,I15815);
or I_7(I15798,I15781,I13767);
and I_8(I15781,I15764,I13755);
DFFARX1 I_9(I13746,I1470,I15611,,,I15928,);
endmodule


