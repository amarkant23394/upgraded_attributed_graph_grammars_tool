module test_I1880(I1477,I1470,I1383,I1880);
input I1477,I1470,I1383;
output I1880;
wire I1518;
not I_0(I1518,I1477);
DFFARX1 I_1(I1383,I1470,I1518,,,I1880,);
endmodule


