module test_I14387(I11296,I1477,I11395,I13214,I11290,I11429,I1470,I13409,I14387);
input I11296,I1477,I11395,I13214,I11290,I11429,I1470,I13409;
output I14387;
wire I11768,I13171,I13601,I13186,I13460,I13197,I11299,I13248,I13231,I13426,I11272,I13508,I13491,I11310;
and I_0(I11768,I11429);
nand I_1(I13171,I13248,I13460);
DFFARX1 I_2(I11299,I1470,I13197,,,I13601,);
nor I_3(I13186,I13601,I13508);
not I_4(I13460,I13426);
nand I_5(I14387,I13171,I13186);
not I_6(I13197,I1477);
nor I_7(I11299,I11395,I11429);
DFFARX1 I_8(I13231,I1470,I13197,,,I13248,);
and I_9(I13231,I13214,I11290);
DFFARX1 I_10(I13409,I1470,I13197,,,I13426,);
DFFARX1 I_11(I11768,I1470,I11310,,,I11272,);
and I_12(I13508,I13491,I11272);
DFFARX1 I_13(I11296,I1470,I13197,,,I13491,);
not I_14(I11310,I1477);
endmodule


