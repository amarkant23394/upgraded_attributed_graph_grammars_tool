module test_I17916(I1477,I1470,I17916);
input I1477,I1470;
output I17916;
wire I14083,I13752,I17413,I13746,I15603,I16052,I15611,I15928,I16069;
DFFARX1 I_0(I1470,,,I14083,);
DFFARX1 I_1(I1470,,,I13752,);
not I_2(I17413,I1477);
DFFARX1 I_3(I15603,I1470,I17413,,,I17916,);
not I_4(I13746,I14083);
nor I_5(I15603,I15928,I16069);
DFFARX1 I_6(I13752,I1470,I15611,,,I16052,);
not I_7(I15611,I1477);
DFFARX1 I_8(I13746,I1470,I15611,,,I15928,);
not I_9(I16069,I16052);
endmodule


