module test_I9337(I1477,I1470,I7221,I9337);
input I1477,I1470,I7221;
output I9337;
wire I9320,I7190,I8896,I6875,I6893,I8913,I7156,I6872,I9303,I8862,I6907,I7269,I7286,I6878;
not I_0(I9320,I9303);
DFFARX1 I_1(I7156,I1470,I6907,,,I7190,);
nor I_2(I8896,I6893,I6872);
DFFARX1 I_3(I7221,I1470,I6907,,,I6875,);
nand I_4(I6893,I7156,I7286);
nand I_5(I8913,I8896,I6878);
DFFARX1 I_6(I1470,I6907,,,I7156,);
DFFARX1 I_7(I7269,I1470,I6907,,,I6872,);
DFFARX1 I_8(I6875,I1470,I8862,,,I9303,);
not I_9(I8862,I1477);
not I_10(I6907,I1477);
DFFARX1 I_11(I1470,I6907,,,I7269,);
nor I_12(I9337,I9320,I8913);
nor I_13(I7286,I7269);
not I_14(I6878,I7190);
endmodule


