module test_I13460(I1477,I1470,I11284,I13460);
input I1477,I1470,I11284;
output I13460;
wire I11287,I13392,I11281,I13197,I11593,I13426,I13409;
DFFARX1 I_0(I1470,,,I11287,);
nand I_1(I13392,I11287,I11284);
not I_2(I11281,I11593);
not I_3(I13197,I1477);
DFFARX1 I_4(I1470,,,I11593,);
DFFARX1 I_5(I13409,I1470,I13197,,,I13426,);
not I_6(I13460,I13426);
and I_7(I13409,I13392,I11281);
endmodule


