module test_I3668(I1477,I1215,I1423,I1470,I1535,I3668);
input I1477,I1215,I1423,I1470,I1535;
output I3668;
wire I3388,I1637,I1507,I1586,I1603;
not I_0(I3388,I1477);
not I_1(I1637,I1215);
DFFARX1 I_2(I1507,I1470,I3388,,,I3668,);
nor I_3(I1507,I1603,I1637);
nor I_4(I1586,I1535,I1215);
nand I_5(I1603,I1586,I1423);
endmodule


