module test_I14732(I1477,I1470,I13635,I13525,I13171,I14732);
input I1477,I1470,I13635,I13525,I13171;
output I14732;
wire I14667,I13189,I13601,I13183,I13197,I14404,I14370,I14421,I14650,I13186,I13165,I14387,I14715;
and I_0(I14667,I14650,I13189);
DFFARX1 I_1(I13635,I1470,I13197,,,I13189,);
DFFARX1 I_2(I1470,I13197,,,I13601,);
nand I_3(I13183,I13601,I13525);
not I_4(I13197,I1477);
and I_5(I14404,I14387,I13183);
not I_6(I14370,I1477);
DFFARX1 I_7(I14404,I1470,I14370,,,I14421,);
DFFARX1 I_8(I13165,I1470,I14370,,,I14650,);
nor I_9(I13186,I13601);
DFFARX1 I_10(I1470,I13197,,,I13165,);
nand I_11(I14387,I13171,I13186);
not I_12(I14715,I14667);
nor I_13(I14732,I14421,I14715);
endmodule


