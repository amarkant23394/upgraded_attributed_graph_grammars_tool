module test_I11542(I9320,I1477,I6992,I7026,I1470,I8879,I8964,I11542);
input I9320,I1477,I6992,I7026,I1470,I8879,I8964;
output I11542;
wire I8824,I11491,I8842,I9179,I8827,I8981,I11508,I8862,I6881,I9083,I6896,I8833,I11525;
nand I_0(I8824,I9083,I8981);
not I_1(I11491,I8827);
nor I_2(I8842,I9320,I9083);
DFFARX1 I_3(I6896,I1470,I8862,,,I9179,);
DFFARX1 I_4(I1470,I8862,,,I8827,);
not I_5(I8981,I8964);
nor I_6(I11508,I11491,I8842);
or I_7(I11542,I11525,I8833);
not I_8(I8862,I1477);
nand I_9(I6881,I6992);
nand I_10(I9083,I8879,I6881);
nor I_11(I6896,I6992,I7026);
not I_12(I8833,I9179);
and I_13(I11525,I11508,I8824);
endmodule


