module test_I16007(I13860,I14066,I15832,I12058,I15798,I1470_clk,I1477_rst,I16007);
input I13860,I14066,I15832,I12058,I15798,I1470_clk,I1477_rst;
output I16007;
wire I15880,I13746,I15863,I15928,I13775_rst,I15611_rst,I13761,I11973_rst,I13891,I15713,I15815,I15897,I12075,I14083,I11944;
nor I_0(I15880,I15815,I15863);
not I_1(I13746,I14083);
not I_2(I15863,I15832);
DFFARX1 I_3 (I13746,I1470_clk,I15611_rst,I15928);
not I_4(I13775_rst,I1477_rst);
not I_5(I15611_rst,I1477_rst);
nand I_6(I13761,I13891,I13860);
not I_7(I11973_rst,I1477_rst);
or I_8(I16007,I15928,I15897);
DFFARX1 I_9 (I11944,I1470_clk,I13775_rst,I13891);
not I_10(I15713,I13761);
DFFARX1 I_11 (I15798,I1470_clk,I15611_rst,I15815);
and I_12(I15897,I15713,I15880);
DFFARX1 I_13 (I12058,I1470_clk,I11973_rst,I12075);
DFFARX1 I_14 (I14066,I1470_clk,I13775_rst,I14083);
not I_15(I11944,I12075);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule