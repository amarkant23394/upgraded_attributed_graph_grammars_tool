module test_I3246(I1301,I3246);
input I1301;
output I3246;
wire ;
not I_0(I3246,I1301);
endmodule


