module test_I2781(I1316,I2138,I2005,I1294,I1988,I1301,I2781);
input I1316,I2138,I2005,I1294,I1988,I1301;
output I2781;
wire I2172,I2764,I2344,I1905,I2313,I1937,I2022,I1923,I2155,I1313;
DFFARX1 I_0(I2155,I1294,I1937,,,I2172,);
not I_1(I2764,I1923);
nor I_2(I2781,I2764,I1905);
nor I_3(I2344,I2313,I1988);
DFFARX1 I_4(I2172,I1294,I1937,,,I1905,);
DFFARX1 I_5(I1294,I1937,,,I2313,);
not I_6(I1937,I1301);
nand I_7(I2022,I2005,I1316);
nand I_8(I1923,I2022,I2344);
or I_9(I2155,I2138,I1313);
DFFARX1 I_10(I1294,,,I1313,);
endmodule


