module test_I1637(I1215,I1637);
input I1215;
output I1637;
wire ;
not I_0(I1637,I1215);
endmodule


