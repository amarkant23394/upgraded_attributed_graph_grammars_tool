module test_I3954(I1447,I2946,I3045,I1477,I1470,I3954);
input I1447,I2946,I3045,I1477,I1470;
output I3954;
wire I2759,I2742,I3155,I3076,I2963,I4068,I2724;
not I_0(I2759,I1477);
or I_1(I2742,I3076,I2963);
not I_2(I3954,I4068);
or I_3(I3155,I3076,I3045);
DFFARX1 I_4(I1447,I1470,I2759,,,I3076,);
DFFARX1 I_5(I2946,I1470,I2759,,,I2963,);
nor I_6(I4068,I2742,I2724);
DFFARX1 I_7(I3155,I1470,I2759,,,I2724,);
endmodule


