module test_final(IN_1_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_6_1_l_12,IN_1_5_l_12,IN_2_5_l_12,IN_3_5_l_12,IN_6_5_l_12,blif_clk_net_3_r_13,blif_reset_net_3_r_13,n_429_or_0_3_r_13,G78_3_r_13,n_576_3_r_13,n_102_3_r_13,n_547_3_r_13,G42_4_r_13,n_572_4_r_13,n_573_4_r_13,n_549_4_r_13,n_569_4_r_13,n_452_4_r_13);
input IN_1_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_6_1_l_12,IN_1_5_l_12,IN_2_5_l_12,IN_3_5_l_12,IN_6_5_l_12,blif_clk_net_3_r_13,blif_reset_net_3_r_13;
output n_429_or_0_3_r_13,G78_3_r_13,n_576_3_r_13,n_102_3_r_13,n_547_3_r_13,G42_4_r_13,n_572_4_r_13,n_573_4_r_13,n_549_4_r_13,n_569_4_r_13,n_452_4_r_13;
wire ACVQN2_0_r_12,n_266_and_0_0_r_12,G199_1_r_12,G214_1_r_12,n_429_or_0_3_r_12,G78_3_r_12,n_576_3_r_12,n_102_3_r_12,n_547_3_r_12,n_42_5_r_12,G199_5_r_12,ACVQN2_0_l_12,n_266_and_0_0_l_12,ACVQN1_0_l_12,N1_1_l_12,G199_1_l_12,G214_1_l_12,n3_1_l_12,n_42_5_l_12,N3_5_l_12,G199_5_l_12,n3_5_l_12,ACVQN1_0_r_12,N1_1_r_12,n3_1_r_12,n12_3_r_12,n_431_3_r_12,n11_3_r_12,n13_3_r_12,n14_3_r_12,n15_3_r_12,n16_3_r_12,N3_5_r_12,n3_5_r_12,n2_3_r_13,ACVQN1_2_l_13,P6_2_l_13,P6_internal_2_l_13,n_429_or_0_3_l_13,n12_3_l_13,n_431_3_l_13,G78_3_l_13,n_576_3_l_13,n11_3_l_13,n_102_3_l_13,n_547_3_l_13,n13_3_l_13,n14_3_l_13,n15_3_l_13,n16_3_l_13,n12_3_r_13,n_431_3_r_13,n11_3_r_13,n13_3_r_13,n14_3_r_13,n15_3_r_13,n16_3_r_13,n4_4_r_13,n_87_4_r_13,n7_4_r_13;
DFFARX1 I_0(G199_1_l_12,blif_clk_net_3_r_13,n2_3_r_13,ACVQN2_0_r_12,);
and I_1(n_266_and_0_0_r_12,ACVQN2_0_l_12,ACVQN1_0_r_12);
DFFARX1 I_2(N1_1_r_12,blif_clk_net_3_r_13,n2_3_r_13,G199_1_r_12,);
DFFARX1 I_3(G214_1_l_12,blif_clk_net_3_r_13,n2_3_r_13,G214_1_r_12,);
nand I_4(n_429_or_0_3_r_12,G199_1_l_12,n12_3_r_12);
DFFARX1 I_5(n_431_3_r_12,blif_clk_net_3_r_13,n2_3_r_13,G78_3_r_12,);
nand I_6(n_576_3_r_12,G214_1_l_12,n11_3_r_12);
not I_7(n_102_3_r_12,ACVQN2_0_l_12);
nand I_8(n_547_3_r_12,n_266_and_0_0_l_12,n13_3_r_12);
nor I_9(n_42_5_r_12,n_266_and_0_0_l_12,n_42_5_l_12);
DFFARX1 I_10(N3_5_r_12,blif_clk_net_3_r_13,n2_3_r_13,G199_5_r_12,);
DFFARX1 I_11(IN_1_0_l_12,blif_clk_net_3_r_13,n2_3_r_13,ACVQN2_0_l_12,);
and I_12(n_266_and_0_0_l_12,IN_4_0_l_12,ACVQN1_0_l_12);
DFFARX1 I_13(IN_2_0_l_12,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_0_l_12,);
and I_14(N1_1_l_12,IN_6_1_l_12,n3_1_l_12);
DFFARX1 I_15(N1_1_l_12,blif_clk_net_3_r_13,n2_3_r_13,G199_1_l_12,);
DFFARX1 I_16(IN_3_1_l_12,blif_clk_net_3_r_13,n2_3_r_13,G214_1_l_12,);
nand I_17(n3_1_l_12,IN_1_1_l_12,IN_2_1_l_12);
nor I_18(n_42_5_l_12,IN_1_5_l_12,IN_3_5_l_12);
and I_19(N3_5_l_12,IN_6_5_l_12,n3_5_l_12);
DFFARX1 I_20(N3_5_l_12,blif_clk_net_3_r_13,n2_3_r_13,G199_5_l_12,);
nand I_21(n3_5_l_12,IN_2_5_l_12,IN_3_5_l_12);
DFFARX1 I_22(ACVQN2_0_l_12,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_0_r_12,);
and I_23(N1_1_r_12,G199_1_l_12,n3_1_r_12);
nand I_24(n3_1_r_12,G214_1_l_12,n_42_5_l_12);
not I_25(n12_3_r_12,n_266_and_0_0_l_12);
or I_26(n_431_3_r_12,n_266_and_0_0_l_12,n14_3_r_12);
nor I_27(n11_3_r_12,G199_5_l_12,n12_3_r_12);
nor I_28(n13_3_r_12,ACVQN2_0_l_12,G199_5_l_12);
and I_29(n14_3_r_12,n_42_5_l_12,n15_3_r_12);
nor I_30(n15_3_r_12,G199_5_l_12,n16_3_r_12);
not I_31(n16_3_r_12,G199_1_l_12);
and I_32(N3_5_r_12,ACVQN2_0_l_12,n3_5_r_12);
nand I_33(n3_5_r_12,n_266_and_0_0_l_12,G199_1_l_12);
nand I_34(n_429_or_0_3_r_13,n_429_or_0_3_l_13,n12_3_r_13);
DFFARX1 I_35(n_431_3_r_13,blif_clk_net_3_r_13,n2_3_r_13,G78_3_r_13,);
nand I_36(n_576_3_r_13,n_547_3_l_13,n11_3_r_13);
not I_37(n_102_3_r_13,ACVQN1_2_l_13);
nand I_38(n_547_3_r_13,P6_2_l_13,n13_3_r_13);
DFFARX1 I_39(n4_4_r_13,blif_clk_net_3_r_13,n2_3_r_13,G42_4_r_13,);
nor I_40(n_572_4_r_13,P6_2_l_13,n_429_or_0_3_l_13);
or I_41(n_573_4_r_13,ACVQN1_2_l_13,G78_3_l_13);
nor I_42(n_549_4_r_13,n_429_or_0_3_l_13,n7_4_r_13);
or I_43(n_569_4_r_13,n_429_or_0_3_l_13,G78_3_l_13);
nor I_44(n_452_4_r_13,ACVQN1_2_l_13,P6_2_l_13);
not I_45(n2_3_r_13,blif_reset_net_3_r_13);
DFFARX1 I_46(n_547_3_r_12,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_2_l_13,);
not I_47(P6_2_l_13,P6_internal_2_l_13);
DFFARX1 I_48(n_42_5_r_12,blif_clk_net_3_r_13,n2_3_r_13,P6_internal_2_l_13,);
nand I_49(n_429_or_0_3_l_13,n12_3_l_13,G199_5_r_12);
not I_50(n12_3_l_13,G214_1_r_12);
or I_51(n_431_3_l_13,n14_3_l_13,ACVQN2_0_r_12);
DFFARX1 I_52(n_431_3_l_13,blif_clk_net_3_r_13,n2_3_r_13,G78_3_l_13,);
nand I_53(n_576_3_l_13,n11_3_l_13,G78_3_r_12);
nor I_54(n11_3_l_13,n12_3_l_13,n_429_or_0_3_r_12);
not I_55(n_102_3_l_13,n_429_or_0_3_r_12);
nand I_56(n_547_3_l_13,n13_3_l_13,G199_1_r_12);
nor I_57(n13_3_l_13,n_429_or_0_3_r_12,n_102_3_r_12);
and I_58(n14_3_l_13,n15_3_l_13,n_266_and_0_0_r_12);
nor I_59(n15_3_l_13,n16_3_l_13,n_576_3_r_12);
not I_60(n16_3_l_13,G199_5_r_12);
not I_61(n12_3_r_13,n_102_3_l_13);
or I_62(n_431_3_r_13,ACVQN1_2_l_13,n14_3_r_13);
nor I_63(n11_3_r_13,ACVQN1_2_l_13,n12_3_r_13);
nor I_64(n13_3_r_13,ACVQN1_2_l_13,n_576_3_l_13);
and I_65(n14_3_r_13,n_102_3_l_13,n15_3_r_13);
nor I_66(n15_3_r_13,G78_3_l_13,n16_3_r_13);
not I_67(n16_3_r_13,n_429_or_0_3_l_13);
nor I_68(n4_4_r_13,P6_2_l_13,n_547_3_l_13);
not I_69(n_87_4_r_13,P6_2_l_13);
and I_70(n7_4_r_13,n_576_3_l_13,n_87_4_r_13);
endmodule


