module test_I8187(I6265,I1477,I5785,I1470,I8187);
input I6265,I1477,I5785,I1470;
output I8187;
wire I8233,I8216,I5751,I5802,I8298,I5719,I5740,I8315,I5722;
DFFARX1 I_0(I8315,I1470,I8216,,,I8187,);
not I_1(I8233,I5722);
not I_2(I8216,I1477);
not I_3(I5751,I1477);
DFFARX1 I_4(I5785,I1470,I5751,,,I5802,);
nor I_5(I8298,I8233,I5719);
DFFARX1 I_6(I6265,I1470,I5751,,,I5719,);
not I_7(I5740,I5802);
nand I_8(I8315,I8298,I5740);
DFFARX1 I_9(I1470,I5751,,,I5722,);
endmodule


