module test_I16801(I14999,I1477,I1470,I15126,I15423,I15502,I16801);
input I14999,I1477,I1470,I15126,I15423,I15502;
output I16801;
wire I14948,I15016,I15211,I14951,I15519,I14965,I15245,I12581,I16886;
DFFARX1 I_0(I15519,I1470,I14965,,,I14948,);
nand I_1(I15016,I14999,I12581);
DFFARX1 I_2(I1470,I14965,,,I15211,);
nand I_3(I14951,I15016,I15245);
not I_4(I16801,I16886);
or I_5(I15519,I15502,I15423);
not I_6(I14965,I1477);
nor I_7(I15245,I15211,I15126);
DFFARX1 I_8(I1470,,,I12581,);
nor I_9(I16886,I14951,I14948);
endmodule


