module test_I12848(I11232,I10797,I1477,I1470,I10732,I12848);
input I11232,I10797,I1477,I1470,I10732;
output I12848;
wire I12619,I10647,I12831,I10624,I10618,I12814,I10896,I10621,I10930;
not I_0(I12619,I1477);
not I_1(I10647,I1477);
and I_2(I12831,I12814,I10618);
DFFARX1 I_3(I11232,I1470,I10647,,,I10624,);
not I_4(I10618,I10930);
nand I_5(I12814,I10624,I10621);
DFFARX1 I_6(I1470,I10647,,,I10896,);
nand I_7(I10621,I10732,I10797);
DFFARX1 I_8(I12831,I1470,I12619,,,I12848,);
DFFARX1 I_9(I10896,I1470,I10647,,,I10930,);
endmodule


