module test_I15815(I14179,I15747,I1477,I13925,I1470,I15815);
input I14179,I15747,I1477,I13925,I1470;
output I15815;
wire I13767,I14004,I15764,I13737,I13775,I15611,I15781,I13755,I15798,I14196;
DFFARX1 I_0(I14196,I1470,I13775,,,I13767,);
DFFARX1 I_1(I1470,I13775,,,I14004,);
nor I_2(I15764,I15747,I13737);
DFFARX1 I_3(I15798,I1470,I15611,,,I15815,);
DFFARX1 I_4(I1470,I13775,,,I13737,);
not I_5(I13775,I1477);
not I_6(I15611,I1477);
and I_7(I15781,I15764,I13755);
nand I_8(I13755,I14004,I13925);
or I_9(I15798,I15781,I13767);
and I_10(I14196,I14004,I14179);
endmodule


