module test_I2946(I1415,I1391,I1263,I1311,I2946);
input I1415,I1391,I1263,I1311;
output I2946;
wire I2929,I2895,I2912;
or I_0(I2946,I2929,I1263);
and I_1(I2929,I2912,I1391);
not I_2(I2895,I1415);
nor I_3(I2912,I2895,I1311);
endmodule


