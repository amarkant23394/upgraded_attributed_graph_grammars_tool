module test_I13749(I1477,I1470,I11990,I13749);
input I1477,I1470,I11990;
output I13749;
wire I13908,I12270,I12239,I14162,I10014,I11938,I12208,I13775,I13891,I11973,I12075,I11944;
not I_0(I13908,I13891);
nand I_1(I12270,I11990,I10014);
DFFARX1 I_2(I12208,I1470,I11973,,,I12239,);
DFFARX1 I_3(I11938,I1470,I13775,,,I14162,);
DFFARX1 I_4(I1470,,,I10014,);
and I_5(I11938,I12270,I12239);
DFFARX1 I_6(I1470,I11973,,,I12208,);
nand I_7(I13749,I14162,I13908);
not I_8(I13775,I1477);
DFFARX1 I_9(I11944,I1470,I13775,,,I13891,);
not I_10(I11973,I1477);
DFFARX1 I_11(I1470,I11973,,,I12075,);
not I_12(I11944,I12075);
endmodule


