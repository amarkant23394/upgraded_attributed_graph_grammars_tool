module test_final(IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_7_r_16,blif_reset_net_7_r_16,N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16);
input IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_7_r_16,blif_reset_net_7_r_16;
output N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16;
wire N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_573_7_r_12,n_549_7_r_12,n_569_7_r_12,n_452_7_r_12,N6147_9_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12,n_549_7_r_16,N3_8_l_16,n8_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16;
nor I_0(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_1(N1508_0_r_12,n30_12,n37_12);
nor I_2(N1507_6_r_12,n25_12,n39_12);
nor I_3(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_4(n1_12,blif_clk_net_7_r_16,n8_16,G42_7_r_12,);
nor I_5(n_572_7_r_12,n23_12,n24_12);
nand I_6(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_7(n_549_7_r_12,n27_12,n28_12);
nand I_8(n_569_7_r_12,n25_12,n26_12);
nand I_9(n_452_7_r_12,IN_1_1_l_12,IN_2_1_l_12);
nand I_10(N6147_9_r_12,n30_12,n31_12);
nor I_11(N6134_9_r_12,n35_12,n36_12);
not I_12(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_13(n1_12,n_573_7_r_12);
not I_14(n23_12,n36_12);
nor I_15(n24_12,IN_3_1_l_12,n_452_7_r_12);
nand I_16(n25_12,n23_12,n40_12);
not I_17(n26_12,n35_12);
not I_18(n27_12,N6134_9_r_12);
nand I_19(n28_12,n26_12,n29_12);
not I_20(n29_12,n24_12);
nand I_21(n30_12,n33_12,n41_12);
nand I_22(n31_12,n32_12,n33_12);
nor I_23(n32_12,n26_12,n34_12);
nor I_24(n33_12,IN_1_2_l_12,IN_2_2_l_12);
nor I_25(n34_12,IN_5_2_l_12,n42_12);
nor I_26(n35_12,IN_1_3_l_12,n38_12);
nand I_27(n36_12,IN_1_10_l_12,IN_2_10_l_12);
nand I_28(n37_12,n23_12,n35_12);
or I_29(n38_12,IN_2_3_l_12,IN_3_3_l_12);
not I_30(n39_12,n30_12);
or I_31(n40_12,IN_3_10_l_12,IN_4_10_l_12);
nor I_32(n41_12,n34_12,n36_12);
nor I_33(n42_12,IN_3_2_l_12,IN_4_2_l_12);
nor I_34(N1371_0_r_16,n35_16,n39_16);
nor I_35(N1508_0_r_16,n39_16,n46_16);
not I_36(N1372_1_r_16,n45_16);
nor I_37(N1508_1_r_16,n53_16,n45_16);
nor I_38(N6147_2_r_16,n37_16,n38_16);
nor I_39(N1507_6_r_16,n44_16,n49_16);
nor I_40(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_41(n4_7_r_16,blif_clk_net_7_r_16,n8_16,G42_7_r_16,);
nor I_42(n_572_7_r_16,n32_16,n33_16);
nand I_43(n_573_7_r_16,n30_16,n31_16);
nand I_44(n_549_7_r_16,n47_16,n_569_7_r_12);
nand I_45(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_46(n_452_7_r_16,n34_16,n35_16);
and I_47(N3_8_l_16,n41_16,N6147_9_r_12);
not I_48(n8_16,blif_reset_net_7_r_16);
DFFARX1 I_49(N3_8_l_16,blif_clk_net_7_r_16,n8_16,n53_16,);
not I_50(n29_16,n53_16);
nor I_51(n4_7_r_16,n35_16,n36_16);
nand I_52(n30_16,N1371_0_r_12,N1508_0_r_12);
not I_53(n31_16,n34_16);
nor I_54(n32_16,n30_16,G42_7_r_12);
not I_55(n33_16,n_549_7_r_16);
nor I_56(n34_16,n48_16,n_572_7_r_12);
and I_57(n35_16,n50_16,n_549_7_r_12);
not I_58(n36_16,n30_16);
nor I_59(n37_16,n31_16,n40_16);
nand I_60(n38_16,n29_16,n39_16);
not I_61(n39_16,n32_16);
nor I_62(n40_16,N1507_6_r_12,N1508_6_r_12);
nand I_63(n41_16,N1507_6_r_12,G42_7_r_12);
nand I_64(n42_16,n35_16,n43_16);
not I_65(n43_16,n44_16);
nor I_66(n44_16,n32_16,n49_16);
nand I_67(n45_16,n36_16,n40_16);
nor I_68(n46_16,n33_16,n34_16);
nand I_69(n47_16,N1508_0_r_12,n_572_7_r_12);
or I_70(n48_16,N1508_6_r_12,N1507_6_r_12);
and I_71(n49_16,n35_16,n36_16);
and I_72(n50_16,n51_16,N1371_0_r_12);
nand I_73(n51_16,n47_16,n52_16);
not I_74(n52_16,n_569_7_r_12);
endmodule


