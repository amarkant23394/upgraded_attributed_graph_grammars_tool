module test_I11953(I10349,I10538,I1477,I1470,I10120,I11953);
input I10349,I10538,I1477,I1470,I10120;
output I11953;
wire I12541,I10038,I12425,I12349,I10041,I12524,I12442,I11973;
nor I_0(I12541,I12349,I12524);
nand I_1(I10038,I10349,I10538);
DFFARX1 I_2(I10038,I1470,I11973,,,I12425,);
nand I_3(I11953,I12442,I12541);
DFFARX1 I_4(I10041,I1470,I11973,,,I12349,);
nor I_5(I10041,I10349,I10120);
not I_6(I12524,I12442);
not I_7(I12442,I12425);
not I_8(I11973,I1477);
endmodule


