module test_final(IN_1_0_l_9,IN_2_0_l_9,IN_4_0_l_9,G18_4_l_9,G15_4_l_9,IN_1_4_l_9,IN_4_4_l_9,IN_5_4_l_9,IN_7_4_l_9,IN_9_4_l_9,IN_10_4_l_9,blif_clk_net_3_r_0,blif_reset_net_3_r_0,n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0);
input IN_1_0_l_9,IN_2_0_l_9,IN_4_0_l_9,G18_4_l_9,G15_4_l_9,IN_1_4_l_9,IN_4_4_l_9,IN_5_4_l_9,IN_7_4_l_9,IN_9_4_l_9,IN_10_4_l_9,blif_clk_net_3_r_0,blif_reset_net_3_r_0;
output n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0;
wire G199_1_r_9,G214_1_r_9,ACVQN1_2_r_9,P6_2_r_9,n_429_or_0_3_r_9,G78_3_r_9,n_576_3_r_9,n_102_3_r_9,n_547_3_r_9,n_42_5_r_9,G199_5_r_9,ACVQN2_0_l_9,n_266_and_0_0_l_9,ACVQN1_0_l_9,n4_4_l_9,G42_4_l_9,n_87_4_l_9,n_572_4_l_9,n_573_4_l_9,n_549_4_l_9,n7_4_l_9,n_569_4_l_9,n_452_4_l_9,N1_1_r_9,n3_1_r_9,P6_internal_2_r_9,n12_3_r_9,n_431_3_r_9,n11_3_r_9,n13_3_r_9,n14_3_r_9,n15_3_r_9,n16_3_r_9,N3_5_r_9,n3_5_r_9,n2_3_r_0,ACVQN2_0_l_0,n_266_and_0_0_l_0,ACVQN1_0_l_0,N1_1_l_0,G199_1_l_0,G214_1_l_0,n3_1_l_0,n_42_5_l_0,N3_5_l_0,G199_5_l_0,n3_5_l_0,n12_3_r_0,n_431_3_r_0,n11_3_r_0,n13_3_r_0,n14_3_r_0,n15_3_r_0,n16_3_r_0,n4_4_r_0,n_87_4_r_0,n7_4_r_0;
DFFARX1 I_0(N1_1_r_9,blif_clk_net_3_r_0,n2_3_r_0,G199_1_r_9,);
DFFARX1 I_1(G42_4_l_9,blif_clk_net_3_r_0,n2_3_r_0,G214_1_r_9,);
DFFARX1 I_2(n_572_4_l_9,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_2_r_9,);
not I_3(P6_2_r_9,P6_internal_2_r_9);
nand I_4(n_429_or_0_3_r_9,n_572_4_l_9,n12_3_r_9);
DFFARX1 I_5(n_431_3_r_9,blif_clk_net_3_r_0,n2_3_r_0,G78_3_r_9,);
nand I_6(n_576_3_r_9,n_573_4_l_9,n11_3_r_9);
not I_7(n_102_3_r_9,n_266_and_0_0_l_9);
nand I_8(n_547_3_r_9,n_549_4_l_9,n13_3_r_9);
nor I_9(n_42_5_r_9,n_569_4_l_9,n_452_4_l_9);
DFFARX1 I_10(N3_5_r_9,blif_clk_net_3_r_0,n2_3_r_0,G199_5_r_9,);
DFFARX1 I_11(IN_1_0_l_9,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_l_9,);
and I_12(n_266_and_0_0_l_9,IN_4_0_l_9,ACVQN1_0_l_9);
DFFARX1 I_13(IN_2_0_l_9,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_l_9,);
nor I_14(n4_4_l_9,G18_4_l_9,IN_1_4_l_9);
DFFARX1 I_15(n4_4_l_9,blif_clk_net_3_r_0,n2_3_r_0,G42_4_l_9,);
not I_16(n_87_4_l_9,G15_4_l_9);
nor I_17(n_572_4_l_9,G15_4_l_9,IN_7_4_l_9);
or I_18(n_573_4_l_9,IN_5_4_l_9,IN_9_4_l_9);
nor I_19(n_549_4_l_9,IN_10_4_l_9,n7_4_l_9);
and I_20(n7_4_l_9,IN_4_4_l_9,n_87_4_l_9);
or I_21(n_569_4_l_9,IN_9_4_l_9,IN_10_4_l_9);
nor I_22(n_452_4_l_9,G18_4_l_9,IN_5_4_l_9);
and I_23(N1_1_r_9,n_266_and_0_0_l_9,n3_1_r_9);
nand I_24(n3_1_r_9,n_572_4_l_9,n_569_4_l_9);
DFFARX1 I_25(n_266_and_0_0_l_9,blif_clk_net_3_r_0,n2_3_r_0,P6_internal_2_r_9,);
not I_26(n12_3_r_9,G42_4_l_9);
or I_27(n_431_3_r_9,n_549_4_l_9,n14_3_r_9);
nor I_28(n11_3_r_9,ACVQN2_0_l_9,n12_3_r_9);
nor I_29(n13_3_r_9,ACVQN2_0_l_9,n_266_and_0_0_l_9);
and I_30(n14_3_r_9,n_452_4_l_9,n15_3_r_9);
nor I_31(n15_3_r_9,G42_4_l_9,n16_3_r_9);
not I_32(n16_3_r_9,n_572_4_l_9);
and I_33(N3_5_r_9,ACVQN2_0_l_9,n3_5_r_9);
nand I_34(n3_5_r_9,n_573_4_l_9,n_452_4_l_9);
nand I_35(n_429_or_0_3_r_0,ACVQN2_0_l_0,n12_3_r_0);
DFFARX1 I_36(n_431_3_r_0,blif_clk_net_3_r_0,n2_3_r_0,G78_3_r_0,);
nand I_37(n_576_3_r_0,n_266_and_0_0_l_0,n11_3_r_0);
not I_38(n_102_3_r_0,n_42_5_l_0);
nand I_39(n_547_3_r_0,ACVQN2_0_l_0,n13_3_r_0);
DFFARX1 I_40(n4_4_r_0,blif_clk_net_3_r_0,n2_3_r_0,G42_4_r_0,);
nor I_41(n_572_4_r_0,G199_1_l_0,G199_5_l_0);
or I_42(n_573_4_r_0,n_42_5_l_0,G199_5_l_0);
nor I_43(n_549_4_r_0,n_266_and_0_0_l_0,n7_4_r_0);
or I_44(n_569_4_r_0,n_266_and_0_0_l_0,n_42_5_l_0);
nor I_45(n_452_4_r_0,ACVQN2_0_l_0,G199_5_l_0);
not I_46(n2_3_r_0,blif_reset_net_3_r_0);
DFFARX1 I_47(n_547_3_r_9,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_l_0,);
and I_48(n_266_and_0_0_l_0,ACVQN1_0_l_0,G199_1_r_9);
DFFARX1 I_49(n_42_5_r_9,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_l_0,);
and I_50(N1_1_l_0,n3_1_l_0,n_576_3_r_9);
DFFARX1 I_51(N1_1_l_0,blif_clk_net_3_r_0,n2_3_r_0,G199_1_l_0,);
DFFARX1 I_52(G78_3_r_9,blif_clk_net_3_r_0,n2_3_r_0,G214_1_l_0,);
nand I_53(n3_1_l_0,G214_1_r_9,P6_2_r_9);
nor I_54(n_42_5_l_0,ACVQN1_2_r_9,n_429_or_0_3_r_9);
and I_55(N3_5_l_0,n3_5_l_0,n_102_3_r_9);
DFFARX1 I_56(N3_5_l_0,blif_clk_net_3_r_0,n2_3_r_0,G199_5_l_0,);
nand I_57(n3_5_l_0,n_429_or_0_3_r_9,G199_5_r_9);
not I_58(n12_3_r_0,G199_1_l_0);
or I_59(n_431_3_r_0,n_266_and_0_0_l_0,n14_3_r_0);
nor I_60(n11_3_r_0,G214_1_l_0,n12_3_r_0);
nor I_61(n13_3_r_0,G214_1_l_0,n_42_5_l_0);
and I_62(n14_3_r_0,n_42_5_l_0,n15_3_r_0);
nor I_63(n15_3_r_0,G199_1_l_0,n16_3_r_0);
not I_64(n16_3_r_0,ACVQN2_0_l_0);
nor I_65(n4_4_r_0,ACVQN2_0_l_0,G214_1_l_0);
not I_66(n_87_4_r_0,G199_5_l_0);
and I_67(n7_4_r_0,ACVQN2_0_l_0,n_87_4_r_0);
endmodule


