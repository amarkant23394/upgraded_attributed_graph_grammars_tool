module test_I3380(I1477,I1849,I1897,I1492,I2038,I1470,I3380);
input I1477,I1849,I1897,I1492,I2038,I1470;
output I3380;
wire I1486,I1801,I3521,I3504,I1495,I3538,I3487,I3747,I3388,I3846,I1489,I1510,I1767,I1518,I1504,I3555,I2103;
DFFARX1 I_0(I1470,I1518,,,I1486,);
DFFARX1 I_1(I1767,I1470,I1518,,,I1801,);
nor I_2(I3521,I3504,I1495);
and I_3(I3504,I3487,I1489);
DFFARX1 I_4(I2103,I1470,I1518,,,I1495,);
nor I_5(I3538,I1492,I1510);
not I_6(I3487,I1486);
DFFARX1 I_7(I1504,I1470,I3388,,,I3747,);
not I_8(I3388,I1477);
nor I_9(I3846,I3747,I3555);
not I_10(I1489,I1801);
DFFARX1 I_11(I1470,I1518,,,I1510,);
DFFARX1 I_12(I1470,I1518,,,I1767,);
not I_13(I1518,I1477);
nand I_14(I1504,I1767,I1897);
nand I_15(I3380,I3521,I3846);
DFFARX1 I_16(I3538,I1470,I3388,,,I3555,);
or I_17(I2103,I2038,I1849);
endmodule


