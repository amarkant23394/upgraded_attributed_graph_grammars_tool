module test_final(IN_1_2_l_5,IN_2_2_l_5,G1_3_l_5,G2_3_l_5,IN_2_3_l_5,IN_4_3_l_5,IN_5_3_l_5,IN_7_3_l_5,IN_8_3_l_5,IN_10_3_l_5,IN_11_3_l_5,blif_clk_net_3_r_13,blif_reset_net_3_r_13,n_429_or_0_3_r_13,G78_3_r_13,n_576_3_r_13,n_102_3_r_13,n_547_3_r_13,G42_4_r_13,n_572_4_r_13,n_573_4_r_13,n_549_4_r_13,n_569_4_r_13,n_452_4_r_13);
input IN_1_2_l_5,IN_2_2_l_5,G1_3_l_5,G2_3_l_5,IN_2_3_l_5,IN_4_3_l_5,IN_5_3_l_5,IN_7_3_l_5,IN_8_3_l_5,IN_10_3_l_5,IN_11_3_l_5,blif_clk_net_3_r_13,blif_reset_net_3_r_13;
output n_429_or_0_3_r_13,G78_3_r_13,n_576_3_r_13,n_102_3_r_13,n_547_3_r_13,G42_4_r_13,n_572_4_r_13,n_573_4_r_13,n_549_4_r_13,n_569_4_r_13,n_452_4_r_13;
wire G199_1_r_5,G214_1_r_5,ACVQN1_2_r_5,P6_2_r_5,n_429_or_0_3_r_5,G78_3_r_5,n_576_3_r_5,n_102_3_r_5,n_547_3_r_5,n_42_5_r_5,G199_5_r_5,ACVQN1_2_l_5,P6_2_l_5,P6_internal_2_l_5,n_429_or_0_3_l_5,n12_3_l_5,n_431_3_l_5,G78_3_l_5,n_576_3_l_5,n11_3_l_5,n_102_3_l_5,n_547_3_l_5,n13_3_l_5,n14_3_l_5,n15_3_l_5,n16_3_l_5,N1_1_r_5,n3_1_r_5,P6_internal_2_r_5,n12_3_r_5,n_431_3_r_5,n11_3_r_5,n13_3_r_5,n14_3_r_5,n15_3_r_5,n16_3_r_5,N3_5_r_5,n3_5_r_5,n2_3_r_13,ACVQN1_2_l_13,P6_2_l_13,P6_internal_2_l_13,n_429_or_0_3_l_13,n12_3_l_13,n_431_3_l_13,G78_3_l_13,n_576_3_l_13,n11_3_l_13,n_102_3_l_13,n_547_3_l_13,n13_3_l_13,n14_3_l_13,n15_3_l_13,n16_3_l_13,n12_3_r_13,n_431_3_r_13,n11_3_r_13,n13_3_r_13,n14_3_r_13,n15_3_r_13,n16_3_r_13,n4_4_r_13,n_87_4_r_13,n7_4_r_13;
DFFARX1 I_0(N1_1_r_5,blif_clk_net_3_r_13,n2_3_r_13,G199_1_r_5,);
DFFARX1 I_1(ACVQN1_2_l_5,blif_clk_net_3_r_13,n2_3_r_13,G214_1_r_5,);
DFFARX1 I_2(n_429_or_0_3_l_5,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_2_r_5,);
not I_3(P6_2_r_5,P6_internal_2_r_5);
nand I_4(n_429_or_0_3_r_5,n_576_3_l_5,n12_3_r_5);
DFFARX1 I_5(n_431_3_r_5,blif_clk_net_3_r_13,n2_3_r_13,G78_3_r_5,);
nand I_6(n_576_3_r_5,P6_2_l_5,n11_3_r_5);
not I_7(n_102_3_r_5,ACVQN1_2_l_5);
nand I_8(n_547_3_r_5,G78_3_l_5,n13_3_r_5);
nor I_9(n_42_5_r_5,n_576_3_l_5,n_102_3_l_5);
DFFARX1 I_10(N3_5_r_5,blif_clk_net_3_r_13,n2_3_r_13,G199_5_r_5,);
DFFARX1 I_11(IN_2_2_l_5,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_2_l_5,);
not I_12(P6_2_l_5,P6_internal_2_l_5);
DFFARX1 I_13(IN_1_2_l_5,blif_clk_net_3_r_13,n2_3_r_13,P6_internal_2_l_5,);
nand I_14(n_429_or_0_3_l_5,G1_3_l_5,n12_3_l_5);
not I_15(n12_3_l_5,IN_5_3_l_5);
or I_16(n_431_3_l_5,IN_8_3_l_5,n14_3_l_5);
DFFARX1 I_17(n_431_3_l_5,blif_clk_net_3_r_13,n2_3_r_13,G78_3_l_5,);
nand I_18(n_576_3_l_5,IN_7_3_l_5,n11_3_l_5);
nor I_19(n11_3_l_5,G2_3_l_5,n12_3_l_5);
not I_20(n_102_3_l_5,G2_3_l_5);
nand I_21(n_547_3_l_5,IN_11_3_l_5,n13_3_l_5);
nor I_22(n13_3_l_5,G2_3_l_5,IN_10_3_l_5);
and I_23(n14_3_l_5,IN_2_3_l_5,n15_3_l_5);
nor I_24(n15_3_l_5,IN_4_3_l_5,n16_3_l_5);
not I_25(n16_3_l_5,G1_3_l_5);
and I_26(N1_1_r_5,n_102_3_l_5,n3_1_r_5);
nand I_27(n3_1_r_5,ACVQN1_2_l_5,n_547_3_l_5);
DFFARX1 I_28(G78_3_l_5,blif_clk_net_3_r_13,n2_3_r_13,P6_internal_2_r_5,);
not I_29(n12_3_r_5,n_102_3_l_5);
or I_30(n_431_3_r_5,P6_2_l_5,n14_3_r_5);
nor I_31(n11_3_r_5,ACVQN1_2_l_5,n12_3_r_5);
nor I_32(n13_3_r_5,ACVQN1_2_l_5,n_576_3_l_5);
and I_33(n14_3_r_5,n_429_or_0_3_l_5,n15_3_r_5);
nor I_34(n15_3_r_5,G78_3_l_5,n16_3_r_5);
not I_35(n16_3_r_5,n_576_3_l_5);
and I_36(N3_5_r_5,n_429_or_0_3_l_5,n3_5_r_5);
nand I_37(n3_5_r_5,P6_2_l_5,n_576_3_l_5);
nand I_38(n_429_or_0_3_r_13,n_429_or_0_3_l_13,n12_3_r_13);
DFFARX1 I_39(n_431_3_r_13,blif_clk_net_3_r_13,n2_3_r_13,G78_3_r_13,);
nand I_40(n_576_3_r_13,n_547_3_l_13,n11_3_r_13);
not I_41(n_102_3_r_13,ACVQN1_2_l_13);
nand I_42(n_547_3_r_13,P6_2_l_13,n13_3_r_13);
DFFARX1 I_43(n4_4_r_13,blif_clk_net_3_r_13,n2_3_r_13,G42_4_r_13,);
nor I_44(n_572_4_r_13,P6_2_l_13,n_429_or_0_3_l_13);
or I_45(n_573_4_r_13,ACVQN1_2_l_13,G78_3_l_13);
nor I_46(n_549_4_r_13,n_429_or_0_3_l_13,n7_4_r_13);
or I_47(n_569_4_r_13,n_429_or_0_3_l_13,G78_3_l_13);
nor I_48(n_452_4_r_13,ACVQN1_2_l_13,P6_2_l_13);
not I_49(n2_3_r_13,blif_reset_net_3_r_13);
DFFARX1 I_50(n_42_5_r_5,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_2_l_13,);
not I_51(P6_2_l_13,P6_internal_2_l_13);
DFFARX1 I_52(ACVQN1_2_r_5,blif_clk_net_3_r_13,n2_3_r_13,P6_internal_2_l_13,);
nand I_53(n_429_or_0_3_l_13,n12_3_l_13,n_429_or_0_3_r_5);
not I_54(n12_3_l_13,n_576_3_r_5);
or I_55(n_431_3_l_13,n14_3_l_13,G199_1_r_5);
DFFARX1 I_56(n_431_3_l_13,blif_clk_net_3_r_13,n2_3_r_13,G78_3_l_13,);
nand I_57(n_576_3_l_13,n11_3_l_13,G78_3_r_5);
nor I_58(n11_3_l_13,n12_3_l_13,n_547_3_r_5);
not I_59(n_102_3_l_13,n_547_3_r_5);
nand I_60(n_547_3_l_13,n13_3_l_13,P6_2_r_5);
nor I_61(n13_3_l_13,G214_1_r_5,n_547_3_r_5);
and I_62(n14_3_l_13,n15_3_l_13,n_102_3_r_5);
nor I_63(n15_3_l_13,n16_3_l_13,G199_5_r_5);
not I_64(n16_3_l_13,n_429_or_0_3_r_5);
not I_65(n12_3_r_13,n_102_3_l_13);
or I_66(n_431_3_r_13,ACVQN1_2_l_13,n14_3_r_13);
nor I_67(n11_3_r_13,ACVQN1_2_l_13,n12_3_r_13);
nor I_68(n13_3_r_13,ACVQN1_2_l_13,n_576_3_l_13);
and I_69(n14_3_r_13,n_102_3_l_13,n15_3_r_13);
nor I_70(n15_3_r_13,G78_3_l_13,n16_3_r_13);
not I_71(n16_3_r_13,n_429_or_0_3_l_13);
nor I_72(n4_4_r_13,P6_2_l_13,n_547_3_l_13);
not I_73(n_87_4_r_13,P6_2_l_13);
and I_74(n7_4_r_13,n_576_3_l_13,n_87_4_r_13);
endmodule


