module test_I1492(I1423,I1215,I1455,I1492);
input I1423,I1215,I1455;
output I1492;
wire I1603,I1637,I1586,I1535,I1668;
nand I_0(I1492,I1603,I1668);
nand I_1(I1603,I1586,I1423);
not I_2(I1637,I1215);
nor I_3(I1586,I1535,I1215);
not I_4(I1535,I1455);
not I_5(I1668,I1637);
endmodule


