module test_final(IN_1_0_l_0,IN_2_0_l_0,IN_4_0_l_0,IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_6_1_l_0,IN_1_5_l_0,IN_2_5_l_0,IN_3_5_l_0,IN_6_5_l_0,blif_reset_net_0_r_14,blif_clk_net_0_r_14,ACVQN2_0_r_14,n_266_and_0_0_r_14,G199_1_r_14,G214_1_r_14,ACVQN1_2_r_14,P6_2_r_14,n_429_or_0_3_r_14,G78_3_r_14,n_576_3_r_14,n_102_3_r_14,n_547_3_r_14);
input IN_1_0_l_0,IN_2_0_l_0,IN_4_0_l_0,IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_6_1_l_0,IN_1_5_l_0,IN_2_5_l_0,IN_3_5_l_0,IN_6_5_l_0,blif_reset_net_0_r_14,blif_clk_net_0_r_14;
output ACVQN2_0_r_14,n_266_and_0_0_r_14,G199_1_r_14,G214_1_r_14,ACVQN1_2_r_14,P6_2_r_14,n_429_or_0_3_r_14,G78_3_r_14,n_576_3_r_14,n_102_3_r_14,n_547_3_r_14;
wire n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0,ACVQN2_0_l_0,n_266_and_0_0_l_0,ACVQN1_0_l_0,N1_1_l_0,G199_1_l_0,G214_1_l_0,n3_1_l_0,n_42_5_l_0,N3_5_l_0,G199_5_l_0,n3_5_l_0,n12_3_r_0,n_431_3_r_0,n11_3_r_0,n13_3_r_0,n14_3_r_0,n15_3_r_0,n16_3_r_0,n4_4_r_0,n_87_4_r_0,n7_4_r_0,n1_0_r_14,ACVQN2_0_l_14,n_266_and_0_0_l_14,ACVQN1_0_l_14,N1_1_l_14,G199_1_l_14,G214_1_l_14,n3_1_l_14,n_42_5_l_14,N3_5_l_14,G199_5_l_14,n3_5_l_14,ACVQN1_0_r_14,N1_1_r_14,n3_1_r_14,P6_internal_2_r_14,n12_3_r_14,n_431_3_r_14,n11_3_r_14,n13_3_r_14,n14_3_r_14,n15_3_r_14,n16_3_r_14;
nand I_0(n_429_or_0_3_r_0,ACVQN2_0_l_0,n12_3_r_0);
DFFARX1 I_1(n_431_3_r_0,blif_clk_net_0_r_14,n1_0_r_14,G78_3_r_0,);
nand I_2(n_576_3_r_0,n_266_and_0_0_l_0,n11_3_r_0);
not I_3(n_102_3_r_0,n_42_5_l_0);
nand I_4(n_547_3_r_0,ACVQN2_0_l_0,n13_3_r_0);
DFFARX1 I_5(n4_4_r_0,blif_clk_net_0_r_14,n1_0_r_14,G42_4_r_0,);
nor I_6(n_572_4_r_0,G199_1_l_0,G199_5_l_0);
or I_7(n_573_4_r_0,n_42_5_l_0,G199_5_l_0);
nor I_8(n_549_4_r_0,n_266_and_0_0_l_0,n7_4_r_0);
or I_9(n_569_4_r_0,n_266_and_0_0_l_0,n_42_5_l_0);
nor I_10(n_452_4_r_0,ACVQN2_0_l_0,G199_5_l_0);
DFFARX1 I_11(IN_1_0_l_0,blif_clk_net_0_r_14,n1_0_r_14,ACVQN2_0_l_0,);
and I_12(n_266_and_0_0_l_0,IN_4_0_l_0,ACVQN1_0_l_0);
DFFARX1 I_13(IN_2_0_l_0,blif_clk_net_0_r_14,n1_0_r_14,ACVQN1_0_l_0,);
and I_14(N1_1_l_0,IN_6_1_l_0,n3_1_l_0);
DFFARX1 I_15(N1_1_l_0,blif_clk_net_0_r_14,n1_0_r_14,G199_1_l_0,);
DFFARX1 I_16(IN_3_1_l_0,blif_clk_net_0_r_14,n1_0_r_14,G214_1_l_0,);
nand I_17(n3_1_l_0,IN_1_1_l_0,IN_2_1_l_0);
nor I_18(n_42_5_l_0,IN_1_5_l_0,IN_3_5_l_0);
and I_19(N3_5_l_0,IN_6_5_l_0,n3_5_l_0);
DFFARX1 I_20(N3_5_l_0,blif_clk_net_0_r_14,n1_0_r_14,G199_5_l_0,);
nand I_21(n3_5_l_0,IN_2_5_l_0,IN_3_5_l_0);
not I_22(n12_3_r_0,G199_1_l_0);
or I_23(n_431_3_r_0,n_266_and_0_0_l_0,n14_3_r_0);
nor I_24(n11_3_r_0,G214_1_l_0,n12_3_r_0);
nor I_25(n13_3_r_0,G214_1_l_0,n_42_5_l_0);
and I_26(n14_3_r_0,n_42_5_l_0,n15_3_r_0);
nor I_27(n15_3_r_0,G199_1_l_0,n16_3_r_0);
not I_28(n16_3_r_0,ACVQN2_0_l_0);
nor I_29(n4_4_r_0,ACVQN2_0_l_0,G214_1_l_0);
not I_30(n_87_4_r_0,G199_5_l_0);
and I_31(n7_4_r_0,ACVQN2_0_l_0,n_87_4_r_0);
DFFARX1 I_32(n_266_and_0_0_l_14,blif_clk_net_0_r_14,n1_0_r_14,ACVQN2_0_r_14,);
and I_33(n_266_and_0_0_r_14,G199_5_l_14,ACVQN1_0_r_14);
DFFARX1 I_34(N1_1_r_14,blif_clk_net_0_r_14,n1_0_r_14,G199_1_r_14,);
DFFARX1 I_35(G199_1_l_14,blif_clk_net_0_r_14,n1_0_r_14,G214_1_r_14,);
DFFARX1 I_36(ACVQN2_0_l_14,blif_clk_net_0_r_14,n1_0_r_14,ACVQN1_2_r_14,);
not I_37(P6_2_r_14,P6_internal_2_r_14);
nand I_38(n_429_or_0_3_r_14,G214_1_l_14,n12_3_r_14);
DFFARX1 I_39(n_431_3_r_14,blif_clk_net_0_r_14,n1_0_r_14,G78_3_r_14,);
nand I_40(n_576_3_r_14,ACVQN2_0_l_14,n11_3_r_14);
not I_41(n_102_3_r_14,G199_5_l_14);
nand I_42(n_547_3_r_14,n_266_and_0_0_l_14,n13_3_r_14);
not I_43(n1_0_r_14,blif_reset_net_0_r_14);
DFFARX1 I_44(n_547_3_r_0,blif_clk_net_0_r_14,n1_0_r_14,ACVQN2_0_l_14,);
and I_45(n_266_and_0_0_l_14,ACVQN1_0_l_14,n_569_4_r_0);
DFFARX1 I_46(G78_3_r_0,blif_clk_net_0_r_14,n1_0_r_14,ACVQN1_0_l_14,);
and I_47(N1_1_l_14,n3_1_l_14,G42_4_r_0);
DFFARX1 I_48(N1_1_l_14,blif_clk_net_0_r_14,n1_0_r_14,G199_1_l_14,);
DFFARX1 I_49(n_573_4_r_0,blif_clk_net_0_r_14,n1_0_r_14,G214_1_l_14,);
nand I_50(n3_1_l_14,n_429_or_0_3_r_0,n_576_3_r_0);
nor I_51(n_42_5_l_14,n_102_3_r_0,n_452_4_r_0);
and I_52(N3_5_l_14,n3_5_l_14,n_572_4_r_0);
DFFARX1 I_53(N3_5_l_14,blif_clk_net_0_r_14,n1_0_r_14,G199_5_l_14,);
nand I_54(n3_5_l_14,n_102_3_r_0,n_549_4_r_0);
DFFARX1 I_55(G214_1_l_14,blif_clk_net_0_r_14,n1_0_r_14,ACVQN1_0_r_14,);
and I_56(N1_1_r_14,G214_1_l_14,n3_1_r_14);
nand I_57(n3_1_r_14,ACVQN2_0_l_14,n_42_5_l_14);
DFFARX1 I_58(G199_5_l_14,blif_clk_net_0_r_14,n1_0_r_14,P6_internal_2_r_14,);
not I_59(n12_3_r_14,n_42_5_l_14);
or I_60(n_431_3_r_14,n_266_and_0_0_l_14,n14_3_r_14);
nor I_61(n11_3_r_14,G199_5_l_14,n12_3_r_14);
nor I_62(n13_3_r_14,G199_1_l_14,G199_5_l_14);
and I_63(n14_3_r_14,n_42_5_l_14,n15_3_r_14);
nor I_64(n15_3_r_14,G199_1_l_14,n16_3_r_14);
not I_65(n16_3_r_14,G214_1_l_14);
endmodule


