module test_I5713(I2167,I2173,I1477,I1470,I5713);
input I2167,I2173,I1477,I1470;
output I5713;
wire I4629,I2143,I5751,I6110,I4544,I6127,I4533,I5013,I4807,I4824,I4509;
nor I_0(I4629,I2167,I2173);
DFFARX1 I_1(I1470,,,I2143,);
not I_2(I5751,I1477);
DFFARX1 I_3(I6127,I1470,I5751,,,I5713,);
DFFARX1 I_4(I4509,I1470,I5751,,,I6110,);
not I_5(I4544,I1477);
and I_6(I6127,I6110,I4533);
or I_7(I4533,I4824,I4629);
or I_8(I5013,I4824);
DFFARX1 I_9(I1470,I4544,,,I4807,);
and I_10(I4824,I4807,I2143);
DFFARX1 I_11(I5013,I1470,I4544,,,I4509,);
endmodule


