module test_final(IN_1_4_l,IN_2_4_l,IN_3_4_l,IN_4_4_l,IN_5_4_l,IN_1_6_l,IN_2_6_l,IN_3_6_l,IN_4_6_l,IN_5_6_l,IN_1_9_l,IN_2_9_l,IN_3_9_l,IN_4_9_l,IN_5_9_l,blif_clk_net_8_r,blif_reset_net_8_r,N1371_0_r,N1508_0_r,N1372_1_r,N1508_1_r,N1507_6_r,N1508_6_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r,N1372_10_r,N1508_10_r);
input IN_1_4_l,IN_2_4_l,IN_3_4_l,IN_4_4_l,IN_5_4_l,IN_1_6_l,IN_2_6_l,IN_3_6_l,IN_4_6_l,IN_5_6_l,IN_1_9_l,IN_2_9_l,IN_3_9_l,IN_4_9_l,IN_5_9_l,blif_clk_net_8_r,blif_reset_net_8_r;
output N1371_0_r,N1508_0_r,N1372_1_r,N1508_1_r,N1507_6_r,N1508_6_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r,N1372_10_r,N1508_10_r;
wire N1372_4_l,N1508_4_l,n6_4_l,n7_4_l,n8_4_l,N1507_6_l,N1508_6_l,n6_6_l,n7_6_l,n8_6_l,n9_6_l,N6150_9_l,N6147_9_l,N6134_9_l,n3_9_l,I_BUFF_1_9_l,n3_0_r,n4_0_r,n4_1_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,N3_8_r,n1_8_r,n3_8_r,N6150_9_r,n3_9_r,n5_10_r,n6_10_r;
not I_0(N1372_4_l,n7_4_l);
nor I_1(N1508_4_l,n6_4_l,n7_4_l);
nor I_2(n6_4_l,IN_5_4_l,n8_4_l);
nand I_3(n7_4_l,IN_1_4_l,IN_2_4_l);
and I_4(n8_4_l,IN_3_4_l,IN_4_4_l);
nor I_5(N1507_6_l,n8_6_l,n9_6_l);
and I_6(N1508_6_l,IN_2_6_l,n6_6_l);
nor I_7(n6_6_l,n7_6_l,n8_6_l);
not I_8(n7_6_l,IN_1_6_l);
nor I_9(n8_6_l,IN_5_6_l,n9_6_l);
and I_10(n9_6_l,IN_3_6_l,IN_4_6_l);
not I_11(N6150_9_l,IN_2_9_l);
nor I_12(N6147_9_l,N6150_9_l,n3_9_l);
nor I_13(N6134_9_l,IN_5_9_l,n3_9_l);
nor I_14(n3_9_l,IN_3_9_l,IN_4_9_l);
buf I_15(I_BUFF_1_9_l,IN_1_9_l);
nor I_16(N1371_0_r,n4_0_r,I_BUFF_1_9_l);
nor I_17(N1508_0_r,n3_0_r,n4_0_r);
nor I_18(n3_0_r,N1372_4_l,N1507_6_l);
not I_19(n4_0_r,N1508_6_l);
not I_20(N1372_1_r,n4_1_r);
nor I_21(N1508_1_r,n4_1_r,I_BUFF_1_9_l);
nand I_22(n4_1_r,N1507_6_l,I_BUFF_1_9_l);
nor I_23(N1507_6_r,n8_6_r,n9_6_r);
and I_24(N1508_6_r,n6_6_r,N1508_6_l);
nor I_25(n6_6_r,n7_6_r,n8_6_r);
not I_26(n7_6_r,N1507_6_l);
nor I_27(n8_6_r,n9_6_r,N6147_9_l);
and I_28(n9_6_r,N1508_4_l,N1508_6_l);
nor I_29(n_42_8_r,N6147_9_l,N6134_9_l);
DFFARX1 I_30(N3_8_r,blif_clk_net_8_r,n1_8_r,G199_8_r,);
and I_31(N3_8_r,n3_8_r,N6134_9_l);
not I_32(n1_8_r,blif_reset_net_8_r);
nand I_33(n3_8_r,N6147_9_l,N1508_6_l);
not I_34(N6150_9_r,N6134_9_l);
nor I_35(N6147_9_r,N6150_9_r,n3_9_r);
nor I_36(N6134_9_r,n3_9_r,N6147_9_l);
nor I_37(n3_9_r,N1372_4_l,N1508_4_l);
buf I_38(I_BUFF_1_9_r,N6147_9_l);
not I_39(N1372_10_r,n6_10_r);
nor I_40(N1508_10_r,n5_10_r,n6_10_r);
nor I_41(n5_10_r,N1508_4_l,N1507_6_l);
nand I_42(n6_10_r,N1372_4_l,N1508_4_l);
endmodule


