module test_I14421(I1477,I11299,I1470,I13508,I14421);
input I1477,I11299,I1470,I13508;
output I14421;
wire I13460,I13601,I13183,I13197,I13248,I13426,I14404,I13186,I13525,I13171,I14387,I14370;
not I_0(I13460,I13426);
DFFARX1 I_1(I11299,I1470,I13197,,,I13601,);
nand I_2(I13183,I13601,I13525);
not I_3(I13197,I1477);
DFFARX1 I_4(I1470,I13197,,,I13248,);
DFFARX1 I_5(I1470,I13197,,,I13426,);
and I_6(I14404,I14387,I13183);
nor I_7(I13186,I13601,I13508);
DFFARX1 I_8(I14404,I1470,I14370,,,I14421,);
nor I_9(I13525,I13508,I13426);
nand I_10(I13171,I13248,I13460);
nand I_11(I14387,I13171,I13186);
not I_12(I14370,I1477);
endmodule


