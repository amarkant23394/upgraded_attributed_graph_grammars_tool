module test_I7444(I1477,I5249,I5204,I1470,I7444);
input I1477,I5249,I5204,I1470;
output I7444;
wire I5368,I6907,I5097,I5481,I6975,I7410,I5073,I6992,I5594,I5625,I5070,I5642,I6924,I5351,I7427,I5082;
nor I_0(I5368,I5351,I5204);
not I_1(I6907,I1477);
nand I_2(I5097,I5642,I5368);
DFFARX1 I_3(I1470,,,I5481,);
nand I_4(I7444,I7427,I6992);
nor I_5(I6975,I6924,I5070);
DFFARX1 I_6(I5082,I1470,I6907,,,I7410,);
DFFARX1 I_7(I1470,,,I5073,);
nand I_8(I6992,I6975,I5097);
DFFARX1 I_9(I1470,,,I5594,);
DFFARX1 I_10(I1470,,,I5625,);
and I_11(I5070,I5249,I5481);
not I_12(I5642,I5625);
not I_13(I6924,I5073);
DFFARX1 I_14(I1470,,,I5351,);
not I_15(I7427,I7410);
not I_16(I5082,I5594);
endmodule


