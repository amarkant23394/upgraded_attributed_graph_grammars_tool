module test_final(IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_7_r_4,blif_reset_net_7_r_4,N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4);
input IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_7_r_4,blif_reset_net_7_r_4;
output N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4;
wire N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_102_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15,n_431_5_r_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15,N1508_0_r_4,n_573_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n6_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4;
and I_0(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_1(N1508_0_r_15,IN_2_0_l_15,n55_15);
nor I_2(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_3(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_4(N1372_4_r_15,n39_15);
nor I_5(N1508_4_r_15,n39_15,n43_15);
nand I_6(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_7(n_431_5_r_15,blif_clk_net_7_r_4,n6_4,G78_5_r_15,);
nand I_8(n_576_5_r_15,n31_15,n32_15);
not I_9(n_102_5_r_15,n33_15);
nand I_10(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_11(N1507_6_r_15,n42_15,n46_15);
nand I_12(N1508_6_r_15,n39_15,n40_15);
nand I_13(n_431_5_r_15,n36_15,n37_15);
nor I_14(n31_15,n33_15,n34_15);
nor I_15(n32_15,IN_1_3_l_15,n44_15);
nor I_16(n33_15,n54_15,n55_15);
nand I_17(n34_15,IN_2_6_l_15,n49_15);
nand I_18(n35_15,IN_1_1_l_15,IN_2_1_l_15);
not I_19(n36_15,n32_15);
nand I_20(n37_15,n34_15,n38_15);
not I_21(n38_15,n46_15);
nand I_22(n39_15,n38_15,n41_15);
nand I_23(n40_15,n41_15,n42_15);
and I_24(n41_15,IN_5_6_l_15,n51_15);
and I_25(n42_15,IN_2_1_l_15,n47_15);
and I_26(n43_15,n34_15,n36_15);
or I_27(n44_15,IN_2_3_l_15,IN_3_3_l_15);
not I_28(n45_15,N1372_1_r_15);
nand I_29(n46_15,IN_2_1_l_15,n53_15);
nor I_30(n47_15,n34_15,n48_15);
not I_31(n48_15,IN_1_1_l_15);
and I_32(n49_15,IN_1_6_l_15,n50_15);
nand I_33(n50_15,n51_15,n52_15);
nand I_34(n51_15,IN_3_6_l_15,IN_4_6_l_15);
not I_35(n52_15,IN_5_6_l_15);
nor I_36(n53_15,IN_3_1_l_15,n48_15);
nor I_37(n54_15,IN_3_0_l_15,IN_4_0_l_15);
not I_38(n55_15,IN_1_0_l_15);
nor I_39(N1371_0_r_4,n25_4,n_576_5_r_15);
not I_40(N1508_0_r_4,n25_4);
nor I_41(N1507_6_r_4,n32_4,n33_4);
nor I_42(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_43(n4_7_r_4,blif_clk_net_7_r_4,n6_4,G42_7_r_4,);
not I_44(n_572_7_r_4,n_573_7_r_4);
nand I_45(n_573_7_r_4,n21_4,n22_4);
nor I_46(n_549_7_r_4,n24_4,n_576_5_r_15);
nand I_47(n_569_7_r_4,n22_4,n23_4);
nor I_48(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_49(N6147_9_r_4,n28_4);
nor I_50(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_51(I_BUFF_1_9_r_4,n21_4);
nor I_52(n4_7_r_4,N6147_9_r_4,n_576_5_r_15);
not I_53(n6_4,blif_reset_net_7_r_4);
nand I_54(n21_4,n39_4,n40_4);
or I_55(n22_4,n31_4,G78_5_r_15);
not I_56(n23_4,n_576_5_r_15);
nor I_57(n24_4,n25_4,n26_4);
nand I_58(n25_4,N1508_6_r_15,G78_5_r_15);
nand I_59(n26_4,n21_4,n27_4);
nand I_60(n27_4,n36_4,n37_4);
nand I_61(n28_4,n38_4,N1508_1_r_15);
nand I_62(n29_4,N1508_0_r_4,n30_4);
nand I_63(n30_4,n34_4,n35_4);
nor I_64(n31_4,n_547_5_r_15,n_429_or_0_5_r_15);
not I_65(n32_4,n30_4);
nor I_66(n33_4,n21_4,n28_4);
nand I_67(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_68(n35_4,N1508_0_r_4,n27_4);
not I_69(n36_4,N1508_1_r_15);
nand I_70(n37_4,N1372_4_r_15,N1508_4_r_15);
or I_71(n38_4,n_547_5_r_15,n_429_or_0_5_r_15);
nor I_72(n39_4,N1508_4_r_15,n_547_5_r_15);
or I_73(n40_4,n41_4,N1507_6_r_15);
nor I_74(n41_4,n_429_or_0_5_r_15,n_576_5_r_15);
endmodule


