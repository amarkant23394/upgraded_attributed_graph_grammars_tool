module Benchmark_testing1000(I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1470,I1477,I5127,I5142,I5139,I5124,I5121,I5148,I5136,I5130,I5145,I5133,I5118,I12080,I12077,I12071,I12101,I12074,I12098,I12095,I12092,I12086,I12089,I12083,I14625,I14628,I14610,I14631,I14622,I14613,I14604,I14634,I14619,I14616,I14607);
input I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1470,I1477;
output I5127,I5142,I5139,I5124,I5121,I5148,I5136,I5130,I5145,I5133,I5118,I12080,I12077,I12071,I12101,I12074,I12098,I12095,I12092,I12086,I12089,I12083,I14625,I14628,I14610,I14631,I14622,I14613,I14604,I14634,I14619,I14616,I14607;
wire I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1470,I1477,I1518,I1535,I15202,I15205,I1552,I15217,I1569,I1586,I1603,I15211,I1501,I1489,I1648,I15214,I1665,I1682,I15208,I15226,I1699,I15229,I1716,I1498,I1747,I1764,I1781,I15199,I1798,I15220,I1507,I1486,I1843,I15223,I1860,I1504,I1891,I1495,I1510,I1936,I1953,I1970,I1987,I1483,I1492,I1480,I2079,I2096,I12747,I12738,I2113,I12741,I2130,I2147,I2164,I12717,I2062,I2050,I2209,I12732,I2226,I2243,I12720,I12735,I2260,I12729,I2277,I2059,I2308,I2325,I2342,I12744,I2359,I12723,I2068,I2047,I2404,I12726,I2421,I2065,I2452,I2056,I2071,I2497,I2514,I2531,I2548,I2044,I2053,I2041,I2640,I2657,I8253,I8256,I2674,I8250,I2691,I2708,I2725,I8241,I2623,I2611,I2770,I8229,I2787,I2804,I8238,I8232,I2821,I8244,I2838,I2620,I2869,I2886,I2903,I8259,I2920,I8247,I2629,I2608,I2965,I8235,I2982,I2626,I3013,I2617,I2632,I3058,I3075,I3092,I3109,I2605,I2614,I2602,I3201,I3218,I4473,I3235,I4461,I4467,I3252,I4476,I3175,I3283,I3300,I4464,I3190,I3172,I3345,I3362,I3379,I4485,I3396,I4458,I3413,I4479,I3430,I4470,I3447,I3464,I3481,I3187,I3512,I3529,I3546,I3169,I3577,I3166,I3608,I4455,I3625,I3642,I3659,I3181,I3690,I3178,I3721,I4482,I3738,I3755,I3184,I3193,I3163,I3847,I3864,I16404,I3881,I16389,I16416,I3898,I16392,I3821,I3929,I3946,I16407,I3836,I3818,I3991,I4008,I4025,I16419,I4042,I16401,I4059,I16410,I4076,I16395,I4093,I4110,I4127,I3833,I4158,I4175,I4192,I3815,I4223,I3812,I4254,I16398,I4271,I4288,I4305,I3827,I4336,I3824,I4367,I16413,I4384,I4401,I3830,I3839,I3809,I4493,I4510,I4527,I4544,I4575,I4592,I4609,I4626,I4643,I4660,I4677,I4694,I4711,I4728,I4773,I4804,I4835,I4852,I4869,I4886,I4903,I4920,I4951,I4996,I5013,I5044,I5061,I5078,I5156,I5173,I16996,I5190,I17002,I17014,I5207,I17005,I5238,I5255,I16984,I5272,I5289,I5306,I16999,I5323,I16987,I5340,I17008,I5357,I16990,I5374,I5391,I5436,I5467,I5498,I5515,I5532,I5549,I17011,I5566,I5583,I5614,I5659,I16993,I5676,I5707,I5724,I5741,I5819,I5836,I5853,I5870,I5790,I5901,I5918,I5935,I5952,I5969,I5986,I6003,I6020,I6037,I6054,I5805,I5802,I6099,I5787,I6130,I5784,I6161,I6178,I6195,I6212,I6229,I6246,I5811,I6277,I5799,I5793,I6322,I6339,I5808,I6370,I6387,I6404,I5796,I5781,I6482,I6499,I11408,I11423,I6516,I11411,I6456,I6547,I11414,I11429,I6564,I6581,I6598,I11417,I6615,I6632,I11420,I11438,I6649,I6666,I6683,I6450,I6714,I6731,I6447,I6762,I11435,I6779,I11426,I6796,I6459,I6444,I6841,I11432,I6858,I6875,I6892,I6909,I6465,I6940,I6474,I6971,I6468,I6471,I6462,I6453,I7077,I7094,I10745,I10760,I7111,I10748,I7051,I7142,I10751,I10766,I7159,I7176,I7193,I10754,I7210,I7227,I10757,I10775,I7244,I7261,I7278,I7045,I7309,I7326,I7042,I7357,I10772,I7374,I10763,I7391,I7054,I7039,I7436,I10769,I7453,I7470,I7487,I7504,I7060,I7535,I7069,I7566,I7063,I7066,I7057,I7048,I7672,I7689,I7706,I7646,I7737,I7754,I7771,I7788,I7805,I7822,I7839,I7856,I7873,I7640,I7904,I7921,I7637,I7952,I7969,I7986,I7649,I7634,I8031,I8048,I8065,I8082,I8099,I7655,I8130,I7664,I8161,I7658,I7661,I7652,I7643,I8267,I8284,I8301,I8332,I8349,I8366,I8383,I8400,I8417,I8434,I8451,I8468,I8499,I8516,I8547,I8564,I8581,I8626,I8643,I8660,I8677,I8694,I8725,I8756,I8862,I8879,I8896,I8836,I8927,I8944,I8961,I8978,I8995,I9012,I9029,I9046,I9063,I8830,I9094,I9111,I8827,I9142,I9159,I9176,I8839,I8824,I9221,I9238,I9255,I9272,I9289,I8845,I9320,I8854,I9351,I8848,I8851,I8842,I8833,I9457,I9474,I9491,I9508,I9525,I9542,I9559,I9576,I9446,I9607,I9431,I9638,I9655,I9672,I9689,I9706,I9723,I9740,I9428,I9771,I9788,I9425,I9819,I9836,I9443,I9867,I9440,I9898,I9915,I9419,I9422,I9960,I9977,I9994,I10011,I9449,I10042,I9434,I9437,I10120,I10137,I10154,I10171,I10188,I10205,I10222,I10239,I10109,I10270,I10094,I10301,I10318,I10335,I10352,I10369,I10386,I10403,I10091,I10434,I10451,I10088,I10482,I10499,I10106,I10530,I10103,I10561,I10578,I10082,I10085,I10623,I10640,I10657,I10674,I10112,I10705,I10097,I10100,I10783,I10800,I13375,I10817,I13372,I13390,I10834,I13393,I10851,I10868,I13378,I10885,I10902,I10933,I10964,I13387,I10981,I13369,I10998,I13363,I11015,I13381,I11032,I11049,I11066,I11097,I11114,I11145,I13366,I11162,I11193,I11224,I11241,I11286,I13384,I11303,I11320,I11337,I11368,I11446,I11463,I11480,I11497,I11514,I11531,I11548,I11565,I11596,I11627,I11644,I11661,I11678,I11695,I11712,I11729,I11760,I11777,I11808,I11825,I11856,I11887,I11904,I11949,I11966,I11983,I12000,I12031,I12109,I12126,I12143,I12160,I12177,I12194,I12211,I12242,I12259,I12276,I12293,I12310,I12327,I12344,I12375,I12406,I12423,I12440,I12485,I12516,I12561,I12578,I12595,I12612,I12629,I12660,I12677,I12755,I12772,I12789,I12806,I12823,I12840,I12857,I12888,I12905,I12922,I12939,I12956,I12973,I12990,I13021,I13052,I13069,I13086,I13131,I13162,I13207,I13224,I13241,I13258,I13275,I13306,I13323,I13401,I13418,I14018,I13435,I14030,I14024,I13452,I14009,I13469,I13486,I14036,I13503,I13534,I13551,I13568,I14033,I13585,I14015,I13602,I14012,I13619,I14039,I13636,I13667,I13698,I13715,I13732,I13777,I14027,I13808,I13853,I14021,I13870,I13887,I13904,I13921,I13952,I13969,I14047,I14064,I17625,I17631,I14081,I17622,I14098,I14115,I17634,I14132,I14163,I17613,I14180,I14197,I14242,I17637,I17619,I14259,I17628,I14276,I14321,I17643,I14338,I17616,I14355,I14386,I14403,I14434,I17640,I14451,I14468,I14499,I14516,I14533,I14550,I14642,I14659,I14676,I14693,I14710,I14727,I14758,I14775,I14792,I14837,I14854,I14871,I14916,I14933,I14950,I14981,I14998,I15029,I15046,I15063,I15094,I15111,I15128,I15145,I15237,I15254,I15271,I15288,I15305,I15322,I15353,I15370,I15387,I15432,I15449,I15466,I15511,I15528,I15545,I15576,I15593,I15624,I15641,I15658,I15689,I15706,I15723,I15740,I15832,I15849,I15866,I15883,I15900,I15917,I15815,I15948,I15965,I15982,I15818,I15800,I16027,I16044,I16061,I15821,I15812,I16106,I16123,I16140,I15803,I16171,I16188,I15794,I16219,I16236,I16253,I15824,I16284,I16301,I16318,I16335,I15809,I15806,I15797,I16427,I16444,I16461,I16478,I16495,I16512,I16529,I16560,I16577,I16594,I16611,I16628,I16645,I16662,I16707,I16724,I16741,I16772,I16789,I16834,I16865,I16882,I16913,I16958,I17022,I17039,I17056,I17073,I17090,I17107,I17124,I17141,I17158,I17175,I17192,I17209,I17226,I17243,I17274,I17291,I17308,I17339,I17370,I17387,I17418,I17463,I17480,I17497,I17556,I17573,I17651,I17668,I17685,I17702,I17733,I17764,I17781,I17798,I17815,I17832,I17863,I17894,I17911,I17928,I17945,I17962,I17979,I18010,I18027,I18044,I18103,I18148,I18165;
not I_0 (I1518,I1477);
nand I_1 (I1535,I15202,I15205);
and I_2 (I1552,I1535,I15217);
DFFARX1 I_3  ( .D(I1552), .CLK(I1470), .RSTB(I1518), .Q(I1569) );
not I_4 (I1586,I1569);
nor I_5 (I1603,I15211,I15205);
or I_6 (I1501,I1603,I1569);
not I_7 (I1489,I1603);
DFFARX1 I_8  ( .D(I15214), .CLK(I1470), .RSTB(I1518), .Q(I1648) );
nor I_9 (I1665,I1648,I1603);
nand I_10 (I1682,I15208,I15226);
and I_11 (I1699,I1682,I15229);
DFFARX1 I_12  ( .D(I1699), .CLK(I1470), .RSTB(I1518), .Q(I1716) );
nor I_13 (I1498,I1716,I1569);
not I_14 (I1747,I1716);
nor I_15 (I1764,I1648,I1747);
DFFARX1 I_16  ( .D(I15199), .CLK(I1470), .RSTB(I1518), .Q(I1781) );
and I_17 (I1798,I1781,I15220);
or I_18 (I1507,I1798,I1603);
nand I_19 (I1486,I1798,I1764);
DFFARX1 I_20  ( .D(I15223), .CLK(I1470), .RSTB(I1518), .Q(I1843) );
and I_21 (I1860,I1843,I1586);
nor I_22 (I1504,I1798,I1860);
nor I_23 (I1891,I1843,I1648);
DFFARX1 I_24  ( .D(I1891), .CLK(I1470), .RSTB(I1518), .Q(I1495) );
nor I_25 (I1510,I1843,I1569);
not I_26 (I1936,I1843);
nor I_27 (I1953,I1716,I1936);
and I_28 (I1970,I1603,I1953);
or I_29 (I1987,I1798,I1970);
DFFARX1 I_30  ( .D(I1987), .CLK(I1470), .RSTB(I1518), .Q(I1483) );
nand I_31 (I1492,I1843,I1665);
nand I_32 (I1480,I1843,I1747);
not I_33 (I2079,I1477);
nand I_34 (I2096,I12747,I12738);
and I_35 (I2113,I2096,I12741);
DFFARX1 I_36  ( .D(I2113), .CLK(I1470), .RSTB(I2079), .Q(I2130) );
not I_37 (I2147,I2130);
nor I_38 (I2164,I12717,I12738);
or I_39 (I2062,I2164,I2130);
not I_40 (I2050,I2164);
DFFARX1 I_41  ( .D(I12732), .CLK(I1470), .RSTB(I2079), .Q(I2209) );
nor I_42 (I2226,I2209,I2164);
nand I_43 (I2243,I12720,I12735);
and I_44 (I2260,I2243,I12729);
DFFARX1 I_45  ( .D(I2260), .CLK(I1470), .RSTB(I2079), .Q(I2277) );
nor I_46 (I2059,I2277,I2130);
not I_47 (I2308,I2277);
nor I_48 (I2325,I2209,I2308);
DFFARX1 I_49  ( .D(I12744), .CLK(I1470), .RSTB(I2079), .Q(I2342) );
and I_50 (I2359,I2342,I12723);
or I_51 (I2068,I2359,I2164);
nand I_52 (I2047,I2359,I2325);
DFFARX1 I_53  ( .D(I12726), .CLK(I1470), .RSTB(I2079), .Q(I2404) );
and I_54 (I2421,I2404,I2147);
nor I_55 (I2065,I2359,I2421);
nor I_56 (I2452,I2404,I2209);
DFFARX1 I_57  ( .D(I2452), .CLK(I1470), .RSTB(I2079), .Q(I2056) );
nor I_58 (I2071,I2404,I2130);
not I_59 (I2497,I2404);
nor I_60 (I2514,I2277,I2497);
and I_61 (I2531,I2164,I2514);
or I_62 (I2548,I2359,I2531);
DFFARX1 I_63  ( .D(I2548), .CLK(I1470), .RSTB(I2079), .Q(I2044) );
nand I_64 (I2053,I2404,I2226);
nand I_65 (I2041,I2404,I2308);
not I_66 (I2640,I1477);
nand I_67 (I2657,I8253,I8256);
and I_68 (I2674,I2657,I8250);
DFFARX1 I_69  ( .D(I2674), .CLK(I1470), .RSTB(I2640), .Q(I2691) );
not I_70 (I2708,I2691);
nor I_71 (I2725,I8241,I8256);
or I_72 (I2623,I2725,I2691);
not I_73 (I2611,I2725);
DFFARX1 I_74  ( .D(I8229), .CLK(I1470), .RSTB(I2640), .Q(I2770) );
nor I_75 (I2787,I2770,I2725);
nand I_76 (I2804,I8238,I8232);
and I_77 (I2821,I2804,I8244);
DFFARX1 I_78  ( .D(I2821), .CLK(I1470), .RSTB(I2640), .Q(I2838) );
nor I_79 (I2620,I2838,I2691);
not I_80 (I2869,I2838);
nor I_81 (I2886,I2770,I2869);
DFFARX1 I_82  ( .D(I8259), .CLK(I1470), .RSTB(I2640), .Q(I2903) );
and I_83 (I2920,I2903,I8247);
or I_84 (I2629,I2920,I2725);
nand I_85 (I2608,I2920,I2886);
DFFARX1 I_86  ( .D(I8235), .CLK(I1470), .RSTB(I2640), .Q(I2965) );
and I_87 (I2982,I2965,I2708);
nor I_88 (I2626,I2920,I2982);
nor I_89 (I3013,I2965,I2770);
DFFARX1 I_90  ( .D(I3013), .CLK(I1470), .RSTB(I2640), .Q(I2617) );
nor I_91 (I2632,I2965,I2691);
not I_92 (I3058,I2965);
nor I_93 (I3075,I2838,I3058);
and I_94 (I3092,I2725,I3075);
or I_95 (I3109,I2920,I3092);
DFFARX1 I_96  ( .D(I3109), .CLK(I1470), .RSTB(I2640), .Q(I2605) );
nand I_97 (I2614,I2965,I2787);
nand I_98 (I2602,I2965,I2869);
not I_99 (I3201,I1477);
not I_100 (I3218,I4473);
nor I_101 (I3235,I4461,I4467);
nand I_102 (I3252,I3235,I4476);
DFFARX1 I_103  ( .D(I3252), .CLK(I1470), .RSTB(I3201), .Q(I3175) );
nor I_104 (I3283,I3218,I4461);
nand I_105 (I3300,I3283,I4464);
not I_106 (I3190,I3300);
DFFARX1 I_107  ( .D(I3300), .CLK(I1470), .RSTB(I3201), .Q(I3172) );
not I_108 (I3345,I4461);
not I_109 (I3362,I3345);
not I_110 (I3379,I4485);
nor I_111 (I3396,I3379,I4458);
and I_112 (I3413,I3396,I4479);
or I_113 (I3430,I3413,I4470);
DFFARX1 I_114  ( .D(I3430), .CLK(I1470), .RSTB(I3201), .Q(I3447) );
nor I_115 (I3464,I3447,I3300);
nor I_116 (I3481,I3447,I3362);
nand I_117 (I3187,I3252,I3481);
nand I_118 (I3512,I3218,I4485);
nand I_119 (I3529,I3512,I3447);
and I_120 (I3546,I3512,I3529);
DFFARX1 I_121  ( .D(I3546), .CLK(I1470), .RSTB(I3201), .Q(I3169) );
DFFARX1 I_122  ( .D(I3512), .CLK(I1470), .RSTB(I3201), .Q(I3577) );
and I_123 (I3166,I3345,I3577);
DFFARX1 I_124  ( .D(I4455), .CLK(I1470), .RSTB(I3201), .Q(I3608) );
not I_125 (I3625,I3608);
nor I_126 (I3642,I3300,I3625);
and I_127 (I3659,I3608,I3642);
nand I_128 (I3181,I3608,I3362);
DFFARX1 I_129  ( .D(I3608), .CLK(I1470), .RSTB(I3201), .Q(I3690) );
not I_130 (I3178,I3690);
DFFARX1 I_131  ( .D(I4482), .CLK(I1470), .RSTB(I3201), .Q(I3721) );
not I_132 (I3738,I3721);
or I_133 (I3755,I3738,I3659);
DFFARX1 I_134  ( .D(I3755), .CLK(I1470), .RSTB(I3201), .Q(I3184) );
nand I_135 (I3193,I3738,I3464);
DFFARX1 I_136  ( .D(I3738), .CLK(I1470), .RSTB(I3201), .Q(I3163) );
not I_137 (I3847,I1477);
not I_138 (I3864,I16404);
nor I_139 (I3881,I16389,I16416);
nand I_140 (I3898,I3881,I16392);
DFFARX1 I_141  ( .D(I3898), .CLK(I1470), .RSTB(I3847), .Q(I3821) );
nor I_142 (I3929,I3864,I16389);
nand I_143 (I3946,I3929,I16407);
not I_144 (I3836,I3946);
DFFARX1 I_145  ( .D(I3946), .CLK(I1470), .RSTB(I3847), .Q(I3818) );
not I_146 (I3991,I16389);
not I_147 (I4008,I3991);
not I_148 (I4025,I16419);
nor I_149 (I4042,I4025,I16401);
and I_150 (I4059,I4042,I16410);
or I_151 (I4076,I4059,I16395);
DFFARX1 I_152  ( .D(I4076), .CLK(I1470), .RSTB(I3847), .Q(I4093) );
nor I_153 (I4110,I4093,I3946);
nor I_154 (I4127,I4093,I4008);
nand I_155 (I3833,I3898,I4127);
nand I_156 (I4158,I3864,I16419);
nand I_157 (I4175,I4158,I4093);
and I_158 (I4192,I4158,I4175);
DFFARX1 I_159  ( .D(I4192), .CLK(I1470), .RSTB(I3847), .Q(I3815) );
DFFARX1 I_160  ( .D(I4158), .CLK(I1470), .RSTB(I3847), .Q(I4223) );
and I_161 (I3812,I3991,I4223);
DFFARX1 I_162  ( .D(I16398), .CLK(I1470), .RSTB(I3847), .Q(I4254) );
not I_163 (I4271,I4254);
nor I_164 (I4288,I3946,I4271);
and I_165 (I4305,I4254,I4288);
nand I_166 (I3827,I4254,I4008);
DFFARX1 I_167  ( .D(I4254), .CLK(I1470), .RSTB(I3847), .Q(I4336) );
not I_168 (I3824,I4336);
DFFARX1 I_169  ( .D(I16413), .CLK(I1470), .RSTB(I3847), .Q(I4367) );
not I_170 (I4384,I4367);
or I_171 (I4401,I4384,I4305);
DFFARX1 I_172  ( .D(I4401), .CLK(I1470), .RSTB(I3847), .Q(I3830) );
nand I_173 (I3839,I4384,I4110);
DFFARX1 I_174  ( .D(I4384), .CLK(I1470), .RSTB(I3847), .Q(I3809) );
not I_175 (I4493,I1477);
not I_176 (I4510,I1207);
nor I_177 (I4527,I1239,I1407);
nand I_178 (I4544,I4527,I1343);
DFFARX1 I_179  ( .D(I4544), .CLK(I1470), .RSTB(I4493), .Q(I4464) );
nor I_180 (I4575,I4510,I1239);
nand I_181 (I4592,I4575,I1327);
nand I_182 (I4609,I4592,I4544);
not I_183 (I4626,I1239);
not I_184 (I4643,I1455);
nor I_185 (I4660,I4643,I1215);
and I_186 (I4677,I4660,I1287);
or I_187 (I4694,I4677,I1447);
DFFARX1 I_188  ( .D(I4694), .CLK(I1470), .RSTB(I4493), .Q(I4711) );
nor I_189 (I4728,I4711,I4592);
nand I_190 (I4479,I4626,I4728);
not I_191 (I4476,I4711);
and I_192 (I4773,I4711,I4609);
DFFARX1 I_193  ( .D(I4773), .CLK(I1470), .RSTB(I4493), .Q(I4461) );
DFFARX1 I_194  ( .D(I4711), .CLK(I1470), .RSTB(I4493), .Q(I4804) );
and I_195 (I4458,I4626,I4804);
nand I_196 (I4835,I4510,I1455);
not I_197 (I4852,I4835);
nor I_198 (I4869,I4711,I4852);
DFFARX1 I_199  ( .D(I1399), .CLK(I1470), .RSTB(I4493), .Q(I4886) );
nand I_200 (I4903,I4886,I4835);
and I_201 (I4920,I4626,I4903);
DFFARX1 I_202  ( .D(I4920), .CLK(I1470), .RSTB(I4493), .Q(I4485) );
not I_203 (I4951,I4886);
nand I_204 (I4473,I4886,I4869);
nand I_205 (I4467,I4886,I4852);
DFFARX1 I_206  ( .D(I1303), .CLK(I1470), .RSTB(I4493), .Q(I4996) );
not I_207 (I5013,I4996);
nor I_208 (I4482,I4886,I5013);
nor I_209 (I5044,I5013,I4951);
and I_210 (I5061,I4592,I5044);
or I_211 (I5078,I4835,I5061);
DFFARX1 I_212  ( .D(I5078), .CLK(I1470), .RSTB(I4493), .Q(I4470) );
DFFARX1 I_213  ( .D(I5013), .CLK(I1470), .RSTB(I4493), .Q(I4455) );
not I_214 (I5156,I1477);
not I_215 (I5173,I16996);
nor I_216 (I5190,I17002,I17014);
nand I_217 (I5207,I5190,I17005);
DFFARX1 I_218  ( .D(I5207), .CLK(I1470), .RSTB(I5156), .Q(I5127) );
nor I_219 (I5238,I5173,I17002);
nand I_220 (I5255,I5238,I16984);
nand I_221 (I5272,I5255,I5207);
not I_222 (I5289,I17002);
not I_223 (I5306,I16999);
nor I_224 (I5323,I5306,I16987);
and I_225 (I5340,I5323,I17008);
or I_226 (I5357,I5340,I16990);
DFFARX1 I_227  ( .D(I5357), .CLK(I1470), .RSTB(I5156), .Q(I5374) );
nor I_228 (I5391,I5374,I5255);
nand I_229 (I5142,I5289,I5391);
not I_230 (I5139,I5374);
and I_231 (I5436,I5374,I5272);
DFFARX1 I_232  ( .D(I5436), .CLK(I1470), .RSTB(I5156), .Q(I5124) );
DFFARX1 I_233  ( .D(I5374), .CLK(I1470), .RSTB(I5156), .Q(I5467) );
and I_234 (I5121,I5289,I5467);
nand I_235 (I5498,I5173,I16999);
not I_236 (I5515,I5498);
nor I_237 (I5532,I5374,I5515);
DFFARX1 I_238  ( .D(I17011), .CLK(I1470), .RSTB(I5156), .Q(I5549) );
nand I_239 (I5566,I5549,I5498);
and I_240 (I5583,I5289,I5566);
DFFARX1 I_241  ( .D(I5583), .CLK(I1470), .RSTB(I5156), .Q(I5148) );
not I_242 (I5614,I5549);
nand I_243 (I5136,I5549,I5532);
nand I_244 (I5130,I5549,I5515);
DFFARX1 I_245  ( .D(I16993), .CLK(I1470), .RSTB(I5156), .Q(I5659) );
not I_246 (I5676,I5659);
nor I_247 (I5145,I5549,I5676);
nor I_248 (I5707,I5676,I5614);
and I_249 (I5724,I5255,I5707);
or I_250 (I5741,I5498,I5724);
DFFARX1 I_251  ( .D(I5741), .CLK(I1470), .RSTB(I5156), .Q(I5133) );
DFFARX1 I_252  ( .D(I5676), .CLK(I1470), .RSTB(I5156), .Q(I5118) );
not I_253 (I5819,I1477);
not I_254 (I5836,I1383);
nor I_255 (I5853,I1431,I1359);
nand I_256 (I5870,I5853,I1423);
DFFARX1 I_257  ( .D(I5870), .CLK(I1470), .RSTB(I5819), .Q(I5790) );
nor I_258 (I5901,I5836,I1431);
nand I_259 (I5918,I5901,I1415);
nand I_260 (I5935,I5918,I5870);
not I_261 (I5952,I1431);
not I_262 (I5969,I1231);
nor I_263 (I5986,I5969,I1271);
and I_264 (I6003,I5986,I1263);
or I_265 (I6020,I6003,I1367);
DFFARX1 I_266  ( .D(I6020), .CLK(I1470), .RSTB(I5819), .Q(I6037) );
nor I_267 (I6054,I6037,I5918);
nand I_268 (I5805,I5952,I6054);
not I_269 (I5802,I6037);
and I_270 (I6099,I6037,I5935);
DFFARX1 I_271  ( .D(I6099), .CLK(I1470), .RSTB(I5819), .Q(I5787) );
DFFARX1 I_272  ( .D(I6037), .CLK(I1470), .RSTB(I5819), .Q(I6130) );
and I_273 (I5784,I5952,I6130);
nand I_274 (I6161,I5836,I1231);
not I_275 (I6178,I6161);
nor I_276 (I6195,I6037,I6178);
DFFARX1 I_277  ( .D(I1247), .CLK(I1470), .RSTB(I5819), .Q(I6212) );
nand I_278 (I6229,I6212,I6161);
and I_279 (I6246,I5952,I6229);
DFFARX1 I_280  ( .D(I6246), .CLK(I1470), .RSTB(I5819), .Q(I5811) );
not I_281 (I6277,I6212);
nand I_282 (I5799,I6212,I6195);
nand I_283 (I5793,I6212,I6178);
DFFARX1 I_284  ( .D(I1391), .CLK(I1470), .RSTB(I5819), .Q(I6322) );
not I_285 (I6339,I6322);
nor I_286 (I5808,I6212,I6339);
nor I_287 (I6370,I6339,I6277);
and I_288 (I6387,I5918,I6370);
or I_289 (I6404,I6161,I6387);
DFFARX1 I_290  ( .D(I6404), .CLK(I1470), .RSTB(I5819), .Q(I5796) );
DFFARX1 I_291  ( .D(I6339), .CLK(I1470), .RSTB(I5819), .Q(I5781) );
not I_292 (I6482,I1477);
or I_293 (I6499,I11408,I11423);
or I_294 (I6516,I11411,I11408);
DFFARX1 I_295  ( .D(I6516), .CLK(I1470), .RSTB(I6482), .Q(I6456) );
nor I_296 (I6547,I11414,I11429);
not I_297 (I6564,I6547);
not I_298 (I6581,I11414);
and I_299 (I6598,I6581,I11417);
nor I_300 (I6615,I6598,I11423);
nor I_301 (I6632,I11420,I11438);
DFFARX1 I_302  ( .D(I6632), .CLK(I1470), .RSTB(I6482), .Q(I6649) );
nand I_303 (I6666,I6649,I6499);
and I_304 (I6683,I6615,I6666);
DFFARX1 I_305  ( .D(I6683), .CLK(I1470), .RSTB(I6482), .Q(I6450) );
nor I_306 (I6714,I11420,I11411);
DFFARX1 I_307  ( .D(I6714), .CLK(I1470), .RSTB(I6482), .Q(I6731) );
and I_308 (I6447,I6547,I6731);
DFFARX1 I_309  ( .D(I11435), .CLK(I1470), .RSTB(I6482), .Q(I6762) );
and I_310 (I6779,I6762,I11426);
DFFARX1 I_311  ( .D(I6779), .CLK(I1470), .RSTB(I6482), .Q(I6796) );
not I_312 (I6459,I6796);
DFFARX1 I_313  ( .D(I6779), .CLK(I1470), .RSTB(I6482), .Q(I6444) );
DFFARX1 I_314  ( .D(I11432), .CLK(I1470), .RSTB(I6482), .Q(I6841) );
not I_315 (I6858,I6841);
nor I_316 (I6875,I6516,I6858);
and I_317 (I6892,I6779,I6875);
or I_318 (I6909,I6499,I6892);
DFFARX1 I_319  ( .D(I6909), .CLK(I1470), .RSTB(I6482), .Q(I6465) );
nor I_320 (I6940,I6841,I6649);
nand I_321 (I6474,I6615,I6940);
nor I_322 (I6971,I6841,I6564);
nand I_323 (I6468,I6714,I6971);
not I_324 (I6471,I6841);
nand I_325 (I6462,I6841,I6564);
DFFARX1 I_326  ( .D(I6841), .CLK(I1470), .RSTB(I6482), .Q(I6453) );
not I_327 (I7077,I1477);
or I_328 (I7094,I10745,I10760);
or I_329 (I7111,I10748,I10745);
DFFARX1 I_330  ( .D(I7111), .CLK(I1470), .RSTB(I7077), .Q(I7051) );
nor I_331 (I7142,I10751,I10766);
not I_332 (I7159,I7142);
not I_333 (I7176,I10751);
and I_334 (I7193,I7176,I10754);
nor I_335 (I7210,I7193,I10760);
nor I_336 (I7227,I10757,I10775);
DFFARX1 I_337  ( .D(I7227), .CLK(I1470), .RSTB(I7077), .Q(I7244) );
nand I_338 (I7261,I7244,I7094);
and I_339 (I7278,I7210,I7261);
DFFARX1 I_340  ( .D(I7278), .CLK(I1470), .RSTB(I7077), .Q(I7045) );
nor I_341 (I7309,I10757,I10748);
DFFARX1 I_342  ( .D(I7309), .CLK(I1470), .RSTB(I7077), .Q(I7326) );
and I_343 (I7042,I7142,I7326);
DFFARX1 I_344  ( .D(I10772), .CLK(I1470), .RSTB(I7077), .Q(I7357) );
and I_345 (I7374,I7357,I10763);
DFFARX1 I_346  ( .D(I7374), .CLK(I1470), .RSTB(I7077), .Q(I7391) );
not I_347 (I7054,I7391);
DFFARX1 I_348  ( .D(I7374), .CLK(I1470), .RSTB(I7077), .Q(I7039) );
DFFARX1 I_349  ( .D(I10769), .CLK(I1470), .RSTB(I7077), .Q(I7436) );
not I_350 (I7453,I7436);
nor I_351 (I7470,I7111,I7453);
and I_352 (I7487,I7374,I7470);
or I_353 (I7504,I7094,I7487);
DFFARX1 I_354  ( .D(I7504), .CLK(I1470), .RSTB(I7077), .Q(I7060) );
nor I_355 (I7535,I7436,I7244);
nand I_356 (I7069,I7210,I7535);
nor I_357 (I7566,I7436,I7159);
nand I_358 (I7063,I7309,I7566);
not I_359 (I7066,I7436);
nand I_360 (I7057,I7436,I7159);
DFFARX1 I_361  ( .D(I7436), .CLK(I1470), .RSTB(I7077), .Q(I7048) );
not I_362 (I7672,I1477);
or I_363 (I7689,I5811,I5796);
or I_364 (I7706,I5793,I5811);
DFFARX1 I_365  ( .D(I7706), .CLK(I1470), .RSTB(I7672), .Q(I7646) );
nor I_366 (I7737,I5781,I5790);
not I_367 (I7754,I7737);
not I_368 (I7771,I5781);
and I_369 (I7788,I7771,I5805);
nor I_370 (I7805,I7788,I5796);
nor I_371 (I7822,I5784,I5799);
DFFARX1 I_372  ( .D(I7822), .CLK(I1470), .RSTB(I7672), .Q(I7839) );
nand I_373 (I7856,I7839,I7689);
and I_374 (I7873,I7805,I7856);
DFFARX1 I_375  ( .D(I7873), .CLK(I1470), .RSTB(I7672), .Q(I7640) );
nor I_376 (I7904,I5784,I5793);
DFFARX1 I_377  ( .D(I7904), .CLK(I1470), .RSTB(I7672), .Q(I7921) );
and I_378 (I7637,I7737,I7921);
DFFARX1 I_379  ( .D(I5787), .CLK(I1470), .RSTB(I7672), .Q(I7952) );
and I_380 (I7969,I7952,I5808);
DFFARX1 I_381  ( .D(I7969), .CLK(I1470), .RSTB(I7672), .Q(I7986) );
not I_382 (I7649,I7986);
DFFARX1 I_383  ( .D(I7969), .CLK(I1470), .RSTB(I7672), .Q(I7634) );
DFFARX1 I_384  ( .D(I5802), .CLK(I1470), .RSTB(I7672), .Q(I8031) );
not I_385 (I8048,I8031);
nor I_386 (I8065,I7706,I8048);
and I_387 (I8082,I7969,I8065);
or I_388 (I8099,I7689,I8082);
DFFARX1 I_389  ( .D(I8099), .CLK(I1470), .RSTB(I7672), .Q(I7655) );
nor I_390 (I8130,I8031,I7839);
nand I_391 (I7664,I7805,I8130);
nor I_392 (I8161,I8031,I7754);
nand I_393 (I7658,I7904,I8161);
not I_394 (I7661,I8031);
nand I_395 (I7652,I8031,I7754);
DFFARX1 I_396  ( .D(I8031), .CLK(I1470), .RSTB(I7672), .Q(I7643) );
not I_397 (I8267,I1477);
or I_398 (I8284,I2062,I2071);
or I_399 (I8301,I2065,I2062);
DFFARX1 I_400  ( .D(I8301), .CLK(I1470), .RSTB(I8267), .Q(I8241) );
nor I_401 (I8332,I2041,I2044);
not I_402 (I8349,I8332);
not I_403 (I8366,I2041);
and I_404 (I8383,I8366,I2053);
nor I_405 (I8400,I8383,I2071);
nor I_406 (I8417,I2059,I2050);
DFFARX1 I_407  ( .D(I8417), .CLK(I1470), .RSTB(I8267), .Q(I8434) );
nand I_408 (I8451,I8434,I8284);
and I_409 (I8468,I8400,I8451);
DFFARX1 I_410  ( .D(I8468), .CLK(I1470), .RSTB(I8267), .Q(I8235) );
nor I_411 (I8499,I2059,I2065);
DFFARX1 I_412  ( .D(I8499), .CLK(I1470), .RSTB(I8267), .Q(I8516) );
and I_413 (I8232,I8332,I8516);
DFFARX1 I_414  ( .D(I2056), .CLK(I1470), .RSTB(I8267), .Q(I8547) );
and I_415 (I8564,I8547,I2047);
DFFARX1 I_416  ( .D(I8564), .CLK(I1470), .RSTB(I8267), .Q(I8581) );
not I_417 (I8244,I8581);
DFFARX1 I_418  ( .D(I8564), .CLK(I1470), .RSTB(I8267), .Q(I8229) );
DFFARX1 I_419  ( .D(I2068), .CLK(I1470), .RSTB(I8267), .Q(I8626) );
not I_420 (I8643,I8626);
nor I_421 (I8660,I8301,I8643);
and I_422 (I8677,I8564,I8660);
or I_423 (I8694,I8284,I8677);
DFFARX1 I_424  ( .D(I8694), .CLK(I1470), .RSTB(I8267), .Q(I8250) );
nor I_425 (I8725,I8626,I8434);
nand I_426 (I8259,I8400,I8725);
nor I_427 (I8756,I8626,I8349);
nand I_428 (I8253,I8499,I8756);
not I_429 (I8256,I8626);
nand I_430 (I8247,I8626,I8349);
DFFARX1 I_431  ( .D(I8626), .CLK(I1470), .RSTB(I8267), .Q(I8238) );
not I_432 (I8862,I1477);
or I_433 (I8879,I1375,I1223);
or I_434 (I8896,I1439,I1375);
DFFARX1 I_435  ( .D(I8896), .CLK(I1470), .RSTB(I8862), .Q(I8836) );
nor I_436 (I8927,I1335,I1319);
not I_437 (I8944,I8927);
not I_438 (I8961,I1335);
and I_439 (I8978,I8961,I1351);
nor I_440 (I8995,I8978,I1223);
nor I_441 (I9012,I1255,I1279);
DFFARX1 I_442  ( .D(I9012), .CLK(I1470), .RSTB(I8862), .Q(I9029) );
nand I_443 (I9046,I9029,I8879);
and I_444 (I9063,I8995,I9046);
DFFARX1 I_445  ( .D(I9063), .CLK(I1470), .RSTB(I8862), .Q(I8830) );
nor I_446 (I9094,I1255,I1439);
DFFARX1 I_447  ( .D(I9094), .CLK(I1470), .RSTB(I8862), .Q(I9111) );
and I_448 (I8827,I8927,I9111);
DFFARX1 I_449  ( .D(I1311), .CLK(I1470), .RSTB(I8862), .Q(I9142) );
and I_450 (I9159,I9142,I1295);
DFFARX1 I_451  ( .D(I9159), .CLK(I1470), .RSTB(I8862), .Q(I9176) );
not I_452 (I8839,I9176);
DFFARX1 I_453  ( .D(I9159), .CLK(I1470), .RSTB(I8862), .Q(I8824) );
DFFARX1 I_454  ( .D(I1463), .CLK(I1470), .RSTB(I8862), .Q(I9221) );
not I_455 (I9238,I9221);
nor I_456 (I9255,I8896,I9238);
and I_457 (I9272,I9159,I9255);
or I_458 (I9289,I8879,I9272);
DFFARX1 I_459  ( .D(I9289), .CLK(I1470), .RSTB(I8862), .Q(I8845) );
nor I_460 (I9320,I9221,I9029);
nand I_461 (I8854,I8995,I9320);
nor I_462 (I9351,I9221,I8944);
nand I_463 (I8848,I9094,I9351);
not I_464 (I8851,I9221);
nand I_465 (I8842,I9221,I8944);
DFFARX1 I_466  ( .D(I9221), .CLK(I1470), .RSTB(I8862), .Q(I8833) );
not I_467 (I9457,I1477);
not I_468 (I9474,I8842);
nor I_469 (I9491,I8836,I8827);
nand I_470 (I9508,I9491,I8839);
nor I_471 (I9525,I9474,I8836);
nand I_472 (I9542,I9525,I8854);
not I_473 (I9559,I9542);
not I_474 (I9576,I8836);
nor I_475 (I9446,I9542,I9576);
not I_476 (I9607,I9576);
nand I_477 (I9431,I9542,I9607);
not I_478 (I9638,I8830);
nor I_479 (I9655,I9638,I8824);
and I_480 (I9672,I9655,I8851);
or I_481 (I9689,I9672,I8848);
DFFARX1 I_482  ( .D(I9689), .CLK(I1470), .RSTB(I9457), .Q(I9706) );
nor I_483 (I9723,I9706,I9559);
DFFARX1 I_484  ( .D(I9706), .CLK(I1470), .RSTB(I9457), .Q(I9740) );
not I_485 (I9428,I9740);
nand I_486 (I9771,I9474,I8830);
and I_487 (I9788,I9771,I9723);
DFFARX1 I_488  ( .D(I9771), .CLK(I1470), .RSTB(I9457), .Q(I9425) );
DFFARX1 I_489  ( .D(I8845), .CLK(I1470), .RSTB(I9457), .Q(I9819) );
nor I_490 (I9836,I9819,I9542);
nand I_491 (I9443,I9706,I9836);
nor I_492 (I9867,I9819,I9607);
not I_493 (I9440,I9819);
nand I_494 (I9898,I9819,I9508);
and I_495 (I9915,I9576,I9898);
DFFARX1 I_496  ( .D(I9915), .CLK(I1470), .RSTB(I9457), .Q(I9419) );
DFFARX1 I_497  ( .D(I9819), .CLK(I1470), .RSTB(I9457), .Q(I9422) );
DFFARX1 I_498  ( .D(I8833), .CLK(I1470), .RSTB(I9457), .Q(I9960) );
not I_499 (I9977,I9960);
nand I_500 (I9994,I9977,I9542);
and I_501 (I10011,I9771,I9994);
DFFARX1 I_502  ( .D(I10011), .CLK(I1470), .RSTB(I9457), .Q(I9449) );
or I_503 (I10042,I9977,I9788);
DFFARX1 I_504  ( .D(I10042), .CLK(I1470), .RSTB(I9457), .Q(I9434) );
nand I_505 (I9437,I9977,I9867);
not I_506 (I10120,I1477);
not I_507 (I10137,I6462);
nor I_508 (I10154,I6456,I6447);
nand I_509 (I10171,I10154,I6459);
nor I_510 (I10188,I10137,I6456);
nand I_511 (I10205,I10188,I6474);
not I_512 (I10222,I10205);
not I_513 (I10239,I6456);
nor I_514 (I10109,I10205,I10239);
not I_515 (I10270,I10239);
nand I_516 (I10094,I10205,I10270);
not I_517 (I10301,I6450);
nor I_518 (I10318,I10301,I6444);
and I_519 (I10335,I10318,I6471);
or I_520 (I10352,I10335,I6468);
DFFARX1 I_521  ( .D(I10352), .CLK(I1470), .RSTB(I10120), .Q(I10369) );
nor I_522 (I10386,I10369,I10222);
DFFARX1 I_523  ( .D(I10369), .CLK(I1470), .RSTB(I10120), .Q(I10403) );
not I_524 (I10091,I10403);
nand I_525 (I10434,I10137,I6450);
and I_526 (I10451,I10434,I10386);
DFFARX1 I_527  ( .D(I10434), .CLK(I1470), .RSTB(I10120), .Q(I10088) );
DFFARX1 I_528  ( .D(I6465), .CLK(I1470), .RSTB(I10120), .Q(I10482) );
nor I_529 (I10499,I10482,I10205);
nand I_530 (I10106,I10369,I10499);
nor I_531 (I10530,I10482,I10270);
not I_532 (I10103,I10482);
nand I_533 (I10561,I10482,I10171);
and I_534 (I10578,I10239,I10561);
DFFARX1 I_535  ( .D(I10578), .CLK(I1470), .RSTB(I10120), .Q(I10082) );
DFFARX1 I_536  ( .D(I10482), .CLK(I1470), .RSTB(I10120), .Q(I10085) );
DFFARX1 I_537  ( .D(I6453), .CLK(I1470), .RSTB(I10120), .Q(I10623) );
not I_538 (I10640,I10623);
nand I_539 (I10657,I10640,I10205);
and I_540 (I10674,I10434,I10657);
DFFARX1 I_541  ( .D(I10674), .CLK(I1470), .RSTB(I10120), .Q(I10112) );
or I_542 (I10705,I10640,I10451);
DFFARX1 I_543  ( .D(I10705), .CLK(I1470), .RSTB(I10120), .Q(I10097) );
nand I_544 (I10100,I10640,I10530);
not I_545 (I10783,I1477);
not I_546 (I10800,I13375);
nor I_547 (I10817,I13372,I13390);
nand I_548 (I10834,I10817,I13393);
nor I_549 (I10851,I10800,I13372);
nand I_550 (I10868,I10851,I13378);
not I_551 (I10885,I10868);
not I_552 (I10902,I13372);
nor I_553 (I10772,I10868,I10902);
not I_554 (I10933,I10902);
nand I_555 (I10757,I10868,I10933);
not I_556 (I10964,I13387);
nor I_557 (I10981,I10964,I13369);
and I_558 (I10998,I10981,I13363);
or I_559 (I11015,I10998,I13381);
DFFARX1 I_560  ( .D(I11015), .CLK(I1470), .RSTB(I10783), .Q(I11032) );
nor I_561 (I11049,I11032,I10885);
DFFARX1 I_562  ( .D(I11032), .CLK(I1470), .RSTB(I10783), .Q(I11066) );
not I_563 (I10754,I11066);
nand I_564 (I11097,I10800,I13387);
and I_565 (I11114,I11097,I11049);
DFFARX1 I_566  ( .D(I11097), .CLK(I1470), .RSTB(I10783), .Q(I10751) );
DFFARX1 I_567  ( .D(I13366), .CLK(I1470), .RSTB(I10783), .Q(I11145) );
nor I_568 (I11162,I11145,I10868);
nand I_569 (I10769,I11032,I11162);
nor I_570 (I11193,I11145,I10933);
not I_571 (I10766,I11145);
nand I_572 (I11224,I11145,I10834);
and I_573 (I11241,I10902,I11224);
DFFARX1 I_574  ( .D(I11241), .CLK(I1470), .RSTB(I10783), .Q(I10745) );
DFFARX1 I_575  ( .D(I11145), .CLK(I1470), .RSTB(I10783), .Q(I10748) );
DFFARX1 I_576  ( .D(I13384), .CLK(I1470), .RSTB(I10783), .Q(I11286) );
not I_577 (I11303,I11286);
nand I_578 (I11320,I11303,I10868);
and I_579 (I11337,I11097,I11320);
DFFARX1 I_580  ( .D(I11337), .CLK(I1470), .RSTB(I10783), .Q(I10775) );
or I_581 (I11368,I11303,I11114);
DFFARX1 I_582  ( .D(I11368), .CLK(I1470), .RSTB(I10783), .Q(I10760) );
nand I_583 (I10763,I11303,I11193);
not I_584 (I11446,I1477);
not I_585 (I11463,I3815);
nor I_586 (I11480,I3812,I3836);
nand I_587 (I11497,I11480,I3833);
nor I_588 (I11514,I11463,I3812);
nand I_589 (I11531,I11514,I3839);
not I_590 (I11548,I11531);
not I_591 (I11565,I3812);
nor I_592 (I11435,I11531,I11565);
not I_593 (I11596,I11565);
nand I_594 (I11420,I11531,I11596);
not I_595 (I11627,I3830);
nor I_596 (I11644,I11627,I3821);
and I_597 (I11661,I11644,I3818);
or I_598 (I11678,I11661,I3827);
DFFARX1 I_599  ( .D(I11678), .CLK(I1470), .RSTB(I11446), .Q(I11695) );
nor I_600 (I11712,I11695,I11548);
DFFARX1 I_601  ( .D(I11695), .CLK(I1470), .RSTB(I11446), .Q(I11729) );
not I_602 (I11417,I11729);
nand I_603 (I11760,I11463,I3830);
and I_604 (I11777,I11760,I11712);
DFFARX1 I_605  ( .D(I11760), .CLK(I1470), .RSTB(I11446), .Q(I11414) );
DFFARX1 I_606  ( .D(I3809), .CLK(I1470), .RSTB(I11446), .Q(I11808) );
nor I_607 (I11825,I11808,I11531);
nand I_608 (I11432,I11695,I11825);
nor I_609 (I11856,I11808,I11596);
not I_610 (I11429,I11808);
nand I_611 (I11887,I11808,I11497);
and I_612 (I11904,I11565,I11887);
DFFARX1 I_613  ( .D(I11904), .CLK(I1470), .RSTB(I11446), .Q(I11408) );
DFFARX1 I_614  ( .D(I11808), .CLK(I1470), .RSTB(I11446), .Q(I11411) );
DFFARX1 I_615  ( .D(I3824), .CLK(I1470), .RSTB(I11446), .Q(I11949) );
not I_616 (I11966,I11949);
nand I_617 (I11983,I11966,I11531);
and I_618 (I12000,I11760,I11983);
DFFARX1 I_619  ( .D(I12000), .CLK(I1470), .RSTB(I11446), .Q(I11438) );
or I_620 (I12031,I11966,I11777);
DFFARX1 I_621  ( .D(I12031), .CLK(I1470), .RSTB(I11446), .Q(I11423) );
nand I_622 (I11426,I11966,I11856);
not I_623 (I12109,I1477);
not I_624 (I12126,I1489);
nor I_625 (I12143,I1504,I1498);
nand I_626 (I12160,I12143,I1507);
nor I_627 (I12177,I12126,I1504);
nand I_628 (I12194,I12177,I1483);
DFFARX1 I_629  ( .D(I12194), .CLK(I1470), .RSTB(I12109), .Q(I12211) );
not I_630 (I12080,I12211);
not I_631 (I12242,I1504);
not I_632 (I12259,I12242);
not I_633 (I12276,I1480);
nor I_634 (I12293,I12276,I1495);
and I_635 (I12310,I12293,I1501);
or I_636 (I12327,I12310,I1510);
DFFARX1 I_637  ( .D(I12327), .CLK(I1470), .RSTB(I12109), .Q(I12344) );
DFFARX1 I_638  ( .D(I12344), .CLK(I1470), .RSTB(I12109), .Q(I12077) );
DFFARX1 I_639  ( .D(I12344), .CLK(I1470), .RSTB(I12109), .Q(I12375) );
DFFARX1 I_640  ( .D(I12344), .CLK(I1470), .RSTB(I12109), .Q(I12071) );
nand I_641 (I12406,I12126,I1480);
nand I_642 (I12423,I12406,I12160);
and I_643 (I12440,I12242,I12423);
DFFARX1 I_644  ( .D(I12440), .CLK(I1470), .RSTB(I12109), .Q(I12101) );
and I_645 (I12074,I12406,I12375);
DFFARX1 I_646  ( .D(I1492), .CLK(I1470), .RSTB(I12109), .Q(I12485) );
nor I_647 (I12098,I12485,I12406);
nor I_648 (I12516,I12485,I12160);
nand I_649 (I12095,I12194,I12516);
not I_650 (I12092,I12485);
DFFARX1 I_651  ( .D(I1486), .CLK(I1470), .RSTB(I12109), .Q(I12561) );
not I_652 (I12578,I12561);
nor I_653 (I12595,I12578,I12259);
and I_654 (I12612,I12485,I12595);
or I_655 (I12629,I12406,I12612);
DFFARX1 I_656  ( .D(I12629), .CLK(I1470), .RSTB(I12109), .Q(I12086) );
not I_657 (I12660,I12578);
nor I_658 (I12677,I12485,I12660);
nand I_659 (I12089,I12578,I12677);
nand I_660 (I12083,I12242,I12660);
not I_661 (I12755,I1477);
not I_662 (I12772,I9443);
nor I_663 (I12789,I9422,I9434);
nand I_664 (I12806,I12789,I9437);
nor I_665 (I12823,I12772,I9422);
nand I_666 (I12840,I12823,I9419);
DFFARX1 I_667  ( .D(I12840), .CLK(I1470), .RSTB(I12755), .Q(I12857) );
not I_668 (I12726,I12857);
not I_669 (I12888,I9422);
not I_670 (I12905,I12888);
not I_671 (I12922,I9440);
nor I_672 (I12939,I12922,I9431);
and I_673 (I12956,I12939,I9425);
or I_674 (I12973,I12956,I9449);
DFFARX1 I_675  ( .D(I12973), .CLK(I1470), .RSTB(I12755), .Q(I12990) );
DFFARX1 I_676  ( .D(I12990), .CLK(I1470), .RSTB(I12755), .Q(I12723) );
DFFARX1 I_677  ( .D(I12990), .CLK(I1470), .RSTB(I12755), .Q(I13021) );
DFFARX1 I_678  ( .D(I12990), .CLK(I1470), .RSTB(I12755), .Q(I12717) );
nand I_679 (I13052,I12772,I9440);
nand I_680 (I13069,I13052,I12806);
and I_681 (I13086,I12888,I13069);
DFFARX1 I_682  ( .D(I13086), .CLK(I1470), .RSTB(I12755), .Q(I12747) );
and I_683 (I12720,I13052,I13021);
DFFARX1 I_684  ( .D(I9446), .CLK(I1470), .RSTB(I12755), .Q(I13131) );
nor I_685 (I12744,I13131,I13052);
nor I_686 (I13162,I13131,I12806);
nand I_687 (I12741,I12840,I13162);
not I_688 (I12738,I13131);
DFFARX1 I_689  ( .D(I9428), .CLK(I1470), .RSTB(I12755), .Q(I13207) );
not I_690 (I13224,I13207);
nor I_691 (I13241,I13224,I12905);
and I_692 (I13258,I13131,I13241);
or I_693 (I13275,I13052,I13258);
DFFARX1 I_694  ( .D(I13275), .CLK(I1470), .RSTB(I12755), .Q(I12732) );
not I_695 (I13306,I13224);
nor I_696 (I13323,I13131,I13306);
nand I_697 (I12735,I13224,I13323);
nand I_698 (I12729,I12888,I13306);
not I_699 (I13401,I1477);
not I_700 (I13418,I14018);
nor I_701 (I13435,I14030,I14024);
nand I_702 (I13452,I13435,I14009);
nor I_703 (I13469,I13418,I14030);
nand I_704 (I13486,I13469,I14036);
DFFARX1 I_705  ( .D(I13486), .CLK(I1470), .RSTB(I13401), .Q(I13503) );
not I_706 (I13372,I13503);
not I_707 (I13534,I14030);
not I_708 (I13551,I13534);
not I_709 (I13568,I14033);
nor I_710 (I13585,I13568,I14015);
and I_711 (I13602,I13585,I14012);
or I_712 (I13619,I13602,I14039);
DFFARX1 I_713  ( .D(I13619), .CLK(I1470), .RSTB(I13401), .Q(I13636) );
DFFARX1 I_714  ( .D(I13636), .CLK(I1470), .RSTB(I13401), .Q(I13369) );
DFFARX1 I_715  ( .D(I13636), .CLK(I1470), .RSTB(I13401), .Q(I13667) );
DFFARX1 I_716  ( .D(I13636), .CLK(I1470), .RSTB(I13401), .Q(I13363) );
nand I_717 (I13698,I13418,I14033);
nand I_718 (I13715,I13698,I13452);
and I_719 (I13732,I13534,I13715);
DFFARX1 I_720  ( .D(I13732), .CLK(I1470), .RSTB(I13401), .Q(I13393) );
and I_721 (I13366,I13698,I13667);
DFFARX1 I_722  ( .D(I14027), .CLK(I1470), .RSTB(I13401), .Q(I13777) );
nor I_723 (I13390,I13777,I13698);
nor I_724 (I13808,I13777,I13452);
nand I_725 (I13387,I13486,I13808);
not I_726 (I13384,I13777);
DFFARX1 I_727  ( .D(I14021), .CLK(I1470), .RSTB(I13401), .Q(I13853) );
not I_728 (I13870,I13853);
nor I_729 (I13887,I13870,I13551);
and I_730 (I13904,I13777,I13887);
or I_731 (I13921,I13698,I13904);
DFFARX1 I_732  ( .D(I13921), .CLK(I1470), .RSTB(I13401), .Q(I13378) );
not I_733 (I13952,I13870);
nor I_734 (I13969,I13777,I13952);
nand I_735 (I13381,I13870,I13969);
nand I_736 (I13375,I13534,I13952);
not I_737 (I14047,I1477);
nand I_738 (I14064,I17625,I17631);
and I_739 (I14081,I14064,I17622);
DFFARX1 I_740  ( .D(I14081), .CLK(I1470), .RSTB(I14047), .Q(I14098) );
nor I_741 (I14115,I17634,I17631);
nor I_742 (I14132,I14115,I14098);
not I_743 (I14030,I14115);
DFFARX1 I_744  ( .D(I17613), .CLK(I1470), .RSTB(I14047), .Q(I14163) );
not I_745 (I14180,I14163);
nor I_746 (I14197,I14115,I14180);
nand I_747 (I14033,I14163,I14132);
DFFARX1 I_748  ( .D(I14163), .CLK(I1470), .RSTB(I14047), .Q(I14015) );
nand I_749 (I14242,I17637,I17619);
and I_750 (I14259,I14242,I17628);
DFFARX1 I_751  ( .D(I14259), .CLK(I1470), .RSTB(I14047), .Q(I14276) );
nor I_752 (I14036,I14276,I14098);
nand I_753 (I14027,I14276,I14197);
DFFARX1 I_754  ( .D(I17643), .CLK(I1470), .RSTB(I14047), .Q(I14321) );
and I_755 (I14338,I14321,I17616);
DFFARX1 I_756  ( .D(I14338), .CLK(I1470), .RSTB(I14047), .Q(I14355) );
not I_757 (I14018,I14355);
nand I_758 (I14386,I14338,I14276);
and I_759 (I14403,I14098,I14386);
DFFARX1 I_760  ( .D(I14403), .CLK(I1470), .RSTB(I14047), .Q(I14009) );
DFFARX1 I_761  ( .D(I17640), .CLK(I1470), .RSTB(I14047), .Q(I14434) );
nand I_762 (I14451,I14434,I14098);
and I_763 (I14468,I14276,I14451);
DFFARX1 I_764  ( .D(I14468), .CLK(I1470), .RSTB(I14047), .Q(I14039) );
not I_765 (I14499,I14434);
nor I_766 (I14516,I14115,I14499);
and I_767 (I14533,I14434,I14516);
or I_768 (I14550,I14338,I14533);
DFFARX1 I_769  ( .D(I14550), .CLK(I1470), .RSTB(I14047), .Q(I14024) );
nand I_770 (I14021,I14434,I14180);
DFFARX1 I_771  ( .D(I14434), .CLK(I1470), .RSTB(I14047), .Q(I14012) );
not I_772 (I14642,I1477);
nand I_773 (I14659,I10100,I10106);
and I_774 (I14676,I14659,I10088);
DFFARX1 I_775  ( .D(I14676), .CLK(I1470), .RSTB(I14642), .Q(I14693) );
nor I_776 (I14710,I10082,I10106);
nor I_777 (I14727,I14710,I14693);
not I_778 (I14625,I14710);
DFFARX1 I_779  ( .D(I10112), .CLK(I1470), .RSTB(I14642), .Q(I14758) );
not I_780 (I14775,I14758);
nor I_781 (I14792,I14710,I14775);
nand I_782 (I14628,I14758,I14727);
DFFARX1 I_783  ( .D(I14758), .CLK(I1470), .RSTB(I14642), .Q(I14610) );
nand I_784 (I14837,I10103,I10094);
and I_785 (I14854,I14837,I10097);
DFFARX1 I_786  ( .D(I14854), .CLK(I1470), .RSTB(I14642), .Q(I14871) );
nor I_787 (I14631,I14871,I14693);
nand I_788 (I14622,I14871,I14792);
DFFARX1 I_789  ( .D(I10109), .CLK(I1470), .RSTB(I14642), .Q(I14916) );
and I_790 (I14933,I14916,I10085);
DFFARX1 I_791  ( .D(I14933), .CLK(I1470), .RSTB(I14642), .Q(I14950) );
not I_792 (I14613,I14950);
nand I_793 (I14981,I14933,I14871);
and I_794 (I14998,I14693,I14981);
DFFARX1 I_795  ( .D(I14998), .CLK(I1470), .RSTB(I14642), .Q(I14604) );
DFFARX1 I_796  ( .D(I10091), .CLK(I1470), .RSTB(I14642), .Q(I15029) );
nand I_797 (I15046,I15029,I14693);
and I_798 (I15063,I14871,I15046);
DFFARX1 I_799  ( .D(I15063), .CLK(I1470), .RSTB(I14642), .Q(I14634) );
not I_800 (I15094,I15029);
nor I_801 (I15111,I14710,I15094);
and I_802 (I15128,I15029,I15111);
or I_803 (I15145,I14933,I15128);
DFFARX1 I_804  ( .D(I15145), .CLK(I1470), .RSTB(I14642), .Q(I14619) );
nand I_805 (I14616,I15029,I14775);
DFFARX1 I_806  ( .D(I15029), .CLK(I1470), .RSTB(I14642), .Q(I14607) );
not I_807 (I15237,I1477);
nand I_808 (I15254,I2605,I2611);
and I_809 (I15271,I15254,I2608);
DFFARX1 I_810  ( .D(I15271), .CLK(I1470), .RSTB(I15237), .Q(I15288) );
nor I_811 (I15305,I2632,I2611);
nor I_812 (I15322,I15305,I15288);
not I_813 (I15220,I15305);
DFFARX1 I_814  ( .D(I2623), .CLK(I1470), .RSTB(I15237), .Q(I15353) );
not I_815 (I15370,I15353);
nor I_816 (I15387,I15305,I15370);
nand I_817 (I15223,I15353,I15322);
DFFARX1 I_818  ( .D(I15353), .CLK(I1470), .RSTB(I15237), .Q(I15205) );
nand I_819 (I15432,I2626,I2629);
and I_820 (I15449,I15432,I2602);
DFFARX1 I_821  ( .D(I15449), .CLK(I1470), .RSTB(I15237), .Q(I15466) );
nor I_822 (I15226,I15466,I15288);
nand I_823 (I15217,I15466,I15387);
DFFARX1 I_824  ( .D(I2620), .CLK(I1470), .RSTB(I15237), .Q(I15511) );
and I_825 (I15528,I15511,I2614);
DFFARX1 I_826  ( .D(I15528), .CLK(I1470), .RSTB(I15237), .Q(I15545) );
not I_827 (I15208,I15545);
nand I_828 (I15576,I15528,I15466);
and I_829 (I15593,I15288,I15576);
DFFARX1 I_830  ( .D(I15593), .CLK(I1470), .RSTB(I15237), .Q(I15199) );
DFFARX1 I_831  ( .D(I2617), .CLK(I1470), .RSTB(I15237), .Q(I15624) );
nand I_832 (I15641,I15624,I15288);
and I_833 (I15658,I15466,I15641);
DFFARX1 I_834  ( .D(I15658), .CLK(I1470), .RSTB(I15237), .Q(I15229) );
not I_835 (I15689,I15624);
nor I_836 (I15706,I15305,I15689);
and I_837 (I15723,I15624,I15706);
or I_838 (I15740,I15528,I15723);
DFFARX1 I_839  ( .D(I15740), .CLK(I1470), .RSTB(I15237), .Q(I15214) );
nand I_840 (I15211,I15624,I15370);
DFFARX1 I_841  ( .D(I15624), .CLK(I1470), .RSTB(I15237), .Q(I15202) );
not I_842 (I15832,I1477);
nand I_843 (I15849,I7649,I7646);
and I_844 (I15866,I15849,I7643);
DFFARX1 I_845  ( .D(I15866), .CLK(I1470), .RSTB(I15832), .Q(I15883) );
nor I_846 (I15900,I7634,I7646);
nor I_847 (I15917,I15900,I15883);
not I_848 (I15815,I15900);
DFFARX1 I_849  ( .D(I7652), .CLK(I1470), .RSTB(I15832), .Q(I15948) );
not I_850 (I15965,I15948);
nor I_851 (I15982,I15900,I15965);
nand I_852 (I15818,I15948,I15917);
DFFARX1 I_853  ( .D(I15948), .CLK(I1470), .RSTB(I15832), .Q(I15800) );
nand I_854 (I16027,I7637,I7661);
and I_855 (I16044,I16027,I7640);
DFFARX1 I_856  ( .D(I16044), .CLK(I1470), .RSTB(I15832), .Q(I16061) );
nor I_857 (I15821,I16061,I15883);
nand I_858 (I15812,I16061,I15982);
DFFARX1 I_859  ( .D(I7658), .CLK(I1470), .RSTB(I15832), .Q(I16106) );
and I_860 (I16123,I16106,I7655);
DFFARX1 I_861  ( .D(I16123), .CLK(I1470), .RSTB(I15832), .Q(I16140) );
not I_862 (I15803,I16140);
nand I_863 (I16171,I16123,I16061);
and I_864 (I16188,I15883,I16171);
DFFARX1 I_865  ( .D(I16188), .CLK(I1470), .RSTB(I15832), .Q(I15794) );
DFFARX1 I_866  ( .D(I7664), .CLK(I1470), .RSTB(I15832), .Q(I16219) );
nand I_867 (I16236,I16219,I15883);
and I_868 (I16253,I16061,I16236);
DFFARX1 I_869  ( .D(I16253), .CLK(I1470), .RSTB(I15832), .Q(I15824) );
not I_870 (I16284,I16219);
nor I_871 (I16301,I15900,I16284);
and I_872 (I16318,I16219,I16301);
or I_873 (I16335,I16123,I16318);
DFFARX1 I_874  ( .D(I16335), .CLK(I1470), .RSTB(I15832), .Q(I15809) );
nand I_875 (I15806,I16219,I15965);
DFFARX1 I_876  ( .D(I16219), .CLK(I1470), .RSTB(I15832), .Q(I15797) );
not I_877 (I16427,I1477);
nand I_878 (I16444,I15809,I15794);
and I_879 (I16461,I16444,I15800);
DFFARX1 I_880  ( .D(I16461), .CLK(I1470), .RSTB(I16427), .Q(I16478) );
nor I_881 (I16495,I15803,I15794);
DFFARX1 I_882  ( .D(I15815), .CLK(I1470), .RSTB(I16427), .Q(I16512) );
nand I_883 (I16529,I16512,I16495);
DFFARX1 I_884  ( .D(I16512), .CLK(I1470), .RSTB(I16427), .Q(I16398) );
nand I_885 (I16560,I15806,I15797);
and I_886 (I16577,I16560,I15824);
DFFARX1 I_887  ( .D(I16577), .CLK(I1470), .RSTB(I16427), .Q(I16594) );
not I_888 (I16611,I16594);
nor I_889 (I16628,I16478,I16611);
and I_890 (I16645,I16495,I16628);
and I_891 (I16662,I16594,I16529);
DFFARX1 I_892  ( .D(I16662), .CLK(I1470), .RSTB(I16427), .Q(I16395) );
DFFARX1 I_893  ( .D(I16594), .CLK(I1470), .RSTB(I16427), .Q(I16389) );
DFFARX1 I_894  ( .D(I15812), .CLK(I1470), .RSTB(I16427), .Q(I16707) );
and I_895 (I16724,I16707,I15818);
nand I_896 (I16741,I16724,I16594);
nor I_897 (I16416,I16724,I16495);
not I_898 (I16772,I16724);
nor I_899 (I16789,I16478,I16772);
nand I_900 (I16407,I16512,I16789);
nand I_901 (I16401,I16594,I16772);
or I_902 (I16834,I16724,I16645);
DFFARX1 I_903  ( .D(I16834), .CLK(I1470), .RSTB(I16427), .Q(I16404) );
DFFARX1 I_904  ( .D(I15821), .CLK(I1470), .RSTB(I16427), .Q(I16865) );
and I_905 (I16882,I16865,I16741);
DFFARX1 I_906  ( .D(I16882), .CLK(I1470), .RSTB(I16427), .Q(I16419) );
nor I_907 (I16913,I16865,I16478);
nand I_908 (I16413,I16724,I16913);
not I_909 (I16410,I16865);
DFFARX1 I_910  ( .D(I16865), .CLK(I1470), .RSTB(I16427), .Q(I16958) );
and I_911 (I16392,I16865,I16958);
not I_912 (I17022,I1477);
not I_913 (I17039,I7069);
nor I_914 (I17056,I7045,I7060);
nand I_915 (I17073,I17056,I7042);
nor I_916 (I17090,I17039,I7045);
nand I_917 (I17107,I17090,I7057);
not I_918 (I17124,I7045);
not I_919 (I17141,I17124);
not I_920 (I17158,I7048);
nor I_921 (I17175,I17158,I7063);
and I_922 (I17192,I17175,I7054);
or I_923 (I17209,I17192,I7039);
DFFARX1 I_924  ( .D(I17209), .CLK(I1470), .RSTB(I17022), .Q(I17226) );
nand I_925 (I17243,I17039,I7048);
or I_926 (I17011,I17243,I17226);
not I_927 (I17274,I17243);
nor I_928 (I17291,I17226,I17274);
and I_929 (I17308,I17124,I17291);
nand I_930 (I16984,I17243,I17141);
DFFARX1 I_931  ( .D(I7051), .CLK(I1470), .RSTB(I17022), .Q(I17339) );
or I_932 (I17005,I17339,I17226);
nor I_933 (I17370,I17339,I17107);
nor I_934 (I17387,I17339,I17141);
nand I_935 (I16990,I17073,I17387);
or I_936 (I17418,I17339,I17308);
DFFARX1 I_937  ( .D(I17418), .CLK(I1470), .RSTB(I17022), .Q(I16987) );
not I_938 (I16993,I17339);
DFFARX1 I_939  ( .D(I7066), .CLK(I1470), .RSTB(I17022), .Q(I17463) );
not I_940 (I17480,I17463);
nor I_941 (I17497,I17480,I17073);
DFFARX1 I_942  ( .D(I17497), .CLK(I1470), .RSTB(I17022), .Q(I16999) );
nor I_943 (I17014,I17339,I17480);
nor I_944 (I17002,I17480,I17243);
not I_945 (I17556,I17480);
and I_946 (I17573,I17107,I17556);
nor I_947 (I17008,I17243,I17573);
nand I_948 (I16996,I17480,I17370);
not I_949 (I17651,I1477);
nand I_950 (I17668,I3184,I3169);
and I_951 (I17685,I17668,I3163);
DFFARX1 I_952  ( .D(I17685), .CLK(I1470), .RSTB(I17651), .Q(I17702) );
not I_953 (I17640,I17702);
DFFARX1 I_954  ( .D(I17702), .CLK(I1470), .RSTB(I17651), .Q(I17733) );
not I_955 (I17628,I17733);
nor I_956 (I17764,I3190,I3169);
not I_957 (I17781,I17764);
nor I_958 (I17798,I17702,I17781);
DFFARX1 I_959  ( .D(I3193), .CLK(I1470), .RSTB(I17651), .Q(I17815) );
not I_960 (I17832,I17815);
nand I_961 (I17631,I17815,I17781);
DFFARX1 I_962  ( .D(I17815), .CLK(I1470), .RSTB(I17651), .Q(I17863) );
and I_963 (I17616,I17702,I17863);
nand I_964 (I17894,I3175,I3178);
and I_965 (I17911,I17894,I3181);
DFFARX1 I_966  ( .D(I17911), .CLK(I1470), .RSTB(I17651), .Q(I17928) );
nor I_967 (I17945,I17928,I17832);
and I_968 (I17962,I17764,I17945);
nor I_969 (I17979,I17928,I17702);
DFFARX1 I_970  ( .D(I17928), .CLK(I1470), .RSTB(I17651), .Q(I17622) );
DFFARX1 I_971  ( .D(I3187), .CLK(I1470), .RSTB(I17651), .Q(I18010) );
and I_972 (I18027,I18010,I3172);
or I_973 (I18044,I18027,I17962);
DFFARX1 I_974  ( .D(I18044), .CLK(I1470), .RSTB(I17651), .Q(I17634) );
nand I_975 (I17643,I18027,I17979);
DFFARX1 I_976  ( .D(I18027), .CLK(I1470), .RSTB(I17651), .Q(I17613) );
DFFARX1 I_977  ( .D(I3166), .CLK(I1470), .RSTB(I17651), .Q(I18103) );
nand I_978 (I17637,I18103,I17798);
DFFARX1 I_979  ( .D(I18103), .CLK(I1470), .RSTB(I17651), .Q(I17625) );
nand I_980 (I18148,I18103,I17764);
and I_981 (I18165,I17815,I18148);
DFFARX1 I_982  ( .D(I18165), .CLK(I1470), .RSTB(I17651), .Q(I17619) );
endmodule


