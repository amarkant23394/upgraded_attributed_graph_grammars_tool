module test_final(G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_3,blif_reset_net_1_r_3,G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3);
input G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_3,blif_reset_net_1_r_3;
output G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3;
wire G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7,n_431_0_l_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n4_1_l_3,n9_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3;
DFFARX1 I_0(n4_1_r_7,blif_clk_net_1_r_3,n9_3,G42_1_r_7,);
nor I_1(n_572_1_r_7,n30_7,n31_7);
nand I_2(n_573_1_r_7,IN_7_0_l_7,n28_7);
nor I_3(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_4(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_5(N1_4_r_7,blif_clk_net_1_r_3,n9_3,G199_4_r_7,);
DFFARX1 I_6(n26_7,blif_clk_net_1_r_3,n9_3,G214_4_r_7,);
DFFARX1 I_7(n5_7,blif_clk_net_1_r_3,n9_3,ACVQN1_5_r_7,);
not I_8(P6_5_r_7,P6_5_r_internal_7);
or I_9(n_431_0_l_7,IN_8_0_l_7,n36_7);
DFFARX1 I_10(n_431_0_l_7,blif_clk_net_1_r_3,n9_3,n43_7,);
not I_11(n27_7,n43_7);
DFFARX1 I_12(IN_2_5_l_7,blif_clk_net_1_r_3,n9_3,ACVQN1_5_l_7,);
DFFARX1 I_13(IN_1_5_l_7,blif_clk_net_1_r_3,n9_3,n44_7,);
nor I_14(n4_1_r_7,n30_7,n38_7);
nor I_15(N1_4_r_7,n27_7,n40_7);
nand I_16(n26_7,IN_11_0_l_7,n39_7);
not I_17(n5_7,G2_0_l_7);
DFFARX1 I_18(ACVQN1_5_l_7,blif_clk_net_1_r_3,n9_3,P6_5_r_internal_7,);
nor I_19(n28_7,n26_7,n29_7);
not I_20(n29_7,IN_5_0_l_7);
not I_21(n30_7,G1_0_l_7);
nand I_22(n31_7,n27_7,n29_7);
nor I_23(n32_7,ACVQN1_5_l_7,n34_7);
nor I_24(n33_7,G2_0_l_7,n29_7);
not I_25(n34_7,IN_7_0_l_7);
nor I_26(n35_7,n43_7,n44_7);
and I_27(n36_7,IN_2_0_l_7,n37_7);
nor I_28(n37_7,IN_4_0_l_7,n30_7);
nand I_29(n38_7,G2_0_l_7,n29_7);
nor I_30(n39_7,G2_0_l_7,IN_10_0_l_7);
nor I_31(n40_7,n44_7,n41_7);
nor I_32(n41_7,n34_7,n42_7);
nand I_33(n42_7,IN_5_0_l_7,n5_7);
DFFARX1 I_34(n4_1_r_3,blif_clk_net_1_r_3,n9_3,G42_1_r_3,);
nor I_35(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_36(n_573_1_r_3,n26_3,n27_3);
nor I_37(n_549_1_r_3,n40_3,n32_3);
nand I_38(n_569_1_r_3,n27_3,n31_3);
and I_39(n_452_1_r_3,n26_3,ACVQN1_5_r_7);
nor I_40(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_41(N3_2_r_3,blif_clk_net_1_r_3,n9_3,G199_2_r_3,);
DFFARX1 I_42(n_572_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_3,);
nor I_43(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_44(n4_1_l_3,G42_1_r_7,ACVQN1_5_r_7);
not I_45(n9_3,blif_reset_net_1_r_3);
DFFARX1 I_46(n4_1_l_3,blif_clk_net_1_r_3,n9_3,G42_1_l_3,);
not I_47(n22_3,G42_1_l_3);
DFFARX1 I_48(G214_4_r_7,blif_clk_net_1_r_3,n9_3,n40_3,);
DFFARX1 I_49(n_569_1_r_7,blif_clk_net_1_r_3,n9_3,n25_internal_3,);
not I_50(n25_3,n25_internal_3);
nor I_51(n4_1_r_3,n40_3,n36_3);
nor I_52(N3_2_r_3,n26_3,n37_3);
nor I_53(n_572_1_l_3,n_549_1_r_7,n_572_1_r_7);
DFFARX1 I_54(G42_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN1_3_r_3,);
nor I_55(n26_3,G199_4_r_7,P6_5_r_7);
not I_56(n27_3,G42_1_r_7);
nor I_57(n28_3,n29_3,G42_1_r_7);
nor I_58(n29_3,n30_3,n_549_1_r_7);
not I_59(n30_3,n_573_1_r_7);
nor I_60(n31_3,n40_3,P6_5_r_7);
nor I_61(n32_3,n25_3,n33_3);
nand I_62(n33_3,n22_3,n_572_1_r_7);
or I_63(n34_3,P6_5_r_7,G42_1_r_7);
nand I_64(n35_3,ACVQN1_3_r_3,n_572_1_r_7);
nor I_65(n36_3,G199_4_r_7,ACVQN1_5_r_7);
nor I_66(n37_3,n38_3,n39_3);
not I_67(n38_3,n_572_1_l_3);
nand I_68(n39_3,n27_3,n30_3);
endmodule


