module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_5_r_15,blif_reset_net_5_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15);
input IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_5_r_15,blif_reset_net_5_r_15;
output N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15;
wire N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14,I_BUFF_1_9_r_14,N3_8_l_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14,N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,n_102_5_r_15,n_431_5_r_15,n9_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15;
nor I_0(N1371_0_r_14,n47_14,n30_14);
nor I_1(N1508_0_r_14,n30_14,n41_14);
nor I_2(N1507_6_r_14,n37_14,n44_14);
nor I_3(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_4(n4_7_r_14,blif_clk_net_5_r_15,n9_15,G42_7_r_14,);
nor I_5(n_572_7_r_14,n28_14,n29_14);
nand I_6(n_573_7_r_14,n26_14,n27_14);
nor I_7(n_549_7_r_14,n31_14,n32_14);
nand I_8(n_569_7_r_14,n26_14,n30_14);
nor I_9(n_452_7_r_14,n47_14,n28_14);
nor I_10(N6147_9_r_14,n36_14,n37_14);
nor I_11(N6134_9_r_14,n28_14,n36_14);
not I_12(I_BUFF_1_9_r_14,n26_14);
and I_13(N3_8_l_14,IN_6_8_l_14,n38_14);
DFFARX1 I_14(N3_8_l_14,blif_clk_net_5_r_15,n9_15,n47_14,);
nor I_15(n4_7_r_14,n47_14,n35_14);
nand I_16(n26_14,IN_1_10_l_14,IN_2_10_l_14);
not I_17(n27_14,n28_14);
nor I_18(n28_14,IN_2_0_l_14,n43_14);
not I_19(n29_14,n33_14);
not I_20(n30_14,n31_14);
nor I_21(n31_14,IN_1_3_l_14,n46_14);
and I_22(n32_14,n33_14,n34_14);
nand I_23(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_24(n34_14,n42_14,n43_14);
nor I_25(n35_14,IN_1_8_l_14,IN_3_8_l_14);
nor I_26(n36_14,n47_14,n34_14);
not I_27(n37_14,n35_14);
nand I_28(n38_14,IN_2_8_l_14,IN_3_8_l_14);
nand I_29(n39_14,n29_14,n40_14);
nand I_30(n40_14,n27_14,n37_14);
nor I_31(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_32(n42_14,IN_3_0_l_14,IN_4_0_l_14);
not I_33(n43_14,IN_1_0_l_14);
nor I_34(n44_14,n27_14,n33_14);
or I_35(n45_14,IN_3_10_l_14,IN_4_10_l_14);
or I_36(n46_14,IN_2_3_l_14,IN_3_3_l_14);
and I_37(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_38(N1508_0_r_15,n55_15,N1508_0_r_14);
nor I_39(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_40(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_41(N1372_4_r_15,n39_15);
nor I_42(N1508_4_r_15,n39_15,n43_15);
nand I_43(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_44(n_431_5_r_15,blif_clk_net_5_r_15,n9_15,G78_5_r_15,);
nand I_45(n_576_5_r_15,n31_15,n32_15);
not I_46(n_102_5_r_15,n33_15);
nand I_47(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_48(N1507_6_r_15,n42_15,n46_15);
nand I_49(N1508_6_r_15,n39_15,n40_15);
nand I_50(n_431_5_r_15,n36_15,n37_15);
not I_51(n9_15,blif_reset_net_5_r_15);
nor I_52(n31_15,n33_15,n34_15);
nor I_53(n32_15,n44_15,n_549_7_r_14);
nor I_54(n33_15,n54_15,n55_15);
nand I_55(n34_15,n49_15,n_569_7_r_14);
nand I_56(n35_15,N1508_0_r_14,N1507_6_r_14);
not I_57(n36_15,n32_15);
nand I_58(n37_15,n34_15,n38_15);
not I_59(n38_15,n46_15);
nand I_60(n39_15,n38_15,n41_15);
nand I_61(n40_15,n41_15,n42_15);
and I_62(n41_15,n51_15,N1507_6_r_14);
and I_63(n42_15,n47_15,N1508_0_r_14);
and I_64(n43_15,n34_15,n36_15);
or I_65(n44_15,N1371_0_r_14,n_573_7_r_14);
not I_66(n45_15,N1372_1_r_15);
nand I_67(n46_15,n53_15,N1508_0_r_14);
nor I_68(n47_15,n34_15,n48_15);
not I_69(n48_15,N1507_6_r_14);
and I_70(n49_15,n50_15,N6134_9_r_14);
nand I_71(n50_15,n51_15,n52_15);
nand I_72(n51_15,N6147_9_r_14,N1371_0_r_14);
not I_73(n52_15,N1507_6_r_14);
nor I_74(n53_15,n48_15,N1508_6_r_14);
nor I_75(n54_15,n_572_7_r_14,n_452_7_r_14);
not I_76(n55_15,G42_7_r_14);
endmodule


