module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_8_r_10,n11_10,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
nor I_35(N1371_0_r_10,n37_10,n38_10);
nor I_36(N1508_0_r_10,n37_10,n58_10);
nand I_37(N6147_2_r_10,n39_10,n40_10);
not I_38(N6147_3_r_10,n39_10);
nor I_39(N1372_4_r_10,n46_10,n49_10);
nor I_40(N1508_4_r_10,n51_10,n52_10);
nor I_41(N1507_6_r_10,n49_10,n60_10);
nor I_42(N1508_6_r_10,n49_10,n50_10);
nor I_43(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_44(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_45(N6147_9_r_10,n36_10,n37_10);
nor I_46(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_47(I_BUFF_1_9_r_10,n48_10);
nor I_48(N3_8_r_10,n44_10,n47_10);
not I_49(n11_10,blif_reset_net_8_r_10);
not I_50(n35_10,n49_10);
nor I_51(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_52(n37_10,G42_7_r_4);
not I_53(n38_10,n46_10);
nand I_54(n39_10,n43_10,n44_10);
nand I_55(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_56(n41_10,n42_10,G42_7_r_4);
not I_57(n42_10,n44_10);
nor I_58(n43_10,n45_10,G42_7_r_4);
nand I_59(n44_10,n54_10,N1371_0_r_4);
nor I_60(n45_10,n59_10,N1508_6_r_4);
nand I_61(n46_10,n61_10,N1371_0_r_4);
nor I_62(n47_10,n46_10,n48_10);
nand I_63(n48_10,n62_10,n63_10);
nand I_64(n49_10,n56_10,n_549_7_r_4);
not I_65(n50_10,n45_10);
nor I_66(n51_10,n42_10,n53_10);
not I_67(n52_10,N1372_4_r_10);
nor I_68(n53_10,n48_10,n50_10);
and I_69(n54_10,n55_10,n_452_7_r_4);
nand I_70(n55_10,n56_10,n57_10);
nand I_71(n56_10,N1507_6_r_4,N1508_6_r_4);
not I_72(n57_10,n_549_7_r_4);
nor I_73(n58_10,n35_10,n45_10);
nor I_74(n59_10,n_572_7_r_4,n_569_7_r_4);
nor I_75(n60_10,n37_10,n46_10);
or I_76(n61_10,n_572_7_r_4,n_569_7_r_4);
nor I_77(n62_10,N1507_6_r_4,n_572_7_r_4);
or I_78(n63_10,n64_10,n_549_7_r_4);
nor I_79(n64_10,N6134_9_r_4,G42_7_r_4);
endmodule


