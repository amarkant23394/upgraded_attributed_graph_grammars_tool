module test_I1304(I1247,I1279,I1294,I1271,I1301,I1304);
input I1247,I1279,I1294,I1271,I1301;
output I1304;
wire I1342,I1475,I1509,I1492;
not I_0(I1342,I1301);
nand I_1(I1475,I1247,I1271);
DFFARX1 I_2(I1492,I1294,I1342,,,I1509,);
DFFARX1 I_3(I1509,I1294,I1342,,,I1304,);
and I_4(I1492,I1475,I1279);
endmodule


