module test_final(G18_1_l_0,G15_1_l_0,IN_1_1_l_0,IN_4_1_l_0,IN_5_1_l_0,IN_7_1_l_0,IN_9_1_l_0,IN_10_1_l_0,IN_1_3_l_0,IN_2_3_l_0,IN_4_3_l_0,blif_clk_net_1_r_17,blif_reset_net_1_r_17,G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17);
input G18_1_l_0,G15_1_l_0,IN_1_1_l_0,IN_4_1_l_0,IN_5_1_l_0,IN_7_1_l_0,IN_9_1_l_0,IN_10_1_l_0,IN_1_3_l_0,IN_2_3_l_0,IN_4_3_l_0,blif_clk_net_1_r_17,blif_reset_net_1_r_17;
output G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17;
wire G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_569_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0,n4_1_l_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n_431_0_l_17,n6_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17;
DFFARX1 I_0(n4_1_r_0,blif_clk_net_1_r_17,n6_17,G42_1_r_0,);
nor I_1(n_572_1_r_0,IN_5_1_l_0,n23_0);
nand I_2(n_573_1_r_0,n21_0,n22_0);
nand I_3(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_4(n_569_1_r_0,n21_0,n26_0);
nor I_5(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_6(N3_2_r_0,blif_clk_net_1_r_17,n6_17,G199_2_r_0,);
DFFARX1 I_7(N1_4_r_0,blif_clk_net_1_r_17,n6_17,G199_4_r_0,);
DFFARX1 I_8(n2_0,blif_clk_net_1_r_17,n6_17,G214_4_r_0,);
nor I_9(n4_1_l_0,G18_1_l_0,IN_1_1_l_0);
DFFARX1 I_10(n4_1_l_0,blif_clk_net_1_r_17,n6_17,n37_0,);
DFFARX1 I_11(IN_1_3_l_0,blif_clk_net_1_r_17,n6_17,n38_0,);
not I_12(n20_0,n38_0);
DFFARX1 I_13(IN_2_3_l_0,blif_clk_net_1_r_17,n6_17,ACVQN1_3_l_0,);
nor I_14(n4_1_r_0,IN_10_1_l_0,n23_0);
nor I_15(N3_2_r_0,n31_0,n32_0);
nor I_16(N1_4_r_0,n29_0,n32_0);
not I_17(n2_0,n31_0);
nor I_18(n21_0,IN_9_1_l_0,n37_0);
not I_19(n22_0,IN_5_1_l_0);
nand I_20(n23_0,n20_0,n30_0);
nand I_21(n24_0,n38_0,n25_0);
nor I_22(n25_0,IN_9_1_l_0,IN_10_1_l_0);
not I_23(n26_0,IN_10_1_l_0);
not I_24(n27_0,n29_0);
nor I_25(n28_0,G15_1_l_0,IN_7_1_l_0);
nand I_26(n29_0,n26_0,n33_0);
not I_27(n30_0,IN_9_1_l_0);
nand I_28(n31_0,IN_4_3_l_0,ACVQN1_3_l_0);
and I_29(n32_0,n35_0,n36_0);
nand I_30(n33_0,IN_4_1_l_0,n34_0);
not I_31(n34_0,G15_1_l_0);
nor I_32(n35_0,G18_1_l_0,G15_1_l_0);
nor I_33(n36_0,IN_5_1_l_0,IN_7_1_l_0);
DFFARX1 I_34(n4_1_r_17,blif_clk_net_1_r_17,n6_17,G42_1_r_17,);
nor I_35(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_36(n_573_1_r_17,n20_17,n21_17);
nand I_37(n_549_1_r_17,n23_17,n24_17);
nand I_38(n_569_1_r_17,n21_17,n22_17);
not I_39(n_452_1_r_17,n23_17);
DFFARX1 I_40(n19_17,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_17,);
nor I_41(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_42(N1_4_r_17,blif_clk_net_1_r_17,n6_17,G199_4_r_17,);
DFFARX1 I_43(n5_17,blif_clk_net_1_r_17,n6_17,G214_4_r_17,);
or I_44(n_431_0_l_17,n26_17,n_549_1_r_0);
not I_45(n6_17,blif_reset_net_1_r_17);
DFFARX1 I_46(n_431_0_l_17,blif_clk_net_1_r_17,n6_17,n20_internal_17,);
not I_47(n20_17,n20_internal_17);
DFFARX1 I_48(n_572_1_r_0,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_17,);
DFFARX1 I_49(G42_1_r_0,blif_clk_net_1_r_17,n6_17,n19_internal_17,);
not I_50(n19_17,n19_internal_17);
nor I_51(n4_1_r_17,n5_17,n25_17);
not I_52(n2_17,n29_17);
DFFARX1 I_53(n2_17,blif_clk_net_1_r_17,n6_17,n17_internal_17,);
not I_54(n17_17,n17_internal_17);
nor I_55(N1_4_r_17,n29_17,n31_17);
not I_56(n5_17,G199_4_r_0);
and I_57(n21_17,n32_17,n_573_1_r_0);
not I_58(n22_17,n25_17);
nand I_59(n23_17,n20_17,n22_17);
nand I_60(n24_17,n19_17,n22_17);
nand I_61(n25_17,n30_17,n_42_2_r_0);
and I_62(n26_17,n27_17,n_573_1_r_0);
nor I_63(n27_17,n28_17,G42_1_r_0);
not I_64(n28_17,G214_4_r_0);
nor I_65(n29_17,n28_17,n_572_1_r_0);
and I_66(n30_17,n5_17,n_572_1_r_0);
nor I_67(n31_17,n21_17,G199_4_r_0);
nor I_68(n32_17,G199_2_r_0,G199_4_r_0);
endmodule


