module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_8_r_8,blif_reset_net_8_r_8,N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_8_r_8,blif_reset_net_8_r_8;
output N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8;
wire N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,I_BUFF_1_9_r_6,N1372_10_r_6,N1508_10_r_6,N3_8_r_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6,N1508_0_r_8,N1372_1_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N3_8_l_8,n8_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8;
nor I_0(N1371_0_r_6,n30_6,n33_6);
nor I_1(N1508_0_r_6,n33_6,n44_6);
not I_2(N1372_1_r_6,n41_6);
nor I_3(N1508_1_r_6,n40_6,n41_6);
nor I_4(N1507_6_r_6,n39_6,n45_6);
nor I_5(N1508_6_r_6,n37_6,n38_6);
nor I_6(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_7(N3_8_r_6,blif_clk_net_8_r_8,n8_8,G199_8_r_6,);
nor I_8(N6147_9_r_6,n32_6,n33_6);
nor I_9(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_10(I_BUFF_1_9_r_6,n37_6);
not I_11(N1372_10_r_6,n43_6);
nor I_12(N1508_10_r_6,n42_6,n43_6);
nor I_13(N3_8_r_6,IN_1_9_l_6,n36_6);
nor I_14(n30_6,IN_5_9_l_6,n53_6);
not I_15(n31_6,n36_6);
nor I_16(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_17(n33_6,IN_1_9_l_6);
not I_18(n34_6,n35_6);
nand I_19(n35_6,IN_2_6_l_6,n49_6);
nand I_20(n36_6,IN_5_6_l_6,n51_6);
nand I_21(n37_6,IN_2_9_l_6,n54_6);
or I_22(n38_6,n35_6,n39_6);
nor I_23(n39_6,n40_6,n45_6);
and I_24(n40_6,n46_6,n47_6);
nand I_25(n41_6,n30_6,n31_6);
nor I_26(n42_6,n34_6,n40_6);
nand I_27(n43_6,IN_1_9_l_6,n30_6);
nor I_28(n44_6,n31_6,n40_6);
nor I_29(n45_6,n35_6,n36_6);
nor I_30(n46_6,IN_1_2_l_6,IN_2_2_l_6);
or I_31(n47_6,IN_5_2_l_6,n48_6);
nor I_32(n48_6,IN_3_2_l_6,IN_4_2_l_6);
and I_33(n49_6,IN_1_6_l_6,n50_6);
nand I_34(n50_6,n51_6,n52_6);
nand I_35(n51_6,IN_3_6_l_6,IN_4_6_l_6);
not I_36(n52_6,IN_5_6_l_6);
nor I_37(n53_6,IN_3_9_l_6,IN_4_9_l_6);
or I_38(n54_6,IN_3_9_l_6,IN_4_9_l_6);
nor I_39(N1371_0_r_8,n46_8,n51_8);
not I_40(N1508_0_r_8,n46_8);
nor I_41(N1372_1_r_8,n37_8,n49_8);
and I_42(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_43(N1507_6_r_8,n47_8,n48_8);
nor I_44(N1508_6_r_8,n37_8,n38_8);
nor I_45(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_46(N3_8_r_8,blif_clk_net_8_r_8,n8_8,G199_8_r_8,);
nor I_47(N6147_9_r_8,n29_8,n30_8);
nor I_48(N6134_9_r_8,n30_8,n31_8);
not I_49(I_BUFF_1_9_r_8,n35_8);
nor I_50(N1372_10_r_8,n46_8,n49_8);
nor I_51(N1508_10_r_8,n40_8,n41_8);
and I_52(N3_8_l_8,n36_8,N1507_6_r_6);
not I_53(n8_8,blif_reset_net_8_r_8);
DFFARX1 I_54(N3_8_l_8,blif_clk_net_8_r_8,n8_8,n53_8,);
not I_55(n29_8,n53_8);
nor I_56(N3_8_r_8,n33_8,n34_8);
and I_57(n30_8,n32_8,n33_8);
nor I_58(n31_8,N1508_1_r_6,N1508_6_r_6);
nand I_59(n32_8,n42_8,G199_8_r_6);
or I_60(n33_8,n46_8,N1371_0_r_6);
nor I_61(n34_8,n32_8,n35_8);
nand I_62(n35_8,n44_8,N1508_0_r_6);
nand I_63(n36_8,N1508_6_r_6,N6147_9_r_6);
not I_64(n37_8,n31_8);
nand I_65(n38_8,N1508_0_r_8,n39_8);
nand I_66(n39_8,n33_8,n50_8);
and I_67(n40_8,n32_8,n35_8);
not I_68(n41_8,N1372_10_r_8);
and I_69(n42_8,n43_8,N6134_9_r_6);
nand I_70(n43_8,n44_8,n45_8);
nand I_71(n44_8,N1508_0_r_6,N1372_10_r_6);
not I_72(n45_8,N1508_0_r_6);
nand I_73(n46_8,N1371_0_r_6,N1372_1_r_6);
not I_74(n47_8,n39_8);
nor I_75(n48_8,n35_8,n49_8);
not I_76(n49_8,n51_8);
nand I_77(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_78(n51_8,n52_8,n_42_8_r_6);
or I_79(n52_8,N1372_1_r_6,N1508_10_r_6);
endmodule


