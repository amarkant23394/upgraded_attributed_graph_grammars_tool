module test_I15730(I1470,I13775,I13843,I11944,I15730);
input I1470,I13775,I13843,I11944;
output I15730;
wire I13826,I13761,I15713,I13860,I13891;
DFFARX1 I_0(I1470,I13775,,,I13826,);
nand I_1(I13761,I13891,I13860);
not I_2(I15713,I13761);
not I_3(I15730,I15713);
nor I_4(I13860,I13843,I13826);
DFFARX1 I_5(I11944,I1470,I13775,,,I13891,);
endmodule


