module test_I6623(I3951,I3945,I1477,I1470,I4068,I4356,I6623);
input I3951,I3945,I1477,I1470,I4068,I4356;
output I6623;
wire I6606,I3960,I6510,I3966,I6589,I6329,I6493,I6572,I4034,I3983;
DFFARX1 I_0(I6589,I1470,I6329,,,I6606,);
DFFARX1 I_1(I4356,I1470,I3983,,,I3960,);
not I_2(I6510,I6493);
or I_3(I3966,I4068,I4034);
and I_4(I6589,I6572,I3960);
not I_5(I6329,I1477);
DFFARX1 I_6(I3966,I1470,I6329,,,I6493,);
nand I_7(I6572,I3951,I3945);
nor I_8(I6623,I6606,I6510);
DFFARX1 I_9(I1470,I3983,,,I4034,);
not I_10(I3983,I1477);
endmodule


