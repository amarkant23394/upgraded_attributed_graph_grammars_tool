module test_I10612(I1477,I1470,I10612);
input I1477,I1470;
output I10612;
wire I10647,I9491,I9816,I9468,I11009,I9621,I9864;
DFFARX1 I_0(I11009,I1470,I10647,,,I10612,);
not I_1(I10647,I1477);
not I_2(I9491,I1477);
DFFARX1 I_3(I1470,I9491,,,I9816,);
DFFARX1 I_4(I9864,I1470,I9491,,,I9468,);
DFFARX1 I_5(I9468,I1470,I10647,,,I11009,);
DFFARX1 I_6(I1470,I9491,,,I9621,);
nor I_7(I9864,I9816,I9621);
endmodule


