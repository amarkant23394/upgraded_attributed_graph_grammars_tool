module test_I6203(I2167,I2173,I1477,I1470,I2695,I6203);
input I2167,I2173,I1477,I1470,I2695;
output I6203;
wire I4629,I4518,I5751,I4869,I2149,I4544,I4674,I2181,I2155,I4691;
nor I_0(I4629,I2167,I2173);
DFFARX1 I_1(I4518,I1470,I5751,,,I6203,);
nand I_2(I4518,I4869,I4691);
not I_3(I5751,I1477);
DFFARX1 I_4(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_5(I2695,I1470,I2181,,,I2149,);
not I_6(I4544,I1477);
DFFARX1 I_7(I2155,I1470,I4544,,,I4674,);
not I_8(I2181,I1477);
DFFARX1 I_9(I1470,I2181,,,I2155,);
nor I_10(I4691,I4674,I4629);
endmodule


