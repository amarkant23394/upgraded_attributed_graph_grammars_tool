module test_I3388_rst(I1477_rst,I3388_rst);
,I3388_rst);
input I1477_rst;
output I3388_rst;
wire ;
not I_0(I3388_rst,I1477_rst);
endmodule


