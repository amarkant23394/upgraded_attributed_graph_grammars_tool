module test_final(G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_12,blif_reset_net_1_r_12,G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12);
input G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_12,blif_reset_net_1_r_12;
output G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12;
wire G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7,n_431_0_l_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n_431_0_l_12,n8_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12;
DFFARX1 I_0(n4_1_r_7,blif_clk_net_1_r_12,n8_12,G42_1_r_7,);
nor I_1(n_572_1_r_7,n30_7,n31_7);
nand I_2(n_573_1_r_7,IN_7_0_l_7,n28_7);
nor I_3(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_4(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_5(N1_4_r_7,blif_clk_net_1_r_12,n8_12,G199_4_r_7,);
DFFARX1 I_6(n26_7,blif_clk_net_1_r_12,n8_12,G214_4_r_7,);
DFFARX1 I_7(n5_7,blif_clk_net_1_r_12,n8_12,ACVQN1_5_r_7,);
not I_8(P6_5_r_7,P6_5_r_internal_7);
or I_9(n_431_0_l_7,IN_8_0_l_7,n36_7);
DFFARX1 I_10(n_431_0_l_7,blif_clk_net_1_r_12,n8_12,n43_7,);
not I_11(n27_7,n43_7);
DFFARX1 I_12(IN_2_5_l_7,blif_clk_net_1_r_12,n8_12,ACVQN1_5_l_7,);
DFFARX1 I_13(IN_1_5_l_7,blif_clk_net_1_r_12,n8_12,n44_7,);
nor I_14(n4_1_r_7,n30_7,n38_7);
nor I_15(N1_4_r_7,n27_7,n40_7);
nand I_16(n26_7,IN_11_0_l_7,n39_7);
not I_17(n5_7,G2_0_l_7);
DFFARX1 I_18(ACVQN1_5_l_7,blif_clk_net_1_r_12,n8_12,P6_5_r_internal_7,);
nor I_19(n28_7,n26_7,n29_7);
not I_20(n29_7,IN_5_0_l_7);
not I_21(n30_7,G1_0_l_7);
nand I_22(n31_7,n27_7,n29_7);
nor I_23(n32_7,ACVQN1_5_l_7,n34_7);
nor I_24(n33_7,G2_0_l_7,n29_7);
not I_25(n34_7,IN_7_0_l_7);
nor I_26(n35_7,n43_7,n44_7);
and I_27(n36_7,IN_2_0_l_7,n37_7);
nor I_28(n37_7,IN_4_0_l_7,n30_7);
nand I_29(n38_7,G2_0_l_7,n29_7);
nor I_30(n39_7,G2_0_l_7,IN_10_0_l_7);
nor I_31(n40_7,n44_7,n41_7);
nor I_32(n41_7,n34_7,n42_7);
nand I_33(n42_7,IN_5_0_l_7,n5_7);
DFFARX1 I_34(n4_1_r_12,blif_clk_net_1_r_12,n8_12,G42_1_r_12,);
nor I_35(n_572_1_r_12,n29_12,n30_12);
nand I_36(n_573_1_r_12,n26_12,n27_12);
nor I_37(n_549_1_r_12,n33_12,n34_12);
and I_38(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_39(N3_2_r_12,blif_clk_net_1_r_12,n8_12,G199_2_r_12,);
DFFARX1 I_40(n3_12,blif_clk_net_1_r_12,n8_12,ACVQN1_5_r_12,);
not I_41(P6_5_r_12,P6_5_r_internal_12);
or I_42(n_431_0_l_12,n36_12,n_572_1_r_7);
not I_43(n8_12,blif_reset_net_1_r_12);
DFFARX1 I_44(n_431_0_l_12,blif_clk_net_1_r_12,n8_12,n41_12,);
DFFARX1 I_45(G214_4_r_7,blif_clk_net_1_r_12,n8_12,ACVQN1_5_l_12,);
not I_46(n22_12,ACVQN1_5_l_12);
DFFARX1 I_47(G199_4_r_7,blif_clk_net_1_r_12,n8_12,n42_12,);
nor I_48(n4_1_r_12,n41_12,n31_12);
nor I_49(N3_2_r_12,n22_12,n40_12);
not I_50(n3_12,n39_12);
DFFARX1 I_51(ACVQN1_5_l_12,blif_clk_net_1_r_12,n8_12,P6_5_r_internal_12,);
and I_52(n26_12,P6_5_r_7,n_572_1_r_7);
nor I_53(n27_12,n28_12,n29_12);
not I_54(n28_12,n_549_1_r_7);
nand I_55(n29_12,n31_12,n32_12);
nand I_56(n30_12,n42_12,n_549_1_r_7);
not I_57(n31_12,G42_1_r_7);
not I_58(n32_12,ACVQN1_5_r_7);
nand I_59(n33_12,n31_12,n35_12);
nand I_60(n34_12,P6_5_r_7,n_572_1_r_7);
nand I_61(n35_12,n41_12,n42_12);
and I_62(n36_12,n37_12,n_569_1_r_7);
nor I_63(n37_12,n38_12,G42_1_r_7);
not I_64(n38_12,n_573_1_r_7);
nor I_65(n39_12,n38_12,P6_5_r_7);
nor I_66(n40_12,n39_12,G42_1_r_7);
endmodule


