module test_I17393(I15597,I1477,I1470,I16069,I17393);
input I15597,I1477,I1470,I16069;
output I17393;
wire I17563,I17413,I17916,I15959,I17775,I17532,I15603,I15585,I17933,I17823,I15928;
not I_0(I17563,I17532);
not I_1(I17413,I1477);
DFFARX1 I_2(I15603,I1470,I17413,,,I17916,);
nor I_3(I15959,I15928);
nand I_4(I17393,I17933,I17823);
DFFARX1 I_5(I15585,I1470,I17413,,,I17775,);
not I_6(I17532,I15597);
nor I_7(I15603,I15928,I16069);
nand I_8(I15585,I16069,I15959);
not I_9(I17933,I17916);
nor I_10(I17823,I17775,I17563);
DFFARX1 I_11(I1470,,,I15928,);
endmodule


