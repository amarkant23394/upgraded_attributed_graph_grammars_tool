module test_final(IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_3_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_4_4_l_2,IN_5_4_l_2,blif_clk_net_8_r_1,blif_reset_net_8_r_1,N6147_3_r_1,N1372_4_r_1,N1508_4_r_1,n_42_8_r_1,G199_8_r_1,N6147_9_r_1,N6134_9_r_1,N1372_10_r_1,N1508_10_r_1);
input IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_3_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_4_4_l_2,IN_5_4_l_2,blif_clk_net_8_r_1,blif_reset_net_8_r_1;
output N6147_3_r_1,N1372_4_r_1,N1508_4_r_1,n_42_8_r_1,G199_8_r_1,N6147_9_r_1,N6134_9_r_1,N1372_10_r_1,N1508_10_r_1;
wire N1371_0_r_2,N1508_0_r_2,N6147_3_r_2,n_429_or_0_5_r_2,G78_5_r_2,n_576_5_r_2,n_102_5_r_2,n_547_5_r_2,N1372_10_r_2,N1508_10_r_2,n_431_5_r_2,n21_2,n22_2,n23_2,n24_2,n25_2,n26_2,n27_2,n28_2,n29_2,n30_2,n31_2,n32_2,I_BUFF_1_9_r_1,N3_8_l_1,n7_1,n38_1,n22_1,N3_8_r_1,n23_1,n24_1,n25_1,n26_1,n27_1,n28_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1;
nor I_0(N1371_0_r_2,n23_2,n24_2);
not I_1(N1508_0_r_2,n24_2);
nor I_2(N6147_3_r_2,n22_2,n26_2);
nand I_3(n_429_or_0_5_r_2,IN_3_1_l_2,n22_2);
DFFARX1 I_4(n_431_5_r_2,blif_clk_net_8_r_1,n7_1,G78_5_r_2,);
nand I_5(n_576_5_r_2,n21_2,n22_2);
not I_6(n_102_5_r_2,n23_2);
nand I_7(n_547_5_r_2,n22_2,n24_2);
not I_8(N1372_10_r_2,n29_2);
nor I_9(N1508_10_r_2,n28_2,n29_2);
nand I_10(n_431_5_r_2,n_102_5_r_2,n25_2);
nor I_11(n21_2,IN_3_1_l_2,n23_2);
and I_12(n22_2,IN_1_1_l_2,IN_2_1_l_2);
nor I_13(n23_2,n24_2,n31_2);
nand I_14(n24_2,IN_1_4_l_2,IN_2_4_l_2);
nand I_15(n25_2,n26_2,n27_2);
nor I_16(n26_2,IN_1_3_l_2,n30_2);
not I_17(n27_2,n_429_or_0_5_r_2);
nor I_18(n28_2,n22_2,n23_2);
nand I_19(n29_2,N1508_0_r_2,n26_2);
or I_20(n30_2,IN_2_3_l_2,IN_3_3_l_2);
nor I_21(n31_2,IN_5_4_l_2,n32_2);
and I_22(n32_2,IN_3_4_l_2,IN_4_4_l_2);
nor I_23(N6147_3_r_1,n26_1,n27_1);
not I_24(N1372_4_r_1,n34_1);
nor I_25(N1508_4_r_1,n30_1,n34_1);
nor I_26(n_42_8_r_1,n23_1,n24_1);
DFFARX1 I_27(N3_8_r_1,blif_clk_net_8_r_1,n7_1,G199_8_r_1,);
nor I_28(N6147_9_r_1,n22_1,n25_1);
nor I_29(N6134_9_r_1,n29_1,n30_1);
not I_30(I_BUFF_1_9_r_1,n32_1);
not I_31(N1372_10_r_1,n36_1);
nor I_32(N1508_10_r_1,n35_1,n36_1);
and I_33(N3_8_l_1,n33_1,N1371_0_r_2);
not I_34(n7_1,blif_reset_net_8_r_1);
DFFARX1 I_35(N3_8_l_1,blif_clk_net_8_r_1,n7_1,n38_1,);
not I_36(n22_1,n38_1);
nor I_37(N3_8_r_1,n31_1,n32_1);
nor I_38(n23_1,n28_1,N6147_3_r_2);
nor I_39(n24_1,n_576_5_r_2,n_547_5_r_2);
nor I_40(n25_1,n23_1,n26_1);
not I_41(n26_1,n30_1);
nand I_42(n27_1,n22_1,n28_1);
nand I_43(n28_1,N1508_10_r_2,n_576_5_r_2);
not I_44(n29_1,n28_1);
nand I_45(n30_1,N1372_10_r_2,N6147_3_r_2);
and I_46(n31_1,n38_1,n24_1);
nand I_47(n32_1,n26_1,n37_1);
nand I_48(n33_1,G78_5_r_2,n_547_5_r_2);
nand I_49(n34_1,n24_1,n29_1);
nor I_50(n35_1,n38_1,n24_1);
nand I_51(n36_1,I_BUFF_1_9_r_1,n23_1);
or I_52(n37_1,N1371_0_r_2,G78_5_r_2);
endmodule


