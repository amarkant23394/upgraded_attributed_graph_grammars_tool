module test_I16145(I1477,I1470,I14278,I16145);
input I1477,I1470,I14278;
output I16145;
wire I13752,I16052,I13775,I15611,I16069;
DFFARX1 I_0(I14278,I1470,I13775,,,I13752,);
not I_1(I16145,I16069);
DFFARX1 I_2(I13752,I1470,I15611,,,I16052,);
not I_3(I13775,I1477);
not I_4(I15611,I1477);
not I_5(I16069,I16052);
endmodule


