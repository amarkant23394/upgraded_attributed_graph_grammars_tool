module test_I15645(I12270,I1477,I1470,I13809,I11959,I15645);
input I12270,I1477,I1470,I13809,I11959;
output I15645;
wire I13826,I13761,I12239,I13860,I14162,I11938,I13891,I13775,I13740,I13843,I12075,I11965,I11944;
DFFARX1 I_0(I13809,I1470,I13775,,,I13826,);
nand I_1(I13761,I13891,I13860);
nor I_2(I15645,I13761,I13740);
DFFARX1 I_3(I1470,,,I12239,);
nor I_4(I13860,I13843,I13826);
DFFARX1 I_5(I11938,I1470,I13775,,,I14162,);
and I_6(I11938,I12270,I12239);
DFFARX1 I_7(I11944,I1470,I13775,,,I13891,);
not I_8(I13775,I1477);
DFFARX1 I_9(I14162,I1470,I13775,,,I13740,);
nor I_10(I13843,I11959,I11965);
DFFARX1 I_11(I1470,,,I12075,);
DFFARX1 I_12(I1470,,,I11965,);
not I_13(I11944,I12075);
endmodule


