module test_final(IN_1_2_l,IN_2_2_l,IN_3_2_l,IN_4_2_l,IN_5_2_l,IN_1_4_l,IN_2_4_l,IN_3_4_l,IN_4_4_l,IN_5_4_l,IN_1_9_l,IN_2_9_l,IN_3_9_l,IN_4_9_l,IN_5_9_l,blif_clk_net_8_r,blif_reset_net_8_r,N1371_0_r,N1508_0_r,N6147_2_r,N6147_3_r,N1372_4_r,N1508_4_r,N1507_6_r,N1508_6_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r);
input IN_1_2_l,IN_2_2_l,IN_3_2_l,IN_4_2_l,IN_5_2_l,IN_1_4_l,IN_2_4_l,IN_3_4_l,IN_4_4_l,IN_5_4_l,IN_1_9_l,IN_2_9_l,IN_3_9_l,IN_4_9_l,IN_5_9_l,blif_clk_net_8_r,blif_reset_net_8_r;
output N1371_0_r,N1508_0_r,N6147_2_r,N6147_3_r,N1372_4_r,N1508_4_r,N1507_6_r,N1508_6_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r;
wire N6147_2_l,n5_2_l,n6_2_l,N6138_2_l,n7_2_l,N1372_4_l,N1508_4_l,n6_4_l,n7_4_l,n8_4_l,N6150_9_l,N6147_9_l,N6134_9_l,n3_9_l,I_BUFF_1_9_l,n3_0_r,n4_0_r,n5_2_r,n6_2_r,N6138_2_r,n7_2_r,n3_3_r,N6138_3_r,n6_4_r,n7_4_r,n8_4_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,N3_8_r,n1_8_r,n3_8_r,N6150_9_r,n3_9_r;
nor I_0(N6147_2_l,n5_2_l,n6_2_l);
nor I_1(n5_2_l,IN_5_2_l,n7_2_l);
not I_2(n6_2_l,N6138_2_l);
nor I_3(N6138_2_l,IN_1_2_l,IN_2_2_l);
nor I_4(n7_2_l,IN_3_2_l,IN_4_2_l);
not I_5(N1372_4_l,n7_4_l);
nor I_6(N1508_4_l,n6_4_l,n7_4_l);
nor I_7(n6_4_l,IN_5_4_l,n8_4_l);
nand I_8(n7_4_l,IN_1_4_l,IN_2_4_l);
and I_9(n8_4_l,IN_3_4_l,IN_4_4_l);
not I_10(N6150_9_l,IN_2_9_l);
nor I_11(N6147_9_l,N6150_9_l,n3_9_l);
nor I_12(N6134_9_l,IN_5_9_l,n3_9_l);
nor I_13(n3_9_l,IN_3_9_l,IN_4_9_l);
buf I_14(I_BUFF_1_9_l,IN_1_9_l);
nor I_15(N1371_0_r,n4_0_r,N6134_9_l);
nor I_16(N1508_0_r,n3_0_r,n4_0_r);
nor I_17(n3_0_r,N1372_4_l,N1508_4_l);
not I_18(n4_0_r,N6147_9_l);
nor I_19(N6147_2_r,n5_2_r,n6_2_r);
nor I_20(n5_2_r,n7_2_r,I_BUFF_1_9_l);
not I_21(n6_2_r,N6138_2_r);
nor I_22(N6138_2_r,N1508_4_l,N6147_9_l);
nor I_23(n7_2_r,N6147_9_l,N6147_2_l);
nor I_24(N6147_3_r,n3_3_r,N6147_2_l);
not I_25(n3_3_r,N6138_3_r);
nor I_26(N6138_3_r,I_BUFF_1_9_l,N6147_2_l);
not I_27(N1372_4_r,n7_4_r);
nor I_28(N1508_4_r,n6_4_r,n7_4_r);
nor I_29(n6_4_r,n8_4_r,N6147_9_l);
nand I_30(n7_4_r,N6134_9_l,N6147_2_l);
and I_31(n8_4_r,I_BUFF_1_9_l,N1508_4_l);
nor I_32(N1507_6_r,n8_6_r,n9_6_r);
and I_33(N1508_6_r,n6_6_r,I_BUFF_1_9_l);
nor I_34(n6_6_r,n7_6_r,n8_6_r);
not I_35(n7_6_r,N6147_9_l);
nor I_36(n8_6_r,n9_6_r,N6147_2_l);
and I_37(n9_6_r,N1508_4_l,N6134_9_l);
nor I_38(n_42_8_r,N6147_2_l,N6134_9_l);
DFFARX1 I_39(N3_8_r,blif_clk_net_8_r,n1_8_r,G199_8_r,);
and I_40(N3_8_r,n3_8_r,N6134_9_l);
not I_41(n1_8_r,blif_reset_net_8_r);
nand I_42(n3_8_r,N6134_9_l,N1372_4_l);
not I_43(N6150_9_r,I_BUFF_1_9_l);
nor I_44(N6147_9_r,N6150_9_r,n3_9_r);
nor I_45(N6134_9_r,n3_9_r,N1372_4_l);
nor I_46(n3_9_r,N1508_4_l,N1372_4_l);
buf I_47(I_BUFF_1_9_r,N1372_4_l);
endmodule


