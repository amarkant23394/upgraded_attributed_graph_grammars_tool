module test_I10020(I1477,I10185,I7535,I1470,I10020);
input I1477,I10185,I7535,I1470;
output I10020;
wire I7538,I10219,I10154,I10137,I7541,I7553,I10052,I10202,I10287,I10120;
DFFARX1 I_0(I1470,,,I7538,);
DFFARX1 I_1(I10202,I1470,I10052,,,I10219,);
nand I_2(I10154,I10137,I10120);
DFFARX1 I_3(I10287,I1470,I10052,,,I10020,);
DFFARX1 I_4(I7553,I1470,I10052,,,I10137,);
DFFARX1 I_5(I1470,,,I7541,);
DFFARX1 I_6(I1470,,,I7553,);
not I_7(I10052,I1477);
and I_8(I10202,I10185,I7541);
and I_9(I10287,I10219,I10154);
nor I_10(I10120,I7538,I7535);
endmodule


