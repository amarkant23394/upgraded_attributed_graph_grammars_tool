module Benchmark_testing100000(I1345,I1353,I1361,I1369,I1377,I1385,I1393,I1401,I1409,I1417,I1425,I1433,I1441,I1449,I1457,I1465,I1473,I1481,I1489,I1497,I1505,I1513,I1521,I1529,I1537,I1545,I1553,I1561,I1569,I1577,I1585,I1593,I1601,I1609,I1617,I1625,I1633,I1641,I1649,I1657,I1665,I1673,I1681,I1689,I1697,I1705,I1713,I1721,I1729,I1737,I1745,I1753,I1761,I1769,I1777,I1785,I1793,I1801,I1809,I1817,I1825,I1833,I1841,I1849,I1857,I1865,I1873,I1881,I1889,I1897,I1905,I1913,I1921,I1929,I1937,I1945,I1953,I1961,I1969,I1977,I1985,I1993,I2001,I2009,I2017,I2025,I2033,I2041,I2049,I2057,I2065,I2073,I2081,I2089,I2097,I2105,I2113,I2121,I2129,I2137,I2145,I2153,I2161,I2169,I2177,I2185,I2193,I2201,I2209,I2217,I2224,I2231,I21929,I21932,I21935,I21938,I21941,I21944,I21947,I21950,I41615,I41618,I41621,I41624,I41627,I41630,I41633,I41636,I61370,I61373,I61376,I61379,I61382,I61385,I61388,I61391,I61394,I61397,I81101,I81104,I81107,I81110,I81113,I81116,I81119,I81122,I81125,I100778,I100781,I100784,I100787,I100790,I100793,I100796,I100799,I120494,I120497,I120500,I120503,I120506,I120509,I120512,I120515,I120518,I120521,I140168,I140171,I140174,I140177,I140180,I140183,I140186,I140189,I140192,I159869,I159872,I159875,I159878,I159881,I159884,I159887,I159890,I159893,I159896,I179561,I179564,I179567,I179570,I179573,I179576,I179579,I179582,I179585,I199241,I199244,I199247,I199250,I199253,I199256,I199259,I199262,I199265,I199268);
input I1345,I1353,I1361,I1369,I1377,I1385,I1393,I1401,I1409,I1417,I1425,I1433,I1441,I1449,I1457,I1465,I1473,I1481,I1489,I1497,I1505,I1513,I1521,I1529,I1537,I1545,I1553,I1561,I1569,I1577,I1585,I1593,I1601,I1609,I1617,I1625,I1633,I1641,I1649,I1657,I1665,I1673,I1681,I1689,I1697,I1705,I1713,I1721,I1729,I1737,I1745,I1753,I1761,I1769,I1777,I1785,I1793,I1801,I1809,I1817,I1825,I1833,I1841,I1849,I1857,I1865,I1873,I1881,I1889,I1897,I1905,I1913,I1921,I1929,I1937,I1945,I1953,I1961,I1969,I1977,I1985,I1993,I2001,I2009,I2017,I2025,I2033,I2041,I2049,I2057,I2065,I2073,I2081,I2089,I2097,I2105,I2113,I2121,I2129,I2137,I2145,I2153,I2161,I2169,I2177,I2185,I2193,I2201,I2209,I2217,I2224,I2231;
output I21929,I21932,I21935,I21938,I21941,I21944,I21947,I21950,I41615,I41618,I41621,I41624,I41627,I41630,I41633,I41636,I61370,I61373,I61376,I61379,I61382,I61385,I61388,I61391,I61394,I61397,I81101,I81104,I81107,I81110,I81113,I81116,I81119,I81122,I81125,I100778,I100781,I100784,I100787,I100790,I100793,I100796,I100799,I120494,I120497,I120500,I120503,I120506,I120509,I120512,I120515,I120518,I120521,I140168,I140171,I140174,I140177,I140180,I140183,I140186,I140189,I140192,I159869,I159872,I159875,I159878,I159881,I159884,I159887,I159890,I159893,I159896,I179561,I179564,I179567,I179570,I179573,I179576,I179579,I179582,I179585,I199241,I199244,I199247,I199250,I199253,I199256,I199259,I199262,I199265,I199268;
wire I1345,I1353,I1361,I1369,I1377,I1385,I1393,I1401,I1409,I1417,I1425,I1433,I1441,I1449,I1457,I1465,I1473,I1481,I1489,I1497,I1505,I1513,I1521,I1529,I1537,I1545,I1553,I1561,I1569,I1577,I1585,I1593,I1601,I1609,I1617,I1625,I1633,I1641,I1649,I1657,I1665,I1673,I1681,I1689,I1697,I1705,I1713,I1721,I1729,I1737,I1745,I1753,I1761,I1769,I1777,I1785,I1793,I1801,I1809,I1817,I1825,I1833,I1841,I1849,I1857,I1865,I1873,I1881,I1889,I1897,I1905,I1913,I1921,I1929,I1937,I1945,I1953,I1961,I1969,I1977,I1985,I1993,I2001,I2009,I2017,I2025,I2033,I2041,I2049,I2057,I2065,I2073,I2081,I2089,I2097,I2105,I2113,I2121,I2129,I2137,I2145,I2153,I2161,I2169,I2177,I2185,I2193,I2201,I2209,I2217,I2224,I2231,I2271,I2274,I2277,I2280,I2283,I2286,I2289,I2292,I2295,I2341,I2344,I2347,I2350,I2353,I2356,I2359,I2362,I2365,I2411,I2414,I2417,I2420,I2423,I2426,I2429,I2432,I2435,I2438,I2484,I2487,I2490,I2493,I2496,I2499,I2502,I2505,I2508,I2554,I2557,I2560,I2563,I2566,I2569,I2572,I2575,I2578,I2624,I2627,I2630,I2633,I2636,I2639,I2642,I2645,I2648,I2694,I2697,I2700,I2703,I2706,I2709,I2712,I2715,I2761,I2764,I2767,I2770,I2773,I2776,I2779,I2782,I2785,I2788,I2834,I2837,I2840,I2843,I2846,I2849,I2852,I2855,I2858,I2904,I2907,I2910,I2913,I2916,I2919,I2922,I2925,I2928,I2931,I2977,I2980,I2983,I2986,I2989,I2992,I2995,I2998,I3001,I3047,I3050,I3053,I3056,I3059,I3062,I3065,I3068,I3114,I3117,I3120,I3123,I3126,I3129,I3132,I3135,I3138,I3184,I3187,I3190,I3193,I3196,I3199,I3202,I3205,I3208,I3211,I3257,I3260,I3263,I3266,I3269,I3272,I3275,I3278,I3281,I3327,I3330,I3333,I3336,I3339,I3342,I3345,I3348,I3351,I3354,I3400,I3403,I3406,I3409,I3412,I3415,I3418,I3421,I3424,I3470,I3473,I3476,I3479,I3482,I3485,I3488,I3491,I3494,I3497,I3543,I3546,I3549,I3552,I3555,I3558,I3561,I3564,I3567,I3613,I3616,I3619,I3622,I3625,I3628,I3631,I3634,I3637,I3640,I3686,I3689,I3692,I3695,I3698,I3701,I3704,I3707,I3710,I3713,I3759,I3762,I3765,I3768,I3771,I3774,I3777,I3780,I3783,I3829,I3832,I3835,I3838,I3841,I3844,I3847,I3850,I3853,I3856,I3902,I3905,I3908,I3911,I3914,I3917,I3920,I3923,I3926,I3972,I3975,I3978,I3981,I3984,I3987,I3990,I3993,I3996,I3999,I4045,I4048,I4051,I4054,I4057,I4060,I4063,I4066,I4069,I4072,I4118,I4121,I4124,I4127,I4130,I4133,I4136,I4139,I4142,I4145,I4191,I4194,I4197,I4200,I4203,I4206,I4209,I4212,I4215,I4218,I4264,I4267,I4270,I4273,I4276,I4279,I4282,I4285,I4288,I4334,I4337,I4340,I4343,I4346,I4349,I4352,I4355,I4358,I4361,I4407,I4410,I4413,I4416,I4419,I4422,I4425,I4428,I4431,I4434,I4480,I4483,I4486,I4489,I4492,I4495,I4498,I4501,I4547,I4550,I4553,I4556,I4559,I4562,I4565,I4568,I4571,I4617,I4620,I4623,I4626,I4629,I4632,I4635,I4638,I4684,I4687,I4690,I4693,I4696,I4699,I4702,I4705,I4708,I4754,I4757,I4760,I4763,I4766,I4769,I4772,I4775,I4821,I4824,I4827,I4830,I4833,I4836,I4839,I4842,I4845,I4891,I4894,I4897,I4900,I4903,I4906,I4909,I4912,I4958,I4961,I4964,I4967,I4970,I4973,I4976,I4979,I4982,I5028,I5031,I5034,I5037,I5040,I5043,I5046,I5049,I5052,I5055,I5101,I5104,I5107,I5110,I5113,I5116,I5119,I5122,I5168,I5171,I5174,I5177,I5180,I5183,I5186,I5189,I5192,I5195,I5241,I5244,I5247,I5250,I5253,I5256,I5259,I5262,I5265,I5268,I5314,I5317,I5320,I5323,I5326,I5329,I5332,I5335,I5338,I5341,I5387,I5390,I5393,I5396,I5399,I5402,I5405,I5408,I5411,I5457,I5460,I5463,I5466,I5469,I5472,I5475,I5478,I5481,I5484,I5530,I5533,I5536,I5539,I5542,I5545,I5548,I5551,I5554,I5600,I5603,I5606,I5609,I5612,I5615,I5618,I5621,I5624,I5627,I5673,I5676,I5679,I5682,I5685,I5688,I5691,I5694,I5740,I5743,I5746,I5749,I5752,I5755,I5758,I5761,I5764,I5767,I5813,I5816,I5819,I5822,I5825,I5828,I5831,I5834,I5837,I5883,I5886,I5889,I5892,I5895,I5898,I5901,I5904,I5907,I5953,I5956,I5959,I5962,I5965,I5968,I5971,I5974,I5977,I6023,I6026,I6029,I6032,I6035,I6038,I6041,I6044,I6047,I6093,I6096,I6099,I6102,I6105,I6108,I6111,I6114,I6160,I6163,I6166,I6169,I6172,I6175,I6178,I6181,I6227,I6230,I6233,I6236,I6239,I6242,I6245,I6248,I6251,I6297,I6300,I6303,I6306,I6309,I6312,I6315,I6318,I6321,I6367,I6370,I6373,I6376,I6379,I6382,I6385,I6388,I6391,I6437,I6440,I6443,I6446,I6449,I6452,I6455,I6458,I6461,I6507,I6510,I6513,I6516,I6519,I6522,I6525,I6528,I6531,I6577,I6580,I6583,I6586,I6589,I6592,I6595,I6598,I6601,I6647,I6650,I6653,I6656,I6659,I6662,I6665,I6668,I6671,I6717,I6720,I6723,I6726,I6729,I6732,I6735,I6738,I6741,I6744,I6790,I6793,I6796,I6799,I6802,I6805,I6808,I6811,I6857,I6860,I6863,I6866,I6869,I6872,I6875,I6878,I6881,I6884,I6930,I6933,I6936,I6939,I6942,I6945,I6948,I6951,I6954,I7000,I7003,I7006,I7009,I7012,I7015,I7018,I7021,I7024,I7027,I7073,I7076,I7079,I7082,I7085,I7088,I7091,I7094,I7140,I7143,I7146,I7149,I7152,I7155,I7158,I7161,I7164,I7210,I7213,I7216,I7219,I7222,I7225,I7228,I7231,I7234,I7280,I7283,I7286,I7289,I7292,I7295,I7298,I7301,I7304,I7350,I7353,I7356,I7359,I7362,I7365,I7368,I7371,I7374,I7420,I7423,I7426,I7429,I7432,I7435,I7438,I7441,I7444,I7490,I7493,I7496,I7499,I7502,I7505,I7508,I7511,I7514,I7517,I7563,I7566,I7569,I7572,I7575,I7578,I7581,I7584,I7587,I7633,I7636,I7639,I7642,I7645,I7648,I7651,I7654,I7700,I7703,I7706,I7709,I7712,I7715,I7718,I7721,I7724,I7770,I7773,I7776,I7779,I7782,I7785,I7788,I7791,I7794,I7840,I7843,I7846,I7849,I7852,I7855,I7858,I7861,I7864,I7867,I7913,I7916,I7919,I7922,I7925,I7928,I7931,I7934,I7937,I7940,I7986,I7989,I7992,I7995,I7998,I8001,I8004,I8007,I8010,I8013,I8059,I8062,I8065,I8068,I8071,I8074,I8077,I8080,I8083,I8129,I8132,I8135,I8138,I8141,I8144,I8147,I8150,I8153,I8156,I8202,I8205,I8208,I8211,I8214,I8217,I8220,I8223,I8226,I8272,I8275,I8278,I8281,I8284,I8287,I8290,I8293,I8296,I8342,I8345,I8348,I8351,I8354,I8357,I8360,I8363,I8366,I8412,I8415,I8418,I8421,I8424,I8427,I8430,I8433,I8436,I8439,I8485,I8488,I8491,I8494,I8497,I8500,I8503,I8506,I8509,I8555,I8558,I8561,I8564,I8567,I8570,I8573,I8576,I8579,I8582,I8628,I8631,I8634,I8637,I8640,I8643,I8646,I8649,I8652,I8655,I8701,I8704,I8707,I8710,I8713,I8716,I8719,I8722,I8725,I8771,I8774,I8777,I8780,I8783,I8786,I8789,I8792,I8795,I8841,I8844,I8847,I8850,I8853,I8856,I8859,I8862,I8865,I8868,I8914,I8917,I8920,I8923,I8926,I8929,I8932,I8935,I8938,I8941,I8987,I8990,I8993,I8996,I8999,I9002,I9005,I9008,I9011,I9014,I9060,I9063,I9066,I9069,I9072,I9075,I9078,I9081,I9084,I9130,I9133,I9136,I9139,I9142,I9145,I9148,I9151,I9154,I9200,I9203,I9206,I9209,I9212,I9215,I9218,I9221,I9267,I9270,I9273,I9276,I9279,I9282,I9285,I9288,I9291,I9294,I9340,I9343,I9346,I9349,I9352,I9355,I9358,I9361,I9364,I9410,I9413,I9416,I9419,I9422,I9425,I9428,I9431,I9434,I9480,I9483,I9486,I9489,I9492,I9495,I9498,I9501,I9504,I9507,I9553,I9556,I9559,I9562,I9565,I9568,I9571,I9574,I9577,I9623,I9626,I9629,I9632,I9635,I9638,I9641,I9644,I9647,I9693,I9696,I9699,I9702,I9705,I9708,I9711,I9714,I9717,I9763,I9766,I9769,I9772,I9775,I9778,I9781,I9784,I9787,I9833,I9836,I9839,I9842,I9845,I9848,I9851,I9854,I9857,I9903,I9906,I9909,I9912,I9915,I9918,I9921,I9924,I9927,I9973,I9976,I9979,I9982,I9985,I9988,I9991,I9994,I9997,I10043,I10046,I10049,I10052,I10055,I10058,I10061,I10064,I10067,I10070,I10116,I10119,I10122,I10125,I10128,I10131,I10134,I10137,I10140,I10186,I10189,I10192,I10195,I10198,I10201,I10204,I10207,I10210,I10213,I10259,I10262,I10265,I10268,I10271,I10274,I10277,I10280,I10283,I10329,I10332,I10335,I10338,I10341,I10344,I10347,I10350,I10353,I10399,I10402,I10405,I10408,I10411,I10414,I10417,I10420,I10423,I10469,I10472,I10475,I10478,I10481,I10484,I10487,I10490,I10493,I10539,I10542,I10545,I10548,I10551,I10554,I10557,I10560,I10606,I10609,I10612,I10615,I10618,I10621,I10624,I10627,I10630,I10633,I10679,I10682,I10685,I10688,I10691,I10694,I10697,I10700,I10703,I10749,I10752,I10755,I10758,I10761,I10764,I10767,I10770,I10773,I10776,I10822,I10825,I10828,I10831,I10834,I10837,I10840,I10843,I10846,I10849,I10895,I10898,I10901,I10904,I10907,I10910,I10913,I10916,I10919,I10965,I10968,I10971,I10974,I10977,I10980,I10983,I10986,I10989,I11035,I11038,I11041,I11044,I11047,I11050,I11053,I11056,I11059,I11062,I11108,I11111,I11114,I11117,I11120,I11123,I11126,I11129,I11132,I11178,I11181,I11184,I11187,I11190,I11193,I11196,I11199,I11202,I11205,I11251,I11254,I11257,I11260,I11263,I11266,I11269,I11272,I11275,I11278,I11324,I11327,I11330,I11333,I11336,I11339,I11342,I11345,I11348,I11351,I11397,I11400,I11403,I11406,I11409,I11412,I11415,I11418,I11421,I11467,I11470,I11473,I11476,I11479,I11482,I11485,I11488,I11534,I11537,I11540,I11543,I11546,I11549,I11552,I11555,I11558,I11604,I11607,I11610,I11613,I11616,I11619,I11622,I11625,I11671,I11674,I11677,I11680,I11683,I11686,I11689,I11692,I11695,I11741,I11744,I11747,I11750,I11753,I11756,I11759,I11762,I11765,I11768,I11814,I11817,I11820,I11823,I11826,I11829,I11832,I11835,I11838,I11884,I11887,I11890,I11893,I11896,I11899,I11902,I11905,I11908,I11954,I11957,I11960,I11963,I11966,I11969,I11972,I11975,I11978,I11981,I12027,I12030,I12033,I12036,I12039,I12042,I12045,I12048,I12051,I12054,I12100,I12103,I12106,I12109,I12112,I12115,I12118,I12121,I12124,I12170,I12173,I12176,I12179,I12182,I12185,I12188,I12191,I12194,I12240,I12243,I12246,I12249,I12252,I12255,I12258,I12261,I12264,I12310,I12313,I12316,I12319,I12322,I12325,I12328,I12331,I12334,I12337,I12383,I12386,I12389,I12392,I12395,I12398,I12401,I12404,I12407,I12410,I12456,I12459,I12462,I12465,I12468,I12471,I12474,I12477,I12480,I12526,I12529,I12532,I12535,I12538,I12541,I12544,I12547,I12550,I12596,I12599,I12602,I12605,I12608,I12611,I12614,I12617,I12620,I12623,I12669,I12672,I12675,I12678,I12681,I12684,I12687,I12690,I12693,I12696,I12742,I12745,I12748,I12751,I12754,I12757,I12760,I12763,I12766,I12769,I12815,I12818,I12821,I12824,I12827,I12830,I12833,I12836,I12839,I12885,I12888,I12891,I12894,I12897,I12900,I12903,I12906,I12909,I12912,I12958,I12961,I12964,I12967,I12970,I12973,I12976,I12979,I12982,I13028,I13031,I13034,I13037,I13040,I13043,I13046,I13049,I13095,I13098,I13101,I13104,I13107,I13110,I13113,I13116,I13119,I13165,I13168,I13171,I13174,I13177,I13180,I13183,I13186,I13189,I13192,I13238,I13241,I13244,I13247,I13250,I13253,I13256,I13259,I13262,I13308,I13311,I13314,I13317,I13320,I13323,I13326,I13329,I13375,I13378,I13381,I13384,I13387,I13390,I13393,I13396,I13399,I13445,I13448,I13451,I13454,I13457,I13460,I13463,I13466,I13469,I13472,I13518,I13521,I13524,I13527,I13530,I13533,I13536,I13539,I13542,I13588,I13591,I13594,I13597,I13600,I13603,I13606,I13609,I13655,I13658,I13661,I13664,I13667,I13670,I13673,I13676,I13679,I13725,I13728,I13731,I13734,I13737,I13740,I13743,I13746,I13749,I13752,I13798,I13801,I13804,I13807,I13810,I13813,I13816,I13819,I13822,I13868,I13871,I13874,I13877,I13880,I13883,I13886,I13889,I13892,I13895,I13941,I13944,I13947,I13950,I13953,I13956,I13959,I13962,I13965,I14011,I14014,I14017,I14020,I14023,I14026,I14029,I14032,I14035,I14038,I14084,I14087,I14090,I14093,I14096,I14099,I14102,I14105,I14151,I14154,I14157,I14160,I14163,I14166,I14169,I14172,I14175,I14178,I14224,I14227,I14230,I14233,I14236,I14239,I14242,I14245,I14248,I14294,I14297,I14300,I14303,I14306,I14309,I14312,I14315,I14318,I14364,I14367,I14370,I14373,I14376,I14379,I14382,I14385,I14388,I14391,I14437,I14440,I14443,I14446,I14449,I14452,I14455,I14458,I14504,I14507,I14510,I14513,I14516,I14519,I14522,I14525,I14528,I14531,I14577,I14580,I14583,I14586,I14589,I14592,I14595,I14598,I14601,I14604,I14650,I14653,I14656,I14659,I14662,I14665,I14668,I14671,I14674,I14720,I14723,I14726,I14729,I14732,I14735,I14738,I14741,I14744,I14790,I14793,I14796,I14799,I14802,I14805,I14808,I14811,I14814,I14860,I14863,I14866,I14869,I14872,I14875,I14878,I14881,I14927,I14930,I14933,I14936,I14939,I14942,I14945,I14948,I14951,I14997,I15000,I15003,I15006,I15009,I15012,I15015,I15018,I15021,I15024,I15070,I15073,I15076,I15079,I15082,I15085,I15088,I15091,I15094,I15097,I15143,I15146,I15149,I15152,I15155,I15158,I15161,I15164,I15167,I15213,I15216,I15219,I15222,I15225,I15228,I15231,I15234,I15237,I15283,I15286,I15289,I15292,I15295,I15298,I15301,I15304,I15307,I15310,I15356,I15359,I15362,I15365,I15368,I15371,I15374,I15377,I15380,I15426,I15429,I15432,I15435,I15438,I15441,I15444,I15447,I15450,I15496,I15499,I15502,I15505,I15508,I15511,I15514,I15517,I15520,I15523,I15569,I15572,I15575,I15578,I15581,I15584,I15587,I15590,I15593,I15639,I15642,I15645,I15648,I15651,I15654,I15657,I15660,I15663,I15666,I15712,I15715,I15718,I15721,I15724,I15727,I15730,I15733,I15736,I15782,I15785,I15788,I15791,I15794,I15797,I15800,I15803,I15849,I15852,I15855,I15858,I15861,I15864,I15867,I15870,I15873,I15876,I15922,I15925,I15928,I15931,I15934,I15937,I15940,I15943,I15946,I15949,I15995,I15998,I16001,I16004,I16007,I16010,I16013,I16016,I16019,I16065,I16068,I16071,I16074,I16077,I16080,I16083,I16086,I16089,I16135,I16138,I16141,I16144,I16147,I16150,I16153,I16156,I16202,I16205,I16208,I16211,I16214,I16217,I16220,I16223,I16226,I16229,I16275,I16278,I16281,I16284,I16287,I16290,I16293,I16296,I16299,I16345,I16348,I16351,I16354,I16357,I16360,I16363,I16366,I16369,I16372,I16418,I16421,I16424,I16427,I16430,I16433,I16436,I16439,I16485,I16488,I16491,I16494,I16497,I16500,I16503,I16506,I16509,I16512,I16558,I16561,I16564,I16567,I16570,I16573,I16576,I16579,I16582,I16628,I16631,I16634,I16637,I16640,I16643,I16646,I16649,I16652,I16655,I16701,I16704,I16707,I16710,I16713,I16716,I16719,I16722,I16725,I16728,I16774,I16777,I16780,I16783,I16786,I16789,I16792,I16795,I16798,I16844,I16847,I16850,I16853,I16856,I16859,I16862,I16865,I16868,I16914,I16917,I16920,I16923,I16926,I16929,I16932,I16935,I16981,I16984,I16987,I16990,I16993,I16996,I16999,I17002,I17005,I17008,I17054,I17057,I17060,I17063,I17066,I17069,I17072,I17075,I17078,I17124,I17127,I17130,I17133,I17136,I17139,I17142,I17145,I17148,I17194,I17197,I17200,I17203,I17206,I17209,I17212,I17215,I17218,I17264,I17267,I17270,I17273,I17276,I17279,I17282,I17285,I17288,I17291,I17337,I17340,I17343,I17346,I17349,I17352,I17355,I17358,I17361,I17407,I17410,I17413,I17416,I17419,I17422,I17425,I17428,I17431,I17434,I17480,I17483,I17486,I17489,I17492,I17495,I17498,I17501,I17504,I17550,I17553,I17556,I17559,I17562,I17565,I17568,I17571,I17574,I17620,I17623,I17626,I17629,I17632,I17635,I17638,I17641,I17644,I17690,I17693,I17696,I17699,I17702,I17705,I17708,I17711,I17714,I17717,I17763,I17766,I17769,I17772,I17775,I17778,I17781,I17784,I17787,I17833,I17836,I17839,I17842,I17845,I17848,I17851,I17854,I17857,I17903,I17906,I17909,I17912,I17915,I17918,I17921,I17924,I17927,I17930,I17976,I17979,I17982,I17985,I17988,I17991,I17994,I17997,I18000,I18046,I18049,I18052,I18055,I18058,I18061,I18064,I18067,I18070,I18116,I18119,I18122,I18125,I18128,I18131,I18134,I18137,I18140,I18186,I18189,I18192,I18195,I18198,I18201,I18204,I18207,I18210,I18213,I18259,I18262,I18265,I18268,I18271,I18274,I18277,I18280,I18283,I18286,I18332,I18335,I18338,I18341,I18344,I18347,I18350,I18353,I18356,I18402,I18405,I18408,I18411,I18414,I18417,I18420,I18423,I18426,I18429,I18475,I18478,I18481,I18484,I18487,I18490,I18493,I18496,I18499,I18545,I18548,I18551,I18554,I18557,I18560,I18563,I18566,I18569,I18615,I18618,I18621,I18624,I18627,I18630,I18633,I18636,I18639,I18685,I18688,I18691,I18694,I18697,I18700,I18703,I18706,I18709,I18712,I18758,I18761,I18764,I18767,I18770,I18773,I18776,I18779,I18782,I18828,I18831,I18834,I18837,I18840,I18843,I18846,I18849,I18852,I18898,I18901,I18904,I18907,I18910,I18913,I18916,I18919,I18922,I18925,I18971,I18974,I18977,I18980,I18983,I18986,I18989,I18992,I18995,I19041,I19044,I19047,I19050,I19053,I19056,I19059,I19062,I19065,I19111,I19114,I19117,I19120,I19123,I19126,I19129,I19132,I19135,I19181,I19184,I19187,I19190,I19193,I19196,I19199,I19202,I19205,I19251,I19254,I19257,I19260,I19263,I19266,I19269,I19272,I19275,I19321,I19324,I19327,I19330,I19333,I19336,I19339,I19342,I19345,I19348,I19394,I19397,I19400,I19403,I19406,I19409,I19412,I19415,I19418,I19421,I19467,I19470,I19473,I19476,I19479,I19482,I19485,I19488,I19491,I19494,I19540,I19543,I19546,I19549,I19552,I19555,I19558,I19561,I19607,I19610,I19613,I19616,I19619,I19622,I19625,I19628,I19631,I19677,I19680,I19683,I19686,I19689,I19692,I19695,I19698,I19701,I19704,I19750,I19753,I19756,I19759,I19762,I19765,I19768,I19771,I19774,I19820,I19823,I19826,I19829,I19832,I19835,I19838,I19841,I19844,I19890,I19893,I19896,I19899,I19902,I19905,I19908,I19911,I19914,I19960,I19963,I19966,I19969,I19972,I19975,I19978,I19981,I20027,I20030,I20033,I20036,I20039,I20042,I20045,I20048,I20051,I20097,I20100,I20103,I20106,I20109,I20112,I20115,I20118,I20121,I20124,I20170,I20173,I20176,I20179,I20182,I20185,I20188,I20191,I20194,I20240,I20243,I20246,I20249,I20252,I20255,I20258,I20261,I20264,I20310,I20313,I20316,I20319,I20322,I20325,I20328,I20331,I20334,I20380,I20383,I20386,I20389,I20392,I20395,I20398,I20401,I20404,I20450,I20453,I20456,I20459,I20462,I20465,I20468,I20471,I20474,I20477,I20523,I20526,I20529,I20532,I20535,I20538,I20541,I20544,I20547,I20593,I20596,I20599,I20602,I20605,I20608,I20611,I20614,I20617,I20663,I20666,I20669,I20672,I20675,I20678,I20681,I20684,I20687,I20733,I20736,I20739,I20742,I20745,I20748,I20751,I20754,I20757,I20760,I20806,I20809,I20812,I20815,I20818,I20821,I20824,I20827,I20830,I20833,I20879,I20882,I20885,I20888,I20891,I20894,I20897,I20900,I20903,I20949,I20952,I20955,I20958,I20961,I20964,I20967,I20970,I20973,I21019,I21022,I21025,I21028,I21031,I21034,I21037,I21040,I21086,I21089,I21092,I21095,I21098,I21101,I21104,I21107,I21110,I21156,I21159,I21162,I21165,I21168,I21171,I21174,I21177,I21180,I21226,I21229,I21232,I21235,I21238,I21241,I21244,I21247,I21250,I21253,I21299,I21302,I21305,I21308,I21311,I21314,I21317,I21320,I21323,I21369,I21372,I21375,I21378,I21381,I21384,I21387,I21390,I21393,I21439,I21442,I21445,I21448,I21451,I21454,I21457,I21460,I21463,I21509,I21512,I21515,I21518,I21521,I21524,I21527,I21530,I21533,I21579,I21582,I21585,I21588,I21591,I21594,I21597,I21600,I21603,I21649,I21652,I21655,I21658,I21661,I21664,I21667,I21670,I21673,I21719,I21722,I21725,I21728,I21731,I21734,I21737,I21740,I21743,I21746,I21792,I21795,I21798,I21801,I21804,I21807,I21810,I21813,I21859,I21862,I21865,I21868,I21871,I21874,I21877,I21880,I21883,I21996,I21999,I22002,I22005,I22008,I22011,I22014,I22017,I22020,I22066,I22069,I22072,I22075,I22078,I22081,I22084,I22087,I22090,I22093,I22139,I22142,I22145,I22148,I22151,I22154,I22157,I22160,I22163,I22209,I22212,I22215,I22218,I22221,I22224,I22227,I22230,I22233,I22279,I22282,I22285,I22288,I22291,I22294,I22297,I22300,I22303,I22306,I22352,I22355,I22358,I22361,I22364,I22367,I22370,I22373,I22376,I22379,I22425,I22428,I22431,I22434,I22437,I22440,I22443,I22446,I22449,I22495,I22498,I22501,I22504,I22507,I22510,I22513,I22516,I22562,I22565,I22568,I22571,I22574,I22577,I22580,I22583,I22586,I22589,I22635,I22638,I22641,I22644,I22647,I22650,I22653,I22656,I22659,I22662,I22708,I22711,I22714,I22717,I22720,I22723,I22726,I22729,I22732,I22735,I22781,I22784,I22787,I22790,I22793,I22796,I22799,I22802,I22805,I22851,I22854,I22857,I22860,I22863,I22866,I22869,I22872,I22875,I22921,I22924,I22927,I22930,I22933,I22936,I22939,I22942,I22945,I22991,I22994,I22997,I23000,I23003,I23006,I23009,I23012,I23015,I23018,I23064,I23067,I23070,I23073,I23076,I23079,I23082,I23085,I23131,I23134,I23137,I23140,I23143,I23146,I23149,I23152,I23155,I23158,I23204,I23207,I23210,I23213,I23216,I23219,I23222,I23225,I23228,I23231,I23277,I23280,I23283,I23286,I23289,I23292,I23295,I23298,I23301,I23347,I23350,I23353,I23356,I23359,I23362,I23365,I23368,I23371,I23417,I23420,I23423,I23426,I23429,I23432,I23435,I23438,I23441,I23487,I23490,I23493,I23496,I23499,I23502,I23505,I23508,I23511,I23557,I23560,I23563,I23566,I23569,I23572,I23575,I23578,I23581,I23584,I23630,I23633,I23636,I23639,I23642,I23645,I23648,I23651,I23654,I23700,I23703,I23706,I23709,I23712,I23715,I23718,I23721,I23724,I23770,I23773,I23776,I23779,I23782,I23785,I23788,I23791,I23794,I23840,I23843,I23846,I23849,I23852,I23855,I23858,I23861,I23864,I23867,I23913,I23916,I23919,I23922,I23925,I23928,I23931,I23934,I23937,I23983,I23986,I23989,I23992,I23995,I23998,I24001,I24004,I24007,I24053,I24056,I24059,I24062,I24065,I24068,I24071,I24074,I24077,I24080,I24126,I24129,I24132,I24135,I24138,I24141,I24144,I24147,I24193,I24196,I24199,I24202,I24205,I24208,I24211,I24214,I24217,I24263,I24266,I24269,I24272,I24275,I24278,I24281,I24284,I24287,I24290,I24336,I24339,I24342,I24345,I24348,I24351,I24354,I24357,I24360,I24406,I24409,I24412,I24415,I24418,I24421,I24424,I24427,I24430,I24433,I24479,I24482,I24485,I24488,I24491,I24494,I24497,I24500,I24503,I24549,I24552,I24555,I24558,I24561,I24564,I24567,I24570,I24573,I24619,I24622,I24625,I24628,I24631,I24634,I24637,I24640,I24643,I24689,I24692,I24695,I24698,I24701,I24704,I24707,I24710,I24713,I24759,I24762,I24765,I24768,I24771,I24774,I24777,I24780,I24783,I24829,I24832,I24835,I24838,I24841,I24844,I24847,I24850,I24853,I24899,I24902,I24905,I24908,I24911,I24914,I24917,I24920,I24923,I24926,I24972,I24975,I24978,I24981,I24984,I24987,I24990,I24993,I25039,I25042,I25045,I25048,I25051,I25054,I25057,I25060,I25063,I25066,I25112,I25115,I25118,I25121,I25124,I25127,I25130,I25133,I25136,I25182,I25185,I25188,I25191,I25194,I25197,I25200,I25203,I25249,I25252,I25255,I25258,I25261,I25264,I25267,I25270,I25273,I25276,I25322,I25325,I25328,I25331,I25334,I25337,I25340,I25343,I25346,I25392,I25395,I25398,I25401,I25404,I25407,I25410,I25413,I25416,I25462,I25465,I25468,I25471,I25474,I25477,I25480,I25483,I25529,I25532,I25535,I25538,I25541,I25544,I25547,I25550,I25553,I25556,I25602,I25605,I25608,I25611,I25614,I25617,I25620,I25623,I25626,I25672,I25675,I25678,I25681,I25684,I25687,I25690,I25693,I25696,I25699,I25745,I25748,I25751,I25754,I25757,I25760,I25763,I25766,I25769,I25815,I25818,I25821,I25824,I25827,I25830,I25833,I25836,I25839,I25885,I25888,I25891,I25894,I25897,I25900,I25903,I25906,I25909,I25912,I25958,I25961,I25964,I25967,I25970,I25973,I25976,I25979,I26025,I26028,I26031,I26034,I26037,I26040,I26043,I26046,I26049,I26095,I26098,I26101,I26104,I26107,I26110,I26113,I26116,I26119,I26165,I26168,I26171,I26174,I26177,I26180,I26183,I26186,I26189,I26192,I26238,I26241,I26244,I26247,I26250,I26253,I26256,I26259,I26262,I26308,I26311,I26314,I26317,I26320,I26323,I26326,I26329,I26332,I26378,I26381,I26384,I26387,I26390,I26393,I26396,I26399,I26402,I26448,I26451,I26454,I26457,I26460,I26463,I26466,I26469,I26472,I26518,I26521,I26524,I26527,I26530,I26533,I26536,I26539,I26542,I26588,I26591,I26594,I26597,I26600,I26603,I26606,I26609,I26612,I26658,I26661,I26664,I26667,I26670,I26673,I26676,I26679,I26682,I26685,I26731,I26734,I26737,I26740,I26743,I26746,I26749,I26752,I26755,I26801,I26804,I26807,I26810,I26813,I26816,I26819,I26822,I26825,I26871,I26874,I26877,I26880,I26883,I26886,I26889,I26892,I26895,I26941,I26944,I26947,I26950,I26953,I26956,I26959,I26962,I26965,I27011,I27014,I27017,I27020,I27023,I27026,I27029,I27032,I27078,I27081,I27084,I27087,I27090,I27093,I27096,I27099,I27102,I27148,I27151,I27154,I27157,I27160,I27163,I27166,I27169,I27172,I27175,I27221,I27224,I27227,I27230,I27233,I27236,I27239,I27242,I27245,I27248,I27294,I27297,I27300,I27303,I27306,I27309,I27312,I27315,I27318,I27364,I27367,I27370,I27373,I27376,I27379,I27382,I27385,I27388,I27434,I27437,I27440,I27443,I27446,I27449,I27452,I27455,I27458,I27504,I27507,I27510,I27513,I27516,I27519,I27522,I27525,I27528,I27574,I27577,I27580,I27583,I27586,I27589,I27592,I27595,I27598,I27644,I27647,I27650,I27653,I27656,I27659,I27662,I27665,I27668,I27714,I27717,I27720,I27723,I27726,I27729,I27732,I27735,I27738,I27784,I27787,I27790,I27793,I27796,I27799,I27802,I27805,I27808,I27854,I27857,I27860,I27863,I27866,I27869,I27872,I27875,I27878,I27924,I27927,I27930,I27933,I27936,I27939,I27942,I27945,I27948,I27951,I27997,I28000,I28003,I28006,I28009,I28012,I28015,I28018,I28021,I28067,I28070,I28073,I28076,I28079,I28082,I28085,I28088,I28091,I28137,I28140,I28143,I28146,I28149,I28152,I28155,I28158,I28161,I28207,I28210,I28213,I28216,I28219,I28222,I28225,I28228,I28231,I28277,I28280,I28283,I28286,I28289,I28292,I28295,I28298,I28301,I28347,I28350,I28353,I28356,I28359,I28362,I28365,I28368,I28371,I28417,I28420,I28423,I28426,I28429,I28432,I28435,I28438,I28441,I28487,I28490,I28493,I28496,I28499,I28502,I28505,I28508,I28511,I28557,I28560,I28563,I28566,I28569,I28572,I28575,I28578,I28581,I28627,I28630,I28633,I28636,I28639,I28642,I28645,I28648,I28651,I28654,I28700,I28703,I28706,I28709,I28712,I28715,I28718,I28721,I28767,I28770,I28773,I28776,I28779,I28782,I28785,I28788,I28791,I28837,I28840,I28843,I28846,I28849,I28852,I28855,I28858,I28904,I28907,I28910,I28913,I28916,I28919,I28922,I28925,I28928,I28974,I28977,I28980,I28983,I28986,I28989,I28992,I28995,I28998,I29044,I29047,I29050,I29053,I29056,I29059,I29062,I29065,I29068,I29114,I29117,I29120,I29123,I29126,I29129,I29132,I29135,I29181,I29184,I29187,I29190,I29193,I29196,I29199,I29202,I29205,I29251,I29254,I29257,I29260,I29263,I29266,I29269,I29272,I29275,I29321,I29324,I29327,I29330,I29333,I29336,I29339,I29342,I29345,I29391,I29394,I29397,I29400,I29403,I29406,I29409,I29412,I29415,I29418,I29464,I29467,I29470,I29473,I29476,I29479,I29482,I29485,I29488,I29534,I29537,I29540,I29543,I29546,I29549,I29552,I29555,I29558,I29561,I29607,I29610,I29613,I29616,I29619,I29622,I29625,I29628,I29631,I29634,I29680,I29683,I29686,I29689,I29692,I29695,I29698,I29701,I29704,I29750,I29753,I29756,I29759,I29762,I29765,I29768,I29771,I29774,I29820,I29823,I29826,I29829,I29832,I29835,I29838,I29841,I29887,I29890,I29893,I29896,I29899,I29902,I29905,I29908,I29911,I29914,I29960,I29963,I29966,I29969,I29972,I29975,I29978,I29981,I29984,I30030,I30033,I30036,I30039,I30042,I30045,I30048,I30051,I30054,I30100,I30103,I30106,I30109,I30112,I30115,I30118,I30121,I30124,I30170,I30173,I30176,I30179,I30182,I30185,I30188,I30191,I30237,I30240,I30243,I30246,I30249,I30252,I30255,I30258,I30261,I30307,I30310,I30313,I30316,I30319,I30322,I30325,I30328,I30331,I30334,I30380,I30383,I30386,I30389,I30392,I30395,I30398,I30401,I30404,I30407,I30453,I30456,I30459,I30462,I30465,I30468,I30471,I30474,I30520,I30523,I30526,I30529,I30532,I30535,I30538,I30541,I30544,I30590,I30593,I30596,I30599,I30602,I30605,I30608,I30611,I30614,I30660,I30663,I30666,I30669,I30672,I30675,I30678,I30681,I30684,I30730,I30733,I30736,I30739,I30742,I30745,I30748,I30751,I30754,I30800,I30803,I30806,I30809,I30812,I30815,I30818,I30821,I30824,I30827,I30873,I30876,I30879,I30882,I30885,I30888,I30891,I30894,I30940,I30943,I30946,I30949,I30952,I30955,I30958,I30961,I30964,I31010,I31013,I31016,I31019,I31022,I31025,I31028,I31031,I31077,I31080,I31083,I31086,I31089,I31092,I31095,I31098,I31101,I31147,I31150,I31153,I31156,I31159,I31162,I31165,I31168,I31171,I31217,I31220,I31223,I31226,I31229,I31232,I31235,I31238,I31241,I31244,I31290,I31293,I31296,I31299,I31302,I31305,I31308,I31311,I31314,I31360,I31363,I31366,I31369,I31372,I31375,I31378,I31381,I31427,I31430,I31433,I31436,I31439,I31442,I31445,I31448,I31451,I31454,I31500,I31503,I31506,I31509,I31512,I31515,I31518,I31521,I31567,I31570,I31573,I31576,I31579,I31582,I31585,I31588,I31591,I31594,I31640,I31643,I31646,I31649,I31652,I31655,I31658,I31661,I31707,I31710,I31713,I31716,I31719,I31722,I31725,I31728,I31731,I31777,I31780,I31783,I31786,I31789,I31792,I31795,I31798,I31801,I31847,I31850,I31853,I31856,I31859,I31862,I31865,I31868,I31914,I31917,I31920,I31923,I31926,I31929,I31932,I31935,I31938,I31941,I31987,I31990,I31993,I31996,I31999,I32002,I32005,I32008,I32011,I32057,I32060,I32063,I32066,I32069,I32072,I32075,I32078,I32081,I32127,I32130,I32133,I32136,I32139,I32142,I32145,I32148,I32151,I32197,I32200,I32203,I32206,I32209,I32212,I32215,I32218,I32221,I32224,I32270,I32273,I32276,I32279,I32282,I32285,I32288,I32291,I32294,I32297,I32343,I32346,I32349,I32352,I32355,I32358,I32361,I32364,I32367,I32370,I32416,I32419,I32422,I32425,I32428,I32431,I32434,I32437,I32440,I32486,I32489,I32492,I32495,I32498,I32501,I32504,I32507,I32510,I32556,I32559,I32562,I32565,I32568,I32571,I32574,I32577,I32580,I32583,I32629,I32632,I32635,I32638,I32641,I32644,I32647,I32650,I32653,I32656,I32702,I32705,I32708,I32711,I32714,I32717,I32720,I32723,I32726,I32772,I32775,I32778,I32781,I32784,I32787,I32790,I32793,I32796,I32842,I32845,I32848,I32851,I32854,I32857,I32860,I32863,I32866,I32912,I32915,I32918,I32921,I32924,I32927,I32930,I32933,I32936,I32939,I32985,I32988,I32991,I32994,I32997,I33000,I33003,I33006,I33009,I33055,I33058,I33061,I33064,I33067,I33070,I33073,I33076,I33122,I33125,I33128,I33131,I33134,I33137,I33140,I33143,I33189,I33192,I33195,I33198,I33201,I33204,I33207,I33210,I33213,I33259,I33262,I33265,I33268,I33271,I33274,I33277,I33280,I33283,I33329,I33332,I33335,I33338,I33341,I33344,I33347,I33350,I33353,I33399,I33402,I33405,I33408,I33411,I33414,I33417,I33420,I33423,I33469,I33472,I33475,I33478,I33481,I33484,I33487,I33490,I33493,I33496,I33542,I33545,I33548,I33551,I33554,I33557,I33560,I33563,I33566,I33612,I33615,I33618,I33621,I33624,I33627,I33630,I33633,I33636,I33639,I33685,I33688,I33691,I33694,I33697,I33700,I33703,I33706,I33709,I33755,I33758,I33761,I33764,I33767,I33770,I33773,I33776,I33779,I33782,I33828,I33831,I33834,I33837,I33840,I33843,I33846,I33849,I33895,I33898,I33901,I33904,I33907,I33910,I33913,I33916,I33919,I33965,I33968,I33971,I33974,I33977,I33980,I33983,I33986,I33989,I34035,I34038,I34041,I34044,I34047,I34050,I34053,I34056,I34059,I34062,I34108,I34111,I34114,I34117,I34120,I34123,I34126,I34129,I34132,I34178,I34181,I34184,I34187,I34190,I34193,I34196,I34199,I34202,I34248,I34251,I34254,I34257,I34260,I34263,I34266,I34269,I34272,I34275,I34321,I34324,I34327,I34330,I34333,I34336,I34339,I34342,I34345,I34391,I34394,I34397,I34400,I34403,I34406,I34409,I34412,I34415,I34418,I34464,I34467,I34470,I34473,I34476,I34479,I34482,I34485,I34488,I34491,I34537,I34540,I34543,I34546,I34549,I34552,I34555,I34558,I34561,I34607,I34610,I34613,I34616,I34619,I34622,I34625,I34628,I34631,I34634,I34680,I34683,I34686,I34689,I34692,I34695,I34698,I34701,I34704,I34750,I34753,I34756,I34759,I34762,I34765,I34768,I34771,I34774,I34777,I34823,I34826,I34829,I34832,I34835,I34838,I34841,I34844,I34847,I34893,I34896,I34899,I34902,I34905,I34908,I34911,I34914,I34917,I34920,I34966,I34969,I34972,I34975,I34978,I34981,I34984,I34987,I34990,I35036,I35039,I35042,I35045,I35048,I35051,I35054,I35057,I35060,I35106,I35109,I35112,I35115,I35118,I35121,I35124,I35127,I35130,I35133,I35179,I35182,I35185,I35188,I35191,I35194,I35197,I35200,I35246,I35249,I35252,I35255,I35258,I35261,I35264,I35267,I35270,I35316,I35319,I35322,I35325,I35328,I35331,I35334,I35337,I35340,I35386,I35389,I35392,I35395,I35398,I35401,I35404,I35407,I35410,I35413,I35459,I35462,I35465,I35468,I35471,I35474,I35477,I35480,I35483,I35486,I35532,I35535,I35538,I35541,I35544,I35547,I35550,I35553,I35556,I35559,I35605,I35608,I35611,I35614,I35617,I35620,I35623,I35626,I35672,I35675,I35678,I35681,I35684,I35687,I35690,I35693,I35696,I35742,I35745,I35748,I35751,I35754,I35757,I35760,I35763,I35766,I35769,I35815,I35818,I35821,I35824,I35827,I35830,I35833,I35836,I35839,I35842,I35888,I35891,I35894,I35897,I35900,I35903,I35906,I35909,I35912,I35915,I35961,I35964,I35967,I35970,I35973,I35976,I35979,I35982,I35985,I35988,I36034,I36037,I36040,I36043,I36046,I36049,I36052,I36055,I36058,I36061,I36107,I36110,I36113,I36116,I36119,I36122,I36125,I36128,I36131,I36177,I36180,I36183,I36186,I36189,I36192,I36195,I36198,I36201,I36247,I36250,I36253,I36256,I36259,I36262,I36265,I36268,I36271,I36317,I36320,I36323,I36326,I36329,I36332,I36335,I36338,I36341,I36387,I36390,I36393,I36396,I36399,I36402,I36405,I36408,I36411,I36414,I36460,I36463,I36466,I36469,I36472,I36475,I36478,I36481,I36484,I36530,I36533,I36536,I36539,I36542,I36545,I36548,I36551,I36554,I36600,I36603,I36606,I36609,I36612,I36615,I36618,I36621,I36624,I36670,I36673,I36676,I36679,I36682,I36685,I36688,I36691,I36694,I36740,I36743,I36746,I36749,I36752,I36755,I36758,I36761,I36764,I36810,I36813,I36816,I36819,I36822,I36825,I36828,I36831,I36834,I36880,I36883,I36886,I36889,I36892,I36895,I36898,I36901,I36904,I36950,I36953,I36956,I36959,I36962,I36965,I36968,I36971,I37017,I37020,I37023,I37026,I37029,I37032,I37035,I37038,I37041,I37044,I37090,I37093,I37096,I37099,I37102,I37105,I37108,I37111,I37114,I37160,I37163,I37166,I37169,I37172,I37175,I37178,I37181,I37184,I37230,I37233,I37236,I37239,I37242,I37245,I37248,I37251,I37254,I37300,I37303,I37306,I37309,I37312,I37315,I37318,I37321,I37324,I37370,I37373,I37376,I37379,I37382,I37385,I37388,I37391,I37394,I37440,I37443,I37446,I37449,I37452,I37455,I37458,I37461,I37464,I37510,I37513,I37516,I37519,I37522,I37525,I37528,I37531,I37534,I37580,I37583,I37586,I37589,I37592,I37595,I37598,I37601,I37604,I37650,I37653,I37656,I37659,I37662,I37665,I37668,I37671,I37674,I37720,I37723,I37726,I37729,I37732,I37735,I37738,I37741,I37787,I37790,I37793,I37796,I37799,I37802,I37805,I37808,I37811,I37857,I37860,I37863,I37866,I37869,I37872,I37875,I37878,I37881,I37884,I37930,I37933,I37936,I37939,I37942,I37945,I37948,I37951,I37954,I38000,I38003,I38006,I38009,I38012,I38015,I38018,I38021,I38067,I38070,I38073,I38076,I38079,I38082,I38085,I38088,I38091,I38137,I38140,I38143,I38146,I38149,I38152,I38155,I38158,I38204,I38207,I38210,I38213,I38216,I38219,I38222,I38225,I38228,I38231,I38277,I38280,I38283,I38286,I38289,I38292,I38295,I38298,I38301,I38347,I38350,I38353,I38356,I38359,I38362,I38365,I38368,I38371,I38374,I38420,I38423,I38426,I38429,I38432,I38435,I38438,I38441,I38444,I38447,I38493,I38496,I38499,I38502,I38505,I38508,I38511,I38514,I38517,I38563,I38566,I38569,I38572,I38575,I38578,I38581,I38584,I38587,I38633,I38636,I38639,I38642,I38645,I38648,I38651,I38654,I38657,I38703,I38706,I38709,I38712,I38715,I38718,I38721,I38724,I38727,I38730,I38776,I38779,I38782,I38785,I38788,I38791,I38794,I38797,I38800,I38803,I38849,I38852,I38855,I38858,I38861,I38864,I38867,I38870,I38873,I38919,I38922,I38925,I38928,I38931,I38934,I38937,I38940,I38943,I38989,I38992,I38995,I38998,I39001,I39004,I39007,I39010,I39013,I39016,I39062,I39065,I39068,I39071,I39074,I39077,I39080,I39083,I39086,I39089,I39135,I39138,I39141,I39144,I39147,I39150,I39153,I39156,I39159,I39205,I39208,I39211,I39214,I39217,I39220,I39223,I39226,I39229,I39275,I39278,I39281,I39284,I39287,I39290,I39293,I39296,I39299,I39302,I39348,I39351,I39354,I39357,I39360,I39363,I39366,I39369,I39372,I39418,I39421,I39424,I39427,I39430,I39433,I39436,I39439,I39442,I39445,I39491,I39494,I39497,I39500,I39503,I39506,I39509,I39512,I39515,I39561,I39564,I39567,I39570,I39573,I39576,I39579,I39582,I39585,I39588,I39634,I39637,I39640,I39643,I39646,I39649,I39652,I39655,I39658,I39661,I39707,I39710,I39713,I39716,I39719,I39722,I39725,I39728,I39731,I39777,I39780,I39783,I39786,I39789,I39792,I39795,I39798,I39801,I39804,I39850,I39853,I39856,I39859,I39862,I39865,I39868,I39871,I39874,I39877,I39923,I39926,I39929,I39932,I39935,I39938,I39941,I39944,I39947,I39993,I39996,I39999,I40002,I40005,I40008,I40011,I40014,I40017,I40020,I40066,I40069,I40072,I40075,I40078,I40081,I40084,I40087,I40133,I40136,I40139,I40142,I40145,I40148,I40151,I40154,I40157,I40203,I40206,I40209,I40212,I40215,I40218,I40221,I40224,I40227,I40273,I40276,I40279,I40282,I40285,I40288,I40291,I40294,I40340,I40343,I40346,I40349,I40352,I40355,I40358,I40361,I40364,I40367,I40413,I40416,I40419,I40422,I40425,I40428,I40431,I40434,I40437,I40483,I40486,I40489,I40492,I40495,I40498,I40501,I40504,I40507,I40510,I40556,I40559,I40562,I40565,I40568,I40571,I40574,I40577,I40623,I40626,I40629,I40632,I40635,I40638,I40641,I40644,I40647,I40693,I40696,I40699,I40702,I40705,I40708,I40711,I40714,I40717,I40720,I40766,I40769,I40772,I40775,I40778,I40781,I40784,I40787,I40790,I40793,I40839,I40842,I40845,I40848,I40851,I40854,I40857,I40860,I40863,I40866,I40912,I40915,I40918,I40921,I40924,I40927,I40930,I40933,I40936,I40982,I40985,I40988,I40991,I40994,I40997,I41000,I41003,I41006,I41052,I41055,I41058,I41061,I41064,I41067,I41070,I41073,I41076,I41079,I41125,I41128,I41131,I41134,I41137,I41140,I41143,I41146,I41149,I41195,I41198,I41201,I41204,I41207,I41210,I41213,I41216,I41219,I41265,I41268,I41271,I41274,I41277,I41280,I41283,I41286,I41289,I41335,I41338,I41341,I41344,I41347,I41350,I41353,I41356,I41402,I41405,I41408,I41411,I41414,I41417,I41420,I41423,I41426,I41429,I41475,I41478,I41481,I41484,I41487,I41490,I41493,I41496,I41499,I41545,I41548,I41551,I41554,I41557,I41560,I41563,I41566,I41569,I41682,I41685,I41688,I41691,I41694,I41697,I41700,I41703,I41706,I41752,I41755,I41758,I41761,I41764,I41767,I41770,I41773,I41776,I41822,I41825,I41828,I41831,I41834,I41837,I41840,I41843,I41846,I41892,I41895,I41898,I41901,I41904,I41907,I41910,I41913,I41916,I41919,I41965,I41968,I41971,I41974,I41977,I41980,I41983,I41986,I41989,I41992,I42038,I42041,I42044,I42047,I42050,I42053,I42056,I42059,I42062,I42108,I42111,I42114,I42117,I42120,I42123,I42126,I42129,I42175,I42178,I42181,I42184,I42187,I42190,I42193,I42196,I42199,I42245,I42248,I42251,I42254,I42257,I42260,I42263,I42266,I42269,I42315,I42318,I42321,I42324,I42327,I42330,I42333,I42336,I42339,I42385,I42388,I42391,I42394,I42397,I42400,I42403,I42406,I42409,I42412,I42458,I42461,I42464,I42467,I42470,I42473,I42476,I42479,I42482,I42528,I42531,I42534,I42537,I42540,I42543,I42546,I42549,I42552,I42555,I42601,I42604,I42607,I42610,I42613,I42616,I42619,I42622,I42625,I42628,I42674,I42677,I42680,I42683,I42686,I42689,I42692,I42695,I42698,I42744,I42747,I42750,I42753,I42756,I42759,I42762,I42765,I42768,I42814,I42817,I42820,I42823,I42826,I42829,I42832,I42835,I42838,I42884,I42887,I42890,I42893,I42896,I42899,I42902,I42905,I42908,I42954,I42957,I42960,I42963,I42966,I42969,I42972,I42975,I42978,I43024,I43027,I43030,I43033,I43036,I43039,I43042,I43045,I43048,I43051,I43097,I43100,I43103,I43106,I43109,I43112,I43115,I43118,I43121,I43124,I43170,I43173,I43176,I43179,I43182,I43185,I43188,I43191,I43194,I43240,I43243,I43246,I43249,I43252,I43255,I43258,I43261,I43264,I43310,I43313,I43316,I43319,I43322,I43325,I43328,I43331,I43334,I43380,I43383,I43386,I43389,I43392,I43395,I43398,I43401,I43404,I43450,I43453,I43456,I43459,I43462,I43465,I43468,I43471,I43474,I43477,I43523,I43526,I43529,I43532,I43535,I43538,I43541,I43544,I43547,I43550,I43596,I43599,I43602,I43605,I43608,I43611,I43614,I43617,I43663,I43666,I43669,I43672,I43675,I43678,I43681,I43684,I43687,I43690,I43736,I43739,I43742,I43745,I43748,I43751,I43754,I43757,I43760,I43806,I43809,I43812,I43815,I43818,I43821,I43824,I43827,I43830,I43833,I43879,I43882,I43885,I43888,I43891,I43894,I43897,I43900,I43946,I43949,I43952,I43955,I43958,I43961,I43964,I43967,I43970,I43973,I44019,I44022,I44025,I44028,I44031,I44034,I44037,I44040,I44043,I44046,I44092,I44095,I44098,I44101,I44104,I44107,I44110,I44113,I44116,I44119,I44165,I44168,I44171,I44174,I44177,I44180,I44183,I44186,I44189,I44235,I44238,I44241,I44244,I44247,I44250,I44253,I44256,I44302,I44305,I44308,I44311,I44314,I44317,I44320,I44323,I44326,I44372,I44375,I44378,I44381,I44384,I44387,I44390,I44393,I44396,I44442,I44445,I44448,I44451,I44454,I44457,I44460,I44463,I44466,I44469,I44515,I44518,I44521,I44524,I44527,I44530,I44533,I44536,I44539,I44542,I44588,I44591,I44594,I44597,I44600,I44603,I44606,I44609,I44612,I44615,I44661,I44664,I44667,I44670,I44673,I44676,I44679,I44682,I44685,I44688,I44734,I44737,I44740,I44743,I44746,I44749,I44752,I44755,I44758,I44804,I44807,I44810,I44813,I44816,I44819,I44822,I44825,I44828,I44831,I44877,I44880,I44883,I44886,I44889,I44892,I44895,I44898,I44901,I44947,I44950,I44953,I44956,I44959,I44962,I44965,I44968,I44971,I45017,I45020,I45023,I45026,I45029,I45032,I45035,I45038,I45041,I45087,I45090,I45093,I45096,I45099,I45102,I45105,I45108,I45111,I45114,I45160,I45163,I45166,I45169,I45172,I45175,I45178,I45181,I45184,I45230,I45233,I45236,I45239,I45242,I45245,I45248,I45251,I45254,I45257,I45303,I45306,I45309,I45312,I45315,I45318,I45321,I45324,I45327,I45330,I45376,I45379,I45382,I45385,I45388,I45391,I45394,I45397,I45400,I45403,I45449,I45452,I45455,I45458,I45461,I45464,I45467,I45470,I45473,I45519,I45522,I45525,I45528,I45531,I45534,I45537,I45540,I45543,I45589,I45592,I45595,I45598,I45601,I45604,I45607,I45610,I45613,I45616,I45662,I45665,I45668,I45671,I45674,I45677,I45680,I45683,I45686,I45689,I45735,I45738,I45741,I45744,I45747,I45750,I45753,I45756,I45759,I45805,I45808,I45811,I45814,I45817,I45820,I45823,I45826,I45829,I45875,I45878,I45881,I45884,I45887,I45890,I45893,I45896,I45899,I45945,I45948,I45951,I45954,I45957,I45960,I45963,I45966,I45969,I46015,I46018,I46021,I46024,I46027,I46030,I46033,I46036,I46039,I46042,I46088,I46091,I46094,I46097,I46100,I46103,I46106,I46109,I46112,I46158,I46161,I46164,I46167,I46170,I46173,I46176,I46179,I46182,I46228,I46231,I46234,I46237,I46240,I46243,I46246,I46249,I46252,I46298,I46301,I46304,I46307,I46310,I46313,I46316,I46319,I46322,I46368,I46371,I46374,I46377,I46380,I46383,I46386,I46389,I46392,I46395,I46441,I46444,I46447,I46450,I46453,I46456,I46459,I46462,I46508,I46511,I46514,I46517,I46520,I46523,I46526,I46529,I46532,I46578,I46581,I46584,I46587,I46590,I46593,I46596,I46599,I46602,I46605,I46651,I46654,I46657,I46660,I46663,I46666,I46669,I46672,I46675,I46721,I46724,I46727,I46730,I46733,I46736,I46739,I46742,I46745,I46791,I46794,I46797,I46800,I46803,I46806,I46809,I46812,I46815,I46861,I46864,I46867,I46870,I46873,I46876,I46879,I46882,I46885,I46888,I46934,I46937,I46940,I46943,I46946,I46949,I46952,I46955,I46958,I47004,I47007,I47010,I47013,I47016,I47019,I47022,I47025,I47028,I47031,I47077,I47080,I47083,I47086,I47089,I47092,I47095,I47098,I47101,I47147,I47150,I47153,I47156,I47159,I47162,I47165,I47168,I47171,I47217,I47220,I47223,I47226,I47229,I47232,I47235,I47238,I47241,I47244,I47290,I47293,I47296,I47299,I47302,I47305,I47308,I47311,I47314,I47360,I47363,I47366,I47369,I47372,I47375,I47378,I47381,I47384,I47430,I47433,I47436,I47439,I47442,I47445,I47448,I47451,I47454,I47500,I47503,I47506,I47509,I47512,I47515,I47518,I47521,I47524,I47570,I47573,I47576,I47579,I47582,I47585,I47588,I47591,I47594,I47640,I47643,I47646,I47649,I47652,I47655,I47658,I47661,I47664,I47667,I47713,I47716,I47719,I47722,I47725,I47728,I47731,I47734,I47737,I47740,I47786,I47789,I47792,I47795,I47798,I47801,I47804,I47807,I47810,I47813,I47859,I47862,I47865,I47868,I47871,I47874,I47877,I47880,I47883,I47929,I47932,I47935,I47938,I47941,I47944,I47947,I47950,I47996,I47999,I48002,I48005,I48008,I48011,I48014,I48017,I48020,I48023,I48069,I48072,I48075,I48078,I48081,I48084,I48087,I48090,I48136,I48139,I48142,I48145,I48148,I48151,I48154,I48157,I48160,I48206,I48209,I48212,I48215,I48218,I48221,I48224,I48227,I48230,I48276,I48279,I48282,I48285,I48288,I48291,I48294,I48297,I48300,I48346,I48349,I48352,I48355,I48358,I48361,I48364,I48367,I48370,I48416,I48419,I48422,I48425,I48428,I48431,I48434,I48437,I48440,I48486,I48489,I48492,I48495,I48498,I48501,I48504,I48507,I48510,I48513,I48559,I48562,I48565,I48568,I48571,I48574,I48577,I48580,I48583,I48629,I48632,I48635,I48638,I48641,I48644,I48647,I48650,I48653,I48656,I48702,I48705,I48708,I48711,I48714,I48717,I48720,I48723,I48726,I48772,I48775,I48778,I48781,I48784,I48787,I48790,I48793,I48796,I48799,I48845,I48848,I48851,I48854,I48857,I48860,I48863,I48866,I48869,I48872,I48918,I48921,I48924,I48927,I48930,I48933,I48936,I48939,I48942,I48988,I48991,I48994,I48997,I49000,I49003,I49006,I49009,I49012,I49015,I49061,I49064,I49067,I49070,I49073,I49076,I49079,I49082,I49085,I49131,I49134,I49137,I49140,I49143,I49146,I49149,I49152,I49155,I49158,I49204,I49207,I49210,I49213,I49216,I49219,I49222,I49225,I49228,I49274,I49277,I49280,I49283,I49286,I49289,I49292,I49295,I49298,I49301,I49347,I49350,I49353,I49356,I49359,I49362,I49365,I49368,I49371,I49374,I49420,I49423,I49426,I49429,I49432,I49435,I49438,I49441,I49487,I49490,I49493,I49496,I49499,I49502,I49505,I49508,I49511,I49514,I49560,I49563,I49566,I49569,I49572,I49575,I49578,I49581,I49584,I49630,I49633,I49636,I49639,I49642,I49645,I49648,I49651,I49654,I49657,I49703,I49706,I49709,I49712,I49715,I49718,I49721,I49724,I49727,I49773,I49776,I49779,I49782,I49785,I49788,I49791,I49794,I49797,I49843,I49846,I49849,I49852,I49855,I49858,I49861,I49864,I49867,I49913,I49916,I49919,I49922,I49925,I49928,I49931,I49934,I49937,I49983,I49986,I49989,I49992,I49995,I49998,I50001,I50004,I50050,I50053,I50056,I50059,I50062,I50065,I50068,I50071,I50074,I50077,I50123,I50126,I50129,I50132,I50135,I50138,I50141,I50144,I50147,I50193,I50196,I50199,I50202,I50205,I50208,I50211,I50214,I50217,I50263,I50266,I50269,I50272,I50275,I50278,I50281,I50284,I50287,I50290,I50336,I50339,I50342,I50345,I50348,I50351,I50354,I50357,I50360,I50406,I50409,I50412,I50415,I50418,I50421,I50424,I50427,I50430,I50433,I50479,I50482,I50485,I50488,I50491,I50494,I50497,I50500,I50503,I50549,I50552,I50555,I50558,I50561,I50564,I50567,I50570,I50573,I50619,I50622,I50625,I50628,I50631,I50634,I50637,I50640,I50643,I50689,I50692,I50695,I50698,I50701,I50704,I50707,I50710,I50713,I50759,I50762,I50765,I50768,I50771,I50774,I50777,I50780,I50783,I50786,I50832,I50835,I50838,I50841,I50844,I50847,I50850,I50853,I50856,I50902,I50905,I50908,I50911,I50914,I50917,I50920,I50923,I50926,I50972,I50975,I50978,I50981,I50984,I50987,I50990,I50993,I50996,I50999,I51045,I51048,I51051,I51054,I51057,I51060,I51063,I51066,I51069,I51115,I51118,I51121,I51124,I51127,I51130,I51133,I51136,I51139,I51185,I51188,I51191,I51194,I51197,I51200,I51203,I51206,I51209,I51255,I51258,I51261,I51264,I51267,I51270,I51273,I51276,I51279,I51325,I51328,I51331,I51334,I51337,I51340,I51343,I51346,I51392,I51395,I51398,I51401,I51404,I51407,I51410,I51413,I51416,I51462,I51465,I51468,I51471,I51474,I51477,I51480,I51483,I51486,I51532,I51535,I51538,I51541,I51544,I51547,I51550,I51553,I51556,I51559,I51605,I51608,I51611,I51614,I51617,I51620,I51623,I51626,I51629,I51632,I51678,I51681,I51684,I51687,I51690,I51693,I51696,I51699,I51702,I51748,I51751,I51754,I51757,I51760,I51763,I51766,I51769,I51772,I51818,I51821,I51824,I51827,I51830,I51833,I51836,I51839,I51842,I51845,I51891,I51894,I51897,I51900,I51903,I51906,I51909,I51912,I51915,I51961,I51964,I51967,I51970,I51973,I51976,I51979,I51982,I51985,I51988,I52034,I52037,I52040,I52043,I52046,I52049,I52052,I52055,I52058,I52104,I52107,I52110,I52113,I52116,I52119,I52122,I52125,I52128,I52174,I52177,I52180,I52183,I52186,I52189,I52192,I52195,I52198,I52244,I52247,I52250,I52253,I52256,I52259,I52262,I52265,I52268,I52271,I52317,I52320,I52323,I52326,I52329,I52332,I52335,I52338,I52341,I52344,I52390,I52393,I52396,I52399,I52402,I52405,I52408,I52411,I52414,I52460,I52463,I52466,I52469,I52472,I52475,I52478,I52481,I52484,I52530,I52533,I52536,I52539,I52542,I52545,I52548,I52551,I52554,I52600,I52603,I52606,I52609,I52612,I52615,I52618,I52621,I52624,I52670,I52673,I52676,I52679,I52682,I52685,I52688,I52691,I52694,I52740,I52743,I52746,I52749,I52752,I52755,I52758,I52761,I52764,I52810,I52813,I52816,I52819,I52822,I52825,I52828,I52831,I52877,I52880,I52883,I52886,I52889,I52892,I52895,I52898,I52901,I52904,I52950,I52953,I52956,I52959,I52962,I52965,I52968,I52971,I52974,I53020,I53023,I53026,I53029,I53032,I53035,I53038,I53041,I53044,I53090,I53093,I53096,I53099,I53102,I53105,I53108,I53111,I53114,I53160,I53163,I53166,I53169,I53172,I53175,I53178,I53181,I53184,I53187,I53233,I53236,I53239,I53242,I53245,I53248,I53251,I53254,I53257,I53260,I53306,I53309,I53312,I53315,I53318,I53321,I53324,I53327,I53330,I53376,I53379,I53382,I53385,I53388,I53391,I53394,I53397,I53400,I53446,I53449,I53452,I53455,I53458,I53461,I53464,I53467,I53470,I53473,I53519,I53522,I53525,I53528,I53531,I53534,I53537,I53540,I53543,I53589,I53592,I53595,I53598,I53601,I53604,I53607,I53610,I53613,I53659,I53662,I53665,I53668,I53671,I53674,I53677,I53680,I53683,I53729,I53732,I53735,I53738,I53741,I53744,I53747,I53750,I53753,I53799,I53802,I53805,I53808,I53811,I53814,I53817,I53820,I53823,I53869,I53872,I53875,I53878,I53881,I53884,I53887,I53890,I53893,I53939,I53942,I53945,I53948,I53951,I53954,I53957,I53960,I54006,I54009,I54012,I54015,I54018,I54021,I54024,I54027,I54030,I54033,I54079,I54082,I54085,I54088,I54091,I54094,I54097,I54100,I54146,I54149,I54152,I54155,I54158,I54161,I54164,I54167,I54170,I54216,I54219,I54222,I54225,I54228,I54231,I54234,I54237,I54240,I54286,I54289,I54292,I54295,I54298,I54301,I54304,I54307,I54310,I54313,I54359,I54362,I54365,I54368,I54371,I54374,I54377,I54380,I54383,I54386,I54432,I54435,I54438,I54441,I54444,I54447,I54450,I54453,I54499,I54502,I54505,I54508,I54511,I54514,I54517,I54520,I54523,I54569,I54572,I54575,I54578,I54581,I54584,I54587,I54590,I54593,I54639,I54642,I54645,I54648,I54651,I54654,I54657,I54660,I54663,I54709,I54712,I54715,I54718,I54721,I54724,I54727,I54730,I54733,I54736,I54782,I54785,I54788,I54791,I54794,I54797,I54800,I54803,I54806,I54809,I54855,I54858,I54861,I54864,I54867,I54870,I54873,I54876,I54879,I54925,I54928,I54931,I54934,I54937,I54940,I54943,I54946,I54949,I54952,I54998,I55001,I55004,I55007,I55010,I55013,I55016,I55019,I55022,I55068,I55071,I55074,I55077,I55080,I55083,I55086,I55089,I55092,I55138,I55141,I55144,I55147,I55150,I55153,I55156,I55159,I55162,I55208,I55211,I55214,I55217,I55220,I55223,I55226,I55229,I55232,I55235,I55281,I55284,I55287,I55290,I55293,I55296,I55299,I55302,I55305,I55351,I55354,I55357,I55360,I55363,I55366,I55369,I55372,I55375,I55421,I55424,I55427,I55430,I55433,I55436,I55439,I55442,I55445,I55448,I55494,I55497,I55500,I55503,I55506,I55509,I55512,I55515,I55561,I55564,I55567,I55570,I55573,I55576,I55579,I55582,I55628,I55631,I55634,I55637,I55640,I55643,I55646,I55649,I55652,I55655,I55701,I55704,I55707,I55710,I55713,I55716,I55719,I55722,I55725,I55771,I55774,I55777,I55780,I55783,I55786,I55789,I55792,I55795,I55798,I55844,I55847,I55850,I55853,I55856,I55859,I55862,I55865,I55868,I55914,I55917,I55920,I55923,I55926,I55929,I55932,I55935,I55938,I55984,I55987,I55990,I55993,I55996,I55999,I56002,I56005,I56008,I56011,I56057,I56060,I56063,I56066,I56069,I56072,I56075,I56078,I56081,I56127,I56130,I56133,I56136,I56139,I56142,I56145,I56148,I56151,I56154,I56200,I56203,I56206,I56209,I56212,I56215,I56218,I56221,I56224,I56270,I56273,I56276,I56279,I56282,I56285,I56288,I56291,I56294,I56297,I56343,I56346,I56349,I56352,I56355,I56358,I56361,I56364,I56367,I56370,I56416,I56419,I56422,I56425,I56428,I56431,I56434,I56437,I56440,I56486,I56489,I56492,I56495,I56498,I56501,I56504,I56507,I56510,I56556,I56559,I56562,I56565,I56568,I56571,I56574,I56577,I56580,I56626,I56629,I56632,I56635,I56638,I56641,I56644,I56647,I56650,I56653,I56699,I56702,I56705,I56708,I56711,I56714,I56717,I56720,I56723,I56726,I56772,I56775,I56778,I56781,I56784,I56787,I56790,I56793,I56796,I56842,I56845,I56848,I56851,I56854,I56857,I56860,I56863,I56866,I56869,I56915,I56918,I56921,I56924,I56927,I56930,I56933,I56936,I56982,I56985,I56988,I56991,I56994,I56997,I57000,I57003,I57006,I57052,I57055,I57058,I57061,I57064,I57067,I57070,I57073,I57076,I57122,I57125,I57128,I57131,I57134,I57137,I57140,I57143,I57146,I57192,I57195,I57198,I57201,I57204,I57207,I57210,I57213,I57216,I57219,I57265,I57268,I57271,I57274,I57277,I57280,I57283,I57286,I57289,I57292,I57338,I57341,I57344,I57347,I57350,I57353,I57356,I57359,I57362,I57408,I57411,I57414,I57417,I57420,I57423,I57426,I57429,I57432,I57478,I57481,I57484,I57487,I57490,I57493,I57496,I57499,I57502,I57505,I57551,I57554,I57557,I57560,I57563,I57566,I57569,I57572,I57575,I57578,I57624,I57627,I57630,I57633,I57636,I57639,I57642,I57645,I57648,I57694,I57697,I57700,I57703,I57706,I57709,I57712,I57715,I57718,I57764,I57767,I57770,I57773,I57776,I57779,I57782,I57785,I57788,I57791,I57837,I57840,I57843,I57846,I57849,I57852,I57855,I57858,I57861,I57864,I57910,I57913,I57916,I57919,I57922,I57925,I57928,I57931,I57934,I57980,I57983,I57986,I57989,I57992,I57995,I57998,I58001,I58004,I58050,I58053,I58056,I58059,I58062,I58065,I58068,I58071,I58074,I58077,I58123,I58126,I58129,I58132,I58135,I58138,I58141,I58144,I58147,I58193,I58196,I58199,I58202,I58205,I58208,I58211,I58214,I58217,I58263,I58266,I58269,I58272,I58275,I58278,I58281,I58284,I58330,I58333,I58336,I58339,I58342,I58345,I58348,I58351,I58354,I58357,I58403,I58406,I58409,I58412,I58415,I58418,I58421,I58424,I58427,I58473,I58476,I58479,I58482,I58485,I58488,I58491,I58494,I58497,I58500,I58546,I58549,I58552,I58555,I58558,I58561,I58564,I58567,I58570,I58573,I58619,I58622,I58625,I58628,I58631,I58634,I58637,I58640,I58643,I58646,I58692,I58695,I58698,I58701,I58704,I58707,I58710,I58713,I58716,I58719,I58765,I58768,I58771,I58774,I58777,I58780,I58783,I58786,I58789,I58835,I58838,I58841,I58844,I58847,I58850,I58853,I58856,I58859,I58862,I58908,I58911,I58914,I58917,I58920,I58923,I58926,I58929,I58932,I58978,I58981,I58984,I58987,I58990,I58993,I58996,I58999,I59045,I59048,I59051,I59054,I59057,I59060,I59063,I59066,I59069,I59115,I59118,I59121,I59124,I59127,I59130,I59133,I59136,I59139,I59185,I59188,I59191,I59194,I59197,I59200,I59203,I59206,I59209,I59212,I59258,I59261,I59264,I59267,I59270,I59273,I59276,I59279,I59325,I59328,I59331,I59334,I59337,I59340,I59343,I59346,I59392,I59395,I59398,I59401,I59404,I59407,I59410,I59413,I59416,I59462,I59465,I59468,I59471,I59474,I59477,I59480,I59483,I59486,I59489,I59535,I59538,I59541,I59544,I59547,I59550,I59553,I59556,I59559,I59605,I59608,I59611,I59614,I59617,I59620,I59623,I59626,I59629,I59675,I59678,I59681,I59684,I59687,I59690,I59693,I59696,I59699,I59702,I59748,I59751,I59754,I59757,I59760,I59763,I59766,I59769,I59772,I59775,I59821,I59824,I59827,I59830,I59833,I59836,I59839,I59842,I59845,I59891,I59894,I59897,I59900,I59903,I59906,I59909,I59912,I59915,I59918,I59964,I59967,I59970,I59973,I59976,I59979,I59982,I59985,I59988,I59991,I60037,I60040,I60043,I60046,I60049,I60052,I60055,I60058,I60061,I60107,I60110,I60113,I60116,I60119,I60122,I60125,I60128,I60131,I60134,I60180,I60183,I60186,I60189,I60192,I60195,I60198,I60201,I60204,I60250,I60253,I60256,I60259,I60262,I60265,I60268,I60271,I60274,I60320,I60323,I60326,I60329,I60332,I60335,I60338,I60341,I60344,I60390,I60393,I60396,I60399,I60402,I60405,I60408,I60411,I60414,I60460,I60463,I60466,I60469,I60472,I60475,I60478,I60481,I60484,I60487,I60533,I60536,I60539,I60542,I60545,I60548,I60551,I60554,I60557,I60603,I60606,I60609,I60612,I60615,I60618,I60621,I60624,I60627,I60673,I60676,I60679,I60682,I60685,I60688,I60691,I60694,I60697,I60743,I60746,I60749,I60752,I60755,I60758,I60761,I60764,I60767,I60813,I60816,I60819,I60822,I60825,I60828,I60831,I60834,I60837,I60883,I60886,I60889,I60892,I60895,I60898,I60901,I60904,I60907,I60910,I60956,I60959,I60962,I60965,I60968,I60971,I60974,I60977,I61023,I61026,I61029,I61032,I61035,I61038,I61041,I61044,I61047,I61093,I61096,I61099,I61102,I61105,I61108,I61111,I61114,I61117,I61163,I61166,I61169,I61172,I61175,I61178,I61181,I61184,I61230,I61233,I61236,I61239,I61242,I61245,I61248,I61251,I61254,I61257,I61303,I61306,I61309,I61312,I61315,I61318,I61321,I61324,I61443,I61446,I61449,I61452,I61455,I61458,I61461,I61464,I61467,I61513,I61516,I61519,I61522,I61525,I61528,I61531,I61534,I61537,I61583,I61586,I61589,I61592,I61595,I61598,I61601,I61604,I61650,I61653,I61656,I61659,I61662,I61665,I61668,I61671,I61674,I61720,I61723,I61726,I61729,I61732,I61735,I61738,I61741,I61744,I61747,I61793,I61796,I61799,I61802,I61805,I61808,I61811,I61814,I61817,I61863,I61866,I61869,I61872,I61875,I61878,I61881,I61884,I61887,I61890,I61936,I61939,I61942,I61945,I61948,I61951,I61954,I61957,I61960,I61963,I62009,I62012,I62015,I62018,I62021,I62024,I62027,I62030,I62033,I62036,I62082,I62085,I62088,I62091,I62094,I62097,I62100,I62103,I62106,I62152,I62155,I62158,I62161,I62164,I62167,I62170,I62173,I62176,I62222,I62225,I62228,I62231,I62234,I62237,I62240,I62243,I62246,I62292,I62295,I62298,I62301,I62304,I62307,I62310,I62313,I62316,I62362,I62365,I62368,I62371,I62374,I62377,I62380,I62383,I62386,I62432,I62435,I62438,I62441,I62444,I62447,I62450,I62453,I62456,I62459,I62505,I62508,I62511,I62514,I62517,I62520,I62523,I62526,I62529,I62575,I62578,I62581,I62584,I62587,I62590,I62593,I62596,I62599,I62645,I62648,I62651,I62654,I62657,I62660,I62663,I62666,I62669,I62715,I62718,I62721,I62724,I62727,I62730,I62733,I62736,I62739,I62785,I62788,I62791,I62794,I62797,I62800,I62803,I62806,I62809,I62855,I62858,I62861,I62864,I62867,I62870,I62873,I62876,I62879,I62882,I62928,I62931,I62934,I62937,I62940,I62943,I62946,I62949,I62952,I62955,I63001,I63004,I63007,I63010,I63013,I63016,I63019,I63022,I63025,I63071,I63074,I63077,I63080,I63083,I63086,I63089,I63092,I63095,I63098,I63144,I63147,I63150,I63153,I63156,I63159,I63162,I63165,I63168,I63171,I63217,I63220,I63223,I63226,I63229,I63232,I63235,I63238,I63241,I63244,I63290,I63293,I63296,I63299,I63302,I63305,I63308,I63311,I63314,I63360,I63363,I63366,I63369,I63372,I63375,I63378,I63381,I63384,I63430,I63433,I63436,I63439,I63442,I63445,I63448,I63451,I63454,I63500,I63503,I63506,I63509,I63512,I63515,I63518,I63521,I63524,I63527,I63573,I63576,I63579,I63582,I63585,I63588,I63591,I63594,I63597,I63643,I63646,I63649,I63652,I63655,I63658,I63661,I63664,I63667,I63670,I63716,I63719,I63722,I63725,I63728,I63731,I63734,I63737,I63740,I63786,I63789,I63792,I63795,I63798,I63801,I63804,I63807,I63810,I63813,I63859,I63862,I63865,I63868,I63871,I63874,I63877,I63880,I63883,I63929,I63932,I63935,I63938,I63941,I63944,I63947,I63950,I63953,I63999,I64002,I64005,I64008,I64011,I64014,I64017,I64020,I64023,I64069,I64072,I64075,I64078,I64081,I64084,I64087,I64090,I64093,I64096,I64142,I64145,I64148,I64151,I64154,I64157,I64160,I64163,I64166,I64169,I64215,I64218,I64221,I64224,I64227,I64230,I64233,I64236,I64282,I64285,I64288,I64291,I64294,I64297,I64300,I64303,I64306,I64352,I64355,I64358,I64361,I64364,I64367,I64370,I64373,I64376,I64422,I64425,I64428,I64431,I64434,I64437,I64440,I64443,I64446,I64449,I64495,I64498,I64501,I64504,I64507,I64510,I64513,I64516,I64562,I64565,I64568,I64571,I64574,I64577,I64580,I64583,I64586,I64589,I64635,I64638,I64641,I64644,I64647,I64650,I64653,I64656,I64659,I64705,I64708,I64711,I64714,I64717,I64720,I64723,I64726,I64729,I64775,I64778,I64781,I64784,I64787,I64790,I64793,I64796,I64799,I64802,I64848,I64851,I64854,I64857,I64860,I64863,I64866,I64869,I64872,I64875,I64921,I64924,I64927,I64930,I64933,I64936,I64939,I64942,I64945,I64991,I64994,I64997,I65000,I65003,I65006,I65009,I65012,I65015,I65061,I65064,I65067,I65070,I65073,I65076,I65079,I65082,I65085,I65131,I65134,I65137,I65140,I65143,I65146,I65149,I65152,I65155,I65201,I65204,I65207,I65210,I65213,I65216,I65219,I65222,I65225,I65228,I65274,I65277,I65280,I65283,I65286,I65289,I65292,I65295,I65298,I65344,I65347,I65350,I65353,I65356,I65359,I65362,I65365,I65368,I65371,I65417,I65420,I65423,I65426,I65429,I65432,I65435,I65438,I65484,I65487,I65490,I65493,I65496,I65499,I65502,I65505,I65508,I65511,I65557,I65560,I65563,I65566,I65569,I65572,I65575,I65578,I65624,I65627,I65630,I65633,I65636,I65639,I65642,I65645,I65648,I65694,I65697,I65700,I65703,I65706,I65709,I65712,I65715,I65718,I65721,I65767,I65770,I65773,I65776,I65779,I65782,I65785,I65788,I65834,I65837,I65840,I65843,I65846,I65849,I65852,I65855,I65858,I65904,I65907,I65910,I65913,I65916,I65919,I65922,I65925,I65928,I65974,I65977,I65980,I65983,I65986,I65989,I65992,I65995,I65998,I66044,I66047,I66050,I66053,I66056,I66059,I66062,I66065,I66068,I66071,I66117,I66120,I66123,I66126,I66129,I66132,I66135,I66138,I66141,I66144,I66190,I66193,I66196,I66199,I66202,I66205,I66208,I66211,I66214,I66260,I66263,I66266,I66269,I66272,I66275,I66278,I66281,I66284,I66330,I66333,I66336,I66339,I66342,I66345,I66348,I66351,I66354,I66400,I66403,I66406,I66409,I66412,I66415,I66418,I66421,I66424,I66427,I66473,I66476,I66479,I66482,I66485,I66488,I66491,I66494,I66497,I66500,I66546,I66549,I66552,I66555,I66558,I66561,I66564,I66567,I66570,I66616,I66619,I66622,I66625,I66628,I66631,I66634,I66637,I66640,I66686,I66689,I66692,I66695,I66698,I66701,I66704,I66707,I66753,I66756,I66759,I66762,I66765,I66768,I66771,I66774,I66777,I66780,I66826,I66829,I66832,I66835,I66838,I66841,I66844,I66847,I66850,I66896,I66899,I66902,I66905,I66908,I66911,I66914,I66917,I66920,I66966,I66969,I66972,I66975,I66978,I66981,I66984,I66987,I67033,I67036,I67039,I67042,I67045,I67048,I67051,I67054,I67057,I67103,I67106,I67109,I67112,I67115,I67118,I67121,I67124,I67127,I67173,I67176,I67179,I67182,I67185,I67188,I67191,I67194,I67197,I67200,I67246,I67249,I67252,I67255,I67258,I67261,I67264,I67267,I67270,I67316,I67319,I67322,I67325,I67328,I67331,I67334,I67337,I67340,I67343,I67389,I67392,I67395,I67398,I67401,I67404,I67407,I67410,I67413,I67459,I67462,I67465,I67468,I67471,I67474,I67477,I67480,I67483,I67529,I67532,I67535,I67538,I67541,I67544,I67547,I67550,I67553,I67556,I67602,I67605,I67608,I67611,I67614,I67617,I67620,I67623,I67669,I67672,I67675,I67678,I67681,I67684,I67687,I67690,I67736,I67739,I67742,I67745,I67748,I67751,I67754,I67757,I67760,I67806,I67809,I67812,I67815,I67818,I67821,I67824,I67827,I67830,I67876,I67879,I67882,I67885,I67888,I67891,I67894,I67897,I67900,I67946,I67949,I67952,I67955,I67958,I67961,I67964,I67967,I67970,I68016,I68019,I68022,I68025,I68028,I68031,I68034,I68037,I68040,I68086,I68089,I68092,I68095,I68098,I68101,I68104,I68107,I68110,I68156,I68159,I68162,I68165,I68168,I68171,I68174,I68177,I68180,I68183,I68229,I68232,I68235,I68238,I68241,I68244,I68247,I68250,I68253,I68256,I68302,I68305,I68308,I68311,I68314,I68317,I68320,I68323,I68326,I68372,I68375,I68378,I68381,I68384,I68387,I68390,I68393,I68396,I68399,I68445,I68448,I68451,I68454,I68457,I68460,I68463,I68466,I68469,I68472,I68518,I68521,I68524,I68527,I68530,I68533,I68536,I68539,I68585,I68588,I68591,I68594,I68597,I68600,I68603,I68606,I68652,I68655,I68658,I68661,I68664,I68667,I68670,I68673,I68676,I68679,I68725,I68728,I68731,I68734,I68737,I68740,I68743,I68746,I68749,I68795,I68798,I68801,I68804,I68807,I68810,I68813,I68816,I68819,I68822,I68868,I68871,I68874,I68877,I68880,I68883,I68886,I68889,I68892,I68938,I68941,I68944,I68947,I68950,I68953,I68956,I68959,I68962,I68965,I69011,I69014,I69017,I69020,I69023,I69026,I69029,I69032,I69035,I69081,I69084,I69087,I69090,I69093,I69096,I69099,I69102,I69105,I69151,I69154,I69157,I69160,I69163,I69166,I69169,I69172,I69175,I69221,I69224,I69227,I69230,I69233,I69236,I69239,I69242,I69245,I69291,I69294,I69297,I69300,I69303,I69306,I69309,I69312,I69315,I69361,I69364,I69367,I69370,I69373,I69376,I69379,I69382,I69428,I69431,I69434,I69437,I69440,I69443,I69446,I69449,I69452,I69455,I69501,I69504,I69507,I69510,I69513,I69516,I69519,I69522,I69525,I69571,I69574,I69577,I69580,I69583,I69586,I69589,I69592,I69638,I69641,I69644,I69647,I69650,I69653,I69656,I69659,I69662,I69708,I69711,I69714,I69717,I69720,I69723,I69726,I69729,I69732,I69778,I69781,I69784,I69787,I69790,I69793,I69796,I69799,I69802,I69848,I69851,I69854,I69857,I69860,I69863,I69866,I69869,I69872,I69875,I69921,I69924,I69927,I69930,I69933,I69936,I69939,I69942,I69945,I69991,I69994,I69997,I70000,I70003,I70006,I70009,I70012,I70015,I70018,I70064,I70067,I70070,I70073,I70076,I70079,I70082,I70085,I70088,I70091,I70137,I70140,I70143,I70146,I70149,I70152,I70155,I70158,I70161,I70207,I70210,I70213,I70216,I70219,I70222,I70225,I70228,I70231,I70277,I70280,I70283,I70286,I70289,I70292,I70295,I70298,I70301,I70347,I70350,I70353,I70356,I70359,I70362,I70365,I70368,I70371,I70374,I70420,I70423,I70426,I70429,I70432,I70435,I70438,I70441,I70444,I70490,I70493,I70496,I70499,I70502,I70505,I70508,I70511,I70514,I70560,I70563,I70566,I70569,I70572,I70575,I70578,I70581,I70627,I70630,I70633,I70636,I70639,I70642,I70645,I70648,I70651,I70697,I70700,I70703,I70706,I70709,I70712,I70715,I70718,I70721,I70724,I70770,I70773,I70776,I70779,I70782,I70785,I70788,I70791,I70794,I70840,I70843,I70846,I70849,I70852,I70855,I70858,I70861,I70864,I70910,I70913,I70916,I70919,I70922,I70925,I70928,I70931,I70977,I70980,I70983,I70986,I70989,I70992,I70995,I70998,I71001,I71047,I71050,I71053,I71056,I71059,I71062,I71065,I71068,I71071,I71117,I71120,I71123,I71126,I71129,I71132,I71135,I71138,I71141,I71187,I71190,I71193,I71196,I71199,I71202,I71205,I71208,I71211,I71257,I71260,I71263,I71266,I71269,I71272,I71275,I71278,I71281,I71284,I71330,I71333,I71336,I71339,I71342,I71345,I71348,I71351,I71354,I71357,I71403,I71406,I71409,I71412,I71415,I71418,I71421,I71424,I71427,I71430,I71476,I71479,I71482,I71485,I71488,I71491,I71494,I71497,I71500,I71503,I71549,I71552,I71555,I71558,I71561,I71564,I71567,I71570,I71573,I71619,I71622,I71625,I71628,I71631,I71634,I71637,I71640,I71643,I71689,I71692,I71695,I71698,I71701,I71704,I71707,I71710,I71713,I71759,I71762,I71765,I71768,I71771,I71774,I71777,I71780,I71783,I71829,I71832,I71835,I71838,I71841,I71844,I71847,I71850,I71896,I71899,I71902,I71905,I71908,I71911,I71914,I71917,I71920,I71966,I71969,I71972,I71975,I71978,I71981,I71984,I71987,I72033,I72036,I72039,I72042,I72045,I72048,I72051,I72054,I72057,I72103,I72106,I72109,I72112,I72115,I72118,I72121,I72124,I72127,I72173,I72176,I72179,I72182,I72185,I72188,I72191,I72194,I72197,I72200,I72246,I72249,I72252,I72255,I72258,I72261,I72264,I72267,I72270,I72316,I72319,I72322,I72325,I72328,I72331,I72334,I72337,I72340,I72343,I72389,I72392,I72395,I72398,I72401,I72404,I72407,I72410,I72413,I72459,I72462,I72465,I72468,I72471,I72474,I72477,I72480,I72483,I72529,I72532,I72535,I72538,I72541,I72544,I72547,I72550,I72553,I72599,I72602,I72605,I72608,I72611,I72614,I72617,I72620,I72623,I72626,I72672,I72675,I72678,I72681,I72684,I72687,I72690,I72693,I72696,I72699,I72745,I72748,I72751,I72754,I72757,I72760,I72763,I72766,I72769,I72772,I72818,I72821,I72824,I72827,I72830,I72833,I72836,I72839,I72842,I72888,I72891,I72894,I72897,I72900,I72903,I72906,I72909,I72912,I72958,I72961,I72964,I72967,I72970,I72973,I72976,I72979,I72982,I72985,I73031,I73034,I73037,I73040,I73043,I73046,I73049,I73052,I73055,I73101,I73104,I73107,I73110,I73113,I73116,I73119,I73122,I73125,I73128,I73174,I73177,I73180,I73183,I73186,I73189,I73192,I73195,I73198,I73244,I73247,I73250,I73253,I73256,I73259,I73262,I73265,I73311,I73314,I73317,I73320,I73323,I73326,I73329,I73332,I73335,I73338,I73384,I73387,I73390,I73393,I73396,I73399,I73402,I73405,I73408,I73454,I73457,I73460,I73463,I73466,I73469,I73472,I73475,I73478,I73524,I73527,I73530,I73533,I73536,I73539,I73542,I73545,I73548,I73594,I73597,I73600,I73603,I73606,I73609,I73612,I73615,I73618,I73664,I73667,I73670,I73673,I73676,I73679,I73682,I73685,I73688,I73734,I73737,I73740,I73743,I73746,I73749,I73752,I73755,I73758,I73761,I73807,I73810,I73813,I73816,I73819,I73822,I73825,I73828,I73874,I73877,I73880,I73883,I73886,I73889,I73892,I73895,I73898,I73944,I73947,I73950,I73953,I73956,I73959,I73962,I73965,I73968,I74014,I74017,I74020,I74023,I74026,I74029,I74032,I74035,I74038,I74084,I74087,I74090,I74093,I74096,I74099,I74102,I74105,I74108,I74154,I74157,I74160,I74163,I74166,I74169,I74172,I74175,I74178,I74181,I74227,I74230,I74233,I74236,I74239,I74242,I74245,I74248,I74294,I74297,I74300,I74303,I74306,I74309,I74312,I74315,I74318,I74364,I74367,I74370,I74373,I74376,I74379,I74382,I74385,I74388,I74391,I74437,I74440,I74443,I74446,I74449,I74452,I74455,I74458,I74461,I74507,I74510,I74513,I74516,I74519,I74522,I74525,I74528,I74531,I74577,I74580,I74583,I74586,I74589,I74592,I74595,I74598,I74601,I74604,I74650,I74653,I74656,I74659,I74662,I74665,I74668,I74671,I74674,I74677,I74723,I74726,I74729,I74732,I74735,I74738,I74741,I74744,I74747,I74793,I74796,I74799,I74802,I74805,I74808,I74811,I74814,I74817,I74863,I74866,I74869,I74872,I74875,I74878,I74881,I74884,I74887,I74890,I74936,I74939,I74942,I74945,I74948,I74951,I74954,I74957,I74960,I75006,I75009,I75012,I75015,I75018,I75021,I75024,I75027,I75030,I75033,I75079,I75082,I75085,I75088,I75091,I75094,I75097,I75100,I75103,I75106,I75152,I75155,I75158,I75161,I75164,I75167,I75170,I75173,I75176,I75222,I75225,I75228,I75231,I75234,I75237,I75240,I75243,I75246,I75292,I75295,I75298,I75301,I75304,I75307,I75310,I75313,I75316,I75362,I75365,I75368,I75371,I75374,I75377,I75380,I75383,I75386,I75389,I75435,I75438,I75441,I75444,I75447,I75450,I75453,I75456,I75459,I75505,I75508,I75511,I75514,I75517,I75520,I75523,I75526,I75529,I75532,I75578,I75581,I75584,I75587,I75590,I75593,I75596,I75599,I75602,I75648,I75651,I75654,I75657,I75660,I75663,I75666,I75669,I75672,I75718,I75721,I75724,I75727,I75730,I75733,I75736,I75739,I75742,I75745,I75791,I75794,I75797,I75800,I75803,I75806,I75809,I75812,I75858,I75861,I75864,I75867,I75870,I75873,I75876,I75879,I75882,I75928,I75931,I75934,I75937,I75940,I75943,I75946,I75949,I75995,I75998,I76001,I76004,I76007,I76010,I76013,I76016,I76019,I76065,I76068,I76071,I76074,I76077,I76080,I76083,I76086,I76089,I76092,I76138,I76141,I76144,I76147,I76150,I76153,I76156,I76159,I76162,I76208,I76211,I76214,I76217,I76220,I76223,I76226,I76229,I76275,I76278,I76281,I76284,I76287,I76290,I76293,I76296,I76299,I76345,I76348,I76351,I76354,I76357,I76360,I76363,I76366,I76369,I76372,I76418,I76421,I76424,I76427,I76430,I76433,I76436,I76439,I76442,I76488,I76491,I76494,I76497,I76500,I76503,I76506,I76509,I76512,I76515,I76561,I76564,I76567,I76570,I76573,I76576,I76579,I76582,I76585,I76631,I76634,I76637,I76640,I76643,I76646,I76649,I76652,I76655,I76658,I76704,I76707,I76710,I76713,I76716,I76719,I76722,I76725,I76728,I76731,I76777,I76780,I76783,I76786,I76789,I76792,I76795,I76798,I76801,I76847,I76850,I76853,I76856,I76859,I76862,I76865,I76868,I76871,I76874,I76920,I76923,I76926,I76929,I76932,I76935,I76938,I76941,I76944,I76990,I76993,I76996,I76999,I77002,I77005,I77008,I77011,I77014,I77017,I77063,I77066,I77069,I77072,I77075,I77078,I77081,I77084,I77087,I77133,I77136,I77139,I77142,I77145,I77148,I77151,I77154,I77157,I77160,I77206,I77209,I77212,I77215,I77218,I77221,I77224,I77227,I77230,I77276,I77279,I77282,I77285,I77288,I77291,I77294,I77297,I77300,I77303,I77349,I77352,I77355,I77358,I77361,I77364,I77367,I77370,I77373,I77419,I77422,I77425,I77428,I77431,I77434,I77437,I77440,I77443,I77446,I77492,I77495,I77498,I77501,I77504,I77507,I77510,I77513,I77559,I77562,I77565,I77568,I77571,I77574,I77577,I77580,I77583,I77629,I77632,I77635,I77638,I77641,I77644,I77647,I77650,I77696,I77699,I77702,I77705,I77708,I77711,I77714,I77717,I77720,I77723,I77769,I77772,I77775,I77778,I77781,I77784,I77787,I77790,I77793,I77796,I77842,I77845,I77848,I77851,I77854,I77857,I77860,I77863,I77866,I77912,I77915,I77918,I77921,I77924,I77927,I77930,I77933,I77936,I77939,I77985,I77988,I77991,I77994,I77997,I78000,I78003,I78006,I78009,I78055,I78058,I78061,I78064,I78067,I78070,I78073,I78076,I78079,I78082,I78128,I78131,I78134,I78137,I78140,I78143,I78146,I78149,I78195,I78198,I78201,I78204,I78207,I78210,I78213,I78216,I78219,I78222,I78268,I78271,I78274,I78277,I78280,I78283,I78286,I78289,I78292,I78338,I78341,I78344,I78347,I78350,I78353,I78356,I78359,I78405,I78408,I78411,I78414,I78417,I78420,I78423,I78426,I78429,I78475,I78478,I78481,I78484,I78487,I78490,I78493,I78496,I78542,I78545,I78548,I78551,I78554,I78557,I78560,I78563,I78566,I78569,I78615,I78618,I78621,I78624,I78627,I78630,I78633,I78636,I78639,I78685,I78688,I78691,I78694,I78697,I78700,I78703,I78706,I78709,I78755,I78758,I78761,I78764,I78767,I78770,I78773,I78776,I78779,I78782,I78828,I78831,I78834,I78837,I78840,I78843,I78846,I78849,I78852,I78898,I78901,I78904,I78907,I78910,I78913,I78916,I78919,I78922,I78968,I78971,I78974,I78977,I78980,I78983,I78986,I78989,I78992,I79038,I79041,I79044,I79047,I79050,I79053,I79056,I79059,I79062,I79108,I79111,I79114,I79117,I79120,I79123,I79126,I79129,I79132,I79135,I79181,I79184,I79187,I79190,I79193,I79196,I79199,I79202,I79205,I79208,I79254,I79257,I79260,I79263,I79266,I79269,I79272,I79275,I79278,I79324,I79327,I79330,I79333,I79336,I79339,I79342,I79345,I79348,I79394,I79397,I79400,I79403,I79406,I79409,I79412,I79415,I79418,I79421,I79467,I79470,I79473,I79476,I79479,I79482,I79485,I79488,I79491,I79537,I79540,I79543,I79546,I79549,I79552,I79555,I79558,I79561,I79607,I79610,I79613,I79616,I79619,I79622,I79625,I79628,I79631,I79677,I79680,I79683,I79686,I79689,I79692,I79695,I79698,I79744,I79747,I79750,I79753,I79756,I79759,I79762,I79765,I79768,I79771,I79817,I79820,I79823,I79826,I79829,I79832,I79835,I79838,I79841,I79887,I79890,I79893,I79896,I79899,I79902,I79905,I79908,I79911,I79914,I79960,I79963,I79966,I79969,I79972,I79975,I79978,I79981,I79984,I79987,I80033,I80036,I80039,I80042,I80045,I80048,I80051,I80054,I80057,I80103,I80106,I80109,I80112,I80115,I80118,I80121,I80124,I80127,I80130,I80176,I80179,I80182,I80185,I80188,I80191,I80194,I80197,I80200,I80246,I80249,I80252,I80255,I80258,I80261,I80264,I80267,I80270,I80273,I80319,I80322,I80325,I80328,I80331,I80334,I80337,I80340,I80343,I80346,I80392,I80395,I80398,I80401,I80404,I80407,I80410,I80413,I80416,I80462,I80465,I80468,I80471,I80474,I80477,I80480,I80483,I80486,I80489,I80535,I80538,I80541,I80544,I80547,I80550,I80553,I80556,I80559,I80605,I80608,I80611,I80614,I80617,I80620,I80623,I80626,I80629,I80675,I80678,I80681,I80684,I80687,I80690,I80693,I80696,I80699,I80702,I80748,I80751,I80754,I80757,I80760,I80763,I80766,I80769,I80815,I80818,I80821,I80824,I80827,I80830,I80833,I80836,I80839,I80885,I80888,I80891,I80894,I80897,I80900,I80903,I80906,I80909,I80912,I80958,I80961,I80964,I80967,I80970,I80973,I80976,I80979,I80982,I80985,I81031,I81034,I81037,I81040,I81043,I81046,I81049,I81052,I81055,I81171,I81174,I81177,I81180,I81183,I81186,I81189,I81192,I81195,I81241,I81244,I81247,I81250,I81253,I81256,I81259,I81262,I81265,I81268,I81314,I81317,I81320,I81323,I81326,I81329,I81332,I81335,I81338,I81341,I81387,I81390,I81393,I81396,I81399,I81402,I81405,I81408,I81454,I81457,I81460,I81463,I81466,I81469,I81472,I81475,I81478,I81524,I81527,I81530,I81533,I81536,I81539,I81542,I81545,I81548,I81594,I81597,I81600,I81603,I81606,I81609,I81612,I81615,I81618,I81621,I81667,I81670,I81673,I81676,I81679,I81682,I81685,I81688,I81691,I81737,I81740,I81743,I81746,I81749,I81752,I81755,I81758,I81761,I81764,I81810,I81813,I81816,I81819,I81822,I81825,I81828,I81831,I81834,I81880,I81883,I81886,I81889,I81892,I81895,I81898,I81901,I81904,I81950,I81953,I81956,I81959,I81962,I81965,I81968,I81971,I81974,I81977,I82023,I82026,I82029,I82032,I82035,I82038,I82041,I82044,I82047,I82093,I82096,I82099,I82102,I82105,I82108,I82111,I82114,I82160,I82163,I82166,I82169,I82172,I82175,I82178,I82181,I82184,I82230,I82233,I82236,I82239,I82242,I82245,I82248,I82251,I82254,I82300,I82303,I82306,I82309,I82312,I82315,I82318,I82321,I82324,I82370,I82373,I82376,I82379,I82382,I82385,I82388,I82391,I82394,I82440,I82443,I82446,I82449,I82452,I82455,I82458,I82461,I82464,I82510,I82513,I82516,I82519,I82522,I82525,I82528,I82531,I82534,I82580,I82583,I82586,I82589,I82592,I82595,I82598,I82601,I82604,I82650,I82653,I82656,I82659,I82662,I82665,I82668,I82671,I82674,I82720,I82723,I82726,I82729,I82732,I82735,I82738,I82741,I82744,I82790,I82793,I82796,I82799,I82802,I82805,I82808,I82811,I82814,I82860,I82863,I82866,I82869,I82872,I82875,I82878,I82881,I82884,I82887,I82933,I82936,I82939,I82942,I82945,I82948,I82951,I82954,I82957,I83003,I83006,I83009,I83012,I83015,I83018,I83021,I83024,I83027,I83073,I83076,I83079,I83082,I83085,I83088,I83091,I83094,I83097,I83100,I83146,I83149,I83152,I83155,I83158,I83161,I83164,I83167,I83170,I83173,I83219,I83222,I83225,I83228,I83231,I83234,I83237,I83240,I83243,I83289,I83292,I83295,I83298,I83301,I83304,I83307,I83310,I83313,I83359,I83362,I83365,I83368,I83371,I83374,I83377,I83380,I83383,I83429,I83432,I83435,I83438,I83441,I83444,I83447,I83450,I83496,I83499,I83502,I83505,I83508,I83511,I83514,I83517,I83520,I83566,I83569,I83572,I83575,I83578,I83581,I83584,I83587,I83590,I83636,I83639,I83642,I83645,I83648,I83651,I83654,I83657,I83703,I83706,I83709,I83712,I83715,I83718,I83721,I83724,I83727,I83730,I83776,I83779,I83782,I83785,I83788,I83791,I83794,I83797,I83800,I83846,I83849,I83852,I83855,I83858,I83861,I83864,I83867,I83870,I83916,I83919,I83922,I83925,I83928,I83931,I83934,I83937,I83940,I83986,I83989,I83992,I83995,I83998,I84001,I84004,I84007,I84010,I84013,I84059,I84062,I84065,I84068,I84071,I84074,I84077,I84080,I84083,I84129,I84132,I84135,I84138,I84141,I84144,I84147,I84150,I84153,I84199,I84202,I84205,I84208,I84211,I84214,I84217,I84220,I84223,I84269,I84272,I84275,I84278,I84281,I84284,I84287,I84290,I84293,I84339,I84342,I84345,I84348,I84351,I84354,I84357,I84360,I84363,I84409,I84412,I84415,I84418,I84421,I84424,I84427,I84430,I84433,I84479,I84482,I84485,I84488,I84491,I84494,I84497,I84500,I84546,I84549,I84552,I84555,I84558,I84561,I84564,I84567,I84570,I84616,I84619,I84622,I84625,I84628,I84631,I84634,I84637,I84683,I84686,I84689,I84692,I84695,I84698,I84701,I84704,I84707,I84753,I84756,I84759,I84762,I84765,I84768,I84771,I84774,I84777,I84780,I84826,I84829,I84832,I84835,I84838,I84841,I84844,I84847,I84850,I84896,I84899,I84902,I84905,I84908,I84911,I84914,I84917,I84920,I84966,I84969,I84972,I84975,I84978,I84981,I84984,I84987,I84990,I84993,I85039,I85042,I85045,I85048,I85051,I85054,I85057,I85060,I85063,I85109,I85112,I85115,I85118,I85121,I85124,I85127,I85130,I85133,I85179,I85182,I85185,I85188,I85191,I85194,I85197,I85200,I85203,I85249,I85252,I85255,I85258,I85261,I85264,I85267,I85270,I85273,I85319,I85322,I85325,I85328,I85331,I85334,I85337,I85340,I85343,I85346,I85392,I85395,I85398,I85401,I85404,I85407,I85410,I85413,I85416,I85419,I85465,I85468,I85471,I85474,I85477,I85480,I85483,I85486,I85489,I85535,I85538,I85541,I85544,I85547,I85550,I85553,I85556,I85559,I85605,I85608,I85611,I85614,I85617,I85620,I85623,I85626,I85629,I85675,I85678,I85681,I85684,I85687,I85690,I85693,I85696,I85699,I85702,I85748,I85751,I85754,I85757,I85760,I85763,I85766,I85769,I85772,I85818,I85821,I85824,I85827,I85830,I85833,I85836,I85839,I85842,I85888,I85891,I85894,I85897,I85900,I85903,I85906,I85909,I85912,I85958,I85961,I85964,I85967,I85970,I85973,I85976,I85979,I85982,I85985,I86031,I86034,I86037,I86040,I86043,I86046,I86049,I86052,I86055,I86101,I86104,I86107,I86110,I86113,I86116,I86119,I86122,I86125,I86171,I86174,I86177,I86180,I86183,I86186,I86189,I86192,I86238,I86241,I86244,I86247,I86250,I86253,I86256,I86259,I86262,I86308,I86311,I86314,I86317,I86320,I86323,I86326,I86329,I86332,I86378,I86381,I86384,I86387,I86390,I86393,I86396,I86399,I86402,I86448,I86451,I86454,I86457,I86460,I86463,I86466,I86469,I86472,I86518,I86521,I86524,I86527,I86530,I86533,I86536,I86539,I86585,I86588,I86591,I86594,I86597,I86600,I86603,I86606,I86609,I86655,I86658,I86661,I86664,I86667,I86670,I86673,I86676,I86722,I86725,I86728,I86731,I86734,I86737,I86740,I86743,I86746,I86792,I86795,I86798,I86801,I86804,I86807,I86810,I86813,I86859,I86862,I86865,I86868,I86871,I86874,I86877,I86880,I86883,I86886,I86932,I86935,I86938,I86941,I86944,I86947,I86950,I86953,I86956,I86959,I87005,I87008,I87011,I87014,I87017,I87020,I87023,I87026,I87072,I87075,I87078,I87081,I87084,I87087,I87090,I87093,I87096,I87142,I87145,I87148,I87151,I87154,I87157,I87160,I87163,I87166,I87212,I87215,I87218,I87221,I87224,I87227,I87230,I87233,I87236,I87239,I87285,I87288,I87291,I87294,I87297,I87300,I87303,I87306,I87309,I87355,I87358,I87361,I87364,I87367,I87370,I87373,I87376,I87379,I87425,I87428,I87431,I87434,I87437,I87440,I87443,I87446,I87449,I87495,I87498,I87501,I87504,I87507,I87510,I87513,I87516,I87519,I87522,I87568,I87571,I87574,I87577,I87580,I87583,I87586,I87589,I87635,I87638,I87641,I87644,I87647,I87650,I87653,I87656,I87659,I87705,I87708,I87711,I87714,I87717,I87720,I87723,I87726,I87729,I87732,I87778,I87781,I87784,I87787,I87790,I87793,I87796,I87799,I87802,I87805,I87851,I87854,I87857,I87860,I87863,I87866,I87869,I87872,I87875,I87921,I87924,I87927,I87930,I87933,I87936,I87939,I87942,I87945,I87948,I87994,I87997,I88000,I88003,I88006,I88009,I88012,I88015,I88018,I88021,I88067,I88070,I88073,I88076,I88079,I88082,I88085,I88088,I88134,I88137,I88140,I88143,I88146,I88149,I88152,I88155,I88158,I88204,I88207,I88210,I88213,I88216,I88219,I88222,I88225,I88228,I88274,I88277,I88280,I88283,I88286,I88289,I88292,I88295,I88298,I88344,I88347,I88350,I88353,I88356,I88359,I88362,I88365,I88368,I88371,I88417,I88420,I88423,I88426,I88429,I88432,I88435,I88438,I88441,I88487,I88490,I88493,I88496,I88499,I88502,I88505,I88508,I88511,I88557,I88560,I88563,I88566,I88569,I88572,I88575,I88578,I88581,I88584,I88630,I88633,I88636,I88639,I88642,I88645,I88648,I88651,I88654,I88700,I88703,I88706,I88709,I88712,I88715,I88718,I88721,I88724,I88770,I88773,I88776,I88779,I88782,I88785,I88788,I88791,I88794,I88840,I88843,I88846,I88849,I88852,I88855,I88858,I88861,I88864,I88867,I88913,I88916,I88919,I88922,I88925,I88928,I88931,I88934,I88937,I88940,I88986,I88989,I88992,I88995,I88998,I89001,I89004,I89007,I89010,I89056,I89059,I89062,I89065,I89068,I89071,I89074,I89077,I89080,I89126,I89129,I89132,I89135,I89138,I89141,I89144,I89147,I89150,I89196,I89199,I89202,I89205,I89208,I89211,I89214,I89217,I89220,I89266,I89269,I89272,I89275,I89278,I89281,I89284,I89287,I89290,I89336,I89339,I89342,I89345,I89348,I89351,I89354,I89357,I89360,I89363,I89409,I89412,I89415,I89418,I89421,I89424,I89427,I89430,I89433,I89479,I89482,I89485,I89488,I89491,I89494,I89497,I89500,I89503,I89506,I89552,I89555,I89558,I89561,I89564,I89567,I89570,I89573,I89576,I89622,I89625,I89628,I89631,I89634,I89637,I89640,I89643,I89646,I89692,I89695,I89698,I89701,I89704,I89707,I89710,I89713,I89716,I89762,I89765,I89768,I89771,I89774,I89777,I89780,I89783,I89786,I89789,I89835,I89838,I89841,I89844,I89847,I89850,I89853,I89856,I89859,I89905,I89908,I89911,I89914,I89917,I89920,I89923,I89926,I89929,I89975,I89978,I89981,I89984,I89987,I89990,I89993,I89996,I89999,I90045,I90048,I90051,I90054,I90057,I90060,I90063,I90066,I90112,I90115,I90118,I90121,I90124,I90127,I90130,I90133,I90136,I90182,I90185,I90188,I90191,I90194,I90197,I90200,I90203,I90206,I90209,I90255,I90258,I90261,I90264,I90267,I90270,I90273,I90276,I90279,I90325,I90328,I90331,I90334,I90337,I90340,I90343,I90346,I90349,I90352,I90398,I90401,I90404,I90407,I90410,I90413,I90416,I90419,I90422,I90468,I90471,I90474,I90477,I90480,I90483,I90486,I90489,I90492,I90538,I90541,I90544,I90547,I90550,I90553,I90556,I90559,I90562,I90608,I90611,I90614,I90617,I90620,I90623,I90626,I90629,I90632,I90678,I90681,I90684,I90687,I90690,I90693,I90696,I90699,I90702,I90705,I90751,I90754,I90757,I90760,I90763,I90766,I90769,I90772,I90775,I90778,I90824,I90827,I90830,I90833,I90836,I90839,I90842,I90845,I90848,I90851,I90897,I90900,I90903,I90906,I90909,I90912,I90915,I90918,I90921,I90967,I90970,I90973,I90976,I90979,I90982,I90985,I90988,I90991,I90994,I91040,I91043,I91046,I91049,I91052,I91055,I91058,I91061,I91107,I91110,I91113,I91116,I91119,I91122,I91125,I91128,I91131,I91177,I91180,I91183,I91186,I91189,I91192,I91195,I91198,I91201,I91247,I91250,I91253,I91256,I91259,I91262,I91265,I91268,I91271,I91274,I91320,I91323,I91326,I91329,I91332,I91335,I91338,I91341,I91344,I91390,I91393,I91396,I91399,I91402,I91405,I91408,I91411,I91414,I91460,I91463,I91466,I91469,I91472,I91475,I91478,I91481,I91527,I91530,I91533,I91536,I91539,I91542,I91545,I91548,I91551,I91554,I91600,I91603,I91606,I91609,I91612,I91615,I91618,I91621,I91624,I91670,I91673,I91676,I91679,I91682,I91685,I91688,I91691,I91694,I91697,I91743,I91746,I91749,I91752,I91755,I91758,I91761,I91764,I91767,I91813,I91816,I91819,I91822,I91825,I91828,I91831,I91834,I91837,I91883,I91886,I91889,I91892,I91895,I91898,I91901,I91904,I91907,I91910,I91956,I91959,I91962,I91965,I91968,I91971,I91974,I91977,I91980,I92026,I92029,I92032,I92035,I92038,I92041,I92044,I92047,I92050,I92053,I92099,I92102,I92105,I92108,I92111,I92114,I92117,I92120,I92123,I92169,I92172,I92175,I92178,I92181,I92184,I92187,I92190,I92193,I92239,I92242,I92245,I92248,I92251,I92254,I92257,I92260,I92263,I92309,I92312,I92315,I92318,I92321,I92324,I92327,I92330,I92333,I92336,I92382,I92385,I92388,I92391,I92394,I92397,I92400,I92403,I92406,I92452,I92455,I92458,I92461,I92464,I92467,I92470,I92473,I92519,I92522,I92525,I92528,I92531,I92534,I92537,I92540,I92543,I92589,I92592,I92595,I92598,I92601,I92604,I92607,I92610,I92613,I92616,I92662,I92665,I92668,I92671,I92674,I92677,I92680,I92683,I92686,I92689,I92735,I92738,I92741,I92744,I92747,I92750,I92753,I92756,I92759,I92805,I92808,I92811,I92814,I92817,I92820,I92823,I92826,I92829,I92832,I92878,I92881,I92884,I92887,I92890,I92893,I92896,I92899,I92902,I92948,I92951,I92954,I92957,I92960,I92963,I92966,I92969,I93015,I93018,I93021,I93024,I93027,I93030,I93033,I93036,I93039,I93042,I93088,I93091,I93094,I93097,I93100,I93103,I93106,I93109,I93112,I93115,I93161,I93164,I93167,I93170,I93173,I93176,I93179,I93182,I93185,I93231,I93234,I93237,I93240,I93243,I93246,I93249,I93252,I93255,I93258,I93304,I93307,I93310,I93313,I93316,I93319,I93322,I93325,I93328,I93374,I93377,I93380,I93383,I93386,I93389,I93392,I93395,I93398,I93444,I93447,I93450,I93453,I93456,I93459,I93462,I93465,I93468,I93514,I93517,I93520,I93523,I93526,I93529,I93532,I93535,I93538,I93584,I93587,I93590,I93593,I93596,I93599,I93602,I93605,I93651,I93654,I93657,I93660,I93663,I93666,I93669,I93672,I93718,I93721,I93724,I93727,I93730,I93733,I93736,I93739,I93742,I93788,I93791,I93794,I93797,I93800,I93803,I93806,I93809,I93812,I93858,I93861,I93864,I93867,I93870,I93873,I93876,I93879,I93882,I93928,I93931,I93934,I93937,I93940,I93943,I93946,I93949,I93952,I93955,I94001,I94004,I94007,I94010,I94013,I94016,I94019,I94022,I94025,I94028,I94074,I94077,I94080,I94083,I94086,I94089,I94092,I94095,I94098,I94101,I94147,I94150,I94153,I94156,I94159,I94162,I94165,I94168,I94214,I94217,I94220,I94223,I94226,I94229,I94232,I94235,I94238,I94284,I94287,I94290,I94293,I94296,I94299,I94302,I94305,I94308,I94354,I94357,I94360,I94363,I94366,I94369,I94372,I94375,I94378,I94381,I94427,I94430,I94433,I94436,I94439,I94442,I94445,I94448,I94451,I94454,I94500,I94503,I94506,I94509,I94512,I94515,I94518,I94521,I94524,I94527,I94573,I94576,I94579,I94582,I94585,I94588,I94591,I94594,I94597,I94643,I94646,I94649,I94652,I94655,I94658,I94661,I94664,I94667,I94713,I94716,I94719,I94722,I94725,I94728,I94731,I94734,I94737,I94783,I94786,I94789,I94792,I94795,I94798,I94801,I94804,I94850,I94853,I94856,I94859,I94862,I94865,I94868,I94871,I94874,I94920,I94923,I94926,I94929,I94932,I94935,I94938,I94941,I94944,I94947,I94993,I94996,I94999,I95002,I95005,I95008,I95011,I95014,I95017,I95063,I95066,I95069,I95072,I95075,I95078,I95081,I95084,I95087,I95090,I95136,I95139,I95142,I95145,I95148,I95151,I95154,I95157,I95160,I95206,I95209,I95212,I95215,I95218,I95221,I95224,I95227,I95230,I95276,I95279,I95282,I95285,I95288,I95291,I95294,I95297,I95343,I95346,I95349,I95352,I95355,I95358,I95361,I95364,I95367,I95413,I95416,I95419,I95422,I95425,I95428,I95431,I95434,I95437,I95483,I95486,I95489,I95492,I95495,I95498,I95501,I95504,I95507,I95553,I95556,I95559,I95562,I95565,I95568,I95571,I95574,I95577,I95580,I95626,I95629,I95632,I95635,I95638,I95641,I95644,I95647,I95650,I95696,I95699,I95702,I95705,I95708,I95711,I95714,I95717,I95763,I95766,I95769,I95772,I95775,I95778,I95781,I95784,I95787,I95833,I95836,I95839,I95842,I95845,I95848,I95851,I95854,I95857,I95860,I95906,I95909,I95912,I95915,I95918,I95921,I95924,I95927,I95973,I95976,I95979,I95982,I95985,I95988,I95991,I95994,I95997,I96043,I96046,I96049,I96052,I96055,I96058,I96061,I96064,I96067,I96113,I96116,I96119,I96122,I96125,I96128,I96131,I96134,I96137,I96183,I96186,I96189,I96192,I96195,I96198,I96201,I96204,I96207,I96253,I96256,I96259,I96262,I96265,I96268,I96271,I96274,I96277,I96280,I96326,I96329,I96332,I96335,I96338,I96341,I96344,I96347,I96350,I96396,I96399,I96402,I96405,I96408,I96411,I96414,I96417,I96463,I96466,I96469,I96472,I96475,I96478,I96481,I96484,I96487,I96533,I96536,I96539,I96542,I96545,I96548,I96551,I96554,I96557,I96560,I96606,I96609,I96612,I96615,I96618,I96621,I96624,I96627,I96630,I96633,I96679,I96682,I96685,I96688,I96691,I96694,I96697,I96700,I96703,I96706,I96752,I96755,I96758,I96761,I96764,I96767,I96770,I96773,I96776,I96822,I96825,I96828,I96831,I96834,I96837,I96840,I96843,I96846,I96892,I96895,I96898,I96901,I96904,I96907,I96910,I96913,I96916,I96962,I96965,I96968,I96971,I96974,I96977,I96980,I96983,I96986,I97032,I97035,I97038,I97041,I97044,I97047,I97050,I97053,I97056,I97102,I97105,I97108,I97111,I97114,I97117,I97120,I97123,I97126,I97172,I97175,I97178,I97181,I97184,I97187,I97190,I97193,I97196,I97242,I97245,I97248,I97251,I97254,I97257,I97260,I97263,I97266,I97312,I97315,I97318,I97321,I97324,I97327,I97330,I97333,I97336,I97382,I97385,I97388,I97391,I97394,I97397,I97400,I97403,I97406,I97409,I97455,I97458,I97461,I97464,I97467,I97470,I97473,I97476,I97479,I97482,I97528,I97531,I97534,I97537,I97540,I97543,I97546,I97549,I97552,I97555,I97601,I97604,I97607,I97610,I97613,I97616,I97619,I97622,I97625,I97628,I97674,I97677,I97680,I97683,I97686,I97689,I97692,I97695,I97698,I97744,I97747,I97750,I97753,I97756,I97759,I97762,I97765,I97768,I97814,I97817,I97820,I97823,I97826,I97829,I97832,I97835,I97838,I97884,I97887,I97890,I97893,I97896,I97899,I97902,I97905,I97908,I97954,I97957,I97960,I97963,I97966,I97969,I97972,I97975,I98021,I98024,I98027,I98030,I98033,I98036,I98039,I98042,I98045,I98091,I98094,I98097,I98100,I98103,I98106,I98109,I98112,I98115,I98118,I98164,I98167,I98170,I98173,I98176,I98179,I98182,I98185,I98188,I98234,I98237,I98240,I98243,I98246,I98249,I98252,I98255,I98258,I98304,I98307,I98310,I98313,I98316,I98319,I98322,I98325,I98328,I98374,I98377,I98380,I98383,I98386,I98389,I98392,I98395,I98441,I98444,I98447,I98450,I98453,I98456,I98459,I98462,I98465,I98511,I98514,I98517,I98520,I98523,I98526,I98529,I98532,I98535,I98538,I98584,I98587,I98590,I98593,I98596,I98599,I98602,I98605,I98608,I98654,I98657,I98660,I98663,I98666,I98669,I98672,I98675,I98678,I98681,I98727,I98730,I98733,I98736,I98739,I98742,I98745,I98748,I98751,I98754,I98800,I98803,I98806,I98809,I98812,I98815,I98818,I98821,I98824,I98870,I98873,I98876,I98879,I98882,I98885,I98888,I98891,I98894,I98897,I98943,I98946,I98949,I98952,I98955,I98958,I98961,I98964,I98967,I98970,I99016,I99019,I99022,I99025,I99028,I99031,I99034,I99037,I99083,I99086,I99089,I99092,I99095,I99098,I99101,I99104,I99107,I99153,I99156,I99159,I99162,I99165,I99168,I99171,I99174,I99177,I99223,I99226,I99229,I99232,I99235,I99238,I99241,I99244,I99247,I99293,I99296,I99299,I99302,I99305,I99308,I99311,I99314,I99317,I99320,I99366,I99369,I99372,I99375,I99378,I99381,I99384,I99387,I99433,I99436,I99439,I99442,I99445,I99448,I99451,I99454,I99457,I99503,I99506,I99509,I99512,I99515,I99518,I99521,I99524,I99527,I99573,I99576,I99579,I99582,I99585,I99588,I99591,I99594,I99597,I99600,I99646,I99649,I99652,I99655,I99658,I99661,I99664,I99667,I99713,I99716,I99719,I99722,I99725,I99728,I99731,I99734,I99737,I99783,I99786,I99789,I99792,I99795,I99798,I99801,I99804,I99807,I99853,I99856,I99859,I99862,I99865,I99868,I99871,I99874,I99877,I99923,I99926,I99929,I99932,I99935,I99938,I99941,I99944,I99947,I99950,I99996,I99999,I100002,I100005,I100008,I100011,I100014,I100017,I100020,I100066,I100069,I100072,I100075,I100078,I100081,I100084,I100087,I100090,I100093,I100139,I100142,I100145,I100148,I100151,I100154,I100157,I100160,I100163,I100166,I100212,I100215,I100218,I100221,I100224,I100227,I100230,I100233,I100236,I100282,I100285,I100288,I100291,I100294,I100297,I100300,I100303,I100306,I100352,I100355,I100358,I100361,I100364,I100367,I100370,I100373,I100376,I100422,I100425,I100428,I100431,I100434,I100437,I100440,I100443,I100446,I100449,I100495,I100498,I100501,I100504,I100507,I100510,I100513,I100516,I100519,I100522,I100568,I100571,I100574,I100577,I100580,I100583,I100586,I100589,I100592,I100638,I100641,I100644,I100647,I100650,I100653,I100656,I100659,I100662,I100708,I100711,I100714,I100717,I100720,I100723,I100726,I100729,I100732,I100845,I100848,I100851,I100854,I100857,I100860,I100863,I100866,I100912,I100915,I100918,I100921,I100924,I100927,I100930,I100933,I100936,I100982,I100985,I100988,I100991,I100994,I100997,I101000,I101003,I101006,I101009,I101055,I101058,I101061,I101064,I101067,I101070,I101073,I101076,I101079,I101125,I101128,I101131,I101134,I101137,I101140,I101143,I101146,I101149,I101195,I101198,I101201,I101204,I101207,I101210,I101213,I101216,I101219,I101265,I101268,I101271,I101274,I101277,I101280,I101283,I101286,I101289,I101292,I101338,I101341,I101344,I101347,I101350,I101353,I101356,I101359,I101362,I101408,I101411,I101414,I101417,I101420,I101423,I101426,I101429,I101432,I101478,I101481,I101484,I101487,I101490,I101493,I101496,I101499,I101502,I101505,I101551,I101554,I101557,I101560,I101563,I101566,I101569,I101572,I101575,I101578,I101624,I101627,I101630,I101633,I101636,I101639,I101642,I101645,I101648,I101694,I101697,I101700,I101703,I101706,I101709,I101712,I101715,I101718,I101764,I101767,I101770,I101773,I101776,I101779,I101782,I101785,I101788,I101791,I101837,I101840,I101843,I101846,I101849,I101852,I101855,I101858,I101861,I101907,I101910,I101913,I101916,I101919,I101922,I101925,I101928,I101931,I101977,I101980,I101983,I101986,I101989,I101992,I101995,I101998,I102001,I102047,I102050,I102053,I102056,I102059,I102062,I102065,I102068,I102071,I102074,I102120,I102123,I102126,I102129,I102132,I102135,I102138,I102141,I102144,I102147,I102193,I102196,I102199,I102202,I102205,I102208,I102211,I102214,I102217,I102263,I102266,I102269,I102272,I102275,I102278,I102281,I102284,I102287,I102290,I102336,I102339,I102342,I102345,I102348,I102351,I102354,I102357,I102360,I102363,I102409,I102412,I102415,I102418,I102421,I102424,I102427,I102430,I102433,I102479,I102482,I102485,I102488,I102491,I102494,I102497,I102500,I102503,I102549,I102552,I102555,I102558,I102561,I102564,I102567,I102570,I102573,I102619,I102622,I102625,I102628,I102631,I102634,I102637,I102640,I102643,I102689,I102692,I102695,I102698,I102701,I102704,I102707,I102710,I102713,I102759,I102762,I102765,I102768,I102771,I102774,I102777,I102780,I102783,I102786,I102832,I102835,I102838,I102841,I102844,I102847,I102850,I102853,I102856,I102902,I102905,I102908,I102911,I102914,I102917,I102920,I102923,I102926,I102972,I102975,I102978,I102981,I102984,I102987,I102990,I102993,I102996,I103042,I103045,I103048,I103051,I103054,I103057,I103060,I103063,I103066,I103112,I103115,I103118,I103121,I103124,I103127,I103130,I103133,I103136,I103139,I103185,I103188,I103191,I103194,I103197,I103200,I103203,I103206,I103209,I103255,I103258,I103261,I103264,I103267,I103270,I103273,I103276,I103279,I103325,I103328,I103331,I103334,I103337,I103340,I103343,I103346,I103349,I103352,I103398,I103401,I103404,I103407,I103410,I103413,I103416,I103419,I103422,I103468,I103471,I103474,I103477,I103480,I103483,I103486,I103489,I103492,I103538,I103541,I103544,I103547,I103550,I103553,I103556,I103559,I103562,I103608,I103611,I103614,I103617,I103620,I103623,I103626,I103629,I103632,I103678,I103681,I103684,I103687,I103690,I103693,I103696,I103699,I103745,I103748,I103751,I103754,I103757,I103760,I103763,I103766,I103769,I103815,I103818,I103821,I103824,I103827,I103830,I103833,I103836,I103839,I103885,I103888,I103891,I103894,I103897,I103900,I103903,I103906,I103909,I103912,I103958,I103961,I103964,I103967,I103970,I103973,I103976,I103979,I103982,I104028,I104031,I104034,I104037,I104040,I104043,I104046,I104049,I104052,I104098,I104101,I104104,I104107,I104110,I104113,I104116,I104119,I104122,I104168,I104171,I104174,I104177,I104180,I104183,I104186,I104189,I104192,I104195,I104241,I104244,I104247,I104250,I104253,I104256,I104259,I104262,I104265,I104268,I104314,I104317,I104320,I104323,I104326,I104329,I104332,I104335,I104338,I104384,I104387,I104390,I104393,I104396,I104399,I104402,I104405,I104408,I104454,I104457,I104460,I104463,I104466,I104469,I104472,I104475,I104478,I104524,I104527,I104530,I104533,I104536,I104539,I104542,I104545,I104548,I104594,I104597,I104600,I104603,I104606,I104609,I104612,I104615,I104618,I104664,I104667,I104670,I104673,I104676,I104679,I104682,I104685,I104688,I104734,I104737,I104740,I104743,I104746,I104749,I104752,I104755,I104758,I104761,I104807,I104810,I104813,I104816,I104819,I104822,I104825,I104828,I104831,I104877,I104880,I104883,I104886,I104889,I104892,I104895,I104898,I104901,I104947,I104950,I104953,I104956,I104959,I104962,I104965,I104968,I104971,I105017,I105020,I105023,I105026,I105029,I105032,I105035,I105038,I105084,I105087,I105090,I105093,I105096,I105099,I105102,I105105,I105108,I105154,I105157,I105160,I105163,I105166,I105169,I105172,I105175,I105178,I105224,I105227,I105230,I105233,I105236,I105239,I105242,I105245,I105248,I105294,I105297,I105300,I105303,I105306,I105309,I105312,I105315,I105318,I105364,I105367,I105370,I105373,I105376,I105379,I105382,I105385,I105431,I105434,I105437,I105440,I105443,I105446,I105449,I105452,I105455,I105458,I105504,I105507,I105510,I105513,I105516,I105519,I105522,I105525,I105571,I105574,I105577,I105580,I105583,I105586,I105589,I105592,I105595,I105641,I105644,I105647,I105650,I105653,I105656,I105659,I105662,I105708,I105711,I105714,I105717,I105720,I105723,I105726,I105729,I105732,I105778,I105781,I105784,I105787,I105790,I105793,I105796,I105799,I105802,I105805,I105851,I105854,I105857,I105860,I105863,I105866,I105869,I105872,I105875,I105921,I105924,I105927,I105930,I105933,I105936,I105939,I105942,I105945,I105991,I105994,I105997,I106000,I106003,I106006,I106009,I106012,I106015,I106061,I106064,I106067,I106070,I106073,I106076,I106079,I106082,I106085,I106131,I106134,I106137,I106140,I106143,I106146,I106149,I106152,I106155,I106158,I106204,I106207,I106210,I106213,I106216,I106219,I106222,I106225,I106271,I106274,I106277,I106280,I106283,I106286,I106289,I106292,I106295,I106341,I106344,I106347,I106350,I106353,I106356,I106359,I106362,I106365,I106411,I106414,I106417,I106420,I106423,I106426,I106429,I106432,I106435,I106438,I106484,I106487,I106490,I106493,I106496,I106499,I106502,I106505,I106508,I106554,I106557,I106560,I106563,I106566,I106569,I106572,I106575,I106578,I106624,I106627,I106630,I106633,I106636,I106639,I106642,I106645,I106648,I106651,I106697,I106700,I106703,I106706,I106709,I106712,I106715,I106718,I106721,I106724,I106770,I106773,I106776,I106779,I106782,I106785,I106788,I106791,I106837,I106840,I106843,I106846,I106849,I106852,I106855,I106858,I106861,I106907,I106910,I106913,I106916,I106919,I106922,I106925,I106928,I106931,I106977,I106980,I106983,I106986,I106989,I106992,I106995,I106998,I107001,I107047,I107050,I107053,I107056,I107059,I107062,I107065,I107068,I107071,I107117,I107120,I107123,I107126,I107129,I107132,I107135,I107138,I107141,I107144,I107190,I107193,I107196,I107199,I107202,I107205,I107208,I107211,I107214,I107260,I107263,I107266,I107269,I107272,I107275,I107278,I107281,I107284,I107330,I107333,I107336,I107339,I107342,I107345,I107348,I107351,I107354,I107400,I107403,I107406,I107409,I107412,I107415,I107418,I107421,I107424,I107427,I107473,I107476,I107479,I107482,I107485,I107488,I107491,I107494,I107497,I107543,I107546,I107549,I107552,I107555,I107558,I107561,I107564,I107567,I107613,I107616,I107619,I107622,I107625,I107628,I107631,I107634,I107637,I107640,I107686,I107689,I107692,I107695,I107698,I107701,I107704,I107707,I107710,I107756,I107759,I107762,I107765,I107768,I107771,I107774,I107777,I107780,I107826,I107829,I107832,I107835,I107838,I107841,I107844,I107847,I107850,I107853,I107899,I107902,I107905,I107908,I107911,I107914,I107917,I107920,I107923,I107969,I107972,I107975,I107978,I107981,I107984,I107987,I107990,I108036,I108039,I108042,I108045,I108048,I108051,I108054,I108057,I108060,I108063,I108109,I108112,I108115,I108118,I108121,I108124,I108127,I108130,I108133,I108179,I108182,I108185,I108188,I108191,I108194,I108197,I108200,I108203,I108206,I108252,I108255,I108258,I108261,I108264,I108267,I108270,I108273,I108276,I108322,I108325,I108328,I108331,I108334,I108337,I108340,I108343,I108346,I108392,I108395,I108398,I108401,I108404,I108407,I108410,I108413,I108416,I108419,I108465,I108468,I108471,I108474,I108477,I108480,I108483,I108486,I108489,I108535,I108538,I108541,I108544,I108547,I108550,I108553,I108556,I108559,I108562,I108608,I108611,I108614,I108617,I108620,I108623,I108626,I108629,I108632,I108678,I108681,I108684,I108687,I108690,I108693,I108696,I108699,I108702,I108748,I108751,I108754,I108757,I108760,I108763,I108766,I108769,I108772,I108775,I108821,I108824,I108827,I108830,I108833,I108836,I108839,I108842,I108845,I108848,I108894,I108897,I108900,I108903,I108906,I108909,I108912,I108915,I108918,I108921,I108967,I108970,I108973,I108976,I108979,I108982,I108985,I108988,I108991,I108994,I109040,I109043,I109046,I109049,I109052,I109055,I109058,I109061,I109064,I109110,I109113,I109116,I109119,I109122,I109125,I109128,I109131,I109177,I109180,I109183,I109186,I109189,I109192,I109195,I109198,I109201,I109247,I109250,I109253,I109256,I109259,I109262,I109265,I109268,I109314,I109317,I109320,I109323,I109326,I109329,I109332,I109335,I109338,I109341,I109387,I109390,I109393,I109396,I109399,I109402,I109405,I109408,I109411,I109457,I109460,I109463,I109466,I109469,I109472,I109475,I109478,I109481,I109484,I109530,I109533,I109536,I109539,I109542,I109545,I109548,I109551,I109554,I109557,I109603,I109606,I109609,I109612,I109615,I109618,I109621,I109624,I109627,I109630,I109676,I109679,I109682,I109685,I109688,I109691,I109694,I109697,I109700,I109746,I109749,I109752,I109755,I109758,I109761,I109764,I109767,I109770,I109816,I109819,I109822,I109825,I109828,I109831,I109834,I109837,I109840,I109843,I109889,I109892,I109895,I109898,I109901,I109904,I109907,I109910,I109913,I109916,I109962,I109965,I109968,I109971,I109974,I109977,I109980,I109983,I109986,I110032,I110035,I110038,I110041,I110044,I110047,I110050,I110053,I110056,I110102,I110105,I110108,I110111,I110114,I110117,I110120,I110123,I110126,I110172,I110175,I110178,I110181,I110184,I110187,I110190,I110193,I110196,I110242,I110245,I110248,I110251,I110254,I110257,I110260,I110263,I110266,I110312,I110315,I110318,I110321,I110324,I110327,I110330,I110333,I110336,I110382,I110385,I110388,I110391,I110394,I110397,I110400,I110403,I110406,I110452,I110455,I110458,I110461,I110464,I110467,I110470,I110473,I110476,I110479,I110525,I110528,I110531,I110534,I110537,I110540,I110543,I110546,I110549,I110595,I110598,I110601,I110604,I110607,I110610,I110613,I110616,I110619,I110622,I110668,I110671,I110674,I110677,I110680,I110683,I110686,I110689,I110692,I110738,I110741,I110744,I110747,I110750,I110753,I110756,I110759,I110762,I110808,I110811,I110814,I110817,I110820,I110823,I110826,I110829,I110875,I110878,I110881,I110884,I110887,I110890,I110893,I110896,I110899,I110945,I110948,I110951,I110954,I110957,I110960,I110963,I110966,I111012,I111015,I111018,I111021,I111024,I111027,I111030,I111033,I111036,I111082,I111085,I111088,I111091,I111094,I111097,I111100,I111103,I111149,I111152,I111155,I111158,I111161,I111164,I111167,I111170,I111173,I111219,I111222,I111225,I111228,I111231,I111234,I111237,I111240,I111243,I111289,I111292,I111295,I111298,I111301,I111304,I111307,I111310,I111313,I111359,I111362,I111365,I111368,I111371,I111374,I111377,I111380,I111426,I111429,I111432,I111435,I111438,I111441,I111444,I111447,I111450,I111496,I111499,I111502,I111505,I111508,I111511,I111514,I111517,I111520,I111523,I111569,I111572,I111575,I111578,I111581,I111584,I111587,I111590,I111593,I111639,I111642,I111645,I111648,I111651,I111654,I111657,I111660,I111663,I111709,I111712,I111715,I111718,I111721,I111724,I111727,I111730,I111733,I111736,I111782,I111785,I111788,I111791,I111794,I111797,I111800,I111803,I111806,I111809,I111855,I111858,I111861,I111864,I111867,I111870,I111873,I111876,I111879,I111925,I111928,I111931,I111934,I111937,I111940,I111943,I111946,I111949,I111952,I111998,I112001,I112004,I112007,I112010,I112013,I112016,I112019,I112022,I112068,I112071,I112074,I112077,I112080,I112083,I112086,I112089,I112092,I112138,I112141,I112144,I112147,I112150,I112153,I112156,I112159,I112162,I112165,I112211,I112214,I112217,I112220,I112223,I112226,I112229,I112232,I112235,I112238,I112284,I112287,I112290,I112293,I112296,I112299,I112302,I112305,I112308,I112354,I112357,I112360,I112363,I112366,I112369,I112372,I112375,I112378,I112424,I112427,I112430,I112433,I112436,I112439,I112442,I112445,I112448,I112451,I112497,I112500,I112503,I112506,I112509,I112512,I112515,I112518,I112521,I112567,I112570,I112573,I112576,I112579,I112582,I112585,I112588,I112591,I112594,I112640,I112643,I112646,I112649,I112652,I112655,I112658,I112661,I112664,I112710,I112713,I112716,I112719,I112722,I112725,I112728,I112731,I112734,I112780,I112783,I112786,I112789,I112792,I112795,I112798,I112801,I112804,I112850,I112853,I112856,I112859,I112862,I112865,I112868,I112871,I112874,I112920,I112923,I112926,I112929,I112932,I112935,I112938,I112941,I112944,I112947,I112993,I112996,I112999,I113002,I113005,I113008,I113011,I113014,I113017,I113063,I113066,I113069,I113072,I113075,I113078,I113081,I113084,I113087,I113090,I113136,I113139,I113142,I113145,I113148,I113151,I113154,I113157,I113160,I113206,I113209,I113212,I113215,I113218,I113221,I113224,I113227,I113230,I113276,I113279,I113282,I113285,I113288,I113291,I113294,I113297,I113300,I113303,I113349,I113352,I113355,I113358,I113361,I113364,I113367,I113370,I113416,I113419,I113422,I113425,I113428,I113431,I113434,I113437,I113440,I113486,I113489,I113492,I113495,I113498,I113501,I113504,I113507,I113510,I113513,I113559,I113562,I113565,I113568,I113571,I113574,I113577,I113580,I113583,I113586,I113632,I113635,I113638,I113641,I113644,I113647,I113650,I113653,I113656,I113659,I113705,I113708,I113711,I113714,I113717,I113720,I113723,I113726,I113729,I113775,I113778,I113781,I113784,I113787,I113790,I113793,I113796,I113799,I113845,I113848,I113851,I113854,I113857,I113860,I113863,I113866,I113869,I113872,I113918,I113921,I113924,I113927,I113930,I113933,I113936,I113939,I113942,I113988,I113991,I113994,I113997,I114000,I114003,I114006,I114009,I114012,I114015,I114061,I114064,I114067,I114070,I114073,I114076,I114079,I114082,I114085,I114088,I114134,I114137,I114140,I114143,I114146,I114149,I114152,I114155,I114201,I114204,I114207,I114210,I114213,I114216,I114219,I114222,I114268,I114271,I114274,I114277,I114280,I114283,I114286,I114289,I114292,I114338,I114341,I114344,I114347,I114350,I114353,I114356,I114359,I114362,I114365,I114411,I114414,I114417,I114420,I114423,I114426,I114429,I114432,I114435,I114438,I114484,I114487,I114490,I114493,I114496,I114499,I114502,I114505,I114508,I114511,I114557,I114560,I114563,I114566,I114569,I114572,I114575,I114578,I114581,I114627,I114630,I114633,I114636,I114639,I114642,I114645,I114648,I114651,I114697,I114700,I114703,I114706,I114709,I114712,I114715,I114718,I114721,I114767,I114770,I114773,I114776,I114779,I114782,I114785,I114788,I114834,I114837,I114840,I114843,I114846,I114849,I114852,I114855,I114858,I114904,I114907,I114910,I114913,I114916,I114919,I114922,I114925,I114928,I114974,I114977,I114980,I114983,I114986,I114989,I114992,I114995,I114998,I115044,I115047,I115050,I115053,I115056,I115059,I115062,I115065,I115068,I115071,I115117,I115120,I115123,I115126,I115129,I115132,I115135,I115138,I115141,I115144,I115190,I115193,I115196,I115199,I115202,I115205,I115208,I115211,I115214,I115260,I115263,I115266,I115269,I115272,I115275,I115278,I115281,I115284,I115330,I115333,I115336,I115339,I115342,I115345,I115348,I115351,I115354,I115357,I115403,I115406,I115409,I115412,I115415,I115418,I115421,I115424,I115470,I115473,I115476,I115479,I115482,I115485,I115488,I115491,I115494,I115540,I115543,I115546,I115549,I115552,I115555,I115558,I115561,I115564,I115567,I115613,I115616,I115619,I115622,I115625,I115628,I115631,I115634,I115637,I115683,I115686,I115689,I115692,I115695,I115698,I115701,I115704,I115707,I115710,I115756,I115759,I115762,I115765,I115768,I115771,I115774,I115777,I115780,I115826,I115829,I115832,I115835,I115838,I115841,I115844,I115847,I115850,I115896,I115899,I115902,I115905,I115908,I115911,I115914,I115917,I115920,I115923,I115969,I115972,I115975,I115978,I115981,I115984,I115987,I115990,I115993,I115996,I116042,I116045,I116048,I116051,I116054,I116057,I116060,I116063,I116066,I116112,I116115,I116118,I116121,I116124,I116127,I116130,I116133,I116136,I116182,I116185,I116188,I116191,I116194,I116197,I116200,I116203,I116206,I116252,I116255,I116258,I116261,I116264,I116267,I116270,I116273,I116319,I116322,I116325,I116328,I116331,I116334,I116337,I116340,I116343,I116346,I116392,I116395,I116398,I116401,I116404,I116407,I116410,I116413,I116416,I116419,I116465,I116468,I116471,I116474,I116477,I116480,I116483,I116486,I116489,I116535,I116538,I116541,I116544,I116547,I116550,I116553,I116556,I116559,I116605,I116608,I116611,I116614,I116617,I116620,I116623,I116626,I116629,I116675,I116678,I116681,I116684,I116687,I116690,I116693,I116696,I116699,I116745,I116748,I116751,I116754,I116757,I116760,I116763,I116766,I116769,I116815,I116818,I116821,I116824,I116827,I116830,I116833,I116836,I116839,I116885,I116888,I116891,I116894,I116897,I116900,I116903,I116906,I116909,I116955,I116958,I116961,I116964,I116967,I116970,I116973,I116976,I116979,I116982,I117028,I117031,I117034,I117037,I117040,I117043,I117046,I117049,I117052,I117098,I117101,I117104,I117107,I117110,I117113,I117116,I117119,I117122,I117125,I117171,I117174,I117177,I117180,I117183,I117186,I117189,I117192,I117195,I117241,I117244,I117247,I117250,I117253,I117256,I117259,I117262,I117308,I117311,I117314,I117317,I117320,I117323,I117326,I117329,I117332,I117335,I117381,I117384,I117387,I117390,I117393,I117396,I117399,I117402,I117448,I117451,I117454,I117457,I117460,I117463,I117466,I117469,I117472,I117518,I117521,I117524,I117527,I117530,I117533,I117536,I117539,I117542,I117588,I117591,I117594,I117597,I117600,I117603,I117606,I117609,I117612,I117615,I117661,I117664,I117667,I117670,I117673,I117676,I117679,I117682,I117685,I117688,I117734,I117737,I117740,I117743,I117746,I117749,I117752,I117755,I117758,I117804,I117807,I117810,I117813,I117816,I117819,I117822,I117825,I117828,I117874,I117877,I117880,I117883,I117886,I117889,I117892,I117895,I117898,I117944,I117947,I117950,I117953,I117956,I117959,I117962,I117965,I117968,I117971,I118017,I118020,I118023,I118026,I118029,I118032,I118035,I118038,I118041,I118087,I118090,I118093,I118096,I118099,I118102,I118105,I118108,I118154,I118157,I118160,I118163,I118166,I118169,I118172,I118175,I118178,I118224,I118227,I118230,I118233,I118236,I118239,I118242,I118245,I118248,I118251,I118297,I118300,I118303,I118306,I118309,I118312,I118315,I118318,I118321,I118367,I118370,I118373,I118376,I118379,I118382,I118385,I118388,I118391,I118437,I118440,I118443,I118446,I118449,I118452,I118455,I118458,I118461,I118507,I118510,I118513,I118516,I118519,I118522,I118525,I118528,I118531,I118577,I118580,I118583,I118586,I118589,I118592,I118595,I118598,I118601,I118604,I118650,I118653,I118656,I118659,I118662,I118665,I118668,I118671,I118674,I118720,I118723,I118726,I118729,I118732,I118735,I118738,I118741,I118787,I118790,I118793,I118796,I118799,I118802,I118805,I118808,I118811,I118857,I118860,I118863,I118866,I118869,I118872,I118875,I118878,I118881,I118927,I118930,I118933,I118936,I118939,I118942,I118945,I118948,I118994,I118997,I119000,I119003,I119006,I119009,I119012,I119015,I119018,I119064,I119067,I119070,I119073,I119076,I119079,I119082,I119085,I119088,I119134,I119137,I119140,I119143,I119146,I119149,I119152,I119155,I119158,I119161,I119207,I119210,I119213,I119216,I119219,I119222,I119225,I119228,I119231,I119277,I119280,I119283,I119286,I119289,I119292,I119295,I119298,I119301,I119304,I119350,I119353,I119356,I119359,I119362,I119365,I119368,I119371,I119374,I119420,I119423,I119426,I119429,I119432,I119435,I119438,I119441,I119444,I119490,I119493,I119496,I119499,I119502,I119505,I119508,I119511,I119514,I119560,I119563,I119566,I119569,I119572,I119575,I119578,I119581,I119584,I119630,I119633,I119636,I119639,I119642,I119645,I119648,I119651,I119654,I119657,I119703,I119706,I119709,I119712,I119715,I119718,I119721,I119724,I119727,I119773,I119776,I119779,I119782,I119785,I119788,I119791,I119794,I119797,I119800,I119846,I119849,I119852,I119855,I119858,I119861,I119864,I119867,I119870,I119873,I119919,I119922,I119925,I119928,I119931,I119934,I119937,I119940,I119943,I119946,I119992,I119995,I119998,I120001,I120004,I120007,I120010,I120013,I120016,I120019,I120065,I120068,I120071,I120074,I120077,I120080,I120083,I120086,I120089,I120135,I120138,I120141,I120144,I120147,I120150,I120153,I120156,I120159,I120205,I120208,I120211,I120214,I120217,I120220,I120223,I120226,I120229,I120232,I120278,I120281,I120284,I120287,I120290,I120293,I120296,I120299,I120302,I120305,I120351,I120354,I120357,I120360,I120363,I120366,I120369,I120372,I120375,I120378,I120424,I120427,I120430,I120433,I120436,I120439,I120442,I120445,I120448,I120567,I120570,I120573,I120576,I120579,I120582,I120585,I120588,I120591,I120637,I120640,I120643,I120646,I120649,I120652,I120655,I120658,I120661,I120664,I120710,I120713,I120716,I120719,I120722,I120725,I120728,I120731,I120734,I120737,I120783,I120786,I120789,I120792,I120795,I120798,I120801,I120804,I120807,I120853,I120856,I120859,I120862,I120865,I120868,I120871,I120874,I120877,I120923,I120926,I120929,I120932,I120935,I120938,I120941,I120944,I120947,I120950,I120996,I120999,I121002,I121005,I121008,I121011,I121014,I121017,I121020,I121066,I121069,I121072,I121075,I121078,I121081,I121084,I121087,I121090,I121093,I121139,I121142,I121145,I121148,I121151,I121154,I121157,I121160,I121163,I121209,I121212,I121215,I121218,I121221,I121224,I121227,I121230,I121233,I121236,I121282,I121285,I121288,I121291,I121294,I121297,I121300,I121303,I121306,I121352,I121355,I121358,I121361,I121364,I121367,I121370,I121373,I121376,I121422,I121425,I121428,I121431,I121434,I121437,I121440,I121443,I121446,I121449,I121495,I121498,I121501,I121504,I121507,I121510,I121513,I121516,I121519,I121565,I121568,I121571,I121574,I121577,I121580,I121583,I121586,I121589,I121635,I121638,I121641,I121644,I121647,I121650,I121653,I121656,I121659,I121662,I121708,I121711,I121714,I121717,I121720,I121723,I121726,I121729,I121732,I121735,I121781,I121784,I121787,I121790,I121793,I121796,I121799,I121802,I121805,I121808,I121854,I121857,I121860,I121863,I121866,I121869,I121872,I121875,I121878,I121924,I121927,I121930,I121933,I121936,I121939,I121942,I121945,I121948,I121994,I121997,I122000,I122003,I122006,I122009,I122012,I122015,I122018,I122021,I122067,I122070,I122073,I122076,I122079,I122082,I122085,I122088,I122091,I122094,I122140,I122143,I122146,I122149,I122152,I122155,I122158,I122161,I122164,I122210,I122213,I122216,I122219,I122222,I122225,I122228,I122231,I122277,I122280,I122283,I122286,I122289,I122292,I122295,I122298,I122301,I122304,I122350,I122353,I122356,I122359,I122362,I122365,I122368,I122371,I122374,I122420,I122423,I122426,I122429,I122432,I122435,I122438,I122441,I122444,I122447,I122493,I122496,I122499,I122502,I122505,I122508,I122511,I122514,I122560,I122563,I122566,I122569,I122572,I122575,I122578,I122581,I122584,I122587,I122633,I122636,I122639,I122642,I122645,I122648,I122651,I122654,I122657,I122703,I122706,I122709,I122712,I122715,I122718,I122721,I122724,I122727,I122773,I122776,I122779,I122782,I122785,I122788,I122791,I122794,I122840,I122843,I122846,I122849,I122852,I122855,I122858,I122861,I122864,I122867,I122913,I122916,I122919,I122922,I122925,I122928,I122931,I122934,I122937,I122983,I122986,I122989,I122992,I122995,I122998,I123001,I123004,I123007,I123010,I123056,I123059,I123062,I123065,I123068,I123071,I123074,I123077,I123080,I123083,I123129,I123132,I123135,I123138,I123141,I123144,I123147,I123150,I123196,I123199,I123202,I123205,I123208,I123211,I123214,I123217,I123220,I123266,I123269,I123272,I123275,I123278,I123281,I123284,I123287,I123290,I123293,I123339,I123342,I123345,I123348,I123351,I123354,I123357,I123360,I123363,I123409,I123412,I123415,I123418,I123421,I123424,I123427,I123430,I123433,I123479,I123482,I123485,I123488,I123491,I123494,I123497,I123500,I123503,I123549,I123552,I123555,I123558,I123561,I123564,I123567,I123570,I123573,I123576,I123622,I123625,I123628,I123631,I123634,I123637,I123640,I123643,I123646,I123649,I123695,I123698,I123701,I123704,I123707,I123710,I123713,I123716,I123719,I123765,I123768,I123771,I123774,I123777,I123780,I123783,I123786,I123789,I123792,I123838,I123841,I123844,I123847,I123850,I123853,I123856,I123859,I123862,I123908,I123911,I123914,I123917,I123920,I123923,I123926,I123929,I123932,I123978,I123981,I123984,I123987,I123990,I123993,I123996,I123999,I124002,I124048,I124051,I124054,I124057,I124060,I124063,I124066,I124069,I124072,I124118,I124121,I124124,I124127,I124130,I124133,I124136,I124139,I124142,I124145,I124191,I124194,I124197,I124200,I124203,I124206,I124209,I124212,I124215,I124261,I124264,I124267,I124270,I124273,I124276,I124279,I124282,I124328,I124331,I124334,I124337,I124340,I124343,I124346,I124349,I124352,I124355,I124401,I124404,I124407,I124410,I124413,I124416,I124419,I124422,I124425,I124471,I124474,I124477,I124480,I124483,I124486,I124489,I124492,I124538,I124541,I124544,I124547,I124550,I124553,I124556,I124559,I124562,I124608,I124611,I124614,I124617,I124620,I124623,I124626,I124629,I124632,I124678,I124681,I124684,I124687,I124690,I124693,I124696,I124699,I124702,I124705,I124751,I124754,I124757,I124760,I124763,I124766,I124769,I124772,I124775,I124821,I124824,I124827,I124830,I124833,I124836,I124839,I124842,I124845,I124848,I124894,I124897,I124900,I124903,I124906,I124909,I124912,I124915,I124918,I124921,I124967,I124970,I124973,I124976,I124979,I124982,I124985,I124988,I124991,I125037,I125040,I125043,I125046,I125049,I125052,I125055,I125058,I125104,I125107,I125110,I125113,I125116,I125119,I125122,I125125,I125128,I125174,I125177,I125180,I125183,I125186,I125189,I125192,I125195,I125198,I125244,I125247,I125250,I125253,I125256,I125259,I125262,I125265,I125268,I125271,I125317,I125320,I125323,I125326,I125329,I125332,I125335,I125338,I125341,I125344,I125390,I125393,I125396,I125399,I125402,I125405,I125408,I125411,I125414,I125460,I125463,I125466,I125469,I125472,I125475,I125478,I125481,I125484,I125487,I125533,I125536,I125539,I125542,I125545,I125548,I125551,I125554,I125557,I125603,I125606,I125609,I125612,I125615,I125618,I125621,I125624,I125627,I125673,I125676,I125679,I125682,I125685,I125688,I125691,I125694,I125740,I125743,I125746,I125749,I125752,I125755,I125758,I125761,I125764,I125767,I125813,I125816,I125819,I125822,I125825,I125828,I125831,I125834,I125880,I125883,I125886,I125889,I125892,I125895,I125898,I125901,I125904,I125950,I125953,I125956,I125959,I125962,I125965,I125968,I125971,I125974,I125977,I126023,I126026,I126029,I126032,I126035,I126038,I126041,I126044,I126090,I126093,I126096,I126099,I126102,I126105,I126108,I126111,I126114,I126160,I126163,I126166,I126169,I126172,I126175,I126178,I126181,I126184,I126230,I126233,I126236,I126239,I126242,I126245,I126248,I126251,I126254,I126300,I126303,I126306,I126309,I126312,I126315,I126318,I126321,I126324,I126327,I126373,I126376,I126379,I126382,I126385,I126388,I126391,I126394,I126397,I126400,I126446,I126449,I126452,I126455,I126458,I126461,I126464,I126467,I126470,I126516,I126519,I126522,I126525,I126528,I126531,I126534,I126537,I126540,I126586,I126589,I126592,I126595,I126598,I126601,I126604,I126607,I126610,I126613,I126659,I126662,I126665,I126668,I126671,I126674,I126677,I126680,I126726,I126729,I126732,I126735,I126738,I126741,I126744,I126747,I126750,I126753,I126799,I126802,I126805,I126808,I126811,I126814,I126817,I126820,I126823,I126826,I126872,I126875,I126878,I126881,I126884,I126887,I126890,I126893,I126896,I126899,I126945,I126948,I126951,I126954,I126957,I126960,I126963,I126966,I126969,I126972,I127018,I127021,I127024,I127027,I127030,I127033,I127036,I127039,I127042,I127088,I127091,I127094,I127097,I127100,I127103,I127106,I127109,I127155,I127158,I127161,I127164,I127167,I127170,I127173,I127176,I127179,I127182,I127228,I127231,I127234,I127237,I127240,I127243,I127246,I127249,I127252,I127298,I127301,I127304,I127307,I127310,I127313,I127316,I127319,I127322,I127368,I127371,I127374,I127377,I127380,I127383,I127386,I127389,I127392,I127395,I127441,I127444,I127447,I127450,I127453,I127456,I127459,I127462,I127465,I127511,I127514,I127517,I127520,I127523,I127526,I127529,I127532,I127535,I127581,I127584,I127587,I127590,I127593,I127596,I127599,I127602,I127648,I127651,I127654,I127657,I127660,I127663,I127666,I127669,I127672,I127718,I127721,I127724,I127727,I127730,I127733,I127736,I127739,I127785,I127788,I127791,I127794,I127797,I127800,I127803,I127806,I127809,I127855,I127858,I127861,I127864,I127867,I127870,I127873,I127876,I127879,I127925,I127928,I127931,I127934,I127937,I127940,I127943,I127946,I127949,I127995,I127998,I128001,I128004,I128007,I128010,I128013,I128016,I128019,I128022,I128068,I128071,I128074,I128077,I128080,I128083,I128086,I128089,I128092,I128138,I128141,I128144,I128147,I128150,I128153,I128156,I128159,I128162,I128208,I128211,I128214,I128217,I128220,I128223,I128226,I128229,I128232,I128235,I128281,I128284,I128287,I128290,I128293,I128296,I128299,I128302,I128305,I128351,I128354,I128357,I128360,I128363,I128366,I128369,I128372,I128375,I128421,I128424,I128427,I128430,I128433,I128436,I128439,I128442,I128488,I128491,I128494,I128497,I128500,I128503,I128506,I128509,I128512,I128558,I128561,I128564,I128567,I128570,I128573,I128576,I128579,I128582,I128585,I128631,I128634,I128637,I128640,I128643,I128646,I128649,I128652,I128655,I128701,I128704,I128707,I128710,I128713,I128716,I128719,I128722,I128725,I128771,I128774,I128777,I128780,I128783,I128786,I128789,I128792,I128838,I128841,I128844,I128847,I128850,I128853,I128856,I128859,I128862,I128865,I128911,I128914,I128917,I128920,I128923,I128926,I128929,I128932,I128935,I128981,I128984,I128987,I128990,I128993,I128996,I128999,I129002,I129005,I129008,I129054,I129057,I129060,I129063,I129066,I129069,I129072,I129075,I129078,I129124,I129127,I129130,I129133,I129136,I129139,I129142,I129145,I129148,I129151,I129197,I129200,I129203,I129206,I129209,I129212,I129215,I129218,I129221,I129224,I129270,I129273,I129276,I129279,I129282,I129285,I129288,I129291,I129294,I129340,I129343,I129346,I129349,I129352,I129355,I129358,I129361,I129364,I129367,I129413,I129416,I129419,I129422,I129425,I129428,I129431,I129434,I129437,I129440,I129486,I129489,I129492,I129495,I129498,I129501,I129504,I129507,I129510,I129556,I129559,I129562,I129565,I129568,I129571,I129574,I129577,I129580,I129583,I129629,I129632,I129635,I129638,I129641,I129644,I129647,I129650,I129653,I129656,I129702,I129705,I129708,I129711,I129714,I129717,I129720,I129723,I129726,I129772,I129775,I129778,I129781,I129784,I129787,I129790,I129793,I129796,I129842,I129845,I129848,I129851,I129854,I129857,I129860,I129863,I129909,I129912,I129915,I129918,I129921,I129924,I129927,I129930,I129933,I129979,I129982,I129985,I129988,I129991,I129994,I129997,I130000,I130003,I130049,I130052,I130055,I130058,I130061,I130064,I130067,I130070,I130073,I130119,I130122,I130125,I130128,I130131,I130134,I130137,I130140,I130143,I130146,I130192,I130195,I130198,I130201,I130204,I130207,I130210,I130213,I130216,I130262,I130265,I130268,I130271,I130274,I130277,I130280,I130283,I130286,I130332,I130335,I130338,I130341,I130344,I130347,I130350,I130353,I130356,I130359,I130405,I130408,I130411,I130414,I130417,I130420,I130423,I130426,I130429,I130475,I130478,I130481,I130484,I130487,I130490,I130493,I130496,I130499,I130545,I130548,I130551,I130554,I130557,I130560,I130563,I130566,I130612,I130615,I130618,I130621,I130624,I130627,I130630,I130633,I130636,I130639,I130685,I130688,I130691,I130694,I130697,I130700,I130703,I130706,I130709,I130755,I130758,I130761,I130764,I130767,I130770,I130773,I130776,I130779,I130825,I130828,I130831,I130834,I130837,I130840,I130843,I130846,I130849,I130895,I130898,I130901,I130904,I130907,I130910,I130913,I130916,I130962,I130965,I130968,I130971,I130974,I130977,I130980,I130983,I130986,I130989,I131035,I131038,I131041,I131044,I131047,I131050,I131053,I131056,I131059,I131062,I131108,I131111,I131114,I131117,I131120,I131123,I131126,I131129,I131132,I131178,I131181,I131184,I131187,I131190,I131193,I131196,I131199,I131202,I131205,I131251,I131254,I131257,I131260,I131263,I131266,I131269,I131272,I131275,I131321,I131324,I131327,I131330,I131333,I131336,I131339,I131342,I131345,I131348,I131394,I131397,I131400,I131403,I131406,I131409,I131412,I131415,I131418,I131464,I131467,I131470,I131473,I131476,I131479,I131482,I131485,I131488,I131534,I131537,I131540,I131543,I131546,I131549,I131552,I131555,I131558,I131604,I131607,I131610,I131613,I131616,I131619,I131622,I131625,I131628,I131674,I131677,I131680,I131683,I131686,I131689,I131692,I131695,I131741,I131744,I131747,I131750,I131753,I131756,I131759,I131762,I131765,I131811,I131814,I131817,I131820,I131823,I131826,I131829,I131832,I131878,I131881,I131884,I131887,I131890,I131893,I131896,I131899,I131902,I131948,I131951,I131954,I131957,I131960,I131963,I131966,I131969,I131972,I132018,I132021,I132024,I132027,I132030,I132033,I132036,I132039,I132042,I132045,I132091,I132094,I132097,I132100,I132103,I132106,I132109,I132112,I132115,I132161,I132164,I132167,I132170,I132173,I132176,I132179,I132182,I132185,I132231,I132234,I132237,I132240,I132243,I132246,I132249,I132252,I132255,I132301,I132304,I132307,I132310,I132313,I132316,I132319,I132322,I132325,I132371,I132374,I132377,I132380,I132383,I132386,I132389,I132392,I132395,I132441,I132444,I132447,I132450,I132453,I132456,I132459,I132462,I132465,I132511,I132514,I132517,I132520,I132523,I132526,I132529,I132532,I132535,I132581,I132584,I132587,I132590,I132593,I132596,I132599,I132602,I132648,I132651,I132654,I132657,I132660,I132663,I132666,I132669,I132672,I132718,I132721,I132724,I132727,I132730,I132733,I132736,I132739,I132742,I132745,I132791,I132794,I132797,I132800,I132803,I132806,I132809,I132812,I132815,I132861,I132864,I132867,I132870,I132873,I132876,I132879,I132882,I132885,I132931,I132934,I132937,I132940,I132943,I132946,I132949,I132952,I132955,I132958,I133004,I133007,I133010,I133013,I133016,I133019,I133022,I133025,I133028,I133074,I133077,I133080,I133083,I133086,I133089,I133092,I133095,I133098,I133101,I133147,I133150,I133153,I133156,I133159,I133162,I133165,I133168,I133171,I133174,I133220,I133223,I133226,I133229,I133232,I133235,I133238,I133241,I133244,I133290,I133293,I133296,I133299,I133302,I133305,I133308,I133311,I133314,I133317,I133363,I133366,I133369,I133372,I133375,I133378,I133381,I133384,I133387,I133433,I133436,I133439,I133442,I133445,I133448,I133451,I133454,I133500,I133503,I133506,I133509,I133512,I133515,I133518,I133521,I133524,I133527,I133573,I133576,I133579,I133582,I133585,I133588,I133591,I133594,I133597,I133643,I133646,I133649,I133652,I133655,I133658,I133661,I133664,I133667,I133713,I133716,I133719,I133722,I133725,I133728,I133731,I133734,I133737,I133740,I133786,I133789,I133792,I133795,I133798,I133801,I133804,I133807,I133810,I133813,I133859,I133862,I133865,I133868,I133871,I133874,I133877,I133880,I133883,I133929,I133932,I133935,I133938,I133941,I133944,I133947,I133950,I133953,I133956,I134002,I134005,I134008,I134011,I134014,I134017,I134020,I134023,I134026,I134072,I134075,I134078,I134081,I134084,I134087,I134090,I134093,I134096,I134142,I134145,I134148,I134151,I134154,I134157,I134160,I134163,I134209,I134212,I134215,I134218,I134221,I134224,I134227,I134230,I134233,I134236,I134282,I134285,I134288,I134291,I134294,I134297,I134300,I134303,I134306,I134352,I134355,I134358,I134361,I134364,I134367,I134370,I134373,I134419,I134422,I134425,I134428,I134431,I134434,I134437,I134440,I134443,I134446,I134492,I134495,I134498,I134501,I134504,I134507,I134510,I134513,I134516,I134519,I134565,I134568,I134571,I134574,I134577,I134580,I134583,I134586,I134589,I134635,I134638,I134641,I134644,I134647,I134650,I134653,I134656,I134702,I134705,I134708,I134711,I134714,I134717,I134720,I134723,I134726,I134772,I134775,I134778,I134781,I134784,I134787,I134790,I134793,I134796,I134842,I134845,I134848,I134851,I134854,I134857,I134860,I134863,I134866,I134912,I134915,I134918,I134921,I134924,I134927,I134930,I134933,I134936,I134982,I134985,I134988,I134991,I134994,I134997,I135000,I135003,I135006,I135009,I135055,I135058,I135061,I135064,I135067,I135070,I135073,I135076,I135079,I135125,I135128,I135131,I135134,I135137,I135140,I135143,I135146,I135149,I135152,I135198,I135201,I135204,I135207,I135210,I135213,I135216,I135219,I135222,I135268,I135271,I135274,I135277,I135280,I135283,I135286,I135289,I135292,I135295,I135341,I135344,I135347,I135350,I135353,I135356,I135359,I135362,I135365,I135411,I135414,I135417,I135420,I135423,I135426,I135429,I135432,I135435,I135481,I135484,I135487,I135490,I135493,I135496,I135499,I135502,I135505,I135508,I135554,I135557,I135560,I135563,I135566,I135569,I135572,I135575,I135621,I135624,I135627,I135630,I135633,I135636,I135639,I135642,I135645,I135648,I135694,I135697,I135700,I135703,I135706,I135709,I135712,I135715,I135718,I135721,I135767,I135770,I135773,I135776,I135779,I135782,I135785,I135788,I135834,I135837,I135840,I135843,I135846,I135849,I135852,I135855,I135858,I135904,I135907,I135910,I135913,I135916,I135919,I135922,I135925,I135971,I135974,I135977,I135980,I135983,I135986,I135989,I135992,I136038,I136041,I136044,I136047,I136050,I136053,I136056,I136059,I136062,I136108,I136111,I136114,I136117,I136120,I136123,I136126,I136129,I136132,I136178,I136181,I136184,I136187,I136190,I136193,I136196,I136199,I136202,I136205,I136251,I136254,I136257,I136260,I136263,I136266,I136269,I136272,I136275,I136321,I136324,I136327,I136330,I136333,I136336,I136339,I136342,I136388,I136391,I136394,I136397,I136400,I136403,I136406,I136409,I136412,I136458,I136461,I136464,I136467,I136470,I136473,I136476,I136479,I136525,I136528,I136531,I136534,I136537,I136540,I136543,I136546,I136592,I136595,I136598,I136601,I136604,I136607,I136610,I136613,I136616,I136619,I136665,I136668,I136671,I136674,I136677,I136680,I136683,I136686,I136689,I136692,I136738,I136741,I136744,I136747,I136750,I136753,I136756,I136759,I136762,I136808,I136811,I136814,I136817,I136820,I136823,I136826,I136829,I136832,I136878,I136881,I136884,I136887,I136890,I136893,I136896,I136899,I136902,I136948,I136951,I136954,I136957,I136960,I136963,I136966,I136969,I137015,I137018,I137021,I137024,I137027,I137030,I137033,I137036,I137082,I137085,I137088,I137091,I137094,I137097,I137100,I137103,I137106,I137109,I137155,I137158,I137161,I137164,I137167,I137170,I137173,I137176,I137179,I137225,I137228,I137231,I137234,I137237,I137240,I137243,I137246,I137249,I137295,I137298,I137301,I137304,I137307,I137310,I137313,I137316,I137362,I137365,I137368,I137371,I137374,I137377,I137380,I137383,I137386,I137432,I137435,I137438,I137441,I137444,I137447,I137450,I137453,I137499,I137502,I137505,I137508,I137511,I137514,I137517,I137520,I137523,I137526,I137572,I137575,I137578,I137581,I137584,I137587,I137590,I137593,I137596,I137642,I137645,I137648,I137651,I137654,I137657,I137660,I137663,I137666,I137669,I137715,I137718,I137721,I137724,I137727,I137730,I137733,I137736,I137739,I137785,I137788,I137791,I137794,I137797,I137800,I137803,I137806,I137809,I137855,I137858,I137861,I137864,I137867,I137870,I137873,I137876,I137922,I137925,I137928,I137931,I137934,I137937,I137940,I137943,I137946,I137949,I137995,I137998,I138001,I138004,I138007,I138010,I138013,I138016,I138019,I138065,I138068,I138071,I138074,I138077,I138080,I138083,I138086,I138089,I138135,I138138,I138141,I138144,I138147,I138150,I138153,I138156,I138159,I138205,I138208,I138211,I138214,I138217,I138220,I138223,I138226,I138229,I138275,I138278,I138281,I138284,I138287,I138290,I138293,I138296,I138299,I138345,I138348,I138351,I138354,I138357,I138360,I138363,I138366,I138412,I138415,I138418,I138421,I138424,I138427,I138430,I138433,I138436,I138439,I138485,I138488,I138491,I138494,I138497,I138500,I138503,I138506,I138552,I138555,I138558,I138561,I138564,I138567,I138570,I138573,I138576,I138579,I138625,I138628,I138631,I138634,I138637,I138640,I138643,I138646,I138649,I138695,I138698,I138701,I138704,I138707,I138710,I138713,I138716,I138719,I138722,I138768,I138771,I138774,I138777,I138780,I138783,I138786,I138789,I138792,I138838,I138841,I138844,I138847,I138850,I138853,I138856,I138859,I138862,I138908,I138911,I138914,I138917,I138920,I138923,I138926,I138929,I138932,I138935,I138981,I138984,I138987,I138990,I138993,I138996,I138999,I139002,I139048,I139051,I139054,I139057,I139060,I139063,I139066,I139069,I139072,I139075,I139121,I139124,I139127,I139130,I139133,I139136,I139139,I139142,I139145,I139191,I139194,I139197,I139200,I139203,I139206,I139209,I139212,I139215,I139261,I139264,I139267,I139270,I139273,I139276,I139279,I139282,I139285,I139331,I139334,I139337,I139340,I139343,I139346,I139349,I139352,I139398,I139401,I139404,I139407,I139410,I139413,I139416,I139419,I139422,I139468,I139471,I139474,I139477,I139480,I139483,I139486,I139489,I139535,I139538,I139541,I139544,I139547,I139550,I139553,I139556,I139559,I139605,I139608,I139611,I139614,I139617,I139620,I139623,I139626,I139629,I139632,I139678,I139681,I139684,I139687,I139690,I139693,I139696,I139699,I139702,I139748,I139751,I139754,I139757,I139760,I139763,I139766,I139769,I139772,I139775,I139821,I139824,I139827,I139830,I139833,I139836,I139839,I139842,I139845,I139891,I139894,I139897,I139900,I139903,I139906,I139909,I139912,I139958,I139961,I139964,I139967,I139970,I139973,I139976,I139979,I139982,I140028,I140031,I140034,I140037,I140040,I140043,I140046,I140049,I140052,I140098,I140101,I140104,I140107,I140110,I140113,I140116,I140119,I140122,I140238,I140241,I140244,I140247,I140250,I140253,I140256,I140259,I140262,I140265,I140311,I140314,I140317,I140320,I140323,I140326,I140329,I140332,I140335,I140381,I140384,I140387,I140390,I140393,I140396,I140399,I140402,I140405,I140408,I140454,I140457,I140460,I140463,I140466,I140469,I140472,I140475,I140478,I140524,I140527,I140530,I140533,I140536,I140539,I140542,I140545,I140591,I140594,I140597,I140600,I140603,I140606,I140609,I140612,I140615,I140618,I140664,I140667,I140670,I140673,I140676,I140679,I140682,I140685,I140688,I140734,I140737,I140740,I140743,I140746,I140749,I140752,I140755,I140801,I140804,I140807,I140810,I140813,I140816,I140819,I140822,I140825,I140871,I140874,I140877,I140880,I140883,I140886,I140889,I140892,I140895,I140941,I140944,I140947,I140950,I140953,I140956,I140959,I140962,I140965,I141011,I141014,I141017,I141020,I141023,I141026,I141029,I141032,I141035,I141081,I141084,I141087,I141090,I141093,I141096,I141099,I141102,I141105,I141108,I141154,I141157,I141160,I141163,I141166,I141169,I141172,I141175,I141178,I141181,I141227,I141230,I141233,I141236,I141239,I141242,I141245,I141248,I141251,I141297,I141300,I141303,I141306,I141309,I141312,I141315,I141318,I141321,I141324,I141370,I141373,I141376,I141379,I141382,I141385,I141388,I141391,I141394,I141397,I141443,I141446,I141449,I141452,I141455,I141458,I141461,I141464,I141467,I141513,I141516,I141519,I141522,I141525,I141528,I141531,I141534,I141537,I141583,I141586,I141589,I141592,I141595,I141598,I141601,I141604,I141607,I141653,I141656,I141659,I141662,I141665,I141668,I141671,I141674,I141677,I141680,I141726,I141729,I141732,I141735,I141738,I141741,I141744,I141747,I141750,I141796,I141799,I141802,I141805,I141808,I141811,I141814,I141817,I141820,I141866,I141869,I141872,I141875,I141878,I141881,I141884,I141887,I141890,I141936,I141939,I141942,I141945,I141948,I141951,I141954,I141957,I141960,I141963,I142009,I142012,I142015,I142018,I142021,I142024,I142027,I142030,I142033,I142079,I142082,I142085,I142088,I142091,I142094,I142097,I142100,I142103,I142106,I142152,I142155,I142158,I142161,I142164,I142167,I142170,I142173,I142176,I142222,I142225,I142228,I142231,I142234,I142237,I142240,I142243,I142246,I142292,I142295,I142298,I142301,I142304,I142307,I142310,I142313,I142316,I142362,I142365,I142368,I142371,I142374,I142377,I142380,I142383,I142429,I142432,I142435,I142438,I142441,I142444,I142447,I142450,I142453,I142456,I142502,I142505,I142508,I142511,I142514,I142517,I142520,I142523,I142569,I142572,I142575,I142578,I142581,I142584,I142587,I142590,I142593,I142639,I142642,I142645,I142648,I142651,I142654,I142657,I142660,I142663,I142666,I142712,I142715,I142718,I142721,I142724,I142727,I142730,I142733,I142736,I142739,I142785,I142788,I142791,I142794,I142797,I142800,I142803,I142806,I142809,I142855,I142858,I142861,I142864,I142867,I142870,I142873,I142876,I142879,I142925,I142928,I142931,I142934,I142937,I142940,I142943,I142946,I142949,I142952,I142998,I143001,I143004,I143007,I143010,I143013,I143016,I143019,I143022,I143068,I143071,I143074,I143077,I143080,I143083,I143086,I143089,I143092,I143138,I143141,I143144,I143147,I143150,I143153,I143156,I143159,I143162,I143165,I143211,I143214,I143217,I143220,I143223,I143226,I143229,I143232,I143235,I143281,I143284,I143287,I143290,I143293,I143296,I143299,I143302,I143305,I143351,I143354,I143357,I143360,I143363,I143366,I143369,I143372,I143375,I143378,I143424,I143427,I143430,I143433,I143436,I143439,I143442,I143445,I143448,I143494,I143497,I143500,I143503,I143506,I143509,I143512,I143515,I143518,I143564,I143567,I143570,I143573,I143576,I143579,I143582,I143585,I143588,I143634,I143637,I143640,I143643,I143646,I143649,I143652,I143655,I143658,I143704,I143707,I143710,I143713,I143716,I143719,I143722,I143725,I143728,I143774,I143777,I143780,I143783,I143786,I143789,I143792,I143795,I143798,I143801,I143847,I143850,I143853,I143856,I143859,I143862,I143865,I143868,I143871,I143917,I143920,I143923,I143926,I143929,I143932,I143935,I143938,I143941,I143987,I143990,I143993,I143996,I143999,I144002,I144005,I144008,I144011,I144014,I144060,I144063,I144066,I144069,I144072,I144075,I144078,I144081,I144084,I144130,I144133,I144136,I144139,I144142,I144145,I144148,I144151,I144154,I144200,I144203,I144206,I144209,I144212,I144215,I144218,I144221,I144224,I144270,I144273,I144276,I144279,I144282,I144285,I144288,I144291,I144294,I144340,I144343,I144346,I144349,I144352,I144355,I144358,I144361,I144364,I144410,I144413,I144416,I144419,I144422,I144425,I144428,I144431,I144434,I144480,I144483,I144486,I144489,I144492,I144495,I144498,I144501,I144504,I144550,I144553,I144556,I144559,I144562,I144565,I144568,I144571,I144574,I144577,I144623,I144626,I144629,I144632,I144635,I144638,I144641,I144644,I144647,I144650,I144696,I144699,I144702,I144705,I144708,I144711,I144714,I144717,I144720,I144766,I144769,I144772,I144775,I144778,I144781,I144784,I144787,I144790,I144836,I144839,I144842,I144845,I144848,I144851,I144854,I144857,I144860,I144863,I144909,I144912,I144915,I144918,I144921,I144924,I144927,I144930,I144933,I144979,I144982,I144985,I144988,I144991,I144994,I144997,I145000,I145046,I145049,I145052,I145055,I145058,I145061,I145064,I145067,I145070,I145116,I145119,I145122,I145125,I145128,I145131,I145134,I145137,I145140,I145186,I145189,I145192,I145195,I145198,I145201,I145204,I145207,I145210,I145213,I145259,I145262,I145265,I145268,I145271,I145274,I145277,I145280,I145283,I145329,I145332,I145335,I145338,I145341,I145344,I145347,I145350,I145353,I145399,I145402,I145405,I145408,I145411,I145414,I145417,I145420,I145423,I145469,I145472,I145475,I145478,I145481,I145484,I145487,I145490,I145493,I145539,I145542,I145545,I145548,I145551,I145554,I145557,I145560,I145563,I145609,I145612,I145615,I145618,I145621,I145624,I145627,I145630,I145633,I145679,I145682,I145685,I145688,I145691,I145694,I145697,I145700,I145703,I145749,I145752,I145755,I145758,I145761,I145764,I145767,I145770,I145816,I145819,I145822,I145825,I145828,I145831,I145834,I145837,I145840,I145843,I145889,I145892,I145895,I145898,I145901,I145904,I145907,I145910,I145956,I145959,I145962,I145965,I145968,I145971,I145974,I145977,I145980,I146026,I146029,I146032,I146035,I146038,I146041,I146044,I146047,I146050,I146053,I146099,I146102,I146105,I146108,I146111,I146114,I146117,I146120,I146123,I146126,I146172,I146175,I146178,I146181,I146184,I146187,I146190,I146193,I146196,I146199,I146245,I146248,I146251,I146254,I146257,I146260,I146263,I146266,I146269,I146315,I146318,I146321,I146324,I146327,I146330,I146333,I146336,I146339,I146385,I146388,I146391,I146394,I146397,I146400,I146403,I146406,I146409,I146412,I146458,I146461,I146464,I146467,I146470,I146473,I146476,I146479,I146482,I146528,I146531,I146534,I146537,I146540,I146543,I146546,I146549,I146552,I146598,I146601,I146604,I146607,I146610,I146613,I146616,I146619,I146665,I146668,I146671,I146674,I146677,I146680,I146683,I146686,I146689,I146735,I146738,I146741,I146744,I146747,I146750,I146753,I146756,I146759,I146805,I146808,I146811,I146814,I146817,I146820,I146823,I146826,I146829,I146832,I146878,I146881,I146884,I146887,I146890,I146893,I146896,I146899,I146902,I146905,I146951,I146954,I146957,I146960,I146963,I146966,I146969,I146972,I146975,I146978,I147024,I147027,I147030,I147033,I147036,I147039,I147042,I147045,I147048,I147094,I147097,I147100,I147103,I147106,I147109,I147112,I147115,I147118,I147164,I147167,I147170,I147173,I147176,I147179,I147182,I147185,I147188,I147191,I147237,I147240,I147243,I147246,I147249,I147252,I147255,I147258,I147261,I147264,I147310,I147313,I147316,I147319,I147322,I147325,I147328,I147331,I147377,I147380,I147383,I147386,I147389,I147392,I147395,I147398,I147401,I147447,I147450,I147453,I147456,I147459,I147462,I147465,I147468,I147471,I147474,I147520,I147523,I147526,I147529,I147532,I147535,I147538,I147541,I147544,I147590,I147593,I147596,I147599,I147602,I147605,I147608,I147611,I147614,I147617,I147663,I147666,I147669,I147672,I147675,I147678,I147681,I147684,I147730,I147733,I147736,I147739,I147742,I147745,I147748,I147751,I147754,I147757,I147803,I147806,I147809,I147812,I147815,I147818,I147821,I147824,I147827,I147873,I147876,I147879,I147882,I147885,I147888,I147891,I147894,I147897,I147943,I147946,I147949,I147952,I147955,I147958,I147961,I147964,I147967,I147970,I148016,I148019,I148022,I148025,I148028,I148031,I148034,I148037,I148040,I148043,I148089,I148092,I148095,I148098,I148101,I148104,I148107,I148110,I148113,I148116,I148162,I148165,I148168,I148171,I148174,I148177,I148180,I148183,I148186,I148232,I148235,I148238,I148241,I148244,I148247,I148250,I148253,I148256,I148302,I148305,I148308,I148311,I148314,I148317,I148320,I148323,I148326,I148372,I148375,I148378,I148381,I148384,I148387,I148390,I148393,I148396,I148442,I148445,I148448,I148451,I148454,I148457,I148460,I148463,I148466,I148469,I148515,I148518,I148521,I148524,I148527,I148530,I148533,I148536,I148539,I148585,I148588,I148591,I148594,I148597,I148600,I148603,I148606,I148609,I148655,I148658,I148661,I148664,I148667,I148670,I148673,I148676,I148679,I148682,I148728,I148731,I148734,I148737,I148740,I148743,I148746,I148749,I148795,I148798,I148801,I148804,I148807,I148810,I148813,I148816,I148819,I148822,I148868,I148871,I148874,I148877,I148880,I148883,I148886,I148889,I148892,I148938,I148941,I148944,I148947,I148950,I148953,I148956,I148959,I148962,I149008,I149011,I149014,I149017,I149020,I149023,I149026,I149029,I149032,I149035,I149081,I149084,I149087,I149090,I149093,I149096,I149099,I149102,I149105,I149151,I149154,I149157,I149160,I149163,I149166,I149169,I149172,I149175,I149221,I149224,I149227,I149230,I149233,I149236,I149239,I149242,I149245,I149291,I149294,I149297,I149300,I149303,I149306,I149309,I149312,I149358,I149361,I149364,I149367,I149370,I149373,I149376,I149379,I149382,I149385,I149431,I149434,I149437,I149440,I149443,I149446,I149449,I149452,I149455,I149501,I149504,I149507,I149510,I149513,I149516,I149519,I149522,I149568,I149571,I149574,I149577,I149580,I149583,I149586,I149589,I149592,I149595,I149641,I149644,I149647,I149650,I149653,I149656,I149659,I149662,I149665,I149668,I149714,I149717,I149720,I149723,I149726,I149729,I149732,I149735,I149738,I149741,I149787,I149790,I149793,I149796,I149799,I149802,I149805,I149808,I149811,I149857,I149860,I149863,I149866,I149869,I149872,I149875,I149878,I149881,I149884,I149930,I149933,I149936,I149939,I149942,I149945,I149948,I149951,I149954,I150000,I150003,I150006,I150009,I150012,I150015,I150018,I150021,I150024,I150070,I150073,I150076,I150079,I150082,I150085,I150088,I150091,I150094,I150140,I150143,I150146,I150149,I150152,I150155,I150158,I150161,I150164,I150167,I150213,I150216,I150219,I150222,I150225,I150228,I150231,I150234,I150237,I150283,I150286,I150289,I150292,I150295,I150298,I150301,I150304,I150307,I150353,I150356,I150359,I150362,I150365,I150368,I150371,I150374,I150377,I150423,I150426,I150429,I150432,I150435,I150438,I150441,I150444,I150447,I150450,I150496,I150499,I150502,I150505,I150508,I150511,I150514,I150517,I150520,I150566,I150569,I150572,I150575,I150578,I150581,I150584,I150587,I150590,I150636,I150639,I150642,I150645,I150648,I150651,I150654,I150657,I150660,I150706,I150709,I150712,I150715,I150718,I150721,I150724,I150727,I150730,I150733,I150779,I150782,I150785,I150788,I150791,I150794,I150797,I150800,I150846,I150849,I150852,I150855,I150858,I150861,I150864,I150867,I150870,I150873,I150919,I150922,I150925,I150928,I150931,I150934,I150937,I150940,I150943,I150989,I150992,I150995,I150998,I151001,I151004,I151007,I151010,I151013,I151016,I151062,I151065,I151068,I151071,I151074,I151077,I151080,I151083,I151086,I151132,I151135,I151138,I151141,I151144,I151147,I151150,I151153,I151199,I151202,I151205,I151208,I151211,I151214,I151217,I151220,I151223,I151269,I151272,I151275,I151278,I151281,I151284,I151287,I151290,I151336,I151339,I151342,I151345,I151348,I151351,I151354,I151357,I151403,I151406,I151409,I151412,I151415,I151418,I151421,I151424,I151427,I151473,I151476,I151479,I151482,I151485,I151488,I151491,I151494,I151497,I151500,I151546,I151549,I151552,I151555,I151558,I151561,I151564,I151567,I151570,I151616,I151619,I151622,I151625,I151628,I151631,I151634,I151637,I151640,I151686,I151689,I151692,I151695,I151698,I151701,I151704,I151707,I151710,I151756,I151759,I151762,I151765,I151768,I151771,I151774,I151777,I151823,I151826,I151829,I151832,I151835,I151838,I151841,I151844,I151847,I151893,I151896,I151899,I151902,I151905,I151908,I151911,I151914,I151960,I151963,I151966,I151969,I151972,I151975,I151978,I151981,I151984,I151987,I152033,I152036,I152039,I152042,I152045,I152048,I152051,I152054,I152057,I152103,I152106,I152109,I152112,I152115,I152118,I152121,I152124,I152127,I152173,I152176,I152179,I152182,I152185,I152188,I152191,I152194,I152197,I152243,I152246,I152249,I152252,I152255,I152258,I152261,I152264,I152267,I152270,I152316,I152319,I152322,I152325,I152328,I152331,I152334,I152337,I152383,I152386,I152389,I152392,I152395,I152398,I152401,I152404,I152407,I152453,I152456,I152459,I152462,I152465,I152468,I152471,I152474,I152477,I152480,I152526,I152529,I152532,I152535,I152538,I152541,I152544,I152547,I152550,I152596,I152599,I152602,I152605,I152608,I152611,I152614,I152617,I152620,I152623,I152669,I152672,I152675,I152678,I152681,I152684,I152687,I152690,I152693,I152739,I152742,I152745,I152748,I152751,I152754,I152757,I152760,I152763,I152809,I152812,I152815,I152818,I152821,I152824,I152827,I152830,I152833,I152879,I152882,I152885,I152888,I152891,I152894,I152897,I152900,I152903,I152949,I152952,I152955,I152958,I152961,I152964,I152967,I152970,I152973,I153019,I153022,I153025,I153028,I153031,I153034,I153037,I153040,I153086,I153089,I153092,I153095,I153098,I153101,I153104,I153107,I153110,I153156,I153159,I153162,I153165,I153168,I153171,I153174,I153177,I153180,I153226,I153229,I153232,I153235,I153238,I153241,I153244,I153247,I153250,I153253,I153299,I153302,I153305,I153308,I153311,I153314,I153317,I153320,I153323,I153369,I153372,I153375,I153378,I153381,I153384,I153387,I153390,I153393,I153439,I153442,I153445,I153448,I153451,I153454,I153457,I153460,I153463,I153509,I153512,I153515,I153518,I153521,I153524,I153527,I153530,I153533,I153536,I153582,I153585,I153588,I153591,I153594,I153597,I153600,I153603,I153649,I153652,I153655,I153658,I153661,I153664,I153667,I153670,I153673,I153719,I153722,I153725,I153728,I153731,I153734,I153737,I153740,I153743,I153789,I153792,I153795,I153798,I153801,I153804,I153807,I153810,I153813,I153859,I153862,I153865,I153868,I153871,I153874,I153877,I153880,I153883,I153886,I153932,I153935,I153938,I153941,I153944,I153947,I153950,I153953,I153956,I153959,I154005,I154008,I154011,I154014,I154017,I154020,I154023,I154026,I154029,I154075,I154078,I154081,I154084,I154087,I154090,I154093,I154096,I154099,I154102,I154148,I154151,I154154,I154157,I154160,I154163,I154166,I154169,I154172,I154218,I154221,I154224,I154227,I154230,I154233,I154236,I154239,I154242,I154288,I154291,I154294,I154297,I154300,I154303,I154306,I154309,I154312,I154358,I154361,I154364,I154367,I154370,I154373,I154376,I154379,I154382,I154385,I154431,I154434,I154437,I154440,I154443,I154446,I154449,I154452,I154455,I154501,I154504,I154507,I154510,I154513,I154516,I154519,I154522,I154525,I154571,I154574,I154577,I154580,I154583,I154586,I154589,I154592,I154595,I154641,I154644,I154647,I154650,I154653,I154656,I154659,I154662,I154665,I154668,I154714,I154717,I154720,I154723,I154726,I154729,I154732,I154735,I154738,I154741,I154787,I154790,I154793,I154796,I154799,I154802,I154805,I154808,I154811,I154814,I154860,I154863,I154866,I154869,I154872,I154875,I154878,I154881,I154884,I154930,I154933,I154936,I154939,I154942,I154945,I154948,I154951,I154997,I155000,I155003,I155006,I155009,I155012,I155015,I155018,I155021,I155067,I155070,I155073,I155076,I155079,I155082,I155085,I155088,I155091,I155094,I155140,I155143,I155146,I155149,I155152,I155155,I155158,I155161,I155164,I155167,I155213,I155216,I155219,I155222,I155225,I155228,I155231,I155234,I155237,I155283,I155286,I155289,I155292,I155295,I155298,I155301,I155304,I155307,I155353,I155356,I155359,I155362,I155365,I155368,I155371,I155374,I155377,I155423,I155426,I155429,I155432,I155435,I155438,I155441,I155444,I155447,I155493,I155496,I155499,I155502,I155505,I155508,I155511,I155514,I155560,I155563,I155566,I155569,I155572,I155575,I155578,I155581,I155584,I155630,I155633,I155636,I155639,I155642,I155645,I155648,I155651,I155654,I155657,I155703,I155706,I155709,I155712,I155715,I155718,I155721,I155724,I155727,I155730,I155776,I155779,I155782,I155785,I155788,I155791,I155794,I155797,I155800,I155846,I155849,I155852,I155855,I155858,I155861,I155864,I155867,I155870,I155916,I155919,I155922,I155925,I155928,I155931,I155934,I155937,I155940,I155986,I155989,I155992,I155995,I155998,I156001,I156004,I156007,I156010,I156056,I156059,I156062,I156065,I156068,I156071,I156074,I156077,I156080,I156083,I156129,I156132,I156135,I156138,I156141,I156144,I156147,I156150,I156153,I156199,I156202,I156205,I156208,I156211,I156214,I156217,I156220,I156223,I156226,I156272,I156275,I156278,I156281,I156284,I156287,I156290,I156293,I156296,I156342,I156345,I156348,I156351,I156354,I156357,I156360,I156363,I156366,I156412,I156415,I156418,I156421,I156424,I156427,I156430,I156433,I156436,I156482,I156485,I156488,I156491,I156494,I156497,I156500,I156503,I156506,I156552,I156555,I156558,I156561,I156564,I156567,I156570,I156573,I156576,I156579,I156625,I156628,I156631,I156634,I156637,I156640,I156643,I156646,I156649,I156695,I156698,I156701,I156704,I156707,I156710,I156713,I156716,I156762,I156765,I156768,I156771,I156774,I156777,I156780,I156783,I156786,I156832,I156835,I156838,I156841,I156844,I156847,I156850,I156853,I156856,I156902,I156905,I156908,I156911,I156914,I156917,I156920,I156923,I156926,I156929,I156975,I156978,I156981,I156984,I156987,I156990,I156993,I156996,I156999,I157002,I157048,I157051,I157054,I157057,I157060,I157063,I157066,I157069,I157072,I157118,I157121,I157124,I157127,I157130,I157133,I157136,I157139,I157142,I157188,I157191,I157194,I157197,I157200,I157203,I157206,I157209,I157212,I157258,I157261,I157264,I157267,I157270,I157273,I157276,I157279,I157282,I157285,I157331,I157334,I157337,I157340,I157343,I157346,I157349,I157352,I157355,I157358,I157404,I157407,I157410,I157413,I157416,I157419,I157422,I157425,I157428,I157474,I157477,I157480,I157483,I157486,I157489,I157492,I157495,I157541,I157544,I157547,I157550,I157553,I157556,I157559,I157562,I157565,I157568,I157614,I157617,I157620,I157623,I157626,I157629,I157632,I157635,I157638,I157684,I157687,I157690,I157693,I157696,I157699,I157702,I157705,I157708,I157711,I157757,I157760,I157763,I157766,I157769,I157772,I157775,I157778,I157781,I157784,I157830,I157833,I157836,I157839,I157842,I157845,I157848,I157851,I157854,I157857,I157903,I157906,I157909,I157912,I157915,I157918,I157921,I157924,I157927,I157973,I157976,I157979,I157982,I157985,I157988,I157991,I157994,I157997,I158000,I158046,I158049,I158052,I158055,I158058,I158061,I158064,I158067,I158113,I158116,I158119,I158122,I158125,I158128,I158131,I158134,I158137,I158183,I158186,I158189,I158192,I158195,I158198,I158201,I158204,I158207,I158210,I158256,I158259,I158262,I158265,I158268,I158271,I158274,I158277,I158280,I158326,I158329,I158332,I158335,I158338,I158341,I158344,I158347,I158350,I158396,I158399,I158402,I158405,I158408,I158411,I158414,I158417,I158420,I158466,I158469,I158472,I158475,I158478,I158481,I158484,I158487,I158490,I158536,I158539,I158542,I158545,I158548,I158551,I158554,I158557,I158603,I158606,I158609,I158612,I158615,I158618,I158621,I158624,I158670,I158673,I158676,I158679,I158682,I158685,I158688,I158691,I158694,I158697,I158743,I158746,I158749,I158752,I158755,I158758,I158761,I158764,I158767,I158813,I158816,I158819,I158822,I158825,I158828,I158831,I158834,I158837,I158840,I158886,I158889,I158892,I158895,I158898,I158901,I158904,I158907,I158953,I158956,I158959,I158962,I158965,I158968,I158971,I158974,I158977,I158980,I159026,I159029,I159032,I159035,I159038,I159041,I159044,I159047,I159050,I159096,I159099,I159102,I159105,I159108,I159111,I159114,I159117,I159120,I159123,I159169,I159172,I159175,I159178,I159181,I159184,I159187,I159190,I159193,I159239,I159242,I159245,I159248,I159251,I159254,I159257,I159260,I159263,I159266,I159312,I159315,I159318,I159321,I159324,I159327,I159330,I159333,I159336,I159382,I159385,I159388,I159391,I159394,I159397,I159400,I159403,I159449,I159452,I159455,I159458,I159461,I159464,I159467,I159470,I159473,I159519,I159522,I159525,I159528,I159531,I159534,I159537,I159540,I159586,I159589,I159592,I159595,I159598,I159601,I159604,I159607,I159610,I159656,I159659,I159662,I159665,I159668,I159671,I159674,I159677,I159680,I159726,I159729,I159732,I159735,I159738,I159741,I159744,I159747,I159750,I159796,I159799,I159802,I159805,I159808,I159811,I159814,I159817,I159820,I159823,I159942,I159945,I159948,I159951,I159954,I159957,I159960,I159963,I159966,I159969,I160015,I160018,I160021,I160024,I160027,I160030,I160033,I160036,I160039,I160085,I160088,I160091,I160094,I160097,I160100,I160103,I160106,I160152,I160155,I160158,I160161,I160164,I160167,I160170,I160173,I160176,I160222,I160225,I160228,I160231,I160234,I160237,I160240,I160243,I160246,I160249,I160295,I160298,I160301,I160304,I160307,I160310,I160313,I160316,I160362,I160365,I160368,I160371,I160374,I160377,I160380,I160383,I160386,I160432,I160435,I160438,I160441,I160444,I160447,I160450,I160453,I160456,I160459,I160505,I160508,I160511,I160514,I160517,I160520,I160523,I160526,I160572,I160575,I160578,I160581,I160584,I160587,I160590,I160593,I160596,I160642,I160645,I160648,I160651,I160654,I160657,I160660,I160663,I160666,I160669,I160715,I160718,I160721,I160724,I160727,I160730,I160733,I160736,I160739,I160785,I160788,I160791,I160794,I160797,I160800,I160803,I160806,I160809,I160855,I160858,I160861,I160864,I160867,I160870,I160873,I160876,I160879,I160925,I160928,I160931,I160934,I160937,I160940,I160943,I160946,I160949,I160952,I160998,I161001,I161004,I161007,I161010,I161013,I161016,I161019,I161022,I161025,I161071,I161074,I161077,I161080,I161083,I161086,I161089,I161092,I161095,I161141,I161144,I161147,I161150,I161153,I161156,I161159,I161162,I161165,I161168,I161214,I161217,I161220,I161223,I161226,I161229,I161232,I161235,I161238,I161284,I161287,I161290,I161293,I161296,I161299,I161302,I161305,I161308,I161354,I161357,I161360,I161363,I161366,I161369,I161372,I161375,I161378,I161424,I161427,I161430,I161433,I161436,I161439,I161442,I161445,I161448,I161494,I161497,I161500,I161503,I161506,I161509,I161512,I161515,I161518,I161521,I161567,I161570,I161573,I161576,I161579,I161582,I161585,I161588,I161591,I161637,I161640,I161643,I161646,I161649,I161652,I161655,I161658,I161661,I161707,I161710,I161713,I161716,I161719,I161722,I161725,I161728,I161731,I161777,I161780,I161783,I161786,I161789,I161792,I161795,I161798,I161844,I161847,I161850,I161853,I161856,I161859,I161862,I161865,I161868,I161914,I161917,I161920,I161923,I161926,I161929,I161932,I161935,I161938,I161984,I161987,I161990,I161993,I161996,I161999,I162002,I162005,I162008,I162011,I162057,I162060,I162063,I162066,I162069,I162072,I162075,I162078,I162081,I162127,I162130,I162133,I162136,I162139,I162142,I162145,I162148,I162151,I162197,I162200,I162203,I162206,I162209,I162212,I162215,I162218,I162221,I162267,I162270,I162273,I162276,I162279,I162282,I162285,I162288,I162291,I162337,I162340,I162343,I162346,I162349,I162352,I162355,I162358,I162404,I162407,I162410,I162413,I162416,I162419,I162422,I162425,I162428,I162431,I162477,I162480,I162483,I162486,I162489,I162492,I162495,I162498,I162501,I162547,I162550,I162553,I162556,I162559,I162562,I162565,I162568,I162571,I162617,I162620,I162623,I162626,I162629,I162632,I162635,I162638,I162641,I162644,I162690,I162693,I162696,I162699,I162702,I162705,I162708,I162711,I162714,I162760,I162763,I162766,I162769,I162772,I162775,I162778,I162781,I162784,I162830,I162833,I162836,I162839,I162842,I162845,I162848,I162851,I162854,I162900,I162903,I162906,I162909,I162912,I162915,I162918,I162921,I162924,I162927,I162973,I162976,I162979,I162982,I162985,I162988,I162991,I162994,I162997,I163043,I163046,I163049,I163052,I163055,I163058,I163061,I163064,I163067,I163070,I163116,I163119,I163122,I163125,I163128,I163131,I163134,I163137,I163140,I163186,I163189,I163192,I163195,I163198,I163201,I163204,I163207,I163210,I163213,I163259,I163262,I163265,I163268,I163271,I163274,I163277,I163280,I163283,I163286,I163332,I163335,I163338,I163341,I163344,I163347,I163350,I163353,I163356,I163359,I163405,I163408,I163411,I163414,I163417,I163420,I163423,I163426,I163429,I163475,I163478,I163481,I163484,I163487,I163490,I163493,I163496,I163542,I163545,I163548,I163551,I163554,I163557,I163560,I163563,I163566,I163612,I163615,I163618,I163621,I163624,I163627,I163630,I163633,I163679,I163682,I163685,I163688,I163691,I163694,I163697,I163700,I163703,I163749,I163752,I163755,I163758,I163761,I163764,I163767,I163770,I163816,I163819,I163822,I163825,I163828,I163831,I163834,I163837,I163840,I163843,I163889,I163892,I163895,I163898,I163901,I163904,I163907,I163910,I163913,I163916,I163962,I163965,I163968,I163971,I163974,I163977,I163980,I163983,I164029,I164032,I164035,I164038,I164041,I164044,I164047,I164050,I164053,I164099,I164102,I164105,I164108,I164111,I164114,I164117,I164120,I164123,I164126,I164172,I164175,I164178,I164181,I164184,I164187,I164190,I164193,I164196,I164242,I164245,I164248,I164251,I164254,I164257,I164260,I164263,I164309,I164312,I164315,I164318,I164321,I164324,I164327,I164330,I164333,I164379,I164382,I164385,I164388,I164391,I164394,I164397,I164400,I164446,I164449,I164452,I164455,I164458,I164461,I164464,I164467,I164470,I164516,I164519,I164522,I164525,I164528,I164531,I164534,I164537,I164540,I164586,I164589,I164592,I164595,I164598,I164601,I164604,I164607,I164610,I164613,I164659,I164662,I164665,I164668,I164671,I164674,I164677,I164680,I164726,I164729,I164732,I164735,I164738,I164741,I164744,I164747,I164750,I164796,I164799,I164802,I164805,I164808,I164811,I164814,I164817,I164820,I164866,I164869,I164872,I164875,I164878,I164881,I164884,I164887,I164933,I164936,I164939,I164942,I164945,I164948,I164951,I164954,I164957,I164960,I165006,I165009,I165012,I165015,I165018,I165021,I165024,I165027,I165030,I165076,I165079,I165082,I165085,I165088,I165091,I165094,I165097,I165100,I165103,I165149,I165152,I165155,I165158,I165161,I165164,I165167,I165170,I165216,I165219,I165222,I165225,I165228,I165231,I165234,I165237,I165240,I165286,I165289,I165292,I165295,I165298,I165301,I165304,I165307,I165310,I165313,I165359,I165362,I165365,I165368,I165371,I165374,I165377,I165380,I165383,I165386,I165432,I165435,I165438,I165441,I165444,I165447,I165450,I165453,I165456,I165459,I165505,I165508,I165511,I165514,I165517,I165520,I165523,I165526,I165529,I165575,I165578,I165581,I165584,I165587,I165590,I165593,I165596,I165599,I165645,I165648,I165651,I165654,I165657,I165660,I165663,I165666,I165669,I165672,I165718,I165721,I165724,I165727,I165730,I165733,I165736,I165739,I165742,I165788,I165791,I165794,I165797,I165800,I165803,I165806,I165809,I165812,I165858,I165861,I165864,I165867,I165870,I165873,I165876,I165879,I165925,I165928,I165931,I165934,I165937,I165940,I165943,I165946,I165949,I165952,I165998,I166001,I166004,I166007,I166010,I166013,I166016,I166019,I166022,I166025,I166071,I166074,I166077,I166080,I166083,I166086,I166089,I166092,I166095,I166141,I166144,I166147,I166150,I166153,I166156,I166159,I166162,I166165,I166211,I166214,I166217,I166220,I166223,I166226,I166229,I166232,I166235,I166281,I166284,I166287,I166290,I166293,I166296,I166299,I166302,I166305,I166351,I166354,I166357,I166360,I166363,I166366,I166369,I166372,I166375,I166378,I166424,I166427,I166430,I166433,I166436,I166439,I166442,I166445,I166448,I166494,I166497,I166500,I166503,I166506,I166509,I166512,I166515,I166518,I166564,I166567,I166570,I166573,I166576,I166579,I166582,I166585,I166588,I166591,I166637,I166640,I166643,I166646,I166649,I166652,I166655,I166658,I166661,I166707,I166710,I166713,I166716,I166719,I166722,I166725,I166728,I166731,I166777,I166780,I166783,I166786,I166789,I166792,I166795,I166798,I166801,I166847,I166850,I166853,I166856,I166859,I166862,I166865,I166868,I166871,I166917,I166920,I166923,I166926,I166929,I166932,I166935,I166938,I166941,I166987,I166990,I166993,I166996,I166999,I167002,I167005,I167008,I167011,I167057,I167060,I167063,I167066,I167069,I167072,I167075,I167078,I167081,I167127,I167130,I167133,I167136,I167139,I167142,I167145,I167148,I167151,I167197,I167200,I167203,I167206,I167209,I167212,I167215,I167218,I167221,I167267,I167270,I167273,I167276,I167279,I167282,I167285,I167288,I167291,I167337,I167340,I167343,I167346,I167349,I167352,I167355,I167358,I167361,I167407,I167410,I167413,I167416,I167419,I167422,I167425,I167428,I167431,I167434,I167480,I167483,I167486,I167489,I167492,I167495,I167498,I167501,I167504,I167507,I167553,I167556,I167559,I167562,I167565,I167568,I167571,I167574,I167577,I167580,I167626,I167629,I167632,I167635,I167638,I167641,I167644,I167647,I167650,I167653,I167699,I167702,I167705,I167708,I167711,I167714,I167717,I167720,I167723,I167726,I167772,I167775,I167778,I167781,I167784,I167787,I167790,I167793,I167796,I167799,I167845,I167848,I167851,I167854,I167857,I167860,I167863,I167866,I167912,I167915,I167918,I167921,I167924,I167927,I167930,I167933,I167979,I167982,I167985,I167988,I167991,I167994,I167997,I168000,I168003,I168049,I168052,I168055,I168058,I168061,I168064,I168067,I168070,I168073,I168119,I168122,I168125,I168128,I168131,I168134,I168137,I168140,I168143,I168189,I168192,I168195,I168198,I168201,I168204,I168207,I168210,I168213,I168216,I168262,I168265,I168268,I168271,I168274,I168277,I168280,I168283,I168329,I168332,I168335,I168338,I168341,I168344,I168347,I168350,I168353,I168399,I168402,I168405,I168408,I168411,I168414,I168417,I168420,I168423,I168426,I168472,I168475,I168478,I168481,I168484,I168487,I168490,I168493,I168496,I168542,I168545,I168548,I168551,I168554,I168557,I168560,I168563,I168566,I168612,I168615,I168618,I168621,I168624,I168627,I168630,I168633,I168636,I168639,I168685,I168688,I168691,I168694,I168697,I168700,I168703,I168706,I168709,I168755,I168758,I168761,I168764,I168767,I168770,I168773,I168776,I168822,I168825,I168828,I168831,I168834,I168837,I168840,I168843,I168846,I168849,I168895,I168898,I168901,I168904,I168907,I168910,I168913,I168916,I168919,I168965,I168968,I168971,I168974,I168977,I168980,I168983,I168986,I169032,I169035,I169038,I169041,I169044,I169047,I169050,I169053,I169056,I169102,I169105,I169108,I169111,I169114,I169117,I169120,I169123,I169169,I169172,I169175,I169178,I169181,I169184,I169187,I169190,I169193,I169239,I169242,I169245,I169248,I169251,I169254,I169257,I169260,I169263,I169309,I169312,I169315,I169318,I169321,I169324,I169327,I169330,I169333,I169379,I169382,I169385,I169388,I169391,I169394,I169397,I169400,I169403,I169449,I169452,I169455,I169458,I169461,I169464,I169467,I169470,I169473,I169476,I169522,I169525,I169528,I169531,I169534,I169537,I169540,I169543,I169546,I169592,I169595,I169598,I169601,I169604,I169607,I169610,I169613,I169616,I169619,I169665,I169668,I169671,I169674,I169677,I169680,I169683,I169686,I169732,I169735,I169738,I169741,I169744,I169747,I169750,I169753,I169756,I169802,I169805,I169808,I169811,I169814,I169817,I169820,I169823,I169826,I169872,I169875,I169878,I169881,I169884,I169887,I169890,I169893,I169896,I169899,I169945,I169948,I169951,I169954,I169957,I169960,I169963,I169966,I169969,I170015,I170018,I170021,I170024,I170027,I170030,I170033,I170036,I170039,I170042,I170088,I170091,I170094,I170097,I170100,I170103,I170106,I170109,I170112,I170115,I170161,I170164,I170167,I170170,I170173,I170176,I170179,I170182,I170185,I170188,I170234,I170237,I170240,I170243,I170246,I170249,I170252,I170255,I170258,I170304,I170307,I170310,I170313,I170316,I170319,I170322,I170325,I170328,I170331,I170377,I170380,I170383,I170386,I170389,I170392,I170395,I170398,I170401,I170404,I170450,I170453,I170456,I170459,I170462,I170465,I170468,I170471,I170474,I170520,I170523,I170526,I170529,I170532,I170535,I170538,I170541,I170544,I170590,I170593,I170596,I170599,I170602,I170605,I170608,I170611,I170614,I170660,I170663,I170666,I170669,I170672,I170675,I170678,I170681,I170684,I170687,I170733,I170736,I170739,I170742,I170745,I170748,I170751,I170754,I170757,I170803,I170806,I170809,I170812,I170815,I170818,I170821,I170824,I170827,I170873,I170876,I170879,I170882,I170885,I170888,I170891,I170894,I170940,I170943,I170946,I170949,I170952,I170955,I170958,I170961,I170964,I171010,I171013,I171016,I171019,I171022,I171025,I171028,I171031,I171077,I171080,I171083,I171086,I171089,I171092,I171095,I171098,I171101,I171104,I171150,I171153,I171156,I171159,I171162,I171165,I171168,I171171,I171174,I171177,I171223,I171226,I171229,I171232,I171235,I171238,I171241,I171244,I171247,I171250,I171296,I171299,I171302,I171305,I171308,I171311,I171314,I171317,I171320,I171323,I171369,I171372,I171375,I171378,I171381,I171384,I171387,I171390,I171393,I171396,I171442,I171445,I171448,I171451,I171454,I171457,I171460,I171463,I171466,I171512,I171515,I171518,I171521,I171524,I171527,I171530,I171533,I171536,I171539,I171585,I171588,I171591,I171594,I171597,I171600,I171603,I171606,I171609,I171655,I171658,I171661,I171664,I171667,I171670,I171673,I171676,I171679,I171725,I171728,I171731,I171734,I171737,I171740,I171743,I171746,I171749,I171795,I171798,I171801,I171804,I171807,I171810,I171813,I171816,I171819,I171865,I171868,I171871,I171874,I171877,I171880,I171883,I171886,I171889,I171892,I171938,I171941,I171944,I171947,I171950,I171953,I171956,I171959,I171962,I171965,I172011,I172014,I172017,I172020,I172023,I172026,I172029,I172032,I172035,I172081,I172084,I172087,I172090,I172093,I172096,I172099,I172102,I172148,I172151,I172154,I172157,I172160,I172163,I172166,I172169,I172172,I172175,I172221,I172224,I172227,I172230,I172233,I172236,I172239,I172242,I172245,I172248,I172294,I172297,I172300,I172303,I172306,I172309,I172312,I172315,I172318,I172321,I172367,I172370,I172373,I172376,I172379,I172382,I172385,I172388,I172391,I172437,I172440,I172443,I172446,I172449,I172452,I172455,I172458,I172461,I172464,I172510,I172513,I172516,I172519,I172522,I172525,I172528,I172531,I172577,I172580,I172583,I172586,I172589,I172592,I172595,I172598,I172601,I172647,I172650,I172653,I172656,I172659,I172662,I172665,I172668,I172671,I172717,I172720,I172723,I172726,I172729,I172732,I172735,I172738,I172741,I172787,I172790,I172793,I172796,I172799,I172802,I172805,I172808,I172811,I172814,I172860,I172863,I172866,I172869,I172872,I172875,I172878,I172881,I172884,I172930,I172933,I172936,I172939,I172942,I172945,I172948,I172951,I172954,I173000,I173003,I173006,I173009,I173012,I173015,I173018,I173021,I173024,I173070,I173073,I173076,I173079,I173082,I173085,I173088,I173091,I173094,I173097,I173143,I173146,I173149,I173152,I173155,I173158,I173161,I173164,I173167,I173213,I173216,I173219,I173222,I173225,I173228,I173231,I173234,I173237,I173283,I173286,I173289,I173292,I173295,I173298,I173301,I173304,I173350,I173353,I173356,I173359,I173362,I173365,I173368,I173371,I173374,I173377,I173423,I173426,I173429,I173432,I173435,I173438,I173441,I173444,I173447,I173493,I173496,I173499,I173502,I173505,I173508,I173511,I173514,I173517,I173563,I173566,I173569,I173572,I173575,I173578,I173581,I173584,I173587,I173590,I173636,I173639,I173642,I173645,I173648,I173651,I173654,I173657,I173660,I173706,I173709,I173712,I173715,I173718,I173721,I173724,I173727,I173730,I173733,I173779,I173782,I173785,I173788,I173791,I173794,I173797,I173800,I173846,I173849,I173852,I173855,I173858,I173861,I173864,I173867,I173870,I173873,I173919,I173922,I173925,I173928,I173931,I173934,I173937,I173940,I173943,I173946,I173992,I173995,I173998,I174001,I174004,I174007,I174010,I174013,I174016,I174062,I174065,I174068,I174071,I174074,I174077,I174080,I174083,I174129,I174132,I174135,I174138,I174141,I174144,I174147,I174150,I174196,I174199,I174202,I174205,I174208,I174211,I174214,I174217,I174220,I174223,I174269,I174272,I174275,I174278,I174281,I174284,I174287,I174290,I174293,I174339,I174342,I174345,I174348,I174351,I174354,I174357,I174360,I174363,I174366,I174412,I174415,I174418,I174421,I174424,I174427,I174430,I174433,I174436,I174482,I174485,I174488,I174491,I174494,I174497,I174500,I174503,I174549,I174552,I174555,I174558,I174561,I174564,I174567,I174570,I174573,I174619,I174622,I174625,I174628,I174631,I174634,I174637,I174640,I174643,I174689,I174692,I174695,I174698,I174701,I174704,I174707,I174710,I174713,I174716,I174762,I174765,I174768,I174771,I174774,I174777,I174780,I174783,I174786,I174789,I174835,I174838,I174841,I174844,I174847,I174850,I174853,I174856,I174859,I174862,I174908,I174911,I174914,I174917,I174920,I174923,I174926,I174929,I174932,I174978,I174981,I174984,I174987,I174990,I174993,I174996,I174999,I175002,I175048,I175051,I175054,I175057,I175060,I175063,I175066,I175069,I175072,I175118,I175121,I175124,I175127,I175130,I175133,I175136,I175139,I175142,I175188,I175191,I175194,I175197,I175200,I175203,I175206,I175209,I175255,I175258,I175261,I175264,I175267,I175270,I175273,I175276,I175279,I175325,I175328,I175331,I175334,I175337,I175340,I175343,I175346,I175349,I175395,I175398,I175401,I175404,I175407,I175410,I175413,I175416,I175419,I175422,I175468,I175471,I175474,I175477,I175480,I175483,I175486,I175489,I175492,I175538,I175541,I175544,I175547,I175550,I175553,I175556,I175559,I175562,I175565,I175611,I175614,I175617,I175620,I175623,I175626,I175629,I175632,I175635,I175638,I175684,I175687,I175690,I175693,I175696,I175699,I175702,I175705,I175708,I175754,I175757,I175760,I175763,I175766,I175769,I175772,I175775,I175778,I175824,I175827,I175830,I175833,I175836,I175839,I175842,I175845,I175848,I175894,I175897,I175900,I175903,I175906,I175909,I175912,I175915,I175961,I175964,I175967,I175970,I175973,I175976,I175979,I175982,I175985,I175988,I176034,I176037,I176040,I176043,I176046,I176049,I176052,I176055,I176058,I176061,I176107,I176110,I176113,I176116,I176119,I176122,I176125,I176128,I176131,I176134,I176180,I176183,I176186,I176189,I176192,I176195,I176198,I176201,I176204,I176207,I176253,I176256,I176259,I176262,I176265,I176268,I176271,I176274,I176320,I176323,I176326,I176329,I176332,I176335,I176338,I176341,I176344,I176390,I176393,I176396,I176399,I176402,I176405,I176408,I176411,I176414,I176417,I176463,I176466,I176469,I176472,I176475,I176478,I176481,I176484,I176487,I176533,I176536,I176539,I176542,I176545,I176548,I176551,I176554,I176557,I176603,I176606,I176609,I176612,I176615,I176618,I176621,I176624,I176627,I176673,I176676,I176679,I176682,I176685,I176688,I176691,I176694,I176697,I176743,I176746,I176749,I176752,I176755,I176758,I176761,I176764,I176767,I176770,I176816,I176819,I176822,I176825,I176828,I176831,I176834,I176837,I176840,I176843,I176889,I176892,I176895,I176898,I176901,I176904,I176907,I176910,I176913,I176959,I176962,I176965,I176968,I176971,I176974,I176977,I176980,I176983,I176986,I177032,I177035,I177038,I177041,I177044,I177047,I177050,I177053,I177099,I177102,I177105,I177108,I177111,I177114,I177117,I177120,I177123,I177169,I177172,I177175,I177178,I177181,I177184,I177187,I177190,I177193,I177239,I177242,I177245,I177248,I177251,I177254,I177257,I177260,I177306,I177309,I177312,I177315,I177318,I177321,I177324,I177327,I177373,I177376,I177379,I177382,I177385,I177388,I177391,I177394,I177397,I177400,I177446,I177449,I177452,I177455,I177458,I177461,I177464,I177467,I177470,I177516,I177519,I177522,I177525,I177528,I177531,I177534,I177537,I177540,I177586,I177589,I177592,I177595,I177598,I177601,I177604,I177607,I177610,I177656,I177659,I177662,I177665,I177668,I177671,I177674,I177677,I177680,I177726,I177729,I177732,I177735,I177738,I177741,I177744,I177747,I177750,I177796,I177799,I177802,I177805,I177808,I177811,I177814,I177817,I177820,I177866,I177869,I177872,I177875,I177878,I177881,I177884,I177887,I177890,I177936,I177939,I177942,I177945,I177948,I177951,I177954,I177957,I177960,I177963,I178009,I178012,I178015,I178018,I178021,I178024,I178027,I178030,I178033,I178079,I178082,I178085,I178088,I178091,I178094,I178097,I178100,I178103,I178149,I178152,I178155,I178158,I178161,I178164,I178167,I178170,I178173,I178219,I178222,I178225,I178228,I178231,I178234,I178237,I178240,I178243,I178289,I178292,I178295,I178298,I178301,I178304,I178307,I178310,I178313,I178359,I178362,I178365,I178368,I178371,I178374,I178377,I178380,I178383,I178386,I178432,I178435,I178438,I178441,I178444,I178447,I178450,I178453,I178456,I178502,I178505,I178508,I178511,I178514,I178517,I178520,I178523,I178526,I178572,I178575,I178578,I178581,I178584,I178587,I178590,I178593,I178596,I178642,I178645,I178648,I178651,I178654,I178657,I178660,I178663,I178666,I178669,I178715,I178718,I178721,I178724,I178727,I178730,I178733,I178736,I178739,I178785,I178788,I178791,I178794,I178797,I178800,I178803,I178806,I178852,I178855,I178858,I178861,I178864,I178867,I178870,I178873,I178876,I178922,I178925,I178928,I178931,I178934,I178937,I178940,I178943,I178989,I178992,I178995,I178998,I179001,I179004,I179007,I179010,I179013,I179016,I179062,I179065,I179068,I179071,I179074,I179077,I179080,I179083,I179086,I179132,I179135,I179138,I179141,I179144,I179147,I179150,I179153,I179156,I179159,I179205,I179208,I179211,I179214,I179217,I179220,I179223,I179226,I179229,I179232,I179278,I179281,I179284,I179287,I179290,I179293,I179296,I179299,I179345,I179348,I179351,I179354,I179357,I179360,I179363,I179366,I179369,I179372,I179418,I179421,I179424,I179427,I179430,I179433,I179436,I179439,I179442,I179488,I179491,I179494,I179497,I179500,I179503,I179506,I179509,I179512,I179515,I179631,I179634,I179637,I179640,I179643,I179646,I179649,I179652,I179655,I179658,I179704,I179707,I179710,I179713,I179716,I179719,I179722,I179725,I179728,I179774,I179777,I179780,I179783,I179786,I179789,I179792,I179795,I179841,I179844,I179847,I179850,I179853,I179856,I179859,I179862,I179865,I179911,I179914,I179917,I179920,I179923,I179926,I179929,I179932,I179935,I179938,I179984,I179987,I179990,I179993,I179996,I179999,I180002,I180005,I180008,I180011,I180057,I180060,I180063,I180066,I180069,I180072,I180075,I180078,I180081,I180127,I180130,I180133,I180136,I180139,I180142,I180145,I180148,I180151,I180197,I180200,I180203,I180206,I180209,I180212,I180215,I180218,I180221,I180224,I180270,I180273,I180276,I180279,I180282,I180285,I180288,I180291,I180294,I180340,I180343,I180346,I180349,I180352,I180355,I180358,I180361,I180364,I180410,I180413,I180416,I180419,I180422,I180425,I180428,I180431,I180434,I180437,I180483,I180486,I180489,I180492,I180495,I180498,I180501,I180504,I180507,I180553,I180556,I180559,I180562,I180565,I180568,I180571,I180574,I180620,I180623,I180626,I180629,I180632,I180635,I180638,I180641,I180644,I180647,I180693,I180696,I180699,I180702,I180705,I180708,I180711,I180714,I180717,I180763,I180766,I180769,I180772,I180775,I180778,I180781,I180784,I180787,I180790,I180836,I180839,I180842,I180845,I180848,I180851,I180854,I180857,I180860,I180906,I180909,I180912,I180915,I180918,I180921,I180924,I180927,I180930,I180976,I180979,I180982,I180985,I180988,I180991,I180994,I180997,I181000,I181046,I181049,I181052,I181055,I181058,I181061,I181064,I181067,I181070,I181116,I181119,I181122,I181125,I181128,I181131,I181134,I181137,I181140,I181143,I181189,I181192,I181195,I181198,I181201,I181204,I181207,I181210,I181256,I181259,I181262,I181265,I181268,I181271,I181274,I181277,I181280,I181326,I181329,I181332,I181335,I181338,I181341,I181344,I181347,I181350,I181353,I181399,I181402,I181405,I181408,I181411,I181414,I181417,I181420,I181423,I181469,I181472,I181475,I181478,I181481,I181484,I181487,I181490,I181493,I181539,I181542,I181545,I181548,I181551,I181554,I181557,I181560,I181563,I181566,I181612,I181615,I181618,I181621,I181624,I181627,I181630,I181633,I181636,I181639,I181685,I181688,I181691,I181694,I181697,I181700,I181703,I181706,I181709,I181755,I181758,I181761,I181764,I181767,I181770,I181773,I181776,I181822,I181825,I181828,I181831,I181834,I181837,I181840,I181843,I181846,I181892,I181895,I181898,I181901,I181904,I181907,I181910,I181913,I181916,I181919,I181965,I181968,I181971,I181974,I181977,I181980,I181983,I181986,I181989,I181992,I182038,I182041,I182044,I182047,I182050,I182053,I182056,I182059,I182062,I182108,I182111,I182114,I182117,I182120,I182123,I182126,I182129,I182132,I182135,I182181,I182184,I182187,I182190,I182193,I182196,I182199,I182202,I182205,I182251,I182254,I182257,I182260,I182263,I182266,I182269,I182272,I182275,I182321,I182324,I182327,I182330,I182333,I182336,I182339,I182342,I182345,I182348,I182394,I182397,I182400,I182403,I182406,I182409,I182412,I182415,I182418,I182464,I182467,I182470,I182473,I182476,I182479,I182482,I182485,I182488,I182491,I182537,I182540,I182543,I182546,I182549,I182552,I182555,I182558,I182561,I182564,I182610,I182613,I182616,I182619,I182622,I182625,I182628,I182631,I182677,I182680,I182683,I182686,I182689,I182692,I182695,I182698,I182744,I182747,I182750,I182753,I182756,I182759,I182762,I182765,I182768,I182814,I182817,I182820,I182823,I182826,I182829,I182832,I182835,I182838,I182884,I182887,I182890,I182893,I182896,I182899,I182902,I182905,I182908,I182911,I182957,I182960,I182963,I182966,I182969,I182972,I182975,I182978,I182981,I183027,I183030,I183033,I183036,I183039,I183042,I183045,I183048,I183051,I183097,I183100,I183103,I183106,I183109,I183112,I183115,I183118,I183121,I183124,I183170,I183173,I183176,I183179,I183182,I183185,I183188,I183191,I183194,I183197,I183243,I183246,I183249,I183252,I183255,I183258,I183261,I183264,I183267,I183313,I183316,I183319,I183322,I183325,I183328,I183331,I183334,I183337,I183340,I183386,I183389,I183392,I183395,I183398,I183401,I183404,I183407,I183410,I183456,I183459,I183462,I183465,I183468,I183471,I183474,I183477,I183480,I183483,I183529,I183532,I183535,I183538,I183541,I183544,I183547,I183550,I183596,I183599,I183602,I183605,I183608,I183611,I183614,I183617,I183620,I183623,I183669,I183672,I183675,I183678,I183681,I183684,I183687,I183690,I183693,I183696,I183742,I183745,I183748,I183751,I183754,I183757,I183760,I183763,I183766,I183769,I183815,I183818,I183821,I183824,I183827,I183830,I183833,I183836,I183839,I183885,I183888,I183891,I183894,I183897,I183900,I183903,I183906,I183909,I183955,I183958,I183961,I183964,I183967,I183970,I183973,I183976,I183979,I184025,I184028,I184031,I184034,I184037,I184040,I184043,I184046,I184049,I184095,I184098,I184101,I184104,I184107,I184110,I184113,I184116,I184119,I184122,I184168,I184171,I184174,I184177,I184180,I184183,I184186,I184189,I184235,I184238,I184241,I184244,I184247,I184250,I184253,I184256,I184259,I184305,I184308,I184311,I184314,I184317,I184320,I184323,I184326,I184329,I184375,I184378,I184381,I184384,I184387,I184390,I184393,I184396,I184399,I184445,I184448,I184451,I184454,I184457,I184460,I184463,I184466,I184469,I184515,I184518,I184521,I184524,I184527,I184530,I184533,I184536,I184539,I184542,I184588,I184591,I184594,I184597,I184600,I184603,I184606,I184609,I184655,I184658,I184661,I184664,I184667,I184670,I184673,I184676,I184722,I184725,I184728,I184731,I184734,I184737,I184740,I184743,I184789,I184792,I184795,I184798,I184801,I184804,I184807,I184810,I184813,I184859,I184862,I184865,I184868,I184871,I184874,I184877,I184880,I184883,I184929,I184932,I184935,I184938,I184941,I184944,I184947,I184950,I184953,I184999,I185002,I185005,I185008,I185011,I185014,I185017,I185020,I185023,I185069,I185072,I185075,I185078,I185081,I185084,I185087,I185090,I185093,I185139,I185142,I185145,I185148,I185151,I185154,I185157,I185160,I185206,I185209,I185212,I185215,I185218,I185221,I185224,I185227,I185230,I185276,I185279,I185282,I185285,I185288,I185291,I185294,I185297,I185300,I185303,I185349,I185352,I185355,I185358,I185361,I185364,I185367,I185370,I185373,I185419,I185422,I185425,I185428,I185431,I185434,I185437,I185440,I185443,I185489,I185492,I185495,I185498,I185501,I185504,I185507,I185510,I185556,I185559,I185562,I185565,I185568,I185571,I185574,I185577,I185580,I185626,I185629,I185632,I185635,I185638,I185641,I185644,I185647,I185650,I185696,I185699,I185702,I185705,I185708,I185711,I185714,I185717,I185720,I185766,I185769,I185772,I185775,I185778,I185781,I185784,I185787,I185790,I185793,I185839,I185842,I185845,I185848,I185851,I185854,I185857,I185860,I185863,I185909,I185912,I185915,I185918,I185921,I185924,I185927,I185930,I185933,I185979,I185982,I185985,I185988,I185991,I185994,I185997,I186000,I186003,I186006,I186052,I186055,I186058,I186061,I186064,I186067,I186070,I186073,I186119,I186122,I186125,I186128,I186131,I186134,I186137,I186140,I186143,I186146,I186192,I186195,I186198,I186201,I186204,I186207,I186210,I186213,I186216,I186262,I186265,I186268,I186271,I186274,I186277,I186280,I186283,I186286,I186289,I186335,I186338,I186341,I186344,I186347,I186350,I186353,I186356,I186359,I186405,I186408,I186411,I186414,I186417,I186420,I186423,I186426,I186429,I186475,I186478,I186481,I186484,I186487,I186490,I186493,I186496,I186499,I186545,I186548,I186551,I186554,I186557,I186560,I186563,I186566,I186612,I186615,I186618,I186621,I186624,I186627,I186630,I186633,I186636,I186639,I186685,I186688,I186691,I186694,I186697,I186700,I186703,I186706,I186709,I186755,I186758,I186761,I186764,I186767,I186770,I186773,I186776,I186779,I186825,I186828,I186831,I186834,I186837,I186840,I186843,I186846,I186849,I186895,I186898,I186901,I186904,I186907,I186910,I186913,I186916,I186919,I186965,I186968,I186971,I186974,I186977,I186980,I186983,I186986,I186989,I187035,I187038,I187041,I187044,I187047,I187050,I187053,I187056,I187059,I187062,I187108,I187111,I187114,I187117,I187120,I187123,I187126,I187129,I187132,I187178,I187181,I187184,I187187,I187190,I187193,I187196,I187199,I187202,I187248,I187251,I187254,I187257,I187260,I187263,I187266,I187269,I187272,I187275,I187321,I187324,I187327,I187330,I187333,I187336,I187339,I187342,I187345,I187391,I187394,I187397,I187400,I187403,I187406,I187409,I187412,I187415,I187418,I187464,I187467,I187470,I187473,I187476,I187479,I187482,I187485,I187488,I187491,I187537,I187540,I187543,I187546,I187549,I187552,I187555,I187558,I187561,I187607,I187610,I187613,I187616,I187619,I187622,I187625,I187628,I187631,I187677,I187680,I187683,I187686,I187689,I187692,I187695,I187698,I187701,I187704,I187750,I187753,I187756,I187759,I187762,I187765,I187768,I187771,I187774,I187820,I187823,I187826,I187829,I187832,I187835,I187838,I187841,I187844,I187890,I187893,I187896,I187899,I187902,I187905,I187908,I187911,I187914,I187917,I187963,I187966,I187969,I187972,I187975,I187978,I187981,I187984,I187987,I188033,I188036,I188039,I188042,I188045,I188048,I188051,I188054,I188057,I188103,I188106,I188109,I188112,I188115,I188118,I188121,I188124,I188127,I188173,I188176,I188179,I188182,I188185,I188188,I188191,I188194,I188197,I188243,I188246,I188249,I188252,I188255,I188258,I188261,I188264,I188267,I188313,I188316,I188319,I188322,I188325,I188328,I188331,I188334,I188337,I188383,I188386,I188389,I188392,I188395,I188398,I188401,I188404,I188450,I188453,I188456,I188459,I188462,I188465,I188468,I188471,I188474,I188520,I188523,I188526,I188529,I188532,I188535,I188538,I188541,I188544,I188547,I188593,I188596,I188599,I188602,I188605,I188608,I188611,I188614,I188617,I188663,I188666,I188669,I188672,I188675,I188678,I188681,I188684,I188687,I188733,I188736,I188739,I188742,I188745,I188748,I188751,I188754,I188757,I188803,I188806,I188809,I188812,I188815,I188818,I188821,I188824,I188827,I188830,I188876,I188879,I188882,I188885,I188888,I188891,I188894,I188897,I188900,I188946,I188949,I188952,I188955,I188958,I188961,I188964,I188967,I189013,I189016,I189019,I189022,I189025,I189028,I189031,I189034,I189037,I189040,I189086,I189089,I189092,I189095,I189098,I189101,I189104,I189107,I189110,I189113,I189159,I189162,I189165,I189168,I189171,I189174,I189177,I189180,I189183,I189229,I189232,I189235,I189238,I189241,I189244,I189247,I189250,I189253,I189299,I189302,I189305,I189308,I189311,I189314,I189317,I189320,I189323,I189369,I189372,I189375,I189378,I189381,I189384,I189387,I189390,I189393,I189396,I189442,I189445,I189448,I189451,I189454,I189457,I189460,I189463,I189466,I189512,I189515,I189518,I189521,I189524,I189527,I189530,I189533,I189579,I189582,I189585,I189588,I189591,I189594,I189597,I189600,I189603,I189649,I189652,I189655,I189658,I189661,I189664,I189667,I189670,I189673,I189676,I189722,I189725,I189728,I189731,I189734,I189737,I189740,I189743,I189789,I189792,I189795,I189798,I189801,I189804,I189807,I189810,I189813,I189859,I189862,I189865,I189868,I189871,I189874,I189877,I189880,I189883,I189886,I189932,I189935,I189938,I189941,I189944,I189947,I189950,I189953,I189956,I190002,I190005,I190008,I190011,I190014,I190017,I190020,I190023,I190026,I190072,I190075,I190078,I190081,I190084,I190087,I190090,I190093,I190096,I190099,I190145,I190148,I190151,I190154,I190157,I190160,I190163,I190166,I190169,I190215,I190218,I190221,I190224,I190227,I190230,I190233,I190236,I190239,I190242,I190288,I190291,I190294,I190297,I190300,I190303,I190306,I190309,I190312,I190315,I190361,I190364,I190367,I190370,I190373,I190376,I190379,I190382,I190385,I190431,I190434,I190437,I190440,I190443,I190446,I190449,I190452,I190455,I190501,I190504,I190507,I190510,I190513,I190516,I190519,I190522,I190525,I190571,I190574,I190577,I190580,I190583,I190586,I190589,I190592,I190595,I190641,I190644,I190647,I190650,I190653,I190656,I190659,I190662,I190665,I190711,I190714,I190717,I190720,I190723,I190726,I190729,I190732,I190735,I190738,I190784,I190787,I190790,I190793,I190796,I190799,I190802,I190805,I190808,I190854,I190857,I190860,I190863,I190866,I190869,I190872,I190875,I190878,I190881,I190927,I190930,I190933,I190936,I190939,I190942,I190945,I190948,I190994,I190997,I191000,I191003,I191006,I191009,I191012,I191015,I191061,I191064,I191067,I191070,I191073,I191076,I191079,I191082,I191085,I191088,I191134,I191137,I191140,I191143,I191146,I191149,I191152,I191155,I191158,I191204,I191207,I191210,I191213,I191216,I191219,I191222,I191225,I191228,I191274,I191277,I191280,I191283,I191286,I191289,I191292,I191295,I191298,I191344,I191347,I191350,I191353,I191356,I191359,I191362,I191365,I191411,I191414,I191417,I191420,I191423,I191426,I191429,I191432,I191435,I191481,I191484,I191487,I191490,I191493,I191496,I191499,I191502,I191505,I191551,I191554,I191557,I191560,I191563,I191566,I191569,I191572,I191575,I191578,I191624,I191627,I191630,I191633,I191636,I191639,I191642,I191645,I191648,I191694,I191697,I191700,I191703,I191706,I191709,I191712,I191715,I191718,I191721,I191767,I191770,I191773,I191776,I191779,I191782,I191785,I191788,I191791,I191837,I191840,I191843,I191846,I191849,I191852,I191855,I191858,I191861,I191907,I191910,I191913,I191916,I191919,I191922,I191925,I191928,I191931,I191977,I191980,I191983,I191986,I191989,I191992,I191995,I191998,I192001,I192047,I192050,I192053,I192056,I192059,I192062,I192065,I192068,I192071,I192074,I192120,I192123,I192126,I192129,I192132,I192135,I192138,I192141,I192144,I192190,I192193,I192196,I192199,I192202,I192205,I192208,I192211,I192257,I192260,I192263,I192266,I192269,I192272,I192275,I192278,I192324,I192327,I192330,I192333,I192336,I192339,I192342,I192345,I192348,I192351,I192397,I192400,I192403,I192406,I192409,I192412,I192415,I192418,I192421,I192467,I192470,I192473,I192476,I192479,I192482,I192485,I192488,I192491,I192537,I192540,I192543,I192546,I192549,I192552,I192555,I192558,I192561,I192564,I192610,I192613,I192616,I192619,I192622,I192625,I192628,I192631,I192634,I192637,I192683,I192686,I192689,I192692,I192695,I192698,I192701,I192704,I192750,I192753,I192756,I192759,I192762,I192765,I192768,I192771,I192774,I192777,I192823,I192826,I192829,I192832,I192835,I192838,I192841,I192844,I192847,I192893,I192896,I192899,I192902,I192905,I192908,I192911,I192914,I192917,I192963,I192966,I192969,I192972,I192975,I192978,I192981,I192984,I192987,I193033,I193036,I193039,I193042,I193045,I193048,I193051,I193054,I193057,I193060,I193106,I193109,I193112,I193115,I193118,I193121,I193124,I193127,I193130,I193176,I193179,I193182,I193185,I193188,I193191,I193194,I193197,I193200,I193246,I193249,I193252,I193255,I193258,I193261,I193264,I193267,I193270,I193316,I193319,I193322,I193325,I193328,I193331,I193334,I193337,I193383,I193386,I193389,I193392,I193395,I193398,I193401,I193404,I193407,I193410,I193456,I193459,I193462,I193465,I193468,I193471,I193474,I193477,I193480,I193526,I193529,I193532,I193535,I193538,I193541,I193544,I193547,I193550,I193596,I193599,I193602,I193605,I193608,I193611,I193614,I193617,I193620,I193666,I193669,I193672,I193675,I193678,I193681,I193684,I193687,I193690,I193736,I193739,I193742,I193745,I193748,I193751,I193754,I193757,I193760,I193806,I193809,I193812,I193815,I193818,I193821,I193824,I193827,I193873,I193876,I193879,I193882,I193885,I193888,I193891,I193894,I193897,I193943,I193946,I193949,I193952,I193955,I193958,I193961,I193964,I193967,I194013,I194016,I194019,I194022,I194025,I194028,I194031,I194034,I194037,I194083,I194086,I194089,I194092,I194095,I194098,I194101,I194104,I194107,I194110,I194156,I194159,I194162,I194165,I194168,I194171,I194174,I194177,I194223,I194226,I194229,I194232,I194235,I194238,I194241,I194244,I194247,I194250,I194296,I194299,I194302,I194305,I194308,I194311,I194314,I194317,I194320,I194366,I194369,I194372,I194375,I194378,I194381,I194384,I194387,I194433,I194436,I194439,I194442,I194445,I194448,I194451,I194454,I194457,I194460,I194506,I194509,I194512,I194515,I194518,I194521,I194524,I194527,I194530,I194576,I194579,I194582,I194585,I194588,I194591,I194594,I194597,I194600,I194646,I194649,I194652,I194655,I194658,I194661,I194664,I194667,I194713,I194716,I194719,I194722,I194725,I194728,I194731,I194734,I194737,I194740,I194786,I194789,I194792,I194795,I194798,I194801,I194804,I194807,I194810,I194856,I194859,I194862,I194865,I194868,I194871,I194874,I194877,I194880,I194926,I194929,I194932,I194935,I194938,I194941,I194944,I194947,I194950,I194953,I194999,I195002,I195005,I195008,I195011,I195014,I195017,I195020,I195023,I195069,I195072,I195075,I195078,I195081,I195084,I195087,I195090,I195093,I195139,I195142,I195145,I195148,I195151,I195154,I195157,I195160,I195163,I195209,I195212,I195215,I195218,I195221,I195224,I195227,I195230,I195276,I195279,I195282,I195285,I195288,I195291,I195294,I195297,I195300,I195346,I195349,I195352,I195355,I195358,I195361,I195364,I195367,I195370,I195416,I195419,I195422,I195425,I195428,I195431,I195434,I195437,I195440,I195486,I195489,I195492,I195495,I195498,I195501,I195504,I195507,I195510,I195513,I195559,I195562,I195565,I195568,I195571,I195574,I195577,I195580,I195583,I195629,I195632,I195635,I195638,I195641,I195644,I195647,I195650,I195653,I195699,I195702,I195705,I195708,I195711,I195714,I195717,I195720,I195723,I195769,I195772,I195775,I195778,I195781,I195784,I195787,I195790,I195793,I195839,I195842,I195845,I195848,I195851,I195854,I195857,I195860,I195863,I195909,I195912,I195915,I195918,I195921,I195924,I195927,I195930,I195933,I195979,I195982,I195985,I195988,I195991,I195994,I195997,I196000,I196003,I196049,I196052,I196055,I196058,I196061,I196064,I196067,I196070,I196073,I196076,I196122,I196125,I196128,I196131,I196134,I196137,I196140,I196143,I196146,I196149,I196195,I196198,I196201,I196204,I196207,I196210,I196213,I196216,I196219,I196265,I196268,I196271,I196274,I196277,I196280,I196283,I196286,I196289,I196335,I196338,I196341,I196344,I196347,I196350,I196353,I196356,I196359,I196362,I196408,I196411,I196414,I196417,I196420,I196423,I196426,I196429,I196432,I196435,I196481,I196484,I196487,I196490,I196493,I196496,I196499,I196502,I196505,I196508,I196554,I196557,I196560,I196563,I196566,I196569,I196572,I196575,I196578,I196581,I196627,I196630,I196633,I196636,I196639,I196642,I196645,I196648,I196651,I196697,I196700,I196703,I196706,I196709,I196712,I196715,I196718,I196721,I196767,I196770,I196773,I196776,I196779,I196782,I196785,I196788,I196791,I196837,I196840,I196843,I196846,I196849,I196852,I196855,I196858,I196861,I196907,I196910,I196913,I196916,I196919,I196922,I196925,I196928,I196931,I196934,I196980,I196983,I196986,I196989,I196992,I196995,I196998,I197001,I197004,I197050,I197053,I197056,I197059,I197062,I197065,I197068,I197071,I197074,I197120,I197123,I197126,I197129,I197132,I197135,I197138,I197141,I197144,I197147,I197193,I197196,I197199,I197202,I197205,I197208,I197211,I197214,I197217,I197220,I197266,I197269,I197272,I197275,I197278,I197281,I197284,I197287,I197290,I197293,I197339,I197342,I197345,I197348,I197351,I197354,I197357,I197360,I197363,I197409,I197412,I197415,I197418,I197421,I197424,I197427,I197430,I197476,I197479,I197482,I197485,I197488,I197491,I197494,I197497,I197500,I197503,I197549,I197552,I197555,I197558,I197561,I197564,I197567,I197570,I197573,I197619,I197622,I197625,I197628,I197631,I197634,I197637,I197640,I197643,I197646,I197692,I197695,I197698,I197701,I197704,I197707,I197710,I197713,I197716,I197762,I197765,I197768,I197771,I197774,I197777,I197780,I197783,I197786,I197832,I197835,I197838,I197841,I197844,I197847,I197850,I197853,I197856,I197902,I197905,I197908,I197911,I197914,I197917,I197920,I197923,I197926,I197972,I197975,I197978,I197981,I197984,I197987,I197990,I197993,I197996,I198042,I198045,I198048,I198051,I198054,I198057,I198060,I198063,I198109,I198112,I198115,I198118,I198121,I198124,I198127,I198130,I198133,I198136,I198182,I198185,I198188,I198191,I198194,I198197,I198200,I198203,I198206,I198209,I198255,I198258,I198261,I198264,I198267,I198270,I198273,I198276,I198279,I198325,I198328,I198331,I198334,I198337,I198340,I198343,I198346,I198349,I198395,I198398,I198401,I198404,I198407,I198410,I198413,I198416,I198419,I198465,I198468,I198471,I198474,I198477,I198480,I198483,I198486,I198489,I198535,I198538,I198541,I198544,I198547,I198550,I198553,I198556,I198559,I198562,I198608,I198611,I198614,I198617,I198620,I198623,I198626,I198629,I198632,I198678,I198681,I198684,I198687,I198690,I198693,I198696,I198699,I198702,I198705,I198751,I198754,I198757,I198760,I198763,I198766,I198769,I198772,I198818,I198821,I198824,I198827,I198830,I198833,I198836,I198839,I198842,I198888,I198891,I198894,I198897,I198900,I198903,I198906,I198909,I198912,I198915,I198961,I198964,I198967,I198970,I198973,I198976,I198979,I198982,I199028,I199031,I199034,I199037,I199040,I199043,I199046,I199049,I199052,I199098,I199101,I199104,I199107,I199110,I199113,I199116,I199119,I199122,I199125,I199171,I199174,I199177,I199180,I199183,I199186,I199189,I199192,I199195;
PAT_8 I_0 (I1385,I1817,I2073,I2121,I1465,I1697,I1905,I2009,I2025,I1721,I1617,I2271,I2274,I2277,I2280,I2283,I2286,I2289,I2292,I2295,I2224,I2231);
PAT_2 I_1 (I2274,I2289,I2295,I2271,I2283,I2286,I2274,I2292,I2277,I2280,I2271,I2341,I2344,I2347,I2350,I2353,I2356,I2359,I2362,I2365,I2224,I2231);
PAT_17 I_2 (I2341,I2341,I2353,I2344,I2347,I2359,I2356,I2365,I2344,I2350,I2362,I2411,I2414,I2417,I2420,I2423,I2426,I2429,I2432,I2435,I2438,I2224,I2231);
PAT_4 I_3 (I2420,I2411,I2429,I2426,I2438,I2435,I2414,I2411,I2417,I2423,I2432,I2484,I2487,I2490,I2493,I2496,I2499,I2502,I2505,I2508,I2224,I2231);
PAT_9 I_4 (I2505,I2487,I2490,I2499,I2502,I2484,I2493,I2487,I2508,I2484,I2496,I2554,I2557,I2560,I2563,I2566,I2569,I2572,I2575,I2578,I2224,I2231);
PAT_2 I_5 (I2569,I2572,I2563,I2578,I2554,I2557,I2560,I2557,I2575,I2566,I2554,I2624,I2627,I2630,I2633,I2636,I2639,I2642,I2645,I2648,I2224,I2231);
PAT_10 I_6 (I2624,I2642,I2639,I2627,I2630,I2645,I2636,I2624,I2633,I2648,I2627,I2694,I2697,I2700,I2703,I2706,I2709,I2712,I2715,I2224,I2231);
PAT_11 I_7 (I2703,I2706,I2715,I2709,I2712,I2694,I2694,I2700,I2697,I2697,I2700,I2761,I2764,I2767,I2770,I2773,I2776,I2779,I2782,I2785,I2788,I2224,I2231);
PAT_9 I_8 (I2767,I2779,I2770,I2782,I2761,I2764,I2773,I2761,I2776,I2785,I2788,I2834,I2837,I2840,I2843,I2846,I2849,I2852,I2855,I2858,I2224,I2231);
PAT_6 I_9 (I2852,I2834,I2846,I2855,I2834,I2843,I2840,I2858,I2849,I2837,I2837,I2904,I2907,I2910,I2913,I2916,I2919,I2922,I2925,I2928,I2931,I2224,I2231);
PAT_4 I_10 (I2904,I2919,I2907,I2910,I2913,I2904,I2931,I2922,I2925,I2916,I2928,I2977,I2980,I2983,I2986,I2989,I2992,I2995,I2998,I3001,I2224,I2231);
PAT_10 I_11 (I2977,I2977,I3001,I2980,I2986,I2995,I2992,I2980,I2998,I2983,I2989,I3047,I3050,I3053,I3056,I3059,I3062,I3065,I3068,I2224,I2231);
PAT_2 I_12 (I3059,I3062,I3053,I3065,I3050,I3047,I3047,I3053,I3068,I3056,I3050,I3114,I3117,I3120,I3123,I3126,I3129,I3132,I3135,I3138,I2224,I2231);
PAT_5 I_13 (I3135,I3114,I3114,I3126,I3123,I3132,I3120,I3129,I3138,I3117,I3117,I3184,I3187,I3190,I3193,I3196,I3199,I3202,I3205,I3208,I3211,I2224,I2231);
PAT_1 I_14 (I3199,I3187,I3205,I3184,I3190,I3184,I3193,I3208,I3202,I3211,I3196,I3257,I3260,I3263,I3266,I3269,I3272,I3275,I3278,I3281,I2224,I2231);
PAT_5 I_15 (I3275,I3278,I3260,I3269,I3266,I3263,I3272,I3281,I3260,I3257,I3257,I3327,I3330,I3333,I3336,I3339,I3342,I3345,I3348,I3351,I3354,I2224,I2231);
PAT_4 I_16 (I3345,I3351,I3354,I3333,I3336,I3348,I3330,I3327,I3339,I3342,I3327,I3400,I3403,I3406,I3409,I3412,I3415,I3418,I3421,I3424,I2224,I2231);
PAT_17 I_17 (I3412,I3409,I3421,I3415,I3400,I3418,I3424,I3403,I3406,I3403,I3400,I3470,I3473,I3476,I3479,I3482,I3485,I3488,I3491,I3494,I3497,I2224,I2231);
PAT_2 I_18 (I3470,I3488,I3485,I3470,I3479,I3494,I3491,I3476,I3497,I3482,I3473,I3543,I3546,I3549,I3552,I3555,I3558,I3561,I3564,I3567,I2224,I2231);
PAT_17 I_19 (I3543,I3543,I3555,I3546,I3549,I3561,I3558,I3567,I3546,I3552,I3564,I3613,I3616,I3619,I3622,I3625,I3628,I3631,I3634,I3637,I3640,I2224,I2231);
PAT_11 I_20 (I3625,I3634,I3640,I3616,I3613,I3631,I3622,I3628,I3619,I3637,I3613,I3686,I3689,I3692,I3695,I3698,I3701,I3704,I3707,I3710,I3713,I2224,I2231);
PAT_15 I_21 (I3710,I3689,I3695,I3704,I3701,I3686,I3698,I3707,I3686,I3692,I3713,I3759,I3762,I3765,I3768,I3771,I3774,I3777,I3780,I3783,I2224,I2231);
PAT_6 I_22 (I3762,I3759,I3765,I3780,I3762,I3783,I3768,I3774,I3771,I3777,I3759,I3829,I3832,I3835,I3838,I3841,I3844,I3847,I3850,I3853,I3856,I2224,I2231);
PAT_15 I_23 (I3847,I3838,I3850,I3853,I3844,I3856,I3829,I3835,I3829,I3832,I3841,I3902,I3905,I3908,I3911,I3914,I3917,I3920,I3923,I3926,I2224,I2231);
PAT_5 I_24 (I3905,I3902,I3908,I3926,I3923,I3911,I3920,I3914,I3905,I3917,I3902,I3972,I3975,I3978,I3981,I3984,I3987,I3990,I3993,I3996,I3999,I2224,I2231);
PAT_17 I_25 (I3999,I3975,I3978,I3981,I3972,I3984,I3972,I3996,I3990,I3987,I3993,I4045,I4048,I4051,I4054,I4057,I4060,I4063,I4066,I4069,I4072,I2224,I2231);
PAT_6 I_26 (I4045,I4063,I4051,I4054,I4060,I4045,I4057,I4048,I4069,I4072,I4066,I4118,I4121,I4124,I4127,I4130,I4133,I4136,I4139,I4142,I4145,I2224,I2231);
PAT_5 I_27 (I4139,I4118,I4124,I4127,I4133,I4136,I4118,I4142,I4121,I4130,I4145,I4191,I4194,I4197,I4200,I4203,I4206,I4209,I4212,I4215,I4218,I2224,I2231);
PAT_9 I_28 (I4206,I4203,I4212,I4209,I4200,I4191,I4197,I4218,I4194,I4215,I4191,I4264,I4267,I4270,I4273,I4276,I4279,I4282,I4285,I4288,I2224,I2231);
PAT_6 I_29 (I4282,I4264,I4276,I4285,I4264,I4273,I4270,I4288,I4279,I4267,I4267,I4334,I4337,I4340,I4343,I4346,I4349,I4352,I4355,I4358,I4361,I2224,I2231);
PAT_17 I_30 (I4346,I4349,I4355,I4343,I4337,I4358,I4352,I4334,I4361,I4340,I4334,I4407,I4410,I4413,I4416,I4419,I4422,I4425,I4428,I4431,I4434,I2224,I2231);
PAT_10 I_31 (I4407,I4413,I4434,I4416,I4431,I4410,I4425,I4419,I4428,I4422,I4407,I4480,I4483,I4486,I4489,I4492,I4495,I4498,I4501,I2224,I2231);
PAT_9 I_32 (I4492,I4480,I4483,I4486,I4480,I4486,I4489,I4483,I4501,I4495,I4498,I4547,I4550,I4553,I4556,I4559,I4562,I4565,I4568,I4571,I2224,I2231);
PAT_0 I_33 (I4556,I4568,I4547,I4550,I4553,I4547,I4562,I4565,I4559,I4571,I4550,I4617,I4620,I4623,I4626,I4629,I4632,I4635,I4638,I2224,I2231);
PAT_4 I_34 (I4626,I4617,I4623,I4638,I4620,I4629,I4617,I4620,I4623,I4632,I4635,I4684,I4687,I4690,I4693,I4696,I4699,I4702,I4705,I4708,I2224,I2231);
PAT_12 I_35 (I4684,I4687,I4705,I4708,I4699,I4690,I4696,I4693,I4684,I4702,I4687,I4754,I4757,I4760,I4763,I4766,I4769,I4772,I4775,I2224,I2231);
PAT_1 I_36 (I4769,I4757,I4772,I4763,I4754,I4757,I4766,I4754,I4775,I4760,I4760,I4821,I4824,I4827,I4830,I4833,I4836,I4839,I4842,I4845,I2224,I2231);
PAT_12 I_37 (I4833,I4827,I4845,I4821,I4830,I4821,I4824,I4842,I4836,I4824,I4839,I4891,I4894,I4897,I4900,I4903,I4906,I4909,I4912,I2224,I2231);
PAT_8 I_38 (I4891,I4900,I4897,I4894,I4906,I4891,I4894,I4897,I4909,I4903,I4912,I4958,I4961,I4964,I4967,I4970,I4973,I4976,I4979,I4982,I2224,I2231);
PAT_11 I_39 (I4979,I4970,I4958,I4961,I4976,I4964,I4967,I4958,I4982,I4973,I4961,I5028,I5031,I5034,I5037,I5040,I5043,I5046,I5049,I5052,I5055,I2224,I2231);
PAT_10 I_40 (I5043,I5049,I5040,I5034,I5052,I5037,I5055,I5046,I5028,I5031,I5028,I5101,I5104,I5107,I5110,I5113,I5116,I5119,I5122,I2224,I2231);
PAT_11 I_41 (I5110,I5113,I5122,I5116,I5119,I5101,I5101,I5107,I5104,I5104,I5107,I5168,I5171,I5174,I5177,I5180,I5183,I5186,I5189,I5192,I5195,I2224,I2231);
PAT_5 I_42 (I5189,I5168,I5195,I5183,I5180,I5192,I5174,I5168,I5186,I5171,I5177,I5241,I5244,I5247,I5250,I5253,I5256,I5259,I5262,I5265,I5268,I2224,I2231);
PAT_11 I_43 (I5253,I5250,I5244,I5262,I5265,I5241,I5259,I5256,I5268,I5247,I5241,I5314,I5317,I5320,I5323,I5326,I5329,I5332,I5335,I5338,I5341,I2224,I2231);
PAT_15 I_44 (I5338,I5317,I5323,I5332,I5329,I5314,I5326,I5335,I5314,I5320,I5341,I5387,I5390,I5393,I5396,I5399,I5402,I5405,I5408,I5411,I2224,I2231);
PAT_6 I_45 (I5390,I5387,I5393,I5408,I5390,I5411,I5396,I5402,I5399,I5405,I5387,I5457,I5460,I5463,I5466,I5469,I5472,I5475,I5478,I5481,I5484,I2224,I2231);
PAT_8 I_46 (I5466,I5472,I5463,I5475,I5457,I5460,I5478,I5457,I5484,I5481,I5469,I5530,I5533,I5536,I5539,I5542,I5545,I5548,I5551,I5554,I2224,I2231);
PAT_5 I_47 (I5536,I5554,I5530,I5551,I5539,I5542,I5533,I5530,I5533,I5545,I5548,I5600,I5603,I5606,I5609,I5612,I5615,I5618,I5621,I5624,I5627,I2224,I2231);
PAT_12 I_48 (I5627,I5615,I5600,I5624,I5603,I5600,I5606,I5609,I5612,I5618,I5621,I5673,I5676,I5679,I5682,I5685,I5688,I5691,I5694,I2224,I2231);
PAT_17 I_49 (I5688,I5682,I5676,I5673,I5673,I5679,I5679,I5691,I5694,I5676,I5685,I5740,I5743,I5746,I5749,I5752,I5755,I5758,I5761,I5764,I5767,I2224,I2231);
PAT_4 I_50 (I5749,I5740,I5758,I5755,I5767,I5764,I5743,I5740,I5746,I5752,I5761,I5813,I5816,I5819,I5822,I5825,I5828,I5831,I5834,I5837,I2224,I2231);
PAT_2 I_51 (I5822,I5816,I5816,I5837,I5813,I5831,I5828,I5819,I5813,I5825,I5834,I5883,I5886,I5889,I5892,I5895,I5898,I5901,I5904,I5907,I2224,I2231);
PAT_9 I_52 (I5898,I5907,I5883,I5889,I5892,I5901,I5886,I5895,I5904,I5886,I5883,I5953,I5956,I5959,I5962,I5965,I5968,I5971,I5974,I5977,I2224,I2231);
PAT_13 I_53 (I5953,I5974,I5956,I5971,I5965,I5962,I5977,I5953,I5959,I5968,I5956,I6023,I6026,I6029,I6032,I6035,I6038,I6041,I6044,I6047,I2224,I2231);
PAT_12 I_54 (I6032,I6023,I6023,I6047,I6044,I6026,I6041,I6035,I6026,I6029,I6038,I6093,I6096,I6099,I6102,I6105,I6108,I6111,I6114,I2224,I2231);
PAT_10 I_55 (I6093,I6114,I6105,I6108,I6099,I6096,I6093,I6111,I6099,I6102,I6096,I6160,I6163,I6166,I6169,I6172,I6175,I6178,I6181,I2224,I2231);
PAT_14 I_56 (I6160,I6181,I6166,I6175,I6172,I6178,I6169,I6163,I6163,I6166,I6160,I6227,I6230,I6233,I6236,I6239,I6242,I6245,I6248,I6251,I2224,I2231);
PAT_9 I_57 (I6236,I6248,I6227,I6245,I6230,I6233,I6251,I6230,I6239,I6227,I6242,I6297,I6300,I6303,I6306,I6309,I6312,I6315,I6318,I6321,I2224,I2231);
PAT_1 I_58 (I6297,I6315,I6297,I6309,I6300,I6306,I6312,I6318,I6321,I6303,I6300,I6367,I6370,I6373,I6376,I6379,I6382,I6385,I6388,I6391,I2224,I2231);
PAT_8 I_59 (I6388,I6370,I6376,I6367,I6385,I6379,I6382,I6367,I6391,I6373,I6370,I6437,I6440,I6443,I6446,I6449,I6452,I6455,I6458,I6461,I2224,I2231);
PAT_13 I_60 (I6449,I6458,I6440,I6461,I6443,I6437,I6437,I6446,I6455,I6452,I6440,I6507,I6510,I6513,I6516,I6519,I6522,I6525,I6528,I6531,I2224,I2231);
PAT_9 I_61 (I6528,I6510,I6510,I6507,I6531,I6513,I6516,I6507,I6519,I6525,I6522,I6577,I6580,I6583,I6586,I6589,I6592,I6595,I6598,I6601,I2224,I2231);
PAT_8 I_62 (I6598,I6586,I6595,I6577,I6580,I6592,I6601,I6580,I6583,I6589,I6577,I6647,I6650,I6653,I6656,I6659,I6662,I6665,I6668,I6671,I2224,I2231);
PAT_11 I_63 (I6668,I6659,I6647,I6650,I6665,I6653,I6656,I6647,I6671,I6662,I6650,I6717,I6720,I6723,I6726,I6729,I6732,I6735,I6738,I6741,I6744,I2224,I2231);
PAT_10 I_64 (I6732,I6738,I6729,I6723,I6741,I6726,I6744,I6735,I6717,I6720,I6717,I6790,I6793,I6796,I6799,I6802,I6805,I6808,I6811,I2224,I2231);
PAT_6 I_65 (I6811,I6805,I6799,I6793,I6790,I6796,I6790,I6796,I6793,I6802,I6808,I6857,I6860,I6863,I6866,I6869,I6872,I6875,I6878,I6881,I6884,I2224,I2231);
PAT_14 I_66 (I6869,I6863,I6857,I6884,I6866,I6860,I6872,I6875,I6857,I6881,I6878,I6930,I6933,I6936,I6939,I6942,I6945,I6948,I6951,I6954,I2224,I2231);
PAT_5 I_67 (I6933,I6936,I6933,I6942,I6930,I6951,I6939,I6930,I6954,I6948,I6945,I7000,I7003,I7006,I7009,I7012,I7015,I7018,I7021,I7024,I7027,I2224,I2231);
PAT_10 I_68 (I7024,I7027,I7006,I7012,I7015,I7021,I7003,I7000,I7000,I7009,I7018,I7073,I7076,I7079,I7082,I7085,I7088,I7091,I7094,I2224,I2231);
PAT_7 I_69 (I7094,I7091,I7088,I7073,I7076,I7079,I7076,I7085,I7073,I7079,I7082,I7140,I7143,I7146,I7149,I7152,I7155,I7158,I7161,I7164,I2224,I2231);
PAT_13 I_70 (I7146,I7164,I7155,I7140,I7152,I7140,I7161,I7143,I7149,I7143,I7158,I7210,I7213,I7216,I7219,I7222,I7225,I7228,I7231,I7234,I2224,I2231);
PAT_7 I_71 (I7219,I7222,I7210,I7225,I7231,I7216,I7213,I7234,I7213,I7210,I7228,I7280,I7283,I7286,I7289,I7292,I7295,I7298,I7301,I7304,I2224,I2231);
PAT_13 I_72 (I7286,I7304,I7295,I7280,I7292,I7280,I7301,I7283,I7289,I7283,I7298,I7350,I7353,I7356,I7359,I7362,I7365,I7368,I7371,I7374,I2224,I2231);
PAT_14 I_73 (I7353,I7368,I7356,I7365,I7359,I7350,I7362,I7371,I7350,I7374,I7353,I7420,I7423,I7426,I7429,I7432,I7435,I7438,I7441,I7444,I2224,I2231);
PAT_11 I_74 (I7432,I7429,I7426,I7420,I7423,I7423,I7435,I7420,I7441,I7444,I7438,I7490,I7493,I7496,I7499,I7502,I7505,I7508,I7511,I7514,I7517,I2224,I2231);
PAT_9 I_75 (I7496,I7508,I7499,I7511,I7490,I7493,I7502,I7490,I7505,I7514,I7517,I7563,I7566,I7569,I7572,I7575,I7578,I7581,I7584,I7587,I2224,I2231);
PAT_12 I_76 (I7584,I7581,I7575,I7563,I7572,I7563,I7566,I7569,I7587,I7578,I7566,I7633,I7636,I7639,I7642,I7645,I7648,I7651,I7654,I2224,I2231);
PAT_15 I_77 (I7654,I7636,I7633,I7633,I7648,I7651,I7645,I7636,I7639,I7642,I7639,I7700,I7703,I7706,I7709,I7712,I7715,I7718,I7721,I7724,I2224,I2231);
PAT_9 I_78 (I7700,I7721,I7709,I7703,I7715,I7703,I7718,I7724,I7706,I7700,I7712,I7770,I7773,I7776,I7779,I7782,I7785,I7788,I7791,I7794,I2224,I2231);
PAT_11 I_79 (I7782,I7788,I7794,I7791,I7779,I7773,I7773,I7770,I7785,I7770,I7776,I7840,I7843,I7846,I7849,I7852,I7855,I7858,I7861,I7864,I7867,I2224,I2231);
PAT_5 I_80 (I7861,I7840,I7867,I7855,I7852,I7864,I7846,I7840,I7858,I7843,I7849,I7913,I7916,I7919,I7922,I7925,I7928,I7931,I7934,I7937,I7940,I2224,I2231);
PAT_11 I_81 (I7925,I7922,I7916,I7934,I7937,I7913,I7931,I7928,I7940,I7919,I7913,I7986,I7989,I7992,I7995,I7998,I8001,I8004,I8007,I8010,I8013,I2224,I2231);
PAT_8 I_82 (I7995,I8001,I8004,I8010,I8007,I7998,I7986,I7986,I8013,I7989,I7992,I8059,I8062,I8065,I8068,I8071,I8074,I8077,I8080,I8083,I2224,I2231);
PAT_17 I_83 (I8083,I8071,I8068,I8062,I8065,I8077,I8059,I8062,I8059,I8074,I8080,I8129,I8132,I8135,I8138,I8141,I8144,I8147,I8150,I8153,I8156,I2224,I2231);
PAT_15 I_84 (I8156,I8150,I8147,I8129,I8138,I8135,I8141,I8132,I8129,I8153,I8144,I8202,I8205,I8208,I8211,I8214,I8217,I8220,I8223,I8226,I2224,I2231);
PAT_13 I_85 (I8211,I8202,I8220,I8205,I8205,I8223,I8214,I8202,I8217,I8226,I8208,I8272,I8275,I8278,I8281,I8284,I8287,I8290,I8293,I8296,I2224,I2231);
PAT_2 I_86 (I8290,I8284,I8281,I8287,I8272,I8296,I8275,I8293,I8272,I8278,I8275,I8342,I8345,I8348,I8351,I8354,I8357,I8360,I8363,I8366,I2224,I2231);
PAT_17 I_87 (I8342,I8342,I8354,I8345,I8348,I8360,I8357,I8366,I8345,I8351,I8363,I8412,I8415,I8418,I8421,I8424,I8427,I8430,I8433,I8436,I8439,I2224,I2231);
PAT_1 I_88 (I8436,I8439,I8418,I8427,I8412,I8433,I8424,I8415,I8421,I8412,I8430,I8485,I8488,I8491,I8494,I8497,I8500,I8503,I8506,I8509,I2224,I2231);
PAT_6 I_89 (I8494,I8485,I8488,I8491,I8506,I8509,I8503,I8485,I8500,I8497,I8488,I8555,I8558,I8561,I8564,I8567,I8570,I8573,I8576,I8579,I8582,I2224,I2231);
PAT_17 I_90 (I8567,I8570,I8576,I8564,I8558,I8579,I8573,I8555,I8582,I8561,I8555,I8628,I8631,I8634,I8637,I8640,I8643,I8646,I8649,I8652,I8655,I2224,I2231);
PAT_4 I_91 (I8637,I8628,I8646,I8643,I8655,I8652,I8631,I8628,I8634,I8640,I8649,I8701,I8704,I8707,I8710,I8713,I8716,I8719,I8722,I8725,I2224,I2231);
PAT_13 I_92 (I8716,I8710,I8722,I8707,I8713,I8701,I8725,I8719,I8704,I8701,I8704,I8771,I8774,I8777,I8780,I8783,I8786,I8789,I8792,I8795,I2224,I2231);
PAT_11 I_93 (I8771,I8783,I8786,I8777,I8774,I8795,I8774,I8792,I8780,I8771,I8789,I8841,I8844,I8847,I8850,I8853,I8856,I8859,I8862,I8865,I8868,I2224,I2231);
PAT_6 I_94 (I8841,I8868,I8856,I8865,I8859,I8853,I8844,I8862,I8850,I8847,I8841,I8914,I8917,I8920,I8923,I8926,I8929,I8932,I8935,I8938,I8941,I2224,I2231);
PAT_17 I_95 (I8926,I8929,I8935,I8923,I8917,I8938,I8932,I8914,I8941,I8920,I8914,I8987,I8990,I8993,I8996,I8999,I9002,I9005,I9008,I9011,I9014,I2224,I2231);
PAT_8 I_96 (I8996,I9008,I9014,I9005,I8990,I8999,I9002,I9011,I8993,I8987,I8987,I9060,I9063,I9066,I9069,I9072,I9075,I9078,I9081,I9084,I2224,I2231);
PAT_4 I_97 (I9078,I9063,I9069,I9060,I9060,I9072,I9063,I9081,I9084,I9066,I9075,I9130,I9133,I9136,I9139,I9142,I9145,I9148,I9151,I9154,I2224,I2231);
PAT_12 I_98 (I9130,I9133,I9151,I9154,I9145,I9136,I9142,I9139,I9130,I9148,I9133,I9200,I9203,I9206,I9209,I9212,I9215,I9218,I9221,I2224,I2231);
PAT_5 I_99 (I9209,I9215,I9221,I9206,I9206,I9200,I9218,I9200,I9203,I9203,I9212,I9267,I9270,I9273,I9276,I9279,I9282,I9285,I9288,I9291,I9294,I2224,I2231);
PAT_7 I_100 (I9285,I9288,I9294,I9291,I9276,I9273,I9267,I9279,I9267,I9270,I9282,I9340,I9343,I9346,I9349,I9352,I9355,I9358,I9361,I9364,I2224,I2231);
PAT_2 I_101 (I9361,I9355,I9346,I9340,I9349,I9343,I9352,I9364,I9358,I9343,I9340,I9410,I9413,I9416,I9419,I9422,I9425,I9428,I9431,I9434,I2224,I2231);
PAT_17 I_102 (I9410,I9410,I9422,I9413,I9416,I9428,I9425,I9434,I9413,I9419,I9431,I9480,I9483,I9486,I9489,I9492,I9495,I9498,I9501,I9504,I9507,I2224,I2231);
PAT_15 I_103 (I9507,I9501,I9498,I9480,I9489,I9486,I9492,I9483,I9480,I9504,I9495,I9553,I9556,I9559,I9562,I9565,I9568,I9571,I9574,I9577,I2224,I2231);
PAT_13 I_104 (I9562,I9553,I9571,I9556,I9556,I9574,I9565,I9553,I9568,I9577,I9559,I9623,I9626,I9629,I9632,I9635,I9638,I9641,I9644,I9647,I2224,I2231);
PAT_9 I_105 (I9644,I9626,I9626,I9623,I9647,I9629,I9632,I9623,I9635,I9641,I9638,I9693,I9696,I9699,I9702,I9705,I9708,I9711,I9714,I9717,I2224,I2231);
PAT_13 I_106 (I9693,I9714,I9696,I9711,I9705,I9702,I9717,I9693,I9699,I9708,I9696,I9763,I9766,I9769,I9772,I9775,I9778,I9781,I9784,I9787,I2224,I2231);
PAT_2 I_107 (I9781,I9775,I9772,I9778,I9763,I9787,I9766,I9784,I9763,I9769,I9766,I9833,I9836,I9839,I9842,I9845,I9848,I9851,I9854,I9857,I2224,I2231);
PAT_13 I_108 (I9842,I9836,I9833,I9854,I9845,I9848,I9836,I9839,I9851,I9857,I9833,I9903,I9906,I9909,I9912,I9915,I9918,I9921,I9924,I9927,I2224,I2231);
PAT_9 I_109 (I9924,I9906,I9906,I9903,I9927,I9909,I9912,I9903,I9915,I9921,I9918,I9973,I9976,I9979,I9982,I9985,I9988,I9991,I9994,I9997,I2224,I2231);
PAT_11 I_110 (I9985,I9991,I9997,I9994,I9982,I9976,I9976,I9973,I9988,I9973,I9979,I10043,I10046,I10049,I10052,I10055,I10058,I10061,I10064,I10067,I10070,I2224,I2231);
PAT_9 I_111 (I10049,I10061,I10052,I10064,I10043,I10046,I10055,I10043,I10058,I10067,I10070,I10116,I10119,I10122,I10125,I10128,I10131,I10134,I10137,I10140,I2224,I2231);
PAT_5 I_112 (I10137,I10116,I10131,I10116,I10122,I10125,I10119,I10119,I10134,I10128,I10140,I10186,I10189,I10192,I10195,I10198,I10201,I10204,I10207,I10210,I10213,I2224,I2231);
PAT_2 I_113 (I10201,I10186,I10198,I10192,I10207,I10189,I10204,I10195,I10210,I10213,I10186,I10259,I10262,I10265,I10268,I10271,I10274,I10277,I10280,I10283,I2224,I2231);
PAT_9 I_114 (I10274,I10283,I10259,I10265,I10268,I10277,I10262,I10271,I10280,I10262,I10259,I10329,I10332,I10335,I10338,I10341,I10344,I10347,I10350,I10353,I2224,I2231);
PAT_13 I_115 (I10329,I10350,I10332,I10347,I10341,I10338,I10353,I10329,I10335,I10344,I10332,I10399,I10402,I10405,I10408,I10411,I10414,I10417,I10420,I10423,I2224,I2231);
PAT_2 I_116 (I10417,I10411,I10408,I10414,I10399,I10423,I10402,I10420,I10399,I10405,I10402,I10469,I10472,I10475,I10478,I10481,I10484,I10487,I10490,I10493,I2224,I2231);
PAT_10 I_117 (I10469,I10487,I10484,I10472,I10475,I10490,I10481,I10469,I10478,I10493,I10472,I10539,I10542,I10545,I10548,I10551,I10554,I10557,I10560,I2224,I2231);
PAT_5 I_118 (I10560,I10539,I10548,I10542,I10557,I10554,I10545,I10545,I10539,I10542,I10551,I10606,I10609,I10612,I10615,I10618,I10621,I10624,I10627,I10630,I10633,I2224,I2231);
PAT_9 I_119 (I10621,I10618,I10627,I10624,I10615,I10606,I10612,I10633,I10609,I10630,I10606,I10679,I10682,I10685,I10688,I10691,I10694,I10697,I10700,I10703,I2224,I2231);
PAT_5 I_120 (I10700,I10679,I10694,I10679,I10685,I10688,I10682,I10682,I10697,I10691,I10703,I10749,I10752,I10755,I10758,I10761,I10764,I10767,I10770,I10773,I10776,I2224,I2231);
PAT_3 I_121 (I10761,I10749,I10776,I10770,I10773,I10749,I10764,I10752,I10755,I10758,I10767,I10822,I10825,I10828,I10831,I10834,I10837,I10840,I10843,I10846,I10849,I2224,I2231);
PAT_13 I_122 (I10843,I10831,I10849,I10828,I10834,I10837,I10825,I10840,I10822,I10822,I10846,I10895,I10898,I10901,I10904,I10907,I10910,I10913,I10916,I10919,I2224,I2231);
PAT_9 I_123 (I10916,I10898,I10898,I10895,I10919,I10901,I10904,I10895,I10907,I10913,I10910,I10965,I10968,I10971,I10974,I10977,I10980,I10983,I10986,I10989,I2224,I2231);
PAT_6 I_124 (I10983,I10965,I10977,I10986,I10965,I10974,I10971,I10989,I10980,I10968,I10968,I11035,I11038,I11041,I11044,I11047,I11050,I11053,I11056,I11059,I11062,I2224,I2231);
PAT_13 I_125 (I11059,I11041,I11056,I11035,I11038,I11044,I11062,I11047,I11053,I11035,I11050,I11108,I11111,I11114,I11117,I11120,I11123,I11126,I11129,I11132,I2224,I2231);
PAT_5 I_126 (I11120,I11111,I11117,I11129,I11111,I11132,I11114,I11123,I11108,I11108,I11126,I11178,I11181,I11184,I11187,I11190,I11193,I11196,I11199,I11202,I11205,I2224,I2231);
PAT_11 I_127 (I11190,I11187,I11181,I11199,I11202,I11178,I11196,I11193,I11205,I11184,I11178,I11251,I11254,I11257,I11260,I11263,I11266,I11269,I11272,I11275,I11278,I2224,I2231);
PAT_5 I_128 (I11272,I11251,I11278,I11266,I11263,I11275,I11257,I11251,I11269,I11254,I11260,I11324,I11327,I11330,I11333,I11336,I11339,I11342,I11345,I11348,I11351,I2224,I2231);
PAT_2 I_129 (I11339,I11324,I11336,I11330,I11345,I11327,I11342,I11333,I11348,I11351,I11324,I11397,I11400,I11403,I11406,I11409,I11412,I11415,I11418,I11421,I2224,I2231);
PAT_12 I_130 (I11406,I11403,I11397,I11400,I11421,I11415,I11418,I11400,I11412,I11397,I11409,I11467,I11470,I11473,I11476,I11479,I11482,I11485,I11488,I2224,I2231);
PAT_13 I_131 (I11479,I11482,I11473,I11488,I11485,I11467,I11470,I11476,I11473,I11470,I11467,I11534,I11537,I11540,I11543,I11546,I11549,I11552,I11555,I11558,I2224,I2231);
PAT_10 I_132 (I11555,I11549,I11543,I11537,I11558,I11537,I11546,I11534,I11534,I11552,I11540,I11604,I11607,I11610,I11613,I11616,I11619,I11622,I11625,I2224,I2231);
PAT_7 I_133 (I11625,I11622,I11619,I11604,I11607,I11610,I11607,I11616,I11604,I11610,I11613,I11671,I11674,I11677,I11680,I11683,I11686,I11689,I11692,I11695,I2224,I2231);
PAT_6 I_134 (I11671,I11689,I11671,I11680,I11686,I11674,I11692,I11677,I11695,I11674,I11683,I11741,I11744,I11747,I11750,I11753,I11756,I11759,I11762,I11765,I11768,I2224,I2231);
PAT_7 I_135 (I11747,I11756,I11759,I11741,I11750,I11744,I11753,I11768,I11762,I11765,I11741,I11814,I11817,I11820,I11823,I11826,I11829,I11832,I11835,I11838,I2224,I2231);
PAT_2 I_136 (I11835,I11829,I11820,I11814,I11823,I11817,I11826,I11838,I11832,I11817,I11814,I11884,I11887,I11890,I11893,I11896,I11899,I11902,I11905,I11908,I2224,I2231);
PAT_17 I_137 (I11884,I11884,I11896,I11887,I11890,I11902,I11899,I11908,I11887,I11893,I11905,I11954,I11957,I11960,I11963,I11966,I11969,I11972,I11975,I11978,I11981,I2224,I2231);
PAT_5 I_138 (I11966,I11960,I11957,I11978,I11963,I11969,I11972,I11954,I11954,I11975,I11981,I12027,I12030,I12033,I12036,I12039,I12042,I12045,I12048,I12051,I12054,I2224,I2231);
PAT_9 I_139 (I12042,I12039,I12048,I12045,I12036,I12027,I12033,I12054,I12030,I12051,I12027,I12100,I12103,I12106,I12109,I12112,I12115,I12118,I12121,I12124,I2224,I2231);
PAT_2 I_140 (I12115,I12118,I12109,I12124,I12100,I12103,I12106,I12103,I12121,I12112,I12100,I12170,I12173,I12176,I12179,I12182,I12185,I12188,I12191,I12194,I2224,I2231);
PAT_13 I_141 (I12179,I12173,I12170,I12191,I12182,I12185,I12173,I12176,I12188,I12194,I12170,I12240,I12243,I12246,I12249,I12252,I12255,I12258,I12261,I12264,I2224,I2231);
PAT_16 I_142 (I12246,I12249,I12258,I12252,I12264,I12240,I12261,I12255,I12243,I12243,I12240,I12310,I12313,I12316,I12319,I12322,I12325,I12328,I12331,I12334,I12337,I2224,I2231);
PAT_5 I_143 (I12328,I12331,I12319,I12325,I12316,I12310,I12334,I12337,I12313,I12310,I12322,I12383,I12386,I12389,I12392,I12395,I12398,I12401,I12404,I12407,I12410,I2224,I2231);
PAT_9 I_144 (I12398,I12395,I12404,I12401,I12392,I12383,I12389,I12410,I12386,I12407,I12383,I12456,I12459,I12462,I12465,I12468,I12471,I12474,I12477,I12480,I2224,I2231);
PAT_2 I_145 (I12471,I12474,I12465,I12480,I12456,I12459,I12462,I12459,I12477,I12468,I12456,I12526,I12529,I12532,I12535,I12538,I12541,I12544,I12547,I12550,I2224,I2231);
PAT_5 I_146 (I12547,I12526,I12526,I12538,I12535,I12544,I12532,I12541,I12550,I12529,I12529,I12596,I12599,I12602,I12605,I12608,I12611,I12614,I12617,I12620,I12623,I2224,I2231);
PAT_16 I_147 (I12614,I12608,I12620,I12623,I12602,I12596,I12599,I12611,I12605,I12617,I12596,I12669,I12672,I12675,I12678,I12681,I12684,I12687,I12690,I12693,I12696,I2224,I2231);
PAT_6 I_148 (I12669,I12672,I12681,I12687,I12675,I12696,I12678,I12690,I12693,I12684,I12669,I12742,I12745,I12748,I12751,I12754,I12757,I12760,I12763,I12766,I12769,I2224,I2231);
PAT_4 I_149 (I12742,I12757,I12745,I12748,I12751,I12742,I12769,I12760,I12763,I12754,I12766,I12815,I12818,I12821,I12824,I12827,I12830,I12833,I12836,I12839,I2224,I2231);
PAT_11 I_150 (I12827,I12836,I12818,I12830,I12815,I12818,I12815,I12824,I12839,I12833,I12821,I12885,I12888,I12891,I12894,I12897,I12900,I12903,I12906,I12909,I12912,I2224,I2231);
PAT_15 I_151 (I12909,I12888,I12894,I12903,I12900,I12885,I12897,I12906,I12885,I12891,I12912,I12958,I12961,I12964,I12967,I12970,I12973,I12976,I12979,I12982,I2224,I2231);
PAT_10 I_152 (I12961,I12970,I12964,I12958,I12979,I12982,I12967,I12958,I12961,I12976,I12973,I13028,I13031,I13034,I13037,I13040,I13043,I13046,I13049,I2224,I2231);
PAT_13 I_153 (I13034,I13040,I13034,I13031,I13046,I13049,I13028,I13028,I13043,I13031,I13037,I13095,I13098,I13101,I13104,I13107,I13110,I13113,I13116,I13119,I2224,I2231);
PAT_17 I_154 (I13119,I13107,I13116,I13113,I13104,I13095,I13098,I13101,I13095,I13110,I13098,I13165,I13168,I13171,I13174,I13177,I13180,I13183,I13186,I13189,I13192,I2224,I2231);
PAT_13 I_155 (I13183,I13186,I13171,I13165,I13177,I13189,I13168,I13180,I13165,I13192,I13174,I13238,I13241,I13244,I13247,I13250,I13253,I13256,I13259,I13262,I2224,I2231);
PAT_10 I_156 (I13259,I13253,I13247,I13241,I13262,I13241,I13250,I13238,I13238,I13256,I13244,I13308,I13311,I13314,I13317,I13320,I13323,I13326,I13329,I2224,I2231);
PAT_8 I_157 (I13329,I13320,I13311,I13308,I13317,I13308,I13323,I13311,I13326,I13314,I13314,I13375,I13378,I13381,I13384,I13387,I13390,I13393,I13396,I13399,I2224,I2231);
PAT_11 I_158 (I13396,I13387,I13375,I13378,I13393,I13381,I13384,I13375,I13399,I13390,I13378,I13445,I13448,I13451,I13454,I13457,I13460,I13463,I13466,I13469,I13472,I2224,I2231);
PAT_2 I_159 (I13445,I13469,I13457,I13451,I13460,I13463,I13448,I13472,I13466,I13454,I13445,I13518,I13521,I13524,I13527,I13530,I13533,I13536,I13539,I13542,I2224,I2231);
PAT_10 I_160 (I13518,I13536,I13533,I13521,I13524,I13539,I13530,I13518,I13527,I13542,I13521,I13588,I13591,I13594,I13597,I13600,I13603,I13606,I13609,I2224,I2231);
PAT_13 I_161 (I13594,I13600,I13594,I13591,I13606,I13609,I13588,I13588,I13603,I13591,I13597,I13655,I13658,I13661,I13664,I13667,I13670,I13673,I13676,I13679,I2224,I2231);
PAT_6 I_162 (I13655,I13667,I13664,I13676,I13673,I13679,I13655,I13670,I13658,I13658,I13661,I13725,I13728,I13731,I13734,I13737,I13740,I13743,I13746,I13749,I13752,I2224,I2231);
PAT_1 I_163 (I13752,I13743,I13731,I13734,I13746,I13737,I13740,I13725,I13728,I13725,I13749,I13798,I13801,I13804,I13807,I13810,I13813,I13816,I13819,I13822,I2224,I2231);
PAT_3 I_164 (I13807,I13801,I13801,I13804,I13816,I13819,I13822,I13810,I13798,I13798,I13813,I13868,I13871,I13874,I13877,I13880,I13883,I13886,I13889,I13892,I13895,I2224,I2231);
PAT_14 I_165 (I13874,I13871,I13877,I13889,I13883,I13892,I13880,I13868,I13886,I13895,I13868,I13941,I13944,I13947,I13950,I13953,I13956,I13959,I13962,I13965,I2224,I2231);
PAT_11 I_166 (I13953,I13950,I13947,I13941,I13944,I13944,I13956,I13941,I13962,I13965,I13959,I14011,I14014,I14017,I14020,I14023,I14026,I14029,I14032,I14035,I14038,I2224,I2231);
PAT_12 I_167 (I14020,I14035,I14017,I14014,I14023,I14026,I14032,I14011,I14029,I14038,I14011,I14084,I14087,I14090,I14093,I14096,I14099,I14102,I14105,I2224,I2231);
PAT_17 I_168 (I14099,I14093,I14087,I14084,I14084,I14090,I14090,I14102,I14105,I14087,I14096,I14151,I14154,I14157,I14160,I14163,I14166,I14169,I14172,I14175,I14178,I2224,I2231);
PAT_8 I_169 (I14160,I14172,I14178,I14169,I14154,I14163,I14166,I14175,I14157,I14151,I14151,I14224,I14227,I14230,I14233,I14236,I14239,I14242,I14245,I14248,I2224,I2231);
PAT_13 I_170 (I14236,I14245,I14227,I14248,I14230,I14224,I14224,I14233,I14242,I14239,I14227,I14294,I14297,I14300,I14303,I14306,I14309,I14312,I14315,I14318,I2224,I2231);
PAT_6 I_171 (I14294,I14306,I14303,I14315,I14312,I14318,I14294,I14309,I14297,I14297,I14300,I14364,I14367,I14370,I14373,I14376,I14379,I14382,I14385,I14388,I14391,I2224,I2231);
PAT_10 I_172 (I14364,I14379,I14382,I14373,I14364,I14388,I14391,I14367,I14376,I14370,I14385,I14437,I14440,I14443,I14446,I14449,I14452,I14455,I14458,I2224,I2231);
PAT_5 I_173 (I14458,I14437,I14446,I14440,I14455,I14452,I14443,I14443,I14437,I14440,I14449,I14504,I14507,I14510,I14513,I14516,I14519,I14522,I14525,I14528,I14531,I2224,I2231);
PAT_6 I_174 (I14522,I14516,I14504,I14510,I14507,I14513,I14519,I14504,I14528,I14525,I14531,I14577,I14580,I14583,I14586,I14589,I14592,I14595,I14598,I14601,I14604,I2224,I2231);
PAT_9 I_175 (I14577,I14604,I14601,I14583,I14589,I14580,I14592,I14577,I14595,I14586,I14598,I14650,I14653,I14656,I14659,I14662,I14665,I14668,I14671,I14674,I2224,I2231);
PAT_4 I_176 (I14650,I14674,I14668,I14656,I14653,I14671,I14653,I14650,I14665,I14659,I14662,I14720,I14723,I14726,I14729,I14732,I14735,I14738,I14741,I14744,I2224,I2231);
PAT_2 I_177 (I14729,I14723,I14723,I14744,I14720,I14738,I14735,I14726,I14720,I14732,I14741,I14790,I14793,I14796,I14799,I14802,I14805,I14808,I14811,I14814,I2224,I2231);
PAT_12 I_178 (I14799,I14796,I14790,I14793,I14814,I14808,I14811,I14793,I14805,I14790,I14802,I14860,I14863,I14866,I14869,I14872,I14875,I14878,I14881,I2224,I2231);
PAT_15 I_179 (I14881,I14863,I14860,I14860,I14875,I14878,I14872,I14863,I14866,I14869,I14866,I14927,I14930,I14933,I14936,I14939,I14942,I14945,I14948,I14951,I2224,I2231);
PAT_5 I_180 (I14930,I14927,I14933,I14951,I14948,I14936,I14945,I14939,I14930,I14942,I14927,I14997,I15000,I15003,I15006,I15009,I15012,I15015,I15018,I15021,I15024,I2224,I2231);
PAT_3 I_181 (I15009,I14997,I15024,I15018,I15021,I14997,I15012,I15000,I15003,I15006,I15015,I15070,I15073,I15076,I15079,I15082,I15085,I15088,I15091,I15094,I15097,I2224,I2231);
PAT_13 I_182 (I15091,I15079,I15097,I15076,I15082,I15085,I15073,I15088,I15070,I15070,I15094,I15143,I15146,I15149,I15152,I15155,I15158,I15161,I15164,I15167,I2224,I2231);
PAT_14 I_183 (I15146,I15161,I15149,I15158,I15152,I15143,I15155,I15164,I15143,I15167,I15146,I15213,I15216,I15219,I15222,I15225,I15228,I15231,I15234,I15237,I2224,I2231);
PAT_5 I_184 (I15216,I15219,I15216,I15225,I15213,I15234,I15222,I15213,I15237,I15231,I15228,I15283,I15286,I15289,I15292,I15295,I15298,I15301,I15304,I15307,I15310,I2224,I2231);
PAT_13 I_185 (I15289,I15298,I15283,I15286,I15307,I15292,I15304,I15283,I15301,I15310,I15295,I15356,I15359,I15362,I15365,I15368,I15371,I15374,I15377,I15380,I2224,I2231);
PAT_14 I_186 (I15359,I15374,I15362,I15371,I15365,I15356,I15368,I15377,I15356,I15380,I15359,I15426,I15429,I15432,I15435,I15438,I15441,I15444,I15447,I15450,I2224,I2231);
PAT_17 I_187 (I15441,I15429,I15450,I15426,I15447,I15435,I15432,I15444,I15438,I15429,I15426,I15496,I15499,I15502,I15505,I15508,I15511,I15514,I15517,I15520,I15523,I2224,I2231);
PAT_7 I_188 (I15514,I15505,I15511,I15499,I15508,I15517,I15523,I15496,I15520,I15502,I15496,I15569,I15572,I15575,I15578,I15581,I15584,I15587,I15590,I15593,I2224,I2231);
PAT_17 I_189 (I15581,I15575,I15584,I15569,I15587,I15590,I15572,I15593,I15578,I15572,I15569,I15639,I15642,I15645,I15648,I15651,I15654,I15657,I15660,I15663,I15666,I2224,I2231);
PAT_1 I_190 (I15663,I15666,I15645,I15654,I15639,I15660,I15651,I15642,I15648,I15639,I15657,I15712,I15715,I15718,I15721,I15724,I15727,I15730,I15733,I15736,I2224,I2231);
PAT_10 I_191 (I15727,I15724,I15715,I15712,I15715,I15730,I15718,I15733,I15736,I15721,I15712,I15782,I15785,I15788,I15791,I15794,I15797,I15800,I15803,I2224,I2231);
PAT_5 I_192 (I15803,I15782,I15791,I15785,I15800,I15797,I15788,I15788,I15782,I15785,I15794,I15849,I15852,I15855,I15858,I15861,I15864,I15867,I15870,I15873,I15876,I2224,I2231);
PAT_6 I_193 (I15867,I15861,I15849,I15855,I15852,I15858,I15864,I15849,I15873,I15870,I15876,I15922,I15925,I15928,I15931,I15934,I15937,I15940,I15943,I15946,I15949,I2224,I2231);
PAT_8 I_194 (I15931,I15937,I15928,I15940,I15922,I15925,I15943,I15922,I15949,I15946,I15934,I15995,I15998,I16001,I16004,I16007,I16010,I16013,I16016,I16019,I2224,I2231);
PAT_7 I_195 (I15995,I16004,I16001,I16007,I16013,I15995,I15998,I16016,I16019,I16010,I15998,I16065,I16068,I16071,I16074,I16077,I16080,I16083,I16086,I16089,I2224,I2231);
PAT_0 I_196 (I16068,I16068,I16074,I16071,I16080,I16089,I16077,I16065,I16083,I16065,I16086,I16135,I16138,I16141,I16144,I16147,I16150,I16153,I16156,I2224,I2231);
PAT_5 I_197 (I16156,I16138,I16153,I16135,I16138,I16141,I16147,I16141,I16144,I16150,I16135,I16202,I16205,I16208,I16211,I16214,I16217,I16220,I16223,I16226,I16229,I2224,I2231);
PAT_2 I_198 (I16217,I16202,I16214,I16208,I16223,I16205,I16220,I16211,I16226,I16229,I16202,I16275,I16278,I16281,I16284,I16287,I16290,I16293,I16296,I16299,I2224,I2231);
PAT_5 I_199 (I16296,I16275,I16275,I16287,I16284,I16293,I16281,I16290,I16299,I16278,I16278,I16345,I16348,I16351,I16354,I16357,I16360,I16363,I16366,I16369,I16372,I2224,I2231);
PAT_10 I_200 (I16369,I16372,I16351,I16357,I16360,I16366,I16348,I16345,I16345,I16354,I16363,I16418,I16421,I16424,I16427,I16430,I16433,I16436,I16439,I2224,I2231);
PAT_6 I_201 (I16439,I16433,I16427,I16421,I16418,I16424,I16418,I16424,I16421,I16430,I16436,I16485,I16488,I16491,I16494,I16497,I16500,I16503,I16506,I16509,I16512,I2224,I2231);
PAT_4 I_202 (I16485,I16500,I16488,I16491,I16494,I16485,I16512,I16503,I16506,I16497,I16509,I16558,I16561,I16564,I16567,I16570,I16573,I16576,I16579,I16582,I2224,I2231);
PAT_11 I_203 (I16570,I16579,I16561,I16573,I16558,I16561,I16558,I16567,I16582,I16576,I16564,I16628,I16631,I16634,I16637,I16640,I16643,I16646,I16649,I16652,I16655,I2224,I2231);
PAT_5 I_204 (I16649,I16628,I16655,I16643,I16640,I16652,I16634,I16628,I16646,I16631,I16637,I16701,I16704,I16707,I16710,I16713,I16716,I16719,I16722,I16725,I16728,I2224,I2231);
PAT_9 I_205 (I16716,I16713,I16722,I16719,I16710,I16701,I16707,I16728,I16704,I16725,I16701,I16774,I16777,I16780,I16783,I16786,I16789,I16792,I16795,I16798,I2224,I2231);
PAT_4 I_206 (I16774,I16798,I16792,I16780,I16777,I16795,I16777,I16774,I16789,I16783,I16786,I16844,I16847,I16850,I16853,I16856,I16859,I16862,I16865,I16868,I2224,I2231);
PAT_12 I_207 (I16844,I16847,I16865,I16868,I16859,I16850,I16856,I16853,I16844,I16862,I16847,I16914,I16917,I16920,I16923,I16926,I16929,I16932,I16935,I2224,I2231);
PAT_5 I_208 (I16923,I16929,I16935,I16920,I16920,I16914,I16932,I16914,I16917,I16917,I16926,I16981,I16984,I16987,I16990,I16993,I16996,I16999,I17002,I17005,I17008,I2224,I2231);
PAT_8 I_209 (I16981,I17008,I16999,I16996,I16990,I16981,I16993,I17005,I16984,I17002,I16987,I17054,I17057,I17060,I17063,I17066,I17069,I17072,I17075,I17078,I2224,I2231);
PAT_4 I_210 (I17072,I17057,I17063,I17054,I17054,I17066,I17057,I17075,I17078,I17060,I17069,I17124,I17127,I17130,I17133,I17136,I17139,I17142,I17145,I17148,I2224,I2231);
PAT_7 I_211 (I17139,I17133,I17130,I17124,I17136,I17142,I17127,I17127,I17145,I17148,I17124,I17194,I17197,I17200,I17203,I17206,I17209,I17212,I17215,I17218,I2224,I2231);
PAT_11 I_212 (I17206,I17200,I17194,I17215,I17218,I17203,I17197,I17212,I17194,I17209,I17197,I17264,I17267,I17270,I17273,I17276,I17279,I17282,I17285,I17288,I17291,I2224,I2231);
PAT_9 I_213 (I17270,I17282,I17273,I17285,I17264,I17267,I17276,I17264,I17279,I17288,I17291,I17337,I17340,I17343,I17346,I17349,I17352,I17355,I17358,I17361,I2224,I2231);
PAT_6 I_214 (I17355,I17337,I17349,I17358,I17337,I17346,I17343,I17361,I17352,I17340,I17340,I17407,I17410,I17413,I17416,I17419,I17422,I17425,I17428,I17431,I17434,I2224,I2231);
PAT_4 I_215 (I17407,I17422,I17410,I17413,I17416,I17407,I17434,I17425,I17428,I17419,I17431,I17480,I17483,I17486,I17489,I17492,I17495,I17498,I17501,I17504,I2224,I2231);
PAT_1 I_216 (I17480,I17501,I17498,I17483,I17495,I17480,I17483,I17504,I17489,I17486,I17492,I17550,I17553,I17556,I17559,I17562,I17565,I17568,I17571,I17574,I2224,I2231);
PAT_4 I_217 (I17562,I17568,I17550,I17553,I17556,I17559,I17571,I17553,I17565,I17550,I17574,I17620,I17623,I17626,I17629,I17632,I17635,I17638,I17641,I17644,I2224,I2231);
PAT_11 I_218 (I17632,I17641,I17623,I17635,I17620,I17623,I17620,I17629,I17644,I17638,I17626,I17690,I17693,I17696,I17699,I17702,I17705,I17708,I17711,I17714,I17717,I2224,I2231);
PAT_15 I_219 (I17714,I17693,I17699,I17708,I17705,I17690,I17702,I17711,I17690,I17696,I17717,I17763,I17766,I17769,I17772,I17775,I17778,I17781,I17784,I17787,I2224,I2231);
PAT_13 I_220 (I17772,I17763,I17781,I17766,I17766,I17784,I17775,I17763,I17778,I17787,I17769,I17833,I17836,I17839,I17842,I17845,I17848,I17851,I17854,I17857,I2224,I2231);
PAT_17 I_221 (I17857,I17845,I17854,I17851,I17842,I17833,I17836,I17839,I17833,I17848,I17836,I17903,I17906,I17909,I17912,I17915,I17918,I17921,I17924,I17927,I17930,I2224,I2231);
PAT_9 I_222 (I17924,I17906,I17912,I17927,I17909,I17921,I17903,I17915,I17903,I17930,I17918,I17976,I17979,I17982,I17985,I17988,I17991,I17994,I17997,I18000,I2224,I2231);
PAT_2 I_223 (I17991,I17994,I17985,I18000,I17976,I17979,I17982,I17979,I17997,I17988,I17976,I18046,I18049,I18052,I18055,I18058,I18061,I18064,I18067,I18070,I2224,I2231);
PAT_9 I_224 (I18061,I18070,I18046,I18052,I18055,I18064,I18049,I18058,I18067,I18049,I18046,I18116,I18119,I18122,I18125,I18128,I18131,I18134,I18137,I18140,I2224,I2231);
PAT_6 I_225 (I18134,I18116,I18128,I18137,I18116,I18125,I18122,I18140,I18131,I18119,I18119,I18186,I18189,I18192,I18195,I18198,I18201,I18204,I18207,I18210,I18213,I2224,I2231);
PAT_3 I_226 (I18189,I18186,I18186,I18198,I18195,I18213,I18192,I18201,I18204,I18210,I18207,I18259,I18262,I18265,I18268,I18271,I18274,I18277,I18280,I18283,I18286,I2224,I2231);
PAT_1 I_227 (I18286,I18283,I18271,I18262,I18280,I18268,I18259,I18277,I18259,I18274,I18265,I18332,I18335,I18338,I18341,I18344,I18347,I18350,I18353,I18356,I2224,I2231);
PAT_17 I_228 (I18344,I18332,I18353,I18356,I18335,I18338,I18335,I18347,I18341,I18332,I18350,I18402,I18405,I18408,I18411,I18414,I18417,I18420,I18423,I18426,I18429,I2224,I2231);
PAT_2 I_229 (I18402,I18420,I18417,I18402,I18411,I18426,I18423,I18408,I18429,I18414,I18405,I18475,I18478,I18481,I18484,I18487,I18490,I18493,I18496,I18499,I2224,I2231);
PAT_14 I_230 (I18481,I18484,I18499,I18490,I18475,I18478,I18493,I18487,I18475,I18496,I18478,I18545,I18548,I18551,I18554,I18557,I18560,I18563,I18566,I18569,I2224,I2231);
PAT_1 I_231 (I18545,I18569,I18554,I18548,I18548,I18551,I18560,I18563,I18557,I18545,I18566,I18615,I18618,I18621,I18624,I18627,I18630,I18633,I18636,I18639,I2224,I2231);
PAT_11 I_232 (I18618,I18633,I18630,I18636,I18639,I18618,I18624,I18627,I18615,I18621,I18615,I18685,I18688,I18691,I18694,I18697,I18700,I18703,I18706,I18709,I18712,I2224,I2231);
PAT_7 I_233 (I18709,I18694,I18691,I18712,I18697,I18685,I18685,I18703,I18706,I18688,I18700,I18758,I18761,I18764,I18767,I18770,I18773,I18776,I18779,I18782,I2224,I2231);
PAT_14 I_234 (I18773,I18767,I18758,I18761,I18770,I18776,I18764,I18779,I18761,I18758,I18782,I18828,I18831,I18834,I18837,I18840,I18843,I18846,I18849,I18852,I2224,I2231);
PAT_17 I_235 (I18843,I18831,I18852,I18828,I18849,I18837,I18834,I18846,I18840,I18831,I18828,I18898,I18901,I18904,I18907,I18910,I18913,I18916,I18919,I18922,I18925,I2224,I2231);
PAT_1 I_236 (I18922,I18925,I18904,I18913,I18898,I18919,I18910,I18901,I18907,I18898,I18916,I18971,I18974,I18977,I18980,I18983,I18986,I18989,I18992,I18995,I2224,I2231);
PAT_9 I_237 (I18986,I18992,I18977,I18995,I18974,I18989,I18974,I18980,I18971,I18983,I18971,I19041,I19044,I19047,I19050,I19053,I19056,I19059,I19062,I19065,I2224,I2231);
PAT_1 I_238 (I19041,I19059,I19041,I19053,I19044,I19050,I19056,I19062,I19065,I19047,I19044,I19111,I19114,I19117,I19120,I19123,I19126,I19129,I19132,I19135,I2224,I2231);
PAT_13 I_239 (I19120,I19129,I19135,I19111,I19126,I19123,I19132,I19117,I19114,I19111,I19114,I19181,I19184,I19187,I19190,I19193,I19196,I19199,I19202,I19205,I2224,I2231);
PAT_2 I_240 (I19199,I19193,I19190,I19196,I19181,I19205,I19184,I19202,I19181,I19187,I19184,I19251,I19254,I19257,I19260,I19263,I19266,I19269,I19272,I19275,I2224,I2231);
PAT_5 I_241 (I19272,I19251,I19251,I19263,I19260,I19269,I19257,I19266,I19275,I19254,I19254,I19321,I19324,I19327,I19330,I19333,I19336,I19339,I19342,I19345,I19348,I2224,I2231);
PAT_6 I_242 (I19339,I19333,I19321,I19327,I19324,I19330,I19336,I19321,I19345,I19342,I19348,I19394,I19397,I19400,I19403,I19406,I19409,I19412,I19415,I19418,I19421,I2224,I2231);
PAT_17 I_243 (I19406,I19409,I19415,I19403,I19397,I19418,I19412,I19394,I19421,I19400,I19394,I19467,I19470,I19473,I19476,I19479,I19482,I19485,I19488,I19491,I19494,I2224,I2231);
PAT_10 I_244 (I19467,I19473,I19494,I19476,I19491,I19470,I19485,I19479,I19488,I19482,I19467,I19540,I19543,I19546,I19549,I19552,I19555,I19558,I19561,I2224,I2231);
PAT_8 I_245 (I19561,I19552,I19543,I19540,I19549,I19540,I19555,I19543,I19558,I19546,I19546,I19607,I19610,I19613,I19616,I19619,I19622,I19625,I19628,I19631,I2224,I2231);
PAT_17 I_246 (I19631,I19619,I19616,I19610,I19613,I19625,I19607,I19610,I19607,I19622,I19628,I19677,I19680,I19683,I19686,I19689,I19692,I19695,I19698,I19701,I19704,I2224,I2231);
PAT_4 I_247 (I19686,I19677,I19695,I19692,I19704,I19701,I19680,I19677,I19683,I19689,I19698,I19750,I19753,I19756,I19759,I19762,I19765,I19768,I19771,I19774,I2224,I2231);
PAT_15 I_248 (I19750,I19753,I19774,I19759,I19768,I19771,I19756,I19765,I19762,I19750,I19753,I19820,I19823,I19826,I19829,I19832,I19835,I19838,I19841,I19844,I2224,I2231);
PAT_13 I_249 (I19829,I19820,I19838,I19823,I19823,I19841,I19832,I19820,I19835,I19844,I19826,I19890,I19893,I19896,I19899,I19902,I19905,I19908,I19911,I19914,I2224,I2231);
PAT_12 I_250 (I19899,I19890,I19890,I19914,I19911,I19893,I19908,I19902,I19893,I19896,I19905,I19960,I19963,I19966,I19969,I19972,I19975,I19978,I19981,I2224,I2231);
PAT_13 I_251 (I19972,I19975,I19966,I19981,I19978,I19960,I19963,I19969,I19966,I19963,I19960,I20027,I20030,I20033,I20036,I20039,I20042,I20045,I20048,I20051,I2224,I2231);
PAT_11 I_252 (I20027,I20039,I20042,I20033,I20030,I20051,I20030,I20048,I20036,I20027,I20045,I20097,I20100,I20103,I20106,I20109,I20112,I20115,I20118,I20121,I20124,I2224,I2231);
PAT_4 I_253 (I20103,I20124,I20097,I20115,I20106,I20097,I20118,I20100,I20109,I20121,I20112,I20170,I20173,I20176,I20179,I20182,I20185,I20188,I20191,I20194,I2224,I2231);
PAT_2 I_254 (I20179,I20173,I20173,I20194,I20170,I20188,I20185,I20176,I20170,I20182,I20191,I20240,I20243,I20246,I20249,I20252,I20255,I20258,I20261,I20264,I2224,I2231);
PAT_4 I_255 (I20240,I20246,I20264,I20258,I20255,I20252,I20243,I20261,I20240,I20243,I20249,I20310,I20313,I20316,I20319,I20322,I20325,I20328,I20331,I20334,I2224,I2231);
PAT_9 I_256 (I20331,I20313,I20316,I20325,I20328,I20310,I20319,I20313,I20334,I20310,I20322,I20380,I20383,I20386,I20389,I20392,I20395,I20398,I20401,I20404,I2224,I2231);
PAT_17 I_257 (I20383,I20389,I20404,I20395,I20398,I20386,I20380,I20392,I20380,I20383,I20401,I20450,I20453,I20456,I20459,I20462,I20465,I20468,I20471,I20474,I20477,I2224,I2231);
PAT_8 I_258 (I20459,I20471,I20477,I20468,I20453,I20462,I20465,I20474,I20456,I20450,I20450,I20523,I20526,I20529,I20532,I20535,I20538,I20541,I20544,I20547,I2224,I2231);
PAT_4 I_259 (I20541,I20526,I20532,I20523,I20523,I20535,I20526,I20544,I20547,I20529,I20538,I20593,I20596,I20599,I20602,I20605,I20608,I20611,I20614,I20617,I2224,I2231);
PAT_1 I_260 (I20593,I20614,I20611,I20596,I20608,I20593,I20596,I20617,I20602,I20599,I20605,I20663,I20666,I20669,I20672,I20675,I20678,I20681,I20684,I20687,I2224,I2231);
PAT_6 I_261 (I20672,I20663,I20666,I20669,I20684,I20687,I20681,I20663,I20678,I20675,I20666,I20733,I20736,I20739,I20742,I20745,I20748,I20751,I20754,I20757,I20760,I2224,I2231);
PAT_11 I_262 (I20733,I20748,I20733,I20745,I20742,I20760,I20757,I20754,I20751,I20736,I20739,I20806,I20809,I20812,I20815,I20818,I20821,I20824,I20827,I20830,I20833,I2224,I2231);
PAT_1 I_263 (I20821,I20812,I20815,I20806,I20827,I20824,I20809,I20806,I20833,I20830,I20818,I20879,I20882,I20885,I20888,I20891,I20894,I20897,I20900,I20903,I2224,I2231);
PAT_4 I_264 (I20891,I20897,I20879,I20882,I20885,I20888,I20900,I20882,I20894,I20879,I20903,I20949,I20952,I20955,I20958,I20961,I20964,I20967,I20970,I20973,I2224,I2231);
PAT_10 I_265 (I20949,I20949,I20973,I20952,I20958,I20967,I20964,I20952,I20970,I20955,I20961,I21019,I21022,I21025,I21028,I21031,I21034,I21037,I21040,I2224,I2231);
PAT_15 I_266 (I21034,I21037,I21025,I21031,I21019,I21019,I21025,I21040,I21028,I21022,I21022,I21086,I21089,I21092,I21095,I21098,I21101,I21104,I21107,I21110,I2224,I2231);
PAT_13 I_267 (I21095,I21086,I21104,I21089,I21089,I21107,I21098,I21086,I21101,I21110,I21092,I21156,I21159,I21162,I21165,I21168,I21171,I21174,I21177,I21180,I2224,I2231);
PAT_17 I_268 (I21180,I21168,I21177,I21174,I21165,I21156,I21159,I21162,I21156,I21171,I21159,I21226,I21229,I21232,I21235,I21238,I21241,I21244,I21247,I21250,I21253,I2224,I2231);
PAT_4 I_269 (I21235,I21226,I21244,I21241,I21253,I21250,I21229,I21226,I21232,I21238,I21247,I21299,I21302,I21305,I21308,I21311,I21314,I21317,I21320,I21323,I2224,I2231);
PAT_8 I_270 (I21311,I21299,I21320,I21305,I21302,I21323,I21308,I21317,I21302,I21299,I21314,I21369,I21372,I21375,I21378,I21381,I21384,I21387,I21390,I21393,I2224,I2231);
PAT_4 I_271 (I21387,I21372,I21378,I21369,I21369,I21381,I21372,I21390,I21393,I21375,I21384,I21439,I21442,I21445,I21448,I21451,I21454,I21457,I21460,I21463,I2224,I2231);
PAT_8 I_272 (I21451,I21439,I21460,I21445,I21442,I21463,I21448,I21457,I21442,I21439,I21454,I21509,I21512,I21515,I21518,I21521,I21524,I21527,I21530,I21533,I2224,I2231);
PAT_2 I_273 (I21512,I21527,I21533,I21509,I21521,I21524,I21512,I21530,I21515,I21518,I21509,I21579,I21582,I21585,I21588,I21591,I21594,I21597,I21600,I21603,I2224,I2231);
PAT_9 I_274 (I21594,I21603,I21579,I21585,I21588,I21597,I21582,I21591,I21600,I21582,I21579,I21649,I21652,I21655,I21658,I21661,I21664,I21667,I21670,I21673,I2224,I2231);
PAT_16 I_275 (I21655,I21658,I21673,I21649,I21661,I21652,I21649,I21664,I21670,I21667,I21652,I21719,I21722,I21725,I21728,I21731,I21734,I21737,I21740,I21743,I21746,I2224,I2231);
PAT_10 I_276 (I21719,I21731,I21746,I21734,I21740,I21743,I21728,I21719,I21737,I21725,I21722,I21792,I21795,I21798,I21801,I21804,I21807,I21810,I21813,I2224,I2231);
PAT_9 I_277 (I21804,I21792,I21795,I21798,I21792,I21798,I21801,I21795,I21813,I21807,I21810,I21859,I21862,I21865,I21868,I21871,I21874,I21877,I21880,I21883,I2224,I2231);
PAT_10 I_278 (I21880,I21877,I21865,I21862,I21883,I21868,I21874,I21862,I21859,I21859,I21871,I21929,I21932,I21935,I21938,I21941,I21944,I21947,I21950,I2224,I2231);
PAT_7 I_279 (I1577,I1889,I1409,I1833,I2081,I2001,I1353,I1345,I1561,I2049,I1609,I21996,I21999,I22002,I22005,I22008,I22011,I22014,I22017,I22020,I2224,I2231);
PAT_5 I_280 (I22002,I21996,I22005,I22014,I22008,I22020,I22017,I21999,I22011,I21999,I21996,I22066,I22069,I22072,I22075,I22078,I22081,I22084,I22087,I22090,I22093,I2224,I2231);
PAT_14 I_281 (I22087,I22072,I22066,I22090,I22093,I22066,I22084,I22069,I22075,I22078,I22081,I22139,I22142,I22145,I22148,I22151,I22154,I22157,I22160,I22163,I2224,I2231);
PAT_9 I_282 (I22148,I22160,I22139,I22157,I22142,I22145,I22163,I22142,I22151,I22139,I22154,I22209,I22212,I22215,I22218,I22221,I22224,I22227,I22230,I22233,I2224,I2231);
PAT_17 I_283 (I22212,I22218,I22233,I22224,I22227,I22215,I22209,I22221,I22209,I22212,I22230,I22279,I22282,I22285,I22288,I22291,I22294,I22297,I22300,I22303,I22306,I2224,I2231);
PAT_3 I_284 (I22291,I22294,I22297,I22300,I22279,I22279,I22285,I22303,I22306,I22288,I22282,I22352,I22355,I22358,I22361,I22364,I22367,I22370,I22373,I22376,I22379,I2224,I2231);
PAT_15 I_285 (I22370,I22379,I22352,I22352,I22361,I22355,I22373,I22364,I22358,I22367,I22376,I22425,I22428,I22431,I22434,I22437,I22440,I22443,I22446,I22449,I2224,I2231);
PAT_12 I_286 (I22443,I22446,I22449,I22437,I22434,I22428,I22425,I22440,I22431,I22425,I22428,I22495,I22498,I22501,I22504,I22507,I22510,I22513,I22516,I2224,I2231);
PAT_11 I_287 (I22501,I22504,I22501,I22513,I22516,I22510,I22498,I22507,I22495,I22498,I22495,I22562,I22565,I22568,I22571,I22574,I22577,I22580,I22583,I22586,I22589,I2224,I2231);
PAT_17 I_288 (I22574,I22565,I22589,I22562,I22571,I22583,I22580,I22577,I22562,I22586,I22568,I22635,I22638,I22641,I22644,I22647,I22650,I22653,I22656,I22659,I22662,I2224,I2231);
PAT_5 I_289 (I22647,I22641,I22638,I22659,I22644,I22650,I22653,I22635,I22635,I22656,I22662,I22708,I22711,I22714,I22717,I22720,I22723,I22726,I22729,I22732,I22735,I2224,I2231);
PAT_1 I_290 (I22723,I22711,I22729,I22708,I22714,I22708,I22717,I22732,I22726,I22735,I22720,I22781,I22784,I22787,I22790,I22793,I22796,I22799,I22802,I22805,I2224,I2231);
PAT_13 I_291 (I22790,I22799,I22805,I22781,I22796,I22793,I22802,I22787,I22784,I22781,I22784,I22851,I22854,I22857,I22860,I22863,I22866,I22869,I22872,I22875,I2224,I2231);
PAT_14 I_292 (I22854,I22869,I22857,I22866,I22860,I22851,I22863,I22872,I22851,I22875,I22854,I22921,I22924,I22927,I22930,I22933,I22936,I22939,I22942,I22945,I2224,I2231);
PAT_16 I_293 (I22936,I22942,I22939,I22945,I22927,I22921,I22930,I22924,I22924,I22933,I22921,I22991,I22994,I22997,I23000,I23003,I23006,I23009,I23012,I23015,I23018,I2224,I2231);
PAT_10 I_294 (I22991,I23003,I23018,I23006,I23012,I23015,I23000,I22991,I23009,I22997,I22994,I23064,I23067,I23070,I23073,I23076,I23079,I23082,I23085,I2224,I2231);
PAT_17 I_295 (I23076,I23085,I23079,I23064,I23070,I23082,I23067,I23067,I23064,I23070,I23073,I23131,I23134,I23137,I23140,I23143,I23146,I23149,I23152,I23155,I23158,I2224,I2231);
PAT_5 I_296 (I23143,I23137,I23134,I23155,I23140,I23146,I23149,I23131,I23131,I23152,I23158,I23204,I23207,I23210,I23213,I23216,I23219,I23222,I23225,I23228,I23231,I2224,I2231);
PAT_9 I_297 (I23219,I23216,I23225,I23222,I23213,I23204,I23210,I23231,I23207,I23228,I23204,I23277,I23280,I23283,I23286,I23289,I23292,I23295,I23298,I23301,I2224,I2231);
PAT_8 I_298 (I23298,I23286,I23295,I23277,I23280,I23292,I23301,I23280,I23283,I23289,I23277,I23347,I23350,I23353,I23356,I23359,I23362,I23365,I23368,I23371,I2224,I2231);
PAT_9 I_299 (I23350,I23359,I23350,I23347,I23362,I23353,I23368,I23356,I23365,I23347,I23371,I23417,I23420,I23423,I23426,I23429,I23432,I23435,I23438,I23441,I2224,I2231);
PAT_13 I_300 (I23417,I23438,I23420,I23435,I23429,I23426,I23441,I23417,I23423,I23432,I23420,I23487,I23490,I23493,I23496,I23499,I23502,I23505,I23508,I23511,I2224,I2231);
PAT_5 I_301 (I23499,I23490,I23496,I23508,I23490,I23511,I23493,I23502,I23487,I23487,I23505,I23557,I23560,I23563,I23566,I23569,I23572,I23575,I23578,I23581,I23584,I2224,I2231);
PAT_2 I_302 (I23572,I23557,I23569,I23563,I23578,I23560,I23575,I23566,I23581,I23584,I23557,I23630,I23633,I23636,I23639,I23642,I23645,I23648,I23651,I23654,I2224,I2231);
PAT_13 I_303 (I23639,I23633,I23630,I23651,I23642,I23645,I23633,I23636,I23648,I23654,I23630,I23700,I23703,I23706,I23709,I23712,I23715,I23718,I23721,I23724,I2224,I2231);
PAT_15 I_304 (I23700,I23712,I23703,I23715,I23700,I23709,I23724,I23721,I23706,I23718,I23703,I23770,I23773,I23776,I23779,I23782,I23785,I23788,I23791,I23794,I2224,I2231);
PAT_17 I_305 (I23770,I23770,I23782,I23773,I23776,I23794,I23791,I23785,I23773,I23779,I23788,I23840,I23843,I23846,I23849,I23852,I23855,I23858,I23861,I23864,I23867,I2224,I2231);
PAT_2 I_306 (I23840,I23858,I23855,I23840,I23849,I23864,I23861,I23846,I23867,I23852,I23843,I23913,I23916,I23919,I23922,I23925,I23928,I23931,I23934,I23937,I2224,I2231);
PAT_14 I_307 (I23919,I23922,I23937,I23928,I23913,I23916,I23931,I23925,I23913,I23934,I23916,I23983,I23986,I23989,I23992,I23995,I23998,I24001,I24004,I24007,I2224,I2231);
PAT_6 I_308 (I23983,I23986,I24007,I23992,I23983,I23989,I23995,I23998,I24001,I23986,I24004,I24053,I24056,I24059,I24062,I24065,I24068,I24071,I24074,I24077,I24080,I2224,I2231);
PAT_12 I_309 (I24053,I24080,I24059,I24062,I24056,I24053,I24074,I24068,I24071,I24065,I24077,I24126,I24129,I24132,I24135,I24138,I24141,I24144,I24147,I2224,I2231);
PAT_9 I_310 (I24135,I24141,I24126,I24132,I24138,I24129,I24126,I24129,I24147,I24132,I24144,I24193,I24196,I24199,I24202,I24205,I24208,I24211,I24214,I24217,I2224,I2231);
PAT_6 I_311 (I24211,I24193,I24205,I24214,I24193,I24202,I24199,I24217,I24208,I24196,I24196,I24263,I24266,I24269,I24272,I24275,I24278,I24281,I24284,I24287,I24290,I2224,I2231);
PAT_4 I_312 (I24263,I24278,I24266,I24269,I24272,I24263,I24290,I24281,I24284,I24275,I24287,I24336,I24339,I24342,I24345,I24348,I24351,I24354,I24357,I24360,I2224,I2231);
PAT_3 I_313 (I24351,I24345,I24339,I24342,I24336,I24357,I24348,I24339,I24354,I24360,I24336,I24406,I24409,I24412,I24415,I24418,I24421,I24424,I24427,I24430,I24433,I2224,I2231);
PAT_14 I_314 (I24412,I24409,I24415,I24427,I24421,I24430,I24418,I24406,I24424,I24433,I24406,I24479,I24482,I24485,I24488,I24491,I24494,I24497,I24500,I24503,I2224,I2231);
PAT_7 I_315 (I24479,I24488,I24485,I24491,I24482,I24503,I24482,I24500,I24497,I24494,I24479,I24549,I24552,I24555,I24558,I24561,I24564,I24567,I24570,I24573,I2224,I2231);
PAT_2 I_316 (I24570,I24564,I24555,I24549,I24558,I24552,I24561,I24573,I24567,I24552,I24549,I24619,I24622,I24625,I24628,I24631,I24634,I24637,I24640,I24643,I2224,I2231);
PAT_13 I_317 (I24628,I24622,I24619,I24640,I24631,I24634,I24622,I24625,I24637,I24643,I24619,I24689,I24692,I24695,I24698,I24701,I24704,I24707,I24710,I24713,I2224,I2231);
PAT_15 I_318 (I24689,I24701,I24692,I24704,I24689,I24698,I24713,I24710,I24695,I24707,I24692,I24759,I24762,I24765,I24768,I24771,I24774,I24777,I24780,I24783,I2224,I2231);
PAT_14 I_319 (I24762,I24762,I24783,I24759,I24765,I24759,I24774,I24771,I24780,I24768,I24777,I24829,I24832,I24835,I24838,I24841,I24844,I24847,I24850,I24853,I2224,I2231);
PAT_5 I_320 (I24832,I24835,I24832,I24841,I24829,I24850,I24838,I24829,I24853,I24847,I24844,I24899,I24902,I24905,I24908,I24911,I24914,I24917,I24920,I24923,I24926,I2224,I2231);
PAT_12 I_321 (I24926,I24914,I24899,I24923,I24902,I24899,I24905,I24908,I24911,I24917,I24920,I24972,I24975,I24978,I24981,I24984,I24987,I24990,I24993,I2224,I2231);
PAT_17 I_322 (I24987,I24981,I24975,I24972,I24972,I24978,I24978,I24990,I24993,I24975,I24984,I25039,I25042,I25045,I25048,I25051,I25054,I25057,I25060,I25063,I25066,I2224,I2231);
PAT_1 I_323 (I25063,I25066,I25045,I25054,I25039,I25060,I25051,I25042,I25048,I25039,I25057,I25112,I25115,I25118,I25121,I25124,I25127,I25130,I25133,I25136,I2224,I2231);
PAT_10 I_324 (I25127,I25124,I25115,I25112,I25115,I25130,I25118,I25133,I25136,I25121,I25112,I25182,I25185,I25188,I25191,I25194,I25197,I25200,I25203,I2224,I2231);
PAT_5 I_325 (I25203,I25182,I25191,I25185,I25200,I25197,I25188,I25188,I25182,I25185,I25194,I25249,I25252,I25255,I25258,I25261,I25264,I25267,I25270,I25273,I25276,I2224,I2231);
PAT_9 I_326 (I25264,I25261,I25270,I25267,I25258,I25249,I25255,I25276,I25252,I25273,I25249,I25322,I25325,I25328,I25331,I25334,I25337,I25340,I25343,I25346,I2224,I2231);
PAT_4 I_327 (I25322,I25346,I25340,I25328,I25325,I25343,I25325,I25322,I25337,I25331,I25334,I25392,I25395,I25398,I25401,I25404,I25407,I25410,I25413,I25416,I2224,I2231);
PAT_10 I_328 (I25392,I25392,I25416,I25395,I25401,I25410,I25407,I25395,I25413,I25398,I25404,I25462,I25465,I25468,I25471,I25474,I25477,I25480,I25483,I2224,I2231);
PAT_6 I_329 (I25483,I25477,I25471,I25465,I25462,I25468,I25462,I25468,I25465,I25474,I25480,I25529,I25532,I25535,I25538,I25541,I25544,I25547,I25550,I25553,I25556,I2224,I2231);
PAT_13 I_330 (I25553,I25535,I25550,I25529,I25532,I25538,I25556,I25541,I25547,I25529,I25544,I25602,I25605,I25608,I25611,I25614,I25617,I25620,I25623,I25626,I2224,I2231);
PAT_5 I_331 (I25614,I25605,I25611,I25623,I25605,I25626,I25608,I25617,I25602,I25602,I25620,I25672,I25675,I25678,I25681,I25684,I25687,I25690,I25693,I25696,I25699,I2224,I2231);
PAT_9 I_332 (I25687,I25684,I25693,I25690,I25681,I25672,I25678,I25699,I25675,I25696,I25672,I25745,I25748,I25751,I25754,I25757,I25760,I25763,I25766,I25769,I2224,I2231);
PAT_13 I_333 (I25745,I25766,I25748,I25763,I25757,I25754,I25769,I25745,I25751,I25760,I25748,I25815,I25818,I25821,I25824,I25827,I25830,I25833,I25836,I25839,I2224,I2231);
PAT_5 I_334 (I25827,I25818,I25824,I25836,I25818,I25839,I25821,I25830,I25815,I25815,I25833,I25885,I25888,I25891,I25894,I25897,I25900,I25903,I25906,I25909,I25912,I2224,I2231);
PAT_12 I_335 (I25912,I25900,I25885,I25909,I25888,I25885,I25891,I25894,I25897,I25903,I25906,I25958,I25961,I25964,I25967,I25970,I25973,I25976,I25979,I2224,I2231);
PAT_4 I_336 (I25964,I25961,I25976,I25979,I25973,I25967,I25958,I25958,I25964,I25970,I25961,I26025,I26028,I26031,I26034,I26037,I26040,I26043,I26046,I26049,I2224,I2231);
PAT_7 I_337 (I26040,I26034,I26031,I26025,I26037,I26043,I26028,I26028,I26046,I26049,I26025,I26095,I26098,I26101,I26104,I26107,I26110,I26113,I26116,I26119,I2224,I2231);
PAT_17 I_338 (I26107,I26101,I26110,I26095,I26113,I26116,I26098,I26119,I26104,I26098,I26095,I26165,I26168,I26171,I26174,I26177,I26180,I26183,I26186,I26189,I26192,I2224,I2231);
PAT_7 I_339 (I26183,I26174,I26180,I26168,I26177,I26186,I26192,I26165,I26189,I26171,I26165,I26238,I26241,I26244,I26247,I26250,I26253,I26256,I26259,I26262,I2224,I2231);
PAT_2 I_340 (I26259,I26253,I26244,I26238,I26247,I26241,I26250,I26262,I26256,I26241,I26238,I26308,I26311,I26314,I26317,I26320,I26323,I26326,I26329,I26332,I2224,I2231);
PAT_14 I_341 (I26314,I26317,I26332,I26323,I26308,I26311,I26326,I26320,I26308,I26329,I26311,I26378,I26381,I26384,I26387,I26390,I26393,I26396,I26399,I26402,I2224,I2231);
PAT_9 I_342 (I26387,I26399,I26378,I26396,I26381,I26384,I26402,I26381,I26390,I26378,I26393,I26448,I26451,I26454,I26457,I26460,I26463,I26466,I26469,I26472,I2224,I2231);
PAT_4 I_343 (I26448,I26472,I26466,I26454,I26451,I26469,I26451,I26448,I26463,I26457,I26460,I26518,I26521,I26524,I26527,I26530,I26533,I26536,I26539,I26542,I2224,I2231);
PAT_2 I_344 (I26527,I26521,I26521,I26542,I26518,I26536,I26533,I26524,I26518,I26530,I26539,I26588,I26591,I26594,I26597,I26600,I26603,I26606,I26609,I26612,I2224,I2231);
PAT_11 I_345 (I26591,I26603,I26588,I26600,I26597,I26609,I26606,I26591,I26612,I26594,I26588,I26658,I26661,I26664,I26667,I26670,I26673,I26676,I26679,I26682,I26685,I2224,I2231);
PAT_15 I_346 (I26682,I26661,I26667,I26676,I26673,I26658,I26670,I26679,I26658,I26664,I26685,I26731,I26734,I26737,I26740,I26743,I26746,I26749,I26752,I26755,I2224,I2231);
PAT_13 I_347 (I26740,I26731,I26749,I26734,I26734,I26752,I26743,I26731,I26746,I26755,I26737,I26801,I26804,I26807,I26810,I26813,I26816,I26819,I26822,I26825,I2224,I2231);
PAT_8 I_348 (I26810,I26822,I26813,I26816,I26825,I26804,I26819,I26801,I26804,I26807,I26801,I26871,I26874,I26877,I26880,I26883,I26886,I26889,I26892,I26895,I2224,I2231);
PAT_13 I_349 (I26883,I26892,I26874,I26895,I26877,I26871,I26871,I26880,I26889,I26886,I26874,I26941,I26944,I26947,I26950,I26953,I26956,I26959,I26962,I26965,I2224,I2231);
PAT_12 I_350 (I26950,I26941,I26941,I26965,I26962,I26944,I26959,I26953,I26944,I26947,I26956,I27011,I27014,I27017,I27020,I27023,I27026,I27029,I27032,I2224,I2231);
PAT_4 I_351 (I27017,I27014,I27029,I27032,I27026,I27020,I27011,I27011,I27017,I27023,I27014,I27078,I27081,I27084,I27087,I27090,I27093,I27096,I27099,I27102,I2224,I2231);
PAT_5 I_352 (I27099,I27081,I27081,I27093,I27096,I27090,I27087,I27078,I27084,I27078,I27102,I27148,I27151,I27154,I27157,I27160,I27163,I27166,I27169,I27172,I27175,I2224,I2231);
PAT_3 I_353 (I27160,I27148,I27175,I27169,I27172,I27148,I27163,I27151,I27154,I27157,I27166,I27221,I27224,I27227,I27230,I27233,I27236,I27239,I27242,I27245,I27248,I2224,I2231);
PAT_13 I_354 (I27242,I27230,I27248,I27227,I27233,I27236,I27224,I27239,I27221,I27221,I27245,I27294,I27297,I27300,I27303,I27306,I27309,I27312,I27315,I27318,I2224,I2231);
PAT_15 I_355 (I27294,I27306,I27297,I27309,I27294,I27303,I27318,I27315,I27300,I27312,I27297,I27364,I27367,I27370,I27373,I27376,I27379,I27382,I27385,I27388,I2224,I2231);
PAT_4 I_356 (I27376,I27382,I27364,I27367,I27370,I27364,I27388,I27385,I27373,I27379,I27367,I27434,I27437,I27440,I27443,I27446,I27449,I27452,I27455,I27458,I2224,I2231);
PAT_7 I_357 (I27449,I27443,I27440,I27434,I27446,I27452,I27437,I27437,I27455,I27458,I27434,I27504,I27507,I27510,I27513,I27516,I27519,I27522,I27525,I27528,I2224,I2231);
PAT_1 I_358 (I27504,I27522,I27525,I27507,I27528,I27516,I27510,I27519,I27507,I27513,I27504,I27574,I27577,I27580,I27583,I27586,I27589,I27592,I27595,I27598,I2224,I2231);
PAT_2 I_359 (I27574,I27580,I27574,I27589,I27577,I27577,I27583,I27586,I27592,I27598,I27595,I27644,I27647,I27650,I27653,I27656,I27659,I27662,I27665,I27668,I2224,I2231);
PAT_4 I_360 (I27644,I27650,I27668,I27662,I27659,I27656,I27647,I27665,I27644,I27647,I27653,I27714,I27717,I27720,I27723,I27726,I27729,I27732,I27735,I27738,I2224,I2231);
PAT_13 I_361 (I27729,I27723,I27735,I27720,I27726,I27714,I27738,I27732,I27717,I27714,I27717,I27784,I27787,I27790,I27793,I27796,I27799,I27802,I27805,I27808,I2224,I2231);
PAT_7 I_362 (I27793,I27796,I27784,I27799,I27805,I27790,I27787,I27808,I27787,I27784,I27802,I27854,I27857,I27860,I27863,I27866,I27869,I27872,I27875,I27878,I2224,I2231);
PAT_5 I_363 (I27860,I27854,I27863,I27872,I27866,I27878,I27875,I27857,I27869,I27857,I27854,I27924,I27927,I27930,I27933,I27936,I27939,I27942,I27945,I27948,I27951,I2224,I2231);
PAT_2 I_364 (I27939,I27924,I27936,I27930,I27945,I27927,I27942,I27933,I27948,I27951,I27924,I27997,I28000,I28003,I28006,I28009,I28012,I28015,I28018,I28021,I2224,I2231);
PAT_13 I_365 (I28006,I28000,I27997,I28018,I28009,I28012,I28000,I28003,I28015,I28021,I27997,I28067,I28070,I28073,I28076,I28079,I28082,I28085,I28088,I28091,I2224,I2231);
PAT_14 I_366 (I28070,I28085,I28073,I28082,I28076,I28067,I28079,I28088,I28067,I28091,I28070,I28137,I28140,I28143,I28146,I28149,I28152,I28155,I28158,I28161,I2224,I2231);
PAT_13 I_367 (I28146,I28161,I28140,I28149,I28137,I28140,I28155,I28143,I28137,I28158,I28152,I28207,I28210,I28213,I28216,I28219,I28222,I28225,I28228,I28231,I2224,I2231);
PAT_14 I_368 (I28210,I28225,I28213,I28222,I28216,I28207,I28219,I28228,I28207,I28231,I28210,I28277,I28280,I28283,I28286,I28289,I28292,I28295,I28298,I28301,I2224,I2231);
PAT_4 I_369 (I28286,I28292,I28283,I28277,I28301,I28289,I28277,I28280,I28298,I28280,I28295,I28347,I28350,I28353,I28356,I28359,I28362,I28365,I28368,I28371,I2224,I2231);
PAT_13 I_370 (I28362,I28356,I28368,I28353,I28359,I28347,I28371,I28365,I28350,I28347,I28350,I28417,I28420,I28423,I28426,I28429,I28432,I28435,I28438,I28441,I2224,I2231);
PAT_7 I_371 (I28426,I28429,I28417,I28432,I28438,I28423,I28420,I28441,I28420,I28417,I28435,I28487,I28490,I28493,I28496,I28499,I28502,I28505,I28508,I28511,I2224,I2231);
PAT_1 I_372 (I28487,I28505,I28508,I28490,I28511,I28499,I28493,I28502,I28490,I28496,I28487,I28557,I28560,I28563,I28566,I28569,I28572,I28575,I28578,I28581,I2224,I2231);
PAT_11 I_373 (I28560,I28575,I28572,I28578,I28581,I28560,I28566,I28569,I28557,I28563,I28557,I28627,I28630,I28633,I28636,I28639,I28642,I28645,I28648,I28651,I28654,I2224,I2231);
PAT_10 I_374 (I28642,I28648,I28639,I28633,I28651,I28636,I28654,I28645,I28627,I28630,I28627,I28700,I28703,I28706,I28709,I28712,I28715,I28718,I28721,I2224,I2231);
PAT_15 I_375 (I28715,I28718,I28706,I28712,I28700,I28700,I28706,I28721,I28709,I28703,I28703,I28767,I28770,I28773,I28776,I28779,I28782,I28785,I28788,I28791,I2224,I2231);
PAT_10 I_376 (I28770,I28779,I28773,I28767,I28788,I28791,I28776,I28767,I28770,I28785,I28782,I28837,I28840,I28843,I28846,I28849,I28852,I28855,I28858,I2224,I2231);
PAT_2 I_377 (I28849,I28852,I28843,I28855,I28840,I28837,I28837,I28843,I28858,I28846,I28840,I28904,I28907,I28910,I28913,I28916,I28919,I28922,I28925,I28928,I2224,I2231);
PAT_4 I_378 (I28904,I28910,I28928,I28922,I28919,I28916,I28907,I28925,I28904,I28907,I28913,I28974,I28977,I28980,I28983,I28986,I28989,I28992,I28995,I28998,I2224,I2231);
PAT_8 I_379 (I28986,I28974,I28995,I28980,I28977,I28998,I28983,I28992,I28977,I28974,I28989,I29044,I29047,I29050,I29053,I29056,I29059,I29062,I29065,I29068,I2224,I2231);
PAT_10 I_380 (I29050,I29044,I29047,I29068,I29062,I29047,I29056,I29044,I29065,I29059,I29053,I29114,I29117,I29120,I29123,I29126,I29129,I29132,I29135,I2224,I2231);
PAT_14 I_381 (I29114,I29135,I29120,I29129,I29126,I29132,I29123,I29117,I29117,I29120,I29114,I29181,I29184,I29187,I29190,I29193,I29196,I29199,I29202,I29205,I2224,I2231);
PAT_9 I_382 (I29190,I29202,I29181,I29199,I29184,I29187,I29205,I29184,I29193,I29181,I29196,I29251,I29254,I29257,I29260,I29263,I29266,I29269,I29272,I29275,I2224,I2231);
PAT_7 I_383 (I29257,I29266,I29251,I29272,I29263,I29251,I29254,I29275,I29269,I29254,I29260,I29321,I29324,I29327,I29330,I29333,I29336,I29339,I29342,I29345,I2224,I2231);
PAT_5 I_384 (I29327,I29321,I29330,I29339,I29333,I29345,I29342,I29324,I29336,I29324,I29321,I29391,I29394,I29397,I29400,I29403,I29406,I29409,I29412,I29415,I29418,I2224,I2231);
PAT_7 I_385 (I29409,I29412,I29418,I29415,I29400,I29397,I29391,I29403,I29391,I29394,I29406,I29464,I29467,I29470,I29473,I29476,I29479,I29482,I29485,I29488,I2224,I2231);
PAT_17 I_386 (I29476,I29470,I29479,I29464,I29482,I29485,I29467,I29488,I29473,I29467,I29464,I29534,I29537,I29540,I29543,I29546,I29549,I29552,I29555,I29558,I29561,I2224,I2231);
PAT_3 I_387 (I29546,I29549,I29552,I29555,I29534,I29534,I29540,I29558,I29561,I29543,I29537,I29607,I29610,I29613,I29616,I29619,I29622,I29625,I29628,I29631,I29634,I2224,I2231);
PAT_14 I_388 (I29613,I29610,I29616,I29628,I29622,I29631,I29619,I29607,I29625,I29634,I29607,I29680,I29683,I29686,I29689,I29692,I29695,I29698,I29701,I29704,I2224,I2231);
PAT_9 I_389 (I29689,I29701,I29680,I29698,I29683,I29686,I29704,I29683,I29692,I29680,I29695,I29750,I29753,I29756,I29759,I29762,I29765,I29768,I29771,I29774,I2224,I2231);
PAT_10 I_390 (I29771,I29768,I29756,I29753,I29774,I29759,I29765,I29753,I29750,I29750,I29762,I29820,I29823,I29826,I29829,I29832,I29835,I29838,I29841,I2224,I2231);
PAT_17 I_391 (I29832,I29841,I29835,I29820,I29826,I29838,I29823,I29823,I29820,I29826,I29829,I29887,I29890,I29893,I29896,I29899,I29902,I29905,I29908,I29911,I29914,I2224,I2231);
PAT_2 I_392 (I29887,I29905,I29902,I29887,I29896,I29911,I29908,I29893,I29914,I29899,I29890,I29960,I29963,I29966,I29969,I29972,I29975,I29978,I29981,I29984,I2224,I2231);
PAT_1 I_393 (I29972,I29960,I29966,I29969,I29960,I29975,I29984,I29963,I29978,I29963,I29981,I30030,I30033,I30036,I30039,I30042,I30045,I30048,I30051,I30054,I2224,I2231);
PAT_4 I_394 (I30042,I30048,I30030,I30033,I30036,I30039,I30051,I30033,I30045,I30030,I30054,I30100,I30103,I30106,I30109,I30112,I30115,I30118,I30121,I30124,I2224,I2231);
PAT_10 I_395 (I30100,I30100,I30124,I30103,I30109,I30118,I30115,I30103,I30121,I30106,I30112,I30170,I30173,I30176,I30179,I30182,I30185,I30188,I30191,I2224,I2231);
PAT_15 I_396 (I30185,I30188,I30176,I30182,I30170,I30170,I30176,I30191,I30179,I30173,I30173,I30237,I30240,I30243,I30246,I30249,I30252,I30255,I30258,I30261,I2224,I2231);
PAT_6 I_397 (I30240,I30237,I30243,I30258,I30240,I30261,I30246,I30252,I30249,I30255,I30237,I30307,I30310,I30313,I30316,I30319,I30322,I30325,I30328,I30331,I30334,I2224,I2231);
PAT_5 I_398 (I30328,I30307,I30313,I30316,I30322,I30325,I30307,I30331,I30310,I30319,I30334,I30380,I30383,I30386,I30389,I30392,I30395,I30398,I30401,I30404,I30407,I2224,I2231);
PAT_12 I_399 (I30407,I30395,I30380,I30404,I30383,I30380,I30386,I30389,I30392,I30398,I30401,I30453,I30456,I30459,I30462,I30465,I30468,I30471,I30474,I2224,I2231);
PAT_4 I_400 (I30459,I30456,I30471,I30474,I30468,I30462,I30453,I30453,I30459,I30465,I30456,I30520,I30523,I30526,I30529,I30532,I30535,I30538,I30541,I30544,I2224,I2231);
PAT_13 I_401 (I30535,I30529,I30541,I30526,I30532,I30520,I30544,I30538,I30523,I30520,I30523,I30590,I30593,I30596,I30599,I30602,I30605,I30608,I30611,I30614,I2224,I2231);
PAT_15 I_402 (I30590,I30602,I30593,I30605,I30590,I30599,I30614,I30611,I30596,I30608,I30593,I30660,I30663,I30666,I30669,I30672,I30675,I30678,I30681,I30684,I2224,I2231);
PAT_13 I_403 (I30669,I30660,I30678,I30663,I30663,I30681,I30672,I30660,I30675,I30684,I30666,I30730,I30733,I30736,I30739,I30742,I30745,I30748,I30751,I30754,I2224,I2231);
PAT_5 I_404 (I30742,I30733,I30739,I30751,I30733,I30754,I30736,I30745,I30730,I30730,I30748,I30800,I30803,I30806,I30809,I30812,I30815,I30818,I30821,I30824,I30827,I2224,I2231);
PAT_10 I_405 (I30824,I30827,I30806,I30812,I30815,I30821,I30803,I30800,I30800,I30809,I30818,I30873,I30876,I30879,I30882,I30885,I30888,I30891,I30894,I2224,I2231);
PAT_4 I_406 (I30888,I30885,I30876,I30894,I30873,I30876,I30882,I30879,I30891,I30873,I30879,I30940,I30943,I30946,I30949,I30952,I30955,I30958,I30961,I30964,I2224,I2231);
PAT_10 I_407 (I30940,I30940,I30964,I30943,I30949,I30958,I30955,I30943,I30961,I30946,I30952,I31010,I31013,I31016,I31019,I31022,I31025,I31028,I31031,I2224,I2231);
PAT_13 I_408 (I31016,I31022,I31016,I31013,I31028,I31031,I31010,I31010,I31025,I31013,I31019,I31077,I31080,I31083,I31086,I31089,I31092,I31095,I31098,I31101,I2224,I2231);
PAT_8 I_409 (I31086,I31098,I31089,I31092,I31101,I31080,I31095,I31077,I31080,I31083,I31077,I31147,I31150,I31153,I31156,I31159,I31162,I31165,I31168,I31171,I2224,I2231);
PAT_17 I_410 (I31171,I31159,I31156,I31150,I31153,I31165,I31147,I31150,I31147,I31162,I31168,I31217,I31220,I31223,I31226,I31229,I31232,I31235,I31238,I31241,I31244,I2224,I2231);
PAT_2 I_411 (I31217,I31235,I31232,I31217,I31226,I31241,I31238,I31223,I31244,I31229,I31220,I31290,I31293,I31296,I31299,I31302,I31305,I31308,I31311,I31314,I2224,I2231);
PAT_10 I_412 (I31290,I31308,I31305,I31293,I31296,I31311,I31302,I31290,I31299,I31314,I31293,I31360,I31363,I31366,I31369,I31372,I31375,I31378,I31381,I2224,I2231);
PAT_11 I_413 (I31369,I31372,I31381,I31375,I31378,I31360,I31360,I31366,I31363,I31363,I31366,I31427,I31430,I31433,I31436,I31439,I31442,I31445,I31448,I31451,I31454,I2224,I2231);
PAT_12 I_414 (I31436,I31451,I31433,I31430,I31439,I31442,I31448,I31427,I31445,I31454,I31427,I31500,I31503,I31506,I31509,I31512,I31515,I31518,I31521,I2224,I2231);
PAT_11 I_415 (I31506,I31509,I31506,I31518,I31521,I31515,I31503,I31512,I31500,I31503,I31500,I31567,I31570,I31573,I31576,I31579,I31582,I31585,I31588,I31591,I31594,I2224,I2231);
PAT_10 I_416 (I31582,I31588,I31579,I31573,I31591,I31576,I31594,I31585,I31567,I31570,I31567,I31640,I31643,I31646,I31649,I31652,I31655,I31658,I31661,I2224,I2231);
PAT_2 I_417 (I31652,I31655,I31646,I31658,I31643,I31640,I31640,I31646,I31661,I31649,I31643,I31707,I31710,I31713,I31716,I31719,I31722,I31725,I31728,I31731,I2224,I2231);
PAT_14 I_418 (I31713,I31716,I31731,I31722,I31707,I31710,I31725,I31719,I31707,I31728,I31710,I31777,I31780,I31783,I31786,I31789,I31792,I31795,I31798,I31801,I2224,I2231);
PAT_10 I_419 (I31780,I31777,I31783,I31801,I31798,I31792,I31780,I31795,I31777,I31789,I31786,I31847,I31850,I31853,I31856,I31859,I31862,I31865,I31868,I2224,I2231);
PAT_6 I_420 (I31868,I31862,I31856,I31850,I31847,I31853,I31847,I31853,I31850,I31859,I31865,I31914,I31917,I31920,I31923,I31926,I31929,I31932,I31935,I31938,I31941,I2224,I2231);
PAT_2 I_421 (I31935,I31941,I31923,I31929,I31914,I31920,I31914,I31926,I31917,I31932,I31938,I31987,I31990,I31993,I31996,I31999,I32002,I32005,I32008,I32011,I2224,I2231);
PAT_14 I_422 (I31993,I31996,I32011,I32002,I31987,I31990,I32005,I31999,I31987,I32008,I31990,I32057,I32060,I32063,I32066,I32069,I32072,I32075,I32078,I32081,I2224,I2231);
PAT_2 I_423 (I32075,I32081,I32066,I32057,I32060,I32060,I32072,I32057,I32078,I32063,I32069,I32127,I32130,I32133,I32136,I32139,I32142,I32145,I32148,I32151,I2224,I2231);
PAT_6 I_424 (I32151,I32127,I32142,I32139,I32145,I32136,I32130,I32148,I32127,I32133,I32130,I32197,I32200,I32203,I32206,I32209,I32212,I32215,I32218,I32221,I32224,I2224,I2231);
PAT_5 I_425 (I32218,I32197,I32203,I32206,I32212,I32215,I32197,I32221,I32200,I32209,I32224,I32270,I32273,I32276,I32279,I32282,I32285,I32288,I32291,I32294,I32297,I2224,I2231);
PAT_6 I_426 (I32288,I32282,I32270,I32276,I32273,I32279,I32285,I32270,I32294,I32291,I32297,I32343,I32346,I32349,I32352,I32355,I32358,I32361,I32364,I32367,I32370,I2224,I2231);
PAT_2 I_427 (I32364,I32370,I32352,I32358,I32343,I32349,I32343,I32355,I32346,I32361,I32367,I32416,I32419,I32422,I32425,I32428,I32431,I32434,I32437,I32440,I2224,I2231);
PAT_14 I_428 (I32422,I32425,I32440,I32431,I32416,I32419,I32434,I32428,I32416,I32437,I32419,I32486,I32489,I32492,I32495,I32498,I32501,I32504,I32507,I32510,I2224,I2231);
PAT_6 I_429 (I32486,I32489,I32510,I32495,I32486,I32492,I32498,I32501,I32504,I32489,I32507,I32556,I32559,I32562,I32565,I32568,I32571,I32574,I32577,I32580,I32583,I2224,I2231);
PAT_17 I_430 (I32568,I32571,I32577,I32565,I32559,I32580,I32574,I32556,I32583,I32562,I32556,I32629,I32632,I32635,I32638,I32641,I32644,I32647,I32650,I32653,I32656,I2224,I2231);
PAT_13 I_431 (I32647,I32650,I32635,I32629,I32641,I32653,I32632,I32644,I32629,I32656,I32638,I32702,I32705,I32708,I32711,I32714,I32717,I32720,I32723,I32726,I2224,I2231);
PAT_2 I_432 (I32720,I32714,I32711,I32717,I32702,I32726,I32705,I32723,I32702,I32708,I32705,I32772,I32775,I32778,I32781,I32784,I32787,I32790,I32793,I32796,I2224,I2231);
PAT_7 I_433 (I32796,I32772,I32778,I32775,I32775,I32784,I32787,I32772,I32790,I32793,I32781,I32842,I32845,I32848,I32851,I32854,I32857,I32860,I32863,I32866,I2224,I2231);
PAT_17 I_434 (I32854,I32848,I32857,I32842,I32860,I32863,I32845,I32866,I32851,I32845,I32842,I32912,I32915,I32918,I32921,I32924,I32927,I32930,I32933,I32936,I32939,I2224,I2231);
PAT_9 I_435 (I32933,I32915,I32921,I32936,I32918,I32930,I32912,I32924,I32912,I32939,I32927,I32985,I32988,I32991,I32994,I32997,I33000,I33003,I33006,I33009,I2224,I2231);
PAT_10 I_436 (I33006,I33003,I32991,I32988,I33009,I32994,I33000,I32988,I32985,I32985,I32997,I33055,I33058,I33061,I33064,I33067,I33070,I33073,I33076,I2224,I2231);
PAT_12 I_437 (I33061,I33055,I33055,I33067,I33070,I33058,I33058,I33073,I33076,I33061,I33064,I33122,I33125,I33128,I33131,I33134,I33137,I33140,I33143,I2224,I2231);
PAT_1 I_438 (I33137,I33125,I33140,I33131,I33122,I33125,I33134,I33122,I33143,I33128,I33128,I33189,I33192,I33195,I33198,I33201,I33204,I33207,I33210,I33213,I2224,I2231);
PAT_15 I_439 (I33192,I33201,I33189,I33204,I33198,I33192,I33213,I33210,I33207,I33195,I33189,I33259,I33262,I33265,I33268,I33271,I33274,I33277,I33280,I33283,I2224,I2231);
PAT_9 I_440 (I33259,I33280,I33268,I33262,I33274,I33262,I33277,I33283,I33265,I33259,I33271,I33329,I33332,I33335,I33338,I33341,I33344,I33347,I33350,I33353,I2224,I2231);
PAT_13 I_441 (I33329,I33350,I33332,I33347,I33341,I33338,I33353,I33329,I33335,I33344,I33332,I33399,I33402,I33405,I33408,I33411,I33414,I33417,I33420,I33423,I2224,I2231);
PAT_5 I_442 (I33411,I33402,I33408,I33420,I33402,I33423,I33405,I33414,I33399,I33399,I33417,I33469,I33472,I33475,I33478,I33481,I33484,I33487,I33490,I33493,I33496,I2224,I2231);
PAT_13 I_443 (I33475,I33484,I33469,I33472,I33493,I33478,I33490,I33469,I33487,I33496,I33481,I33542,I33545,I33548,I33551,I33554,I33557,I33560,I33563,I33566,I2224,I2231);
PAT_11 I_444 (I33542,I33554,I33557,I33548,I33545,I33566,I33545,I33563,I33551,I33542,I33560,I33612,I33615,I33618,I33621,I33624,I33627,I33630,I33633,I33636,I33639,I2224,I2231);
PAT_4 I_445 (I33618,I33639,I33612,I33630,I33621,I33612,I33633,I33615,I33624,I33636,I33627,I33685,I33688,I33691,I33694,I33697,I33700,I33703,I33706,I33709,I2224,I2231);
PAT_5 I_446 (I33706,I33688,I33688,I33700,I33703,I33697,I33694,I33685,I33691,I33685,I33709,I33755,I33758,I33761,I33764,I33767,I33770,I33773,I33776,I33779,I33782,I2224,I2231);
PAT_10 I_447 (I33779,I33782,I33761,I33767,I33770,I33776,I33758,I33755,I33755,I33764,I33773,I33828,I33831,I33834,I33837,I33840,I33843,I33846,I33849,I2224,I2231);
PAT_14 I_448 (I33828,I33849,I33834,I33843,I33840,I33846,I33837,I33831,I33831,I33834,I33828,I33895,I33898,I33901,I33904,I33907,I33910,I33913,I33916,I33919,I2224,I2231);
PAT_9 I_449 (I33904,I33916,I33895,I33913,I33898,I33901,I33919,I33898,I33907,I33895,I33910,I33965,I33968,I33971,I33974,I33977,I33980,I33983,I33986,I33989,I2224,I2231);
PAT_11 I_450 (I33977,I33983,I33989,I33986,I33974,I33968,I33968,I33965,I33980,I33965,I33971,I34035,I34038,I34041,I34044,I34047,I34050,I34053,I34056,I34059,I34062,I2224,I2231);
PAT_13 I_451 (I34035,I34038,I34047,I34059,I34062,I34050,I34056,I34044,I34053,I34041,I34035,I34108,I34111,I34114,I34117,I34120,I34123,I34126,I34129,I34132,I2224,I2231);
PAT_7 I_452 (I34117,I34120,I34108,I34123,I34129,I34114,I34111,I34132,I34111,I34108,I34126,I34178,I34181,I34184,I34187,I34190,I34193,I34196,I34199,I34202,I2224,I2231);
PAT_5 I_453 (I34184,I34178,I34187,I34196,I34190,I34202,I34199,I34181,I34193,I34181,I34178,I34248,I34251,I34254,I34257,I34260,I34263,I34266,I34269,I34272,I34275,I2224,I2231);
PAT_4 I_454 (I34266,I34272,I34275,I34254,I34257,I34269,I34251,I34248,I34260,I34263,I34248,I34321,I34324,I34327,I34330,I34333,I34336,I34339,I34342,I34345,I2224,I2231);
PAT_6 I_455 (I34321,I34327,I34324,I34336,I34339,I34333,I34345,I34342,I34321,I34330,I34324,I34391,I34394,I34397,I34400,I34403,I34406,I34409,I34412,I34415,I34418,I2224,I2231);
PAT_11 I_456 (I34391,I34406,I34391,I34403,I34400,I34418,I34415,I34412,I34409,I34394,I34397,I34464,I34467,I34470,I34473,I34476,I34479,I34482,I34485,I34488,I34491,I2224,I2231);
PAT_2 I_457 (I34464,I34488,I34476,I34470,I34479,I34482,I34467,I34491,I34485,I34473,I34464,I34537,I34540,I34543,I34546,I34549,I34552,I34555,I34558,I34561,I2224,I2231);
PAT_11 I_458 (I34540,I34552,I34537,I34549,I34546,I34558,I34555,I34540,I34561,I34543,I34537,I34607,I34610,I34613,I34616,I34619,I34622,I34625,I34628,I34631,I34634,I2224,I2231);
PAT_14 I_459 (I34628,I34616,I34610,I34631,I34622,I34625,I34613,I34634,I34619,I34607,I34607,I34680,I34683,I34686,I34689,I34692,I34695,I34698,I34701,I34704,I2224,I2231);
PAT_17 I_460 (I34695,I34683,I34704,I34680,I34701,I34689,I34686,I34698,I34692,I34683,I34680,I34750,I34753,I34756,I34759,I34762,I34765,I34768,I34771,I34774,I34777,I2224,I2231);
PAT_2 I_461 (I34750,I34768,I34765,I34750,I34759,I34774,I34771,I34756,I34777,I34762,I34753,I34823,I34826,I34829,I34832,I34835,I34838,I34841,I34844,I34847,I2224,I2231);
PAT_11 I_462 (I34826,I34838,I34823,I34835,I34832,I34844,I34841,I34826,I34847,I34829,I34823,I34893,I34896,I34899,I34902,I34905,I34908,I34911,I34914,I34917,I34920,I2224,I2231);
PAT_4 I_463 (I34899,I34920,I34893,I34911,I34902,I34893,I34914,I34896,I34905,I34917,I34908,I34966,I34969,I34972,I34975,I34978,I34981,I34984,I34987,I34990,I2224,I2231);
PAT_9 I_464 (I34987,I34969,I34972,I34981,I34984,I34966,I34975,I34969,I34990,I34966,I34978,I35036,I35039,I35042,I35045,I35048,I35051,I35054,I35057,I35060,I2224,I2231);
PAT_5 I_465 (I35057,I35036,I35051,I35036,I35042,I35045,I35039,I35039,I35054,I35048,I35060,I35106,I35109,I35112,I35115,I35118,I35121,I35124,I35127,I35130,I35133,I2224,I2231);
PAT_10 I_466 (I35130,I35133,I35112,I35118,I35121,I35127,I35109,I35106,I35106,I35115,I35124,I35179,I35182,I35185,I35188,I35191,I35194,I35197,I35200,I2224,I2231);
PAT_9 I_467 (I35191,I35179,I35182,I35185,I35179,I35185,I35188,I35182,I35200,I35194,I35197,I35246,I35249,I35252,I35255,I35258,I35261,I35264,I35267,I35270,I2224,I2231);
PAT_4 I_468 (I35246,I35270,I35264,I35252,I35249,I35267,I35249,I35246,I35261,I35255,I35258,I35316,I35319,I35322,I35325,I35328,I35331,I35334,I35337,I35340,I2224,I2231);
PAT_5 I_469 (I35337,I35319,I35319,I35331,I35334,I35328,I35325,I35316,I35322,I35316,I35340,I35386,I35389,I35392,I35395,I35398,I35401,I35404,I35407,I35410,I35413,I2224,I2231);
PAT_17 I_470 (I35413,I35389,I35392,I35395,I35386,I35398,I35386,I35410,I35404,I35401,I35407,I35459,I35462,I35465,I35468,I35471,I35474,I35477,I35480,I35483,I35486,I2224,I2231);
PAT_11 I_471 (I35471,I35480,I35486,I35462,I35459,I35477,I35468,I35474,I35465,I35483,I35459,I35532,I35535,I35538,I35541,I35544,I35547,I35550,I35553,I35556,I35559,I2224,I2231);
PAT_12 I_472 (I35541,I35556,I35538,I35535,I35544,I35547,I35553,I35532,I35550,I35559,I35532,I35605,I35608,I35611,I35614,I35617,I35620,I35623,I35626,I2224,I2231);
PAT_1 I_473 (I35620,I35608,I35623,I35614,I35605,I35608,I35617,I35605,I35626,I35611,I35611,I35672,I35675,I35678,I35681,I35684,I35687,I35690,I35693,I35696,I2224,I2231);
PAT_3 I_474 (I35681,I35675,I35675,I35678,I35690,I35693,I35696,I35684,I35672,I35672,I35687,I35742,I35745,I35748,I35751,I35754,I35757,I35760,I35763,I35766,I35769,I2224,I2231);
PAT_17 I_475 (I35754,I35769,I35748,I35757,I35745,I35760,I35742,I35751,I35763,I35742,I35766,I35815,I35818,I35821,I35824,I35827,I35830,I35833,I35836,I35839,I35842,I2224,I2231);
PAT_11 I_476 (I35827,I35836,I35842,I35818,I35815,I35833,I35824,I35830,I35821,I35839,I35815,I35888,I35891,I35894,I35897,I35900,I35903,I35906,I35909,I35912,I35915,I2224,I2231);
PAT_6 I_477 (I35888,I35915,I35903,I35912,I35906,I35900,I35891,I35909,I35897,I35894,I35888,I35961,I35964,I35967,I35970,I35973,I35976,I35979,I35982,I35985,I35988,I2224,I2231);
PAT_17 I_478 (I35973,I35976,I35982,I35970,I35964,I35985,I35979,I35961,I35988,I35967,I35961,I36034,I36037,I36040,I36043,I36046,I36049,I36052,I36055,I36058,I36061,I2224,I2231);
PAT_2 I_479 (I36034,I36052,I36049,I36034,I36043,I36058,I36055,I36040,I36061,I36046,I36037,I36107,I36110,I36113,I36116,I36119,I36122,I36125,I36128,I36131,I2224,I2231);
PAT_4 I_480 (I36107,I36113,I36131,I36125,I36122,I36119,I36110,I36128,I36107,I36110,I36116,I36177,I36180,I36183,I36186,I36189,I36192,I36195,I36198,I36201,I2224,I2231);
PAT_14 I_481 (I36180,I36195,I36192,I36177,I36189,I36180,I36177,I36183,I36198,I36186,I36201,I36247,I36250,I36253,I36256,I36259,I36262,I36265,I36268,I36271,I2224,I2231);
PAT_9 I_482 (I36256,I36268,I36247,I36265,I36250,I36253,I36271,I36250,I36259,I36247,I36262,I36317,I36320,I36323,I36326,I36329,I36332,I36335,I36338,I36341,I2224,I2231);
PAT_5 I_483 (I36338,I36317,I36332,I36317,I36323,I36326,I36320,I36320,I36335,I36329,I36341,I36387,I36390,I36393,I36396,I36399,I36402,I36405,I36408,I36411,I36414,I2224,I2231);
PAT_9 I_484 (I36402,I36399,I36408,I36405,I36396,I36387,I36393,I36414,I36390,I36411,I36387,I36460,I36463,I36466,I36469,I36472,I36475,I36478,I36481,I36484,I2224,I2231);
PAT_1 I_485 (I36460,I36478,I36460,I36472,I36463,I36469,I36475,I36481,I36484,I36466,I36463,I36530,I36533,I36536,I36539,I36542,I36545,I36548,I36551,I36554,I2224,I2231);
PAT_8 I_486 (I36551,I36533,I36539,I36530,I36548,I36542,I36545,I36530,I36554,I36536,I36533,I36600,I36603,I36606,I36609,I36612,I36615,I36618,I36621,I36624,I2224,I2231);
PAT_2 I_487 (I36603,I36618,I36624,I36600,I36612,I36615,I36603,I36621,I36606,I36609,I36600,I36670,I36673,I36676,I36679,I36682,I36685,I36688,I36691,I36694,I2224,I2231);
PAT_9 I_488 (I36685,I36694,I36670,I36676,I36679,I36688,I36673,I36682,I36691,I36673,I36670,I36740,I36743,I36746,I36749,I36752,I36755,I36758,I36761,I36764,I2224,I2231);
PAT_2 I_489 (I36755,I36758,I36749,I36764,I36740,I36743,I36746,I36743,I36761,I36752,I36740,I36810,I36813,I36816,I36819,I36822,I36825,I36828,I36831,I36834,I2224,I2231);
PAT_7 I_490 (I36834,I36810,I36816,I36813,I36813,I36822,I36825,I36810,I36828,I36831,I36819,I36880,I36883,I36886,I36889,I36892,I36895,I36898,I36901,I36904,I2224,I2231);
PAT_10 I_491 (I36880,I36883,I36880,I36901,I36889,I36892,I36883,I36904,I36895,I36886,I36898,I36950,I36953,I36956,I36959,I36962,I36965,I36968,I36971,I2224,I2231);
PAT_6 I_492 (I36971,I36965,I36959,I36953,I36950,I36956,I36950,I36956,I36953,I36962,I36968,I37017,I37020,I37023,I37026,I37029,I37032,I37035,I37038,I37041,I37044,I2224,I2231);
PAT_9 I_493 (I37017,I37044,I37041,I37023,I37029,I37020,I37032,I37017,I37035,I37026,I37038,I37090,I37093,I37096,I37099,I37102,I37105,I37108,I37111,I37114,I2224,I2231);
PAT_15 I_494 (I37102,I37111,I37114,I37093,I37108,I37096,I37099,I37090,I37105,I37090,I37093,I37160,I37163,I37166,I37169,I37172,I37175,I37178,I37181,I37184,I2224,I2231);
PAT_2 I_495 (I37163,I37163,I37166,I37172,I37160,I37160,I37169,I37184,I37178,I37181,I37175,I37230,I37233,I37236,I37239,I37242,I37245,I37248,I37251,I37254,I2224,I2231);
PAT_13 I_496 (I37239,I37233,I37230,I37251,I37242,I37245,I37233,I37236,I37248,I37254,I37230,I37300,I37303,I37306,I37309,I37312,I37315,I37318,I37321,I37324,I2224,I2231);
PAT_2 I_497 (I37318,I37312,I37309,I37315,I37300,I37324,I37303,I37321,I37300,I37306,I37303,I37370,I37373,I37376,I37379,I37382,I37385,I37388,I37391,I37394,I2224,I2231);
PAT_4 I_498 (I37370,I37376,I37394,I37388,I37385,I37382,I37373,I37391,I37370,I37373,I37379,I37440,I37443,I37446,I37449,I37452,I37455,I37458,I37461,I37464,I2224,I2231);
PAT_9 I_499 (I37461,I37443,I37446,I37455,I37458,I37440,I37449,I37443,I37464,I37440,I37452,I37510,I37513,I37516,I37519,I37522,I37525,I37528,I37531,I37534,I2224,I2231);
PAT_1 I_500 (I37510,I37528,I37510,I37522,I37513,I37519,I37525,I37531,I37534,I37516,I37513,I37580,I37583,I37586,I37589,I37592,I37595,I37598,I37601,I37604,I2224,I2231);
PAT_2 I_501 (I37580,I37586,I37580,I37595,I37583,I37583,I37589,I37592,I37598,I37604,I37601,I37650,I37653,I37656,I37659,I37662,I37665,I37668,I37671,I37674,I2224,I2231);
PAT_10 I_502 (I37650,I37668,I37665,I37653,I37656,I37671,I37662,I37650,I37659,I37674,I37653,I37720,I37723,I37726,I37729,I37732,I37735,I37738,I37741,I2224,I2231);
PAT_4 I_503 (I37735,I37732,I37723,I37741,I37720,I37723,I37729,I37726,I37738,I37720,I37726,I37787,I37790,I37793,I37796,I37799,I37802,I37805,I37808,I37811,I2224,I2231);
PAT_5 I_504 (I37808,I37790,I37790,I37802,I37805,I37799,I37796,I37787,I37793,I37787,I37811,I37857,I37860,I37863,I37866,I37869,I37872,I37875,I37878,I37881,I37884,I2224,I2231);
PAT_15 I_505 (I37875,I37860,I37857,I37857,I37872,I37869,I37881,I37866,I37878,I37863,I37884,I37930,I37933,I37936,I37939,I37942,I37945,I37948,I37951,I37954,I2224,I2231);
PAT_12 I_506 (I37948,I37951,I37954,I37942,I37939,I37933,I37930,I37945,I37936,I37930,I37933,I38000,I38003,I38006,I38009,I38012,I38015,I38018,I38021,I2224,I2231);
PAT_2 I_507 (I38018,I38012,I38021,I38015,I38009,I38006,I38000,I38000,I38006,I38003,I38003,I38067,I38070,I38073,I38076,I38079,I38082,I38085,I38088,I38091,I2224,I2231);
PAT_10 I_508 (I38067,I38085,I38082,I38070,I38073,I38088,I38079,I38067,I38076,I38091,I38070,I38137,I38140,I38143,I38146,I38149,I38152,I38155,I38158,I2224,I2231);
PAT_11 I_509 (I38146,I38149,I38158,I38152,I38155,I38137,I38137,I38143,I38140,I38140,I38143,I38204,I38207,I38210,I38213,I38216,I38219,I38222,I38225,I38228,I38231,I2224,I2231);
PAT_2 I_510 (I38204,I38228,I38216,I38210,I38219,I38222,I38207,I38231,I38225,I38213,I38204,I38277,I38280,I38283,I38286,I38289,I38292,I38295,I38298,I38301,I2224,I2231);
PAT_11 I_511 (I38280,I38292,I38277,I38289,I38286,I38298,I38295,I38280,I38301,I38283,I38277,I38347,I38350,I38353,I38356,I38359,I38362,I38365,I38368,I38371,I38374,I2224,I2231);
PAT_6 I_512 (I38347,I38374,I38362,I38371,I38365,I38359,I38350,I38368,I38356,I38353,I38347,I38420,I38423,I38426,I38429,I38432,I38435,I38438,I38441,I38444,I38447,I2224,I2231);
PAT_8 I_513 (I38429,I38435,I38426,I38438,I38420,I38423,I38441,I38420,I38447,I38444,I38432,I38493,I38496,I38499,I38502,I38505,I38508,I38511,I38514,I38517,I2224,I2231);
PAT_13 I_514 (I38505,I38514,I38496,I38517,I38499,I38493,I38493,I38502,I38511,I38508,I38496,I38563,I38566,I38569,I38572,I38575,I38578,I38581,I38584,I38587,I2224,I2231);
PAT_8 I_515 (I38572,I38584,I38575,I38578,I38587,I38566,I38581,I38563,I38566,I38569,I38563,I38633,I38636,I38639,I38642,I38645,I38648,I38651,I38654,I38657,I2224,I2231);
PAT_17 I_516 (I38657,I38645,I38642,I38636,I38639,I38651,I38633,I38636,I38633,I38648,I38654,I38703,I38706,I38709,I38712,I38715,I38718,I38721,I38724,I38727,I38730,I2224,I2231);
PAT_6 I_517 (I38703,I38721,I38709,I38712,I38718,I38703,I38715,I38706,I38727,I38730,I38724,I38776,I38779,I38782,I38785,I38788,I38791,I38794,I38797,I38800,I38803,I2224,I2231);
PAT_9 I_518 (I38776,I38803,I38800,I38782,I38788,I38779,I38791,I38776,I38794,I38785,I38797,I38849,I38852,I38855,I38858,I38861,I38864,I38867,I38870,I38873,I2224,I2231);
PAT_4 I_519 (I38849,I38873,I38867,I38855,I38852,I38870,I38852,I38849,I38864,I38858,I38861,I38919,I38922,I38925,I38928,I38931,I38934,I38937,I38940,I38943,I2224,I2231);
PAT_11 I_520 (I38931,I38940,I38922,I38934,I38919,I38922,I38919,I38928,I38943,I38937,I38925,I38989,I38992,I38995,I38998,I39001,I39004,I39007,I39010,I39013,I39016,I2224,I2231);
PAT_5 I_521 (I39010,I38989,I39016,I39004,I39001,I39013,I38995,I38989,I39007,I38992,I38998,I39062,I39065,I39068,I39071,I39074,I39077,I39080,I39083,I39086,I39089,I2224,I2231);
PAT_13 I_522 (I39068,I39077,I39062,I39065,I39086,I39071,I39083,I39062,I39080,I39089,I39074,I39135,I39138,I39141,I39144,I39147,I39150,I39153,I39156,I39159,I2224,I2231);
PAT_8 I_523 (I39144,I39156,I39147,I39150,I39159,I39138,I39153,I39135,I39138,I39141,I39135,I39205,I39208,I39211,I39214,I39217,I39220,I39223,I39226,I39229,I2224,I2231);
PAT_11 I_524 (I39226,I39217,I39205,I39208,I39223,I39211,I39214,I39205,I39229,I39220,I39208,I39275,I39278,I39281,I39284,I39287,I39290,I39293,I39296,I39299,I39302,I2224,I2231);
PAT_13 I_525 (I39275,I39278,I39287,I39299,I39302,I39290,I39296,I39284,I39293,I39281,I39275,I39348,I39351,I39354,I39357,I39360,I39363,I39366,I39369,I39372,I2224,I2231);
PAT_3 I_526 (I39372,I39351,I39366,I39354,I39360,I39369,I39348,I39357,I39348,I39351,I39363,I39418,I39421,I39424,I39427,I39430,I39433,I39436,I39439,I39442,I39445,I2224,I2231);
PAT_9 I_527 (I39418,I39442,I39424,I39439,I39427,I39421,I39436,I39445,I39418,I39430,I39433,I39491,I39494,I39497,I39500,I39503,I39506,I39509,I39512,I39515,I2224,I2231);
PAT_3 I_528 (I39515,I39494,I39497,I39509,I39500,I39494,I39503,I39491,I39512,I39491,I39506,I39561,I39564,I39567,I39570,I39573,I39576,I39579,I39582,I39585,I39588,I2224,I2231);
PAT_5 I_529 (I39582,I39573,I39564,I39561,I39567,I39588,I39579,I39570,I39561,I39585,I39576,I39634,I39637,I39640,I39643,I39646,I39649,I39652,I39655,I39658,I39661,I2224,I2231);
PAT_7 I_530 (I39652,I39655,I39661,I39658,I39643,I39640,I39634,I39646,I39634,I39637,I39649,I39707,I39710,I39713,I39716,I39719,I39722,I39725,I39728,I39731,I2224,I2231);
PAT_5 I_531 (I39713,I39707,I39716,I39725,I39719,I39731,I39728,I39710,I39722,I39710,I39707,I39777,I39780,I39783,I39786,I39789,I39792,I39795,I39798,I39801,I39804,I2224,I2231);
PAT_3 I_532 (I39789,I39777,I39804,I39798,I39801,I39777,I39792,I39780,I39783,I39786,I39795,I39850,I39853,I39856,I39859,I39862,I39865,I39868,I39871,I39874,I39877,I2224,I2231);
PAT_2 I_533 (I39877,I39862,I39853,I39850,I39874,I39865,I39859,I39868,I39850,I39871,I39856,I39923,I39926,I39929,I39932,I39935,I39938,I39941,I39944,I39947,I2224,I2231);
PAT_5 I_534 (I39944,I39923,I39923,I39935,I39932,I39941,I39929,I39938,I39947,I39926,I39926,I39993,I39996,I39999,I40002,I40005,I40008,I40011,I40014,I40017,I40020,I2224,I2231);
PAT_10 I_535 (I40017,I40020,I39999,I40005,I40008,I40014,I39996,I39993,I39993,I40002,I40011,I40066,I40069,I40072,I40075,I40078,I40081,I40084,I40087,I2224,I2231);
PAT_4 I_536 (I40081,I40078,I40069,I40087,I40066,I40069,I40075,I40072,I40084,I40066,I40072,I40133,I40136,I40139,I40142,I40145,I40148,I40151,I40154,I40157,I2224,I2231);
PAT_8 I_537 (I40145,I40133,I40154,I40139,I40136,I40157,I40142,I40151,I40136,I40133,I40148,I40203,I40206,I40209,I40212,I40215,I40218,I40221,I40224,I40227,I2224,I2231);
PAT_10 I_538 (I40209,I40203,I40206,I40227,I40221,I40206,I40215,I40203,I40224,I40218,I40212,I40273,I40276,I40279,I40282,I40285,I40288,I40291,I40294,I2224,I2231);
PAT_6 I_539 (I40294,I40288,I40282,I40276,I40273,I40279,I40273,I40279,I40276,I40285,I40291,I40340,I40343,I40346,I40349,I40352,I40355,I40358,I40361,I40364,I40367,I2224,I2231);
PAT_2 I_540 (I40361,I40367,I40349,I40355,I40340,I40346,I40340,I40352,I40343,I40358,I40364,I40413,I40416,I40419,I40422,I40425,I40428,I40431,I40434,I40437,I2224,I2231);
PAT_11 I_541 (I40416,I40428,I40413,I40425,I40422,I40434,I40431,I40416,I40437,I40419,I40413,I40483,I40486,I40489,I40492,I40495,I40498,I40501,I40504,I40507,I40510,I2224,I2231);
PAT_12 I_542 (I40492,I40507,I40489,I40486,I40495,I40498,I40504,I40483,I40501,I40510,I40483,I40556,I40559,I40562,I40565,I40568,I40571,I40574,I40577,I2224,I2231);
PAT_9 I_543 (I40565,I40571,I40556,I40562,I40568,I40559,I40556,I40559,I40577,I40562,I40574,I40623,I40626,I40629,I40632,I40635,I40638,I40641,I40644,I40647,I2224,I2231);
PAT_11 I_544 (I40635,I40641,I40647,I40644,I40632,I40626,I40626,I40623,I40638,I40623,I40629,I40693,I40696,I40699,I40702,I40705,I40708,I40711,I40714,I40717,I40720,I2224,I2231);
PAT_6 I_545 (I40693,I40720,I40708,I40717,I40711,I40705,I40696,I40714,I40702,I40699,I40693,I40766,I40769,I40772,I40775,I40778,I40781,I40784,I40787,I40790,I40793,I2224,I2231);
PAT_5 I_546 (I40787,I40766,I40772,I40775,I40781,I40784,I40766,I40790,I40769,I40778,I40793,I40839,I40842,I40845,I40848,I40851,I40854,I40857,I40860,I40863,I40866,I2224,I2231);
PAT_13 I_547 (I40845,I40854,I40839,I40842,I40863,I40848,I40860,I40839,I40857,I40866,I40851,I40912,I40915,I40918,I40921,I40924,I40927,I40930,I40933,I40936,I2224,I2231);
PAT_8 I_548 (I40921,I40933,I40924,I40927,I40936,I40915,I40930,I40912,I40915,I40918,I40912,I40982,I40985,I40988,I40991,I40994,I40997,I41000,I41003,I41006,I2224,I2231);
PAT_5 I_549 (I40988,I41006,I40982,I41003,I40991,I40994,I40985,I40982,I40985,I40997,I41000,I41052,I41055,I41058,I41061,I41064,I41067,I41070,I41073,I41076,I41079,I2224,I2231);
PAT_14 I_550 (I41073,I41058,I41052,I41076,I41079,I41052,I41070,I41055,I41061,I41064,I41067,I41125,I41128,I41131,I41134,I41137,I41140,I41143,I41146,I41149,I2224,I2231);
PAT_13 I_551 (I41134,I41149,I41128,I41137,I41125,I41128,I41143,I41131,I41125,I41146,I41140,I41195,I41198,I41201,I41204,I41207,I41210,I41213,I41216,I41219,I2224,I2231);
PAT_4 I_552 (I41204,I41207,I41219,I41201,I41216,I41213,I41198,I41210,I41198,I41195,I41195,I41265,I41268,I41271,I41274,I41277,I41280,I41283,I41286,I41289,I2224,I2231);
PAT_10 I_553 (I41265,I41265,I41289,I41268,I41274,I41283,I41280,I41268,I41286,I41271,I41277,I41335,I41338,I41341,I41344,I41347,I41350,I41353,I41356,I2224,I2231);
PAT_16 I_554 (I41338,I41347,I41353,I41341,I41341,I41335,I41350,I41344,I41335,I41338,I41356,I41402,I41405,I41408,I41411,I41414,I41417,I41420,I41423,I41426,I41429,I2224,I2231);
PAT_9 I_555 (I41420,I41402,I41402,I41411,I41408,I41426,I41429,I41405,I41423,I41417,I41414,I41475,I41478,I41481,I41484,I41487,I41490,I41493,I41496,I41499,I2224,I2231);
PAT_13 I_556 (I41475,I41496,I41478,I41493,I41487,I41484,I41499,I41475,I41481,I41490,I41478,I41545,I41548,I41551,I41554,I41557,I41560,I41563,I41566,I41569,I2224,I2231);
PAT_10 I_557 (I41566,I41560,I41554,I41548,I41569,I41548,I41557,I41545,I41545,I41563,I41551,I41615,I41618,I41621,I41624,I41627,I41630,I41633,I41636,I2224,I2231);
PAT_9 I_558 (I1825,I1769,I1625,I2033,I2057,I1649,I1985,I1497,I1681,I2105,I1457,I41682,I41685,I41688,I41691,I41694,I41697,I41700,I41703,I41706,I2224,I2231);
PAT_2 I_559 (I41697,I41700,I41691,I41706,I41682,I41685,I41688,I41685,I41703,I41694,I41682,I41752,I41755,I41758,I41761,I41764,I41767,I41770,I41773,I41776,I2224,I2231);
PAT_9 I_560 (I41767,I41776,I41752,I41758,I41761,I41770,I41755,I41764,I41773,I41755,I41752,I41822,I41825,I41828,I41831,I41834,I41837,I41840,I41843,I41846,I2224,I2231);
PAT_17 I_561 (I41825,I41831,I41846,I41837,I41840,I41828,I41822,I41834,I41822,I41825,I41843,I41892,I41895,I41898,I41901,I41904,I41907,I41910,I41913,I41916,I41919,I2224,I2231);
PAT_6 I_562 (I41892,I41910,I41898,I41901,I41907,I41892,I41904,I41895,I41916,I41919,I41913,I41965,I41968,I41971,I41974,I41977,I41980,I41983,I41986,I41989,I41992,I2224,I2231);
PAT_4 I_563 (I41965,I41980,I41968,I41971,I41974,I41965,I41992,I41983,I41986,I41977,I41989,I42038,I42041,I42044,I42047,I42050,I42053,I42056,I42059,I42062,I2224,I2231);
PAT_12 I_564 (I42038,I42041,I42059,I42062,I42053,I42044,I42050,I42047,I42038,I42056,I42041,I42108,I42111,I42114,I42117,I42120,I42123,I42126,I42129,I2224,I2231);
PAT_4 I_565 (I42114,I42111,I42126,I42129,I42123,I42117,I42108,I42108,I42114,I42120,I42111,I42175,I42178,I42181,I42184,I42187,I42190,I42193,I42196,I42199,I2224,I2231);
PAT_14 I_566 (I42178,I42193,I42190,I42175,I42187,I42178,I42175,I42181,I42196,I42184,I42199,I42245,I42248,I42251,I42254,I42257,I42260,I42263,I42266,I42269,I2224,I2231);
PAT_8 I_567 (I42251,I42254,I42248,I42260,I42269,I42248,I42245,I42266,I42245,I42257,I42263,I42315,I42318,I42321,I42324,I42327,I42330,I42333,I42336,I42339,I2224,I2231);
PAT_11 I_568 (I42336,I42327,I42315,I42318,I42333,I42321,I42324,I42315,I42339,I42330,I42318,I42385,I42388,I42391,I42394,I42397,I42400,I42403,I42406,I42409,I42412,I2224,I2231);
PAT_13 I_569 (I42385,I42388,I42397,I42409,I42412,I42400,I42406,I42394,I42403,I42391,I42385,I42458,I42461,I42464,I42467,I42470,I42473,I42476,I42479,I42482,I2224,I2231);
PAT_17 I_570 (I42482,I42470,I42479,I42476,I42467,I42458,I42461,I42464,I42458,I42473,I42461,I42528,I42531,I42534,I42537,I42540,I42543,I42546,I42549,I42552,I42555,I2224,I2231);
PAT_5 I_571 (I42540,I42534,I42531,I42552,I42537,I42543,I42546,I42528,I42528,I42549,I42555,I42601,I42604,I42607,I42610,I42613,I42616,I42619,I42622,I42625,I42628,I2224,I2231);
PAT_2 I_572 (I42616,I42601,I42613,I42607,I42622,I42604,I42619,I42610,I42625,I42628,I42601,I42674,I42677,I42680,I42683,I42686,I42689,I42692,I42695,I42698,I2224,I2231);
PAT_9 I_573 (I42689,I42698,I42674,I42680,I42683,I42692,I42677,I42686,I42695,I42677,I42674,I42744,I42747,I42750,I42753,I42756,I42759,I42762,I42765,I42768,I2224,I2231);
PAT_4 I_574 (I42744,I42768,I42762,I42750,I42747,I42765,I42747,I42744,I42759,I42753,I42756,I42814,I42817,I42820,I42823,I42826,I42829,I42832,I42835,I42838,I2224,I2231);
PAT_13 I_575 (I42829,I42823,I42835,I42820,I42826,I42814,I42838,I42832,I42817,I42814,I42817,I42884,I42887,I42890,I42893,I42896,I42899,I42902,I42905,I42908,I2224,I2231);
PAT_9 I_576 (I42905,I42887,I42887,I42884,I42908,I42890,I42893,I42884,I42896,I42902,I42899,I42954,I42957,I42960,I42963,I42966,I42969,I42972,I42975,I42978,I2224,I2231);
PAT_11 I_577 (I42966,I42972,I42978,I42975,I42963,I42957,I42957,I42954,I42969,I42954,I42960,I43024,I43027,I43030,I43033,I43036,I43039,I43042,I43045,I43048,I43051,I2224,I2231);
PAT_17 I_578 (I43036,I43027,I43051,I43024,I43033,I43045,I43042,I43039,I43024,I43048,I43030,I43097,I43100,I43103,I43106,I43109,I43112,I43115,I43118,I43121,I43124,I2224,I2231);
PAT_4 I_579 (I43106,I43097,I43115,I43112,I43124,I43121,I43100,I43097,I43103,I43109,I43118,I43170,I43173,I43176,I43179,I43182,I43185,I43188,I43191,I43194,I2224,I2231);
PAT_13 I_580 (I43185,I43179,I43191,I43176,I43182,I43170,I43194,I43188,I43173,I43170,I43173,I43240,I43243,I43246,I43249,I43252,I43255,I43258,I43261,I43264,I2224,I2231);
PAT_15 I_581 (I43240,I43252,I43243,I43255,I43240,I43249,I43264,I43261,I43246,I43258,I43243,I43310,I43313,I43316,I43319,I43322,I43325,I43328,I43331,I43334,I2224,I2231);
PAT_14 I_582 (I43313,I43313,I43334,I43310,I43316,I43310,I43325,I43322,I43331,I43319,I43328,I43380,I43383,I43386,I43389,I43392,I43395,I43398,I43401,I43404,I2224,I2231);
PAT_11 I_583 (I43392,I43389,I43386,I43380,I43383,I43383,I43395,I43380,I43401,I43404,I43398,I43450,I43453,I43456,I43459,I43462,I43465,I43468,I43471,I43474,I43477,I2224,I2231);
PAT_6 I_584 (I43450,I43477,I43465,I43474,I43468,I43462,I43453,I43471,I43459,I43456,I43450,I43523,I43526,I43529,I43532,I43535,I43538,I43541,I43544,I43547,I43550,I2224,I2231);
PAT_12 I_585 (I43523,I43550,I43529,I43532,I43526,I43523,I43544,I43538,I43541,I43535,I43547,I43596,I43599,I43602,I43605,I43608,I43611,I43614,I43617,I2224,I2231);
PAT_6 I_586 (I43605,I43599,I43617,I43602,I43599,I43602,I43611,I43596,I43614,I43596,I43608,I43663,I43666,I43669,I43672,I43675,I43678,I43681,I43684,I43687,I43690,I2224,I2231);
PAT_15 I_587 (I43681,I43672,I43684,I43687,I43678,I43690,I43663,I43669,I43663,I43666,I43675,I43736,I43739,I43742,I43745,I43748,I43751,I43754,I43757,I43760,I2224,I2231);
PAT_17 I_588 (I43736,I43736,I43748,I43739,I43742,I43760,I43757,I43751,I43739,I43745,I43754,I43806,I43809,I43812,I43815,I43818,I43821,I43824,I43827,I43830,I43833,I2224,I2231);
PAT_10 I_589 (I43806,I43812,I43833,I43815,I43830,I43809,I43824,I43818,I43827,I43821,I43806,I43879,I43882,I43885,I43888,I43891,I43894,I43897,I43900,I2224,I2231);
PAT_5 I_590 (I43900,I43879,I43888,I43882,I43897,I43894,I43885,I43885,I43879,I43882,I43891,I43946,I43949,I43952,I43955,I43958,I43961,I43964,I43967,I43970,I43973,I2224,I2231);
PAT_17 I_591 (I43973,I43949,I43952,I43955,I43946,I43958,I43946,I43970,I43964,I43961,I43967,I44019,I44022,I44025,I44028,I44031,I44034,I44037,I44040,I44043,I44046,I2224,I2231);
PAT_16 I_592 (I44019,I44043,I44019,I44040,I44037,I44025,I44031,I44022,I44046,I44034,I44028,I44092,I44095,I44098,I44101,I44104,I44107,I44110,I44113,I44116,I44119,I2224,I2231);
PAT_13 I_593 (I44104,I44095,I44092,I44098,I44107,I44116,I44113,I44110,I44101,I44092,I44119,I44165,I44168,I44171,I44174,I44177,I44180,I44183,I44186,I44189,I2224,I2231);
PAT_10 I_594 (I44186,I44180,I44174,I44168,I44189,I44168,I44177,I44165,I44165,I44183,I44171,I44235,I44238,I44241,I44244,I44247,I44250,I44253,I44256,I2224,I2231);
PAT_2 I_595 (I44247,I44250,I44241,I44253,I44238,I44235,I44235,I44241,I44256,I44244,I44238,I44302,I44305,I44308,I44311,I44314,I44317,I44320,I44323,I44326,I2224,I2231);
PAT_9 I_596 (I44317,I44326,I44302,I44308,I44311,I44320,I44305,I44314,I44323,I44305,I44302,I44372,I44375,I44378,I44381,I44384,I44387,I44390,I44393,I44396,I2224,I2231);
PAT_11 I_597 (I44384,I44390,I44396,I44393,I44381,I44375,I44375,I44372,I44387,I44372,I44378,I44442,I44445,I44448,I44451,I44454,I44457,I44460,I44463,I44466,I44469,I2224,I2231);
PAT_5 I_598 (I44463,I44442,I44469,I44457,I44454,I44466,I44448,I44442,I44460,I44445,I44451,I44515,I44518,I44521,I44524,I44527,I44530,I44533,I44536,I44539,I44542,I2224,I2231);
PAT_6 I_599 (I44533,I44527,I44515,I44521,I44518,I44524,I44530,I44515,I44539,I44536,I44542,I44588,I44591,I44594,I44597,I44600,I44603,I44606,I44609,I44612,I44615,I2224,I2231);
PAT_11 I_600 (I44588,I44603,I44588,I44600,I44597,I44615,I44612,I44609,I44606,I44591,I44594,I44661,I44664,I44667,I44670,I44673,I44676,I44679,I44682,I44685,I44688,I2224,I2231);
PAT_1 I_601 (I44676,I44667,I44670,I44661,I44682,I44679,I44664,I44661,I44688,I44685,I44673,I44734,I44737,I44740,I44743,I44746,I44749,I44752,I44755,I44758,I2224,I2231);
PAT_6 I_602 (I44743,I44734,I44737,I44740,I44755,I44758,I44752,I44734,I44749,I44746,I44737,I44804,I44807,I44810,I44813,I44816,I44819,I44822,I44825,I44828,I44831,I2224,I2231);
PAT_9 I_603 (I44804,I44831,I44828,I44810,I44816,I44807,I44819,I44804,I44822,I44813,I44825,I44877,I44880,I44883,I44886,I44889,I44892,I44895,I44898,I44901,I2224,I2231);
PAT_2 I_604 (I44892,I44895,I44886,I44901,I44877,I44880,I44883,I44880,I44898,I44889,I44877,I44947,I44950,I44953,I44956,I44959,I44962,I44965,I44968,I44971,I2224,I2231);
PAT_14 I_605 (I44953,I44956,I44971,I44962,I44947,I44950,I44965,I44959,I44947,I44968,I44950,I45017,I45020,I45023,I45026,I45029,I45032,I45035,I45038,I45041,I2224,I2231);
PAT_5 I_606 (I45020,I45023,I45020,I45029,I45017,I45038,I45026,I45017,I45041,I45035,I45032,I45087,I45090,I45093,I45096,I45099,I45102,I45105,I45108,I45111,I45114,I2224,I2231);
PAT_13 I_607 (I45093,I45102,I45087,I45090,I45111,I45096,I45108,I45087,I45105,I45114,I45099,I45160,I45163,I45166,I45169,I45172,I45175,I45178,I45181,I45184,I2224,I2231);
PAT_6 I_608 (I45160,I45172,I45169,I45181,I45178,I45184,I45160,I45175,I45163,I45163,I45166,I45230,I45233,I45236,I45239,I45242,I45245,I45248,I45251,I45254,I45257,I2224,I2231);
PAT_11 I_609 (I45230,I45245,I45230,I45242,I45239,I45257,I45254,I45251,I45248,I45233,I45236,I45303,I45306,I45309,I45312,I45315,I45318,I45321,I45324,I45327,I45330,I2224,I2231);
PAT_6 I_610 (I45303,I45330,I45318,I45327,I45321,I45315,I45306,I45324,I45312,I45309,I45303,I45376,I45379,I45382,I45385,I45388,I45391,I45394,I45397,I45400,I45403,I2224,I2231);
PAT_7 I_611 (I45382,I45391,I45394,I45376,I45385,I45379,I45388,I45403,I45397,I45400,I45376,I45449,I45452,I45455,I45458,I45461,I45464,I45467,I45470,I45473,I2224,I2231);
PAT_9 I_612 (I45470,I45458,I45467,I45473,I45455,I45461,I45452,I45464,I45449,I45449,I45452,I45519,I45522,I45525,I45528,I45531,I45534,I45537,I45540,I45543,I2224,I2231);
PAT_6 I_613 (I45537,I45519,I45531,I45540,I45519,I45528,I45525,I45543,I45534,I45522,I45522,I45589,I45592,I45595,I45598,I45601,I45604,I45607,I45610,I45613,I45616,I2224,I2231);
PAT_11 I_614 (I45589,I45604,I45589,I45601,I45598,I45616,I45613,I45610,I45607,I45592,I45595,I45662,I45665,I45668,I45671,I45674,I45677,I45680,I45683,I45686,I45689,I2224,I2231);
PAT_13 I_615 (I45662,I45665,I45674,I45686,I45689,I45677,I45683,I45671,I45680,I45668,I45662,I45735,I45738,I45741,I45744,I45747,I45750,I45753,I45756,I45759,I2224,I2231);
PAT_1 I_616 (I45735,I45744,I45738,I45756,I45750,I45741,I45753,I45747,I45738,I45759,I45735,I45805,I45808,I45811,I45814,I45817,I45820,I45823,I45826,I45829,I2224,I2231);
PAT_7 I_617 (I45808,I45814,I45811,I45817,I45823,I45820,I45829,I45826,I45808,I45805,I45805,I45875,I45878,I45881,I45884,I45887,I45890,I45893,I45896,I45899,I2224,I2231);
PAT_15 I_618 (I45893,I45878,I45878,I45890,I45875,I45899,I45881,I45887,I45896,I45875,I45884,I45945,I45948,I45951,I45954,I45957,I45960,I45963,I45966,I45969,I2224,I2231);
PAT_11 I_619 (I45966,I45948,I45945,I45960,I45951,I45945,I45963,I45969,I45957,I45948,I45954,I46015,I46018,I46021,I46024,I46027,I46030,I46033,I46036,I46039,I46042,I2224,I2231);
PAT_13 I_620 (I46015,I46018,I46027,I46039,I46042,I46030,I46036,I46024,I46033,I46021,I46015,I46088,I46091,I46094,I46097,I46100,I46103,I46106,I46109,I46112,I2224,I2231);
PAT_15 I_621 (I46088,I46100,I46091,I46103,I46088,I46097,I46112,I46109,I46094,I46106,I46091,I46158,I46161,I46164,I46167,I46170,I46173,I46176,I46179,I46182,I2224,I2231);
PAT_8 I_622 (I46179,I46158,I46158,I46167,I46164,I46161,I46176,I46173,I46161,I46182,I46170,I46228,I46231,I46234,I46237,I46240,I46243,I46246,I46249,I46252,I2224,I2231);
PAT_2 I_623 (I46231,I46246,I46252,I46228,I46240,I46243,I46231,I46249,I46234,I46237,I46228,I46298,I46301,I46304,I46307,I46310,I46313,I46316,I46319,I46322,I2224,I2231);
PAT_5 I_624 (I46319,I46298,I46298,I46310,I46307,I46316,I46304,I46313,I46322,I46301,I46301,I46368,I46371,I46374,I46377,I46380,I46383,I46386,I46389,I46392,I46395,I2224,I2231);
PAT_10 I_625 (I46392,I46395,I46374,I46380,I46383,I46389,I46371,I46368,I46368,I46377,I46386,I46441,I46444,I46447,I46450,I46453,I46456,I46459,I46462,I2224,I2231);
PAT_13 I_626 (I46447,I46453,I46447,I46444,I46459,I46462,I46441,I46441,I46456,I46444,I46450,I46508,I46511,I46514,I46517,I46520,I46523,I46526,I46529,I46532,I2224,I2231);
PAT_5 I_627 (I46520,I46511,I46517,I46529,I46511,I46532,I46514,I46523,I46508,I46508,I46526,I46578,I46581,I46584,I46587,I46590,I46593,I46596,I46599,I46602,I46605,I2224,I2231);
PAT_7 I_628 (I46596,I46599,I46605,I46602,I46587,I46584,I46578,I46590,I46578,I46581,I46593,I46651,I46654,I46657,I46660,I46663,I46666,I46669,I46672,I46675,I2224,I2231);
PAT_2 I_629 (I46672,I46666,I46657,I46651,I46660,I46654,I46663,I46675,I46669,I46654,I46651,I46721,I46724,I46727,I46730,I46733,I46736,I46739,I46742,I46745,I2224,I2231);
PAT_7 I_630 (I46745,I46721,I46727,I46724,I46724,I46733,I46736,I46721,I46739,I46742,I46730,I46791,I46794,I46797,I46800,I46803,I46806,I46809,I46812,I46815,I2224,I2231);
PAT_17 I_631 (I46803,I46797,I46806,I46791,I46809,I46812,I46794,I46815,I46800,I46794,I46791,I46861,I46864,I46867,I46870,I46873,I46876,I46879,I46882,I46885,I46888,I2224,I2231);
PAT_9 I_632 (I46882,I46864,I46870,I46885,I46867,I46879,I46861,I46873,I46861,I46888,I46876,I46934,I46937,I46940,I46943,I46946,I46949,I46952,I46955,I46958,I2224,I2231);
PAT_6 I_633 (I46952,I46934,I46946,I46955,I46934,I46943,I46940,I46958,I46949,I46937,I46937,I47004,I47007,I47010,I47013,I47016,I47019,I47022,I47025,I47028,I47031,I2224,I2231);
PAT_9 I_634 (I47004,I47031,I47028,I47010,I47016,I47007,I47019,I47004,I47022,I47013,I47025,I47077,I47080,I47083,I47086,I47089,I47092,I47095,I47098,I47101,I2224,I2231);
PAT_7 I_635 (I47083,I47092,I47077,I47098,I47089,I47077,I47080,I47101,I47095,I47080,I47086,I47147,I47150,I47153,I47156,I47159,I47162,I47165,I47168,I47171,I2224,I2231);
PAT_6 I_636 (I47147,I47165,I47147,I47156,I47162,I47150,I47168,I47153,I47171,I47150,I47159,I47217,I47220,I47223,I47226,I47229,I47232,I47235,I47238,I47241,I47244,I2224,I2231);
PAT_9 I_637 (I47217,I47244,I47241,I47223,I47229,I47220,I47232,I47217,I47235,I47226,I47238,I47290,I47293,I47296,I47299,I47302,I47305,I47308,I47311,I47314,I2224,I2231);
PAT_13 I_638 (I47290,I47311,I47293,I47308,I47302,I47299,I47314,I47290,I47296,I47305,I47293,I47360,I47363,I47366,I47369,I47372,I47375,I47378,I47381,I47384,I2224,I2231);
PAT_4 I_639 (I47369,I47372,I47384,I47366,I47381,I47378,I47363,I47375,I47363,I47360,I47360,I47430,I47433,I47436,I47439,I47442,I47445,I47448,I47451,I47454,I2224,I2231);
PAT_9 I_640 (I47451,I47433,I47436,I47445,I47448,I47430,I47439,I47433,I47454,I47430,I47442,I47500,I47503,I47506,I47509,I47512,I47515,I47518,I47521,I47524,I2224,I2231);
PAT_4 I_641 (I47500,I47524,I47518,I47506,I47503,I47521,I47503,I47500,I47515,I47509,I47512,I47570,I47573,I47576,I47579,I47582,I47585,I47588,I47591,I47594,I2224,I2231);
PAT_17 I_642 (I47582,I47579,I47591,I47585,I47570,I47588,I47594,I47573,I47576,I47573,I47570,I47640,I47643,I47646,I47649,I47652,I47655,I47658,I47661,I47664,I47667,I2224,I2231);
PAT_5 I_643 (I47652,I47646,I47643,I47664,I47649,I47655,I47658,I47640,I47640,I47661,I47667,I47713,I47716,I47719,I47722,I47725,I47728,I47731,I47734,I47737,I47740,I2224,I2231);
PAT_6 I_644 (I47731,I47725,I47713,I47719,I47716,I47722,I47728,I47713,I47737,I47734,I47740,I47786,I47789,I47792,I47795,I47798,I47801,I47804,I47807,I47810,I47813,I2224,I2231);
PAT_13 I_645 (I47810,I47792,I47807,I47786,I47789,I47795,I47813,I47798,I47804,I47786,I47801,I47859,I47862,I47865,I47868,I47871,I47874,I47877,I47880,I47883,I2224,I2231);
PAT_10 I_646 (I47880,I47874,I47868,I47862,I47883,I47862,I47871,I47859,I47859,I47877,I47865,I47929,I47932,I47935,I47938,I47941,I47944,I47947,I47950,I2224,I2231);
PAT_6 I_647 (I47950,I47944,I47938,I47932,I47929,I47935,I47929,I47935,I47932,I47941,I47947,I47996,I47999,I48002,I48005,I48008,I48011,I48014,I48017,I48020,I48023,I2224,I2231);
PAT_12 I_648 (I47996,I48023,I48002,I48005,I47999,I47996,I48017,I48011,I48014,I48008,I48020,I48069,I48072,I48075,I48078,I48081,I48084,I48087,I48090,I2224,I2231);
PAT_13 I_649 (I48081,I48084,I48075,I48090,I48087,I48069,I48072,I48078,I48075,I48072,I48069,I48136,I48139,I48142,I48145,I48148,I48151,I48154,I48157,I48160,I2224,I2231);
PAT_1 I_650 (I48136,I48145,I48139,I48157,I48151,I48142,I48154,I48148,I48139,I48160,I48136,I48206,I48209,I48212,I48215,I48218,I48221,I48224,I48227,I48230,I2224,I2231);
PAT_9 I_651 (I48221,I48227,I48212,I48230,I48209,I48224,I48209,I48215,I48206,I48218,I48206,I48276,I48279,I48282,I48285,I48288,I48291,I48294,I48297,I48300,I2224,I2231);
PAT_7 I_652 (I48282,I48291,I48276,I48297,I48288,I48276,I48279,I48300,I48294,I48279,I48285,I48346,I48349,I48352,I48355,I48358,I48361,I48364,I48367,I48370,I2224,I2231);
PAT_4 I_653 (I48370,I48346,I48346,I48361,I48355,I48349,I48349,I48364,I48367,I48352,I48358,I48416,I48419,I48422,I48425,I48428,I48431,I48434,I48437,I48440,I2224,I2231);
PAT_5 I_654 (I48437,I48419,I48419,I48431,I48434,I48428,I48425,I48416,I48422,I48416,I48440,I48486,I48489,I48492,I48495,I48498,I48501,I48504,I48507,I48510,I48513,I2224,I2231);
PAT_14 I_655 (I48507,I48492,I48486,I48510,I48513,I48486,I48504,I48489,I48495,I48498,I48501,I48559,I48562,I48565,I48568,I48571,I48574,I48577,I48580,I48583,I2224,I2231);
PAT_11 I_656 (I48571,I48568,I48565,I48559,I48562,I48562,I48574,I48559,I48580,I48583,I48577,I48629,I48632,I48635,I48638,I48641,I48644,I48647,I48650,I48653,I48656,I2224,I2231);
PAT_13 I_657 (I48629,I48632,I48641,I48653,I48656,I48644,I48650,I48638,I48647,I48635,I48629,I48702,I48705,I48708,I48711,I48714,I48717,I48720,I48723,I48726,I2224,I2231);
PAT_6 I_658 (I48702,I48714,I48711,I48723,I48720,I48726,I48702,I48717,I48705,I48705,I48708,I48772,I48775,I48778,I48781,I48784,I48787,I48790,I48793,I48796,I48799,I2224,I2231);
PAT_11 I_659 (I48772,I48787,I48772,I48784,I48781,I48799,I48796,I48793,I48790,I48775,I48778,I48845,I48848,I48851,I48854,I48857,I48860,I48863,I48866,I48869,I48872,I2224,I2231);
PAT_2 I_660 (I48845,I48869,I48857,I48851,I48860,I48863,I48848,I48872,I48866,I48854,I48845,I48918,I48921,I48924,I48927,I48930,I48933,I48936,I48939,I48942,I2224,I2231);
PAT_6 I_661 (I48942,I48918,I48933,I48930,I48936,I48927,I48921,I48939,I48918,I48924,I48921,I48988,I48991,I48994,I48997,I49000,I49003,I49006,I49009,I49012,I49015,I2224,I2231);
PAT_4 I_662 (I48988,I49003,I48991,I48994,I48997,I48988,I49015,I49006,I49009,I49000,I49012,I49061,I49064,I49067,I49070,I49073,I49076,I49079,I49082,I49085,I2224,I2231);
PAT_5 I_663 (I49082,I49064,I49064,I49076,I49079,I49073,I49070,I49061,I49067,I49061,I49085,I49131,I49134,I49137,I49140,I49143,I49146,I49149,I49152,I49155,I49158,I2224,I2231);
PAT_8 I_664 (I49131,I49158,I49149,I49146,I49140,I49131,I49143,I49155,I49134,I49152,I49137,I49204,I49207,I49210,I49213,I49216,I49219,I49222,I49225,I49228,I2224,I2231);
PAT_17 I_665 (I49228,I49216,I49213,I49207,I49210,I49222,I49204,I49207,I49204,I49219,I49225,I49274,I49277,I49280,I49283,I49286,I49289,I49292,I49295,I49298,I49301,I2224,I2231);
PAT_11 I_666 (I49286,I49295,I49301,I49277,I49274,I49292,I49283,I49289,I49280,I49298,I49274,I49347,I49350,I49353,I49356,I49359,I49362,I49365,I49368,I49371,I49374,I2224,I2231);
PAT_12 I_667 (I49356,I49371,I49353,I49350,I49359,I49362,I49368,I49347,I49365,I49374,I49347,I49420,I49423,I49426,I49429,I49432,I49435,I49438,I49441,I2224,I2231);
PAT_5 I_668 (I49429,I49435,I49441,I49426,I49426,I49420,I49438,I49420,I49423,I49423,I49432,I49487,I49490,I49493,I49496,I49499,I49502,I49505,I49508,I49511,I49514,I2224,I2231);
PAT_2 I_669 (I49502,I49487,I49499,I49493,I49508,I49490,I49505,I49496,I49511,I49514,I49487,I49560,I49563,I49566,I49569,I49572,I49575,I49578,I49581,I49584,I2224,I2231);
PAT_6 I_670 (I49584,I49560,I49575,I49572,I49578,I49569,I49563,I49581,I49560,I49566,I49563,I49630,I49633,I49636,I49639,I49642,I49645,I49648,I49651,I49654,I49657,I2224,I2231);
PAT_9 I_671 (I49630,I49657,I49654,I49636,I49642,I49633,I49645,I49630,I49648,I49639,I49651,I49703,I49706,I49709,I49712,I49715,I49718,I49721,I49724,I49727,I2224,I2231);
PAT_14 I_672 (I49712,I49703,I49727,I49709,I49706,I49703,I49718,I49724,I49715,I49706,I49721,I49773,I49776,I49779,I49782,I49785,I49788,I49791,I49794,I49797,I2224,I2231);
PAT_9 I_673 (I49782,I49794,I49773,I49791,I49776,I49779,I49797,I49776,I49785,I49773,I49788,I49843,I49846,I49849,I49852,I49855,I49858,I49861,I49864,I49867,I2224,I2231);
PAT_8 I_674 (I49864,I49852,I49861,I49843,I49846,I49858,I49867,I49846,I49849,I49855,I49843,I49913,I49916,I49919,I49922,I49925,I49928,I49931,I49934,I49937,I2224,I2231);
PAT_10 I_675 (I49919,I49913,I49916,I49937,I49931,I49916,I49925,I49913,I49934,I49928,I49922,I49983,I49986,I49989,I49992,I49995,I49998,I50001,I50004,I2224,I2231);
PAT_5 I_676 (I50004,I49983,I49992,I49986,I50001,I49998,I49989,I49989,I49983,I49986,I49995,I50050,I50053,I50056,I50059,I50062,I50065,I50068,I50071,I50074,I50077,I2224,I2231);
PAT_4 I_677 (I50068,I50074,I50077,I50056,I50059,I50071,I50053,I50050,I50062,I50065,I50050,I50123,I50126,I50129,I50132,I50135,I50138,I50141,I50144,I50147,I2224,I2231);
PAT_13 I_678 (I50138,I50132,I50144,I50129,I50135,I50123,I50147,I50141,I50126,I50123,I50126,I50193,I50196,I50199,I50202,I50205,I50208,I50211,I50214,I50217,I2224,I2231);
PAT_11 I_679 (I50193,I50205,I50208,I50199,I50196,I50217,I50196,I50214,I50202,I50193,I50211,I50263,I50266,I50269,I50272,I50275,I50278,I50281,I50284,I50287,I50290,I2224,I2231);
PAT_4 I_680 (I50269,I50290,I50263,I50281,I50272,I50263,I50284,I50266,I50275,I50287,I50278,I50336,I50339,I50342,I50345,I50348,I50351,I50354,I50357,I50360,I2224,I2231);
PAT_17 I_681 (I50348,I50345,I50357,I50351,I50336,I50354,I50360,I50339,I50342,I50339,I50336,I50406,I50409,I50412,I50415,I50418,I50421,I50424,I50427,I50430,I50433,I2224,I2231);
PAT_9 I_682 (I50427,I50409,I50415,I50430,I50412,I50424,I50406,I50418,I50406,I50433,I50421,I50479,I50482,I50485,I50488,I50491,I50494,I50497,I50500,I50503,I2224,I2231);
PAT_7 I_683 (I50485,I50494,I50479,I50500,I50491,I50479,I50482,I50503,I50497,I50482,I50488,I50549,I50552,I50555,I50558,I50561,I50564,I50567,I50570,I50573,I2224,I2231);
PAT_13 I_684 (I50555,I50573,I50564,I50549,I50561,I50549,I50570,I50552,I50558,I50552,I50567,I50619,I50622,I50625,I50628,I50631,I50634,I50637,I50640,I50643,I2224,I2231);
PAT_1 I_685 (I50619,I50628,I50622,I50640,I50634,I50625,I50637,I50631,I50622,I50643,I50619,I50689,I50692,I50695,I50698,I50701,I50704,I50707,I50710,I50713,I2224,I2231);
PAT_17 I_686 (I50701,I50689,I50710,I50713,I50692,I50695,I50692,I50704,I50698,I50689,I50707,I50759,I50762,I50765,I50768,I50771,I50774,I50777,I50780,I50783,I50786,I2224,I2231);
PAT_9 I_687 (I50780,I50762,I50768,I50783,I50765,I50777,I50759,I50771,I50759,I50786,I50774,I50832,I50835,I50838,I50841,I50844,I50847,I50850,I50853,I50856,I2224,I2231);
PAT_7 I_688 (I50838,I50847,I50832,I50853,I50844,I50832,I50835,I50856,I50850,I50835,I50841,I50902,I50905,I50908,I50911,I50914,I50917,I50920,I50923,I50926,I2224,I2231);
PAT_11 I_689 (I50914,I50908,I50902,I50923,I50926,I50911,I50905,I50920,I50902,I50917,I50905,I50972,I50975,I50978,I50981,I50984,I50987,I50990,I50993,I50996,I50999,I2224,I2231);
PAT_1 I_690 (I50987,I50978,I50981,I50972,I50993,I50990,I50975,I50972,I50999,I50996,I50984,I51045,I51048,I51051,I51054,I51057,I51060,I51063,I51066,I51069,I2224,I2231);
PAT_13 I_691 (I51054,I51063,I51069,I51045,I51060,I51057,I51066,I51051,I51048,I51045,I51048,I51115,I51118,I51121,I51124,I51127,I51130,I51133,I51136,I51139,I2224,I2231);
PAT_9 I_692 (I51136,I51118,I51118,I51115,I51139,I51121,I51124,I51115,I51127,I51133,I51130,I51185,I51188,I51191,I51194,I51197,I51200,I51203,I51206,I51209,I2224,I2231);
PAT_8 I_693 (I51206,I51194,I51203,I51185,I51188,I51200,I51209,I51188,I51191,I51197,I51185,I51255,I51258,I51261,I51264,I51267,I51270,I51273,I51276,I51279,I2224,I2231);
PAT_10 I_694 (I51261,I51255,I51258,I51279,I51273,I51258,I51267,I51255,I51276,I51270,I51264,I51325,I51328,I51331,I51334,I51337,I51340,I51343,I51346,I2224,I2231);
PAT_1 I_695 (I51331,I51331,I51340,I51325,I51337,I51328,I51343,I51325,I51346,I51334,I51328,I51392,I51395,I51398,I51401,I51404,I51407,I51410,I51413,I51416,I2224,I2231);
PAT_15 I_696 (I51395,I51404,I51392,I51407,I51401,I51395,I51416,I51413,I51410,I51398,I51392,I51462,I51465,I51468,I51471,I51474,I51477,I51480,I51483,I51486,I2224,I2231);
PAT_6 I_697 (I51465,I51462,I51468,I51483,I51465,I51486,I51471,I51477,I51474,I51480,I51462,I51532,I51535,I51538,I51541,I51544,I51547,I51550,I51553,I51556,I51559,I2224,I2231);
PAT_17 I_698 (I51544,I51547,I51553,I51541,I51535,I51556,I51550,I51532,I51559,I51538,I51532,I51605,I51608,I51611,I51614,I51617,I51620,I51623,I51626,I51629,I51632,I2224,I2231);
PAT_13 I_699 (I51623,I51626,I51611,I51605,I51617,I51629,I51608,I51620,I51605,I51632,I51614,I51678,I51681,I51684,I51687,I51690,I51693,I51696,I51699,I51702,I2224,I2231);
PAT_14 I_700 (I51681,I51696,I51684,I51693,I51687,I51678,I51690,I51699,I51678,I51702,I51681,I51748,I51751,I51754,I51757,I51760,I51763,I51766,I51769,I51772,I2224,I2231);
PAT_16 I_701 (I51763,I51769,I51766,I51772,I51754,I51748,I51757,I51751,I51751,I51760,I51748,I51818,I51821,I51824,I51827,I51830,I51833,I51836,I51839,I51842,I51845,I2224,I2231);
PAT_8 I_702 (I51818,I51821,I51830,I51839,I51827,I51842,I51845,I51833,I51824,I51836,I51818,I51891,I51894,I51897,I51900,I51903,I51906,I51909,I51912,I51915,I2224,I2231);
PAT_5 I_703 (I51897,I51915,I51891,I51912,I51900,I51903,I51894,I51891,I51894,I51906,I51909,I51961,I51964,I51967,I51970,I51973,I51976,I51979,I51982,I51985,I51988,I2224,I2231);
PAT_1 I_704 (I51976,I51964,I51982,I51961,I51967,I51961,I51970,I51985,I51979,I51988,I51973,I52034,I52037,I52040,I52043,I52046,I52049,I52052,I52055,I52058,I2224,I2231);
PAT_9 I_705 (I52049,I52055,I52040,I52058,I52037,I52052,I52037,I52043,I52034,I52046,I52034,I52104,I52107,I52110,I52113,I52116,I52119,I52122,I52125,I52128,I2224,I2231);
PAT_4 I_706 (I52104,I52128,I52122,I52110,I52107,I52125,I52107,I52104,I52119,I52113,I52116,I52174,I52177,I52180,I52183,I52186,I52189,I52192,I52195,I52198,I2224,I2231);
PAT_6 I_707 (I52174,I52180,I52177,I52189,I52192,I52186,I52198,I52195,I52174,I52183,I52177,I52244,I52247,I52250,I52253,I52256,I52259,I52262,I52265,I52268,I52271,I2224,I2231);
PAT_11 I_708 (I52244,I52259,I52244,I52256,I52253,I52271,I52268,I52265,I52262,I52247,I52250,I52317,I52320,I52323,I52326,I52329,I52332,I52335,I52338,I52341,I52344,I2224,I2231);
PAT_8 I_709 (I52326,I52332,I52335,I52341,I52338,I52329,I52317,I52317,I52344,I52320,I52323,I52390,I52393,I52396,I52399,I52402,I52405,I52408,I52411,I52414,I2224,I2231);
PAT_1 I_710 (I52393,I52414,I52396,I52411,I52393,I52399,I52390,I52390,I52408,I52405,I52402,I52460,I52463,I52466,I52469,I52472,I52475,I52478,I52481,I52484,I2224,I2231);
PAT_14 I_711 (I52463,I52478,I52475,I52466,I52460,I52460,I52472,I52481,I52484,I52469,I52463,I52530,I52533,I52536,I52539,I52542,I52545,I52548,I52551,I52554,I2224,I2231);
PAT_9 I_712 (I52539,I52551,I52530,I52548,I52533,I52536,I52554,I52533,I52542,I52530,I52545,I52600,I52603,I52606,I52609,I52612,I52615,I52618,I52621,I52624,I2224,I2231);
PAT_13 I_713 (I52600,I52621,I52603,I52618,I52612,I52609,I52624,I52600,I52606,I52615,I52603,I52670,I52673,I52676,I52679,I52682,I52685,I52688,I52691,I52694,I2224,I2231);
PAT_4 I_714 (I52679,I52682,I52694,I52676,I52691,I52688,I52673,I52685,I52673,I52670,I52670,I52740,I52743,I52746,I52749,I52752,I52755,I52758,I52761,I52764,I2224,I2231);
PAT_10 I_715 (I52740,I52740,I52764,I52743,I52749,I52758,I52755,I52743,I52761,I52746,I52752,I52810,I52813,I52816,I52819,I52822,I52825,I52828,I52831,I2224,I2231);
PAT_11 I_716 (I52819,I52822,I52831,I52825,I52828,I52810,I52810,I52816,I52813,I52813,I52816,I52877,I52880,I52883,I52886,I52889,I52892,I52895,I52898,I52901,I52904,I2224,I2231);
PAT_9 I_717 (I52883,I52895,I52886,I52898,I52877,I52880,I52889,I52877,I52892,I52901,I52904,I52950,I52953,I52956,I52959,I52962,I52965,I52968,I52971,I52974,I2224,I2231);
PAT_4 I_718 (I52950,I52974,I52968,I52956,I52953,I52971,I52953,I52950,I52965,I52959,I52962,I53020,I53023,I53026,I53029,I53032,I53035,I53038,I53041,I53044,I2224,I2231);
PAT_7 I_719 (I53035,I53029,I53026,I53020,I53032,I53038,I53023,I53023,I53041,I53044,I53020,I53090,I53093,I53096,I53099,I53102,I53105,I53108,I53111,I53114,I2224,I2231);
PAT_17 I_720 (I53102,I53096,I53105,I53090,I53108,I53111,I53093,I53114,I53099,I53093,I53090,I53160,I53163,I53166,I53169,I53172,I53175,I53178,I53181,I53184,I53187,I2224,I2231);
PAT_5 I_721 (I53172,I53166,I53163,I53184,I53169,I53175,I53178,I53160,I53160,I53181,I53187,I53233,I53236,I53239,I53242,I53245,I53248,I53251,I53254,I53257,I53260,I2224,I2231);
PAT_13 I_722 (I53239,I53248,I53233,I53236,I53257,I53242,I53254,I53233,I53251,I53260,I53245,I53306,I53309,I53312,I53315,I53318,I53321,I53324,I53327,I53330,I2224,I2231);
PAT_4 I_723 (I53315,I53318,I53330,I53312,I53327,I53324,I53309,I53321,I53309,I53306,I53306,I53376,I53379,I53382,I53385,I53388,I53391,I53394,I53397,I53400,I2224,I2231);
PAT_17 I_724 (I53388,I53385,I53397,I53391,I53376,I53394,I53400,I53379,I53382,I53379,I53376,I53446,I53449,I53452,I53455,I53458,I53461,I53464,I53467,I53470,I53473,I2224,I2231);
PAT_13 I_725 (I53464,I53467,I53452,I53446,I53458,I53470,I53449,I53461,I53446,I53473,I53455,I53519,I53522,I53525,I53528,I53531,I53534,I53537,I53540,I53543,I2224,I2231);
PAT_9 I_726 (I53540,I53522,I53522,I53519,I53543,I53525,I53528,I53519,I53531,I53537,I53534,I53589,I53592,I53595,I53598,I53601,I53604,I53607,I53610,I53613,I2224,I2231);
PAT_2 I_727 (I53604,I53607,I53598,I53613,I53589,I53592,I53595,I53592,I53610,I53601,I53589,I53659,I53662,I53665,I53668,I53671,I53674,I53677,I53680,I53683,I2224,I2231);
PAT_4 I_728 (I53659,I53665,I53683,I53677,I53674,I53671,I53662,I53680,I53659,I53662,I53668,I53729,I53732,I53735,I53738,I53741,I53744,I53747,I53750,I53753,I2224,I2231);
PAT_13 I_729 (I53744,I53738,I53750,I53735,I53741,I53729,I53753,I53747,I53732,I53729,I53732,I53799,I53802,I53805,I53808,I53811,I53814,I53817,I53820,I53823,I2224,I2231);
PAT_2 I_730 (I53817,I53811,I53808,I53814,I53799,I53823,I53802,I53820,I53799,I53805,I53802,I53869,I53872,I53875,I53878,I53881,I53884,I53887,I53890,I53893,I2224,I2231);
PAT_10 I_731 (I53869,I53887,I53884,I53872,I53875,I53890,I53881,I53869,I53878,I53893,I53872,I53939,I53942,I53945,I53948,I53951,I53954,I53957,I53960,I2224,I2231);
PAT_5 I_732 (I53960,I53939,I53948,I53942,I53957,I53954,I53945,I53945,I53939,I53942,I53951,I54006,I54009,I54012,I54015,I54018,I54021,I54024,I54027,I54030,I54033,I2224,I2231);
PAT_10 I_733 (I54030,I54033,I54012,I54018,I54021,I54027,I54009,I54006,I54006,I54015,I54024,I54079,I54082,I54085,I54088,I54091,I54094,I54097,I54100,I2224,I2231);
PAT_13 I_734 (I54085,I54091,I54085,I54082,I54097,I54100,I54079,I54079,I54094,I54082,I54088,I54146,I54149,I54152,I54155,I54158,I54161,I54164,I54167,I54170,I2224,I2231);
PAT_9 I_735 (I54167,I54149,I54149,I54146,I54170,I54152,I54155,I54146,I54158,I54164,I54161,I54216,I54219,I54222,I54225,I54228,I54231,I54234,I54237,I54240,I2224,I2231);
PAT_17 I_736 (I54219,I54225,I54240,I54231,I54234,I54222,I54216,I54228,I54216,I54219,I54237,I54286,I54289,I54292,I54295,I54298,I54301,I54304,I54307,I54310,I54313,I2224,I2231);
PAT_11 I_737 (I54298,I54307,I54313,I54289,I54286,I54304,I54295,I54301,I54292,I54310,I54286,I54359,I54362,I54365,I54368,I54371,I54374,I54377,I54380,I54383,I54386,I2224,I2231);
PAT_12 I_738 (I54368,I54383,I54365,I54362,I54371,I54374,I54380,I54359,I54377,I54386,I54359,I54432,I54435,I54438,I54441,I54444,I54447,I54450,I54453,I2224,I2231);
PAT_13 I_739 (I54444,I54447,I54438,I54453,I54450,I54432,I54435,I54441,I54438,I54435,I54432,I54499,I54502,I54505,I54508,I54511,I54514,I54517,I54520,I54523,I2224,I2231);
PAT_9 I_740 (I54520,I54502,I54502,I54499,I54523,I54505,I54508,I54499,I54511,I54517,I54514,I54569,I54572,I54575,I54578,I54581,I54584,I54587,I54590,I54593,I2224,I2231);
PAT_13 I_741 (I54569,I54590,I54572,I54587,I54581,I54578,I54593,I54569,I54575,I54584,I54572,I54639,I54642,I54645,I54648,I54651,I54654,I54657,I54660,I54663,I2224,I2231);
PAT_11 I_742 (I54639,I54651,I54654,I54645,I54642,I54663,I54642,I54660,I54648,I54639,I54657,I54709,I54712,I54715,I54718,I54721,I54724,I54727,I54730,I54733,I54736,I2224,I2231);
PAT_17 I_743 (I54721,I54712,I54736,I54709,I54718,I54730,I54727,I54724,I54709,I54733,I54715,I54782,I54785,I54788,I54791,I54794,I54797,I54800,I54803,I54806,I54809,I2224,I2231);
PAT_9 I_744 (I54803,I54785,I54791,I54806,I54788,I54800,I54782,I54794,I54782,I54809,I54797,I54855,I54858,I54861,I54864,I54867,I54870,I54873,I54876,I54879,I2224,I2231);
PAT_5 I_745 (I54876,I54855,I54870,I54855,I54861,I54864,I54858,I54858,I54873,I54867,I54879,I54925,I54928,I54931,I54934,I54937,I54940,I54943,I54946,I54949,I54952,I2224,I2231);
PAT_4 I_746 (I54943,I54949,I54952,I54931,I54934,I54946,I54928,I54925,I54937,I54940,I54925,I54998,I55001,I55004,I55007,I55010,I55013,I55016,I55019,I55022,I2224,I2231);
PAT_9 I_747 (I55019,I55001,I55004,I55013,I55016,I54998,I55007,I55001,I55022,I54998,I55010,I55068,I55071,I55074,I55077,I55080,I55083,I55086,I55089,I55092,I2224,I2231);
PAT_2 I_748 (I55083,I55086,I55077,I55092,I55068,I55071,I55074,I55071,I55089,I55080,I55068,I55138,I55141,I55144,I55147,I55150,I55153,I55156,I55159,I55162,I2224,I2231);
PAT_11 I_749 (I55141,I55153,I55138,I55150,I55147,I55159,I55156,I55141,I55162,I55144,I55138,I55208,I55211,I55214,I55217,I55220,I55223,I55226,I55229,I55232,I55235,I2224,I2231);
PAT_9 I_750 (I55214,I55226,I55217,I55229,I55208,I55211,I55220,I55208,I55223,I55232,I55235,I55281,I55284,I55287,I55290,I55293,I55296,I55299,I55302,I55305,I2224,I2231);
PAT_14 I_751 (I55290,I55281,I55305,I55287,I55284,I55281,I55296,I55302,I55293,I55284,I55299,I55351,I55354,I55357,I55360,I55363,I55366,I55369,I55372,I55375,I2224,I2231);
PAT_5 I_752 (I55354,I55357,I55354,I55363,I55351,I55372,I55360,I55351,I55375,I55369,I55366,I55421,I55424,I55427,I55430,I55433,I55436,I55439,I55442,I55445,I55448,I2224,I2231);
PAT_12 I_753 (I55448,I55436,I55421,I55445,I55424,I55421,I55427,I55430,I55433,I55439,I55442,I55494,I55497,I55500,I55503,I55506,I55509,I55512,I55515,I2224,I2231);
PAT_10 I_754 (I55494,I55515,I55506,I55509,I55500,I55497,I55494,I55512,I55500,I55503,I55497,I55561,I55564,I55567,I55570,I55573,I55576,I55579,I55582,I2224,I2231);
PAT_5 I_755 (I55582,I55561,I55570,I55564,I55579,I55576,I55567,I55567,I55561,I55564,I55573,I55628,I55631,I55634,I55637,I55640,I55643,I55646,I55649,I55652,I55655,I2224,I2231);
PAT_7 I_756 (I55646,I55649,I55655,I55652,I55637,I55634,I55628,I55640,I55628,I55631,I55643,I55701,I55704,I55707,I55710,I55713,I55716,I55719,I55722,I55725,I2224,I2231);
PAT_6 I_757 (I55701,I55719,I55701,I55710,I55716,I55704,I55722,I55707,I55725,I55704,I55713,I55771,I55774,I55777,I55780,I55783,I55786,I55789,I55792,I55795,I55798,I2224,I2231);
PAT_13 I_758 (I55795,I55777,I55792,I55771,I55774,I55780,I55798,I55783,I55789,I55771,I55786,I55844,I55847,I55850,I55853,I55856,I55859,I55862,I55865,I55868,I2224,I2231);
PAT_1 I_759 (I55844,I55853,I55847,I55865,I55859,I55850,I55862,I55856,I55847,I55868,I55844,I55914,I55917,I55920,I55923,I55926,I55929,I55932,I55935,I55938,I2224,I2231);
PAT_17 I_760 (I55926,I55914,I55935,I55938,I55917,I55920,I55917,I55929,I55923,I55914,I55932,I55984,I55987,I55990,I55993,I55996,I55999,I56002,I56005,I56008,I56011,I2224,I2231);
PAT_4 I_761 (I55993,I55984,I56002,I55999,I56011,I56008,I55987,I55984,I55990,I55996,I56005,I56057,I56060,I56063,I56066,I56069,I56072,I56075,I56078,I56081,I2224,I2231);
PAT_11 I_762 (I56069,I56078,I56060,I56072,I56057,I56060,I56057,I56066,I56081,I56075,I56063,I56127,I56130,I56133,I56136,I56139,I56142,I56145,I56148,I56151,I56154,I2224,I2231);
PAT_4 I_763 (I56133,I56154,I56127,I56145,I56136,I56127,I56148,I56130,I56139,I56151,I56142,I56200,I56203,I56206,I56209,I56212,I56215,I56218,I56221,I56224,I2224,I2231);
PAT_17 I_764 (I56212,I56209,I56221,I56215,I56200,I56218,I56224,I56203,I56206,I56203,I56200,I56270,I56273,I56276,I56279,I56282,I56285,I56288,I56291,I56294,I56297,I2224,I2231);
PAT_6 I_765 (I56270,I56288,I56276,I56279,I56285,I56270,I56282,I56273,I56294,I56297,I56291,I56343,I56346,I56349,I56352,I56355,I56358,I56361,I56364,I56367,I56370,I2224,I2231);
PAT_13 I_766 (I56367,I56349,I56364,I56343,I56346,I56352,I56370,I56355,I56361,I56343,I56358,I56416,I56419,I56422,I56425,I56428,I56431,I56434,I56437,I56440,I2224,I2231);
PAT_15 I_767 (I56416,I56428,I56419,I56431,I56416,I56425,I56440,I56437,I56422,I56434,I56419,I56486,I56489,I56492,I56495,I56498,I56501,I56504,I56507,I56510,I2224,I2231);
PAT_2 I_768 (I56489,I56489,I56492,I56498,I56486,I56486,I56495,I56510,I56504,I56507,I56501,I56556,I56559,I56562,I56565,I56568,I56571,I56574,I56577,I56580,I2224,I2231);
PAT_16 I_769 (I56574,I56556,I56577,I56565,I56556,I56568,I56562,I56559,I56559,I56580,I56571,I56626,I56629,I56632,I56635,I56638,I56641,I56644,I56647,I56650,I56653,I2224,I2231);
PAT_5 I_770 (I56644,I56647,I56635,I56641,I56632,I56626,I56650,I56653,I56629,I56626,I56638,I56699,I56702,I56705,I56708,I56711,I56714,I56717,I56720,I56723,I56726,I2224,I2231);
PAT_13 I_771 (I56705,I56714,I56699,I56702,I56723,I56708,I56720,I56699,I56717,I56726,I56711,I56772,I56775,I56778,I56781,I56784,I56787,I56790,I56793,I56796,I2224,I2231);
PAT_6 I_772 (I56772,I56784,I56781,I56793,I56790,I56796,I56772,I56787,I56775,I56775,I56778,I56842,I56845,I56848,I56851,I56854,I56857,I56860,I56863,I56866,I56869,I2224,I2231);
PAT_10 I_773 (I56842,I56857,I56860,I56851,I56842,I56866,I56869,I56845,I56854,I56848,I56863,I56915,I56918,I56921,I56924,I56927,I56930,I56933,I56936,I2224,I2231);
PAT_8 I_774 (I56936,I56927,I56918,I56915,I56924,I56915,I56930,I56918,I56933,I56921,I56921,I56982,I56985,I56988,I56991,I56994,I56997,I57000,I57003,I57006,I2224,I2231);
PAT_9 I_775 (I56985,I56994,I56985,I56982,I56997,I56988,I57003,I56991,I57000,I56982,I57006,I57052,I57055,I57058,I57061,I57064,I57067,I57070,I57073,I57076,I2224,I2231);
PAT_4 I_776 (I57052,I57076,I57070,I57058,I57055,I57073,I57055,I57052,I57067,I57061,I57064,I57122,I57125,I57128,I57131,I57134,I57137,I57140,I57143,I57146,I2224,I2231);
PAT_6 I_777 (I57122,I57128,I57125,I57137,I57140,I57134,I57146,I57143,I57122,I57131,I57125,I57192,I57195,I57198,I57201,I57204,I57207,I57210,I57213,I57216,I57219,I2224,I2231);
PAT_17 I_778 (I57204,I57207,I57213,I57201,I57195,I57216,I57210,I57192,I57219,I57198,I57192,I57265,I57268,I57271,I57274,I57277,I57280,I57283,I57286,I57289,I57292,I2224,I2231);
PAT_13 I_779 (I57283,I57286,I57271,I57265,I57277,I57289,I57268,I57280,I57265,I57292,I57274,I57338,I57341,I57344,I57347,I57350,I57353,I57356,I57359,I57362,I2224,I2231);
PAT_1 I_780 (I57338,I57347,I57341,I57359,I57353,I57344,I57356,I57350,I57341,I57362,I57338,I57408,I57411,I57414,I57417,I57420,I57423,I57426,I57429,I57432,I2224,I2231);
PAT_11 I_781 (I57411,I57426,I57423,I57429,I57432,I57411,I57417,I57420,I57408,I57414,I57408,I57478,I57481,I57484,I57487,I57490,I57493,I57496,I57499,I57502,I57505,I2224,I2231);
PAT_5 I_782 (I57499,I57478,I57505,I57493,I57490,I57502,I57484,I57478,I57496,I57481,I57487,I57551,I57554,I57557,I57560,I57563,I57566,I57569,I57572,I57575,I57578,I2224,I2231);
PAT_13 I_783 (I57557,I57566,I57551,I57554,I57575,I57560,I57572,I57551,I57569,I57578,I57563,I57624,I57627,I57630,I57633,I57636,I57639,I57642,I57645,I57648,I2224,I2231);
PAT_4 I_784 (I57633,I57636,I57648,I57630,I57645,I57642,I57627,I57639,I57627,I57624,I57624,I57694,I57697,I57700,I57703,I57706,I57709,I57712,I57715,I57718,I2224,I2231);
PAT_11 I_785 (I57706,I57715,I57697,I57709,I57694,I57697,I57694,I57703,I57718,I57712,I57700,I57764,I57767,I57770,I57773,I57776,I57779,I57782,I57785,I57788,I57791,I2224,I2231);
PAT_5 I_786 (I57785,I57764,I57791,I57779,I57776,I57788,I57770,I57764,I57782,I57767,I57773,I57837,I57840,I57843,I57846,I57849,I57852,I57855,I57858,I57861,I57864,I2224,I2231);
PAT_1 I_787 (I57852,I57840,I57858,I57837,I57843,I57837,I57846,I57861,I57855,I57864,I57849,I57910,I57913,I57916,I57919,I57922,I57925,I57928,I57931,I57934,I2224,I2231);
PAT_9 I_788 (I57925,I57931,I57916,I57934,I57913,I57928,I57913,I57919,I57910,I57922,I57910,I57980,I57983,I57986,I57989,I57992,I57995,I57998,I58001,I58004,I2224,I2231);
PAT_5 I_789 (I58001,I57980,I57995,I57980,I57986,I57989,I57983,I57983,I57998,I57992,I58004,I58050,I58053,I58056,I58059,I58062,I58065,I58068,I58071,I58074,I58077,I2224,I2231);
PAT_7 I_790 (I58068,I58071,I58077,I58074,I58059,I58056,I58050,I58062,I58050,I58053,I58065,I58123,I58126,I58129,I58132,I58135,I58138,I58141,I58144,I58147,I2224,I2231);
PAT_14 I_791 (I58138,I58132,I58123,I58126,I58135,I58141,I58129,I58144,I58126,I58123,I58147,I58193,I58196,I58199,I58202,I58205,I58208,I58211,I58214,I58217,I2224,I2231);
PAT_10 I_792 (I58196,I58193,I58199,I58217,I58214,I58208,I58196,I58211,I58193,I58205,I58202,I58263,I58266,I58269,I58272,I58275,I58278,I58281,I58284,I2224,I2231);
PAT_5 I_793 (I58284,I58263,I58272,I58266,I58281,I58278,I58269,I58269,I58263,I58266,I58275,I58330,I58333,I58336,I58339,I58342,I58345,I58348,I58351,I58354,I58357,I2224,I2231);
PAT_15 I_794 (I58348,I58333,I58330,I58330,I58345,I58342,I58354,I58339,I58351,I58336,I58357,I58403,I58406,I58409,I58412,I58415,I58418,I58421,I58424,I58427,I2224,I2231);
PAT_5 I_795 (I58406,I58403,I58409,I58427,I58424,I58412,I58421,I58415,I58406,I58418,I58403,I58473,I58476,I58479,I58482,I58485,I58488,I58491,I58494,I58497,I58500,I2224,I2231);
PAT_6 I_796 (I58491,I58485,I58473,I58479,I58476,I58482,I58488,I58473,I58497,I58494,I58500,I58546,I58549,I58552,I58555,I58558,I58561,I58564,I58567,I58570,I58573,I2224,I2231);
PAT_11 I_797 (I58546,I58561,I58546,I58558,I58555,I58573,I58570,I58567,I58564,I58549,I58552,I58619,I58622,I58625,I58628,I58631,I58634,I58637,I58640,I58643,I58646,I2224,I2231);
PAT_5 I_798 (I58640,I58619,I58646,I58634,I58631,I58643,I58625,I58619,I58637,I58622,I58628,I58692,I58695,I58698,I58701,I58704,I58707,I58710,I58713,I58716,I58719,I2224,I2231);
PAT_9 I_799 (I58707,I58704,I58713,I58710,I58701,I58692,I58698,I58719,I58695,I58716,I58692,I58765,I58768,I58771,I58774,I58777,I58780,I58783,I58786,I58789,I2224,I2231);
PAT_6 I_800 (I58783,I58765,I58777,I58786,I58765,I58774,I58771,I58789,I58780,I58768,I58768,I58835,I58838,I58841,I58844,I58847,I58850,I58853,I58856,I58859,I58862,I2224,I2231);
PAT_9 I_801 (I58835,I58862,I58859,I58841,I58847,I58838,I58850,I58835,I58853,I58844,I58856,I58908,I58911,I58914,I58917,I58920,I58923,I58926,I58929,I58932,I2224,I2231);
PAT_10 I_802 (I58929,I58926,I58914,I58911,I58932,I58917,I58923,I58911,I58908,I58908,I58920,I58978,I58981,I58984,I58987,I58990,I58993,I58996,I58999,I2224,I2231);
PAT_2 I_803 (I58990,I58993,I58984,I58996,I58981,I58978,I58978,I58984,I58999,I58987,I58981,I59045,I59048,I59051,I59054,I59057,I59060,I59063,I59066,I59069,I2224,I2231);
PAT_8 I_804 (I59057,I59048,I59054,I59045,I59051,I59066,I59063,I59045,I59060,I59048,I59069,I59115,I59118,I59121,I59124,I59127,I59130,I59133,I59136,I59139,I2224,I2231);
PAT_17 I_805 (I59139,I59127,I59124,I59118,I59121,I59133,I59115,I59118,I59115,I59130,I59136,I59185,I59188,I59191,I59194,I59197,I59200,I59203,I59206,I59209,I59212,I2224,I2231);
PAT_12 I_806 (I59209,I59191,I59185,I59203,I59197,I59206,I59188,I59212,I59185,I59194,I59200,I59258,I59261,I59264,I59267,I59270,I59273,I59276,I59279,I2224,I2231);
PAT_0 I_807 (I59270,I59273,I59279,I59258,I59267,I59261,I59258,I59264,I59261,I59264,I59276,I59325,I59328,I59331,I59334,I59337,I59340,I59343,I59346,I2224,I2231);
PAT_13 I_808 (I59334,I59343,I59325,I59328,I59328,I59331,I59337,I59331,I59325,I59340,I59346,I59392,I59395,I59398,I59401,I59404,I59407,I59410,I59413,I59416,I2224,I2231);
PAT_5 I_809 (I59404,I59395,I59401,I59413,I59395,I59416,I59398,I59407,I59392,I59392,I59410,I59462,I59465,I59468,I59471,I59474,I59477,I59480,I59483,I59486,I59489,I2224,I2231);
PAT_1 I_810 (I59477,I59465,I59483,I59462,I59468,I59462,I59471,I59486,I59480,I59489,I59474,I59535,I59538,I59541,I59544,I59547,I59550,I59553,I59556,I59559,I2224,I2231);
PAT_13 I_811 (I59544,I59553,I59559,I59535,I59550,I59547,I59556,I59541,I59538,I59535,I59538,I59605,I59608,I59611,I59614,I59617,I59620,I59623,I59626,I59629,I2224,I2231);
PAT_5 I_812 (I59617,I59608,I59614,I59626,I59608,I59629,I59611,I59620,I59605,I59605,I59623,I59675,I59678,I59681,I59684,I59687,I59690,I59693,I59696,I59699,I59702,I2224,I2231);
PAT_17 I_813 (I59702,I59678,I59681,I59684,I59675,I59687,I59675,I59699,I59693,I59690,I59696,I59748,I59751,I59754,I59757,I59760,I59763,I59766,I59769,I59772,I59775,I2224,I2231);
PAT_13 I_814 (I59766,I59769,I59754,I59748,I59760,I59772,I59751,I59763,I59748,I59775,I59757,I59821,I59824,I59827,I59830,I59833,I59836,I59839,I59842,I59845,I2224,I2231);
PAT_6 I_815 (I59821,I59833,I59830,I59842,I59839,I59845,I59821,I59836,I59824,I59824,I59827,I59891,I59894,I59897,I59900,I59903,I59906,I59909,I59912,I59915,I59918,I2224,I2231);
PAT_11 I_816 (I59891,I59906,I59891,I59903,I59900,I59918,I59915,I59912,I59909,I59894,I59897,I59964,I59967,I59970,I59973,I59976,I59979,I59982,I59985,I59988,I59991,I2224,I2231);
PAT_13 I_817 (I59964,I59967,I59976,I59988,I59991,I59979,I59985,I59973,I59982,I59970,I59964,I60037,I60040,I60043,I60046,I60049,I60052,I60055,I60058,I60061,I2224,I2231);
PAT_6 I_818 (I60037,I60049,I60046,I60058,I60055,I60061,I60037,I60052,I60040,I60040,I60043,I60107,I60110,I60113,I60116,I60119,I60122,I60125,I60128,I60131,I60134,I2224,I2231);
PAT_13 I_819 (I60131,I60113,I60128,I60107,I60110,I60116,I60134,I60119,I60125,I60107,I60122,I60180,I60183,I60186,I60189,I60192,I60195,I60198,I60201,I60204,I2224,I2231);
PAT_15 I_820 (I60180,I60192,I60183,I60195,I60180,I60189,I60204,I60201,I60186,I60198,I60183,I60250,I60253,I60256,I60259,I60262,I60265,I60268,I60271,I60274,I2224,I2231);
PAT_2 I_821 (I60253,I60253,I60256,I60262,I60250,I60250,I60259,I60274,I60268,I60271,I60265,I60320,I60323,I60326,I60329,I60332,I60335,I60338,I60341,I60344,I2224,I2231);
PAT_9 I_822 (I60335,I60344,I60320,I60326,I60329,I60338,I60323,I60332,I60341,I60323,I60320,I60390,I60393,I60396,I60399,I60402,I60405,I60408,I60411,I60414,I2224,I2231);
PAT_11 I_823 (I60402,I60408,I60414,I60411,I60399,I60393,I60393,I60390,I60405,I60390,I60396,I60460,I60463,I60466,I60469,I60472,I60475,I60478,I60481,I60484,I60487,I2224,I2231);
PAT_13 I_824 (I60460,I60463,I60472,I60484,I60487,I60475,I60481,I60469,I60478,I60466,I60460,I60533,I60536,I60539,I60542,I60545,I60548,I60551,I60554,I60557,I2224,I2231);
PAT_9 I_825 (I60554,I60536,I60536,I60533,I60557,I60539,I60542,I60533,I60545,I60551,I60548,I60603,I60606,I60609,I60612,I60615,I60618,I60621,I60624,I60627,I2224,I2231);
PAT_4 I_826 (I60603,I60627,I60621,I60609,I60606,I60624,I60606,I60603,I60618,I60612,I60615,I60673,I60676,I60679,I60682,I60685,I60688,I60691,I60694,I60697,I2224,I2231);
PAT_2 I_827 (I60682,I60676,I60676,I60697,I60673,I60691,I60688,I60679,I60673,I60685,I60694,I60743,I60746,I60749,I60752,I60755,I60758,I60761,I60764,I60767,I2224,I2231);
PAT_7 I_828 (I60767,I60743,I60749,I60746,I60746,I60755,I60758,I60743,I60761,I60764,I60752,I60813,I60816,I60819,I60822,I60825,I60828,I60831,I60834,I60837,I2224,I2231);
PAT_5 I_829 (I60819,I60813,I60822,I60831,I60825,I60837,I60834,I60816,I60828,I60816,I60813,I60883,I60886,I60889,I60892,I60895,I60898,I60901,I60904,I60907,I60910,I2224,I2231);
PAT_12 I_830 (I60910,I60898,I60883,I60907,I60886,I60883,I60889,I60892,I60895,I60901,I60904,I60956,I60959,I60962,I60965,I60968,I60971,I60974,I60977,I2224,I2231);
PAT_2 I_831 (I60974,I60968,I60977,I60971,I60965,I60962,I60956,I60956,I60962,I60959,I60959,I61023,I61026,I61029,I61032,I61035,I61038,I61041,I61044,I61047,I2224,I2231);
PAT_9 I_832 (I61038,I61047,I61023,I61029,I61032,I61041,I61026,I61035,I61044,I61026,I61023,I61093,I61096,I61099,I61102,I61105,I61108,I61111,I61114,I61117,I2224,I2231);
PAT_0 I_833 (I61102,I61114,I61093,I61096,I61099,I61093,I61108,I61111,I61105,I61117,I61096,I61163,I61166,I61169,I61172,I61175,I61178,I61181,I61184,I2224,I2231);
PAT_6 I_834 (I61175,I61169,I61166,I61163,I61169,I61166,I61163,I61184,I61172,I61181,I61178,I61230,I61233,I61236,I61239,I61242,I61245,I61248,I61251,I61254,I61257,I2224,I2231);
PAT_12 I_835 (I61230,I61257,I61236,I61239,I61233,I61230,I61251,I61245,I61248,I61242,I61254,I61303,I61306,I61309,I61312,I61315,I61318,I61321,I61324,I2224,I2231);
PAT_6 I_836 (I61312,I61306,I61324,I61309,I61306,I61309,I61318,I61303,I61321,I61303,I61315,I61370,I61373,I61376,I61379,I61382,I61385,I61388,I61391,I61394,I61397,I2224,I2231);
PAT_13 I_837 (I1745,I2177,I2153,I1361,I1785,I2169,I1377,I1529,I1401,I1425,I1753,I61443,I61446,I61449,I61452,I61455,I61458,I61461,I61464,I61467,I2224,I2231);
PAT_14 I_838 (I61446,I61461,I61449,I61458,I61452,I61443,I61455,I61464,I61443,I61467,I61446,I61513,I61516,I61519,I61522,I61525,I61528,I61531,I61534,I61537,I2224,I2231);
PAT_10 I_839 (I61516,I61513,I61519,I61537,I61534,I61528,I61516,I61531,I61513,I61525,I61522,I61583,I61586,I61589,I61592,I61595,I61598,I61601,I61604,I2224,I2231);
PAT_8 I_840 (I61604,I61595,I61586,I61583,I61592,I61583,I61598,I61586,I61601,I61589,I61589,I61650,I61653,I61656,I61659,I61662,I61665,I61668,I61671,I61674,I2224,I2231);
PAT_6 I_841 (I61653,I61650,I61656,I61668,I61665,I61659,I61662,I61650,I61671,I61653,I61674,I61720,I61723,I61726,I61729,I61732,I61735,I61738,I61741,I61744,I61747,I2224,I2231);
PAT_9 I_842 (I61720,I61747,I61744,I61726,I61732,I61723,I61735,I61720,I61738,I61729,I61741,I61793,I61796,I61799,I61802,I61805,I61808,I61811,I61814,I61817,I2224,I2231);
PAT_11 I_843 (I61805,I61811,I61817,I61814,I61802,I61796,I61796,I61793,I61808,I61793,I61799,I61863,I61866,I61869,I61872,I61875,I61878,I61881,I61884,I61887,I61890,I2224,I2231);
PAT_5 I_844 (I61884,I61863,I61890,I61878,I61875,I61887,I61869,I61863,I61881,I61866,I61872,I61936,I61939,I61942,I61945,I61948,I61951,I61954,I61957,I61960,I61963,I2224,I2231);
PAT_6 I_845 (I61954,I61948,I61936,I61942,I61939,I61945,I61951,I61936,I61960,I61957,I61963,I62009,I62012,I62015,I62018,I62021,I62024,I62027,I62030,I62033,I62036,I2224,I2231);
PAT_2 I_846 (I62030,I62036,I62018,I62024,I62009,I62015,I62009,I62021,I62012,I62027,I62033,I62082,I62085,I62088,I62091,I62094,I62097,I62100,I62103,I62106,I2224,I2231);
PAT_13 I_847 (I62091,I62085,I62082,I62103,I62094,I62097,I62085,I62088,I62100,I62106,I62082,I62152,I62155,I62158,I62161,I62164,I62167,I62170,I62173,I62176,I2224,I2231);
PAT_9 I_848 (I62173,I62155,I62155,I62152,I62176,I62158,I62161,I62152,I62164,I62170,I62167,I62222,I62225,I62228,I62231,I62234,I62237,I62240,I62243,I62246,I2224,I2231);
PAT_4 I_849 (I62222,I62246,I62240,I62228,I62225,I62243,I62225,I62222,I62237,I62231,I62234,I62292,I62295,I62298,I62301,I62304,I62307,I62310,I62313,I62316,I2224,I2231);
PAT_7 I_850 (I62307,I62301,I62298,I62292,I62304,I62310,I62295,I62295,I62313,I62316,I62292,I62362,I62365,I62368,I62371,I62374,I62377,I62380,I62383,I62386,I2224,I2231);
PAT_16 I_851 (I62386,I62362,I62380,I62368,I62377,I62371,I62362,I62383,I62365,I62374,I62365,I62432,I62435,I62438,I62441,I62444,I62447,I62450,I62453,I62456,I62459,I2224,I2231);
PAT_9 I_852 (I62450,I62432,I62432,I62441,I62438,I62456,I62459,I62435,I62453,I62447,I62444,I62505,I62508,I62511,I62514,I62517,I62520,I62523,I62526,I62529,I2224,I2231);
PAT_4 I_853 (I62505,I62529,I62523,I62511,I62508,I62526,I62508,I62505,I62520,I62514,I62517,I62575,I62578,I62581,I62584,I62587,I62590,I62593,I62596,I62599,I2224,I2231);
PAT_14 I_854 (I62578,I62593,I62590,I62575,I62587,I62578,I62575,I62581,I62596,I62584,I62599,I62645,I62648,I62651,I62654,I62657,I62660,I62663,I62666,I62669,I2224,I2231);
PAT_15 I_855 (I62657,I62651,I62648,I62666,I62663,I62654,I62645,I62648,I62645,I62660,I62669,I62715,I62718,I62721,I62724,I62727,I62730,I62733,I62736,I62739,I2224,I2231);
PAT_8 I_856 (I62736,I62715,I62715,I62724,I62721,I62718,I62733,I62730,I62718,I62739,I62727,I62785,I62788,I62791,I62794,I62797,I62800,I62803,I62806,I62809,I2224,I2231);
PAT_16 I_857 (I62806,I62785,I62785,I62794,I62791,I62803,I62788,I62797,I62800,I62809,I62788,I62855,I62858,I62861,I62864,I62867,I62870,I62873,I62876,I62879,I62882,I2224,I2231);
PAT_6 I_858 (I62855,I62858,I62867,I62873,I62861,I62882,I62864,I62876,I62879,I62870,I62855,I62928,I62931,I62934,I62937,I62940,I62943,I62946,I62949,I62952,I62955,I2224,I2231);
PAT_8 I_859 (I62937,I62943,I62934,I62946,I62928,I62931,I62949,I62928,I62955,I62952,I62940,I63001,I63004,I63007,I63010,I63013,I63016,I63019,I63022,I63025,I2224,I2231);
PAT_17 I_860 (I63025,I63013,I63010,I63004,I63007,I63019,I63001,I63004,I63001,I63016,I63022,I63071,I63074,I63077,I63080,I63083,I63086,I63089,I63092,I63095,I63098,I2224,I2231);
PAT_11 I_861 (I63083,I63092,I63098,I63074,I63071,I63089,I63080,I63086,I63077,I63095,I63071,I63144,I63147,I63150,I63153,I63156,I63159,I63162,I63165,I63168,I63171,I2224,I2231);
PAT_5 I_862 (I63165,I63144,I63171,I63159,I63156,I63168,I63150,I63144,I63162,I63147,I63153,I63217,I63220,I63223,I63226,I63229,I63232,I63235,I63238,I63241,I63244,I2224,I2231);
PAT_7 I_863 (I63235,I63238,I63244,I63241,I63226,I63223,I63217,I63229,I63217,I63220,I63232,I63290,I63293,I63296,I63299,I63302,I63305,I63308,I63311,I63314,I2224,I2231);
PAT_4 I_864 (I63314,I63290,I63290,I63305,I63299,I63293,I63293,I63308,I63311,I63296,I63302,I63360,I63363,I63366,I63369,I63372,I63375,I63378,I63381,I63384,I2224,I2231);
PAT_2 I_865 (I63369,I63363,I63363,I63384,I63360,I63378,I63375,I63366,I63360,I63372,I63381,I63430,I63433,I63436,I63439,I63442,I63445,I63448,I63451,I63454,I2224,I2231);
PAT_11 I_866 (I63433,I63445,I63430,I63442,I63439,I63451,I63448,I63433,I63454,I63436,I63430,I63500,I63503,I63506,I63509,I63512,I63515,I63518,I63521,I63524,I63527,I2224,I2231);
PAT_2 I_867 (I63500,I63524,I63512,I63506,I63515,I63518,I63503,I63527,I63521,I63509,I63500,I63573,I63576,I63579,I63582,I63585,I63588,I63591,I63594,I63597,I2224,I2231);
PAT_11 I_868 (I63576,I63588,I63573,I63585,I63582,I63594,I63591,I63576,I63597,I63579,I63573,I63643,I63646,I63649,I63652,I63655,I63658,I63661,I63664,I63667,I63670,I2224,I2231);
PAT_9 I_869 (I63649,I63661,I63652,I63664,I63643,I63646,I63655,I63643,I63658,I63667,I63670,I63716,I63719,I63722,I63725,I63728,I63731,I63734,I63737,I63740,I2224,I2231);
PAT_5 I_870 (I63737,I63716,I63731,I63716,I63722,I63725,I63719,I63719,I63734,I63728,I63740,I63786,I63789,I63792,I63795,I63798,I63801,I63804,I63807,I63810,I63813,I2224,I2231);
PAT_2 I_871 (I63801,I63786,I63798,I63792,I63807,I63789,I63804,I63795,I63810,I63813,I63786,I63859,I63862,I63865,I63868,I63871,I63874,I63877,I63880,I63883,I2224,I2231);
PAT_9 I_872 (I63874,I63883,I63859,I63865,I63868,I63877,I63862,I63871,I63880,I63862,I63859,I63929,I63932,I63935,I63938,I63941,I63944,I63947,I63950,I63953,I2224,I2231);
PAT_14 I_873 (I63938,I63929,I63953,I63935,I63932,I63929,I63944,I63950,I63941,I63932,I63947,I63999,I64002,I64005,I64008,I64011,I64014,I64017,I64020,I64023,I2224,I2231);
PAT_17 I_874 (I64014,I64002,I64023,I63999,I64020,I64008,I64005,I64017,I64011,I64002,I63999,I64069,I64072,I64075,I64078,I64081,I64084,I64087,I64090,I64093,I64096,I2224,I2231);
PAT_11 I_875 (I64081,I64090,I64096,I64072,I64069,I64087,I64078,I64084,I64075,I64093,I64069,I64142,I64145,I64148,I64151,I64154,I64157,I64160,I64163,I64166,I64169,I2224,I2231);
PAT_10 I_876 (I64157,I64163,I64154,I64148,I64166,I64151,I64169,I64160,I64142,I64145,I64142,I64215,I64218,I64221,I64224,I64227,I64230,I64233,I64236,I2224,I2231);
PAT_4 I_877 (I64230,I64227,I64218,I64236,I64215,I64218,I64224,I64221,I64233,I64215,I64221,I64282,I64285,I64288,I64291,I64294,I64297,I64300,I64303,I64306,I2224,I2231);
PAT_9 I_878 (I64303,I64285,I64288,I64297,I64300,I64282,I64291,I64285,I64306,I64282,I64294,I64352,I64355,I64358,I64361,I64364,I64367,I64370,I64373,I64376,I2224,I2231);
PAT_6 I_879 (I64370,I64352,I64364,I64373,I64352,I64361,I64358,I64376,I64367,I64355,I64355,I64422,I64425,I64428,I64431,I64434,I64437,I64440,I64443,I64446,I64449,I2224,I2231);
PAT_12 I_880 (I64422,I64449,I64428,I64431,I64425,I64422,I64443,I64437,I64440,I64434,I64446,I64495,I64498,I64501,I64504,I64507,I64510,I64513,I64516,I2224,I2231);
PAT_5 I_881 (I64504,I64510,I64516,I64501,I64501,I64495,I64513,I64495,I64498,I64498,I64507,I64562,I64565,I64568,I64571,I64574,I64577,I64580,I64583,I64586,I64589,I2224,I2231);
PAT_2 I_882 (I64577,I64562,I64574,I64568,I64583,I64565,I64580,I64571,I64586,I64589,I64562,I64635,I64638,I64641,I64644,I64647,I64650,I64653,I64656,I64659,I2224,I2231);
PAT_13 I_883 (I64644,I64638,I64635,I64656,I64647,I64650,I64638,I64641,I64653,I64659,I64635,I64705,I64708,I64711,I64714,I64717,I64720,I64723,I64726,I64729,I2224,I2231);
PAT_5 I_884 (I64717,I64708,I64714,I64726,I64708,I64729,I64711,I64720,I64705,I64705,I64723,I64775,I64778,I64781,I64784,I64787,I64790,I64793,I64796,I64799,I64802,I2224,I2231);
PAT_17 I_885 (I64802,I64778,I64781,I64784,I64775,I64787,I64775,I64799,I64793,I64790,I64796,I64848,I64851,I64854,I64857,I64860,I64863,I64866,I64869,I64872,I64875,I2224,I2231);
PAT_9 I_886 (I64869,I64851,I64857,I64872,I64854,I64866,I64848,I64860,I64848,I64875,I64863,I64921,I64924,I64927,I64930,I64933,I64936,I64939,I64942,I64945,I2224,I2231);
PAT_2 I_887 (I64936,I64939,I64930,I64945,I64921,I64924,I64927,I64924,I64942,I64933,I64921,I64991,I64994,I64997,I65000,I65003,I65006,I65009,I65012,I65015,I2224,I2231);
PAT_9 I_888 (I65006,I65015,I64991,I64997,I65000,I65009,I64994,I65003,I65012,I64994,I64991,I65061,I65064,I65067,I65070,I65073,I65076,I65079,I65082,I65085,I2224,I2231);
PAT_4 I_889 (I65061,I65085,I65079,I65067,I65064,I65082,I65064,I65061,I65076,I65070,I65073,I65131,I65134,I65137,I65140,I65143,I65146,I65149,I65152,I65155,I2224,I2231);
PAT_6 I_890 (I65131,I65137,I65134,I65146,I65149,I65143,I65155,I65152,I65131,I65140,I65134,I65201,I65204,I65207,I65210,I65213,I65216,I65219,I65222,I65225,I65228,I2224,I2231);
PAT_13 I_891 (I65225,I65207,I65222,I65201,I65204,I65210,I65228,I65213,I65219,I65201,I65216,I65274,I65277,I65280,I65283,I65286,I65289,I65292,I65295,I65298,I2224,I2231);
PAT_11 I_892 (I65274,I65286,I65289,I65280,I65277,I65298,I65277,I65295,I65283,I65274,I65292,I65344,I65347,I65350,I65353,I65356,I65359,I65362,I65365,I65368,I65371,I2224,I2231);
PAT_10 I_893 (I65359,I65365,I65356,I65350,I65368,I65353,I65371,I65362,I65344,I65347,I65344,I65417,I65420,I65423,I65426,I65429,I65432,I65435,I65438,I2224,I2231);
PAT_5 I_894 (I65438,I65417,I65426,I65420,I65435,I65432,I65423,I65423,I65417,I65420,I65429,I65484,I65487,I65490,I65493,I65496,I65499,I65502,I65505,I65508,I65511,I2224,I2231);
PAT_10 I_895 (I65508,I65511,I65490,I65496,I65499,I65505,I65487,I65484,I65484,I65493,I65502,I65557,I65560,I65563,I65566,I65569,I65572,I65575,I65578,I2224,I2231);
PAT_13 I_896 (I65563,I65569,I65563,I65560,I65575,I65578,I65557,I65557,I65572,I65560,I65566,I65624,I65627,I65630,I65633,I65636,I65639,I65642,I65645,I65648,I2224,I2231);
PAT_5 I_897 (I65636,I65627,I65633,I65645,I65627,I65648,I65630,I65639,I65624,I65624,I65642,I65694,I65697,I65700,I65703,I65706,I65709,I65712,I65715,I65718,I65721,I2224,I2231);
PAT_10 I_898 (I65718,I65721,I65700,I65706,I65709,I65715,I65697,I65694,I65694,I65703,I65712,I65767,I65770,I65773,I65776,I65779,I65782,I65785,I65788,I2224,I2231);
PAT_13 I_899 (I65773,I65779,I65773,I65770,I65785,I65788,I65767,I65767,I65782,I65770,I65776,I65834,I65837,I65840,I65843,I65846,I65849,I65852,I65855,I65858,I2224,I2231);
PAT_9 I_900 (I65855,I65837,I65837,I65834,I65858,I65840,I65843,I65834,I65846,I65852,I65849,I65904,I65907,I65910,I65913,I65916,I65919,I65922,I65925,I65928,I2224,I2231);
PAT_1 I_901 (I65904,I65922,I65904,I65916,I65907,I65913,I65919,I65925,I65928,I65910,I65907,I65974,I65977,I65980,I65983,I65986,I65989,I65992,I65995,I65998,I2224,I2231);
PAT_6 I_902 (I65983,I65974,I65977,I65980,I65995,I65998,I65992,I65974,I65989,I65986,I65977,I66044,I66047,I66050,I66053,I66056,I66059,I66062,I66065,I66068,I66071,I2224,I2231);
PAT_5 I_903 (I66065,I66044,I66050,I66053,I66059,I66062,I66044,I66068,I66047,I66056,I66071,I66117,I66120,I66123,I66126,I66129,I66132,I66135,I66138,I66141,I66144,I2224,I2231);
PAT_7 I_904 (I66135,I66138,I66144,I66141,I66126,I66123,I66117,I66129,I66117,I66120,I66132,I66190,I66193,I66196,I66199,I66202,I66205,I66208,I66211,I66214,I2224,I2231);
PAT_14 I_905 (I66205,I66199,I66190,I66193,I66202,I66208,I66196,I66211,I66193,I66190,I66214,I66260,I66263,I66266,I66269,I66272,I66275,I66278,I66281,I66284,I2224,I2231);
PAT_9 I_906 (I66269,I66281,I66260,I66278,I66263,I66266,I66284,I66263,I66272,I66260,I66275,I66330,I66333,I66336,I66339,I66342,I66345,I66348,I66351,I66354,I2224,I2231);
PAT_11 I_907 (I66342,I66348,I66354,I66351,I66339,I66333,I66333,I66330,I66345,I66330,I66336,I66400,I66403,I66406,I66409,I66412,I66415,I66418,I66421,I66424,I66427,I2224,I2231);
PAT_16 I_908 (I66409,I66415,I66421,I66427,I66412,I66403,I66400,I66400,I66418,I66424,I66406,I66473,I66476,I66479,I66482,I66485,I66488,I66491,I66494,I66497,I66500,I2224,I2231);
PAT_8 I_909 (I66473,I66476,I66485,I66494,I66482,I66497,I66500,I66488,I66479,I66491,I66473,I66546,I66549,I66552,I66555,I66558,I66561,I66564,I66567,I66570,I2224,I2231);
PAT_7 I_910 (I66546,I66555,I66552,I66558,I66564,I66546,I66549,I66567,I66570,I66561,I66549,I66616,I66619,I66622,I66625,I66628,I66631,I66634,I66637,I66640,I2224,I2231);
PAT_10 I_911 (I66616,I66619,I66616,I66637,I66625,I66628,I66619,I66640,I66631,I66622,I66634,I66686,I66689,I66692,I66695,I66698,I66701,I66704,I66707,I2224,I2231);
PAT_11 I_912 (I66695,I66698,I66707,I66701,I66704,I66686,I66686,I66692,I66689,I66689,I66692,I66753,I66756,I66759,I66762,I66765,I66768,I66771,I66774,I66777,I66780,I2224,I2231);
PAT_13 I_913 (I66753,I66756,I66765,I66777,I66780,I66768,I66774,I66762,I66771,I66759,I66753,I66826,I66829,I66832,I66835,I66838,I66841,I66844,I66847,I66850,I2224,I2231);
PAT_9 I_914 (I66847,I66829,I66829,I66826,I66850,I66832,I66835,I66826,I66838,I66844,I66841,I66896,I66899,I66902,I66905,I66908,I66911,I66914,I66917,I66920,I2224,I2231);
PAT_10 I_915 (I66917,I66914,I66902,I66899,I66920,I66905,I66911,I66899,I66896,I66896,I66908,I66966,I66969,I66972,I66975,I66978,I66981,I66984,I66987,I2224,I2231);
PAT_2 I_916 (I66978,I66981,I66972,I66984,I66969,I66966,I66966,I66972,I66987,I66975,I66969,I67033,I67036,I67039,I67042,I67045,I67048,I67051,I67054,I67057,I2224,I2231);
PAT_14 I_917 (I67039,I67042,I67057,I67048,I67033,I67036,I67051,I67045,I67033,I67054,I67036,I67103,I67106,I67109,I67112,I67115,I67118,I67121,I67124,I67127,I2224,I2231);
PAT_5 I_918 (I67106,I67109,I67106,I67115,I67103,I67124,I67112,I67103,I67127,I67121,I67118,I67173,I67176,I67179,I67182,I67185,I67188,I67191,I67194,I67197,I67200,I2224,I2231);
PAT_9 I_919 (I67188,I67185,I67194,I67191,I67182,I67173,I67179,I67200,I67176,I67197,I67173,I67246,I67249,I67252,I67255,I67258,I67261,I67264,I67267,I67270,I2224,I2231);
PAT_17 I_920 (I67249,I67255,I67270,I67261,I67264,I67252,I67246,I67258,I67246,I67249,I67267,I67316,I67319,I67322,I67325,I67328,I67331,I67334,I67337,I67340,I67343,I2224,I2231);
PAT_2 I_921 (I67316,I67334,I67331,I67316,I67325,I67340,I67337,I67322,I67343,I67328,I67319,I67389,I67392,I67395,I67398,I67401,I67404,I67407,I67410,I67413,I2224,I2231);
PAT_9 I_922 (I67404,I67413,I67389,I67395,I67398,I67407,I67392,I67401,I67410,I67392,I67389,I67459,I67462,I67465,I67468,I67471,I67474,I67477,I67480,I67483,I2224,I2231);
PAT_17 I_923 (I67462,I67468,I67483,I67474,I67477,I67465,I67459,I67471,I67459,I67462,I67480,I67529,I67532,I67535,I67538,I67541,I67544,I67547,I67550,I67553,I67556,I2224,I2231);
PAT_12 I_924 (I67553,I67535,I67529,I67547,I67541,I67550,I67532,I67556,I67529,I67538,I67544,I67602,I67605,I67608,I67611,I67614,I67617,I67620,I67623,I2224,I2231);
PAT_10 I_925 (I67602,I67623,I67614,I67617,I67608,I67605,I67602,I67620,I67608,I67611,I67605,I67669,I67672,I67675,I67678,I67681,I67684,I67687,I67690,I2224,I2231);
PAT_9 I_926 (I67681,I67669,I67672,I67675,I67669,I67675,I67678,I67672,I67690,I67684,I67687,I67736,I67739,I67742,I67745,I67748,I67751,I67754,I67757,I67760,I2224,I2231);
PAT_15 I_927 (I67748,I67757,I67760,I67739,I67754,I67742,I67745,I67736,I67751,I67736,I67739,I67806,I67809,I67812,I67815,I67818,I67821,I67824,I67827,I67830,I2224,I2231);
PAT_4 I_928 (I67818,I67824,I67806,I67809,I67812,I67806,I67830,I67827,I67815,I67821,I67809,I67876,I67879,I67882,I67885,I67888,I67891,I67894,I67897,I67900,I2224,I2231);
PAT_9 I_929 (I67897,I67879,I67882,I67891,I67894,I67876,I67885,I67879,I67900,I67876,I67888,I67946,I67949,I67952,I67955,I67958,I67961,I67964,I67967,I67970,I2224,I2231);
PAT_14 I_930 (I67955,I67946,I67970,I67952,I67949,I67946,I67961,I67967,I67958,I67949,I67964,I68016,I68019,I68022,I68025,I68028,I68031,I68034,I68037,I68040,I2224,I2231);
PAT_8 I_931 (I68022,I68025,I68019,I68031,I68040,I68019,I68016,I68037,I68016,I68028,I68034,I68086,I68089,I68092,I68095,I68098,I68101,I68104,I68107,I68110,I2224,I2231);
PAT_11 I_932 (I68107,I68098,I68086,I68089,I68104,I68092,I68095,I68086,I68110,I68101,I68089,I68156,I68159,I68162,I68165,I68168,I68171,I68174,I68177,I68180,I68183,I2224,I2231);
PAT_17 I_933 (I68168,I68159,I68183,I68156,I68165,I68177,I68174,I68171,I68156,I68180,I68162,I68229,I68232,I68235,I68238,I68241,I68244,I68247,I68250,I68253,I68256,I2224,I2231);
PAT_7 I_934 (I68247,I68238,I68244,I68232,I68241,I68250,I68256,I68229,I68253,I68235,I68229,I68302,I68305,I68308,I68311,I68314,I68317,I68320,I68323,I68326,I2224,I2231);
PAT_17 I_935 (I68314,I68308,I68317,I68302,I68320,I68323,I68305,I68326,I68311,I68305,I68302,I68372,I68375,I68378,I68381,I68384,I68387,I68390,I68393,I68396,I68399,I2224,I2231);
PAT_6 I_936 (I68372,I68390,I68378,I68381,I68387,I68372,I68384,I68375,I68396,I68399,I68393,I68445,I68448,I68451,I68454,I68457,I68460,I68463,I68466,I68469,I68472,I2224,I2231);
PAT_12 I_937 (I68445,I68472,I68451,I68454,I68448,I68445,I68466,I68460,I68463,I68457,I68469,I68518,I68521,I68524,I68527,I68530,I68533,I68536,I68539,I2224,I2231);
PAT_10 I_938 (I68518,I68539,I68530,I68533,I68524,I68521,I68518,I68536,I68524,I68527,I68521,I68585,I68588,I68591,I68594,I68597,I68600,I68603,I68606,I2224,I2231);
PAT_11 I_939 (I68594,I68597,I68606,I68600,I68603,I68585,I68585,I68591,I68588,I68588,I68591,I68652,I68655,I68658,I68661,I68664,I68667,I68670,I68673,I68676,I68679,I2224,I2231);
PAT_13 I_940 (I68652,I68655,I68664,I68676,I68679,I68667,I68673,I68661,I68670,I68658,I68652,I68725,I68728,I68731,I68734,I68737,I68740,I68743,I68746,I68749,I2224,I2231);
PAT_11 I_941 (I68725,I68737,I68740,I68731,I68728,I68749,I68728,I68746,I68734,I68725,I68743,I68795,I68798,I68801,I68804,I68807,I68810,I68813,I68816,I68819,I68822,I2224,I2231);
PAT_4 I_942 (I68801,I68822,I68795,I68813,I68804,I68795,I68816,I68798,I68807,I68819,I68810,I68868,I68871,I68874,I68877,I68880,I68883,I68886,I68889,I68892,I2224,I2231);
PAT_6 I_943 (I68868,I68874,I68871,I68883,I68886,I68880,I68892,I68889,I68868,I68877,I68871,I68938,I68941,I68944,I68947,I68950,I68953,I68956,I68959,I68962,I68965,I2224,I2231);
PAT_9 I_944 (I68938,I68965,I68962,I68944,I68950,I68941,I68953,I68938,I68956,I68947,I68959,I69011,I69014,I69017,I69020,I69023,I69026,I69029,I69032,I69035,I2224,I2231);
PAT_8 I_945 (I69032,I69020,I69029,I69011,I69014,I69026,I69035,I69014,I69017,I69023,I69011,I69081,I69084,I69087,I69090,I69093,I69096,I69099,I69102,I69105,I2224,I2231);
PAT_4 I_946 (I69099,I69084,I69090,I69081,I69081,I69093,I69084,I69102,I69105,I69087,I69096,I69151,I69154,I69157,I69160,I69163,I69166,I69169,I69172,I69175,I2224,I2231);
PAT_2 I_947 (I69160,I69154,I69154,I69175,I69151,I69169,I69166,I69157,I69151,I69163,I69172,I69221,I69224,I69227,I69230,I69233,I69236,I69239,I69242,I69245,I2224,I2231);
PAT_8 I_948 (I69233,I69224,I69230,I69221,I69227,I69242,I69239,I69221,I69236,I69224,I69245,I69291,I69294,I69297,I69300,I69303,I69306,I69309,I69312,I69315,I2224,I2231);
PAT_10 I_949 (I69297,I69291,I69294,I69315,I69309,I69294,I69303,I69291,I69312,I69306,I69300,I69361,I69364,I69367,I69370,I69373,I69376,I69379,I69382,I2224,I2231);
PAT_5 I_950 (I69382,I69361,I69370,I69364,I69379,I69376,I69367,I69367,I69361,I69364,I69373,I69428,I69431,I69434,I69437,I69440,I69443,I69446,I69449,I69452,I69455,I2224,I2231);
PAT_9 I_951 (I69443,I69440,I69449,I69446,I69437,I69428,I69434,I69455,I69431,I69452,I69428,I69501,I69504,I69507,I69510,I69513,I69516,I69519,I69522,I69525,I2224,I2231);
PAT_12 I_952 (I69522,I69519,I69513,I69501,I69510,I69501,I69504,I69507,I69525,I69516,I69504,I69571,I69574,I69577,I69580,I69583,I69586,I69589,I69592,I2224,I2231);
PAT_9 I_953 (I69580,I69586,I69571,I69577,I69583,I69574,I69571,I69574,I69592,I69577,I69589,I69638,I69641,I69644,I69647,I69650,I69653,I69656,I69659,I69662,I2224,I2231);
PAT_1 I_954 (I69638,I69656,I69638,I69650,I69641,I69647,I69653,I69659,I69662,I69644,I69641,I69708,I69711,I69714,I69717,I69720,I69723,I69726,I69729,I69732,I2224,I2231);
PAT_9 I_955 (I69723,I69729,I69714,I69732,I69711,I69726,I69711,I69717,I69708,I69720,I69708,I69778,I69781,I69784,I69787,I69790,I69793,I69796,I69799,I69802,I2224,I2231);
PAT_11 I_956 (I69790,I69796,I69802,I69799,I69787,I69781,I69781,I69778,I69793,I69778,I69784,I69848,I69851,I69854,I69857,I69860,I69863,I69866,I69869,I69872,I69875,I2224,I2231);
PAT_8 I_957 (I69857,I69863,I69866,I69872,I69869,I69860,I69848,I69848,I69875,I69851,I69854,I69921,I69924,I69927,I69930,I69933,I69936,I69939,I69942,I69945,I2224,I2231);
PAT_5 I_958 (I69927,I69945,I69921,I69942,I69930,I69933,I69924,I69921,I69924,I69936,I69939,I69991,I69994,I69997,I70000,I70003,I70006,I70009,I70012,I70015,I70018,I2224,I2231);
PAT_6 I_959 (I70009,I70003,I69991,I69997,I69994,I70000,I70006,I69991,I70015,I70012,I70018,I70064,I70067,I70070,I70073,I70076,I70079,I70082,I70085,I70088,I70091,I2224,I2231);
PAT_7 I_960 (I70070,I70079,I70082,I70064,I70073,I70067,I70076,I70091,I70085,I70088,I70064,I70137,I70140,I70143,I70146,I70149,I70152,I70155,I70158,I70161,I2224,I2231);
PAT_2 I_961 (I70158,I70152,I70143,I70137,I70146,I70140,I70149,I70161,I70155,I70140,I70137,I70207,I70210,I70213,I70216,I70219,I70222,I70225,I70228,I70231,I2224,I2231);
PAT_9 I_962 (I70222,I70231,I70207,I70213,I70216,I70225,I70210,I70219,I70228,I70210,I70207,I70277,I70280,I70283,I70286,I70289,I70292,I70295,I70298,I70301,I2224,I2231);
PAT_17 I_963 (I70280,I70286,I70301,I70292,I70295,I70283,I70277,I70289,I70277,I70280,I70298,I70347,I70350,I70353,I70356,I70359,I70362,I70365,I70368,I70371,I70374,I2224,I2231);
PAT_4 I_964 (I70356,I70347,I70365,I70362,I70374,I70371,I70350,I70347,I70353,I70359,I70368,I70420,I70423,I70426,I70429,I70432,I70435,I70438,I70441,I70444,I2224,I2231);
PAT_13 I_965 (I70435,I70429,I70441,I70426,I70432,I70420,I70444,I70438,I70423,I70420,I70423,I70490,I70493,I70496,I70499,I70502,I70505,I70508,I70511,I70514,I2224,I2231);
PAT_10 I_966 (I70511,I70505,I70499,I70493,I70514,I70493,I70502,I70490,I70490,I70508,I70496,I70560,I70563,I70566,I70569,I70572,I70575,I70578,I70581,I2224,I2231);
PAT_15 I_967 (I70575,I70578,I70566,I70572,I70560,I70560,I70566,I70581,I70569,I70563,I70563,I70627,I70630,I70633,I70636,I70639,I70642,I70645,I70648,I70651,I2224,I2231);
PAT_11 I_968 (I70648,I70630,I70627,I70642,I70633,I70627,I70645,I70651,I70639,I70630,I70636,I70697,I70700,I70703,I70706,I70709,I70712,I70715,I70718,I70721,I70724,I2224,I2231);
PAT_4 I_969 (I70703,I70724,I70697,I70715,I70706,I70697,I70718,I70700,I70709,I70721,I70712,I70770,I70773,I70776,I70779,I70782,I70785,I70788,I70791,I70794,I2224,I2231);
PAT_13 I_970 (I70785,I70779,I70791,I70776,I70782,I70770,I70794,I70788,I70773,I70770,I70773,I70840,I70843,I70846,I70849,I70852,I70855,I70858,I70861,I70864,I2224,I2231);
PAT_10 I_971 (I70861,I70855,I70849,I70843,I70864,I70843,I70852,I70840,I70840,I70858,I70846,I70910,I70913,I70916,I70919,I70922,I70925,I70928,I70931,I2224,I2231);
PAT_9 I_972 (I70922,I70910,I70913,I70916,I70910,I70916,I70919,I70913,I70931,I70925,I70928,I70977,I70980,I70983,I70986,I70989,I70992,I70995,I70998,I71001,I2224,I2231);
PAT_7 I_973 (I70983,I70992,I70977,I70998,I70989,I70977,I70980,I71001,I70995,I70980,I70986,I71047,I71050,I71053,I71056,I71059,I71062,I71065,I71068,I71071,I2224,I2231);
PAT_13 I_974 (I71053,I71071,I71062,I71047,I71059,I71047,I71068,I71050,I71056,I71050,I71065,I71117,I71120,I71123,I71126,I71129,I71132,I71135,I71138,I71141,I2224,I2231);
PAT_9 I_975 (I71138,I71120,I71120,I71117,I71141,I71123,I71126,I71117,I71129,I71135,I71132,I71187,I71190,I71193,I71196,I71199,I71202,I71205,I71208,I71211,I2224,I2231);
PAT_17 I_976 (I71190,I71196,I71211,I71202,I71205,I71193,I71187,I71199,I71187,I71190,I71208,I71257,I71260,I71263,I71266,I71269,I71272,I71275,I71278,I71281,I71284,I2224,I2231);
PAT_16 I_977 (I71257,I71281,I71257,I71278,I71275,I71263,I71269,I71260,I71284,I71272,I71266,I71330,I71333,I71336,I71339,I71342,I71345,I71348,I71351,I71354,I71357,I2224,I2231);
PAT_11 I_978 (I71333,I71330,I71357,I71336,I71351,I71354,I71348,I71330,I71339,I71342,I71345,I71403,I71406,I71409,I71412,I71415,I71418,I71421,I71424,I71427,I71430,I2224,I2231);
PAT_16 I_979 (I71412,I71418,I71424,I71430,I71415,I71406,I71403,I71403,I71421,I71427,I71409,I71476,I71479,I71482,I71485,I71488,I71491,I71494,I71497,I71500,I71503,I2224,I2231);
PAT_9 I_980 (I71494,I71476,I71476,I71485,I71482,I71500,I71503,I71479,I71497,I71491,I71488,I71549,I71552,I71555,I71558,I71561,I71564,I71567,I71570,I71573,I2224,I2231);
PAT_13 I_981 (I71549,I71570,I71552,I71567,I71561,I71558,I71573,I71549,I71555,I71564,I71552,I71619,I71622,I71625,I71628,I71631,I71634,I71637,I71640,I71643,I2224,I2231);
PAT_2 I_982 (I71637,I71631,I71628,I71634,I71619,I71643,I71622,I71640,I71619,I71625,I71622,I71689,I71692,I71695,I71698,I71701,I71704,I71707,I71710,I71713,I2224,I2231);
PAT_7 I_983 (I71713,I71689,I71695,I71692,I71692,I71701,I71704,I71689,I71707,I71710,I71698,I71759,I71762,I71765,I71768,I71771,I71774,I71777,I71780,I71783,I2224,I2231);
PAT_10 I_984 (I71759,I71762,I71759,I71780,I71768,I71771,I71762,I71783,I71774,I71765,I71777,I71829,I71832,I71835,I71838,I71841,I71844,I71847,I71850,I2224,I2231);
PAT_13 I_985 (I71835,I71841,I71835,I71832,I71847,I71850,I71829,I71829,I71844,I71832,I71838,I71896,I71899,I71902,I71905,I71908,I71911,I71914,I71917,I71920,I2224,I2231);
PAT_10 I_986 (I71917,I71911,I71905,I71899,I71920,I71899,I71908,I71896,I71896,I71914,I71902,I71966,I71969,I71972,I71975,I71978,I71981,I71984,I71987,I2224,I2231);
PAT_2 I_987 (I71978,I71981,I71972,I71984,I71969,I71966,I71966,I71972,I71987,I71975,I71969,I72033,I72036,I72039,I72042,I72045,I72048,I72051,I72054,I72057,I2224,I2231);
PAT_9 I_988 (I72048,I72057,I72033,I72039,I72042,I72051,I72036,I72045,I72054,I72036,I72033,I72103,I72106,I72109,I72112,I72115,I72118,I72121,I72124,I72127,I2224,I2231);
PAT_17 I_989 (I72106,I72112,I72127,I72118,I72121,I72109,I72103,I72115,I72103,I72106,I72124,I72173,I72176,I72179,I72182,I72185,I72188,I72191,I72194,I72197,I72200,I2224,I2231);
PAT_13 I_990 (I72191,I72194,I72179,I72173,I72185,I72197,I72176,I72188,I72173,I72200,I72182,I72246,I72249,I72252,I72255,I72258,I72261,I72264,I72267,I72270,I2224,I2231);
PAT_11 I_991 (I72246,I72258,I72261,I72252,I72249,I72270,I72249,I72267,I72255,I72246,I72264,I72316,I72319,I72322,I72325,I72328,I72331,I72334,I72337,I72340,I72343,I2224,I2231);
PAT_13 I_992 (I72316,I72319,I72328,I72340,I72343,I72331,I72337,I72325,I72334,I72322,I72316,I72389,I72392,I72395,I72398,I72401,I72404,I72407,I72410,I72413,I2224,I2231);
PAT_2 I_993 (I72407,I72401,I72398,I72404,I72389,I72413,I72392,I72410,I72389,I72395,I72392,I72459,I72462,I72465,I72468,I72471,I72474,I72477,I72480,I72483,I2224,I2231);
PAT_14 I_994 (I72465,I72468,I72483,I72474,I72459,I72462,I72477,I72471,I72459,I72480,I72462,I72529,I72532,I72535,I72538,I72541,I72544,I72547,I72550,I72553,I2224,I2231);
PAT_5 I_995 (I72532,I72535,I72532,I72541,I72529,I72550,I72538,I72529,I72553,I72547,I72544,I72599,I72602,I72605,I72608,I72611,I72614,I72617,I72620,I72623,I72626,I2224,I2231);
PAT_6 I_996 (I72617,I72611,I72599,I72605,I72602,I72608,I72614,I72599,I72623,I72620,I72626,I72672,I72675,I72678,I72681,I72684,I72687,I72690,I72693,I72696,I72699,I2224,I2231);
PAT_11 I_997 (I72672,I72687,I72672,I72684,I72681,I72699,I72696,I72693,I72690,I72675,I72678,I72745,I72748,I72751,I72754,I72757,I72760,I72763,I72766,I72769,I72772,I2224,I2231);
PAT_13 I_998 (I72745,I72748,I72757,I72769,I72772,I72760,I72766,I72754,I72763,I72751,I72745,I72818,I72821,I72824,I72827,I72830,I72833,I72836,I72839,I72842,I2224,I2231);
PAT_8 I_999 (I72827,I72839,I72830,I72833,I72842,I72821,I72836,I72818,I72821,I72824,I72818,I72888,I72891,I72894,I72897,I72900,I72903,I72906,I72909,I72912,I2224,I2231);
PAT_5 I_1000 (I72894,I72912,I72888,I72909,I72897,I72900,I72891,I72888,I72891,I72903,I72906,I72958,I72961,I72964,I72967,I72970,I72973,I72976,I72979,I72982,I72985,I2224,I2231);
PAT_13 I_1001 (I72964,I72973,I72958,I72961,I72982,I72967,I72979,I72958,I72976,I72985,I72970,I73031,I73034,I73037,I73040,I73043,I73046,I73049,I73052,I73055,I2224,I2231);
PAT_5 I_1002 (I73043,I73034,I73040,I73052,I73034,I73055,I73037,I73046,I73031,I73031,I73049,I73101,I73104,I73107,I73110,I73113,I73116,I73119,I73122,I73125,I73128,I2224,I2231);
PAT_8 I_1003 (I73101,I73128,I73119,I73116,I73110,I73101,I73113,I73125,I73104,I73122,I73107,I73174,I73177,I73180,I73183,I73186,I73189,I73192,I73195,I73198,I2224,I2231);
PAT_12 I_1004 (I73174,I73177,I73177,I73198,I73183,I73192,I73195,I73186,I73180,I73189,I73174,I73244,I73247,I73250,I73253,I73256,I73259,I73262,I73265,I2224,I2231);
PAT_16 I_1005 (I73253,I73247,I73250,I73244,I73244,I73250,I73265,I73262,I73247,I73256,I73259,I73311,I73314,I73317,I73320,I73323,I73326,I73329,I73332,I73335,I73338,I2224,I2231);
PAT_15 I_1006 (I73335,I73311,I73332,I73326,I73317,I73320,I73311,I73314,I73338,I73329,I73323,I73384,I73387,I73390,I73393,I73396,I73399,I73402,I73405,I73408,I2224,I2231);
PAT_9 I_1007 (I73384,I73405,I73393,I73387,I73399,I73387,I73402,I73408,I73390,I73384,I73396,I73454,I73457,I73460,I73463,I73466,I73469,I73472,I73475,I73478,I2224,I2231);
PAT_2 I_1008 (I73469,I73472,I73463,I73478,I73454,I73457,I73460,I73457,I73475,I73466,I73454,I73524,I73527,I73530,I73533,I73536,I73539,I73542,I73545,I73548,I2224,I2231);
PAT_9 I_1009 (I73539,I73548,I73524,I73530,I73533,I73542,I73527,I73536,I73545,I73527,I73524,I73594,I73597,I73600,I73603,I73606,I73609,I73612,I73615,I73618,I2224,I2231);
PAT_4 I_1010 (I73594,I73618,I73612,I73600,I73597,I73615,I73597,I73594,I73609,I73603,I73606,I73664,I73667,I73670,I73673,I73676,I73679,I73682,I73685,I73688,I2224,I2231);
PAT_11 I_1011 (I73676,I73685,I73667,I73679,I73664,I73667,I73664,I73673,I73688,I73682,I73670,I73734,I73737,I73740,I73743,I73746,I73749,I73752,I73755,I73758,I73761,I2224,I2231);
PAT_10 I_1012 (I73749,I73755,I73746,I73740,I73758,I73743,I73761,I73752,I73734,I73737,I73734,I73807,I73810,I73813,I73816,I73819,I73822,I73825,I73828,I2224,I2231);
PAT_14 I_1013 (I73807,I73828,I73813,I73822,I73819,I73825,I73816,I73810,I73810,I73813,I73807,I73874,I73877,I73880,I73883,I73886,I73889,I73892,I73895,I73898,I2224,I2231);
PAT_2 I_1014 (I73892,I73898,I73883,I73874,I73877,I73877,I73889,I73874,I73895,I73880,I73886,I73944,I73947,I73950,I73953,I73956,I73959,I73962,I73965,I73968,I2224,I2231);
PAT_13 I_1015 (I73953,I73947,I73944,I73965,I73956,I73959,I73947,I73950,I73962,I73968,I73944,I74014,I74017,I74020,I74023,I74026,I74029,I74032,I74035,I74038,I2224,I2231);
PAT_7 I_1016 (I74023,I74026,I74014,I74029,I74035,I74020,I74017,I74038,I74017,I74014,I74032,I74084,I74087,I74090,I74093,I74096,I74099,I74102,I74105,I74108,I2224,I2231);
PAT_11 I_1017 (I74096,I74090,I74084,I74105,I74108,I74093,I74087,I74102,I74084,I74099,I74087,I74154,I74157,I74160,I74163,I74166,I74169,I74172,I74175,I74178,I74181,I2224,I2231);
PAT_10 I_1018 (I74169,I74175,I74166,I74160,I74178,I74163,I74181,I74172,I74154,I74157,I74154,I74227,I74230,I74233,I74236,I74239,I74242,I74245,I74248,I2224,I2231);
PAT_13 I_1019 (I74233,I74239,I74233,I74230,I74245,I74248,I74227,I74227,I74242,I74230,I74236,I74294,I74297,I74300,I74303,I74306,I74309,I74312,I74315,I74318,I2224,I2231);
PAT_11 I_1020 (I74294,I74306,I74309,I74300,I74297,I74318,I74297,I74315,I74303,I74294,I74312,I74364,I74367,I74370,I74373,I74376,I74379,I74382,I74385,I74388,I74391,I2224,I2231);
PAT_1 I_1021 (I74379,I74370,I74373,I74364,I74385,I74382,I74367,I74364,I74391,I74388,I74376,I74437,I74440,I74443,I74446,I74449,I74452,I74455,I74458,I74461,I2224,I2231);
PAT_8 I_1022 (I74458,I74440,I74446,I74437,I74455,I74449,I74452,I74437,I74461,I74443,I74440,I74507,I74510,I74513,I74516,I74519,I74522,I74525,I74528,I74531,I2224,I2231);
PAT_6 I_1023 (I74510,I74507,I74513,I74525,I74522,I74516,I74519,I74507,I74528,I74510,I74531,I74577,I74580,I74583,I74586,I74589,I74592,I74595,I74598,I74601,I74604,I2224,I2231);
PAT_11 I_1024 (I74577,I74592,I74577,I74589,I74586,I74604,I74601,I74598,I74595,I74580,I74583,I74650,I74653,I74656,I74659,I74662,I74665,I74668,I74671,I74674,I74677,I2224,I2231);
PAT_9 I_1025 (I74656,I74668,I74659,I74671,I74650,I74653,I74662,I74650,I74665,I74674,I74677,I74723,I74726,I74729,I74732,I74735,I74738,I74741,I74744,I74747,I2224,I2231);
PAT_8 I_1026 (I74744,I74732,I74741,I74723,I74726,I74738,I74747,I74726,I74729,I74735,I74723,I74793,I74796,I74799,I74802,I74805,I74808,I74811,I74814,I74817,I2224,I2231);
PAT_17 I_1027 (I74817,I74805,I74802,I74796,I74799,I74811,I74793,I74796,I74793,I74808,I74814,I74863,I74866,I74869,I74872,I74875,I74878,I74881,I74884,I74887,I74890,I2224,I2231);
PAT_9 I_1028 (I74884,I74866,I74872,I74887,I74869,I74881,I74863,I74875,I74863,I74890,I74878,I74936,I74939,I74942,I74945,I74948,I74951,I74954,I74957,I74960,I2224,I2231);
PAT_17 I_1029 (I74939,I74945,I74960,I74951,I74954,I74942,I74936,I74948,I74936,I74939,I74957,I75006,I75009,I75012,I75015,I75018,I75021,I75024,I75027,I75030,I75033,I2224,I2231);
PAT_3 I_1030 (I75018,I75021,I75024,I75027,I75006,I75006,I75012,I75030,I75033,I75015,I75009,I75079,I75082,I75085,I75088,I75091,I75094,I75097,I75100,I75103,I75106,I2224,I2231);
PAT_9 I_1031 (I75079,I75103,I75085,I75100,I75088,I75082,I75097,I75106,I75079,I75091,I75094,I75152,I75155,I75158,I75161,I75164,I75167,I75170,I75173,I75176,I2224,I2231);
PAT_14 I_1032 (I75161,I75152,I75176,I75158,I75155,I75152,I75167,I75173,I75164,I75155,I75170,I75222,I75225,I75228,I75231,I75234,I75237,I75240,I75243,I75246,I2224,I2231);
PAT_9 I_1033 (I75231,I75243,I75222,I75240,I75225,I75228,I75246,I75225,I75234,I75222,I75237,I75292,I75295,I75298,I75301,I75304,I75307,I75310,I75313,I75316,I2224,I2231);
PAT_5 I_1034 (I75313,I75292,I75307,I75292,I75298,I75301,I75295,I75295,I75310,I75304,I75316,I75362,I75365,I75368,I75371,I75374,I75377,I75380,I75383,I75386,I75389,I2224,I2231);
PAT_13 I_1035 (I75368,I75377,I75362,I75365,I75386,I75371,I75383,I75362,I75380,I75389,I75374,I75435,I75438,I75441,I75444,I75447,I75450,I75453,I75456,I75459,I2224,I2231);
PAT_11 I_1036 (I75435,I75447,I75450,I75441,I75438,I75459,I75438,I75456,I75444,I75435,I75453,I75505,I75508,I75511,I75514,I75517,I75520,I75523,I75526,I75529,I75532,I2224,I2231);
PAT_9 I_1037 (I75511,I75523,I75514,I75526,I75505,I75508,I75517,I75505,I75520,I75529,I75532,I75578,I75581,I75584,I75587,I75590,I75593,I75596,I75599,I75602,I2224,I2231);
PAT_1 I_1038 (I75578,I75596,I75578,I75590,I75581,I75587,I75593,I75599,I75602,I75584,I75581,I75648,I75651,I75654,I75657,I75660,I75663,I75666,I75669,I75672,I2224,I2231);
PAT_16 I_1039 (I75669,I75672,I75663,I75648,I75666,I75648,I75651,I75657,I75651,I75660,I75654,I75718,I75721,I75724,I75727,I75730,I75733,I75736,I75739,I75742,I75745,I2224,I2231);
PAT_12 I_1040 (I75721,I75718,I75736,I75718,I75745,I75742,I75730,I75727,I75733,I75724,I75739,I75791,I75794,I75797,I75800,I75803,I75806,I75809,I75812,I2224,I2231);
PAT_2 I_1041 (I75809,I75803,I75812,I75806,I75800,I75797,I75791,I75791,I75797,I75794,I75794,I75858,I75861,I75864,I75867,I75870,I75873,I75876,I75879,I75882,I2224,I2231);
PAT_10 I_1042 (I75858,I75876,I75873,I75861,I75864,I75879,I75870,I75858,I75867,I75882,I75861,I75928,I75931,I75934,I75937,I75940,I75943,I75946,I75949,I2224,I2231);
PAT_9 I_1043 (I75940,I75928,I75931,I75934,I75928,I75934,I75937,I75931,I75949,I75943,I75946,I75995,I75998,I76001,I76004,I76007,I76010,I76013,I76016,I76019,I2224,I2231);
PAT_11 I_1044 (I76007,I76013,I76019,I76016,I76004,I75998,I75998,I75995,I76010,I75995,I76001,I76065,I76068,I76071,I76074,I76077,I76080,I76083,I76086,I76089,I76092,I2224,I2231);
PAT_9 I_1045 (I76071,I76083,I76074,I76086,I76065,I76068,I76077,I76065,I76080,I76089,I76092,I76138,I76141,I76144,I76147,I76150,I76153,I76156,I76159,I76162,I2224,I2231);
PAT_10 I_1046 (I76159,I76156,I76144,I76141,I76162,I76147,I76153,I76141,I76138,I76138,I76150,I76208,I76211,I76214,I76217,I76220,I76223,I76226,I76229,I2224,I2231);
PAT_13 I_1047 (I76214,I76220,I76214,I76211,I76226,I76229,I76208,I76208,I76223,I76211,I76217,I76275,I76278,I76281,I76284,I76287,I76290,I76293,I76296,I76299,I2224,I2231);
PAT_17 I_1048 (I76299,I76287,I76296,I76293,I76284,I76275,I76278,I76281,I76275,I76290,I76278,I76345,I76348,I76351,I76354,I76357,I76360,I76363,I76366,I76369,I76372,I2224,I2231);
PAT_4 I_1049 (I76354,I76345,I76363,I76360,I76372,I76369,I76348,I76345,I76351,I76357,I76366,I76418,I76421,I76424,I76427,I76430,I76433,I76436,I76439,I76442,I2224,I2231);
PAT_11 I_1050 (I76430,I76439,I76421,I76433,I76418,I76421,I76418,I76427,I76442,I76436,I76424,I76488,I76491,I76494,I76497,I76500,I76503,I76506,I76509,I76512,I76515,I2224,I2231);
PAT_2 I_1051 (I76488,I76512,I76500,I76494,I76503,I76506,I76491,I76515,I76509,I76497,I76488,I76561,I76564,I76567,I76570,I76573,I76576,I76579,I76582,I76585,I2224,I2231);
PAT_17 I_1052 (I76561,I76561,I76573,I76564,I76567,I76579,I76576,I76585,I76564,I76570,I76582,I76631,I76634,I76637,I76640,I76643,I76646,I76649,I76652,I76655,I76658,I2224,I2231);
PAT_5 I_1053 (I76643,I76637,I76634,I76655,I76640,I76646,I76649,I76631,I76631,I76652,I76658,I76704,I76707,I76710,I76713,I76716,I76719,I76722,I76725,I76728,I76731,I2224,I2231);
PAT_13 I_1054 (I76710,I76719,I76704,I76707,I76728,I76713,I76725,I76704,I76722,I76731,I76716,I76777,I76780,I76783,I76786,I76789,I76792,I76795,I76798,I76801,I2224,I2231);
PAT_5 I_1055 (I76789,I76780,I76786,I76798,I76780,I76801,I76783,I76792,I76777,I76777,I76795,I76847,I76850,I76853,I76856,I76859,I76862,I76865,I76868,I76871,I76874,I2224,I2231);
PAT_13 I_1056 (I76853,I76862,I76847,I76850,I76871,I76856,I76868,I76847,I76865,I76874,I76859,I76920,I76923,I76926,I76929,I76932,I76935,I76938,I76941,I76944,I2224,I2231);
PAT_5 I_1057 (I76932,I76923,I76929,I76941,I76923,I76944,I76926,I76935,I76920,I76920,I76938,I76990,I76993,I76996,I76999,I77002,I77005,I77008,I77011,I77014,I77017,I2224,I2231);
PAT_1 I_1058 (I77005,I76993,I77011,I76990,I76996,I76990,I76999,I77014,I77008,I77017,I77002,I77063,I77066,I77069,I77072,I77075,I77078,I77081,I77084,I77087,I2224,I2231);
PAT_5 I_1059 (I77081,I77084,I77066,I77075,I77072,I77069,I77078,I77087,I77066,I77063,I77063,I77133,I77136,I77139,I77142,I77145,I77148,I77151,I77154,I77157,I77160,I2224,I2231);
PAT_2 I_1060 (I77148,I77133,I77145,I77139,I77154,I77136,I77151,I77142,I77157,I77160,I77133,I77206,I77209,I77212,I77215,I77218,I77221,I77224,I77227,I77230,I2224,I2231);
PAT_5 I_1061 (I77227,I77206,I77206,I77218,I77215,I77224,I77212,I77221,I77230,I77209,I77209,I77276,I77279,I77282,I77285,I77288,I77291,I77294,I77297,I77300,I77303,I2224,I2231);
PAT_13 I_1062 (I77282,I77291,I77276,I77279,I77300,I77285,I77297,I77276,I77294,I77303,I77288,I77349,I77352,I77355,I77358,I77361,I77364,I77367,I77370,I77373,I2224,I2231);
PAT_5 I_1063 (I77361,I77352,I77358,I77370,I77352,I77373,I77355,I77364,I77349,I77349,I77367,I77419,I77422,I77425,I77428,I77431,I77434,I77437,I77440,I77443,I77446,I2224,I2231);
PAT_10 I_1064 (I77443,I77446,I77425,I77431,I77434,I77440,I77422,I77419,I77419,I77428,I77437,I77492,I77495,I77498,I77501,I77504,I77507,I77510,I77513,I2224,I2231);
PAT_9 I_1065 (I77504,I77492,I77495,I77498,I77492,I77498,I77501,I77495,I77513,I77507,I77510,I77559,I77562,I77565,I77568,I77571,I77574,I77577,I77580,I77583,I2224,I2231);
PAT_10 I_1066 (I77580,I77577,I77565,I77562,I77583,I77568,I77574,I77562,I77559,I77559,I77571,I77629,I77632,I77635,I77638,I77641,I77644,I77647,I77650,I2224,I2231);
PAT_17 I_1067 (I77641,I77650,I77644,I77629,I77635,I77647,I77632,I77632,I77629,I77635,I77638,I77696,I77699,I77702,I77705,I77708,I77711,I77714,I77717,I77720,I77723,I2224,I2231);
PAT_11 I_1068 (I77708,I77717,I77723,I77699,I77696,I77714,I77705,I77711,I77702,I77720,I77696,I77769,I77772,I77775,I77778,I77781,I77784,I77787,I77790,I77793,I77796,I2224,I2231);
PAT_9 I_1069 (I77775,I77787,I77778,I77790,I77769,I77772,I77781,I77769,I77784,I77793,I77796,I77842,I77845,I77848,I77851,I77854,I77857,I77860,I77863,I77866,I2224,I2231);
PAT_5 I_1070 (I77863,I77842,I77857,I77842,I77848,I77851,I77845,I77845,I77860,I77854,I77866,I77912,I77915,I77918,I77921,I77924,I77927,I77930,I77933,I77936,I77939,I2224,I2231);
PAT_13 I_1071 (I77918,I77927,I77912,I77915,I77936,I77921,I77933,I77912,I77930,I77939,I77924,I77985,I77988,I77991,I77994,I77997,I78000,I78003,I78006,I78009,I2224,I2231);
PAT_5 I_1072 (I77997,I77988,I77994,I78006,I77988,I78009,I77991,I78000,I77985,I77985,I78003,I78055,I78058,I78061,I78064,I78067,I78070,I78073,I78076,I78079,I78082,I2224,I2231);
PAT_10 I_1073 (I78079,I78082,I78061,I78067,I78070,I78076,I78058,I78055,I78055,I78064,I78073,I78128,I78131,I78134,I78137,I78140,I78143,I78146,I78149,I2224,I2231);
PAT_11 I_1074 (I78137,I78140,I78149,I78143,I78146,I78128,I78128,I78134,I78131,I78131,I78134,I78195,I78198,I78201,I78204,I78207,I78210,I78213,I78216,I78219,I78222,I2224,I2231);
PAT_4 I_1075 (I78201,I78222,I78195,I78213,I78204,I78195,I78216,I78198,I78207,I78219,I78210,I78268,I78271,I78274,I78277,I78280,I78283,I78286,I78289,I78292,I2224,I2231);
PAT_10 I_1076 (I78268,I78268,I78292,I78271,I78277,I78286,I78283,I78271,I78289,I78274,I78280,I78338,I78341,I78344,I78347,I78350,I78353,I78356,I78359,I2224,I2231);
PAT_13 I_1077 (I78344,I78350,I78344,I78341,I78356,I78359,I78338,I78338,I78353,I78341,I78347,I78405,I78408,I78411,I78414,I78417,I78420,I78423,I78426,I78429,I2224,I2231);
PAT_12 I_1078 (I78414,I78405,I78405,I78429,I78426,I78408,I78423,I78417,I78408,I78411,I78420,I78475,I78478,I78481,I78484,I78487,I78490,I78493,I78496,I2224,I2231);
PAT_16 I_1079 (I78484,I78478,I78481,I78475,I78475,I78481,I78496,I78493,I78478,I78487,I78490,I78542,I78545,I78548,I78551,I78554,I78557,I78560,I78563,I78566,I78569,I2224,I2231);
PAT_13 I_1080 (I78554,I78545,I78542,I78548,I78557,I78566,I78563,I78560,I78551,I78542,I78569,I78615,I78618,I78621,I78624,I78627,I78630,I78633,I78636,I78639,I2224,I2231);
PAT_8 I_1081 (I78624,I78636,I78627,I78630,I78639,I78618,I78633,I78615,I78618,I78621,I78615,I78685,I78688,I78691,I78694,I78697,I78700,I78703,I78706,I78709,I2224,I2231);
PAT_6 I_1082 (I78688,I78685,I78691,I78703,I78700,I78694,I78697,I78685,I78706,I78688,I78709,I78755,I78758,I78761,I78764,I78767,I78770,I78773,I78776,I78779,I78782,I2224,I2231);
PAT_13 I_1083 (I78779,I78761,I78776,I78755,I78758,I78764,I78782,I78767,I78773,I78755,I78770,I78828,I78831,I78834,I78837,I78840,I78843,I78846,I78849,I78852,I2224,I2231);
PAT_9 I_1084 (I78849,I78831,I78831,I78828,I78852,I78834,I78837,I78828,I78840,I78846,I78843,I78898,I78901,I78904,I78907,I78910,I78913,I78916,I78919,I78922,I2224,I2231);
PAT_13 I_1085 (I78898,I78919,I78901,I78916,I78910,I78907,I78922,I78898,I78904,I78913,I78901,I78968,I78971,I78974,I78977,I78980,I78983,I78986,I78989,I78992,I2224,I2231);
PAT_7 I_1086 (I78977,I78980,I78968,I78983,I78989,I78974,I78971,I78992,I78971,I78968,I78986,I79038,I79041,I79044,I79047,I79050,I79053,I79056,I79059,I79062,I2224,I2231);
PAT_6 I_1087 (I79038,I79056,I79038,I79047,I79053,I79041,I79059,I79044,I79062,I79041,I79050,I79108,I79111,I79114,I79117,I79120,I79123,I79126,I79129,I79132,I79135,I2224,I2231);
PAT_5 I_1088 (I79129,I79108,I79114,I79117,I79123,I79126,I79108,I79132,I79111,I79120,I79135,I79181,I79184,I79187,I79190,I79193,I79196,I79199,I79202,I79205,I79208,I2224,I2231);
PAT_1 I_1089 (I79196,I79184,I79202,I79181,I79187,I79181,I79190,I79205,I79199,I79208,I79193,I79254,I79257,I79260,I79263,I79266,I79269,I79272,I79275,I79278,I2224,I2231);
PAT_9 I_1090 (I79269,I79275,I79260,I79278,I79257,I79272,I79257,I79263,I79254,I79266,I79254,I79324,I79327,I79330,I79333,I79336,I79339,I79342,I79345,I79348,I2224,I2231);
PAT_17 I_1091 (I79327,I79333,I79348,I79339,I79342,I79330,I79324,I79336,I79324,I79327,I79345,I79394,I79397,I79400,I79403,I79406,I79409,I79412,I79415,I79418,I79421,I2224,I2231);
PAT_13 I_1092 (I79412,I79415,I79400,I79394,I79406,I79418,I79397,I79409,I79394,I79421,I79403,I79467,I79470,I79473,I79476,I79479,I79482,I79485,I79488,I79491,I2224,I2231);
PAT_4 I_1093 (I79476,I79479,I79491,I79473,I79488,I79485,I79470,I79482,I79470,I79467,I79467,I79537,I79540,I79543,I79546,I79549,I79552,I79555,I79558,I79561,I2224,I2231);
PAT_9 I_1094 (I79558,I79540,I79543,I79552,I79555,I79537,I79546,I79540,I79561,I79537,I79549,I79607,I79610,I79613,I79616,I79619,I79622,I79625,I79628,I79631,I2224,I2231);
PAT_10 I_1095 (I79628,I79625,I79613,I79610,I79631,I79616,I79622,I79610,I79607,I79607,I79619,I79677,I79680,I79683,I79686,I79689,I79692,I79695,I79698,I2224,I2231);
PAT_6 I_1096 (I79698,I79692,I79686,I79680,I79677,I79683,I79677,I79683,I79680,I79689,I79695,I79744,I79747,I79750,I79753,I79756,I79759,I79762,I79765,I79768,I79771,I2224,I2231);
PAT_8 I_1097 (I79753,I79759,I79750,I79762,I79744,I79747,I79765,I79744,I79771,I79768,I79756,I79817,I79820,I79823,I79826,I79829,I79832,I79835,I79838,I79841,I2224,I2231);
PAT_17 I_1098 (I79841,I79829,I79826,I79820,I79823,I79835,I79817,I79820,I79817,I79832,I79838,I79887,I79890,I79893,I79896,I79899,I79902,I79905,I79908,I79911,I79914,I2224,I2231);
PAT_11 I_1099 (I79899,I79908,I79914,I79890,I79887,I79905,I79896,I79902,I79893,I79911,I79887,I79960,I79963,I79966,I79969,I79972,I79975,I79978,I79981,I79984,I79987,I2224,I2231);
PAT_4 I_1100 (I79966,I79987,I79960,I79978,I79969,I79960,I79981,I79963,I79972,I79984,I79975,I80033,I80036,I80039,I80042,I80045,I80048,I80051,I80054,I80057,I2224,I2231);
PAT_17 I_1101 (I80045,I80042,I80054,I80048,I80033,I80051,I80057,I80036,I80039,I80036,I80033,I80103,I80106,I80109,I80112,I80115,I80118,I80121,I80124,I80127,I80130,I2224,I2231);
PAT_14 I_1102 (I80106,I80121,I80103,I80127,I80112,I80118,I80103,I80124,I80109,I80130,I80115,I80176,I80179,I80182,I80185,I80188,I80191,I80194,I80197,I80200,I2224,I2231);
PAT_17 I_1103 (I80191,I80179,I80200,I80176,I80197,I80185,I80182,I80194,I80188,I80179,I80176,I80246,I80249,I80252,I80255,I80258,I80261,I80264,I80267,I80270,I80273,I2224,I2231);
PAT_6 I_1104 (I80246,I80264,I80252,I80255,I80261,I80246,I80258,I80249,I80270,I80273,I80267,I80319,I80322,I80325,I80328,I80331,I80334,I80337,I80340,I80343,I80346,I2224,I2231);
PAT_13 I_1105 (I80343,I80325,I80340,I80319,I80322,I80328,I80346,I80331,I80337,I80319,I80334,I80392,I80395,I80398,I80401,I80404,I80407,I80410,I80413,I80416,I2224,I2231);
PAT_17 I_1106 (I80416,I80404,I80413,I80410,I80401,I80392,I80395,I80398,I80392,I80407,I80395,I80462,I80465,I80468,I80471,I80474,I80477,I80480,I80483,I80486,I80489,I2224,I2231);
PAT_2 I_1107 (I80462,I80480,I80477,I80462,I80471,I80486,I80483,I80468,I80489,I80474,I80465,I80535,I80538,I80541,I80544,I80547,I80550,I80553,I80556,I80559,I2224,I2231);
PAT_13 I_1108 (I80544,I80538,I80535,I80556,I80547,I80550,I80538,I80541,I80553,I80559,I80535,I80605,I80608,I80611,I80614,I80617,I80620,I80623,I80626,I80629,I2224,I2231);
PAT_6 I_1109 (I80605,I80617,I80614,I80626,I80623,I80629,I80605,I80620,I80608,I80608,I80611,I80675,I80678,I80681,I80684,I80687,I80690,I80693,I80696,I80699,I80702,I2224,I2231);
PAT_10 I_1110 (I80675,I80690,I80693,I80684,I80675,I80699,I80702,I80678,I80687,I80681,I80696,I80748,I80751,I80754,I80757,I80760,I80763,I80766,I80769,I2224,I2231);
PAT_13 I_1111 (I80754,I80760,I80754,I80751,I80766,I80769,I80748,I80748,I80763,I80751,I80757,I80815,I80818,I80821,I80824,I80827,I80830,I80833,I80836,I80839,I2224,I2231);
PAT_11 I_1112 (I80815,I80827,I80830,I80821,I80818,I80839,I80818,I80836,I80824,I80815,I80833,I80885,I80888,I80891,I80894,I80897,I80900,I80903,I80906,I80909,I80912,I2224,I2231);
PAT_5 I_1113 (I80906,I80885,I80912,I80900,I80897,I80909,I80891,I80885,I80903,I80888,I80894,I80958,I80961,I80964,I80967,I80970,I80973,I80976,I80979,I80982,I80985,I2224,I2231);
PAT_4 I_1114 (I80976,I80982,I80985,I80964,I80967,I80979,I80961,I80958,I80970,I80973,I80958,I81031,I81034,I81037,I81040,I81043,I81046,I81049,I81052,I81055,I2224,I2231);
PAT_13 I_1115 (I81046,I81040,I81052,I81037,I81043,I81031,I81055,I81049,I81034,I81031,I81034,I81101,I81104,I81107,I81110,I81113,I81116,I81119,I81122,I81125,I2224,I2231);
PAT_4 I_1116 (I1473,I2041,I1569,I1441,I1393,I1777,I1537,I1881,I1737,I1729,I1809,I81171,I81174,I81177,I81180,I81183,I81186,I81189,I81192,I81195,I2224,I2231);
PAT_6 I_1117 (I81171,I81177,I81174,I81186,I81189,I81183,I81195,I81192,I81171,I81180,I81174,I81241,I81244,I81247,I81250,I81253,I81256,I81259,I81262,I81265,I81268,I2224,I2231);
PAT_5 I_1118 (I81262,I81241,I81247,I81250,I81256,I81259,I81241,I81265,I81244,I81253,I81268,I81314,I81317,I81320,I81323,I81326,I81329,I81332,I81335,I81338,I81341,I2224,I2231);
PAT_10 I_1119 (I81338,I81341,I81320,I81326,I81329,I81335,I81317,I81314,I81314,I81323,I81332,I81387,I81390,I81393,I81396,I81399,I81402,I81405,I81408,I2224,I2231);
PAT_13 I_1120 (I81393,I81399,I81393,I81390,I81405,I81408,I81387,I81387,I81402,I81390,I81396,I81454,I81457,I81460,I81463,I81466,I81469,I81472,I81475,I81478,I2224,I2231);
PAT_8 I_1121 (I81463,I81475,I81466,I81469,I81478,I81457,I81472,I81454,I81457,I81460,I81454,I81524,I81527,I81530,I81533,I81536,I81539,I81542,I81545,I81548,I2224,I2231);
PAT_11 I_1122 (I81545,I81536,I81524,I81527,I81542,I81530,I81533,I81524,I81548,I81539,I81527,I81594,I81597,I81600,I81603,I81606,I81609,I81612,I81615,I81618,I81621,I2224,I2231);
PAT_8 I_1123 (I81603,I81609,I81612,I81618,I81615,I81606,I81594,I81594,I81621,I81597,I81600,I81667,I81670,I81673,I81676,I81679,I81682,I81685,I81688,I81691,I2224,I2231);
PAT_5 I_1124 (I81673,I81691,I81667,I81688,I81676,I81679,I81670,I81667,I81670,I81682,I81685,I81737,I81740,I81743,I81746,I81749,I81752,I81755,I81758,I81761,I81764,I2224,I2231);
PAT_9 I_1125 (I81752,I81749,I81758,I81755,I81746,I81737,I81743,I81764,I81740,I81761,I81737,I81810,I81813,I81816,I81819,I81822,I81825,I81828,I81831,I81834,I2224,I2231);
PAT_14 I_1126 (I81819,I81810,I81834,I81816,I81813,I81810,I81825,I81831,I81822,I81813,I81828,I81880,I81883,I81886,I81889,I81892,I81895,I81898,I81901,I81904,I2224,I2231);
PAT_11 I_1127 (I81892,I81889,I81886,I81880,I81883,I81883,I81895,I81880,I81901,I81904,I81898,I81950,I81953,I81956,I81959,I81962,I81965,I81968,I81971,I81974,I81977,I2224,I2231);
PAT_9 I_1128 (I81956,I81968,I81959,I81971,I81950,I81953,I81962,I81950,I81965,I81974,I81977,I82023,I82026,I82029,I82032,I82035,I82038,I82041,I82044,I82047,I2224,I2231);
PAT_10 I_1129 (I82044,I82041,I82029,I82026,I82047,I82032,I82038,I82026,I82023,I82023,I82035,I82093,I82096,I82099,I82102,I82105,I82108,I82111,I82114,I2224,I2231);
PAT_2 I_1130 (I82105,I82108,I82099,I82111,I82096,I82093,I82093,I82099,I82114,I82102,I82096,I82160,I82163,I82166,I82169,I82172,I82175,I82178,I82181,I82184,I2224,I2231);
PAT_8 I_1131 (I82172,I82163,I82169,I82160,I82166,I82181,I82178,I82160,I82175,I82163,I82184,I82230,I82233,I82236,I82239,I82242,I82245,I82248,I82251,I82254,I2224,I2231);
PAT_9 I_1132 (I82233,I82242,I82233,I82230,I82245,I82236,I82251,I82239,I82248,I82230,I82254,I82300,I82303,I82306,I82309,I82312,I82315,I82318,I82321,I82324,I2224,I2231);
PAT_2 I_1133 (I82315,I82318,I82309,I82324,I82300,I82303,I82306,I82303,I82321,I82312,I82300,I82370,I82373,I82376,I82379,I82382,I82385,I82388,I82391,I82394,I2224,I2231);
PAT_8 I_1134 (I82382,I82373,I82379,I82370,I82376,I82391,I82388,I82370,I82385,I82373,I82394,I82440,I82443,I82446,I82449,I82452,I82455,I82458,I82461,I82464,I2224,I2231);
PAT_13 I_1135 (I82452,I82461,I82443,I82464,I82446,I82440,I82440,I82449,I82458,I82455,I82443,I82510,I82513,I82516,I82519,I82522,I82525,I82528,I82531,I82534,I2224,I2231);
PAT_8 I_1136 (I82519,I82531,I82522,I82525,I82534,I82513,I82528,I82510,I82513,I82516,I82510,I82580,I82583,I82586,I82589,I82592,I82595,I82598,I82601,I82604,I2224,I2231);
PAT_13 I_1137 (I82592,I82601,I82583,I82604,I82586,I82580,I82580,I82589,I82598,I82595,I82583,I82650,I82653,I82656,I82659,I82662,I82665,I82668,I82671,I82674,I2224,I2231);
PAT_9 I_1138 (I82671,I82653,I82653,I82650,I82674,I82656,I82659,I82650,I82662,I82668,I82665,I82720,I82723,I82726,I82729,I82732,I82735,I82738,I82741,I82744,I2224,I2231);
PAT_8 I_1139 (I82741,I82729,I82738,I82720,I82723,I82735,I82744,I82723,I82726,I82732,I82720,I82790,I82793,I82796,I82799,I82802,I82805,I82808,I82811,I82814,I2224,I2231);
PAT_16 I_1140 (I82811,I82790,I82790,I82799,I82796,I82808,I82793,I82802,I82805,I82814,I82793,I82860,I82863,I82866,I82869,I82872,I82875,I82878,I82881,I82884,I82887,I2224,I2231);
PAT_2 I_1141 (I82869,I82875,I82863,I82887,I82860,I82878,I82872,I82866,I82884,I82860,I82881,I82933,I82936,I82939,I82942,I82945,I82948,I82951,I82954,I82957,I2224,I2231);
PAT_13 I_1142 (I82942,I82936,I82933,I82954,I82945,I82948,I82936,I82939,I82951,I82957,I82933,I83003,I83006,I83009,I83012,I83015,I83018,I83021,I83024,I83027,I2224,I2231);
PAT_17 I_1143 (I83027,I83015,I83024,I83021,I83012,I83003,I83006,I83009,I83003,I83018,I83006,I83073,I83076,I83079,I83082,I83085,I83088,I83091,I83094,I83097,I83100,I2224,I2231);
PAT_11 I_1144 (I83085,I83094,I83100,I83076,I83073,I83091,I83082,I83088,I83079,I83097,I83073,I83146,I83149,I83152,I83155,I83158,I83161,I83164,I83167,I83170,I83173,I2224,I2231);
PAT_1 I_1145 (I83161,I83152,I83155,I83146,I83167,I83164,I83149,I83146,I83173,I83170,I83158,I83219,I83222,I83225,I83228,I83231,I83234,I83237,I83240,I83243,I2224,I2231);
PAT_7 I_1146 (I83222,I83228,I83225,I83231,I83237,I83234,I83243,I83240,I83222,I83219,I83219,I83289,I83292,I83295,I83298,I83301,I83304,I83307,I83310,I83313,I2224,I2231);
PAT_13 I_1147 (I83295,I83313,I83304,I83289,I83301,I83289,I83310,I83292,I83298,I83292,I83307,I83359,I83362,I83365,I83368,I83371,I83374,I83377,I83380,I83383,I2224,I2231);
PAT_10 I_1148 (I83380,I83374,I83368,I83362,I83383,I83362,I83371,I83359,I83359,I83377,I83365,I83429,I83432,I83435,I83438,I83441,I83444,I83447,I83450,I2224,I2231);
PAT_4 I_1149 (I83444,I83441,I83432,I83450,I83429,I83432,I83438,I83435,I83447,I83429,I83435,I83496,I83499,I83502,I83505,I83508,I83511,I83514,I83517,I83520,I2224,I2231);
PAT_9 I_1150 (I83517,I83499,I83502,I83511,I83514,I83496,I83505,I83499,I83520,I83496,I83508,I83566,I83569,I83572,I83575,I83578,I83581,I83584,I83587,I83590,I2224,I2231);
PAT_10 I_1151 (I83587,I83584,I83572,I83569,I83590,I83575,I83581,I83569,I83566,I83566,I83578,I83636,I83639,I83642,I83645,I83648,I83651,I83654,I83657,I2224,I2231);
PAT_5 I_1152 (I83657,I83636,I83645,I83639,I83654,I83651,I83642,I83642,I83636,I83639,I83648,I83703,I83706,I83709,I83712,I83715,I83718,I83721,I83724,I83727,I83730,I2224,I2231);
PAT_4 I_1153 (I83721,I83727,I83730,I83709,I83712,I83724,I83706,I83703,I83715,I83718,I83703,I83776,I83779,I83782,I83785,I83788,I83791,I83794,I83797,I83800,I2224,I2231);
PAT_7 I_1154 (I83791,I83785,I83782,I83776,I83788,I83794,I83779,I83779,I83797,I83800,I83776,I83846,I83849,I83852,I83855,I83858,I83861,I83864,I83867,I83870,I2224,I2231);
PAT_4 I_1155 (I83870,I83846,I83846,I83861,I83855,I83849,I83849,I83864,I83867,I83852,I83858,I83916,I83919,I83922,I83925,I83928,I83931,I83934,I83937,I83940,I2224,I2231);
PAT_5 I_1156 (I83937,I83919,I83919,I83931,I83934,I83928,I83925,I83916,I83922,I83916,I83940,I83986,I83989,I83992,I83995,I83998,I84001,I84004,I84007,I84010,I84013,I2224,I2231);
PAT_14 I_1157 (I84007,I83992,I83986,I84010,I84013,I83986,I84004,I83989,I83995,I83998,I84001,I84059,I84062,I84065,I84068,I84071,I84074,I84077,I84080,I84083,I2224,I2231);
PAT_13 I_1158 (I84068,I84083,I84062,I84071,I84059,I84062,I84077,I84065,I84059,I84080,I84074,I84129,I84132,I84135,I84138,I84141,I84144,I84147,I84150,I84153,I2224,I2231);
PAT_7 I_1159 (I84138,I84141,I84129,I84144,I84150,I84135,I84132,I84153,I84132,I84129,I84147,I84199,I84202,I84205,I84208,I84211,I84214,I84217,I84220,I84223,I2224,I2231);
PAT_2 I_1160 (I84220,I84214,I84205,I84199,I84208,I84202,I84211,I84223,I84217,I84202,I84199,I84269,I84272,I84275,I84278,I84281,I84284,I84287,I84290,I84293,I2224,I2231);
PAT_1 I_1161 (I84281,I84269,I84275,I84278,I84269,I84284,I84293,I84272,I84287,I84272,I84290,I84339,I84342,I84345,I84348,I84351,I84354,I84357,I84360,I84363,I2224,I2231);
PAT_2 I_1162 (I84339,I84345,I84339,I84354,I84342,I84342,I84348,I84351,I84357,I84363,I84360,I84409,I84412,I84415,I84418,I84421,I84424,I84427,I84430,I84433,I2224,I2231);
PAT_10 I_1163 (I84409,I84427,I84424,I84412,I84415,I84430,I84421,I84409,I84418,I84433,I84412,I84479,I84482,I84485,I84488,I84491,I84494,I84497,I84500,I2224,I2231);
PAT_8 I_1164 (I84500,I84491,I84482,I84479,I84488,I84479,I84494,I84482,I84497,I84485,I84485,I84546,I84549,I84552,I84555,I84558,I84561,I84564,I84567,I84570,I2224,I2231);
PAT_0 I_1165 (I84546,I84564,I84555,I84570,I84558,I84546,I84549,I84552,I84561,I84549,I84567,I84616,I84619,I84622,I84625,I84628,I84631,I84634,I84637,I2224,I2231);
PAT_8 I_1166 (I84637,I84631,I84634,I84619,I84619,I84622,I84616,I84625,I84622,I84616,I84628,I84683,I84686,I84689,I84692,I84695,I84698,I84701,I84704,I84707,I2224,I2231);
PAT_11 I_1167 (I84704,I84695,I84683,I84686,I84701,I84689,I84692,I84683,I84707,I84698,I84686,I84753,I84756,I84759,I84762,I84765,I84768,I84771,I84774,I84777,I84780,I2224,I2231);
PAT_13 I_1168 (I84753,I84756,I84765,I84777,I84780,I84768,I84774,I84762,I84771,I84759,I84753,I84826,I84829,I84832,I84835,I84838,I84841,I84844,I84847,I84850,I2224,I2231);
PAT_8 I_1169 (I84835,I84847,I84838,I84841,I84850,I84829,I84844,I84826,I84829,I84832,I84826,I84896,I84899,I84902,I84905,I84908,I84911,I84914,I84917,I84920,I2224,I2231);
PAT_6 I_1170 (I84899,I84896,I84902,I84914,I84911,I84905,I84908,I84896,I84917,I84899,I84920,I84966,I84969,I84972,I84975,I84978,I84981,I84984,I84987,I84990,I84993,I2224,I2231);
PAT_8 I_1171 (I84975,I84981,I84972,I84984,I84966,I84969,I84987,I84966,I84993,I84990,I84978,I85039,I85042,I85045,I85048,I85051,I85054,I85057,I85060,I85063,I2224,I2231);
PAT_7 I_1172 (I85039,I85048,I85045,I85051,I85057,I85039,I85042,I85060,I85063,I85054,I85042,I85109,I85112,I85115,I85118,I85121,I85124,I85127,I85130,I85133,I2224,I2231);
PAT_8 I_1173 (I85115,I85127,I85109,I85112,I85118,I85109,I85133,I85130,I85121,I85124,I85112,I85179,I85182,I85185,I85188,I85191,I85194,I85197,I85200,I85203,I2224,I2231);
PAT_13 I_1174 (I85191,I85200,I85182,I85203,I85185,I85179,I85179,I85188,I85197,I85194,I85182,I85249,I85252,I85255,I85258,I85261,I85264,I85267,I85270,I85273,I2224,I2231);
PAT_11 I_1175 (I85249,I85261,I85264,I85255,I85252,I85273,I85252,I85270,I85258,I85249,I85267,I85319,I85322,I85325,I85328,I85331,I85334,I85337,I85340,I85343,I85346,I2224,I2231);
PAT_6 I_1176 (I85319,I85346,I85334,I85343,I85337,I85331,I85322,I85340,I85328,I85325,I85319,I85392,I85395,I85398,I85401,I85404,I85407,I85410,I85413,I85416,I85419,I2224,I2231);
PAT_13 I_1177 (I85416,I85398,I85413,I85392,I85395,I85401,I85419,I85404,I85410,I85392,I85407,I85465,I85468,I85471,I85474,I85477,I85480,I85483,I85486,I85489,I2224,I2231);
PAT_4 I_1178 (I85474,I85477,I85489,I85471,I85486,I85483,I85468,I85480,I85468,I85465,I85465,I85535,I85538,I85541,I85544,I85547,I85550,I85553,I85556,I85559,I2224,I2231);
PAT_1 I_1179 (I85535,I85556,I85553,I85538,I85550,I85535,I85538,I85559,I85544,I85541,I85547,I85605,I85608,I85611,I85614,I85617,I85620,I85623,I85626,I85629,I2224,I2231);
PAT_3 I_1180 (I85614,I85608,I85608,I85611,I85623,I85626,I85629,I85617,I85605,I85605,I85620,I85675,I85678,I85681,I85684,I85687,I85690,I85693,I85696,I85699,I85702,I2224,I2231);
PAT_13 I_1181 (I85696,I85684,I85702,I85681,I85687,I85690,I85678,I85693,I85675,I85675,I85699,I85748,I85751,I85754,I85757,I85760,I85763,I85766,I85769,I85772,I2224,I2231);
PAT_9 I_1182 (I85769,I85751,I85751,I85748,I85772,I85754,I85757,I85748,I85760,I85766,I85763,I85818,I85821,I85824,I85827,I85830,I85833,I85836,I85839,I85842,I2224,I2231);
PAT_1 I_1183 (I85818,I85836,I85818,I85830,I85821,I85827,I85833,I85839,I85842,I85824,I85821,I85888,I85891,I85894,I85897,I85900,I85903,I85906,I85909,I85912,I2224,I2231);
PAT_6 I_1184 (I85897,I85888,I85891,I85894,I85909,I85912,I85906,I85888,I85903,I85900,I85891,I85958,I85961,I85964,I85967,I85970,I85973,I85976,I85979,I85982,I85985,I2224,I2231);
PAT_14 I_1185 (I85970,I85964,I85958,I85985,I85967,I85961,I85973,I85976,I85958,I85982,I85979,I86031,I86034,I86037,I86040,I86043,I86046,I86049,I86052,I86055,I2224,I2231);
PAT_13 I_1186 (I86040,I86055,I86034,I86043,I86031,I86034,I86049,I86037,I86031,I86052,I86046,I86101,I86104,I86107,I86110,I86113,I86116,I86119,I86122,I86125,I2224,I2231);
PAT_10 I_1187 (I86122,I86116,I86110,I86104,I86125,I86104,I86113,I86101,I86101,I86119,I86107,I86171,I86174,I86177,I86180,I86183,I86186,I86189,I86192,I2224,I2231);
PAT_13 I_1188 (I86177,I86183,I86177,I86174,I86189,I86192,I86171,I86171,I86186,I86174,I86180,I86238,I86241,I86244,I86247,I86250,I86253,I86256,I86259,I86262,I2224,I2231);
PAT_9 I_1189 (I86259,I86241,I86241,I86238,I86262,I86244,I86247,I86238,I86250,I86256,I86253,I86308,I86311,I86314,I86317,I86320,I86323,I86326,I86329,I86332,I2224,I2231);
PAT_4 I_1190 (I86308,I86332,I86326,I86314,I86311,I86329,I86311,I86308,I86323,I86317,I86320,I86378,I86381,I86384,I86387,I86390,I86393,I86396,I86399,I86402,I2224,I2231);
PAT_2 I_1191 (I86387,I86381,I86381,I86402,I86378,I86396,I86393,I86384,I86378,I86390,I86399,I86448,I86451,I86454,I86457,I86460,I86463,I86466,I86469,I86472,I2224,I2231);
PAT_10 I_1192 (I86448,I86466,I86463,I86451,I86454,I86469,I86460,I86448,I86457,I86472,I86451,I86518,I86521,I86524,I86527,I86530,I86533,I86536,I86539,I2224,I2231);
PAT_8 I_1193 (I86539,I86530,I86521,I86518,I86527,I86518,I86533,I86521,I86536,I86524,I86524,I86585,I86588,I86591,I86594,I86597,I86600,I86603,I86606,I86609,I2224,I2231);
PAT_12 I_1194 (I86585,I86588,I86588,I86609,I86594,I86603,I86606,I86597,I86591,I86600,I86585,I86655,I86658,I86661,I86664,I86667,I86670,I86673,I86676,I2224,I2231);
PAT_4 I_1195 (I86661,I86658,I86673,I86676,I86670,I86664,I86655,I86655,I86661,I86667,I86658,I86722,I86725,I86728,I86731,I86734,I86737,I86740,I86743,I86746,I2224,I2231);
PAT_10 I_1196 (I86722,I86722,I86746,I86725,I86731,I86740,I86737,I86725,I86743,I86728,I86734,I86792,I86795,I86798,I86801,I86804,I86807,I86810,I86813,I2224,I2231);
PAT_5 I_1197 (I86813,I86792,I86801,I86795,I86810,I86807,I86798,I86798,I86792,I86795,I86804,I86859,I86862,I86865,I86868,I86871,I86874,I86877,I86880,I86883,I86886,I2224,I2231);
PAT_6 I_1198 (I86877,I86871,I86859,I86865,I86862,I86868,I86874,I86859,I86883,I86880,I86886,I86932,I86935,I86938,I86941,I86944,I86947,I86950,I86953,I86956,I86959,I2224,I2231);
PAT_10 I_1199 (I86932,I86947,I86950,I86941,I86932,I86956,I86959,I86935,I86944,I86938,I86953,I87005,I87008,I87011,I87014,I87017,I87020,I87023,I87026,I2224,I2231);
PAT_2 I_1200 (I87017,I87020,I87011,I87023,I87008,I87005,I87005,I87011,I87026,I87014,I87008,I87072,I87075,I87078,I87081,I87084,I87087,I87090,I87093,I87096,I2224,I2231);
PAT_7 I_1201 (I87096,I87072,I87078,I87075,I87075,I87084,I87087,I87072,I87090,I87093,I87081,I87142,I87145,I87148,I87151,I87154,I87157,I87160,I87163,I87166,I2224,I2231);
PAT_11 I_1202 (I87154,I87148,I87142,I87163,I87166,I87151,I87145,I87160,I87142,I87157,I87145,I87212,I87215,I87218,I87221,I87224,I87227,I87230,I87233,I87236,I87239,I2224,I2231);
PAT_9 I_1203 (I87218,I87230,I87221,I87233,I87212,I87215,I87224,I87212,I87227,I87236,I87239,I87285,I87288,I87291,I87294,I87297,I87300,I87303,I87306,I87309,I2224,I2231);
PAT_13 I_1204 (I87285,I87306,I87288,I87303,I87297,I87294,I87309,I87285,I87291,I87300,I87288,I87355,I87358,I87361,I87364,I87367,I87370,I87373,I87376,I87379,I2224,I2231);
PAT_9 I_1205 (I87376,I87358,I87358,I87355,I87379,I87361,I87364,I87355,I87367,I87373,I87370,I87425,I87428,I87431,I87434,I87437,I87440,I87443,I87446,I87449,I2224,I2231);
PAT_11 I_1206 (I87437,I87443,I87449,I87446,I87434,I87428,I87428,I87425,I87440,I87425,I87431,I87495,I87498,I87501,I87504,I87507,I87510,I87513,I87516,I87519,I87522,I2224,I2231);
PAT_10 I_1207 (I87510,I87516,I87507,I87501,I87519,I87504,I87522,I87513,I87495,I87498,I87495,I87568,I87571,I87574,I87577,I87580,I87583,I87586,I87589,I2224,I2231);
PAT_7 I_1208 (I87589,I87586,I87583,I87568,I87571,I87574,I87571,I87580,I87568,I87574,I87577,I87635,I87638,I87641,I87644,I87647,I87650,I87653,I87656,I87659,I2224,I2231);
PAT_5 I_1209 (I87641,I87635,I87644,I87653,I87647,I87659,I87656,I87638,I87650,I87638,I87635,I87705,I87708,I87711,I87714,I87717,I87720,I87723,I87726,I87729,I87732,I2224,I2231);
PAT_11 I_1210 (I87717,I87714,I87708,I87726,I87729,I87705,I87723,I87720,I87732,I87711,I87705,I87778,I87781,I87784,I87787,I87790,I87793,I87796,I87799,I87802,I87805,I2224,I2231);
PAT_2 I_1211 (I87778,I87802,I87790,I87784,I87793,I87796,I87781,I87805,I87799,I87787,I87778,I87851,I87854,I87857,I87860,I87863,I87866,I87869,I87872,I87875,I2224,I2231);
PAT_5 I_1212 (I87872,I87851,I87851,I87863,I87860,I87869,I87857,I87866,I87875,I87854,I87854,I87921,I87924,I87927,I87930,I87933,I87936,I87939,I87942,I87945,I87948,I2224,I2231);
PAT_17 I_1213 (I87948,I87924,I87927,I87930,I87921,I87933,I87921,I87945,I87939,I87936,I87942,I87994,I87997,I88000,I88003,I88006,I88009,I88012,I88015,I88018,I88021,I2224,I2231);
PAT_10 I_1214 (I87994,I88000,I88021,I88003,I88018,I87997,I88012,I88006,I88015,I88009,I87994,I88067,I88070,I88073,I88076,I88079,I88082,I88085,I88088,I2224,I2231);
PAT_8 I_1215 (I88088,I88079,I88070,I88067,I88076,I88067,I88082,I88070,I88085,I88073,I88073,I88134,I88137,I88140,I88143,I88146,I88149,I88152,I88155,I88158,I2224,I2231);
PAT_13 I_1216 (I88146,I88155,I88137,I88158,I88140,I88134,I88134,I88143,I88152,I88149,I88137,I88204,I88207,I88210,I88213,I88216,I88219,I88222,I88225,I88228,I2224,I2231);
PAT_14 I_1217 (I88207,I88222,I88210,I88219,I88213,I88204,I88216,I88225,I88204,I88228,I88207,I88274,I88277,I88280,I88283,I88286,I88289,I88292,I88295,I88298,I2224,I2231);
PAT_17 I_1218 (I88289,I88277,I88298,I88274,I88295,I88283,I88280,I88292,I88286,I88277,I88274,I88344,I88347,I88350,I88353,I88356,I88359,I88362,I88365,I88368,I88371,I2224,I2231);
PAT_2 I_1219 (I88344,I88362,I88359,I88344,I88353,I88368,I88365,I88350,I88371,I88356,I88347,I88417,I88420,I88423,I88426,I88429,I88432,I88435,I88438,I88441,I2224,I2231);
PAT_15 I_1220 (I88420,I88432,I88438,I88441,I88423,I88435,I88417,I88426,I88417,I88429,I88420,I88487,I88490,I88493,I88496,I88499,I88502,I88505,I88508,I88511,I2224,I2231);
PAT_17 I_1221 (I88487,I88487,I88499,I88490,I88493,I88511,I88508,I88502,I88490,I88496,I88505,I88557,I88560,I88563,I88566,I88569,I88572,I88575,I88578,I88581,I88584,I2224,I2231);
PAT_13 I_1222 (I88575,I88578,I88563,I88557,I88569,I88581,I88560,I88572,I88557,I88584,I88566,I88630,I88633,I88636,I88639,I88642,I88645,I88648,I88651,I88654,I2224,I2231);
PAT_9 I_1223 (I88651,I88633,I88633,I88630,I88654,I88636,I88639,I88630,I88642,I88648,I88645,I88700,I88703,I88706,I88709,I88712,I88715,I88718,I88721,I88724,I2224,I2231);
PAT_1 I_1224 (I88700,I88718,I88700,I88712,I88703,I88709,I88715,I88721,I88724,I88706,I88703,I88770,I88773,I88776,I88779,I88782,I88785,I88788,I88791,I88794,I2224,I2231);
PAT_11 I_1225 (I88773,I88788,I88785,I88791,I88794,I88773,I88779,I88782,I88770,I88776,I88770,I88840,I88843,I88846,I88849,I88852,I88855,I88858,I88861,I88864,I88867,I2224,I2231);
PAT_17 I_1226 (I88852,I88843,I88867,I88840,I88849,I88861,I88858,I88855,I88840,I88864,I88846,I88913,I88916,I88919,I88922,I88925,I88928,I88931,I88934,I88937,I88940,I2224,I2231);
PAT_13 I_1227 (I88931,I88934,I88919,I88913,I88925,I88937,I88916,I88928,I88913,I88940,I88922,I88986,I88989,I88992,I88995,I88998,I89001,I89004,I89007,I89010,I2224,I2231);
PAT_7 I_1228 (I88995,I88998,I88986,I89001,I89007,I88992,I88989,I89010,I88989,I88986,I89004,I89056,I89059,I89062,I89065,I89068,I89071,I89074,I89077,I89080,I2224,I2231);
PAT_8 I_1229 (I89062,I89074,I89056,I89059,I89065,I89056,I89080,I89077,I89068,I89071,I89059,I89126,I89129,I89132,I89135,I89138,I89141,I89144,I89147,I89150,I2224,I2231);
PAT_9 I_1230 (I89129,I89138,I89129,I89126,I89141,I89132,I89147,I89135,I89144,I89126,I89150,I89196,I89199,I89202,I89205,I89208,I89211,I89214,I89217,I89220,I2224,I2231);
PAT_14 I_1231 (I89205,I89196,I89220,I89202,I89199,I89196,I89211,I89217,I89208,I89199,I89214,I89266,I89269,I89272,I89275,I89278,I89281,I89284,I89287,I89290,I2224,I2231);
PAT_11 I_1232 (I89278,I89275,I89272,I89266,I89269,I89269,I89281,I89266,I89287,I89290,I89284,I89336,I89339,I89342,I89345,I89348,I89351,I89354,I89357,I89360,I89363,I2224,I2231);
PAT_13 I_1233 (I89336,I89339,I89348,I89360,I89363,I89351,I89357,I89345,I89354,I89342,I89336,I89409,I89412,I89415,I89418,I89421,I89424,I89427,I89430,I89433,I2224,I2231);
PAT_5 I_1234 (I89421,I89412,I89418,I89430,I89412,I89433,I89415,I89424,I89409,I89409,I89427,I89479,I89482,I89485,I89488,I89491,I89494,I89497,I89500,I89503,I89506,I2224,I2231);
PAT_9 I_1235 (I89494,I89491,I89500,I89497,I89488,I89479,I89485,I89506,I89482,I89503,I89479,I89552,I89555,I89558,I89561,I89564,I89567,I89570,I89573,I89576,I2224,I2231);
PAT_8 I_1236 (I89573,I89561,I89570,I89552,I89555,I89567,I89576,I89555,I89558,I89564,I89552,I89622,I89625,I89628,I89631,I89634,I89637,I89640,I89643,I89646,I2224,I2231);
PAT_9 I_1237 (I89625,I89634,I89625,I89622,I89637,I89628,I89643,I89631,I89640,I89622,I89646,I89692,I89695,I89698,I89701,I89704,I89707,I89710,I89713,I89716,I2224,I2231);
PAT_17 I_1238 (I89695,I89701,I89716,I89707,I89710,I89698,I89692,I89704,I89692,I89695,I89713,I89762,I89765,I89768,I89771,I89774,I89777,I89780,I89783,I89786,I89789,I2224,I2231);
PAT_8 I_1239 (I89771,I89783,I89789,I89780,I89765,I89774,I89777,I89786,I89768,I89762,I89762,I89835,I89838,I89841,I89844,I89847,I89850,I89853,I89856,I89859,I2224,I2231);
PAT_9 I_1240 (I89838,I89847,I89838,I89835,I89850,I89841,I89856,I89844,I89853,I89835,I89859,I89905,I89908,I89911,I89914,I89917,I89920,I89923,I89926,I89929,I2224,I2231);
PAT_1 I_1241 (I89905,I89923,I89905,I89917,I89908,I89914,I89920,I89926,I89929,I89911,I89908,I89975,I89978,I89981,I89984,I89987,I89990,I89993,I89996,I89999,I2224,I2231);
PAT_12 I_1242 (I89987,I89981,I89999,I89975,I89984,I89975,I89978,I89996,I89990,I89978,I89993,I90045,I90048,I90051,I90054,I90057,I90060,I90063,I90066,I2224,I2231);
PAT_9 I_1243 (I90054,I90060,I90045,I90051,I90057,I90048,I90045,I90048,I90066,I90051,I90063,I90112,I90115,I90118,I90121,I90124,I90127,I90130,I90133,I90136,I2224,I2231);
PAT_5 I_1244 (I90133,I90112,I90127,I90112,I90118,I90121,I90115,I90115,I90130,I90124,I90136,I90182,I90185,I90188,I90191,I90194,I90197,I90200,I90203,I90206,I90209,I2224,I2231);
PAT_9 I_1245 (I90197,I90194,I90203,I90200,I90191,I90182,I90188,I90209,I90185,I90206,I90182,I90255,I90258,I90261,I90264,I90267,I90270,I90273,I90276,I90279,I2224,I2231);
PAT_5 I_1246 (I90276,I90255,I90270,I90255,I90261,I90264,I90258,I90258,I90273,I90267,I90279,I90325,I90328,I90331,I90334,I90337,I90340,I90343,I90346,I90349,I90352,I2224,I2231);
PAT_7 I_1247 (I90343,I90346,I90352,I90349,I90334,I90331,I90325,I90337,I90325,I90328,I90340,I90398,I90401,I90404,I90407,I90410,I90413,I90416,I90419,I90422,I2224,I2231);
PAT_9 I_1248 (I90419,I90407,I90416,I90422,I90404,I90410,I90401,I90413,I90398,I90398,I90401,I90468,I90471,I90474,I90477,I90480,I90483,I90486,I90489,I90492,I2224,I2231);
PAT_8 I_1249 (I90489,I90477,I90486,I90468,I90471,I90483,I90492,I90471,I90474,I90480,I90468,I90538,I90541,I90544,I90547,I90550,I90553,I90556,I90559,I90562,I2224,I2231);
PAT_9 I_1250 (I90541,I90550,I90541,I90538,I90553,I90544,I90559,I90547,I90556,I90538,I90562,I90608,I90611,I90614,I90617,I90620,I90623,I90626,I90629,I90632,I2224,I2231);
PAT_17 I_1251 (I90611,I90617,I90632,I90623,I90626,I90614,I90608,I90620,I90608,I90611,I90629,I90678,I90681,I90684,I90687,I90690,I90693,I90696,I90699,I90702,I90705,I2224,I2231);
PAT_11 I_1252 (I90690,I90699,I90705,I90681,I90678,I90696,I90687,I90693,I90684,I90702,I90678,I90751,I90754,I90757,I90760,I90763,I90766,I90769,I90772,I90775,I90778,I2224,I2231);
PAT_6 I_1253 (I90751,I90778,I90766,I90775,I90769,I90763,I90754,I90772,I90760,I90757,I90751,I90824,I90827,I90830,I90833,I90836,I90839,I90842,I90845,I90848,I90851,I2224,I2231);
PAT_13 I_1254 (I90848,I90830,I90845,I90824,I90827,I90833,I90851,I90836,I90842,I90824,I90839,I90897,I90900,I90903,I90906,I90909,I90912,I90915,I90918,I90921,I2224,I2231);
PAT_6 I_1255 (I90897,I90909,I90906,I90918,I90915,I90921,I90897,I90912,I90900,I90900,I90903,I90967,I90970,I90973,I90976,I90979,I90982,I90985,I90988,I90991,I90994,I2224,I2231);
PAT_10 I_1256 (I90967,I90982,I90985,I90976,I90967,I90991,I90994,I90970,I90979,I90973,I90988,I91040,I91043,I91046,I91049,I91052,I91055,I91058,I91061,I2224,I2231);
PAT_2 I_1257 (I91052,I91055,I91046,I91058,I91043,I91040,I91040,I91046,I91061,I91049,I91043,I91107,I91110,I91113,I91116,I91119,I91122,I91125,I91128,I91131,I2224,I2231);
PAT_13 I_1258 (I91116,I91110,I91107,I91128,I91119,I91122,I91110,I91113,I91125,I91131,I91107,I91177,I91180,I91183,I91186,I91189,I91192,I91195,I91198,I91201,I2224,I2231);
PAT_11 I_1259 (I91177,I91189,I91192,I91183,I91180,I91201,I91180,I91198,I91186,I91177,I91195,I91247,I91250,I91253,I91256,I91259,I91262,I91265,I91268,I91271,I91274,I2224,I2231);
PAT_2 I_1260 (I91247,I91271,I91259,I91253,I91262,I91265,I91250,I91274,I91268,I91256,I91247,I91320,I91323,I91326,I91329,I91332,I91335,I91338,I91341,I91344,I2224,I2231);
PAT_4 I_1261 (I91320,I91326,I91344,I91338,I91335,I91332,I91323,I91341,I91320,I91323,I91329,I91390,I91393,I91396,I91399,I91402,I91405,I91408,I91411,I91414,I2224,I2231);
PAT_10 I_1262 (I91390,I91390,I91414,I91393,I91399,I91408,I91405,I91393,I91411,I91396,I91402,I91460,I91463,I91466,I91469,I91472,I91475,I91478,I91481,I2224,I2231);
PAT_5 I_1263 (I91481,I91460,I91469,I91463,I91478,I91475,I91466,I91466,I91460,I91463,I91472,I91527,I91530,I91533,I91536,I91539,I91542,I91545,I91548,I91551,I91554,I2224,I2231);
PAT_4 I_1264 (I91545,I91551,I91554,I91533,I91536,I91548,I91530,I91527,I91539,I91542,I91527,I91600,I91603,I91606,I91609,I91612,I91615,I91618,I91621,I91624,I2224,I2231);
PAT_11 I_1265 (I91612,I91621,I91603,I91615,I91600,I91603,I91600,I91609,I91624,I91618,I91606,I91670,I91673,I91676,I91679,I91682,I91685,I91688,I91691,I91694,I91697,I2224,I2231);
PAT_13 I_1266 (I91670,I91673,I91682,I91694,I91697,I91685,I91691,I91679,I91688,I91676,I91670,I91743,I91746,I91749,I91752,I91755,I91758,I91761,I91764,I91767,I2224,I2231);
PAT_4 I_1267 (I91752,I91755,I91767,I91749,I91764,I91761,I91746,I91758,I91746,I91743,I91743,I91813,I91816,I91819,I91822,I91825,I91828,I91831,I91834,I91837,I2224,I2231);
PAT_11 I_1268 (I91825,I91834,I91816,I91828,I91813,I91816,I91813,I91822,I91837,I91831,I91819,I91883,I91886,I91889,I91892,I91895,I91898,I91901,I91904,I91907,I91910,I2224,I2231);
PAT_13 I_1269 (I91883,I91886,I91895,I91907,I91910,I91898,I91904,I91892,I91901,I91889,I91883,I91956,I91959,I91962,I91965,I91968,I91971,I91974,I91977,I91980,I2224,I2231);
PAT_6 I_1270 (I91956,I91968,I91965,I91977,I91974,I91980,I91956,I91971,I91959,I91959,I91962,I92026,I92029,I92032,I92035,I92038,I92041,I92044,I92047,I92050,I92053,I2224,I2231);
PAT_8 I_1271 (I92035,I92041,I92032,I92044,I92026,I92029,I92047,I92026,I92053,I92050,I92038,I92099,I92102,I92105,I92108,I92111,I92114,I92117,I92120,I92123,I2224,I2231);
PAT_13 I_1272 (I92111,I92120,I92102,I92123,I92105,I92099,I92099,I92108,I92117,I92114,I92102,I92169,I92172,I92175,I92178,I92181,I92184,I92187,I92190,I92193,I2224,I2231);
PAT_2 I_1273 (I92187,I92181,I92178,I92184,I92169,I92193,I92172,I92190,I92169,I92175,I92172,I92239,I92242,I92245,I92248,I92251,I92254,I92257,I92260,I92263,I2224,I2231);
PAT_11 I_1274 (I92242,I92254,I92239,I92251,I92248,I92260,I92257,I92242,I92263,I92245,I92239,I92309,I92312,I92315,I92318,I92321,I92324,I92327,I92330,I92333,I92336,I2224,I2231);
PAT_13 I_1275 (I92309,I92312,I92321,I92333,I92336,I92324,I92330,I92318,I92327,I92315,I92309,I92382,I92385,I92388,I92391,I92394,I92397,I92400,I92403,I92406,I2224,I2231);
PAT_10 I_1276 (I92403,I92397,I92391,I92385,I92406,I92385,I92394,I92382,I92382,I92400,I92388,I92452,I92455,I92458,I92461,I92464,I92467,I92470,I92473,I2224,I2231);
PAT_13 I_1277 (I92458,I92464,I92458,I92455,I92470,I92473,I92452,I92452,I92467,I92455,I92461,I92519,I92522,I92525,I92528,I92531,I92534,I92537,I92540,I92543,I2224,I2231);
PAT_6 I_1278 (I92519,I92531,I92528,I92540,I92537,I92543,I92519,I92534,I92522,I92522,I92525,I92589,I92592,I92595,I92598,I92601,I92604,I92607,I92610,I92613,I92616,I2224,I2231);
PAT_17 I_1279 (I92601,I92604,I92610,I92598,I92592,I92613,I92607,I92589,I92616,I92595,I92589,I92662,I92665,I92668,I92671,I92674,I92677,I92680,I92683,I92686,I92689,I2224,I2231);
PAT_14 I_1280 (I92665,I92680,I92662,I92686,I92671,I92677,I92662,I92683,I92668,I92689,I92674,I92735,I92738,I92741,I92744,I92747,I92750,I92753,I92756,I92759,I2224,I2231);
PAT_11 I_1281 (I92747,I92744,I92741,I92735,I92738,I92738,I92750,I92735,I92756,I92759,I92753,I92805,I92808,I92811,I92814,I92817,I92820,I92823,I92826,I92829,I92832,I2224,I2231);
PAT_4 I_1282 (I92811,I92832,I92805,I92823,I92814,I92805,I92826,I92808,I92817,I92829,I92820,I92878,I92881,I92884,I92887,I92890,I92893,I92896,I92899,I92902,I2224,I2231);
PAT_10 I_1283 (I92878,I92878,I92902,I92881,I92887,I92896,I92893,I92881,I92899,I92884,I92890,I92948,I92951,I92954,I92957,I92960,I92963,I92966,I92969,I2224,I2231);
PAT_5 I_1284 (I92969,I92948,I92957,I92951,I92966,I92963,I92954,I92954,I92948,I92951,I92960,I93015,I93018,I93021,I93024,I93027,I93030,I93033,I93036,I93039,I93042,I2224,I2231);
PAT_6 I_1285 (I93033,I93027,I93015,I93021,I93018,I93024,I93030,I93015,I93039,I93036,I93042,I93088,I93091,I93094,I93097,I93100,I93103,I93106,I93109,I93112,I93115,I2224,I2231);
PAT_13 I_1286 (I93112,I93094,I93109,I93088,I93091,I93097,I93115,I93100,I93106,I93088,I93103,I93161,I93164,I93167,I93170,I93173,I93176,I93179,I93182,I93185,I2224,I2231);
PAT_5 I_1287 (I93173,I93164,I93170,I93182,I93164,I93185,I93167,I93176,I93161,I93161,I93179,I93231,I93234,I93237,I93240,I93243,I93246,I93249,I93252,I93255,I93258,I2224,I2231);
PAT_9 I_1288 (I93246,I93243,I93252,I93249,I93240,I93231,I93237,I93258,I93234,I93255,I93231,I93304,I93307,I93310,I93313,I93316,I93319,I93322,I93325,I93328,I2224,I2231);
PAT_4 I_1289 (I93304,I93328,I93322,I93310,I93307,I93325,I93307,I93304,I93319,I93313,I93316,I93374,I93377,I93380,I93383,I93386,I93389,I93392,I93395,I93398,I2224,I2231);
PAT_13 I_1290 (I93389,I93383,I93395,I93380,I93386,I93374,I93398,I93392,I93377,I93374,I93377,I93444,I93447,I93450,I93453,I93456,I93459,I93462,I93465,I93468,I2224,I2231);
PAT_4 I_1291 (I93453,I93456,I93468,I93450,I93465,I93462,I93447,I93459,I93447,I93444,I93444,I93514,I93517,I93520,I93523,I93526,I93529,I93532,I93535,I93538,I2224,I2231);
PAT_12 I_1292 (I93514,I93517,I93535,I93538,I93529,I93520,I93526,I93523,I93514,I93532,I93517,I93584,I93587,I93590,I93593,I93596,I93599,I93602,I93605,I2224,I2231);
PAT_10 I_1293 (I93584,I93605,I93596,I93599,I93590,I93587,I93584,I93602,I93590,I93593,I93587,I93651,I93654,I93657,I93660,I93663,I93666,I93669,I93672,I2224,I2231);
PAT_8 I_1294 (I93672,I93663,I93654,I93651,I93660,I93651,I93666,I93654,I93669,I93657,I93657,I93718,I93721,I93724,I93727,I93730,I93733,I93736,I93739,I93742,I2224,I2231);
PAT_14 I_1295 (I93724,I93736,I93721,I93718,I93721,I93742,I93718,I93730,I93733,I93739,I93727,I93788,I93791,I93794,I93797,I93800,I93803,I93806,I93809,I93812,I2224,I2231);
PAT_2 I_1296 (I93806,I93812,I93797,I93788,I93791,I93791,I93803,I93788,I93809,I93794,I93800,I93858,I93861,I93864,I93867,I93870,I93873,I93876,I93879,I93882,I2224,I2231);
PAT_11 I_1297 (I93861,I93873,I93858,I93870,I93867,I93879,I93876,I93861,I93882,I93864,I93858,I93928,I93931,I93934,I93937,I93940,I93943,I93946,I93949,I93952,I93955,I2224,I2231);
PAT_17 I_1298 (I93940,I93931,I93955,I93928,I93937,I93949,I93946,I93943,I93928,I93952,I93934,I94001,I94004,I94007,I94010,I94013,I94016,I94019,I94022,I94025,I94028,I2224,I2231);
PAT_6 I_1299 (I94001,I94019,I94007,I94010,I94016,I94001,I94013,I94004,I94025,I94028,I94022,I94074,I94077,I94080,I94083,I94086,I94089,I94092,I94095,I94098,I94101,I2224,I2231);
PAT_0 I_1300 (I94074,I94092,I94086,I94098,I94080,I94101,I94083,I94074,I94089,I94095,I94077,I94147,I94150,I94153,I94156,I94159,I94162,I94165,I94168,I2224,I2231);
PAT_2 I_1301 (I94153,I94156,I94165,I94150,I94153,I94150,I94159,I94147,I94147,I94162,I94168,I94214,I94217,I94220,I94223,I94226,I94229,I94232,I94235,I94238,I2224,I2231);
PAT_4 I_1302 (I94214,I94220,I94238,I94232,I94229,I94226,I94217,I94235,I94214,I94217,I94223,I94284,I94287,I94290,I94293,I94296,I94299,I94302,I94305,I94308,I2224,I2231);
PAT_17 I_1303 (I94296,I94293,I94305,I94299,I94284,I94302,I94308,I94287,I94290,I94287,I94284,I94354,I94357,I94360,I94363,I94366,I94369,I94372,I94375,I94378,I94381,I2224,I2231);
PAT_6 I_1304 (I94354,I94372,I94360,I94363,I94369,I94354,I94366,I94357,I94378,I94381,I94375,I94427,I94430,I94433,I94436,I94439,I94442,I94445,I94448,I94451,I94454,I2224,I2231);
PAT_11 I_1305 (I94427,I94442,I94427,I94439,I94436,I94454,I94451,I94448,I94445,I94430,I94433,I94500,I94503,I94506,I94509,I94512,I94515,I94518,I94521,I94524,I94527,I2224,I2231);
PAT_13 I_1306 (I94500,I94503,I94512,I94524,I94527,I94515,I94521,I94509,I94518,I94506,I94500,I94573,I94576,I94579,I94582,I94585,I94588,I94591,I94594,I94597,I2224,I2231);
PAT_9 I_1307 (I94594,I94576,I94576,I94573,I94597,I94579,I94582,I94573,I94585,I94591,I94588,I94643,I94646,I94649,I94652,I94655,I94658,I94661,I94664,I94667,I2224,I2231);
PAT_13 I_1308 (I94643,I94664,I94646,I94661,I94655,I94652,I94667,I94643,I94649,I94658,I94646,I94713,I94716,I94719,I94722,I94725,I94728,I94731,I94734,I94737,I2224,I2231);
PAT_10 I_1309 (I94734,I94728,I94722,I94716,I94737,I94716,I94725,I94713,I94713,I94731,I94719,I94783,I94786,I94789,I94792,I94795,I94798,I94801,I94804,I2224,I2231);
PAT_9 I_1310 (I94795,I94783,I94786,I94789,I94783,I94789,I94792,I94786,I94804,I94798,I94801,I94850,I94853,I94856,I94859,I94862,I94865,I94868,I94871,I94874,I2224,I2231);
PAT_5 I_1311 (I94871,I94850,I94865,I94850,I94856,I94859,I94853,I94853,I94868,I94862,I94874,I94920,I94923,I94926,I94929,I94932,I94935,I94938,I94941,I94944,I94947,I2224,I2231);
PAT_4 I_1312 (I94938,I94944,I94947,I94926,I94929,I94941,I94923,I94920,I94932,I94935,I94920,I94993,I94996,I94999,I95002,I95005,I95008,I95011,I95014,I95017,I2224,I2231);
PAT_11 I_1313 (I95005,I95014,I94996,I95008,I94993,I94996,I94993,I95002,I95017,I95011,I94999,I95063,I95066,I95069,I95072,I95075,I95078,I95081,I95084,I95087,I95090,I2224,I2231);
PAT_13 I_1314 (I95063,I95066,I95075,I95087,I95090,I95078,I95084,I95072,I95081,I95069,I95063,I95136,I95139,I95142,I95145,I95148,I95151,I95154,I95157,I95160,I2224,I2231);
PAT_7 I_1315 (I95145,I95148,I95136,I95151,I95157,I95142,I95139,I95160,I95139,I95136,I95154,I95206,I95209,I95212,I95215,I95218,I95221,I95224,I95227,I95230,I2224,I2231);
PAT_12 I_1316 (I95212,I95206,I95218,I95206,I95230,I95209,I95209,I95227,I95215,I95221,I95224,I95276,I95279,I95282,I95285,I95288,I95291,I95294,I95297,I2224,I2231);
PAT_2 I_1317 (I95294,I95288,I95297,I95291,I95285,I95282,I95276,I95276,I95282,I95279,I95279,I95343,I95346,I95349,I95352,I95355,I95358,I95361,I95364,I95367,I2224,I2231);
PAT_8 I_1318 (I95355,I95346,I95352,I95343,I95349,I95364,I95361,I95343,I95358,I95346,I95367,I95413,I95416,I95419,I95422,I95425,I95428,I95431,I95434,I95437,I2224,I2231);
PAT_1 I_1319 (I95416,I95437,I95419,I95434,I95416,I95422,I95413,I95413,I95431,I95428,I95425,I95483,I95486,I95489,I95492,I95495,I95498,I95501,I95504,I95507,I2224,I2231);
PAT_11 I_1320 (I95486,I95501,I95498,I95504,I95507,I95486,I95492,I95495,I95483,I95489,I95483,I95553,I95556,I95559,I95562,I95565,I95568,I95571,I95574,I95577,I95580,I2224,I2231);
PAT_4 I_1321 (I95559,I95580,I95553,I95571,I95562,I95553,I95574,I95556,I95565,I95577,I95568,I95626,I95629,I95632,I95635,I95638,I95641,I95644,I95647,I95650,I2224,I2231);
PAT_10 I_1322 (I95626,I95626,I95650,I95629,I95635,I95644,I95641,I95629,I95647,I95632,I95638,I95696,I95699,I95702,I95705,I95708,I95711,I95714,I95717,I2224,I2231);
PAT_9 I_1323 (I95708,I95696,I95699,I95702,I95696,I95702,I95705,I95699,I95717,I95711,I95714,I95763,I95766,I95769,I95772,I95775,I95778,I95781,I95784,I95787,I2224,I2231);
PAT_6 I_1324 (I95781,I95763,I95775,I95784,I95763,I95772,I95769,I95787,I95778,I95766,I95766,I95833,I95836,I95839,I95842,I95845,I95848,I95851,I95854,I95857,I95860,I2224,I2231);
PAT_10 I_1325 (I95833,I95848,I95851,I95842,I95833,I95857,I95860,I95836,I95845,I95839,I95854,I95906,I95909,I95912,I95915,I95918,I95921,I95924,I95927,I2224,I2231);
PAT_1 I_1326 (I95912,I95912,I95921,I95906,I95918,I95909,I95924,I95906,I95927,I95915,I95909,I95973,I95976,I95979,I95982,I95985,I95988,I95991,I95994,I95997,I2224,I2231);
PAT_7 I_1327 (I95976,I95982,I95979,I95985,I95991,I95988,I95997,I95994,I95976,I95973,I95973,I96043,I96046,I96049,I96052,I96055,I96058,I96061,I96064,I96067,I2224,I2231);
PAT_9 I_1328 (I96064,I96052,I96061,I96067,I96049,I96055,I96046,I96058,I96043,I96043,I96046,I96113,I96116,I96119,I96122,I96125,I96128,I96131,I96134,I96137,I2224,I2231);
PAT_2 I_1329 (I96128,I96131,I96122,I96137,I96113,I96116,I96119,I96116,I96134,I96125,I96113,I96183,I96186,I96189,I96192,I96195,I96198,I96201,I96204,I96207,I2224,I2231);
PAT_11 I_1330 (I96186,I96198,I96183,I96195,I96192,I96204,I96201,I96186,I96207,I96189,I96183,I96253,I96256,I96259,I96262,I96265,I96268,I96271,I96274,I96277,I96280,I2224,I2231);
PAT_9 I_1331 (I96259,I96271,I96262,I96274,I96253,I96256,I96265,I96253,I96268,I96277,I96280,I96326,I96329,I96332,I96335,I96338,I96341,I96344,I96347,I96350,I2224,I2231);
PAT_10 I_1332 (I96347,I96344,I96332,I96329,I96350,I96335,I96341,I96329,I96326,I96326,I96338,I96396,I96399,I96402,I96405,I96408,I96411,I96414,I96417,I2224,I2231);
PAT_15 I_1333 (I96411,I96414,I96402,I96408,I96396,I96396,I96402,I96417,I96405,I96399,I96399,I96463,I96466,I96469,I96472,I96475,I96478,I96481,I96484,I96487,I2224,I2231);
PAT_6 I_1334 (I96466,I96463,I96469,I96484,I96466,I96487,I96472,I96478,I96475,I96481,I96463,I96533,I96536,I96539,I96542,I96545,I96548,I96551,I96554,I96557,I96560,I2224,I2231);
PAT_5 I_1335 (I96554,I96533,I96539,I96542,I96548,I96551,I96533,I96557,I96536,I96545,I96560,I96606,I96609,I96612,I96615,I96618,I96621,I96624,I96627,I96630,I96633,I2224,I2231);
PAT_17 I_1336 (I96633,I96609,I96612,I96615,I96606,I96618,I96606,I96630,I96624,I96621,I96627,I96679,I96682,I96685,I96688,I96691,I96694,I96697,I96700,I96703,I96706,I2224,I2231);
PAT_9 I_1337 (I96700,I96682,I96688,I96703,I96685,I96697,I96679,I96691,I96679,I96706,I96694,I96752,I96755,I96758,I96761,I96764,I96767,I96770,I96773,I96776,I2224,I2231);
PAT_4 I_1338 (I96752,I96776,I96770,I96758,I96755,I96773,I96755,I96752,I96767,I96761,I96764,I96822,I96825,I96828,I96831,I96834,I96837,I96840,I96843,I96846,I2224,I2231);
PAT_9 I_1339 (I96843,I96825,I96828,I96837,I96840,I96822,I96831,I96825,I96846,I96822,I96834,I96892,I96895,I96898,I96901,I96904,I96907,I96910,I96913,I96916,I2224,I2231);
PAT_8 I_1340 (I96913,I96901,I96910,I96892,I96895,I96907,I96916,I96895,I96898,I96904,I96892,I96962,I96965,I96968,I96971,I96974,I96977,I96980,I96983,I96986,I2224,I2231);
PAT_15 I_1341 (I96974,I96983,I96977,I96986,I96962,I96968,I96965,I96971,I96962,I96965,I96980,I97032,I97035,I97038,I97041,I97044,I97047,I97050,I97053,I97056,I2224,I2231);
PAT_7 I_1342 (I97032,I97044,I97032,I97056,I97038,I97035,I97050,I97035,I97053,I97047,I97041,I97102,I97105,I97108,I97111,I97114,I97117,I97120,I97123,I97126,I2224,I2231);
PAT_8 I_1343 (I97108,I97120,I97102,I97105,I97111,I97102,I97126,I97123,I97114,I97117,I97105,I97172,I97175,I97178,I97181,I97184,I97187,I97190,I97193,I97196,I2224,I2231);
PAT_13 I_1344 (I97184,I97193,I97175,I97196,I97178,I97172,I97172,I97181,I97190,I97187,I97175,I97242,I97245,I97248,I97251,I97254,I97257,I97260,I97263,I97266,I2224,I2231);
PAT_2 I_1345 (I97260,I97254,I97251,I97257,I97242,I97266,I97245,I97263,I97242,I97248,I97245,I97312,I97315,I97318,I97321,I97324,I97327,I97330,I97333,I97336,I2224,I2231);
PAT_11 I_1346 (I97315,I97327,I97312,I97324,I97321,I97333,I97330,I97315,I97336,I97318,I97312,I97382,I97385,I97388,I97391,I97394,I97397,I97400,I97403,I97406,I97409,I2224,I2231);
PAT_5 I_1347 (I97403,I97382,I97409,I97397,I97394,I97406,I97388,I97382,I97400,I97385,I97391,I97455,I97458,I97461,I97464,I97467,I97470,I97473,I97476,I97479,I97482,I2224,I2231);
PAT_6 I_1348 (I97473,I97467,I97455,I97461,I97458,I97464,I97470,I97455,I97479,I97476,I97482,I97528,I97531,I97534,I97537,I97540,I97543,I97546,I97549,I97552,I97555,I2224,I2231);
PAT_3 I_1349 (I97531,I97528,I97528,I97540,I97537,I97555,I97534,I97543,I97546,I97552,I97549,I97601,I97604,I97607,I97610,I97613,I97616,I97619,I97622,I97625,I97628,I2224,I2231);
PAT_2 I_1350 (I97628,I97613,I97604,I97601,I97625,I97616,I97610,I97619,I97601,I97622,I97607,I97674,I97677,I97680,I97683,I97686,I97689,I97692,I97695,I97698,I2224,I2231);
PAT_8 I_1351 (I97686,I97677,I97683,I97674,I97680,I97695,I97692,I97674,I97689,I97677,I97698,I97744,I97747,I97750,I97753,I97756,I97759,I97762,I97765,I97768,I2224,I2231);
PAT_13 I_1352 (I97756,I97765,I97747,I97768,I97750,I97744,I97744,I97753,I97762,I97759,I97747,I97814,I97817,I97820,I97823,I97826,I97829,I97832,I97835,I97838,I2224,I2231);
PAT_15 I_1353 (I97814,I97826,I97817,I97829,I97814,I97823,I97838,I97835,I97820,I97832,I97817,I97884,I97887,I97890,I97893,I97896,I97899,I97902,I97905,I97908,I2224,I2231);
PAT_10 I_1354 (I97887,I97896,I97890,I97884,I97905,I97908,I97893,I97884,I97887,I97902,I97899,I97954,I97957,I97960,I97963,I97966,I97969,I97972,I97975,I2224,I2231);
PAT_2 I_1355 (I97966,I97969,I97960,I97972,I97957,I97954,I97954,I97960,I97975,I97963,I97957,I98021,I98024,I98027,I98030,I98033,I98036,I98039,I98042,I98045,I2224,I2231);
PAT_6 I_1356 (I98045,I98021,I98036,I98033,I98039,I98030,I98024,I98042,I98021,I98027,I98024,I98091,I98094,I98097,I98100,I98103,I98106,I98109,I98112,I98115,I98118,I2224,I2231);
PAT_9 I_1357 (I98091,I98118,I98115,I98097,I98103,I98094,I98106,I98091,I98109,I98100,I98112,I98164,I98167,I98170,I98173,I98176,I98179,I98182,I98185,I98188,I2224,I2231);
PAT_13 I_1358 (I98164,I98185,I98167,I98182,I98176,I98173,I98188,I98164,I98170,I98179,I98167,I98234,I98237,I98240,I98243,I98246,I98249,I98252,I98255,I98258,I2224,I2231);
PAT_1 I_1359 (I98234,I98243,I98237,I98255,I98249,I98240,I98252,I98246,I98237,I98258,I98234,I98304,I98307,I98310,I98313,I98316,I98319,I98322,I98325,I98328,I2224,I2231);
PAT_0 I_1360 (I98304,I98307,I98307,I98325,I98310,I98316,I98304,I98322,I98328,I98319,I98313,I98374,I98377,I98380,I98383,I98386,I98389,I98392,I98395,I2224,I2231);
PAT_2 I_1361 (I98380,I98383,I98392,I98377,I98380,I98377,I98386,I98374,I98374,I98389,I98395,I98441,I98444,I98447,I98450,I98453,I98456,I98459,I98462,I98465,I2224,I2231);
PAT_17 I_1362 (I98441,I98441,I98453,I98444,I98447,I98459,I98456,I98465,I98444,I98450,I98462,I98511,I98514,I98517,I98520,I98523,I98526,I98529,I98532,I98535,I98538,I2224,I2231);
PAT_8 I_1363 (I98520,I98532,I98538,I98529,I98514,I98523,I98526,I98535,I98517,I98511,I98511,I98584,I98587,I98590,I98593,I98596,I98599,I98602,I98605,I98608,I2224,I2231);
PAT_11 I_1364 (I98605,I98596,I98584,I98587,I98602,I98590,I98593,I98584,I98608,I98599,I98587,I98654,I98657,I98660,I98663,I98666,I98669,I98672,I98675,I98678,I98681,I2224,I2231);
PAT_17 I_1365 (I98666,I98657,I98681,I98654,I98663,I98675,I98672,I98669,I98654,I98678,I98660,I98727,I98730,I98733,I98736,I98739,I98742,I98745,I98748,I98751,I98754,I2224,I2231);
PAT_7 I_1366 (I98745,I98736,I98742,I98730,I98739,I98748,I98754,I98727,I98751,I98733,I98727,I98800,I98803,I98806,I98809,I98812,I98815,I98818,I98821,I98824,I2224,I2231);
PAT_5 I_1367 (I98806,I98800,I98809,I98818,I98812,I98824,I98821,I98803,I98815,I98803,I98800,I98870,I98873,I98876,I98879,I98882,I98885,I98888,I98891,I98894,I98897,I2224,I2231);
PAT_6 I_1368 (I98888,I98882,I98870,I98876,I98873,I98879,I98885,I98870,I98894,I98891,I98897,I98943,I98946,I98949,I98952,I98955,I98958,I98961,I98964,I98967,I98970,I2224,I2231);
PAT_10 I_1369 (I98943,I98958,I98961,I98952,I98943,I98967,I98970,I98946,I98955,I98949,I98964,I99016,I99019,I99022,I99025,I99028,I99031,I99034,I99037,I2224,I2231);
PAT_9 I_1370 (I99028,I99016,I99019,I99022,I99016,I99022,I99025,I99019,I99037,I99031,I99034,I99083,I99086,I99089,I99092,I99095,I99098,I99101,I99104,I99107,I2224,I2231);
PAT_4 I_1371 (I99083,I99107,I99101,I99089,I99086,I99104,I99086,I99083,I99098,I99092,I99095,I99153,I99156,I99159,I99162,I99165,I99168,I99171,I99174,I99177,I2224,I2231);
PAT_8 I_1372 (I99165,I99153,I99174,I99159,I99156,I99177,I99162,I99171,I99156,I99153,I99168,I99223,I99226,I99229,I99232,I99235,I99238,I99241,I99244,I99247,I2224,I2231);
PAT_6 I_1373 (I99226,I99223,I99229,I99241,I99238,I99232,I99235,I99223,I99244,I99226,I99247,I99293,I99296,I99299,I99302,I99305,I99308,I99311,I99314,I99317,I99320,I2224,I2231);
PAT_10 I_1374 (I99293,I99308,I99311,I99302,I99293,I99317,I99320,I99296,I99305,I99299,I99314,I99366,I99369,I99372,I99375,I99378,I99381,I99384,I99387,I2224,I2231);
PAT_8 I_1375 (I99387,I99378,I99369,I99366,I99375,I99366,I99381,I99369,I99384,I99372,I99372,I99433,I99436,I99439,I99442,I99445,I99448,I99451,I99454,I99457,I2224,I2231);
PAT_15 I_1376 (I99445,I99454,I99448,I99457,I99433,I99439,I99436,I99442,I99433,I99436,I99451,I99503,I99506,I99509,I99512,I99515,I99518,I99521,I99524,I99527,I2224,I2231);
PAT_5 I_1377 (I99506,I99503,I99509,I99527,I99524,I99512,I99521,I99515,I99506,I99518,I99503,I99573,I99576,I99579,I99582,I99585,I99588,I99591,I99594,I99597,I99600,I2224,I2231);
PAT_10 I_1378 (I99597,I99600,I99579,I99585,I99588,I99594,I99576,I99573,I99573,I99582,I99591,I99646,I99649,I99652,I99655,I99658,I99661,I99664,I99667,I2224,I2231);
PAT_14 I_1379 (I99646,I99667,I99652,I99661,I99658,I99664,I99655,I99649,I99649,I99652,I99646,I99713,I99716,I99719,I99722,I99725,I99728,I99731,I99734,I99737,I2224,I2231);
PAT_9 I_1380 (I99722,I99734,I99713,I99731,I99716,I99719,I99737,I99716,I99725,I99713,I99728,I99783,I99786,I99789,I99792,I99795,I99798,I99801,I99804,I99807,I2224,I2231);
PAT_13 I_1381 (I99783,I99804,I99786,I99801,I99795,I99792,I99807,I99783,I99789,I99798,I99786,I99853,I99856,I99859,I99862,I99865,I99868,I99871,I99874,I99877,I2224,I2231);
PAT_6 I_1382 (I99853,I99865,I99862,I99874,I99871,I99877,I99853,I99868,I99856,I99856,I99859,I99923,I99926,I99929,I99932,I99935,I99938,I99941,I99944,I99947,I99950,I2224,I2231);
PAT_15 I_1383 (I99941,I99932,I99944,I99947,I99938,I99950,I99923,I99929,I99923,I99926,I99935,I99996,I99999,I100002,I100005,I100008,I100011,I100014,I100017,I100020,I2224,I2231);
PAT_5 I_1384 (I99999,I99996,I100002,I100020,I100017,I100005,I100014,I100008,I99999,I100011,I99996,I100066,I100069,I100072,I100075,I100078,I100081,I100084,I100087,I100090,I100093,I2224,I2231);
PAT_6 I_1385 (I100084,I100078,I100066,I100072,I100069,I100075,I100081,I100066,I100090,I100087,I100093,I100139,I100142,I100145,I100148,I100151,I100154,I100157,I100160,I100163,I100166,I2224,I2231);
PAT_7 I_1386 (I100145,I100154,I100157,I100139,I100148,I100142,I100151,I100166,I100160,I100163,I100139,I100212,I100215,I100218,I100221,I100224,I100227,I100230,I100233,I100236,I2224,I2231);
PAT_8 I_1387 (I100218,I100230,I100212,I100215,I100221,I100212,I100236,I100233,I100224,I100227,I100215,I100282,I100285,I100288,I100291,I100294,I100297,I100300,I100303,I100306,I2224,I2231);
PAT_1 I_1388 (I100285,I100306,I100288,I100303,I100285,I100291,I100282,I100282,I100300,I100297,I100294,I100352,I100355,I100358,I100361,I100364,I100367,I100370,I100373,I100376,I2224,I2231);
PAT_11 I_1389 (I100355,I100370,I100367,I100373,I100376,I100355,I100361,I100364,I100352,I100358,I100352,I100422,I100425,I100428,I100431,I100434,I100437,I100440,I100443,I100446,I100449,I2224,I2231);
PAT_5 I_1390 (I100443,I100422,I100449,I100437,I100434,I100446,I100428,I100422,I100440,I100425,I100431,I100495,I100498,I100501,I100504,I100507,I100510,I100513,I100516,I100519,I100522,I2224,I2231);
PAT_9 I_1391 (I100510,I100507,I100516,I100513,I100504,I100495,I100501,I100522,I100498,I100519,I100495,I100568,I100571,I100574,I100577,I100580,I100583,I100586,I100589,I100592,I2224,I2231);
PAT_8 I_1392 (I100589,I100577,I100586,I100568,I100571,I100583,I100592,I100571,I100574,I100580,I100568,I100638,I100641,I100644,I100647,I100650,I100653,I100656,I100659,I100662,I2224,I2231);
PAT_9 I_1393 (I100641,I100650,I100641,I100638,I100653,I100644,I100659,I100647,I100656,I100638,I100662,I100708,I100711,I100714,I100717,I100720,I100723,I100726,I100729,I100732,I2224,I2231);
PAT_12 I_1394 (I100729,I100726,I100720,I100708,I100717,I100708,I100711,I100714,I100732,I100723,I100711,I100778,I100781,I100784,I100787,I100790,I100793,I100796,I100799,I2224,I2231);
PAT_10 I_1395 (I1593,I1489,I1865,I1897,I1929,I1977,I1993,I1761,I1969,I1369,I1601,I100845,I100848,I100851,I100854,I100857,I100860,I100863,I100866,I2224,I2231);
PAT_9 I_1396 (I100857,I100845,I100848,I100851,I100845,I100851,I100854,I100848,I100866,I100860,I100863,I100912,I100915,I100918,I100921,I100924,I100927,I100930,I100933,I100936,I2224,I2231);
PAT_11 I_1397 (I100924,I100930,I100936,I100933,I100921,I100915,I100915,I100912,I100927,I100912,I100918,I100982,I100985,I100988,I100991,I100994,I100997,I101000,I101003,I101006,I101009,I2224,I2231);
PAT_13 I_1398 (I100982,I100985,I100994,I101006,I101009,I100997,I101003,I100991,I101000,I100988,I100982,I101055,I101058,I101061,I101064,I101067,I101070,I101073,I101076,I101079,I2224,I2231);
PAT_4 I_1399 (I101064,I101067,I101079,I101061,I101076,I101073,I101058,I101070,I101058,I101055,I101055,I101125,I101128,I101131,I101134,I101137,I101140,I101143,I101146,I101149,I2224,I2231);
PAT_13 I_1400 (I101140,I101134,I101146,I101131,I101137,I101125,I101149,I101143,I101128,I101125,I101128,I101195,I101198,I101201,I101204,I101207,I101210,I101213,I101216,I101219,I2224,I2231);
PAT_11 I_1401 (I101195,I101207,I101210,I101201,I101198,I101219,I101198,I101216,I101204,I101195,I101213,I101265,I101268,I101271,I101274,I101277,I101280,I101283,I101286,I101289,I101292,I2224,I2231);
PAT_4 I_1402 (I101271,I101292,I101265,I101283,I101274,I101265,I101286,I101268,I101277,I101289,I101280,I101338,I101341,I101344,I101347,I101350,I101353,I101356,I101359,I101362,I2224,I2231);
PAT_7 I_1403 (I101353,I101347,I101344,I101338,I101350,I101356,I101341,I101341,I101359,I101362,I101338,I101408,I101411,I101414,I101417,I101420,I101423,I101426,I101429,I101432,I2224,I2231);
PAT_5 I_1404 (I101414,I101408,I101417,I101426,I101420,I101432,I101429,I101411,I101423,I101411,I101408,I101478,I101481,I101484,I101487,I101490,I101493,I101496,I101499,I101502,I101505,I2224,I2231);
PAT_3 I_1405 (I101490,I101478,I101505,I101499,I101502,I101478,I101493,I101481,I101484,I101487,I101496,I101551,I101554,I101557,I101560,I101563,I101566,I101569,I101572,I101575,I101578,I2224,I2231);
PAT_4 I_1406 (I101557,I101563,I101551,I101560,I101551,I101578,I101572,I101566,I101575,I101554,I101569,I101624,I101627,I101630,I101633,I101636,I101639,I101642,I101645,I101648,I2224,I2231);
PAT_14 I_1407 (I101627,I101642,I101639,I101624,I101636,I101627,I101624,I101630,I101645,I101633,I101648,I101694,I101697,I101700,I101703,I101706,I101709,I101712,I101715,I101718,I2224,I2231);
PAT_17 I_1408 (I101709,I101697,I101718,I101694,I101715,I101703,I101700,I101712,I101706,I101697,I101694,I101764,I101767,I101770,I101773,I101776,I101779,I101782,I101785,I101788,I101791,I2224,I2231);
PAT_14 I_1409 (I101767,I101782,I101764,I101788,I101773,I101779,I101764,I101785,I101770,I101791,I101776,I101837,I101840,I101843,I101846,I101849,I101852,I101855,I101858,I101861,I2224,I2231);
PAT_8 I_1410 (I101843,I101846,I101840,I101852,I101861,I101840,I101837,I101858,I101837,I101849,I101855,I101907,I101910,I101913,I101916,I101919,I101922,I101925,I101928,I101931,I2224,I2231);
PAT_4 I_1411 (I101925,I101910,I101916,I101907,I101907,I101919,I101910,I101928,I101931,I101913,I101922,I101977,I101980,I101983,I101986,I101989,I101992,I101995,I101998,I102001,I2224,I2231);
PAT_5 I_1412 (I101998,I101980,I101980,I101992,I101995,I101989,I101986,I101977,I101983,I101977,I102001,I102047,I102050,I102053,I102056,I102059,I102062,I102065,I102068,I102071,I102074,I2224,I2231);
PAT_11 I_1413 (I102059,I102056,I102050,I102068,I102071,I102047,I102065,I102062,I102074,I102053,I102047,I102120,I102123,I102126,I102129,I102132,I102135,I102138,I102141,I102144,I102147,I2224,I2231);
PAT_2 I_1414 (I102120,I102144,I102132,I102126,I102135,I102138,I102123,I102147,I102141,I102129,I102120,I102193,I102196,I102199,I102202,I102205,I102208,I102211,I102214,I102217,I2224,I2231);
PAT_5 I_1415 (I102214,I102193,I102193,I102205,I102202,I102211,I102199,I102208,I102217,I102196,I102196,I102263,I102266,I102269,I102272,I102275,I102278,I102281,I102284,I102287,I102290,I2224,I2231);
PAT_6 I_1416 (I102281,I102275,I102263,I102269,I102266,I102272,I102278,I102263,I102287,I102284,I102290,I102336,I102339,I102342,I102345,I102348,I102351,I102354,I102357,I102360,I102363,I2224,I2231);
PAT_7 I_1417 (I102342,I102351,I102354,I102336,I102345,I102339,I102348,I102363,I102357,I102360,I102336,I102409,I102412,I102415,I102418,I102421,I102424,I102427,I102430,I102433,I2224,I2231);
PAT_1 I_1418 (I102409,I102427,I102430,I102412,I102433,I102421,I102415,I102424,I102412,I102418,I102409,I102479,I102482,I102485,I102488,I102491,I102494,I102497,I102500,I102503,I2224,I2231);
PAT_13 I_1419 (I102488,I102497,I102503,I102479,I102494,I102491,I102500,I102485,I102482,I102479,I102482,I102549,I102552,I102555,I102558,I102561,I102564,I102567,I102570,I102573,I2224,I2231);
PAT_2 I_1420 (I102567,I102561,I102558,I102564,I102549,I102573,I102552,I102570,I102549,I102555,I102552,I102619,I102622,I102625,I102628,I102631,I102634,I102637,I102640,I102643,I2224,I2231);
PAT_4 I_1421 (I102619,I102625,I102643,I102637,I102634,I102631,I102622,I102640,I102619,I102622,I102628,I102689,I102692,I102695,I102698,I102701,I102704,I102707,I102710,I102713,I2224,I2231);
PAT_11 I_1422 (I102701,I102710,I102692,I102704,I102689,I102692,I102689,I102698,I102713,I102707,I102695,I102759,I102762,I102765,I102768,I102771,I102774,I102777,I102780,I102783,I102786,I2224,I2231);
PAT_9 I_1423 (I102765,I102777,I102768,I102780,I102759,I102762,I102771,I102759,I102774,I102783,I102786,I102832,I102835,I102838,I102841,I102844,I102847,I102850,I102853,I102856,I2224,I2231);
PAT_4 I_1424 (I102832,I102856,I102850,I102838,I102835,I102853,I102835,I102832,I102847,I102841,I102844,I102902,I102905,I102908,I102911,I102914,I102917,I102920,I102923,I102926,I2224,I2231);
PAT_9 I_1425 (I102923,I102905,I102908,I102917,I102920,I102902,I102911,I102905,I102926,I102902,I102914,I102972,I102975,I102978,I102981,I102984,I102987,I102990,I102993,I102996,I2224,I2231);
PAT_4 I_1426 (I102972,I102996,I102990,I102978,I102975,I102993,I102975,I102972,I102987,I102981,I102984,I103042,I103045,I103048,I103051,I103054,I103057,I103060,I103063,I103066,I2224,I2231);
PAT_5 I_1427 (I103063,I103045,I103045,I103057,I103060,I103054,I103051,I103042,I103048,I103042,I103066,I103112,I103115,I103118,I103121,I103124,I103127,I103130,I103133,I103136,I103139,I2224,I2231);
PAT_8 I_1428 (I103112,I103139,I103130,I103127,I103121,I103112,I103124,I103136,I103115,I103133,I103118,I103185,I103188,I103191,I103194,I103197,I103200,I103203,I103206,I103209,I2224,I2231);
PAT_7 I_1429 (I103185,I103194,I103191,I103197,I103203,I103185,I103188,I103206,I103209,I103200,I103188,I103255,I103258,I103261,I103264,I103267,I103270,I103273,I103276,I103279,I2224,I2231);
PAT_17 I_1430 (I103267,I103261,I103270,I103255,I103273,I103276,I103258,I103279,I103264,I103258,I103255,I103325,I103328,I103331,I103334,I103337,I103340,I103343,I103346,I103349,I103352,I2224,I2231);
PAT_13 I_1431 (I103343,I103346,I103331,I103325,I103337,I103349,I103328,I103340,I103325,I103352,I103334,I103398,I103401,I103404,I103407,I103410,I103413,I103416,I103419,I103422,I2224,I2231);
PAT_2 I_1432 (I103416,I103410,I103407,I103413,I103398,I103422,I103401,I103419,I103398,I103404,I103401,I103468,I103471,I103474,I103477,I103480,I103483,I103486,I103489,I103492,I2224,I2231);
PAT_7 I_1433 (I103492,I103468,I103474,I103471,I103471,I103480,I103483,I103468,I103486,I103489,I103477,I103538,I103541,I103544,I103547,I103550,I103553,I103556,I103559,I103562,I2224,I2231);
PAT_2 I_1434 (I103559,I103553,I103544,I103538,I103547,I103541,I103550,I103562,I103556,I103541,I103538,I103608,I103611,I103614,I103617,I103620,I103623,I103626,I103629,I103632,I2224,I2231);
PAT_12 I_1435 (I103617,I103614,I103608,I103611,I103632,I103626,I103629,I103611,I103623,I103608,I103620,I103678,I103681,I103684,I103687,I103690,I103693,I103696,I103699,I2224,I2231);
PAT_7 I_1436 (I103684,I103687,I103678,I103690,I103696,I103684,I103699,I103693,I103681,I103681,I103678,I103745,I103748,I103751,I103754,I103757,I103760,I103763,I103766,I103769,I2224,I2231);
PAT_15 I_1437 (I103763,I103748,I103748,I103760,I103745,I103769,I103751,I103757,I103766,I103745,I103754,I103815,I103818,I103821,I103824,I103827,I103830,I103833,I103836,I103839,I2224,I2231);
PAT_6 I_1438 (I103818,I103815,I103821,I103836,I103818,I103839,I103824,I103830,I103827,I103833,I103815,I103885,I103888,I103891,I103894,I103897,I103900,I103903,I103906,I103909,I103912,I2224,I2231);
PAT_9 I_1439 (I103885,I103912,I103909,I103891,I103897,I103888,I103900,I103885,I103903,I103894,I103906,I103958,I103961,I103964,I103967,I103970,I103973,I103976,I103979,I103982,I2224,I2231);
PAT_2 I_1440 (I103973,I103976,I103967,I103982,I103958,I103961,I103964,I103961,I103979,I103970,I103958,I104028,I104031,I104034,I104037,I104040,I104043,I104046,I104049,I104052,I2224,I2231);
PAT_13 I_1441 (I104037,I104031,I104028,I104049,I104040,I104043,I104031,I104034,I104046,I104052,I104028,I104098,I104101,I104104,I104107,I104110,I104113,I104116,I104119,I104122,I2224,I2231);
PAT_17 I_1442 (I104122,I104110,I104119,I104116,I104107,I104098,I104101,I104104,I104098,I104113,I104101,I104168,I104171,I104174,I104177,I104180,I104183,I104186,I104189,I104192,I104195,I2224,I2231);
PAT_5 I_1443 (I104180,I104174,I104171,I104192,I104177,I104183,I104186,I104168,I104168,I104189,I104195,I104241,I104244,I104247,I104250,I104253,I104256,I104259,I104262,I104265,I104268,I2224,I2231);
PAT_9 I_1444 (I104256,I104253,I104262,I104259,I104250,I104241,I104247,I104268,I104244,I104265,I104241,I104314,I104317,I104320,I104323,I104326,I104329,I104332,I104335,I104338,I2224,I2231);
PAT_13 I_1445 (I104314,I104335,I104317,I104332,I104326,I104323,I104338,I104314,I104320,I104329,I104317,I104384,I104387,I104390,I104393,I104396,I104399,I104402,I104405,I104408,I2224,I2231);
PAT_9 I_1446 (I104405,I104387,I104387,I104384,I104408,I104390,I104393,I104384,I104396,I104402,I104399,I104454,I104457,I104460,I104463,I104466,I104469,I104472,I104475,I104478,I2224,I2231);
PAT_8 I_1447 (I104475,I104463,I104472,I104454,I104457,I104469,I104478,I104457,I104460,I104466,I104454,I104524,I104527,I104530,I104533,I104536,I104539,I104542,I104545,I104548,I2224,I2231);
PAT_2 I_1448 (I104527,I104542,I104548,I104524,I104536,I104539,I104527,I104545,I104530,I104533,I104524,I104594,I104597,I104600,I104603,I104606,I104609,I104612,I104615,I104618,I2224,I2231);
PAT_7 I_1449 (I104618,I104594,I104600,I104597,I104597,I104606,I104609,I104594,I104612,I104615,I104603,I104664,I104667,I104670,I104673,I104676,I104679,I104682,I104685,I104688,I2224,I2231);
PAT_5 I_1450 (I104670,I104664,I104673,I104682,I104676,I104688,I104685,I104667,I104679,I104667,I104664,I104734,I104737,I104740,I104743,I104746,I104749,I104752,I104755,I104758,I104761,I2224,I2231);
PAT_8 I_1451 (I104734,I104761,I104752,I104749,I104743,I104734,I104746,I104758,I104737,I104755,I104740,I104807,I104810,I104813,I104816,I104819,I104822,I104825,I104828,I104831,I2224,I2231);
PAT_9 I_1452 (I104810,I104819,I104810,I104807,I104822,I104813,I104828,I104816,I104825,I104807,I104831,I104877,I104880,I104883,I104886,I104889,I104892,I104895,I104898,I104901,I2224,I2231);
PAT_4 I_1453 (I104877,I104901,I104895,I104883,I104880,I104898,I104880,I104877,I104892,I104886,I104889,I104947,I104950,I104953,I104956,I104959,I104962,I104965,I104968,I104971,I2224,I2231);
PAT_10 I_1454 (I104947,I104947,I104971,I104950,I104956,I104965,I104962,I104950,I104968,I104953,I104959,I105017,I105020,I105023,I105026,I105029,I105032,I105035,I105038,I2224,I2231);
PAT_15 I_1455 (I105032,I105035,I105023,I105029,I105017,I105017,I105023,I105038,I105026,I105020,I105020,I105084,I105087,I105090,I105093,I105096,I105099,I105102,I105105,I105108,I2224,I2231);
PAT_8 I_1456 (I105105,I105084,I105084,I105093,I105090,I105087,I105102,I105099,I105087,I105108,I105096,I105154,I105157,I105160,I105163,I105166,I105169,I105172,I105175,I105178,I2224,I2231);
PAT_13 I_1457 (I105166,I105175,I105157,I105178,I105160,I105154,I105154,I105163,I105172,I105169,I105157,I105224,I105227,I105230,I105233,I105236,I105239,I105242,I105245,I105248,I2224,I2231);
PAT_7 I_1458 (I105233,I105236,I105224,I105239,I105245,I105230,I105227,I105248,I105227,I105224,I105242,I105294,I105297,I105300,I105303,I105306,I105309,I105312,I105315,I105318,I2224,I2231);
PAT_10 I_1459 (I105294,I105297,I105294,I105315,I105303,I105306,I105297,I105318,I105309,I105300,I105312,I105364,I105367,I105370,I105373,I105376,I105379,I105382,I105385,I2224,I2231);
PAT_5 I_1460 (I105385,I105364,I105373,I105367,I105382,I105379,I105370,I105370,I105364,I105367,I105376,I105431,I105434,I105437,I105440,I105443,I105446,I105449,I105452,I105455,I105458,I2224,I2231);
PAT_12 I_1461 (I105458,I105446,I105431,I105455,I105434,I105431,I105437,I105440,I105443,I105449,I105452,I105504,I105507,I105510,I105513,I105516,I105519,I105522,I105525,I2224,I2231);
PAT_8 I_1462 (I105504,I105513,I105510,I105507,I105519,I105504,I105507,I105510,I105522,I105516,I105525,I105571,I105574,I105577,I105580,I105583,I105586,I105589,I105592,I105595,I2224,I2231);
PAT_0 I_1463 (I105571,I105589,I105580,I105595,I105583,I105571,I105574,I105577,I105586,I105574,I105592,I105641,I105644,I105647,I105650,I105653,I105656,I105659,I105662,I2224,I2231);
PAT_13 I_1464 (I105650,I105659,I105641,I105644,I105644,I105647,I105653,I105647,I105641,I105656,I105662,I105708,I105711,I105714,I105717,I105720,I105723,I105726,I105729,I105732,I2224,I2231);
PAT_5 I_1465 (I105720,I105711,I105717,I105729,I105711,I105732,I105714,I105723,I105708,I105708,I105726,I105778,I105781,I105784,I105787,I105790,I105793,I105796,I105799,I105802,I105805,I2224,I2231);
PAT_9 I_1466 (I105793,I105790,I105799,I105796,I105787,I105778,I105784,I105805,I105781,I105802,I105778,I105851,I105854,I105857,I105860,I105863,I105866,I105869,I105872,I105875,I2224,I2231);
PAT_4 I_1467 (I105851,I105875,I105869,I105857,I105854,I105872,I105854,I105851,I105866,I105860,I105863,I105921,I105924,I105927,I105930,I105933,I105936,I105939,I105942,I105945,I2224,I2231);
PAT_9 I_1468 (I105942,I105924,I105927,I105936,I105939,I105921,I105930,I105924,I105945,I105921,I105933,I105991,I105994,I105997,I106000,I106003,I106006,I106009,I106012,I106015,I2224,I2231);
PAT_13 I_1469 (I105991,I106012,I105994,I106009,I106003,I106000,I106015,I105991,I105997,I106006,I105994,I106061,I106064,I106067,I106070,I106073,I106076,I106079,I106082,I106085,I2224,I2231);
PAT_5 I_1470 (I106073,I106064,I106070,I106082,I106064,I106085,I106067,I106076,I106061,I106061,I106079,I106131,I106134,I106137,I106140,I106143,I106146,I106149,I106152,I106155,I106158,I2224,I2231);
PAT_12 I_1471 (I106158,I106146,I106131,I106155,I106134,I106131,I106137,I106140,I106143,I106149,I106152,I106204,I106207,I106210,I106213,I106216,I106219,I106222,I106225,I2224,I2231);
PAT_13 I_1472 (I106216,I106219,I106210,I106225,I106222,I106204,I106207,I106213,I106210,I106207,I106204,I106271,I106274,I106277,I106280,I106283,I106286,I106289,I106292,I106295,I2224,I2231);
PAT_4 I_1473 (I106280,I106283,I106295,I106277,I106292,I106289,I106274,I106286,I106274,I106271,I106271,I106341,I106344,I106347,I106350,I106353,I106356,I106359,I106362,I106365,I2224,I2231);
PAT_17 I_1474 (I106353,I106350,I106362,I106356,I106341,I106359,I106365,I106344,I106347,I106344,I106341,I106411,I106414,I106417,I106420,I106423,I106426,I106429,I106432,I106435,I106438,I2224,I2231);
PAT_13 I_1475 (I106429,I106432,I106417,I106411,I106423,I106435,I106414,I106426,I106411,I106438,I106420,I106484,I106487,I106490,I106493,I106496,I106499,I106502,I106505,I106508,I2224,I2231);
PAT_8 I_1476 (I106493,I106505,I106496,I106499,I106508,I106487,I106502,I106484,I106487,I106490,I106484,I106554,I106557,I106560,I106563,I106566,I106569,I106572,I106575,I106578,I2224,I2231);
PAT_6 I_1477 (I106557,I106554,I106560,I106572,I106569,I106563,I106566,I106554,I106575,I106557,I106578,I106624,I106627,I106630,I106633,I106636,I106639,I106642,I106645,I106648,I106651,I2224,I2231);
PAT_17 I_1478 (I106636,I106639,I106645,I106633,I106627,I106648,I106642,I106624,I106651,I106630,I106624,I106697,I106700,I106703,I106706,I106709,I106712,I106715,I106718,I106721,I106724,I2224,I2231);
PAT_12 I_1479 (I106721,I106703,I106697,I106715,I106709,I106718,I106700,I106724,I106697,I106706,I106712,I106770,I106773,I106776,I106779,I106782,I106785,I106788,I106791,I2224,I2231);
PAT_1 I_1480 (I106785,I106773,I106788,I106779,I106770,I106773,I106782,I106770,I106791,I106776,I106776,I106837,I106840,I106843,I106846,I106849,I106852,I106855,I106858,I106861,I2224,I2231);
PAT_9 I_1481 (I106852,I106858,I106843,I106861,I106840,I106855,I106840,I106846,I106837,I106849,I106837,I106907,I106910,I106913,I106916,I106919,I106922,I106925,I106928,I106931,I2224,I2231);
PAT_7 I_1482 (I106913,I106922,I106907,I106928,I106919,I106907,I106910,I106931,I106925,I106910,I106916,I106977,I106980,I106983,I106986,I106989,I106992,I106995,I106998,I107001,I2224,I2231);
PAT_9 I_1483 (I106998,I106986,I106995,I107001,I106983,I106989,I106980,I106992,I106977,I106977,I106980,I107047,I107050,I107053,I107056,I107059,I107062,I107065,I107068,I107071,I2224,I2231);
PAT_5 I_1484 (I107068,I107047,I107062,I107047,I107053,I107056,I107050,I107050,I107065,I107059,I107071,I107117,I107120,I107123,I107126,I107129,I107132,I107135,I107138,I107141,I107144,I2224,I2231);
PAT_1 I_1485 (I107132,I107120,I107138,I107117,I107123,I107117,I107126,I107141,I107135,I107144,I107129,I107190,I107193,I107196,I107199,I107202,I107205,I107208,I107211,I107214,I2224,I2231);
PAT_4 I_1486 (I107202,I107208,I107190,I107193,I107196,I107199,I107211,I107193,I107205,I107190,I107214,I107260,I107263,I107266,I107269,I107272,I107275,I107278,I107281,I107284,I2224,I2231);
PAT_13 I_1487 (I107275,I107269,I107281,I107266,I107272,I107260,I107284,I107278,I107263,I107260,I107263,I107330,I107333,I107336,I107339,I107342,I107345,I107348,I107351,I107354,I2224,I2231);
PAT_17 I_1488 (I107354,I107342,I107351,I107348,I107339,I107330,I107333,I107336,I107330,I107345,I107333,I107400,I107403,I107406,I107409,I107412,I107415,I107418,I107421,I107424,I107427,I2224,I2231);
PAT_2 I_1489 (I107400,I107418,I107415,I107400,I107409,I107424,I107421,I107406,I107427,I107412,I107403,I107473,I107476,I107479,I107482,I107485,I107488,I107491,I107494,I107497,I2224,I2231);
PAT_4 I_1490 (I107473,I107479,I107497,I107491,I107488,I107485,I107476,I107494,I107473,I107476,I107482,I107543,I107546,I107549,I107552,I107555,I107558,I107561,I107564,I107567,I2224,I2231);
PAT_17 I_1491 (I107555,I107552,I107564,I107558,I107543,I107561,I107567,I107546,I107549,I107546,I107543,I107613,I107616,I107619,I107622,I107625,I107628,I107631,I107634,I107637,I107640,I2224,I2231);
PAT_1 I_1492 (I107637,I107640,I107619,I107628,I107613,I107634,I107625,I107616,I107622,I107613,I107631,I107686,I107689,I107692,I107695,I107698,I107701,I107704,I107707,I107710,I2224,I2231);
PAT_2 I_1493 (I107686,I107692,I107686,I107701,I107689,I107689,I107695,I107698,I107704,I107710,I107707,I107756,I107759,I107762,I107765,I107768,I107771,I107774,I107777,I107780,I2224,I2231);
PAT_11 I_1494 (I107759,I107771,I107756,I107768,I107765,I107777,I107774,I107759,I107780,I107762,I107756,I107826,I107829,I107832,I107835,I107838,I107841,I107844,I107847,I107850,I107853,I2224,I2231);
PAT_4 I_1495 (I107832,I107853,I107826,I107844,I107835,I107826,I107847,I107829,I107838,I107850,I107841,I107899,I107902,I107905,I107908,I107911,I107914,I107917,I107920,I107923,I2224,I2231);
PAT_10 I_1496 (I107899,I107899,I107923,I107902,I107908,I107917,I107914,I107902,I107920,I107905,I107911,I107969,I107972,I107975,I107978,I107981,I107984,I107987,I107990,I2224,I2231);
PAT_5 I_1497 (I107990,I107969,I107978,I107972,I107987,I107984,I107975,I107975,I107969,I107972,I107981,I108036,I108039,I108042,I108045,I108048,I108051,I108054,I108057,I108060,I108063,I2224,I2231);
PAT_1 I_1498 (I108051,I108039,I108057,I108036,I108042,I108036,I108045,I108060,I108054,I108063,I108048,I108109,I108112,I108115,I108118,I108121,I108124,I108127,I108130,I108133,I2224,I2231);
PAT_17 I_1499 (I108121,I108109,I108130,I108133,I108112,I108115,I108112,I108124,I108118,I108109,I108127,I108179,I108182,I108185,I108188,I108191,I108194,I108197,I108200,I108203,I108206,I2224,I2231);
PAT_13 I_1500 (I108197,I108200,I108185,I108179,I108191,I108203,I108182,I108194,I108179,I108206,I108188,I108252,I108255,I108258,I108261,I108264,I108267,I108270,I108273,I108276,I2224,I2231);
PAT_2 I_1501 (I108270,I108264,I108261,I108267,I108252,I108276,I108255,I108273,I108252,I108258,I108255,I108322,I108325,I108328,I108331,I108334,I108337,I108340,I108343,I108346,I2224,I2231);
PAT_11 I_1502 (I108325,I108337,I108322,I108334,I108331,I108343,I108340,I108325,I108346,I108328,I108322,I108392,I108395,I108398,I108401,I108404,I108407,I108410,I108413,I108416,I108419,I2224,I2231);
PAT_8 I_1503 (I108401,I108407,I108410,I108416,I108413,I108404,I108392,I108392,I108419,I108395,I108398,I108465,I108468,I108471,I108474,I108477,I108480,I108483,I108486,I108489,I2224,I2231);
PAT_6 I_1504 (I108468,I108465,I108471,I108483,I108480,I108474,I108477,I108465,I108486,I108468,I108489,I108535,I108538,I108541,I108544,I108547,I108550,I108553,I108556,I108559,I108562,I2224,I2231);
PAT_13 I_1505 (I108559,I108541,I108556,I108535,I108538,I108544,I108562,I108547,I108553,I108535,I108550,I108608,I108611,I108614,I108617,I108620,I108623,I108626,I108629,I108632,I2224,I2231);
PAT_7 I_1506 (I108617,I108620,I108608,I108623,I108629,I108614,I108611,I108632,I108611,I108608,I108626,I108678,I108681,I108684,I108687,I108690,I108693,I108696,I108699,I108702,I2224,I2231);
PAT_17 I_1507 (I108690,I108684,I108693,I108678,I108696,I108699,I108681,I108702,I108687,I108681,I108678,I108748,I108751,I108754,I108757,I108760,I108763,I108766,I108769,I108772,I108775,I2224,I2231);
PAT_6 I_1508 (I108748,I108766,I108754,I108757,I108763,I108748,I108760,I108751,I108772,I108775,I108769,I108821,I108824,I108827,I108830,I108833,I108836,I108839,I108842,I108845,I108848,I2224,I2231);
PAT_5 I_1509 (I108842,I108821,I108827,I108830,I108836,I108839,I108821,I108845,I108824,I108833,I108848,I108894,I108897,I108900,I108903,I108906,I108909,I108912,I108915,I108918,I108921,I2224,I2231);
PAT_11 I_1510 (I108906,I108903,I108897,I108915,I108918,I108894,I108912,I108909,I108921,I108900,I108894,I108967,I108970,I108973,I108976,I108979,I108982,I108985,I108988,I108991,I108994,I2224,I2231);
PAT_2 I_1511 (I108967,I108991,I108979,I108973,I108982,I108985,I108970,I108994,I108988,I108976,I108967,I109040,I109043,I109046,I109049,I109052,I109055,I109058,I109061,I109064,I2224,I2231);
PAT_10 I_1512 (I109040,I109058,I109055,I109043,I109046,I109061,I109052,I109040,I109049,I109064,I109043,I109110,I109113,I109116,I109119,I109122,I109125,I109128,I109131,I2224,I2231);
PAT_8 I_1513 (I109131,I109122,I109113,I109110,I109119,I109110,I109125,I109113,I109128,I109116,I109116,I109177,I109180,I109183,I109186,I109189,I109192,I109195,I109198,I109201,I2224,I2231);
PAT_12 I_1514 (I109177,I109180,I109180,I109201,I109186,I109195,I109198,I109189,I109183,I109192,I109177,I109247,I109250,I109253,I109256,I109259,I109262,I109265,I109268,I2224,I2231);
PAT_5 I_1515 (I109256,I109262,I109268,I109253,I109253,I109247,I109265,I109247,I109250,I109250,I109259,I109314,I109317,I109320,I109323,I109326,I109329,I109332,I109335,I109338,I109341,I2224,I2231);
PAT_13 I_1516 (I109320,I109329,I109314,I109317,I109338,I109323,I109335,I109314,I109332,I109341,I109326,I109387,I109390,I109393,I109396,I109399,I109402,I109405,I109408,I109411,I2224,I2231);
PAT_11 I_1517 (I109387,I109399,I109402,I109393,I109390,I109411,I109390,I109408,I109396,I109387,I109405,I109457,I109460,I109463,I109466,I109469,I109472,I109475,I109478,I109481,I109484,I2224,I2231);
PAT_6 I_1518 (I109457,I109484,I109472,I109481,I109475,I109469,I109460,I109478,I109466,I109463,I109457,I109530,I109533,I109536,I109539,I109542,I109545,I109548,I109551,I109554,I109557,I2224,I2231);
PAT_11 I_1519 (I109530,I109545,I109530,I109542,I109539,I109557,I109554,I109551,I109548,I109533,I109536,I109603,I109606,I109609,I109612,I109615,I109618,I109621,I109624,I109627,I109630,I2224,I2231);
PAT_2 I_1520 (I109603,I109627,I109615,I109609,I109618,I109621,I109606,I109630,I109624,I109612,I109603,I109676,I109679,I109682,I109685,I109688,I109691,I109694,I109697,I109700,I2224,I2231);
PAT_7 I_1521 (I109700,I109676,I109682,I109679,I109679,I109688,I109691,I109676,I109694,I109697,I109685,I109746,I109749,I109752,I109755,I109758,I109761,I109764,I109767,I109770,I2224,I2231);
PAT_6 I_1522 (I109746,I109764,I109746,I109755,I109761,I109749,I109767,I109752,I109770,I109749,I109758,I109816,I109819,I109822,I109825,I109828,I109831,I109834,I109837,I109840,I109843,I2224,I2231);
PAT_11 I_1523 (I109816,I109831,I109816,I109828,I109825,I109843,I109840,I109837,I109834,I109819,I109822,I109889,I109892,I109895,I109898,I109901,I109904,I109907,I109910,I109913,I109916,I2224,I2231);
PAT_4 I_1524 (I109895,I109916,I109889,I109907,I109898,I109889,I109910,I109892,I109901,I109913,I109904,I109962,I109965,I109968,I109971,I109974,I109977,I109980,I109983,I109986,I2224,I2231);
PAT_7 I_1525 (I109977,I109971,I109968,I109962,I109974,I109980,I109965,I109965,I109983,I109986,I109962,I110032,I110035,I110038,I110041,I110044,I110047,I110050,I110053,I110056,I2224,I2231);
PAT_9 I_1526 (I110053,I110041,I110050,I110056,I110038,I110044,I110035,I110047,I110032,I110032,I110035,I110102,I110105,I110108,I110111,I110114,I110117,I110120,I110123,I110126,I2224,I2231);
PAT_1 I_1527 (I110102,I110120,I110102,I110114,I110105,I110111,I110117,I110123,I110126,I110108,I110105,I110172,I110175,I110178,I110181,I110184,I110187,I110190,I110193,I110196,I2224,I2231);
PAT_14 I_1528 (I110175,I110190,I110187,I110178,I110172,I110172,I110184,I110193,I110196,I110181,I110175,I110242,I110245,I110248,I110251,I110254,I110257,I110260,I110263,I110266,I2224,I2231);
PAT_2 I_1529 (I110260,I110266,I110251,I110242,I110245,I110245,I110257,I110242,I110263,I110248,I110254,I110312,I110315,I110318,I110321,I110324,I110327,I110330,I110333,I110336,I2224,I2231);
PAT_9 I_1530 (I110327,I110336,I110312,I110318,I110321,I110330,I110315,I110324,I110333,I110315,I110312,I110382,I110385,I110388,I110391,I110394,I110397,I110400,I110403,I110406,I2224,I2231);
PAT_5 I_1531 (I110403,I110382,I110397,I110382,I110388,I110391,I110385,I110385,I110400,I110394,I110406,I110452,I110455,I110458,I110461,I110464,I110467,I110470,I110473,I110476,I110479,I2224,I2231);
PAT_13 I_1532 (I110458,I110467,I110452,I110455,I110476,I110461,I110473,I110452,I110470,I110479,I110464,I110525,I110528,I110531,I110534,I110537,I110540,I110543,I110546,I110549,I2224,I2231);
PAT_11 I_1533 (I110525,I110537,I110540,I110531,I110528,I110549,I110528,I110546,I110534,I110525,I110543,I110595,I110598,I110601,I110604,I110607,I110610,I110613,I110616,I110619,I110622,I2224,I2231);
PAT_7 I_1534 (I110619,I110604,I110601,I110622,I110607,I110595,I110595,I110613,I110616,I110598,I110610,I110668,I110671,I110674,I110677,I110680,I110683,I110686,I110689,I110692,I2224,I2231);
PAT_13 I_1535 (I110674,I110692,I110683,I110668,I110680,I110668,I110689,I110671,I110677,I110671,I110686,I110738,I110741,I110744,I110747,I110750,I110753,I110756,I110759,I110762,I2224,I2231);
PAT_10 I_1536 (I110759,I110753,I110747,I110741,I110762,I110741,I110750,I110738,I110738,I110756,I110744,I110808,I110811,I110814,I110817,I110820,I110823,I110826,I110829,I2224,I2231);
PAT_9 I_1537 (I110820,I110808,I110811,I110814,I110808,I110814,I110817,I110811,I110829,I110823,I110826,I110875,I110878,I110881,I110884,I110887,I110890,I110893,I110896,I110899,I2224,I2231);
PAT_12 I_1538 (I110896,I110893,I110887,I110875,I110884,I110875,I110878,I110881,I110899,I110890,I110878,I110945,I110948,I110951,I110954,I110957,I110960,I110963,I110966,I2224,I2231);
PAT_1 I_1539 (I110960,I110948,I110963,I110954,I110945,I110948,I110957,I110945,I110966,I110951,I110951,I111012,I111015,I111018,I111021,I111024,I111027,I111030,I111033,I111036,I2224,I2231);
PAT_10 I_1540 (I111027,I111024,I111015,I111012,I111015,I111030,I111018,I111033,I111036,I111021,I111012,I111082,I111085,I111088,I111091,I111094,I111097,I111100,I111103,I2224,I2231);
PAT_9 I_1541 (I111094,I111082,I111085,I111088,I111082,I111088,I111091,I111085,I111103,I111097,I111100,I111149,I111152,I111155,I111158,I111161,I111164,I111167,I111170,I111173,I2224,I2231);
PAT_4 I_1542 (I111149,I111173,I111167,I111155,I111152,I111170,I111152,I111149,I111164,I111158,I111161,I111219,I111222,I111225,I111228,I111231,I111234,I111237,I111240,I111243,I2224,I2231);
PAT_13 I_1543 (I111234,I111228,I111240,I111225,I111231,I111219,I111243,I111237,I111222,I111219,I111222,I111289,I111292,I111295,I111298,I111301,I111304,I111307,I111310,I111313,I2224,I2231);
PAT_12 I_1544 (I111298,I111289,I111289,I111313,I111310,I111292,I111307,I111301,I111292,I111295,I111304,I111359,I111362,I111365,I111368,I111371,I111374,I111377,I111380,I2224,I2231);
PAT_8 I_1545 (I111359,I111368,I111365,I111362,I111374,I111359,I111362,I111365,I111377,I111371,I111380,I111426,I111429,I111432,I111435,I111438,I111441,I111444,I111447,I111450,I2224,I2231);
PAT_5 I_1546 (I111432,I111450,I111426,I111447,I111435,I111438,I111429,I111426,I111429,I111441,I111444,I111496,I111499,I111502,I111505,I111508,I111511,I111514,I111517,I111520,I111523,I2224,I2231);
PAT_9 I_1547 (I111511,I111508,I111517,I111514,I111505,I111496,I111502,I111523,I111499,I111520,I111496,I111569,I111572,I111575,I111578,I111581,I111584,I111587,I111590,I111593,I2224,I2231);
PAT_7 I_1548 (I111575,I111584,I111569,I111590,I111581,I111569,I111572,I111593,I111587,I111572,I111578,I111639,I111642,I111645,I111648,I111651,I111654,I111657,I111660,I111663,I2224,I2231);
PAT_6 I_1549 (I111639,I111657,I111639,I111648,I111654,I111642,I111660,I111645,I111663,I111642,I111651,I111709,I111712,I111715,I111718,I111721,I111724,I111727,I111730,I111733,I111736,I2224,I2231);
PAT_17 I_1550 (I111721,I111724,I111730,I111718,I111712,I111733,I111727,I111709,I111736,I111715,I111709,I111782,I111785,I111788,I111791,I111794,I111797,I111800,I111803,I111806,I111809,I2224,I2231);
PAT_2 I_1551 (I111782,I111800,I111797,I111782,I111791,I111806,I111803,I111788,I111809,I111794,I111785,I111855,I111858,I111861,I111864,I111867,I111870,I111873,I111876,I111879,I2224,I2231);
PAT_5 I_1552 (I111876,I111855,I111855,I111867,I111864,I111873,I111861,I111870,I111879,I111858,I111858,I111925,I111928,I111931,I111934,I111937,I111940,I111943,I111946,I111949,I111952,I2224,I2231);
PAT_1 I_1553 (I111940,I111928,I111946,I111925,I111931,I111925,I111934,I111949,I111943,I111952,I111937,I111998,I112001,I112004,I112007,I112010,I112013,I112016,I112019,I112022,I2224,I2231);
PAT_8 I_1554 (I112019,I112001,I112007,I111998,I112016,I112010,I112013,I111998,I112022,I112004,I112001,I112068,I112071,I112074,I112077,I112080,I112083,I112086,I112089,I112092,I2224,I2231);
PAT_5 I_1555 (I112074,I112092,I112068,I112089,I112077,I112080,I112071,I112068,I112071,I112083,I112086,I112138,I112141,I112144,I112147,I112150,I112153,I112156,I112159,I112162,I112165,I2224,I2231);
PAT_17 I_1556 (I112165,I112141,I112144,I112147,I112138,I112150,I112138,I112162,I112156,I112153,I112159,I112211,I112214,I112217,I112220,I112223,I112226,I112229,I112232,I112235,I112238,I2224,I2231);
PAT_9 I_1557 (I112232,I112214,I112220,I112235,I112217,I112229,I112211,I112223,I112211,I112238,I112226,I112284,I112287,I112290,I112293,I112296,I112299,I112302,I112305,I112308,I2224,I2231);
PAT_8 I_1558 (I112305,I112293,I112302,I112284,I112287,I112299,I112308,I112287,I112290,I112296,I112284,I112354,I112357,I112360,I112363,I112366,I112369,I112372,I112375,I112378,I2224,I2231);
PAT_5 I_1559 (I112360,I112378,I112354,I112375,I112363,I112366,I112357,I112354,I112357,I112369,I112372,I112424,I112427,I112430,I112433,I112436,I112439,I112442,I112445,I112448,I112451,I2224,I2231);
PAT_9 I_1560 (I112439,I112436,I112445,I112442,I112433,I112424,I112430,I112451,I112427,I112448,I112424,I112497,I112500,I112503,I112506,I112509,I112512,I112515,I112518,I112521,I2224,I2231);
PAT_17 I_1561 (I112500,I112506,I112521,I112512,I112515,I112503,I112497,I112509,I112497,I112500,I112518,I112567,I112570,I112573,I112576,I112579,I112582,I112585,I112588,I112591,I112594,I2224,I2231);
PAT_7 I_1562 (I112585,I112576,I112582,I112570,I112579,I112588,I112594,I112567,I112591,I112573,I112567,I112640,I112643,I112646,I112649,I112652,I112655,I112658,I112661,I112664,I2224,I2231);
PAT_14 I_1563 (I112655,I112649,I112640,I112643,I112652,I112658,I112646,I112661,I112643,I112640,I112664,I112710,I112713,I112716,I112719,I112722,I112725,I112728,I112731,I112734,I2224,I2231);
PAT_9 I_1564 (I112719,I112731,I112710,I112728,I112713,I112716,I112734,I112713,I112722,I112710,I112725,I112780,I112783,I112786,I112789,I112792,I112795,I112798,I112801,I112804,I2224,I2231);
PAT_14 I_1565 (I112789,I112780,I112804,I112786,I112783,I112780,I112795,I112801,I112792,I112783,I112798,I112850,I112853,I112856,I112859,I112862,I112865,I112868,I112871,I112874,I2224,I2231);
PAT_5 I_1566 (I112853,I112856,I112853,I112862,I112850,I112871,I112859,I112850,I112874,I112868,I112865,I112920,I112923,I112926,I112929,I112932,I112935,I112938,I112941,I112944,I112947,I2224,I2231);
PAT_8 I_1567 (I112920,I112947,I112938,I112935,I112929,I112920,I112932,I112944,I112923,I112941,I112926,I112993,I112996,I112999,I113002,I113005,I113008,I113011,I113014,I113017,I2224,I2231);
PAT_6 I_1568 (I112996,I112993,I112999,I113011,I113008,I113002,I113005,I112993,I113014,I112996,I113017,I113063,I113066,I113069,I113072,I113075,I113078,I113081,I113084,I113087,I113090,I2224,I2231);
PAT_13 I_1569 (I113087,I113069,I113084,I113063,I113066,I113072,I113090,I113075,I113081,I113063,I113078,I113136,I113139,I113142,I113145,I113148,I113151,I113154,I113157,I113160,I2224,I2231);
PAT_2 I_1570 (I113154,I113148,I113145,I113151,I113136,I113160,I113139,I113157,I113136,I113142,I113139,I113206,I113209,I113212,I113215,I113218,I113221,I113224,I113227,I113230,I2224,I2231);
PAT_6 I_1571 (I113230,I113206,I113221,I113218,I113224,I113215,I113209,I113227,I113206,I113212,I113209,I113276,I113279,I113282,I113285,I113288,I113291,I113294,I113297,I113300,I113303,I2224,I2231);
PAT_10 I_1572 (I113276,I113291,I113294,I113285,I113276,I113300,I113303,I113279,I113288,I113282,I113297,I113349,I113352,I113355,I113358,I113361,I113364,I113367,I113370,I2224,I2231);
PAT_9 I_1573 (I113361,I113349,I113352,I113355,I113349,I113355,I113358,I113352,I113370,I113364,I113367,I113416,I113419,I113422,I113425,I113428,I113431,I113434,I113437,I113440,I2224,I2231);
PAT_11 I_1574 (I113428,I113434,I113440,I113437,I113425,I113419,I113419,I113416,I113431,I113416,I113422,I113486,I113489,I113492,I113495,I113498,I113501,I113504,I113507,I113510,I113513,I2224,I2231);
PAT_17 I_1575 (I113498,I113489,I113513,I113486,I113495,I113507,I113504,I113501,I113486,I113510,I113492,I113559,I113562,I113565,I113568,I113571,I113574,I113577,I113580,I113583,I113586,I2224,I2231);
PAT_11 I_1576 (I113571,I113580,I113586,I113562,I113559,I113577,I113568,I113574,I113565,I113583,I113559,I113632,I113635,I113638,I113641,I113644,I113647,I113650,I113653,I113656,I113659,I2224,I2231);
PAT_9 I_1577 (I113638,I113650,I113641,I113653,I113632,I113635,I113644,I113632,I113647,I113656,I113659,I113705,I113708,I113711,I113714,I113717,I113720,I113723,I113726,I113729,I2224,I2231);
PAT_8 I_1578 (I113726,I113714,I113723,I113705,I113708,I113720,I113729,I113708,I113711,I113717,I113705,I113775,I113778,I113781,I113784,I113787,I113790,I113793,I113796,I113799,I2224,I2231);
PAT_6 I_1579 (I113778,I113775,I113781,I113793,I113790,I113784,I113787,I113775,I113796,I113778,I113799,I113845,I113848,I113851,I113854,I113857,I113860,I113863,I113866,I113869,I113872,I2224,I2231);
PAT_9 I_1580 (I113845,I113872,I113869,I113851,I113857,I113848,I113860,I113845,I113863,I113854,I113866,I113918,I113921,I113924,I113927,I113930,I113933,I113936,I113939,I113942,I2224,I2231);
PAT_5 I_1581 (I113939,I113918,I113933,I113918,I113924,I113927,I113921,I113921,I113936,I113930,I113942,I113988,I113991,I113994,I113997,I114000,I114003,I114006,I114009,I114012,I114015,I2224,I2231);
PAT_6 I_1582 (I114006,I114000,I113988,I113994,I113991,I113997,I114003,I113988,I114012,I114009,I114015,I114061,I114064,I114067,I114070,I114073,I114076,I114079,I114082,I114085,I114088,I2224,I2231);
PAT_10 I_1583 (I114061,I114076,I114079,I114070,I114061,I114085,I114088,I114064,I114073,I114067,I114082,I114134,I114137,I114140,I114143,I114146,I114149,I114152,I114155,I2224,I2231);
PAT_12 I_1584 (I114140,I114134,I114134,I114146,I114149,I114137,I114137,I114152,I114155,I114140,I114143,I114201,I114204,I114207,I114210,I114213,I114216,I114219,I114222,I2224,I2231);
PAT_4 I_1585 (I114207,I114204,I114219,I114222,I114216,I114210,I114201,I114201,I114207,I114213,I114204,I114268,I114271,I114274,I114277,I114280,I114283,I114286,I114289,I114292,I2224,I2231);
PAT_6 I_1586 (I114268,I114274,I114271,I114283,I114286,I114280,I114292,I114289,I114268,I114277,I114271,I114338,I114341,I114344,I114347,I114350,I114353,I114356,I114359,I114362,I114365,I2224,I2231);
PAT_17 I_1587 (I114350,I114353,I114359,I114347,I114341,I114362,I114356,I114338,I114365,I114344,I114338,I114411,I114414,I114417,I114420,I114423,I114426,I114429,I114432,I114435,I114438,I2224,I2231);
PAT_11 I_1588 (I114423,I114432,I114438,I114414,I114411,I114429,I114420,I114426,I114417,I114435,I114411,I114484,I114487,I114490,I114493,I114496,I114499,I114502,I114505,I114508,I114511,I2224,I2231);
PAT_9 I_1589 (I114490,I114502,I114493,I114505,I114484,I114487,I114496,I114484,I114499,I114508,I114511,I114557,I114560,I114563,I114566,I114569,I114572,I114575,I114578,I114581,I2224,I2231);
PAT_4 I_1590 (I114557,I114581,I114575,I114563,I114560,I114578,I114560,I114557,I114572,I114566,I114569,I114627,I114630,I114633,I114636,I114639,I114642,I114645,I114648,I114651,I2224,I2231);
PAT_9 I_1591 (I114648,I114630,I114633,I114642,I114645,I114627,I114636,I114630,I114651,I114627,I114639,I114697,I114700,I114703,I114706,I114709,I114712,I114715,I114718,I114721,I2224,I2231);
PAT_12 I_1592 (I114718,I114715,I114709,I114697,I114706,I114697,I114700,I114703,I114721,I114712,I114700,I114767,I114770,I114773,I114776,I114779,I114782,I114785,I114788,I2224,I2231);
PAT_13 I_1593 (I114779,I114782,I114773,I114788,I114785,I114767,I114770,I114776,I114773,I114770,I114767,I114834,I114837,I114840,I114843,I114846,I114849,I114852,I114855,I114858,I2224,I2231);
PAT_2 I_1594 (I114852,I114846,I114843,I114849,I114834,I114858,I114837,I114855,I114834,I114840,I114837,I114904,I114907,I114910,I114913,I114916,I114919,I114922,I114925,I114928,I2224,I2231);
PAT_9 I_1595 (I114919,I114928,I114904,I114910,I114913,I114922,I114907,I114916,I114925,I114907,I114904,I114974,I114977,I114980,I114983,I114986,I114989,I114992,I114995,I114998,I2224,I2231);
PAT_17 I_1596 (I114977,I114983,I114998,I114989,I114992,I114980,I114974,I114986,I114974,I114977,I114995,I115044,I115047,I115050,I115053,I115056,I115059,I115062,I115065,I115068,I115071,I2224,I2231);
PAT_11 I_1597 (I115056,I115065,I115071,I115047,I115044,I115062,I115053,I115059,I115050,I115068,I115044,I115117,I115120,I115123,I115126,I115129,I115132,I115135,I115138,I115141,I115144,I2224,I2231);
PAT_7 I_1598 (I115141,I115126,I115123,I115144,I115129,I115117,I115117,I115135,I115138,I115120,I115132,I115190,I115193,I115196,I115199,I115202,I115205,I115208,I115211,I115214,I2224,I2231);
PAT_9 I_1599 (I115211,I115199,I115208,I115214,I115196,I115202,I115193,I115205,I115190,I115190,I115193,I115260,I115263,I115266,I115269,I115272,I115275,I115278,I115281,I115284,I2224,I2231);
PAT_5 I_1600 (I115281,I115260,I115275,I115260,I115266,I115269,I115263,I115263,I115278,I115272,I115284,I115330,I115333,I115336,I115339,I115342,I115345,I115348,I115351,I115354,I115357,I2224,I2231);
PAT_0 I_1601 (I115351,I115330,I115357,I115354,I115330,I115348,I115342,I115333,I115339,I115345,I115336,I115403,I115406,I115409,I115412,I115415,I115418,I115421,I115424,I2224,I2231);
PAT_1 I_1602 (I115406,I115403,I115403,I115421,I115406,I115415,I115409,I115418,I115412,I115424,I115409,I115470,I115473,I115476,I115479,I115482,I115485,I115488,I115491,I115494,I2224,I2231);
PAT_17 I_1603 (I115482,I115470,I115491,I115494,I115473,I115476,I115473,I115485,I115479,I115470,I115488,I115540,I115543,I115546,I115549,I115552,I115555,I115558,I115561,I115564,I115567,I2224,I2231);
PAT_13 I_1604 (I115558,I115561,I115546,I115540,I115552,I115564,I115543,I115555,I115540,I115567,I115549,I115613,I115616,I115619,I115622,I115625,I115628,I115631,I115634,I115637,I2224,I2231);
PAT_5 I_1605 (I115625,I115616,I115622,I115634,I115616,I115637,I115619,I115628,I115613,I115613,I115631,I115683,I115686,I115689,I115692,I115695,I115698,I115701,I115704,I115707,I115710,I2224,I2231);
PAT_7 I_1606 (I115701,I115704,I115710,I115707,I115692,I115689,I115683,I115695,I115683,I115686,I115698,I115756,I115759,I115762,I115765,I115768,I115771,I115774,I115777,I115780,I2224,I2231);
PAT_9 I_1607 (I115777,I115765,I115774,I115780,I115762,I115768,I115759,I115771,I115756,I115756,I115759,I115826,I115829,I115832,I115835,I115838,I115841,I115844,I115847,I115850,I2224,I2231);
PAT_5 I_1608 (I115847,I115826,I115841,I115826,I115832,I115835,I115829,I115829,I115844,I115838,I115850,I115896,I115899,I115902,I115905,I115908,I115911,I115914,I115917,I115920,I115923,I2224,I2231);
PAT_17 I_1609 (I115923,I115899,I115902,I115905,I115896,I115908,I115896,I115920,I115914,I115911,I115917,I115969,I115972,I115975,I115978,I115981,I115984,I115987,I115990,I115993,I115996,I2224,I2231);
PAT_2 I_1610 (I115969,I115987,I115984,I115969,I115978,I115993,I115990,I115975,I115996,I115981,I115972,I116042,I116045,I116048,I116051,I116054,I116057,I116060,I116063,I116066,I2224,I2231);
PAT_9 I_1611 (I116057,I116066,I116042,I116048,I116051,I116060,I116045,I116054,I116063,I116045,I116042,I116112,I116115,I116118,I116121,I116124,I116127,I116130,I116133,I116136,I2224,I2231);
PAT_15 I_1612 (I116124,I116133,I116136,I116115,I116130,I116118,I116121,I116112,I116127,I116112,I116115,I116182,I116185,I116188,I116191,I116194,I116197,I116200,I116203,I116206,I2224,I2231);
PAT_12 I_1613 (I116200,I116203,I116206,I116194,I116191,I116185,I116182,I116197,I116188,I116182,I116185,I116252,I116255,I116258,I116261,I116264,I116267,I116270,I116273,I2224,I2231);
PAT_6 I_1614 (I116261,I116255,I116273,I116258,I116255,I116258,I116267,I116252,I116270,I116252,I116264,I116319,I116322,I116325,I116328,I116331,I116334,I116337,I116340,I116343,I116346,I2224,I2231);
PAT_11 I_1615 (I116319,I116334,I116319,I116331,I116328,I116346,I116343,I116340,I116337,I116322,I116325,I116392,I116395,I116398,I116401,I116404,I116407,I116410,I116413,I116416,I116419,I2224,I2231);
PAT_2 I_1616 (I116392,I116416,I116404,I116398,I116407,I116410,I116395,I116419,I116413,I116401,I116392,I116465,I116468,I116471,I116474,I116477,I116480,I116483,I116486,I116489,I2224,I2231);
PAT_9 I_1617 (I116480,I116489,I116465,I116471,I116474,I116483,I116468,I116477,I116486,I116468,I116465,I116535,I116538,I116541,I116544,I116547,I116550,I116553,I116556,I116559,I2224,I2231);
PAT_4 I_1618 (I116535,I116559,I116553,I116541,I116538,I116556,I116538,I116535,I116550,I116544,I116547,I116605,I116608,I116611,I116614,I116617,I116620,I116623,I116626,I116629,I2224,I2231);
PAT_2 I_1619 (I116614,I116608,I116608,I116629,I116605,I116623,I116620,I116611,I116605,I116617,I116626,I116675,I116678,I116681,I116684,I116687,I116690,I116693,I116696,I116699,I2224,I2231);
PAT_1 I_1620 (I116687,I116675,I116681,I116684,I116675,I116690,I116699,I116678,I116693,I116678,I116696,I116745,I116748,I116751,I116754,I116757,I116760,I116763,I116766,I116769,I2224,I2231);
PAT_13 I_1621 (I116754,I116763,I116769,I116745,I116760,I116757,I116766,I116751,I116748,I116745,I116748,I116815,I116818,I116821,I116824,I116827,I116830,I116833,I116836,I116839,I2224,I2231);
PAT_2 I_1622 (I116833,I116827,I116824,I116830,I116815,I116839,I116818,I116836,I116815,I116821,I116818,I116885,I116888,I116891,I116894,I116897,I116900,I116903,I116906,I116909,I2224,I2231);
PAT_6 I_1623 (I116909,I116885,I116900,I116897,I116903,I116894,I116888,I116906,I116885,I116891,I116888,I116955,I116958,I116961,I116964,I116967,I116970,I116973,I116976,I116979,I116982,I2224,I2231);
PAT_9 I_1624 (I116955,I116982,I116979,I116961,I116967,I116958,I116970,I116955,I116973,I116964,I116976,I117028,I117031,I117034,I117037,I117040,I117043,I117046,I117049,I117052,I2224,I2231);
PAT_5 I_1625 (I117049,I117028,I117043,I117028,I117034,I117037,I117031,I117031,I117046,I117040,I117052,I117098,I117101,I117104,I117107,I117110,I117113,I117116,I117119,I117122,I117125,I2224,I2231);
PAT_13 I_1626 (I117104,I117113,I117098,I117101,I117122,I117107,I117119,I117098,I117116,I117125,I117110,I117171,I117174,I117177,I117180,I117183,I117186,I117189,I117192,I117195,I2224,I2231);
PAT_12 I_1627 (I117180,I117171,I117171,I117195,I117192,I117174,I117189,I117183,I117174,I117177,I117186,I117241,I117244,I117247,I117250,I117253,I117256,I117259,I117262,I2224,I2231);
PAT_11 I_1628 (I117247,I117250,I117247,I117259,I117262,I117256,I117244,I117253,I117241,I117244,I117241,I117308,I117311,I117314,I117317,I117320,I117323,I117326,I117329,I117332,I117335,I2224,I2231);
PAT_10 I_1629 (I117323,I117329,I117320,I117314,I117332,I117317,I117335,I117326,I117308,I117311,I117308,I117381,I117384,I117387,I117390,I117393,I117396,I117399,I117402,I2224,I2231);
PAT_14 I_1630 (I117381,I117402,I117387,I117396,I117393,I117399,I117390,I117384,I117384,I117387,I117381,I117448,I117451,I117454,I117457,I117460,I117463,I117466,I117469,I117472,I2224,I2231);
PAT_13 I_1631 (I117457,I117472,I117451,I117460,I117448,I117451,I117466,I117454,I117448,I117469,I117463,I117518,I117521,I117524,I117527,I117530,I117533,I117536,I117539,I117542,I2224,I2231);
PAT_5 I_1632 (I117530,I117521,I117527,I117539,I117521,I117542,I117524,I117533,I117518,I117518,I117536,I117588,I117591,I117594,I117597,I117600,I117603,I117606,I117609,I117612,I117615,I2224,I2231);
PAT_11 I_1633 (I117600,I117597,I117591,I117609,I117612,I117588,I117606,I117603,I117615,I117594,I117588,I117661,I117664,I117667,I117670,I117673,I117676,I117679,I117682,I117685,I117688,I2224,I2231);
PAT_13 I_1634 (I117661,I117664,I117673,I117685,I117688,I117676,I117682,I117670,I117679,I117667,I117661,I117734,I117737,I117740,I117743,I117746,I117749,I117752,I117755,I117758,I2224,I2231);
PAT_4 I_1635 (I117743,I117746,I117758,I117740,I117755,I117752,I117737,I117749,I117737,I117734,I117734,I117804,I117807,I117810,I117813,I117816,I117819,I117822,I117825,I117828,I2224,I2231);
PAT_2 I_1636 (I117813,I117807,I117807,I117828,I117804,I117822,I117819,I117810,I117804,I117816,I117825,I117874,I117877,I117880,I117883,I117886,I117889,I117892,I117895,I117898,I2224,I2231);
PAT_5 I_1637 (I117895,I117874,I117874,I117886,I117883,I117892,I117880,I117889,I117898,I117877,I117877,I117944,I117947,I117950,I117953,I117956,I117959,I117962,I117965,I117968,I117971,I2224,I2231);
PAT_15 I_1638 (I117962,I117947,I117944,I117944,I117959,I117956,I117968,I117953,I117965,I117950,I117971,I118017,I118020,I118023,I118026,I118029,I118032,I118035,I118038,I118041,I2224,I2231);
PAT_10 I_1639 (I118020,I118029,I118023,I118017,I118038,I118041,I118026,I118017,I118020,I118035,I118032,I118087,I118090,I118093,I118096,I118099,I118102,I118105,I118108,I2224,I2231);
PAT_2 I_1640 (I118099,I118102,I118093,I118105,I118090,I118087,I118087,I118093,I118108,I118096,I118090,I118154,I118157,I118160,I118163,I118166,I118169,I118172,I118175,I118178,I2224,I2231);
PAT_17 I_1641 (I118154,I118154,I118166,I118157,I118160,I118172,I118169,I118178,I118157,I118163,I118175,I118224,I118227,I118230,I118233,I118236,I118239,I118242,I118245,I118248,I118251,I2224,I2231);
PAT_13 I_1642 (I118242,I118245,I118230,I118224,I118236,I118248,I118227,I118239,I118224,I118251,I118233,I118297,I118300,I118303,I118306,I118309,I118312,I118315,I118318,I118321,I2224,I2231);
PAT_2 I_1643 (I118315,I118309,I118306,I118312,I118297,I118321,I118300,I118318,I118297,I118303,I118300,I118367,I118370,I118373,I118376,I118379,I118382,I118385,I118388,I118391,I2224,I2231);
PAT_4 I_1644 (I118367,I118373,I118391,I118385,I118382,I118379,I118370,I118388,I118367,I118370,I118376,I118437,I118440,I118443,I118446,I118449,I118452,I118455,I118458,I118461,I2224,I2231);
PAT_7 I_1645 (I118452,I118446,I118443,I118437,I118449,I118455,I118440,I118440,I118458,I118461,I118437,I118507,I118510,I118513,I118516,I118519,I118522,I118525,I118528,I118531,I2224,I2231);
PAT_5 I_1646 (I118513,I118507,I118516,I118525,I118519,I118531,I118528,I118510,I118522,I118510,I118507,I118577,I118580,I118583,I118586,I118589,I118592,I118595,I118598,I118601,I118604,I2224,I2231);
PAT_9 I_1647 (I118592,I118589,I118598,I118595,I118586,I118577,I118583,I118604,I118580,I118601,I118577,I118650,I118653,I118656,I118659,I118662,I118665,I118668,I118671,I118674,I2224,I2231);
PAT_10 I_1648 (I118671,I118668,I118656,I118653,I118674,I118659,I118665,I118653,I118650,I118650,I118662,I118720,I118723,I118726,I118729,I118732,I118735,I118738,I118741,I2224,I2231);
PAT_2 I_1649 (I118732,I118735,I118726,I118738,I118723,I118720,I118720,I118726,I118741,I118729,I118723,I118787,I118790,I118793,I118796,I118799,I118802,I118805,I118808,I118811,I2224,I2231);
PAT_9 I_1650 (I118802,I118811,I118787,I118793,I118796,I118805,I118790,I118799,I118808,I118790,I118787,I118857,I118860,I118863,I118866,I118869,I118872,I118875,I118878,I118881,I2224,I2231);
PAT_10 I_1651 (I118878,I118875,I118863,I118860,I118881,I118866,I118872,I118860,I118857,I118857,I118869,I118927,I118930,I118933,I118936,I118939,I118942,I118945,I118948,I2224,I2231);
PAT_15 I_1652 (I118942,I118945,I118933,I118939,I118927,I118927,I118933,I118948,I118936,I118930,I118930,I118994,I118997,I119000,I119003,I119006,I119009,I119012,I119015,I119018,I2224,I2231);
PAT_1 I_1653 (I119000,I118997,I118997,I118994,I118994,I119003,I119018,I119012,I119006,I119009,I119015,I119064,I119067,I119070,I119073,I119076,I119079,I119082,I119085,I119088,I2224,I2231);
PAT_6 I_1654 (I119073,I119064,I119067,I119070,I119085,I119088,I119082,I119064,I119079,I119076,I119067,I119134,I119137,I119140,I119143,I119146,I119149,I119152,I119155,I119158,I119161,I2224,I2231);
PAT_13 I_1655 (I119158,I119140,I119155,I119134,I119137,I119143,I119161,I119146,I119152,I119134,I119149,I119207,I119210,I119213,I119216,I119219,I119222,I119225,I119228,I119231,I2224,I2231);
PAT_5 I_1656 (I119219,I119210,I119216,I119228,I119210,I119231,I119213,I119222,I119207,I119207,I119225,I119277,I119280,I119283,I119286,I119289,I119292,I119295,I119298,I119301,I119304,I2224,I2231);
PAT_15 I_1657 (I119295,I119280,I119277,I119277,I119292,I119289,I119301,I119286,I119298,I119283,I119304,I119350,I119353,I119356,I119359,I119362,I119365,I119368,I119371,I119374,I2224,I2231);
PAT_8 I_1658 (I119371,I119350,I119350,I119359,I119356,I119353,I119368,I119365,I119353,I119374,I119362,I119420,I119423,I119426,I119429,I119432,I119435,I119438,I119441,I119444,I2224,I2231);
PAT_13 I_1659 (I119432,I119441,I119423,I119444,I119426,I119420,I119420,I119429,I119438,I119435,I119423,I119490,I119493,I119496,I119499,I119502,I119505,I119508,I119511,I119514,I2224,I2231);
PAT_2 I_1660 (I119508,I119502,I119499,I119505,I119490,I119514,I119493,I119511,I119490,I119496,I119493,I119560,I119563,I119566,I119569,I119572,I119575,I119578,I119581,I119584,I2224,I2231);
PAT_17 I_1661 (I119560,I119560,I119572,I119563,I119566,I119578,I119575,I119584,I119563,I119569,I119581,I119630,I119633,I119636,I119639,I119642,I119645,I119648,I119651,I119654,I119657,I2224,I2231);
PAT_13 I_1662 (I119648,I119651,I119636,I119630,I119642,I119654,I119633,I119645,I119630,I119657,I119639,I119703,I119706,I119709,I119712,I119715,I119718,I119721,I119724,I119727,I2224,I2231);
PAT_5 I_1663 (I119715,I119706,I119712,I119724,I119706,I119727,I119709,I119718,I119703,I119703,I119721,I119773,I119776,I119779,I119782,I119785,I119788,I119791,I119794,I119797,I119800,I2224,I2231);
PAT_6 I_1664 (I119791,I119785,I119773,I119779,I119776,I119782,I119788,I119773,I119797,I119794,I119800,I119846,I119849,I119852,I119855,I119858,I119861,I119864,I119867,I119870,I119873,I2224,I2231);
PAT_11 I_1665 (I119846,I119861,I119846,I119858,I119855,I119873,I119870,I119867,I119864,I119849,I119852,I119919,I119922,I119925,I119928,I119931,I119934,I119937,I119940,I119943,I119946,I2224,I2231);
PAT_6 I_1666 (I119919,I119946,I119934,I119943,I119937,I119931,I119922,I119940,I119928,I119925,I119919,I119992,I119995,I119998,I120001,I120004,I120007,I120010,I120013,I120016,I120019,I2224,I2231);
PAT_15 I_1667 (I120010,I120001,I120013,I120016,I120007,I120019,I119992,I119998,I119992,I119995,I120004,I120065,I120068,I120071,I120074,I120077,I120080,I120083,I120086,I120089,I2224,I2231);
PAT_1 I_1668 (I120071,I120068,I120068,I120065,I120065,I120074,I120089,I120083,I120077,I120080,I120086,I120135,I120138,I120141,I120144,I120147,I120150,I120153,I120156,I120159,I2224,I2231);
PAT_6 I_1669 (I120144,I120135,I120138,I120141,I120156,I120159,I120153,I120135,I120150,I120147,I120138,I120205,I120208,I120211,I120214,I120217,I120220,I120223,I120226,I120229,I120232,I2224,I2231);
PAT_5 I_1670 (I120226,I120205,I120211,I120214,I120220,I120223,I120205,I120229,I120208,I120217,I120232,I120278,I120281,I120284,I120287,I120290,I120293,I120296,I120299,I120302,I120305,I2224,I2231);
PAT_17 I_1671 (I120305,I120281,I120284,I120287,I120278,I120290,I120278,I120302,I120296,I120293,I120299,I120351,I120354,I120357,I120360,I120363,I120366,I120369,I120372,I120375,I120378,I2224,I2231);
PAT_9 I_1672 (I120372,I120354,I120360,I120375,I120357,I120369,I120351,I120363,I120351,I120378,I120366,I120424,I120427,I120430,I120433,I120436,I120439,I120442,I120445,I120448,I2224,I2231);
PAT_5 I_1673 (I120445,I120424,I120439,I120424,I120430,I120433,I120427,I120427,I120442,I120436,I120448,I120494,I120497,I120500,I120503,I120506,I120509,I120512,I120515,I120518,I120521,I2224,I2231);
PAT_4 I_1674 (I1689,I1801,I1513,I1937,I1793,I2137,I1921,I2217,I2201,I1665,I2161,I120567,I120570,I120573,I120576,I120579,I120582,I120585,I120588,I120591,I2224,I2231);
PAT_17 I_1675 (I120579,I120576,I120588,I120582,I120567,I120585,I120591,I120570,I120573,I120570,I120567,I120637,I120640,I120643,I120646,I120649,I120652,I120655,I120658,I120661,I120664,I2224,I2231);
PAT_6 I_1676 (I120637,I120655,I120643,I120646,I120652,I120637,I120649,I120640,I120661,I120664,I120658,I120710,I120713,I120716,I120719,I120722,I120725,I120728,I120731,I120734,I120737,I2224,I2231);
PAT_9 I_1677 (I120710,I120737,I120734,I120716,I120722,I120713,I120725,I120710,I120728,I120719,I120731,I120783,I120786,I120789,I120792,I120795,I120798,I120801,I120804,I120807,I2224,I2231);
PAT_13 I_1678 (I120783,I120804,I120786,I120801,I120795,I120792,I120807,I120783,I120789,I120798,I120786,I120853,I120856,I120859,I120862,I120865,I120868,I120871,I120874,I120877,I2224,I2231);
PAT_17 I_1679 (I120877,I120865,I120874,I120871,I120862,I120853,I120856,I120859,I120853,I120868,I120856,I120923,I120926,I120929,I120932,I120935,I120938,I120941,I120944,I120947,I120950,I2224,I2231);
PAT_14 I_1680 (I120926,I120941,I120923,I120947,I120932,I120938,I120923,I120944,I120929,I120950,I120935,I120996,I120999,I121002,I121005,I121008,I121011,I121014,I121017,I121020,I2224,I2231);
PAT_5 I_1681 (I120999,I121002,I120999,I121008,I120996,I121017,I121005,I120996,I121020,I121014,I121011,I121066,I121069,I121072,I121075,I121078,I121081,I121084,I121087,I121090,I121093,I2224,I2231);
PAT_2 I_1682 (I121081,I121066,I121078,I121072,I121087,I121069,I121084,I121075,I121090,I121093,I121066,I121139,I121142,I121145,I121148,I121151,I121154,I121157,I121160,I121163,I2224,I2231);
PAT_11 I_1683 (I121142,I121154,I121139,I121151,I121148,I121160,I121157,I121142,I121163,I121145,I121139,I121209,I121212,I121215,I121218,I121221,I121224,I121227,I121230,I121233,I121236,I2224,I2231);
PAT_8 I_1684 (I121218,I121224,I121227,I121233,I121230,I121221,I121209,I121209,I121236,I121212,I121215,I121282,I121285,I121288,I121291,I121294,I121297,I121300,I121303,I121306,I2224,I2231);
PAT_13 I_1685 (I121294,I121303,I121285,I121306,I121288,I121282,I121282,I121291,I121300,I121297,I121285,I121352,I121355,I121358,I121361,I121364,I121367,I121370,I121373,I121376,I2224,I2231);
PAT_17 I_1686 (I121376,I121364,I121373,I121370,I121361,I121352,I121355,I121358,I121352,I121367,I121355,I121422,I121425,I121428,I121431,I121434,I121437,I121440,I121443,I121446,I121449,I2224,I2231);
PAT_9 I_1687 (I121443,I121425,I121431,I121446,I121428,I121440,I121422,I121434,I121422,I121449,I121437,I121495,I121498,I121501,I121504,I121507,I121510,I121513,I121516,I121519,I2224,I2231);
PAT_4 I_1688 (I121495,I121519,I121513,I121501,I121498,I121516,I121498,I121495,I121510,I121504,I121507,I121565,I121568,I121571,I121574,I121577,I121580,I121583,I121586,I121589,I2224,I2231);
PAT_17 I_1689 (I121577,I121574,I121586,I121580,I121565,I121583,I121589,I121568,I121571,I121568,I121565,I121635,I121638,I121641,I121644,I121647,I121650,I121653,I121656,I121659,I121662,I2224,I2231);
PAT_6 I_1690 (I121635,I121653,I121641,I121644,I121650,I121635,I121647,I121638,I121659,I121662,I121656,I121708,I121711,I121714,I121717,I121720,I121723,I121726,I121729,I121732,I121735,I2224,I2231);
PAT_11 I_1691 (I121708,I121723,I121708,I121720,I121717,I121735,I121732,I121729,I121726,I121711,I121714,I121781,I121784,I121787,I121790,I121793,I121796,I121799,I121802,I121805,I121808,I2224,I2231);
PAT_7 I_1692 (I121805,I121790,I121787,I121808,I121793,I121781,I121781,I121799,I121802,I121784,I121796,I121854,I121857,I121860,I121863,I121866,I121869,I121872,I121875,I121878,I2224,I2231);
PAT_8 I_1693 (I121860,I121872,I121854,I121857,I121863,I121854,I121878,I121875,I121866,I121869,I121857,I121924,I121927,I121930,I121933,I121936,I121939,I121942,I121945,I121948,I2224,I2231);
PAT_17 I_1694 (I121948,I121936,I121933,I121927,I121930,I121942,I121924,I121927,I121924,I121939,I121945,I121994,I121997,I122000,I122003,I122006,I122009,I122012,I122015,I122018,I122021,I2224,I2231);
PAT_5 I_1695 (I122006,I122000,I121997,I122018,I122003,I122009,I122012,I121994,I121994,I122015,I122021,I122067,I122070,I122073,I122076,I122079,I122082,I122085,I122088,I122091,I122094,I2224,I2231);
PAT_4 I_1696 (I122085,I122091,I122094,I122073,I122076,I122088,I122070,I122067,I122079,I122082,I122067,I122140,I122143,I122146,I122149,I122152,I122155,I122158,I122161,I122164,I2224,I2231);
PAT_12 I_1697 (I122140,I122143,I122161,I122164,I122155,I122146,I122152,I122149,I122140,I122158,I122143,I122210,I122213,I122216,I122219,I122222,I122225,I122228,I122231,I2224,I2231);
PAT_5 I_1698 (I122219,I122225,I122231,I122216,I122216,I122210,I122228,I122210,I122213,I122213,I122222,I122277,I122280,I122283,I122286,I122289,I122292,I122295,I122298,I122301,I122304,I2224,I2231);
PAT_2 I_1699 (I122292,I122277,I122289,I122283,I122298,I122280,I122295,I122286,I122301,I122304,I122277,I122350,I122353,I122356,I122359,I122362,I122365,I122368,I122371,I122374,I2224,I2231);
PAT_5 I_1700 (I122371,I122350,I122350,I122362,I122359,I122368,I122356,I122365,I122374,I122353,I122353,I122420,I122423,I122426,I122429,I122432,I122435,I122438,I122441,I122444,I122447,I2224,I2231);
PAT_12 I_1701 (I122447,I122435,I122420,I122444,I122423,I122420,I122426,I122429,I122432,I122438,I122441,I122493,I122496,I122499,I122502,I122505,I122508,I122511,I122514,I2224,I2231);
PAT_16 I_1702 (I122502,I122496,I122499,I122493,I122493,I122499,I122514,I122511,I122496,I122505,I122508,I122560,I122563,I122566,I122569,I122572,I122575,I122578,I122581,I122584,I122587,I2224,I2231);
PAT_2 I_1703 (I122569,I122575,I122563,I122587,I122560,I122578,I122572,I122566,I122584,I122560,I122581,I122633,I122636,I122639,I122642,I122645,I122648,I122651,I122654,I122657,I2224,I2231);
PAT_4 I_1704 (I122633,I122639,I122657,I122651,I122648,I122645,I122636,I122654,I122633,I122636,I122642,I122703,I122706,I122709,I122712,I122715,I122718,I122721,I122724,I122727,I2224,I2231);
PAT_12 I_1705 (I122703,I122706,I122724,I122727,I122718,I122709,I122715,I122712,I122703,I122721,I122706,I122773,I122776,I122779,I122782,I122785,I122788,I122791,I122794,I2224,I2231);
PAT_11 I_1706 (I122779,I122782,I122779,I122791,I122794,I122788,I122776,I122785,I122773,I122776,I122773,I122840,I122843,I122846,I122849,I122852,I122855,I122858,I122861,I122864,I122867,I2224,I2231);
PAT_15 I_1707 (I122864,I122843,I122849,I122858,I122855,I122840,I122852,I122861,I122840,I122846,I122867,I122913,I122916,I122919,I122922,I122925,I122928,I122931,I122934,I122937,I2224,I2231);
PAT_6 I_1708 (I122916,I122913,I122919,I122934,I122916,I122937,I122922,I122928,I122925,I122931,I122913,I122983,I122986,I122989,I122992,I122995,I122998,I123001,I123004,I123007,I123010,I2224,I2231);
PAT_5 I_1709 (I123004,I122983,I122989,I122992,I122998,I123001,I122983,I123007,I122986,I122995,I123010,I123056,I123059,I123062,I123065,I123068,I123071,I123074,I123077,I123080,I123083,I2224,I2231);
PAT_12 I_1710 (I123083,I123071,I123056,I123080,I123059,I123056,I123062,I123065,I123068,I123074,I123077,I123129,I123132,I123135,I123138,I123141,I123144,I123147,I123150,I2224,I2231);
PAT_4 I_1711 (I123135,I123132,I123147,I123150,I123144,I123138,I123129,I123129,I123135,I123141,I123132,I123196,I123199,I123202,I123205,I123208,I123211,I123214,I123217,I123220,I2224,I2231);
PAT_5 I_1712 (I123217,I123199,I123199,I123211,I123214,I123208,I123205,I123196,I123202,I123196,I123220,I123266,I123269,I123272,I123275,I123278,I123281,I123284,I123287,I123290,I123293,I2224,I2231);
PAT_9 I_1713 (I123281,I123278,I123287,I123284,I123275,I123266,I123272,I123293,I123269,I123290,I123266,I123339,I123342,I123345,I123348,I123351,I123354,I123357,I123360,I123363,I2224,I2231);
PAT_13 I_1714 (I123339,I123360,I123342,I123357,I123351,I123348,I123363,I123339,I123345,I123354,I123342,I123409,I123412,I123415,I123418,I123421,I123424,I123427,I123430,I123433,I2224,I2231);
PAT_9 I_1715 (I123430,I123412,I123412,I123409,I123433,I123415,I123418,I123409,I123421,I123427,I123424,I123479,I123482,I123485,I123488,I123491,I123494,I123497,I123500,I123503,I2224,I2231);
PAT_3 I_1716 (I123503,I123482,I123485,I123497,I123488,I123482,I123491,I123479,I123500,I123479,I123494,I123549,I123552,I123555,I123558,I123561,I123564,I123567,I123570,I123573,I123576,I2224,I2231);
PAT_17 I_1717 (I123561,I123576,I123555,I123564,I123552,I123567,I123549,I123558,I123570,I123549,I123573,I123622,I123625,I123628,I123631,I123634,I123637,I123640,I123643,I123646,I123649,I2224,I2231);
PAT_13 I_1718 (I123640,I123643,I123628,I123622,I123634,I123646,I123625,I123637,I123622,I123649,I123631,I123695,I123698,I123701,I123704,I123707,I123710,I123713,I123716,I123719,I2224,I2231);
PAT_3 I_1719 (I123719,I123698,I123713,I123701,I123707,I123716,I123695,I123704,I123695,I123698,I123710,I123765,I123768,I123771,I123774,I123777,I123780,I123783,I123786,I123789,I123792,I2224,I2231);
PAT_15 I_1720 (I123783,I123792,I123765,I123765,I123774,I123768,I123786,I123777,I123771,I123780,I123789,I123838,I123841,I123844,I123847,I123850,I123853,I123856,I123859,I123862,I2224,I2231);
PAT_2 I_1721 (I123841,I123841,I123844,I123850,I123838,I123838,I123847,I123862,I123856,I123859,I123853,I123908,I123911,I123914,I123917,I123920,I123923,I123926,I123929,I123932,I2224,I2231);
PAT_8 I_1722 (I123920,I123911,I123917,I123908,I123914,I123929,I123926,I123908,I123923,I123911,I123932,I123978,I123981,I123984,I123987,I123990,I123993,I123996,I123999,I124002,I2224,I2231);
PAT_14 I_1723 (I123984,I123996,I123981,I123978,I123981,I124002,I123978,I123990,I123993,I123999,I123987,I124048,I124051,I124054,I124057,I124060,I124063,I124066,I124069,I124072,I2224,I2231);
PAT_6 I_1724 (I124048,I124051,I124072,I124057,I124048,I124054,I124060,I124063,I124066,I124051,I124069,I124118,I124121,I124124,I124127,I124130,I124133,I124136,I124139,I124142,I124145,I2224,I2231);
PAT_9 I_1725 (I124118,I124145,I124142,I124124,I124130,I124121,I124133,I124118,I124136,I124127,I124139,I124191,I124194,I124197,I124200,I124203,I124206,I124209,I124212,I124215,I2224,I2231);
PAT_12 I_1726 (I124212,I124209,I124203,I124191,I124200,I124191,I124194,I124197,I124215,I124206,I124194,I124261,I124264,I124267,I124270,I124273,I124276,I124279,I124282,I2224,I2231);
PAT_5 I_1727 (I124270,I124276,I124282,I124267,I124267,I124261,I124279,I124261,I124264,I124264,I124273,I124328,I124331,I124334,I124337,I124340,I124343,I124346,I124349,I124352,I124355,I2224,I2231);
PAT_13 I_1728 (I124334,I124343,I124328,I124331,I124352,I124337,I124349,I124328,I124346,I124355,I124340,I124401,I124404,I124407,I124410,I124413,I124416,I124419,I124422,I124425,I2224,I2231);
PAT_10 I_1729 (I124422,I124416,I124410,I124404,I124425,I124404,I124413,I124401,I124401,I124419,I124407,I124471,I124474,I124477,I124480,I124483,I124486,I124489,I124492,I2224,I2231);
PAT_2 I_1730 (I124483,I124486,I124477,I124489,I124474,I124471,I124471,I124477,I124492,I124480,I124474,I124538,I124541,I124544,I124547,I124550,I124553,I124556,I124559,I124562,I2224,I2231);
PAT_9 I_1731 (I124553,I124562,I124538,I124544,I124547,I124556,I124541,I124550,I124559,I124541,I124538,I124608,I124611,I124614,I124617,I124620,I124623,I124626,I124629,I124632,I2224,I2231);
PAT_6 I_1732 (I124626,I124608,I124620,I124629,I124608,I124617,I124614,I124632,I124623,I124611,I124611,I124678,I124681,I124684,I124687,I124690,I124693,I124696,I124699,I124702,I124705,I2224,I2231);
PAT_9 I_1733 (I124678,I124705,I124702,I124684,I124690,I124681,I124693,I124678,I124696,I124687,I124699,I124751,I124754,I124757,I124760,I124763,I124766,I124769,I124772,I124775,I2224,I2231);
PAT_11 I_1734 (I124763,I124769,I124775,I124772,I124760,I124754,I124754,I124751,I124766,I124751,I124757,I124821,I124824,I124827,I124830,I124833,I124836,I124839,I124842,I124845,I124848,I2224,I2231);
PAT_5 I_1735 (I124842,I124821,I124848,I124836,I124833,I124845,I124827,I124821,I124839,I124824,I124830,I124894,I124897,I124900,I124903,I124906,I124909,I124912,I124915,I124918,I124921,I2224,I2231);
PAT_9 I_1736 (I124909,I124906,I124915,I124912,I124903,I124894,I124900,I124921,I124897,I124918,I124894,I124967,I124970,I124973,I124976,I124979,I124982,I124985,I124988,I124991,I2224,I2231);
PAT_10 I_1737 (I124988,I124985,I124973,I124970,I124991,I124976,I124982,I124970,I124967,I124967,I124979,I125037,I125040,I125043,I125046,I125049,I125052,I125055,I125058,I2224,I2231);
PAT_4 I_1738 (I125052,I125049,I125040,I125058,I125037,I125040,I125046,I125043,I125055,I125037,I125043,I125104,I125107,I125110,I125113,I125116,I125119,I125122,I125125,I125128,I2224,I2231);
PAT_15 I_1739 (I125104,I125107,I125128,I125113,I125122,I125125,I125110,I125119,I125116,I125104,I125107,I125174,I125177,I125180,I125183,I125186,I125189,I125192,I125195,I125198,I2224,I2231);
PAT_17 I_1740 (I125174,I125174,I125186,I125177,I125180,I125198,I125195,I125189,I125177,I125183,I125192,I125244,I125247,I125250,I125253,I125256,I125259,I125262,I125265,I125268,I125271,I2224,I2231);
PAT_5 I_1741 (I125256,I125250,I125247,I125268,I125253,I125259,I125262,I125244,I125244,I125265,I125271,I125317,I125320,I125323,I125326,I125329,I125332,I125335,I125338,I125341,I125344,I2224,I2231);
PAT_15 I_1742 (I125335,I125320,I125317,I125317,I125332,I125329,I125341,I125326,I125338,I125323,I125344,I125390,I125393,I125396,I125399,I125402,I125405,I125408,I125411,I125414,I2224,I2231);
PAT_6 I_1743 (I125393,I125390,I125396,I125411,I125393,I125414,I125399,I125405,I125402,I125408,I125390,I125460,I125463,I125466,I125469,I125472,I125475,I125478,I125481,I125484,I125487,I2224,I2231);
PAT_15 I_1744 (I125478,I125469,I125481,I125484,I125475,I125487,I125460,I125466,I125460,I125463,I125472,I125533,I125536,I125539,I125542,I125545,I125548,I125551,I125554,I125557,I2224,I2231);
PAT_4 I_1745 (I125545,I125551,I125533,I125536,I125539,I125533,I125557,I125554,I125542,I125548,I125536,I125603,I125606,I125609,I125612,I125615,I125618,I125621,I125624,I125627,I2224,I2231);
PAT_10 I_1746 (I125603,I125603,I125627,I125606,I125612,I125621,I125618,I125606,I125624,I125609,I125615,I125673,I125676,I125679,I125682,I125685,I125688,I125691,I125694,I2224,I2231);
PAT_6 I_1747 (I125694,I125688,I125682,I125676,I125673,I125679,I125673,I125679,I125676,I125685,I125691,I125740,I125743,I125746,I125749,I125752,I125755,I125758,I125761,I125764,I125767,I2224,I2231);
PAT_10 I_1748 (I125740,I125755,I125758,I125749,I125740,I125764,I125767,I125743,I125752,I125746,I125761,I125813,I125816,I125819,I125822,I125825,I125828,I125831,I125834,I2224,I2231);
PAT_9 I_1749 (I125825,I125813,I125816,I125819,I125813,I125819,I125822,I125816,I125834,I125828,I125831,I125880,I125883,I125886,I125889,I125892,I125895,I125898,I125901,I125904,I2224,I2231);
PAT_11 I_1750 (I125892,I125898,I125904,I125901,I125889,I125883,I125883,I125880,I125895,I125880,I125886,I125950,I125953,I125956,I125959,I125962,I125965,I125968,I125971,I125974,I125977,I2224,I2231);
PAT_12 I_1751 (I125959,I125974,I125956,I125953,I125962,I125965,I125971,I125950,I125968,I125977,I125950,I126023,I126026,I126029,I126032,I126035,I126038,I126041,I126044,I2224,I2231);
PAT_13 I_1752 (I126035,I126038,I126029,I126044,I126041,I126023,I126026,I126032,I126029,I126026,I126023,I126090,I126093,I126096,I126099,I126102,I126105,I126108,I126111,I126114,I2224,I2231);
PAT_2 I_1753 (I126108,I126102,I126099,I126105,I126090,I126114,I126093,I126111,I126090,I126096,I126093,I126160,I126163,I126166,I126169,I126172,I126175,I126178,I126181,I126184,I2224,I2231);
PAT_8 I_1754 (I126172,I126163,I126169,I126160,I126166,I126181,I126178,I126160,I126175,I126163,I126184,I126230,I126233,I126236,I126239,I126242,I126245,I126248,I126251,I126254,I2224,I2231);
PAT_5 I_1755 (I126236,I126254,I126230,I126251,I126239,I126242,I126233,I126230,I126233,I126245,I126248,I126300,I126303,I126306,I126309,I126312,I126315,I126318,I126321,I126324,I126327,I2224,I2231);
PAT_11 I_1756 (I126312,I126309,I126303,I126321,I126324,I126300,I126318,I126315,I126327,I126306,I126300,I126373,I126376,I126379,I126382,I126385,I126388,I126391,I126394,I126397,I126400,I2224,I2231);
PAT_4 I_1757 (I126379,I126400,I126373,I126391,I126382,I126373,I126394,I126376,I126385,I126397,I126388,I126446,I126449,I126452,I126455,I126458,I126461,I126464,I126467,I126470,I2224,I2231);
PAT_13 I_1758 (I126461,I126455,I126467,I126452,I126458,I126446,I126470,I126464,I126449,I126446,I126449,I126516,I126519,I126522,I126525,I126528,I126531,I126534,I126537,I126540,I2224,I2231);
PAT_11 I_1759 (I126516,I126528,I126531,I126522,I126519,I126540,I126519,I126537,I126525,I126516,I126534,I126586,I126589,I126592,I126595,I126598,I126601,I126604,I126607,I126610,I126613,I2224,I2231);
PAT_12 I_1760 (I126595,I126610,I126592,I126589,I126598,I126601,I126607,I126586,I126604,I126613,I126586,I126659,I126662,I126665,I126668,I126671,I126674,I126677,I126680,I2224,I2231);
PAT_3 I_1761 (I126659,I126659,I126665,I126671,I126665,I126677,I126680,I126662,I126662,I126668,I126674,I126726,I126729,I126732,I126735,I126738,I126741,I126744,I126747,I126750,I126753,I2224,I2231);
PAT_11 I_1762 (I126729,I126750,I126726,I126738,I126735,I126753,I126741,I126726,I126732,I126747,I126744,I126799,I126802,I126805,I126808,I126811,I126814,I126817,I126820,I126823,I126826,I2224,I2231);
PAT_6 I_1763 (I126799,I126826,I126814,I126823,I126817,I126811,I126802,I126820,I126808,I126805,I126799,I126872,I126875,I126878,I126881,I126884,I126887,I126890,I126893,I126896,I126899,I2224,I2231);
PAT_5 I_1764 (I126893,I126872,I126878,I126881,I126887,I126890,I126872,I126896,I126875,I126884,I126899,I126945,I126948,I126951,I126954,I126957,I126960,I126963,I126966,I126969,I126972,I2224,I2231);
PAT_4 I_1765 (I126963,I126969,I126972,I126951,I126954,I126966,I126948,I126945,I126957,I126960,I126945,I127018,I127021,I127024,I127027,I127030,I127033,I127036,I127039,I127042,I2224,I2231);
PAT_10 I_1766 (I127018,I127018,I127042,I127021,I127027,I127036,I127033,I127021,I127039,I127024,I127030,I127088,I127091,I127094,I127097,I127100,I127103,I127106,I127109,I2224,I2231);
PAT_11 I_1767 (I127097,I127100,I127109,I127103,I127106,I127088,I127088,I127094,I127091,I127091,I127094,I127155,I127158,I127161,I127164,I127167,I127170,I127173,I127176,I127179,I127182,I2224,I2231);
PAT_2 I_1768 (I127155,I127179,I127167,I127161,I127170,I127173,I127158,I127182,I127176,I127164,I127155,I127228,I127231,I127234,I127237,I127240,I127243,I127246,I127249,I127252,I2224,I2231);
PAT_4 I_1769 (I127228,I127234,I127252,I127246,I127243,I127240,I127231,I127249,I127228,I127231,I127237,I127298,I127301,I127304,I127307,I127310,I127313,I127316,I127319,I127322,I2224,I2231);
PAT_5 I_1770 (I127319,I127301,I127301,I127313,I127316,I127310,I127307,I127298,I127304,I127298,I127322,I127368,I127371,I127374,I127377,I127380,I127383,I127386,I127389,I127392,I127395,I2224,I2231);
PAT_9 I_1771 (I127383,I127380,I127389,I127386,I127377,I127368,I127374,I127395,I127371,I127392,I127368,I127441,I127444,I127447,I127450,I127453,I127456,I127459,I127462,I127465,I2224,I2231);
PAT_2 I_1772 (I127456,I127459,I127450,I127465,I127441,I127444,I127447,I127444,I127462,I127453,I127441,I127511,I127514,I127517,I127520,I127523,I127526,I127529,I127532,I127535,I2224,I2231);
PAT_10 I_1773 (I127511,I127529,I127526,I127514,I127517,I127532,I127523,I127511,I127520,I127535,I127514,I127581,I127584,I127587,I127590,I127593,I127596,I127599,I127602,I2224,I2231);
PAT_14 I_1774 (I127581,I127602,I127587,I127596,I127593,I127599,I127590,I127584,I127584,I127587,I127581,I127648,I127651,I127654,I127657,I127660,I127663,I127666,I127669,I127672,I2224,I2231);
PAT_10 I_1775 (I127651,I127648,I127654,I127672,I127669,I127663,I127651,I127666,I127648,I127660,I127657,I127718,I127721,I127724,I127727,I127730,I127733,I127736,I127739,I2224,I2231);
PAT_13 I_1776 (I127724,I127730,I127724,I127721,I127736,I127739,I127718,I127718,I127733,I127721,I127727,I127785,I127788,I127791,I127794,I127797,I127800,I127803,I127806,I127809,I2224,I2231);
PAT_8 I_1777 (I127794,I127806,I127797,I127800,I127809,I127788,I127803,I127785,I127788,I127791,I127785,I127855,I127858,I127861,I127864,I127867,I127870,I127873,I127876,I127879,I2224,I2231);
PAT_9 I_1778 (I127858,I127867,I127858,I127855,I127870,I127861,I127876,I127864,I127873,I127855,I127879,I127925,I127928,I127931,I127934,I127937,I127940,I127943,I127946,I127949,I2224,I2231);
PAT_17 I_1779 (I127928,I127934,I127949,I127940,I127943,I127931,I127925,I127937,I127925,I127928,I127946,I127995,I127998,I128001,I128004,I128007,I128010,I128013,I128016,I128019,I128022,I2224,I2231);
PAT_1 I_1780 (I128019,I128022,I128001,I128010,I127995,I128016,I128007,I127998,I128004,I127995,I128013,I128068,I128071,I128074,I128077,I128080,I128083,I128086,I128089,I128092,I2224,I2231);
PAT_13 I_1781 (I128077,I128086,I128092,I128068,I128083,I128080,I128089,I128074,I128071,I128068,I128071,I128138,I128141,I128144,I128147,I128150,I128153,I128156,I128159,I128162,I2224,I2231);
PAT_5 I_1782 (I128150,I128141,I128147,I128159,I128141,I128162,I128144,I128153,I128138,I128138,I128156,I128208,I128211,I128214,I128217,I128220,I128223,I128226,I128229,I128232,I128235,I2224,I2231);
PAT_9 I_1783 (I128223,I128220,I128229,I128226,I128217,I128208,I128214,I128235,I128211,I128232,I128208,I128281,I128284,I128287,I128290,I128293,I128296,I128299,I128302,I128305,I2224,I2231);
PAT_13 I_1784 (I128281,I128302,I128284,I128299,I128293,I128290,I128305,I128281,I128287,I128296,I128284,I128351,I128354,I128357,I128360,I128363,I128366,I128369,I128372,I128375,I2224,I2231);
PAT_12 I_1785 (I128360,I128351,I128351,I128375,I128372,I128354,I128369,I128363,I128354,I128357,I128366,I128421,I128424,I128427,I128430,I128433,I128436,I128439,I128442,I2224,I2231);
PAT_4 I_1786 (I128427,I128424,I128439,I128442,I128436,I128430,I128421,I128421,I128427,I128433,I128424,I128488,I128491,I128494,I128497,I128500,I128503,I128506,I128509,I128512,I2224,I2231);
PAT_5 I_1787 (I128509,I128491,I128491,I128503,I128506,I128500,I128497,I128488,I128494,I128488,I128512,I128558,I128561,I128564,I128567,I128570,I128573,I128576,I128579,I128582,I128585,I2224,I2231);
PAT_2 I_1788 (I128573,I128558,I128570,I128564,I128579,I128561,I128576,I128567,I128582,I128585,I128558,I128631,I128634,I128637,I128640,I128643,I128646,I128649,I128652,I128655,I2224,I2231);
PAT_15 I_1789 (I128634,I128646,I128652,I128655,I128637,I128649,I128631,I128640,I128631,I128643,I128634,I128701,I128704,I128707,I128710,I128713,I128716,I128719,I128722,I128725,I2224,I2231);
PAT_10 I_1790 (I128704,I128713,I128707,I128701,I128722,I128725,I128710,I128701,I128704,I128719,I128716,I128771,I128774,I128777,I128780,I128783,I128786,I128789,I128792,I2224,I2231);
PAT_17 I_1791 (I128783,I128792,I128786,I128771,I128777,I128789,I128774,I128774,I128771,I128777,I128780,I128838,I128841,I128844,I128847,I128850,I128853,I128856,I128859,I128862,I128865,I2224,I2231);
PAT_1 I_1792 (I128862,I128865,I128844,I128853,I128838,I128859,I128850,I128841,I128847,I128838,I128856,I128911,I128914,I128917,I128920,I128923,I128926,I128929,I128932,I128935,I2224,I2231);
PAT_11 I_1793 (I128914,I128929,I128926,I128932,I128935,I128914,I128920,I128923,I128911,I128917,I128911,I128981,I128984,I128987,I128990,I128993,I128996,I128999,I129002,I129005,I129008,I2224,I2231);
PAT_9 I_1794 (I128987,I128999,I128990,I129002,I128981,I128984,I128993,I128981,I128996,I129005,I129008,I129054,I129057,I129060,I129063,I129066,I129069,I129072,I129075,I129078,I2224,I2231);
PAT_11 I_1795 (I129066,I129072,I129078,I129075,I129063,I129057,I129057,I129054,I129069,I129054,I129060,I129124,I129127,I129130,I129133,I129136,I129139,I129142,I129145,I129148,I129151,I2224,I2231);
PAT_17 I_1796 (I129136,I129127,I129151,I129124,I129133,I129145,I129142,I129139,I129124,I129148,I129130,I129197,I129200,I129203,I129206,I129209,I129212,I129215,I129218,I129221,I129224,I2224,I2231);
PAT_9 I_1797 (I129218,I129200,I129206,I129221,I129203,I129215,I129197,I129209,I129197,I129224,I129212,I129270,I129273,I129276,I129279,I129282,I129285,I129288,I129291,I129294,I2224,I2231);
PAT_6 I_1798 (I129288,I129270,I129282,I129291,I129270,I129279,I129276,I129294,I129285,I129273,I129273,I129340,I129343,I129346,I129349,I129352,I129355,I129358,I129361,I129364,I129367,I2224,I2231);
PAT_5 I_1799 (I129361,I129340,I129346,I129349,I129355,I129358,I129340,I129364,I129343,I129352,I129367,I129413,I129416,I129419,I129422,I129425,I129428,I129431,I129434,I129437,I129440,I2224,I2231);
PAT_4 I_1800 (I129431,I129437,I129440,I129419,I129422,I129434,I129416,I129413,I129425,I129428,I129413,I129486,I129489,I129492,I129495,I129498,I129501,I129504,I129507,I129510,I2224,I2231);
PAT_17 I_1801 (I129498,I129495,I129507,I129501,I129486,I129504,I129510,I129489,I129492,I129489,I129486,I129556,I129559,I129562,I129565,I129568,I129571,I129574,I129577,I129580,I129583,I2224,I2231);
PAT_11 I_1802 (I129568,I129577,I129583,I129559,I129556,I129574,I129565,I129571,I129562,I129580,I129556,I129629,I129632,I129635,I129638,I129641,I129644,I129647,I129650,I129653,I129656,I2224,I2231);
PAT_13 I_1803 (I129629,I129632,I129641,I129653,I129656,I129644,I129650,I129638,I129647,I129635,I129629,I129702,I129705,I129708,I129711,I129714,I129717,I129720,I129723,I129726,I2224,I2231);
PAT_1 I_1804 (I129702,I129711,I129705,I129723,I129717,I129708,I129720,I129714,I129705,I129726,I129702,I129772,I129775,I129778,I129781,I129784,I129787,I129790,I129793,I129796,I2224,I2231);
PAT_12 I_1805 (I129784,I129778,I129796,I129772,I129781,I129772,I129775,I129793,I129787,I129775,I129790,I129842,I129845,I129848,I129851,I129854,I129857,I129860,I129863,I2224,I2231);
PAT_4 I_1806 (I129848,I129845,I129860,I129863,I129857,I129851,I129842,I129842,I129848,I129854,I129845,I129909,I129912,I129915,I129918,I129921,I129924,I129927,I129930,I129933,I2224,I2231);
PAT_15 I_1807 (I129909,I129912,I129933,I129918,I129927,I129930,I129915,I129924,I129921,I129909,I129912,I129979,I129982,I129985,I129988,I129991,I129994,I129997,I130000,I130003,I2224,I2231);
PAT_9 I_1808 (I129979,I130000,I129988,I129982,I129994,I129982,I129997,I130003,I129985,I129979,I129991,I130049,I130052,I130055,I130058,I130061,I130064,I130067,I130070,I130073,I2224,I2231);
PAT_5 I_1809 (I130070,I130049,I130064,I130049,I130055,I130058,I130052,I130052,I130067,I130061,I130073,I130119,I130122,I130125,I130128,I130131,I130134,I130137,I130140,I130143,I130146,I2224,I2231);
PAT_4 I_1810 (I130137,I130143,I130146,I130125,I130128,I130140,I130122,I130119,I130131,I130134,I130119,I130192,I130195,I130198,I130201,I130204,I130207,I130210,I130213,I130216,I2224,I2231);
PAT_13 I_1811 (I130207,I130201,I130213,I130198,I130204,I130192,I130216,I130210,I130195,I130192,I130195,I130262,I130265,I130268,I130271,I130274,I130277,I130280,I130283,I130286,I2224,I2231);
PAT_16 I_1812 (I130268,I130271,I130280,I130274,I130286,I130262,I130283,I130277,I130265,I130265,I130262,I130332,I130335,I130338,I130341,I130344,I130347,I130350,I130353,I130356,I130359,I2224,I2231);
PAT_15 I_1813 (I130356,I130332,I130353,I130347,I130338,I130341,I130332,I130335,I130359,I130350,I130344,I130405,I130408,I130411,I130414,I130417,I130420,I130423,I130426,I130429,I2224,I2231);
PAT_1 I_1814 (I130411,I130408,I130408,I130405,I130405,I130414,I130429,I130423,I130417,I130420,I130426,I130475,I130478,I130481,I130484,I130487,I130490,I130493,I130496,I130499,I2224,I2231);
PAT_12 I_1815 (I130487,I130481,I130499,I130475,I130484,I130475,I130478,I130496,I130490,I130478,I130493,I130545,I130548,I130551,I130554,I130557,I130560,I130563,I130566,I2224,I2231);
PAT_17 I_1816 (I130560,I130554,I130548,I130545,I130545,I130551,I130551,I130563,I130566,I130548,I130557,I130612,I130615,I130618,I130621,I130624,I130627,I130630,I130633,I130636,I130639,I2224,I2231);
PAT_9 I_1817 (I130633,I130615,I130621,I130636,I130618,I130630,I130612,I130624,I130612,I130639,I130627,I130685,I130688,I130691,I130694,I130697,I130700,I130703,I130706,I130709,I2224,I2231);
PAT_4 I_1818 (I130685,I130709,I130703,I130691,I130688,I130706,I130688,I130685,I130700,I130694,I130697,I130755,I130758,I130761,I130764,I130767,I130770,I130773,I130776,I130779,I2224,I2231);
PAT_9 I_1819 (I130776,I130758,I130761,I130770,I130773,I130755,I130764,I130758,I130779,I130755,I130767,I130825,I130828,I130831,I130834,I130837,I130840,I130843,I130846,I130849,I2224,I2231);
PAT_10 I_1820 (I130846,I130843,I130831,I130828,I130849,I130834,I130840,I130828,I130825,I130825,I130837,I130895,I130898,I130901,I130904,I130907,I130910,I130913,I130916,I2224,I2231);
PAT_11 I_1821 (I130904,I130907,I130916,I130910,I130913,I130895,I130895,I130901,I130898,I130898,I130901,I130962,I130965,I130968,I130971,I130974,I130977,I130980,I130983,I130986,I130989,I2224,I2231);
PAT_6 I_1822 (I130962,I130989,I130977,I130986,I130980,I130974,I130965,I130983,I130971,I130968,I130962,I131035,I131038,I131041,I131044,I131047,I131050,I131053,I131056,I131059,I131062,I2224,I2231);
PAT_13 I_1823 (I131059,I131041,I131056,I131035,I131038,I131044,I131062,I131047,I131053,I131035,I131050,I131108,I131111,I131114,I131117,I131120,I131123,I131126,I131129,I131132,I2224,I2231);
PAT_17 I_1824 (I131132,I131120,I131129,I131126,I131117,I131108,I131111,I131114,I131108,I131123,I131111,I131178,I131181,I131184,I131187,I131190,I131193,I131196,I131199,I131202,I131205,I2224,I2231);
PAT_9 I_1825 (I131199,I131181,I131187,I131202,I131184,I131196,I131178,I131190,I131178,I131205,I131193,I131251,I131254,I131257,I131260,I131263,I131266,I131269,I131272,I131275,I2224,I2231);
PAT_6 I_1826 (I131269,I131251,I131263,I131272,I131251,I131260,I131257,I131275,I131266,I131254,I131254,I131321,I131324,I131327,I131330,I131333,I131336,I131339,I131342,I131345,I131348,I2224,I2231);
PAT_9 I_1827 (I131321,I131348,I131345,I131327,I131333,I131324,I131336,I131321,I131339,I131330,I131342,I131394,I131397,I131400,I131403,I131406,I131409,I131412,I131415,I131418,I2224,I2231);
PAT_4 I_1828 (I131394,I131418,I131412,I131400,I131397,I131415,I131397,I131394,I131409,I131403,I131406,I131464,I131467,I131470,I131473,I131476,I131479,I131482,I131485,I131488,I2224,I2231);
PAT_13 I_1829 (I131479,I131473,I131485,I131470,I131476,I131464,I131488,I131482,I131467,I131464,I131467,I131534,I131537,I131540,I131543,I131546,I131549,I131552,I131555,I131558,I2224,I2231);
PAT_2 I_1830 (I131552,I131546,I131543,I131549,I131534,I131558,I131537,I131555,I131534,I131540,I131537,I131604,I131607,I131610,I131613,I131616,I131619,I131622,I131625,I131628,I2224,I2231);
PAT_12 I_1831 (I131613,I131610,I131604,I131607,I131628,I131622,I131625,I131607,I131619,I131604,I131616,I131674,I131677,I131680,I131683,I131686,I131689,I131692,I131695,I2224,I2231);
PAT_4 I_1832 (I131680,I131677,I131692,I131695,I131689,I131683,I131674,I131674,I131680,I131686,I131677,I131741,I131744,I131747,I131750,I131753,I131756,I131759,I131762,I131765,I2224,I2231);
PAT_10 I_1833 (I131741,I131741,I131765,I131744,I131750,I131759,I131756,I131744,I131762,I131747,I131753,I131811,I131814,I131817,I131820,I131823,I131826,I131829,I131832,I2224,I2231);
PAT_4 I_1834 (I131826,I131823,I131814,I131832,I131811,I131814,I131820,I131817,I131829,I131811,I131817,I131878,I131881,I131884,I131887,I131890,I131893,I131896,I131899,I131902,I2224,I2231);
PAT_2 I_1835 (I131887,I131881,I131881,I131902,I131878,I131896,I131893,I131884,I131878,I131890,I131899,I131948,I131951,I131954,I131957,I131960,I131963,I131966,I131969,I131972,I2224,I2231);
PAT_17 I_1836 (I131948,I131948,I131960,I131951,I131954,I131966,I131963,I131972,I131951,I131957,I131969,I132018,I132021,I132024,I132027,I132030,I132033,I132036,I132039,I132042,I132045,I2224,I2231);
PAT_2 I_1837 (I132018,I132036,I132033,I132018,I132027,I132042,I132039,I132024,I132045,I132030,I132021,I132091,I132094,I132097,I132100,I132103,I132106,I132109,I132112,I132115,I2224,I2231);
PAT_8 I_1838 (I132103,I132094,I132100,I132091,I132097,I132112,I132109,I132091,I132106,I132094,I132115,I132161,I132164,I132167,I132170,I132173,I132176,I132179,I132182,I132185,I2224,I2231);
PAT_13 I_1839 (I132173,I132182,I132164,I132185,I132167,I132161,I132161,I132170,I132179,I132176,I132164,I132231,I132234,I132237,I132240,I132243,I132246,I132249,I132252,I132255,I2224,I2231);
PAT_4 I_1840 (I132240,I132243,I132255,I132237,I132252,I132249,I132234,I132246,I132234,I132231,I132231,I132301,I132304,I132307,I132310,I132313,I132316,I132319,I132322,I132325,I2224,I2231);
PAT_15 I_1841 (I132301,I132304,I132325,I132310,I132319,I132322,I132307,I132316,I132313,I132301,I132304,I132371,I132374,I132377,I132380,I132383,I132386,I132389,I132392,I132395,I2224,I2231);
PAT_2 I_1842 (I132374,I132374,I132377,I132383,I132371,I132371,I132380,I132395,I132389,I132392,I132386,I132441,I132444,I132447,I132450,I132453,I132456,I132459,I132462,I132465,I2224,I2231);
PAT_9 I_1843 (I132456,I132465,I132441,I132447,I132450,I132459,I132444,I132453,I132462,I132444,I132441,I132511,I132514,I132517,I132520,I132523,I132526,I132529,I132532,I132535,I2224,I2231);
PAT_12 I_1844 (I132532,I132529,I132523,I132511,I132520,I132511,I132514,I132517,I132535,I132526,I132514,I132581,I132584,I132587,I132590,I132593,I132596,I132599,I132602,I2224,I2231);
PAT_2 I_1845 (I132599,I132593,I132602,I132596,I132590,I132587,I132581,I132581,I132587,I132584,I132584,I132648,I132651,I132654,I132657,I132660,I132663,I132666,I132669,I132672,I2224,I2231);
PAT_6 I_1846 (I132672,I132648,I132663,I132660,I132666,I132657,I132651,I132669,I132648,I132654,I132651,I132718,I132721,I132724,I132727,I132730,I132733,I132736,I132739,I132742,I132745,I2224,I2231);
PAT_9 I_1847 (I132718,I132745,I132742,I132724,I132730,I132721,I132733,I132718,I132736,I132727,I132739,I132791,I132794,I132797,I132800,I132803,I132806,I132809,I132812,I132815,I2224,I2231);
PAT_2 I_1848 (I132806,I132809,I132800,I132815,I132791,I132794,I132797,I132794,I132812,I132803,I132791,I132861,I132864,I132867,I132870,I132873,I132876,I132879,I132882,I132885,I2224,I2231);
PAT_17 I_1849 (I132861,I132861,I132873,I132864,I132867,I132879,I132876,I132885,I132864,I132870,I132882,I132931,I132934,I132937,I132940,I132943,I132946,I132949,I132952,I132955,I132958,I2224,I2231);
PAT_4 I_1850 (I132940,I132931,I132949,I132946,I132958,I132955,I132934,I132931,I132937,I132943,I132952,I133004,I133007,I133010,I133013,I133016,I133019,I133022,I133025,I133028,I2224,I2231);
PAT_5 I_1851 (I133025,I133007,I133007,I133019,I133022,I133016,I133013,I133004,I133010,I133004,I133028,I133074,I133077,I133080,I133083,I133086,I133089,I133092,I133095,I133098,I133101,I2224,I2231);
PAT_16 I_1852 (I133092,I133086,I133098,I133101,I133080,I133074,I133077,I133089,I133083,I133095,I133074,I133147,I133150,I133153,I133156,I133159,I133162,I133165,I133168,I133171,I133174,I2224,I2231);
PAT_4 I_1853 (I133159,I133165,I133150,I133162,I133147,I133153,I133156,I133168,I133171,I133147,I133174,I133220,I133223,I133226,I133229,I133232,I133235,I133238,I133241,I133244,I2224,I2231);
PAT_6 I_1854 (I133220,I133226,I133223,I133235,I133238,I133232,I133244,I133241,I133220,I133229,I133223,I133290,I133293,I133296,I133299,I133302,I133305,I133308,I133311,I133314,I133317,I2224,I2231);
PAT_8 I_1855 (I133299,I133305,I133296,I133308,I133290,I133293,I133311,I133290,I133317,I133314,I133302,I133363,I133366,I133369,I133372,I133375,I133378,I133381,I133384,I133387,I2224,I2231);
PAT_10 I_1856 (I133369,I133363,I133366,I133387,I133381,I133366,I133375,I133363,I133384,I133378,I133372,I133433,I133436,I133439,I133442,I133445,I133448,I133451,I133454,I2224,I2231);
PAT_11 I_1857 (I133442,I133445,I133454,I133448,I133451,I133433,I133433,I133439,I133436,I133436,I133439,I133500,I133503,I133506,I133509,I133512,I133515,I133518,I133521,I133524,I133527,I2224,I2231);
PAT_9 I_1858 (I133506,I133518,I133509,I133521,I133500,I133503,I133512,I133500,I133515,I133524,I133527,I133573,I133576,I133579,I133582,I133585,I133588,I133591,I133594,I133597,I2224,I2231);
PAT_13 I_1859 (I133573,I133594,I133576,I133591,I133585,I133582,I133597,I133573,I133579,I133588,I133576,I133643,I133646,I133649,I133652,I133655,I133658,I133661,I133664,I133667,I2224,I2231);
PAT_5 I_1860 (I133655,I133646,I133652,I133664,I133646,I133667,I133649,I133658,I133643,I133643,I133661,I133713,I133716,I133719,I133722,I133725,I133728,I133731,I133734,I133737,I133740,I2224,I2231);
PAT_11 I_1861 (I133725,I133722,I133716,I133734,I133737,I133713,I133731,I133728,I133740,I133719,I133713,I133786,I133789,I133792,I133795,I133798,I133801,I133804,I133807,I133810,I133813,I2224,I2231);
PAT_13 I_1862 (I133786,I133789,I133798,I133810,I133813,I133801,I133807,I133795,I133804,I133792,I133786,I133859,I133862,I133865,I133868,I133871,I133874,I133877,I133880,I133883,I2224,I2231);
PAT_3 I_1863 (I133883,I133862,I133877,I133865,I133871,I133880,I133859,I133868,I133859,I133862,I133874,I133929,I133932,I133935,I133938,I133941,I133944,I133947,I133950,I133953,I133956,I2224,I2231);
PAT_13 I_1864 (I133950,I133938,I133956,I133935,I133941,I133944,I133932,I133947,I133929,I133929,I133953,I134002,I134005,I134008,I134011,I134014,I134017,I134020,I134023,I134026,I2224,I2231);
PAT_9 I_1865 (I134023,I134005,I134005,I134002,I134026,I134008,I134011,I134002,I134014,I134020,I134017,I134072,I134075,I134078,I134081,I134084,I134087,I134090,I134093,I134096,I2224,I2231);
PAT_10 I_1866 (I134093,I134090,I134078,I134075,I134096,I134081,I134087,I134075,I134072,I134072,I134084,I134142,I134145,I134148,I134151,I134154,I134157,I134160,I134163,I2224,I2231);
PAT_17 I_1867 (I134154,I134163,I134157,I134142,I134148,I134160,I134145,I134145,I134142,I134148,I134151,I134209,I134212,I134215,I134218,I134221,I134224,I134227,I134230,I134233,I134236,I2224,I2231);
PAT_8 I_1868 (I134218,I134230,I134236,I134227,I134212,I134221,I134224,I134233,I134215,I134209,I134209,I134282,I134285,I134288,I134291,I134294,I134297,I134300,I134303,I134306,I2224,I2231);
PAT_10 I_1869 (I134288,I134282,I134285,I134306,I134300,I134285,I134294,I134282,I134303,I134297,I134291,I134352,I134355,I134358,I134361,I134364,I134367,I134370,I134373,I2224,I2231);
PAT_6 I_1870 (I134373,I134367,I134361,I134355,I134352,I134358,I134352,I134358,I134355,I134364,I134370,I134419,I134422,I134425,I134428,I134431,I134434,I134437,I134440,I134443,I134446,I2224,I2231);
PAT_16 I_1871 (I134437,I134446,I134443,I134434,I134428,I134431,I134425,I134419,I134419,I134440,I134422,I134492,I134495,I134498,I134501,I134504,I134507,I134510,I134513,I134516,I134519,I2224,I2231);
PAT_9 I_1872 (I134510,I134492,I134492,I134501,I134498,I134516,I134519,I134495,I134513,I134507,I134504,I134565,I134568,I134571,I134574,I134577,I134580,I134583,I134586,I134589,I2224,I2231);
PAT_10 I_1873 (I134586,I134583,I134571,I134568,I134589,I134574,I134580,I134568,I134565,I134565,I134577,I134635,I134638,I134641,I134644,I134647,I134650,I134653,I134656,I2224,I2231);
PAT_8 I_1874 (I134656,I134647,I134638,I134635,I134644,I134635,I134650,I134638,I134653,I134641,I134641,I134702,I134705,I134708,I134711,I134714,I134717,I134720,I134723,I134726,I2224,I2231);
PAT_9 I_1875 (I134705,I134714,I134705,I134702,I134717,I134708,I134723,I134711,I134720,I134702,I134726,I134772,I134775,I134778,I134781,I134784,I134787,I134790,I134793,I134796,I2224,I2231);
PAT_8 I_1876 (I134793,I134781,I134790,I134772,I134775,I134787,I134796,I134775,I134778,I134784,I134772,I134842,I134845,I134848,I134851,I134854,I134857,I134860,I134863,I134866,I2224,I2231);
PAT_2 I_1877 (I134845,I134860,I134866,I134842,I134854,I134857,I134845,I134863,I134848,I134851,I134842,I134912,I134915,I134918,I134921,I134924,I134927,I134930,I134933,I134936,I2224,I2231);
PAT_11 I_1878 (I134915,I134927,I134912,I134924,I134921,I134933,I134930,I134915,I134936,I134918,I134912,I134982,I134985,I134988,I134991,I134994,I134997,I135000,I135003,I135006,I135009,I2224,I2231);
PAT_9 I_1879 (I134988,I135000,I134991,I135003,I134982,I134985,I134994,I134982,I134997,I135006,I135009,I135055,I135058,I135061,I135064,I135067,I135070,I135073,I135076,I135079,I2224,I2231);
PAT_6 I_1880 (I135073,I135055,I135067,I135076,I135055,I135064,I135061,I135079,I135070,I135058,I135058,I135125,I135128,I135131,I135134,I135137,I135140,I135143,I135146,I135149,I135152,I2224,I2231);
PAT_8 I_1881 (I135134,I135140,I135131,I135143,I135125,I135128,I135146,I135125,I135152,I135149,I135137,I135198,I135201,I135204,I135207,I135210,I135213,I135216,I135219,I135222,I2224,I2231);
PAT_5 I_1882 (I135204,I135222,I135198,I135219,I135207,I135210,I135201,I135198,I135201,I135213,I135216,I135268,I135271,I135274,I135277,I135280,I135283,I135286,I135289,I135292,I135295,I2224,I2231);
PAT_4 I_1883 (I135286,I135292,I135295,I135274,I135277,I135289,I135271,I135268,I135280,I135283,I135268,I135341,I135344,I135347,I135350,I135353,I135356,I135359,I135362,I135365,I2224,I2231);
PAT_13 I_1884 (I135356,I135350,I135362,I135347,I135353,I135341,I135365,I135359,I135344,I135341,I135344,I135411,I135414,I135417,I135420,I135423,I135426,I135429,I135432,I135435,I2224,I2231);
PAT_11 I_1885 (I135411,I135423,I135426,I135417,I135414,I135435,I135414,I135432,I135420,I135411,I135429,I135481,I135484,I135487,I135490,I135493,I135496,I135499,I135502,I135505,I135508,I2224,I2231);
PAT_10 I_1886 (I135496,I135502,I135493,I135487,I135505,I135490,I135508,I135499,I135481,I135484,I135481,I135554,I135557,I135560,I135563,I135566,I135569,I135572,I135575,I2224,I2231);
PAT_6 I_1887 (I135575,I135569,I135563,I135557,I135554,I135560,I135554,I135560,I135557,I135566,I135572,I135621,I135624,I135627,I135630,I135633,I135636,I135639,I135642,I135645,I135648,I2224,I2231);
PAT_17 I_1888 (I135633,I135636,I135642,I135630,I135624,I135645,I135639,I135621,I135648,I135627,I135621,I135694,I135697,I135700,I135703,I135706,I135709,I135712,I135715,I135718,I135721,I2224,I2231);
PAT_10 I_1889 (I135694,I135700,I135721,I135703,I135718,I135697,I135712,I135706,I135715,I135709,I135694,I135767,I135770,I135773,I135776,I135779,I135782,I135785,I135788,I2224,I2231);
PAT_4 I_1890 (I135782,I135779,I135770,I135788,I135767,I135770,I135776,I135773,I135785,I135767,I135773,I135834,I135837,I135840,I135843,I135846,I135849,I135852,I135855,I135858,I2224,I2231);
PAT_10 I_1891 (I135834,I135834,I135858,I135837,I135843,I135852,I135849,I135837,I135855,I135840,I135846,I135904,I135907,I135910,I135913,I135916,I135919,I135922,I135925,I2224,I2231);
PAT_12 I_1892 (I135910,I135904,I135904,I135916,I135919,I135907,I135907,I135922,I135925,I135910,I135913,I135971,I135974,I135977,I135980,I135983,I135986,I135989,I135992,I2224,I2231);
PAT_13 I_1893 (I135983,I135986,I135977,I135992,I135989,I135971,I135974,I135980,I135977,I135974,I135971,I136038,I136041,I136044,I136047,I136050,I136053,I136056,I136059,I136062,I2224,I2231);
PAT_2 I_1894 (I136056,I136050,I136047,I136053,I136038,I136062,I136041,I136059,I136038,I136044,I136041,I136108,I136111,I136114,I136117,I136120,I136123,I136126,I136129,I136132,I2224,I2231);
PAT_5 I_1895 (I136129,I136108,I136108,I136120,I136117,I136126,I136114,I136123,I136132,I136111,I136111,I136178,I136181,I136184,I136187,I136190,I136193,I136196,I136199,I136202,I136205,I2224,I2231);
PAT_13 I_1896 (I136184,I136193,I136178,I136181,I136202,I136187,I136199,I136178,I136196,I136205,I136190,I136251,I136254,I136257,I136260,I136263,I136266,I136269,I136272,I136275,I2224,I2231);
PAT_0 I_1897 (I136257,I136260,I136251,I136251,I136263,I136272,I136275,I136266,I136269,I136254,I136254,I136321,I136324,I136327,I136330,I136333,I136336,I136339,I136342,I2224,I2231);
PAT_9 I_1898 (I136327,I136339,I136324,I136333,I136336,I136324,I136321,I136330,I136342,I136327,I136321,I136388,I136391,I136394,I136397,I136400,I136403,I136406,I136409,I136412,I2224,I2231);
PAT_12 I_1899 (I136409,I136406,I136400,I136388,I136397,I136388,I136391,I136394,I136412,I136403,I136391,I136458,I136461,I136464,I136467,I136470,I136473,I136476,I136479,I2224,I2231);
PAT_10 I_1900 (I136458,I136479,I136470,I136473,I136464,I136461,I136458,I136476,I136464,I136467,I136461,I136525,I136528,I136531,I136534,I136537,I136540,I136543,I136546,I2224,I2231);
PAT_5 I_1901 (I136546,I136525,I136534,I136528,I136543,I136540,I136531,I136531,I136525,I136528,I136537,I136592,I136595,I136598,I136601,I136604,I136607,I136610,I136613,I136616,I136619,I2224,I2231);
PAT_11 I_1902 (I136604,I136601,I136595,I136613,I136616,I136592,I136610,I136607,I136619,I136598,I136592,I136665,I136668,I136671,I136674,I136677,I136680,I136683,I136686,I136689,I136692,I2224,I2231);
PAT_2 I_1903 (I136665,I136689,I136677,I136671,I136680,I136683,I136668,I136692,I136686,I136674,I136665,I136738,I136741,I136744,I136747,I136750,I136753,I136756,I136759,I136762,I2224,I2231);
PAT_9 I_1904 (I136753,I136762,I136738,I136744,I136747,I136756,I136741,I136750,I136759,I136741,I136738,I136808,I136811,I136814,I136817,I136820,I136823,I136826,I136829,I136832,I2224,I2231);
PAT_4 I_1905 (I136808,I136832,I136826,I136814,I136811,I136829,I136811,I136808,I136823,I136817,I136820,I136878,I136881,I136884,I136887,I136890,I136893,I136896,I136899,I136902,I2224,I2231);
PAT_10 I_1906 (I136878,I136878,I136902,I136881,I136887,I136896,I136893,I136881,I136899,I136884,I136890,I136948,I136951,I136954,I136957,I136960,I136963,I136966,I136969,I2224,I2231);
PAT_0 I_1907 (I136951,I136954,I136963,I136951,I136969,I136966,I136960,I136948,I136954,I136957,I136948,I137015,I137018,I137021,I137024,I137027,I137030,I137033,I137036,I2224,I2231);
PAT_11 I_1908 (I137021,I137030,I137036,I137015,I137033,I137021,I137018,I137024,I137027,I137015,I137018,I137082,I137085,I137088,I137091,I137094,I137097,I137100,I137103,I137106,I137109,I2224,I2231);
PAT_2 I_1909 (I137082,I137106,I137094,I137088,I137097,I137100,I137085,I137109,I137103,I137091,I137082,I137155,I137158,I137161,I137164,I137167,I137170,I137173,I137176,I137179,I2224,I2231);
PAT_4 I_1910 (I137155,I137161,I137179,I137173,I137170,I137167,I137158,I137176,I137155,I137158,I137164,I137225,I137228,I137231,I137234,I137237,I137240,I137243,I137246,I137249,I2224,I2231);
PAT_10 I_1911 (I137225,I137225,I137249,I137228,I137234,I137243,I137240,I137228,I137246,I137231,I137237,I137295,I137298,I137301,I137304,I137307,I137310,I137313,I137316,I2224,I2231);
PAT_9 I_1912 (I137307,I137295,I137298,I137301,I137295,I137301,I137304,I137298,I137316,I137310,I137313,I137362,I137365,I137368,I137371,I137374,I137377,I137380,I137383,I137386,I2224,I2231);
PAT_12 I_1913 (I137383,I137380,I137374,I137362,I137371,I137362,I137365,I137368,I137386,I137377,I137365,I137432,I137435,I137438,I137441,I137444,I137447,I137450,I137453,I2224,I2231);
PAT_5 I_1914 (I137441,I137447,I137453,I137438,I137438,I137432,I137450,I137432,I137435,I137435,I137444,I137499,I137502,I137505,I137508,I137511,I137514,I137517,I137520,I137523,I137526,I2224,I2231);
PAT_9 I_1915 (I137514,I137511,I137520,I137517,I137508,I137499,I137505,I137526,I137502,I137523,I137499,I137572,I137575,I137578,I137581,I137584,I137587,I137590,I137593,I137596,I2224,I2231);
PAT_11 I_1916 (I137584,I137590,I137596,I137593,I137581,I137575,I137575,I137572,I137587,I137572,I137578,I137642,I137645,I137648,I137651,I137654,I137657,I137660,I137663,I137666,I137669,I2224,I2231);
PAT_1 I_1917 (I137657,I137648,I137651,I137642,I137663,I137660,I137645,I137642,I137669,I137666,I137654,I137715,I137718,I137721,I137724,I137727,I137730,I137733,I137736,I137739,I2224,I2231);
PAT_9 I_1918 (I137730,I137736,I137721,I137739,I137718,I137733,I137718,I137724,I137715,I137727,I137715,I137785,I137788,I137791,I137794,I137797,I137800,I137803,I137806,I137809,I2224,I2231);
PAT_0 I_1919 (I137794,I137806,I137785,I137788,I137791,I137785,I137800,I137803,I137797,I137809,I137788,I137855,I137858,I137861,I137864,I137867,I137870,I137873,I137876,I2224,I2231);
PAT_17 I_1920 (I137876,I137873,I137861,I137855,I137858,I137867,I137864,I137870,I137861,I137855,I137858,I137922,I137925,I137928,I137931,I137934,I137937,I137940,I137943,I137946,I137949,I2224,I2231);
PAT_9 I_1921 (I137943,I137925,I137931,I137946,I137928,I137940,I137922,I137934,I137922,I137949,I137937,I137995,I137998,I138001,I138004,I138007,I138010,I138013,I138016,I138019,I2224,I2231);
PAT_7 I_1922 (I138001,I138010,I137995,I138016,I138007,I137995,I137998,I138019,I138013,I137998,I138004,I138065,I138068,I138071,I138074,I138077,I138080,I138083,I138086,I138089,I2224,I2231);
PAT_9 I_1923 (I138086,I138074,I138083,I138089,I138071,I138077,I138068,I138080,I138065,I138065,I138068,I138135,I138138,I138141,I138144,I138147,I138150,I138153,I138156,I138159,I2224,I2231);
PAT_14 I_1924 (I138144,I138135,I138159,I138141,I138138,I138135,I138150,I138156,I138147,I138138,I138153,I138205,I138208,I138211,I138214,I138217,I138220,I138223,I138226,I138229,I2224,I2231);
PAT_15 I_1925 (I138217,I138211,I138208,I138226,I138223,I138214,I138205,I138208,I138205,I138220,I138229,I138275,I138278,I138281,I138284,I138287,I138290,I138293,I138296,I138299,I2224,I2231);
PAT_10 I_1926 (I138278,I138287,I138281,I138275,I138296,I138299,I138284,I138275,I138278,I138293,I138290,I138345,I138348,I138351,I138354,I138357,I138360,I138363,I138366,I2224,I2231);
PAT_17 I_1927 (I138357,I138366,I138360,I138345,I138351,I138363,I138348,I138348,I138345,I138351,I138354,I138412,I138415,I138418,I138421,I138424,I138427,I138430,I138433,I138436,I138439,I2224,I2231);
PAT_12 I_1928 (I138436,I138418,I138412,I138430,I138424,I138433,I138415,I138439,I138412,I138421,I138427,I138485,I138488,I138491,I138494,I138497,I138500,I138503,I138506,I2224,I2231);
PAT_6 I_1929 (I138494,I138488,I138506,I138491,I138488,I138491,I138500,I138485,I138503,I138485,I138497,I138552,I138555,I138558,I138561,I138564,I138567,I138570,I138573,I138576,I138579,I2224,I2231);
PAT_8 I_1930 (I138561,I138567,I138558,I138570,I138552,I138555,I138573,I138552,I138579,I138576,I138564,I138625,I138628,I138631,I138634,I138637,I138640,I138643,I138646,I138649,I2224,I2231);
PAT_3 I_1931 (I138646,I138637,I138628,I138634,I138631,I138643,I138628,I138649,I138625,I138640,I138625,I138695,I138698,I138701,I138704,I138707,I138710,I138713,I138716,I138719,I138722,I2224,I2231);
PAT_13 I_1932 (I138716,I138704,I138722,I138701,I138707,I138710,I138698,I138713,I138695,I138695,I138719,I138768,I138771,I138774,I138777,I138780,I138783,I138786,I138789,I138792,I2224,I2231);
PAT_9 I_1933 (I138789,I138771,I138771,I138768,I138792,I138774,I138777,I138768,I138780,I138786,I138783,I138838,I138841,I138844,I138847,I138850,I138853,I138856,I138859,I138862,I2224,I2231);
PAT_17 I_1934 (I138841,I138847,I138862,I138853,I138856,I138844,I138838,I138850,I138838,I138841,I138859,I138908,I138911,I138914,I138917,I138920,I138923,I138926,I138929,I138932,I138935,I2224,I2231);
PAT_10 I_1935 (I138908,I138914,I138935,I138917,I138932,I138911,I138926,I138920,I138929,I138923,I138908,I138981,I138984,I138987,I138990,I138993,I138996,I138999,I139002,I2224,I2231);
PAT_5 I_1936 (I139002,I138981,I138990,I138984,I138999,I138996,I138987,I138987,I138981,I138984,I138993,I139048,I139051,I139054,I139057,I139060,I139063,I139066,I139069,I139072,I139075,I2224,I2231);
PAT_8 I_1937 (I139048,I139075,I139066,I139063,I139057,I139048,I139060,I139072,I139051,I139069,I139054,I139121,I139124,I139127,I139130,I139133,I139136,I139139,I139142,I139145,I2224,I2231);
PAT_9 I_1938 (I139124,I139133,I139124,I139121,I139136,I139127,I139142,I139130,I139139,I139121,I139145,I139191,I139194,I139197,I139200,I139203,I139206,I139209,I139212,I139215,I2224,I2231);
PAT_15 I_1939 (I139203,I139212,I139215,I139194,I139209,I139197,I139200,I139191,I139206,I139191,I139194,I139261,I139264,I139267,I139270,I139273,I139276,I139279,I139282,I139285,I2224,I2231);
PAT_12 I_1940 (I139279,I139282,I139285,I139273,I139270,I139264,I139261,I139276,I139267,I139261,I139264,I139331,I139334,I139337,I139340,I139343,I139346,I139349,I139352,I2224,I2231);
PAT_8 I_1941 (I139331,I139340,I139337,I139334,I139346,I139331,I139334,I139337,I139349,I139343,I139352,I139398,I139401,I139404,I139407,I139410,I139413,I139416,I139419,I139422,I2224,I2231);
PAT_10 I_1942 (I139404,I139398,I139401,I139422,I139416,I139401,I139410,I139398,I139419,I139413,I139407,I139468,I139471,I139474,I139477,I139480,I139483,I139486,I139489,I2224,I2231);
PAT_4 I_1943 (I139483,I139480,I139471,I139489,I139468,I139471,I139477,I139474,I139486,I139468,I139474,I139535,I139538,I139541,I139544,I139547,I139550,I139553,I139556,I139559,I2224,I2231);
PAT_17 I_1944 (I139547,I139544,I139556,I139550,I139535,I139553,I139559,I139538,I139541,I139538,I139535,I139605,I139608,I139611,I139614,I139617,I139620,I139623,I139626,I139629,I139632,I2224,I2231);
PAT_13 I_1945 (I139623,I139626,I139611,I139605,I139617,I139629,I139608,I139620,I139605,I139632,I139614,I139678,I139681,I139684,I139687,I139690,I139693,I139696,I139699,I139702,I2224,I2231);
PAT_16 I_1946 (I139684,I139687,I139696,I139690,I139702,I139678,I139699,I139693,I139681,I139681,I139678,I139748,I139751,I139754,I139757,I139760,I139763,I139766,I139769,I139772,I139775,I2224,I2231);
PAT_15 I_1947 (I139772,I139748,I139769,I139763,I139754,I139757,I139748,I139751,I139775,I139766,I139760,I139821,I139824,I139827,I139830,I139833,I139836,I139839,I139842,I139845,I2224,I2231);
PAT_10 I_1948 (I139824,I139833,I139827,I139821,I139842,I139845,I139830,I139821,I139824,I139839,I139836,I139891,I139894,I139897,I139900,I139903,I139906,I139909,I139912,I2224,I2231);
PAT_2 I_1949 (I139903,I139906,I139897,I139909,I139894,I139891,I139891,I139897,I139912,I139900,I139894,I139958,I139961,I139964,I139967,I139970,I139973,I139976,I139979,I139982,I2224,I2231);
PAT_4 I_1950 (I139958,I139964,I139982,I139976,I139973,I139970,I139961,I139979,I139958,I139961,I139967,I140028,I140031,I140034,I140037,I140040,I140043,I140046,I140049,I140052,I2224,I2231);
PAT_13 I_1951 (I140043,I140037,I140049,I140034,I140040,I140028,I140052,I140046,I140031,I140028,I140031,I140098,I140101,I140104,I140107,I140110,I140113,I140116,I140119,I140122,I2224,I2231);
PAT_14 I_1952 (I140101,I140116,I140104,I140113,I140107,I140098,I140110,I140119,I140098,I140122,I140101,I140168,I140171,I140174,I140177,I140180,I140183,I140186,I140189,I140192,I2224,I2231);
PAT_6 I_1953 (I1849,I2209,I1449,I2145,I1521,I2113,I2129,I1953,I2193,I1873,I1945,I140238,I140241,I140244,I140247,I140250,I140253,I140256,I140259,I140262,I140265,I2224,I2231);
PAT_2 I_1954 (I140259,I140265,I140247,I140253,I140238,I140244,I140238,I140250,I140241,I140256,I140262,I140311,I140314,I140317,I140320,I140323,I140326,I140329,I140332,I140335,I2224,I2231);
PAT_6 I_1955 (I140335,I140311,I140326,I140323,I140329,I140320,I140314,I140332,I140311,I140317,I140314,I140381,I140384,I140387,I140390,I140393,I140396,I140399,I140402,I140405,I140408,I2224,I2231);
PAT_14 I_1956 (I140393,I140387,I140381,I140408,I140390,I140384,I140396,I140399,I140381,I140405,I140402,I140454,I140457,I140460,I140463,I140466,I140469,I140472,I140475,I140478,I2224,I2231);
PAT_10 I_1957 (I140457,I140454,I140460,I140478,I140475,I140469,I140457,I140472,I140454,I140466,I140463,I140524,I140527,I140530,I140533,I140536,I140539,I140542,I140545,I2224,I2231);
PAT_5 I_1958 (I140545,I140524,I140533,I140527,I140542,I140539,I140530,I140530,I140524,I140527,I140536,I140591,I140594,I140597,I140600,I140603,I140606,I140609,I140612,I140615,I140618,I2224,I2231);
PAT_4 I_1959 (I140609,I140615,I140618,I140597,I140600,I140612,I140594,I140591,I140603,I140606,I140591,I140664,I140667,I140670,I140673,I140676,I140679,I140682,I140685,I140688,I2224,I2231);
PAT_10 I_1960 (I140664,I140664,I140688,I140667,I140673,I140682,I140679,I140667,I140685,I140670,I140676,I140734,I140737,I140740,I140743,I140746,I140749,I140752,I140755,I2224,I2231);
PAT_9 I_1961 (I140746,I140734,I140737,I140740,I140734,I140740,I140743,I140737,I140755,I140749,I140752,I140801,I140804,I140807,I140810,I140813,I140816,I140819,I140822,I140825,I2224,I2231);
PAT_13 I_1962 (I140801,I140822,I140804,I140819,I140813,I140810,I140825,I140801,I140807,I140816,I140804,I140871,I140874,I140877,I140880,I140883,I140886,I140889,I140892,I140895,I2224,I2231);
PAT_1 I_1963 (I140871,I140880,I140874,I140892,I140886,I140877,I140889,I140883,I140874,I140895,I140871,I140941,I140944,I140947,I140950,I140953,I140956,I140959,I140962,I140965,I2224,I2231);
PAT_8 I_1964 (I140962,I140944,I140950,I140941,I140959,I140953,I140956,I140941,I140965,I140947,I140944,I141011,I141014,I141017,I141020,I141023,I141026,I141029,I141032,I141035,I2224,I2231);
PAT_11 I_1965 (I141032,I141023,I141011,I141014,I141029,I141017,I141020,I141011,I141035,I141026,I141014,I141081,I141084,I141087,I141090,I141093,I141096,I141099,I141102,I141105,I141108,I2224,I2231);
PAT_17 I_1966 (I141093,I141084,I141108,I141081,I141090,I141102,I141099,I141096,I141081,I141105,I141087,I141154,I141157,I141160,I141163,I141166,I141169,I141172,I141175,I141178,I141181,I2224,I2231);
PAT_13 I_1967 (I141172,I141175,I141160,I141154,I141166,I141178,I141157,I141169,I141154,I141181,I141163,I141227,I141230,I141233,I141236,I141239,I141242,I141245,I141248,I141251,I2224,I2231);
PAT_5 I_1968 (I141239,I141230,I141236,I141248,I141230,I141251,I141233,I141242,I141227,I141227,I141245,I141297,I141300,I141303,I141306,I141309,I141312,I141315,I141318,I141321,I141324,I2224,I2231);
PAT_11 I_1969 (I141309,I141306,I141300,I141318,I141321,I141297,I141315,I141312,I141324,I141303,I141297,I141370,I141373,I141376,I141379,I141382,I141385,I141388,I141391,I141394,I141397,I2224,I2231);
PAT_13 I_1970 (I141370,I141373,I141382,I141394,I141397,I141385,I141391,I141379,I141388,I141376,I141370,I141443,I141446,I141449,I141452,I141455,I141458,I141461,I141464,I141467,I2224,I2231);
PAT_14 I_1971 (I141446,I141461,I141449,I141458,I141452,I141443,I141455,I141464,I141443,I141467,I141446,I141513,I141516,I141519,I141522,I141525,I141528,I141531,I141534,I141537,I2224,I2231);
PAT_4 I_1972 (I141522,I141528,I141519,I141513,I141537,I141525,I141513,I141516,I141534,I141516,I141531,I141583,I141586,I141589,I141592,I141595,I141598,I141601,I141604,I141607,I2224,I2231);
PAT_11 I_1973 (I141595,I141604,I141586,I141598,I141583,I141586,I141583,I141592,I141607,I141601,I141589,I141653,I141656,I141659,I141662,I141665,I141668,I141671,I141674,I141677,I141680,I2224,I2231);
PAT_8 I_1974 (I141662,I141668,I141671,I141677,I141674,I141665,I141653,I141653,I141680,I141656,I141659,I141726,I141729,I141732,I141735,I141738,I141741,I141744,I141747,I141750,I2224,I2231);
PAT_2 I_1975 (I141729,I141744,I141750,I141726,I141738,I141741,I141729,I141747,I141732,I141735,I141726,I141796,I141799,I141802,I141805,I141808,I141811,I141814,I141817,I141820,I2224,I2231);
PAT_13 I_1976 (I141805,I141799,I141796,I141817,I141808,I141811,I141799,I141802,I141814,I141820,I141796,I141866,I141869,I141872,I141875,I141878,I141881,I141884,I141887,I141890,I2224,I2231);
PAT_11 I_1977 (I141866,I141878,I141881,I141872,I141869,I141890,I141869,I141887,I141875,I141866,I141884,I141936,I141939,I141942,I141945,I141948,I141951,I141954,I141957,I141960,I141963,I2224,I2231);
PAT_9 I_1978 (I141942,I141954,I141945,I141957,I141936,I141939,I141948,I141936,I141951,I141960,I141963,I142009,I142012,I142015,I142018,I142021,I142024,I142027,I142030,I142033,I2224,I2231);
PAT_5 I_1979 (I142030,I142009,I142024,I142009,I142015,I142018,I142012,I142012,I142027,I142021,I142033,I142079,I142082,I142085,I142088,I142091,I142094,I142097,I142100,I142103,I142106,I2224,I2231);
PAT_15 I_1980 (I142097,I142082,I142079,I142079,I142094,I142091,I142103,I142088,I142100,I142085,I142106,I142152,I142155,I142158,I142161,I142164,I142167,I142170,I142173,I142176,I2224,I2231);
PAT_9 I_1981 (I142152,I142173,I142161,I142155,I142167,I142155,I142170,I142176,I142158,I142152,I142164,I142222,I142225,I142228,I142231,I142234,I142237,I142240,I142243,I142246,I2224,I2231);
PAT_13 I_1982 (I142222,I142243,I142225,I142240,I142234,I142231,I142246,I142222,I142228,I142237,I142225,I142292,I142295,I142298,I142301,I142304,I142307,I142310,I142313,I142316,I2224,I2231);
PAT_10 I_1983 (I142313,I142307,I142301,I142295,I142316,I142295,I142304,I142292,I142292,I142310,I142298,I142362,I142365,I142368,I142371,I142374,I142377,I142380,I142383,I2224,I2231);
PAT_6 I_1984 (I142383,I142377,I142371,I142365,I142362,I142368,I142362,I142368,I142365,I142374,I142380,I142429,I142432,I142435,I142438,I142441,I142444,I142447,I142450,I142453,I142456,I2224,I2231);
PAT_10 I_1985 (I142429,I142444,I142447,I142438,I142429,I142453,I142456,I142432,I142441,I142435,I142450,I142502,I142505,I142508,I142511,I142514,I142517,I142520,I142523,I2224,I2231);
PAT_2 I_1986 (I142514,I142517,I142508,I142520,I142505,I142502,I142502,I142508,I142523,I142511,I142505,I142569,I142572,I142575,I142578,I142581,I142584,I142587,I142590,I142593,I2224,I2231);
PAT_5 I_1987 (I142590,I142569,I142569,I142581,I142578,I142587,I142575,I142584,I142593,I142572,I142572,I142639,I142642,I142645,I142648,I142651,I142654,I142657,I142660,I142663,I142666,I2224,I2231);
PAT_17 I_1988 (I142666,I142642,I142645,I142648,I142639,I142651,I142639,I142663,I142657,I142654,I142660,I142712,I142715,I142718,I142721,I142724,I142727,I142730,I142733,I142736,I142739,I2224,I2231);
PAT_9 I_1989 (I142733,I142715,I142721,I142736,I142718,I142730,I142712,I142724,I142712,I142739,I142727,I142785,I142788,I142791,I142794,I142797,I142800,I142803,I142806,I142809,I2224,I2231);
PAT_13 I_1990 (I142785,I142806,I142788,I142803,I142797,I142794,I142809,I142785,I142791,I142800,I142788,I142855,I142858,I142861,I142864,I142867,I142870,I142873,I142876,I142879,I2224,I2231);
PAT_11 I_1991 (I142855,I142867,I142870,I142861,I142858,I142879,I142858,I142876,I142864,I142855,I142873,I142925,I142928,I142931,I142934,I142937,I142940,I142943,I142946,I142949,I142952,I2224,I2231);
PAT_9 I_1992 (I142931,I142943,I142934,I142946,I142925,I142928,I142937,I142925,I142940,I142949,I142952,I142998,I143001,I143004,I143007,I143010,I143013,I143016,I143019,I143022,I2224,I2231);
PAT_13 I_1993 (I142998,I143019,I143001,I143016,I143010,I143007,I143022,I142998,I143004,I143013,I143001,I143068,I143071,I143074,I143077,I143080,I143083,I143086,I143089,I143092,I2224,I2231);
PAT_5 I_1994 (I143080,I143071,I143077,I143089,I143071,I143092,I143074,I143083,I143068,I143068,I143086,I143138,I143141,I143144,I143147,I143150,I143153,I143156,I143159,I143162,I143165,I2224,I2231);
PAT_1 I_1995 (I143153,I143141,I143159,I143138,I143144,I143138,I143147,I143162,I143156,I143165,I143150,I143211,I143214,I143217,I143220,I143223,I143226,I143229,I143232,I143235,I2224,I2231);
PAT_2 I_1996 (I143211,I143217,I143211,I143226,I143214,I143214,I143220,I143223,I143229,I143235,I143232,I143281,I143284,I143287,I143290,I143293,I143296,I143299,I143302,I143305,I2224,I2231);
PAT_5 I_1997 (I143302,I143281,I143281,I143293,I143290,I143299,I143287,I143296,I143305,I143284,I143284,I143351,I143354,I143357,I143360,I143363,I143366,I143369,I143372,I143375,I143378,I2224,I2231);
PAT_15 I_1998 (I143369,I143354,I143351,I143351,I143366,I143363,I143375,I143360,I143372,I143357,I143378,I143424,I143427,I143430,I143433,I143436,I143439,I143442,I143445,I143448,I2224,I2231);
PAT_4 I_1999 (I143436,I143442,I143424,I143427,I143430,I143424,I143448,I143445,I143433,I143439,I143427,I143494,I143497,I143500,I143503,I143506,I143509,I143512,I143515,I143518,I2224,I2231);
PAT_8 I_2000 (I143506,I143494,I143515,I143500,I143497,I143518,I143503,I143512,I143497,I143494,I143509,I143564,I143567,I143570,I143573,I143576,I143579,I143582,I143585,I143588,I2224,I2231);
PAT_13 I_2001 (I143576,I143585,I143567,I143588,I143570,I143564,I143564,I143573,I143582,I143579,I143567,I143634,I143637,I143640,I143643,I143646,I143649,I143652,I143655,I143658,I2224,I2231);
PAT_9 I_2002 (I143655,I143637,I143637,I143634,I143658,I143640,I143643,I143634,I143646,I143652,I143649,I143704,I143707,I143710,I143713,I143716,I143719,I143722,I143725,I143728,I2224,I2231);
PAT_6 I_2003 (I143722,I143704,I143716,I143725,I143704,I143713,I143710,I143728,I143719,I143707,I143707,I143774,I143777,I143780,I143783,I143786,I143789,I143792,I143795,I143798,I143801,I2224,I2231);
PAT_2 I_2004 (I143795,I143801,I143783,I143789,I143774,I143780,I143774,I143786,I143777,I143792,I143798,I143847,I143850,I143853,I143856,I143859,I143862,I143865,I143868,I143871,I2224,I2231);
PAT_4 I_2005 (I143847,I143853,I143871,I143865,I143862,I143859,I143850,I143868,I143847,I143850,I143856,I143917,I143920,I143923,I143926,I143929,I143932,I143935,I143938,I143941,I2224,I2231);
PAT_5 I_2006 (I143938,I143920,I143920,I143932,I143935,I143929,I143926,I143917,I143923,I143917,I143941,I143987,I143990,I143993,I143996,I143999,I144002,I144005,I144008,I144011,I144014,I2224,I2231);
PAT_13 I_2007 (I143993,I144002,I143987,I143990,I144011,I143996,I144008,I143987,I144005,I144014,I143999,I144060,I144063,I144066,I144069,I144072,I144075,I144078,I144081,I144084,I2224,I2231);
PAT_2 I_2008 (I144078,I144072,I144069,I144075,I144060,I144084,I144063,I144081,I144060,I144066,I144063,I144130,I144133,I144136,I144139,I144142,I144145,I144148,I144151,I144154,I2224,I2231);
PAT_4 I_2009 (I144130,I144136,I144154,I144148,I144145,I144142,I144133,I144151,I144130,I144133,I144139,I144200,I144203,I144206,I144209,I144212,I144215,I144218,I144221,I144224,I2224,I2231);
PAT_8 I_2010 (I144212,I144200,I144221,I144206,I144203,I144224,I144209,I144218,I144203,I144200,I144215,I144270,I144273,I144276,I144279,I144282,I144285,I144288,I144291,I144294,I2224,I2231);
PAT_2 I_2011 (I144273,I144288,I144294,I144270,I144282,I144285,I144273,I144291,I144276,I144279,I144270,I144340,I144343,I144346,I144349,I144352,I144355,I144358,I144361,I144364,I2224,I2231);
PAT_4 I_2012 (I144340,I144346,I144364,I144358,I144355,I144352,I144343,I144361,I144340,I144343,I144349,I144410,I144413,I144416,I144419,I144422,I144425,I144428,I144431,I144434,I2224,I2231);
PAT_1 I_2013 (I144410,I144431,I144428,I144413,I144425,I144410,I144413,I144434,I144419,I144416,I144422,I144480,I144483,I144486,I144489,I144492,I144495,I144498,I144501,I144504,I2224,I2231);
PAT_5 I_2014 (I144498,I144501,I144483,I144492,I144489,I144486,I144495,I144504,I144483,I144480,I144480,I144550,I144553,I144556,I144559,I144562,I144565,I144568,I144571,I144574,I144577,I2224,I2231);
PAT_17 I_2015 (I144577,I144553,I144556,I144559,I144550,I144562,I144550,I144574,I144568,I144565,I144571,I144623,I144626,I144629,I144632,I144635,I144638,I144641,I144644,I144647,I144650,I2224,I2231);
PAT_2 I_2016 (I144623,I144641,I144638,I144623,I144632,I144647,I144644,I144629,I144650,I144635,I144626,I144696,I144699,I144702,I144705,I144708,I144711,I144714,I144717,I144720,I2224,I2231);
PAT_9 I_2017 (I144711,I144720,I144696,I144702,I144705,I144714,I144699,I144708,I144717,I144699,I144696,I144766,I144769,I144772,I144775,I144778,I144781,I144784,I144787,I144790,I2224,I2231);
PAT_11 I_2018 (I144778,I144784,I144790,I144787,I144775,I144769,I144769,I144766,I144781,I144766,I144772,I144836,I144839,I144842,I144845,I144848,I144851,I144854,I144857,I144860,I144863,I2224,I2231);
PAT_9 I_2019 (I144842,I144854,I144845,I144857,I144836,I144839,I144848,I144836,I144851,I144860,I144863,I144909,I144912,I144915,I144918,I144921,I144924,I144927,I144930,I144933,I2224,I2231);
PAT_12 I_2020 (I144930,I144927,I144921,I144909,I144918,I144909,I144912,I144915,I144933,I144924,I144912,I144979,I144982,I144985,I144988,I144991,I144994,I144997,I145000,I2224,I2231);
PAT_8 I_2021 (I144979,I144988,I144985,I144982,I144994,I144979,I144982,I144985,I144997,I144991,I145000,I145046,I145049,I145052,I145055,I145058,I145061,I145064,I145067,I145070,I2224,I2231);
PAT_14 I_2022 (I145052,I145064,I145049,I145046,I145049,I145070,I145046,I145058,I145061,I145067,I145055,I145116,I145119,I145122,I145125,I145128,I145131,I145134,I145137,I145140,I2224,I2231);
PAT_6 I_2023 (I145116,I145119,I145140,I145125,I145116,I145122,I145128,I145131,I145134,I145119,I145137,I145186,I145189,I145192,I145195,I145198,I145201,I145204,I145207,I145210,I145213,I2224,I2231);
PAT_13 I_2024 (I145210,I145192,I145207,I145186,I145189,I145195,I145213,I145198,I145204,I145186,I145201,I145259,I145262,I145265,I145268,I145271,I145274,I145277,I145280,I145283,I2224,I2231);
PAT_4 I_2025 (I145268,I145271,I145283,I145265,I145280,I145277,I145262,I145274,I145262,I145259,I145259,I145329,I145332,I145335,I145338,I145341,I145344,I145347,I145350,I145353,I2224,I2231);
PAT_2 I_2026 (I145338,I145332,I145332,I145353,I145329,I145347,I145344,I145335,I145329,I145341,I145350,I145399,I145402,I145405,I145408,I145411,I145414,I145417,I145420,I145423,I2224,I2231);
PAT_9 I_2027 (I145414,I145423,I145399,I145405,I145408,I145417,I145402,I145411,I145420,I145402,I145399,I145469,I145472,I145475,I145478,I145481,I145484,I145487,I145490,I145493,I2224,I2231);
PAT_13 I_2028 (I145469,I145490,I145472,I145487,I145481,I145478,I145493,I145469,I145475,I145484,I145472,I145539,I145542,I145545,I145548,I145551,I145554,I145557,I145560,I145563,I2224,I2231);
PAT_8 I_2029 (I145548,I145560,I145551,I145554,I145563,I145542,I145557,I145539,I145542,I145545,I145539,I145609,I145612,I145615,I145618,I145621,I145624,I145627,I145630,I145633,I2224,I2231);
PAT_14 I_2030 (I145615,I145627,I145612,I145609,I145612,I145633,I145609,I145621,I145624,I145630,I145618,I145679,I145682,I145685,I145688,I145691,I145694,I145697,I145700,I145703,I2224,I2231);
PAT_12 I_2031 (I145688,I145694,I145679,I145703,I145682,I145682,I145697,I145679,I145700,I145691,I145685,I145749,I145752,I145755,I145758,I145761,I145764,I145767,I145770,I2224,I2231);
PAT_6 I_2032 (I145758,I145752,I145770,I145755,I145752,I145755,I145764,I145749,I145767,I145749,I145761,I145816,I145819,I145822,I145825,I145828,I145831,I145834,I145837,I145840,I145843,I2224,I2231);
PAT_12 I_2033 (I145816,I145843,I145822,I145825,I145819,I145816,I145837,I145831,I145834,I145828,I145840,I145889,I145892,I145895,I145898,I145901,I145904,I145907,I145910,I2224,I2231);
PAT_9 I_2034 (I145898,I145904,I145889,I145895,I145901,I145892,I145889,I145892,I145910,I145895,I145907,I145956,I145959,I145962,I145965,I145968,I145971,I145974,I145977,I145980,I2224,I2231);
PAT_6 I_2035 (I145974,I145956,I145968,I145977,I145956,I145965,I145962,I145980,I145971,I145959,I145959,I146026,I146029,I146032,I146035,I146038,I146041,I146044,I146047,I146050,I146053,I2224,I2231);
PAT_17 I_2036 (I146038,I146041,I146047,I146035,I146029,I146050,I146044,I146026,I146053,I146032,I146026,I146099,I146102,I146105,I146108,I146111,I146114,I146117,I146120,I146123,I146126,I2224,I2231);
PAT_5 I_2037 (I146111,I146105,I146102,I146123,I146108,I146114,I146117,I146099,I146099,I146120,I146126,I146172,I146175,I146178,I146181,I146184,I146187,I146190,I146193,I146196,I146199,I2224,I2231);
PAT_9 I_2038 (I146187,I146184,I146193,I146190,I146181,I146172,I146178,I146199,I146175,I146196,I146172,I146245,I146248,I146251,I146254,I146257,I146260,I146263,I146266,I146269,I2224,I2231);
PAT_13 I_2039 (I146245,I146266,I146248,I146263,I146257,I146254,I146269,I146245,I146251,I146260,I146248,I146315,I146318,I146321,I146324,I146327,I146330,I146333,I146336,I146339,I2224,I2231);
PAT_11 I_2040 (I146315,I146327,I146330,I146321,I146318,I146339,I146318,I146336,I146324,I146315,I146333,I146385,I146388,I146391,I146394,I146397,I146400,I146403,I146406,I146409,I146412,I2224,I2231);
PAT_4 I_2041 (I146391,I146412,I146385,I146403,I146394,I146385,I146406,I146388,I146397,I146409,I146400,I146458,I146461,I146464,I146467,I146470,I146473,I146476,I146479,I146482,I2224,I2231);
PAT_9 I_2042 (I146479,I146461,I146464,I146473,I146476,I146458,I146467,I146461,I146482,I146458,I146470,I146528,I146531,I146534,I146537,I146540,I146543,I146546,I146549,I146552,I2224,I2231);
PAT_10 I_2043 (I146549,I146546,I146534,I146531,I146552,I146537,I146543,I146531,I146528,I146528,I146540,I146598,I146601,I146604,I146607,I146610,I146613,I146616,I146619,I2224,I2231);
PAT_4 I_2044 (I146613,I146610,I146601,I146619,I146598,I146601,I146607,I146604,I146616,I146598,I146604,I146665,I146668,I146671,I146674,I146677,I146680,I146683,I146686,I146689,I2224,I2231);
PAT_13 I_2045 (I146680,I146674,I146686,I146671,I146677,I146665,I146689,I146683,I146668,I146665,I146668,I146735,I146738,I146741,I146744,I146747,I146750,I146753,I146756,I146759,I2224,I2231);
PAT_17 I_2046 (I146759,I146747,I146756,I146753,I146744,I146735,I146738,I146741,I146735,I146750,I146738,I146805,I146808,I146811,I146814,I146817,I146820,I146823,I146826,I146829,I146832,I2224,I2231);
PAT_11 I_2047 (I146817,I146826,I146832,I146808,I146805,I146823,I146814,I146820,I146811,I146829,I146805,I146878,I146881,I146884,I146887,I146890,I146893,I146896,I146899,I146902,I146905,I2224,I2231);
PAT_17 I_2048 (I146890,I146881,I146905,I146878,I146887,I146899,I146896,I146893,I146878,I146902,I146884,I146951,I146954,I146957,I146960,I146963,I146966,I146969,I146972,I146975,I146978,I2224,I2231);
PAT_9 I_2049 (I146972,I146954,I146960,I146975,I146957,I146969,I146951,I146963,I146951,I146978,I146966,I147024,I147027,I147030,I147033,I147036,I147039,I147042,I147045,I147048,I2224,I2231);
PAT_13 I_2050 (I147024,I147045,I147027,I147042,I147036,I147033,I147048,I147024,I147030,I147039,I147027,I147094,I147097,I147100,I147103,I147106,I147109,I147112,I147115,I147118,I2224,I2231);
PAT_17 I_2051 (I147118,I147106,I147115,I147112,I147103,I147094,I147097,I147100,I147094,I147109,I147097,I147164,I147167,I147170,I147173,I147176,I147179,I147182,I147185,I147188,I147191,I2224,I2231);
PAT_6 I_2052 (I147164,I147182,I147170,I147173,I147179,I147164,I147176,I147167,I147188,I147191,I147185,I147237,I147240,I147243,I147246,I147249,I147252,I147255,I147258,I147261,I147264,I2224,I2231);
PAT_0 I_2053 (I147237,I147255,I147249,I147261,I147243,I147264,I147246,I147237,I147252,I147258,I147240,I147310,I147313,I147316,I147319,I147322,I147325,I147328,I147331,I2224,I2231);
PAT_8 I_2054 (I147331,I147325,I147328,I147313,I147313,I147316,I147310,I147319,I147316,I147310,I147322,I147377,I147380,I147383,I147386,I147389,I147392,I147395,I147398,I147401,I2224,I2231);
PAT_6 I_2055 (I147380,I147377,I147383,I147395,I147392,I147386,I147389,I147377,I147398,I147380,I147401,I147447,I147450,I147453,I147456,I147459,I147462,I147465,I147468,I147471,I147474,I2224,I2231);
PAT_13 I_2056 (I147471,I147453,I147468,I147447,I147450,I147456,I147474,I147459,I147465,I147447,I147462,I147520,I147523,I147526,I147529,I147532,I147535,I147538,I147541,I147544,I2224,I2231);
PAT_5 I_2057 (I147532,I147523,I147529,I147541,I147523,I147544,I147526,I147535,I147520,I147520,I147538,I147590,I147593,I147596,I147599,I147602,I147605,I147608,I147611,I147614,I147617,I2224,I2231);
PAT_10 I_2058 (I147614,I147617,I147596,I147602,I147605,I147611,I147593,I147590,I147590,I147599,I147608,I147663,I147666,I147669,I147672,I147675,I147678,I147681,I147684,I2224,I2231);
PAT_6 I_2059 (I147684,I147678,I147672,I147666,I147663,I147669,I147663,I147669,I147666,I147675,I147681,I147730,I147733,I147736,I147739,I147742,I147745,I147748,I147751,I147754,I147757,I2224,I2231);
PAT_2 I_2060 (I147751,I147757,I147739,I147745,I147730,I147736,I147730,I147742,I147733,I147748,I147754,I147803,I147806,I147809,I147812,I147815,I147818,I147821,I147824,I147827,I2224,I2231);
PAT_13 I_2061 (I147812,I147806,I147803,I147824,I147815,I147818,I147806,I147809,I147821,I147827,I147803,I147873,I147876,I147879,I147882,I147885,I147888,I147891,I147894,I147897,I2224,I2231);
PAT_5 I_2062 (I147885,I147876,I147882,I147894,I147876,I147897,I147879,I147888,I147873,I147873,I147891,I147943,I147946,I147949,I147952,I147955,I147958,I147961,I147964,I147967,I147970,I2224,I2231);
PAT_11 I_2063 (I147955,I147952,I147946,I147964,I147967,I147943,I147961,I147958,I147970,I147949,I147943,I148016,I148019,I148022,I148025,I148028,I148031,I148034,I148037,I148040,I148043,I2224,I2231);
PAT_6 I_2064 (I148016,I148043,I148031,I148040,I148034,I148028,I148019,I148037,I148025,I148022,I148016,I148089,I148092,I148095,I148098,I148101,I148104,I148107,I148110,I148113,I148116,I2224,I2231);
PAT_1 I_2065 (I148116,I148107,I148095,I148098,I148110,I148101,I148104,I148089,I148092,I148089,I148113,I148162,I148165,I148168,I148171,I148174,I148177,I148180,I148183,I148186,I2224,I2231);
PAT_9 I_2066 (I148177,I148183,I148168,I148186,I148165,I148180,I148165,I148171,I148162,I148174,I148162,I148232,I148235,I148238,I148241,I148244,I148247,I148250,I148253,I148256,I2224,I2231);
PAT_15 I_2067 (I148244,I148253,I148256,I148235,I148250,I148238,I148241,I148232,I148247,I148232,I148235,I148302,I148305,I148308,I148311,I148314,I148317,I148320,I148323,I148326,I2224,I2231);
PAT_1 I_2068 (I148308,I148305,I148305,I148302,I148302,I148311,I148326,I148320,I148314,I148317,I148323,I148372,I148375,I148378,I148381,I148384,I148387,I148390,I148393,I148396,I2224,I2231);
PAT_11 I_2069 (I148375,I148390,I148387,I148393,I148396,I148375,I148381,I148384,I148372,I148378,I148372,I148442,I148445,I148448,I148451,I148454,I148457,I148460,I148463,I148466,I148469,I2224,I2231);
PAT_14 I_2070 (I148463,I148451,I148445,I148466,I148457,I148460,I148448,I148469,I148454,I148442,I148442,I148515,I148518,I148521,I148524,I148527,I148530,I148533,I148536,I148539,I2224,I2231);
PAT_1 I_2071 (I148515,I148539,I148524,I148518,I148518,I148521,I148530,I148533,I148527,I148515,I148536,I148585,I148588,I148591,I148594,I148597,I148600,I148603,I148606,I148609,I2224,I2231);
PAT_6 I_2072 (I148594,I148585,I148588,I148591,I148606,I148609,I148603,I148585,I148600,I148597,I148588,I148655,I148658,I148661,I148664,I148667,I148670,I148673,I148676,I148679,I148682,I2224,I2231);
PAT_12 I_2073 (I148655,I148682,I148661,I148664,I148658,I148655,I148676,I148670,I148673,I148667,I148679,I148728,I148731,I148734,I148737,I148740,I148743,I148746,I148749,I2224,I2231);
PAT_6 I_2074 (I148737,I148731,I148749,I148734,I148731,I148734,I148743,I148728,I148746,I148728,I148740,I148795,I148798,I148801,I148804,I148807,I148810,I148813,I148816,I148819,I148822,I2224,I2231);
PAT_2 I_2075 (I148816,I148822,I148804,I148810,I148795,I148801,I148795,I148807,I148798,I148813,I148819,I148868,I148871,I148874,I148877,I148880,I148883,I148886,I148889,I148892,I2224,I2231);
PAT_13 I_2076 (I148877,I148871,I148868,I148889,I148880,I148883,I148871,I148874,I148886,I148892,I148868,I148938,I148941,I148944,I148947,I148950,I148953,I148956,I148959,I148962,I2224,I2231);
PAT_6 I_2077 (I148938,I148950,I148947,I148959,I148956,I148962,I148938,I148953,I148941,I148941,I148944,I149008,I149011,I149014,I149017,I149020,I149023,I149026,I149029,I149032,I149035,I2224,I2231);
PAT_9 I_2078 (I149008,I149035,I149032,I149014,I149020,I149011,I149023,I149008,I149026,I149017,I149029,I149081,I149084,I149087,I149090,I149093,I149096,I149099,I149102,I149105,I2224,I2231);
PAT_13 I_2079 (I149081,I149102,I149084,I149099,I149093,I149090,I149105,I149081,I149087,I149096,I149084,I149151,I149154,I149157,I149160,I149163,I149166,I149169,I149172,I149175,I2224,I2231);
PAT_4 I_2080 (I149160,I149163,I149175,I149157,I149172,I149169,I149154,I149166,I149154,I149151,I149151,I149221,I149224,I149227,I149230,I149233,I149236,I149239,I149242,I149245,I2224,I2231);
PAT_10 I_2081 (I149221,I149221,I149245,I149224,I149230,I149239,I149236,I149224,I149242,I149227,I149233,I149291,I149294,I149297,I149300,I149303,I149306,I149309,I149312,I2224,I2231);
PAT_5 I_2082 (I149312,I149291,I149300,I149294,I149309,I149306,I149297,I149297,I149291,I149294,I149303,I149358,I149361,I149364,I149367,I149370,I149373,I149376,I149379,I149382,I149385,I2224,I2231);
PAT_15 I_2083 (I149376,I149361,I149358,I149358,I149373,I149370,I149382,I149367,I149379,I149364,I149385,I149431,I149434,I149437,I149440,I149443,I149446,I149449,I149452,I149455,I2224,I2231);
PAT_10 I_2084 (I149434,I149443,I149437,I149431,I149452,I149455,I149440,I149431,I149434,I149449,I149446,I149501,I149504,I149507,I149510,I149513,I149516,I149519,I149522,I2224,I2231);
PAT_11 I_2085 (I149510,I149513,I149522,I149516,I149519,I149501,I149501,I149507,I149504,I149504,I149507,I149568,I149571,I149574,I149577,I149580,I149583,I149586,I149589,I149592,I149595,I2224,I2231);
PAT_5 I_2086 (I149589,I149568,I149595,I149583,I149580,I149592,I149574,I149568,I149586,I149571,I149577,I149641,I149644,I149647,I149650,I149653,I149656,I149659,I149662,I149665,I149668,I2224,I2231);
PAT_11 I_2087 (I149653,I149650,I149644,I149662,I149665,I149641,I149659,I149656,I149668,I149647,I149641,I149714,I149717,I149720,I149723,I149726,I149729,I149732,I149735,I149738,I149741,I2224,I2231);
PAT_2 I_2088 (I149714,I149738,I149726,I149720,I149729,I149732,I149717,I149741,I149735,I149723,I149714,I149787,I149790,I149793,I149796,I149799,I149802,I149805,I149808,I149811,I2224,I2231);
PAT_5 I_2089 (I149808,I149787,I149787,I149799,I149796,I149805,I149793,I149802,I149811,I149790,I149790,I149857,I149860,I149863,I149866,I149869,I149872,I149875,I149878,I149881,I149884,I2224,I2231);
PAT_2 I_2090 (I149872,I149857,I149869,I149863,I149878,I149860,I149875,I149866,I149881,I149884,I149857,I149930,I149933,I149936,I149939,I149942,I149945,I149948,I149951,I149954,I2224,I2231);
PAT_4 I_2091 (I149930,I149936,I149954,I149948,I149945,I149942,I149933,I149951,I149930,I149933,I149939,I150000,I150003,I150006,I150009,I150012,I150015,I150018,I150021,I150024,I2224,I2231);
PAT_2 I_2092 (I150009,I150003,I150003,I150024,I150000,I150018,I150015,I150006,I150000,I150012,I150021,I150070,I150073,I150076,I150079,I150082,I150085,I150088,I150091,I150094,I2224,I2231);
PAT_5 I_2093 (I150091,I150070,I150070,I150082,I150079,I150088,I150076,I150085,I150094,I150073,I150073,I150140,I150143,I150146,I150149,I150152,I150155,I150158,I150161,I150164,I150167,I2224,I2231);
PAT_2 I_2094 (I150155,I150140,I150152,I150146,I150161,I150143,I150158,I150149,I150164,I150167,I150140,I150213,I150216,I150219,I150222,I150225,I150228,I150231,I150234,I150237,I2224,I2231);
PAT_7 I_2095 (I150237,I150213,I150219,I150216,I150216,I150225,I150228,I150213,I150231,I150234,I150222,I150283,I150286,I150289,I150292,I150295,I150298,I150301,I150304,I150307,I2224,I2231);
PAT_13 I_2096 (I150289,I150307,I150298,I150283,I150295,I150283,I150304,I150286,I150292,I150286,I150301,I150353,I150356,I150359,I150362,I150365,I150368,I150371,I150374,I150377,I2224,I2231);
PAT_11 I_2097 (I150353,I150365,I150368,I150359,I150356,I150377,I150356,I150374,I150362,I150353,I150371,I150423,I150426,I150429,I150432,I150435,I150438,I150441,I150444,I150447,I150450,I2224,I2231);
PAT_13 I_2098 (I150423,I150426,I150435,I150447,I150450,I150438,I150444,I150432,I150441,I150429,I150423,I150496,I150499,I150502,I150505,I150508,I150511,I150514,I150517,I150520,I2224,I2231);
PAT_9 I_2099 (I150517,I150499,I150499,I150496,I150520,I150502,I150505,I150496,I150508,I150514,I150511,I150566,I150569,I150572,I150575,I150578,I150581,I150584,I150587,I150590,I2224,I2231);
PAT_1 I_2100 (I150566,I150584,I150566,I150578,I150569,I150575,I150581,I150587,I150590,I150572,I150569,I150636,I150639,I150642,I150645,I150648,I150651,I150654,I150657,I150660,I2224,I2231);
PAT_5 I_2101 (I150654,I150657,I150639,I150648,I150645,I150642,I150651,I150660,I150639,I150636,I150636,I150706,I150709,I150712,I150715,I150718,I150721,I150724,I150727,I150730,I150733,I2224,I2231);
PAT_10 I_2102 (I150730,I150733,I150712,I150718,I150721,I150727,I150709,I150706,I150706,I150715,I150724,I150779,I150782,I150785,I150788,I150791,I150794,I150797,I150800,I2224,I2231);
PAT_5 I_2103 (I150800,I150779,I150788,I150782,I150797,I150794,I150785,I150785,I150779,I150782,I150791,I150846,I150849,I150852,I150855,I150858,I150861,I150864,I150867,I150870,I150873,I2224,I2231);
PAT_13 I_2104 (I150852,I150861,I150846,I150849,I150870,I150855,I150867,I150846,I150864,I150873,I150858,I150919,I150922,I150925,I150928,I150931,I150934,I150937,I150940,I150943,I2224,I2231);
PAT_11 I_2105 (I150919,I150931,I150934,I150925,I150922,I150943,I150922,I150940,I150928,I150919,I150937,I150989,I150992,I150995,I150998,I151001,I151004,I151007,I151010,I151013,I151016,I2224,I2231);
PAT_2 I_2106 (I150989,I151013,I151001,I150995,I151004,I151007,I150992,I151016,I151010,I150998,I150989,I151062,I151065,I151068,I151071,I151074,I151077,I151080,I151083,I151086,I2224,I2231);
PAT_10 I_2107 (I151062,I151080,I151077,I151065,I151068,I151083,I151074,I151062,I151071,I151086,I151065,I151132,I151135,I151138,I151141,I151144,I151147,I151150,I151153,I2224,I2231);
PAT_9 I_2108 (I151144,I151132,I151135,I151138,I151132,I151138,I151141,I151135,I151153,I151147,I151150,I151199,I151202,I151205,I151208,I151211,I151214,I151217,I151220,I151223,I2224,I2231);
PAT_12 I_2109 (I151220,I151217,I151211,I151199,I151208,I151199,I151202,I151205,I151223,I151214,I151202,I151269,I151272,I151275,I151278,I151281,I151284,I151287,I151290,I2224,I2231);
PAT_10 I_2110 (I151269,I151290,I151281,I151284,I151275,I151272,I151269,I151287,I151275,I151278,I151272,I151336,I151339,I151342,I151345,I151348,I151351,I151354,I151357,I2224,I2231);
PAT_4 I_2111 (I151351,I151348,I151339,I151357,I151336,I151339,I151345,I151342,I151354,I151336,I151342,I151403,I151406,I151409,I151412,I151415,I151418,I151421,I151424,I151427,I2224,I2231);
PAT_11 I_2112 (I151415,I151424,I151406,I151418,I151403,I151406,I151403,I151412,I151427,I151421,I151409,I151473,I151476,I151479,I151482,I151485,I151488,I151491,I151494,I151497,I151500,I2224,I2231);
PAT_4 I_2113 (I151479,I151500,I151473,I151491,I151482,I151473,I151494,I151476,I151485,I151497,I151488,I151546,I151549,I151552,I151555,I151558,I151561,I151564,I151567,I151570,I2224,I2231);
PAT_13 I_2114 (I151561,I151555,I151567,I151552,I151558,I151546,I151570,I151564,I151549,I151546,I151549,I151616,I151619,I151622,I151625,I151628,I151631,I151634,I151637,I151640,I2224,I2231);
PAT_4 I_2115 (I151625,I151628,I151640,I151622,I151637,I151634,I151619,I151631,I151619,I151616,I151616,I151686,I151689,I151692,I151695,I151698,I151701,I151704,I151707,I151710,I2224,I2231);
PAT_10 I_2116 (I151686,I151686,I151710,I151689,I151695,I151704,I151701,I151689,I151707,I151692,I151698,I151756,I151759,I151762,I151765,I151768,I151771,I151774,I151777,I2224,I2231);
PAT_8 I_2117 (I151777,I151768,I151759,I151756,I151765,I151756,I151771,I151759,I151774,I151762,I151762,I151823,I151826,I151829,I151832,I151835,I151838,I151841,I151844,I151847,I2224,I2231);
PAT_12 I_2118 (I151823,I151826,I151826,I151847,I151832,I151841,I151844,I151835,I151829,I151838,I151823,I151893,I151896,I151899,I151902,I151905,I151908,I151911,I151914,I2224,I2231);
PAT_11 I_2119 (I151899,I151902,I151899,I151911,I151914,I151908,I151896,I151905,I151893,I151896,I151893,I151960,I151963,I151966,I151969,I151972,I151975,I151978,I151981,I151984,I151987,I2224,I2231);
PAT_8 I_2120 (I151969,I151975,I151978,I151984,I151981,I151972,I151960,I151960,I151987,I151963,I151966,I152033,I152036,I152039,I152042,I152045,I152048,I152051,I152054,I152057,I2224,I2231);
PAT_4 I_2121 (I152051,I152036,I152042,I152033,I152033,I152045,I152036,I152054,I152057,I152039,I152048,I152103,I152106,I152109,I152112,I152115,I152118,I152121,I152124,I152127,I2224,I2231);
PAT_7 I_2122 (I152118,I152112,I152109,I152103,I152115,I152121,I152106,I152106,I152124,I152127,I152103,I152173,I152176,I152179,I152182,I152185,I152188,I152191,I152194,I152197,I2224,I2231);
PAT_5 I_2123 (I152179,I152173,I152182,I152191,I152185,I152197,I152194,I152176,I152188,I152176,I152173,I152243,I152246,I152249,I152252,I152255,I152258,I152261,I152264,I152267,I152270,I2224,I2231);
PAT_10 I_2124 (I152267,I152270,I152249,I152255,I152258,I152264,I152246,I152243,I152243,I152252,I152261,I152316,I152319,I152322,I152325,I152328,I152331,I152334,I152337,I2224,I2231);
PAT_13 I_2125 (I152322,I152328,I152322,I152319,I152334,I152337,I152316,I152316,I152331,I152319,I152325,I152383,I152386,I152389,I152392,I152395,I152398,I152401,I152404,I152407,I2224,I2231);
PAT_6 I_2126 (I152383,I152395,I152392,I152404,I152401,I152407,I152383,I152398,I152386,I152386,I152389,I152453,I152456,I152459,I152462,I152465,I152468,I152471,I152474,I152477,I152480,I2224,I2231);
PAT_15 I_2127 (I152471,I152462,I152474,I152477,I152468,I152480,I152453,I152459,I152453,I152456,I152465,I152526,I152529,I152532,I152535,I152538,I152541,I152544,I152547,I152550,I2224,I2231);
PAT_6 I_2128 (I152529,I152526,I152532,I152547,I152529,I152550,I152535,I152541,I152538,I152544,I152526,I152596,I152599,I152602,I152605,I152608,I152611,I152614,I152617,I152620,I152623,I2224,I2231);
PAT_1 I_2129 (I152623,I152614,I152602,I152605,I152617,I152608,I152611,I152596,I152599,I152596,I152620,I152669,I152672,I152675,I152678,I152681,I152684,I152687,I152690,I152693,I2224,I2231);
PAT_9 I_2130 (I152684,I152690,I152675,I152693,I152672,I152687,I152672,I152678,I152669,I152681,I152669,I152739,I152742,I152745,I152748,I152751,I152754,I152757,I152760,I152763,I2224,I2231);
PAT_7 I_2131 (I152745,I152754,I152739,I152760,I152751,I152739,I152742,I152763,I152757,I152742,I152748,I152809,I152812,I152815,I152818,I152821,I152824,I152827,I152830,I152833,I2224,I2231);
PAT_13 I_2132 (I152815,I152833,I152824,I152809,I152821,I152809,I152830,I152812,I152818,I152812,I152827,I152879,I152882,I152885,I152888,I152891,I152894,I152897,I152900,I152903,I2224,I2231);
PAT_15 I_2133 (I152879,I152891,I152882,I152894,I152879,I152888,I152903,I152900,I152885,I152897,I152882,I152949,I152952,I152955,I152958,I152961,I152964,I152967,I152970,I152973,I2224,I2231);
PAT_12 I_2134 (I152967,I152970,I152973,I152961,I152958,I152952,I152949,I152964,I152955,I152949,I152952,I153019,I153022,I153025,I153028,I153031,I153034,I153037,I153040,I2224,I2231);
PAT_1 I_2135 (I153034,I153022,I153037,I153028,I153019,I153022,I153031,I153019,I153040,I153025,I153025,I153086,I153089,I153092,I153095,I153098,I153101,I153104,I153107,I153110,I2224,I2231);
PAT_4 I_2136 (I153098,I153104,I153086,I153089,I153092,I153095,I153107,I153089,I153101,I153086,I153110,I153156,I153159,I153162,I153165,I153168,I153171,I153174,I153177,I153180,I2224,I2231);
PAT_5 I_2137 (I153177,I153159,I153159,I153171,I153174,I153168,I153165,I153156,I153162,I153156,I153180,I153226,I153229,I153232,I153235,I153238,I153241,I153244,I153247,I153250,I153253,I2224,I2231);
PAT_7 I_2138 (I153244,I153247,I153253,I153250,I153235,I153232,I153226,I153238,I153226,I153229,I153241,I153299,I153302,I153305,I153308,I153311,I153314,I153317,I153320,I153323,I2224,I2231);
PAT_14 I_2139 (I153314,I153308,I153299,I153302,I153311,I153317,I153305,I153320,I153302,I153299,I153323,I153369,I153372,I153375,I153378,I153381,I153384,I153387,I153390,I153393,I2224,I2231);
PAT_15 I_2140 (I153381,I153375,I153372,I153390,I153387,I153378,I153369,I153372,I153369,I153384,I153393,I153439,I153442,I153445,I153448,I153451,I153454,I153457,I153460,I153463,I2224,I2231);
PAT_6 I_2141 (I153442,I153439,I153445,I153460,I153442,I153463,I153448,I153454,I153451,I153457,I153439,I153509,I153512,I153515,I153518,I153521,I153524,I153527,I153530,I153533,I153536,I2224,I2231);
PAT_10 I_2142 (I153509,I153524,I153527,I153518,I153509,I153533,I153536,I153512,I153521,I153515,I153530,I153582,I153585,I153588,I153591,I153594,I153597,I153600,I153603,I2224,I2231);
PAT_13 I_2143 (I153588,I153594,I153588,I153585,I153600,I153603,I153582,I153582,I153597,I153585,I153591,I153649,I153652,I153655,I153658,I153661,I153664,I153667,I153670,I153673,I2224,I2231);
PAT_2 I_2144 (I153667,I153661,I153658,I153664,I153649,I153673,I153652,I153670,I153649,I153655,I153652,I153719,I153722,I153725,I153728,I153731,I153734,I153737,I153740,I153743,I2224,I2231);
PAT_9 I_2145 (I153734,I153743,I153719,I153725,I153728,I153737,I153722,I153731,I153740,I153722,I153719,I153789,I153792,I153795,I153798,I153801,I153804,I153807,I153810,I153813,I2224,I2231);
PAT_11 I_2146 (I153801,I153807,I153813,I153810,I153798,I153792,I153792,I153789,I153804,I153789,I153795,I153859,I153862,I153865,I153868,I153871,I153874,I153877,I153880,I153883,I153886,I2224,I2231);
PAT_5 I_2147 (I153880,I153859,I153886,I153874,I153871,I153883,I153865,I153859,I153877,I153862,I153868,I153932,I153935,I153938,I153941,I153944,I153947,I153950,I153953,I153956,I153959,I2224,I2231);
PAT_4 I_2148 (I153950,I153956,I153959,I153938,I153941,I153953,I153935,I153932,I153944,I153947,I153932,I154005,I154008,I154011,I154014,I154017,I154020,I154023,I154026,I154029,I2224,I2231);
PAT_6 I_2149 (I154005,I154011,I154008,I154020,I154023,I154017,I154029,I154026,I154005,I154014,I154008,I154075,I154078,I154081,I154084,I154087,I154090,I154093,I154096,I154099,I154102,I2224,I2231);
PAT_13 I_2150 (I154099,I154081,I154096,I154075,I154078,I154084,I154102,I154087,I154093,I154075,I154090,I154148,I154151,I154154,I154157,I154160,I154163,I154166,I154169,I154172,I2224,I2231);
PAT_2 I_2151 (I154166,I154160,I154157,I154163,I154148,I154172,I154151,I154169,I154148,I154154,I154151,I154218,I154221,I154224,I154227,I154230,I154233,I154236,I154239,I154242,I2224,I2231);
PAT_1 I_2152 (I154230,I154218,I154224,I154227,I154218,I154233,I154242,I154221,I154236,I154221,I154239,I154288,I154291,I154294,I154297,I154300,I154303,I154306,I154309,I154312,I2224,I2231);
PAT_6 I_2153 (I154297,I154288,I154291,I154294,I154309,I154312,I154306,I154288,I154303,I154300,I154291,I154358,I154361,I154364,I154367,I154370,I154373,I154376,I154379,I154382,I154385,I2224,I2231);
PAT_13 I_2154 (I154382,I154364,I154379,I154358,I154361,I154367,I154385,I154370,I154376,I154358,I154373,I154431,I154434,I154437,I154440,I154443,I154446,I154449,I154452,I154455,I2224,I2231);
PAT_8 I_2155 (I154440,I154452,I154443,I154446,I154455,I154434,I154449,I154431,I154434,I154437,I154431,I154501,I154504,I154507,I154510,I154513,I154516,I154519,I154522,I154525,I2224,I2231);
PAT_9 I_2156 (I154504,I154513,I154504,I154501,I154516,I154507,I154522,I154510,I154519,I154501,I154525,I154571,I154574,I154577,I154580,I154583,I154586,I154589,I154592,I154595,I2224,I2231);
PAT_11 I_2157 (I154583,I154589,I154595,I154592,I154580,I154574,I154574,I154571,I154586,I154571,I154577,I154641,I154644,I154647,I154650,I154653,I154656,I154659,I154662,I154665,I154668,I2224,I2231);
PAT_16 I_2158 (I154650,I154656,I154662,I154668,I154653,I154644,I154641,I154641,I154659,I154665,I154647,I154714,I154717,I154720,I154723,I154726,I154729,I154732,I154735,I154738,I154741,I2224,I2231);
PAT_5 I_2159 (I154732,I154735,I154723,I154729,I154720,I154714,I154738,I154741,I154717,I154714,I154726,I154787,I154790,I154793,I154796,I154799,I154802,I154805,I154808,I154811,I154814,I2224,I2231);
PAT_9 I_2160 (I154802,I154799,I154808,I154805,I154796,I154787,I154793,I154814,I154790,I154811,I154787,I154860,I154863,I154866,I154869,I154872,I154875,I154878,I154881,I154884,I2224,I2231);
PAT_10 I_2161 (I154881,I154878,I154866,I154863,I154884,I154869,I154875,I154863,I154860,I154860,I154872,I154930,I154933,I154936,I154939,I154942,I154945,I154948,I154951,I2224,I2231);
PAT_14 I_2162 (I154930,I154951,I154936,I154945,I154942,I154948,I154939,I154933,I154933,I154936,I154930,I154997,I155000,I155003,I155006,I155009,I155012,I155015,I155018,I155021,I2224,I2231);
PAT_6 I_2163 (I154997,I155000,I155021,I155006,I154997,I155003,I155009,I155012,I155015,I155000,I155018,I155067,I155070,I155073,I155076,I155079,I155082,I155085,I155088,I155091,I155094,I2224,I2231);
PAT_5 I_2164 (I155088,I155067,I155073,I155076,I155082,I155085,I155067,I155091,I155070,I155079,I155094,I155140,I155143,I155146,I155149,I155152,I155155,I155158,I155161,I155164,I155167,I2224,I2231);
PAT_2 I_2165 (I155155,I155140,I155152,I155146,I155161,I155143,I155158,I155149,I155164,I155167,I155140,I155213,I155216,I155219,I155222,I155225,I155228,I155231,I155234,I155237,I2224,I2231);
PAT_15 I_2166 (I155216,I155228,I155234,I155237,I155219,I155231,I155213,I155222,I155213,I155225,I155216,I155283,I155286,I155289,I155292,I155295,I155298,I155301,I155304,I155307,I2224,I2231);
PAT_2 I_2167 (I155286,I155286,I155289,I155295,I155283,I155283,I155292,I155307,I155301,I155304,I155298,I155353,I155356,I155359,I155362,I155365,I155368,I155371,I155374,I155377,I2224,I2231);
PAT_8 I_2168 (I155365,I155356,I155362,I155353,I155359,I155374,I155371,I155353,I155368,I155356,I155377,I155423,I155426,I155429,I155432,I155435,I155438,I155441,I155444,I155447,I2224,I2231);
PAT_10 I_2169 (I155429,I155423,I155426,I155447,I155441,I155426,I155435,I155423,I155444,I155438,I155432,I155493,I155496,I155499,I155502,I155505,I155508,I155511,I155514,I2224,I2231);
PAT_13 I_2170 (I155499,I155505,I155499,I155496,I155511,I155514,I155493,I155493,I155508,I155496,I155502,I155560,I155563,I155566,I155569,I155572,I155575,I155578,I155581,I155584,I2224,I2231);
PAT_11 I_2171 (I155560,I155572,I155575,I155566,I155563,I155584,I155563,I155581,I155569,I155560,I155578,I155630,I155633,I155636,I155639,I155642,I155645,I155648,I155651,I155654,I155657,I2224,I2231);
PAT_5 I_2172 (I155651,I155630,I155657,I155645,I155642,I155654,I155636,I155630,I155648,I155633,I155639,I155703,I155706,I155709,I155712,I155715,I155718,I155721,I155724,I155727,I155730,I2224,I2231);
PAT_9 I_2173 (I155718,I155715,I155724,I155721,I155712,I155703,I155709,I155730,I155706,I155727,I155703,I155776,I155779,I155782,I155785,I155788,I155791,I155794,I155797,I155800,I2224,I2231);
PAT_4 I_2174 (I155776,I155800,I155794,I155782,I155779,I155797,I155779,I155776,I155791,I155785,I155788,I155846,I155849,I155852,I155855,I155858,I155861,I155864,I155867,I155870,I2224,I2231);
PAT_13 I_2175 (I155861,I155855,I155867,I155852,I155858,I155846,I155870,I155864,I155849,I155846,I155849,I155916,I155919,I155922,I155925,I155928,I155931,I155934,I155937,I155940,I2224,I2231);
PAT_8 I_2176 (I155925,I155937,I155928,I155931,I155940,I155919,I155934,I155916,I155919,I155922,I155916,I155986,I155989,I155992,I155995,I155998,I156001,I156004,I156007,I156010,I2224,I2231);
PAT_5 I_2177 (I155992,I156010,I155986,I156007,I155995,I155998,I155989,I155986,I155989,I156001,I156004,I156056,I156059,I156062,I156065,I156068,I156071,I156074,I156077,I156080,I156083,I2224,I2231);
PAT_4 I_2178 (I156074,I156080,I156083,I156062,I156065,I156077,I156059,I156056,I156068,I156071,I156056,I156129,I156132,I156135,I156138,I156141,I156144,I156147,I156150,I156153,I2224,I2231);
PAT_6 I_2179 (I156129,I156135,I156132,I156144,I156147,I156141,I156153,I156150,I156129,I156138,I156132,I156199,I156202,I156205,I156208,I156211,I156214,I156217,I156220,I156223,I156226,I2224,I2231);
PAT_2 I_2180 (I156220,I156226,I156208,I156214,I156199,I156205,I156199,I156211,I156202,I156217,I156223,I156272,I156275,I156278,I156281,I156284,I156287,I156290,I156293,I156296,I2224,I2231);
PAT_1 I_2181 (I156284,I156272,I156278,I156281,I156272,I156287,I156296,I156275,I156290,I156275,I156293,I156342,I156345,I156348,I156351,I156354,I156357,I156360,I156363,I156366,I2224,I2231);
PAT_9 I_2182 (I156357,I156363,I156348,I156366,I156345,I156360,I156345,I156351,I156342,I156354,I156342,I156412,I156415,I156418,I156421,I156424,I156427,I156430,I156433,I156436,I2224,I2231);
PAT_14 I_2183 (I156421,I156412,I156436,I156418,I156415,I156412,I156427,I156433,I156424,I156415,I156430,I156482,I156485,I156488,I156491,I156494,I156497,I156500,I156503,I156506,I2224,I2231);
PAT_17 I_2184 (I156497,I156485,I156506,I156482,I156503,I156491,I156488,I156500,I156494,I156485,I156482,I156552,I156555,I156558,I156561,I156564,I156567,I156570,I156573,I156576,I156579,I2224,I2231);
PAT_1 I_2185 (I156576,I156579,I156558,I156567,I156552,I156573,I156564,I156555,I156561,I156552,I156570,I156625,I156628,I156631,I156634,I156637,I156640,I156643,I156646,I156649,I2224,I2231);
PAT_12 I_2186 (I156637,I156631,I156649,I156625,I156634,I156625,I156628,I156646,I156640,I156628,I156643,I156695,I156698,I156701,I156704,I156707,I156710,I156713,I156716,I2224,I2231);
PAT_7 I_2187 (I156701,I156704,I156695,I156707,I156713,I156701,I156716,I156710,I156698,I156698,I156695,I156762,I156765,I156768,I156771,I156774,I156777,I156780,I156783,I156786,I2224,I2231);
PAT_9 I_2188 (I156783,I156771,I156780,I156786,I156768,I156774,I156765,I156777,I156762,I156762,I156765,I156832,I156835,I156838,I156841,I156844,I156847,I156850,I156853,I156856,I2224,I2231);
PAT_11 I_2189 (I156844,I156850,I156856,I156853,I156841,I156835,I156835,I156832,I156847,I156832,I156838,I156902,I156905,I156908,I156911,I156914,I156917,I156920,I156923,I156926,I156929,I2224,I2231);
PAT_5 I_2190 (I156923,I156902,I156929,I156917,I156914,I156926,I156908,I156902,I156920,I156905,I156911,I156975,I156978,I156981,I156984,I156987,I156990,I156993,I156996,I156999,I157002,I2224,I2231);
PAT_7 I_2191 (I156993,I156996,I157002,I156999,I156984,I156981,I156975,I156987,I156975,I156978,I156990,I157048,I157051,I157054,I157057,I157060,I157063,I157066,I157069,I157072,I2224,I2231);
PAT_4 I_2192 (I157072,I157048,I157048,I157063,I157057,I157051,I157051,I157066,I157069,I157054,I157060,I157118,I157121,I157124,I157127,I157130,I157133,I157136,I157139,I157142,I2224,I2231);
PAT_9 I_2193 (I157139,I157121,I157124,I157133,I157136,I157118,I157127,I157121,I157142,I157118,I157130,I157188,I157191,I157194,I157197,I157200,I157203,I157206,I157209,I157212,I2224,I2231);
PAT_5 I_2194 (I157209,I157188,I157203,I157188,I157194,I157197,I157191,I157191,I157206,I157200,I157212,I157258,I157261,I157264,I157267,I157270,I157273,I157276,I157279,I157282,I157285,I2224,I2231);
PAT_11 I_2195 (I157270,I157267,I157261,I157279,I157282,I157258,I157276,I157273,I157285,I157264,I157258,I157331,I157334,I157337,I157340,I157343,I157346,I157349,I157352,I157355,I157358,I2224,I2231);
PAT_2 I_2196 (I157331,I157355,I157343,I157337,I157346,I157349,I157334,I157358,I157352,I157340,I157331,I157404,I157407,I157410,I157413,I157416,I157419,I157422,I157425,I157428,I2224,I2231);
PAT_10 I_2197 (I157404,I157422,I157419,I157407,I157410,I157425,I157416,I157404,I157413,I157428,I157407,I157474,I157477,I157480,I157483,I157486,I157489,I157492,I157495,I2224,I2231);
PAT_11 I_2198 (I157483,I157486,I157495,I157489,I157492,I157474,I157474,I157480,I157477,I157477,I157480,I157541,I157544,I157547,I157550,I157553,I157556,I157559,I157562,I157565,I157568,I2224,I2231);
PAT_8 I_2199 (I157550,I157556,I157559,I157565,I157562,I157553,I157541,I157541,I157568,I157544,I157547,I157614,I157617,I157620,I157623,I157626,I157629,I157632,I157635,I157638,I2224,I2231);
PAT_11 I_2200 (I157635,I157626,I157614,I157617,I157632,I157620,I157623,I157614,I157638,I157629,I157617,I157684,I157687,I157690,I157693,I157696,I157699,I157702,I157705,I157708,I157711,I2224,I2231);
PAT_6 I_2201 (I157684,I157711,I157699,I157708,I157702,I157696,I157687,I157705,I157693,I157690,I157684,I157757,I157760,I157763,I157766,I157769,I157772,I157775,I157778,I157781,I157784,I2224,I2231);
PAT_5 I_2202 (I157778,I157757,I157763,I157766,I157772,I157775,I157757,I157781,I157760,I157769,I157784,I157830,I157833,I157836,I157839,I157842,I157845,I157848,I157851,I157854,I157857,I2224,I2231);
PAT_15 I_2203 (I157848,I157833,I157830,I157830,I157845,I157842,I157854,I157839,I157851,I157836,I157857,I157903,I157906,I157909,I157912,I157915,I157918,I157921,I157924,I157927,I2224,I2231);
PAT_11 I_2204 (I157924,I157906,I157903,I157918,I157909,I157903,I157921,I157927,I157915,I157906,I157912,I157973,I157976,I157979,I157982,I157985,I157988,I157991,I157994,I157997,I158000,I2224,I2231);
PAT_10 I_2205 (I157988,I157994,I157985,I157979,I157997,I157982,I158000,I157991,I157973,I157976,I157973,I158046,I158049,I158052,I158055,I158058,I158061,I158064,I158067,I2224,I2231);
PAT_9 I_2206 (I158058,I158046,I158049,I158052,I158046,I158052,I158055,I158049,I158067,I158061,I158064,I158113,I158116,I158119,I158122,I158125,I158128,I158131,I158134,I158137,I2224,I2231);
PAT_17 I_2207 (I158116,I158122,I158137,I158128,I158131,I158119,I158113,I158125,I158113,I158116,I158134,I158183,I158186,I158189,I158192,I158195,I158198,I158201,I158204,I158207,I158210,I2224,I2231);
PAT_9 I_2208 (I158204,I158186,I158192,I158207,I158189,I158201,I158183,I158195,I158183,I158210,I158198,I158256,I158259,I158262,I158265,I158268,I158271,I158274,I158277,I158280,I2224,I2231);
PAT_13 I_2209 (I158256,I158277,I158259,I158274,I158268,I158265,I158280,I158256,I158262,I158271,I158259,I158326,I158329,I158332,I158335,I158338,I158341,I158344,I158347,I158350,I2224,I2231);
PAT_9 I_2210 (I158347,I158329,I158329,I158326,I158350,I158332,I158335,I158326,I158338,I158344,I158341,I158396,I158399,I158402,I158405,I158408,I158411,I158414,I158417,I158420,I2224,I2231);
PAT_4 I_2211 (I158396,I158420,I158414,I158402,I158399,I158417,I158399,I158396,I158411,I158405,I158408,I158466,I158469,I158472,I158475,I158478,I158481,I158484,I158487,I158490,I2224,I2231);
PAT_12 I_2212 (I158466,I158469,I158487,I158490,I158481,I158472,I158478,I158475,I158466,I158484,I158469,I158536,I158539,I158542,I158545,I158548,I158551,I158554,I158557,I2224,I2231);
PAT_10 I_2213 (I158536,I158557,I158548,I158551,I158542,I158539,I158536,I158554,I158542,I158545,I158539,I158603,I158606,I158609,I158612,I158615,I158618,I158621,I158624,I2224,I2231);
PAT_11 I_2214 (I158612,I158615,I158624,I158618,I158621,I158603,I158603,I158609,I158606,I158606,I158609,I158670,I158673,I158676,I158679,I158682,I158685,I158688,I158691,I158694,I158697,I2224,I2231);
PAT_13 I_2215 (I158670,I158673,I158682,I158694,I158697,I158685,I158691,I158679,I158688,I158676,I158670,I158743,I158746,I158749,I158752,I158755,I158758,I158761,I158764,I158767,I2224,I2231);
PAT_6 I_2216 (I158743,I158755,I158752,I158764,I158761,I158767,I158743,I158758,I158746,I158746,I158749,I158813,I158816,I158819,I158822,I158825,I158828,I158831,I158834,I158837,I158840,I2224,I2231);
PAT_12 I_2217 (I158813,I158840,I158819,I158822,I158816,I158813,I158834,I158828,I158831,I158825,I158837,I158886,I158889,I158892,I158895,I158898,I158901,I158904,I158907,I2224,I2231);
PAT_6 I_2218 (I158895,I158889,I158907,I158892,I158889,I158892,I158901,I158886,I158904,I158886,I158898,I158953,I158956,I158959,I158962,I158965,I158968,I158971,I158974,I158977,I158980,I2224,I2231);
PAT_9 I_2219 (I158953,I158980,I158977,I158959,I158965,I158956,I158968,I158953,I158971,I158962,I158974,I159026,I159029,I159032,I159035,I159038,I159041,I159044,I159047,I159050,I2224,I2231);
PAT_17 I_2220 (I159029,I159035,I159050,I159041,I159044,I159032,I159026,I159038,I159026,I159029,I159047,I159096,I159099,I159102,I159105,I159108,I159111,I159114,I159117,I159120,I159123,I2224,I2231);
PAT_8 I_2221 (I159105,I159117,I159123,I159114,I159099,I159108,I159111,I159120,I159102,I159096,I159096,I159169,I159172,I159175,I159178,I159181,I159184,I159187,I159190,I159193,I2224,I2231);
PAT_11 I_2222 (I159190,I159181,I159169,I159172,I159187,I159175,I159178,I159169,I159193,I159184,I159172,I159239,I159242,I159245,I159248,I159251,I159254,I159257,I159260,I159263,I159266,I2224,I2231);
PAT_9 I_2223 (I159245,I159257,I159248,I159260,I159239,I159242,I159251,I159239,I159254,I159263,I159266,I159312,I159315,I159318,I159321,I159324,I159327,I159330,I159333,I159336,I2224,I2231);
PAT_10 I_2224 (I159333,I159330,I159318,I159315,I159336,I159321,I159327,I159315,I159312,I159312,I159324,I159382,I159385,I159388,I159391,I159394,I159397,I159400,I159403,I2224,I2231);
PAT_9 I_2225 (I159394,I159382,I159385,I159388,I159382,I159388,I159391,I159385,I159403,I159397,I159400,I159449,I159452,I159455,I159458,I159461,I159464,I159467,I159470,I159473,I2224,I2231);
PAT_12 I_2226 (I159470,I159467,I159461,I159449,I159458,I159449,I159452,I159455,I159473,I159464,I159452,I159519,I159522,I159525,I159528,I159531,I159534,I159537,I159540,I2224,I2231);
PAT_9 I_2227 (I159528,I159534,I159519,I159525,I159531,I159522,I159519,I159522,I159540,I159525,I159537,I159586,I159589,I159592,I159595,I159598,I159601,I159604,I159607,I159610,I2224,I2231);
PAT_2 I_2228 (I159601,I159604,I159595,I159610,I159586,I159589,I159592,I159589,I159607,I159598,I159586,I159656,I159659,I159662,I159665,I159668,I159671,I159674,I159677,I159680,I2224,I2231);
PAT_4 I_2229 (I159656,I159662,I159680,I159674,I159671,I159668,I159659,I159677,I159656,I159659,I159665,I159726,I159729,I159732,I159735,I159738,I159741,I159744,I159747,I159750,I2224,I2231);
PAT_5 I_2230 (I159747,I159729,I159729,I159741,I159744,I159738,I159735,I159726,I159732,I159726,I159750,I159796,I159799,I159802,I159805,I159808,I159811,I159814,I159817,I159820,I159823,I2224,I2231);
PAT_11 I_2231 (I159808,I159805,I159799,I159817,I159820,I159796,I159814,I159811,I159823,I159802,I159796,I159869,I159872,I159875,I159878,I159881,I159884,I159887,I159890,I159893,I159896,I2224,I2231);
PAT_17 I_2232 (I1713,I1657,I1673,I1505,I1417,I1433,I1481,I1633,I1841,I2097,I1857,I159942,I159945,I159948,I159951,I159954,I159957,I159960,I159963,I159966,I159969,I2224,I2231);
PAT_13 I_2233 (I159960,I159963,I159948,I159942,I159954,I159966,I159945,I159957,I159942,I159969,I159951,I160015,I160018,I160021,I160024,I160027,I160030,I160033,I160036,I160039,I2224,I2231);
PAT_12 I_2234 (I160024,I160015,I160015,I160039,I160036,I160018,I160033,I160027,I160018,I160021,I160030,I160085,I160088,I160091,I160094,I160097,I160100,I160103,I160106,I2224,I2231);
PAT_7 I_2235 (I160091,I160094,I160085,I160097,I160103,I160091,I160106,I160100,I160088,I160088,I160085,I160152,I160155,I160158,I160161,I160164,I160167,I160170,I160173,I160176,I2224,I2231);
PAT_3 I_2236 (I160173,I160161,I160152,I160158,I160167,I160155,I160176,I160152,I160170,I160164,I160155,I160222,I160225,I160228,I160231,I160234,I160237,I160240,I160243,I160246,I160249,I2224,I2231);
PAT_12 I_2237 (I160237,I160243,I160222,I160249,I160240,I160231,I160234,I160225,I160222,I160228,I160246,I160295,I160298,I160301,I160304,I160307,I160310,I160313,I160316,I2224,I2231);
PAT_9 I_2238 (I160304,I160310,I160295,I160301,I160307,I160298,I160295,I160298,I160316,I160301,I160313,I160362,I160365,I160368,I160371,I160374,I160377,I160380,I160383,I160386,I2224,I2231);
PAT_17 I_2239 (I160365,I160371,I160386,I160377,I160380,I160368,I160362,I160374,I160362,I160365,I160383,I160432,I160435,I160438,I160441,I160444,I160447,I160450,I160453,I160456,I160459,I2224,I2231);
PAT_10 I_2240 (I160432,I160438,I160459,I160441,I160456,I160435,I160450,I160444,I160453,I160447,I160432,I160505,I160508,I160511,I160514,I160517,I160520,I160523,I160526,I2224,I2231);
PAT_4 I_2241 (I160520,I160517,I160508,I160526,I160505,I160508,I160514,I160511,I160523,I160505,I160511,I160572,I160575,I160578,I160581,I160584,I160587,I160590,I160593,I160596,I2224,I2231);
PAT_6 I_2242 (I160572,I160578,I160575,I160587,I160590,I160584,I160596,I160593,I160572,I160581,I160575,I160642,I160645,I160648,I160651,I160654,I160657,I160660,I160663,I160666,I160669,I2224,I2231);
PAT_8 I_2243 (I160651,I160657,I160648,I160660,I160642,I160645,I160663,I160642,I160669,I160666,I160654,I160715,I160718,I160721,I160724,I160727,I160730,I160733,I160736,I160739,I2224,I2231);
PAT_4 I_2244 (I160733,I160718,I160724,I160715,I160715,I160727,I160718,I160736,I160739,I160721,I160730,I160785,I160788,I160791,I160794,I160797,I160800,I160803,I160806,I160809,I2224,I2231);
PAT_9 I_2245 (I160806,I160788,I160791,I160800,I160803,I160785,I160794,I160788,I160809,I160785,I160797,I160855,I160858,I160861,I160864,I160867,I160870,I160873,I160876,I160879,I2224,I2231);
PAT_17 I_2246 (I160858,I160864,I160879,I160870,I160873,I160861,I160855,I160867,I160855,I160858,I160876,I160925,I160928,I160931,I160934,I160937,I160940,I160943,I160946,I160949,I160952,I2224,I2231);
PAT_6 I_2247 (I160925,I160943,I160931,I160934,I160940,I160925,I160937,I160928,I160949,I160952,I160946,I160998,I161001,I161004,I161007,I161010,I161013,I161016,I161019,I161022,I161025,I2224,I2231);
PAT_9 I_2248 (I160998,I161025,I161022,I161004,I161010,I161001,I161013,I160998,I161016,I161007,I161019,I161071,I161074,I161077,I161080,I161083,I161086,I161089,I161092,I161095,I2224,I2231);
PAT_11 I_2249 (I161083,I161089,I161095,I161092,I161080,I161074,I161074,I161071,I161086,I161071,I161077,I161141,I161144,I161147,I161150,I161153,I161156,I161159,I161162,I161165,I161168,I2224,I2231);
PAT_15 I_2250 (I161165,I161144,I161150,I161159,I161156,I161141,I161153,I161162,I161141,I161147,I161168,I161214,I161217,I161220,I161223,I161226,I161229,I161232,I161235,I161238,I2224,I2231);
PAT_8 I_2251 (I161235,I161214,I161214,I161223,I161220,I161217,I161232,I161229,I161217,I161238,I161226,I161284,I161287,I161290,I161293,I161296,I161299,I161302,I161305,I161308,I2224,I2231);
PAT_4 I_2252 (I161302,I161287,I161293,I161284,I161284,I161296,I161287,I161305,I161308,I161290,I161299,I161354,I161357,I161360,I161363,I161366,I161369,I161372,I161375,I161378,I2224,I2231);
PAT_15 I_2253 (I161354,I161357,I161378,I161363,I161372,I161375,I161360,I161369,I161366,I161354,I161357,I161424,I161427,I161430,I161433,I161436,I161439,I161442,I161445,I161448,I2224,I2231);
PAT_17 I_2254 (I161424,I161424,I161436,I161427,I161430,I161448,I161445,I161439,I161427,I161433,I161442,I161494,I161497,I161500,I161503,I161506,I161509,I161512,I161515,I161518,I161521,I2224,I2231);
PAT_4 I_2255 (I161503,I161494,I161512,I161509,I161521,I161518,I161497,I161494,I161500,I161506,I161515,I161567,I161570,I161573,I161576,I161579,I161582,I161585,I161588,I161591,I2224,I2231);
PAT_7 I_2256 (I161582,I161576,I161573,I161567,I161579,I161585,I161570,I161570,I161588,I161591,I161567,I161637,I161640,I161643,I161646,I161649,I161652,I161655,I161658,I161661,I2224,I2231);
PAT_9 I_2257 (I161658,I161646,I161655,I161661,I161643,I161649,I161640,I161652,I161637,I161637,I161640,I161707,I161710,I161713,I161716,I161719,I161722,I161725,I161728,I161731,I2224,I2231);
PAT_10 I_2258 (I161728,I161725,I161713,I161710,I161731,I161716,I161722,I161710,I161707,I161707,I161719,I161777,I161780,I161783,I161786,I161789,I161792,I161795,I161798,I2224,I2231);
PAT_13 I_2259 (I161783,I161789,I161783,I161780,I161795,I161798,I161777,I161777,I161792,I161780,I161786,I161844,I161847,I161850,I161853,I161856,I161859,I161862,I161865,I161868,I2224,I2231);
PAT_15 I_2260 (I161844,I161856,I161847,I161859,I161844,I161853,I161868,I161865,I161850,I161862,I161847,I161914,I161917,I161920,I161923,I161926,I161929,I161932,I161935,I161938,I2224,I2231);
PAT_3 I_2261 (I161935,I161923,I161914,I161917,I161920,I161929,I161926,I161932,I161914,I161917,I161938,I161984,I161987,I161990,I161993,I161996,I161999,I162002,I162005,I162008,I162011,I2224,I2231);
PAT_2 I_2262 (I162011,I161996,I161987,I161984,I162008,I161999,I161993,I162002,I161984,I162005,I161990,I162057,I162060,I162063,I162066,I162069,I162072,I162075,I162078,I162081,I2224,I2231);
PAT_4 I_2263 (I162057,I162063,I162081,I162075,I162072,I162069,I162060,I162078,I162057,I162060,I162066,I162127,I162130,I162133,I162136,I162139,I162142,I162145,I162148,I162151,I2224,I2231);
PAT_2 I_2264 (I162136,I162130,I162130,I162151,I162127,I162145,I162142,I162133,I162127,I162139,I162148,I162197,I162200,I162203,I162206,I162209,I162212,I162215,I162218,I162221,I2224,I2231);
PAT_13 I_2265 (I162206,I162200,I162197,I162218,I162209,I162212,I162200,I162203,I162215,I162221,I162197,I162267,I162270,I162273,I162276,I162279,I162282,I162285,I162288,I162291,I2224,I2231);
PAT_10 I_2266 (I162288,I162282,I162276,I162270,I162291,I162270,I162279,I162267,I162267,I162285,I162273,I162337,I162340,I162343,I162346,I162349,I162352,I162355,I162358,I2224,I2231);
PAT_6 I_2267 (I162358,I162352,I162346,I162340,I162337,I162343,I162337,I162343,I162340,I162349,I162355,I162404,I162407,I162410,I162413,I162416,I162419,I162422,I162425,I162428,I162431,I2224,I2231);
PAT_13 I_2268 (I162428,I162410,I162425,I162404,I162407,I162413,I162431,I162416,I162422,I162404,I162419,I162477,I162480,I162483,I162486,I162489,I162492,I162495,I162498,I162501,I2224,I2231);
PAT_9 I_2269 (I162498,I162480,I162480,I162477,I162501,I162483,I162486,I162477,I162489,I162495,I162492,I162547,I162550,I162553,I162556,I162559,I162562,I162565,I162568,I162571,I2224,I2231);
PAT_17 I_2270 (I162550,I162556,I162571,I162562,I162565,I162553,I162547,I162559,I162547,I162550,I162568,I162617,I162620,I162623,I162626,I162629,I162632,I162635,I162638,I162641,I162644,I2224,I2231);
PAT_8 I_2271 (I162626,I162638,I162644,I162635,I162620,I162629,I162632,I162641,I162623,I162617,I162617,I162690,I162693,I162696,I162699,I162702,I162705,I162708,I162711,I162714,I2224,I2231);
PAT_4 I_2272 (I162708,I162693,I162699,I162690,I162690,I162702,I162693,I162711,I162714,I162696,I162705,I162760,I162763,I162766,I162769,I162772,I162775,I162778,I162781,I162784,I2224,I2231);
PAT_13 I_2273 (I162775,I162769,I162781,I162766,I162772,I162760,I162784,I162778,I162763,I162760,I162763,I162830,I162833,I162836,I162839,I162842,I162845,I162848,I162851,I162854,I2224,I2231);
PAT_6 I_2274 (I162830,I162842,I162839,I162851,I162848,I162854,I162830,I162845,I162833,I162833,I162836,I162900,I162903,I162906,I162909,I162912,I162915,I162918,I162921,I162924,I162927,I2224,I2231);
PAT_9 I_2275 (I162900,I162927,I162924,I162906,I162912,I162903,I162915,I162900,I162918,I162909,I162921,I162973,I162976,I162979,I162982,I162985,I162988,I162991,I162994,I162997,I2224,I2231);
PAT_11 I_2276 (I162985,I162991,I162997,I162994,I162982,I162976,I162976,I162973,I162988,I162973,I162979,I163043,I163046,I163049,I163052,I163055,I163058,I163061,I163064,I163067,I163070,I2224,I2231);
PAT_9 I_2277 (I163049,I163061,I163052,I163064,I163043,I163046,I163055,I163043,I163058,I163067,I163070,I163116,I163119,I163122,I163125,I163128,I163131,I163134,I163137,I163140,I2224,I2231);
PAT_11 I_2278 (I163128,I163134,I163140,I163137,I163125,I163119,I163119,I163116,I163131,I163116,I163122,I163186,I163189,I163192,I163195,I163198,I163201,I163204,I163207,I163210,I163213,I2224,I2231);
PAT_17 I_2279 (I163198,I163189,I163213,I163186,I163195,I163207,I163204,I163201,I163186,I163210,I163192,I163259,I163262,I163265,I163268,I163271,I163274,I163277,I163280,I163283,I163286,I2224,I2231);
PAT_6 I_2280 (I163259,I163277,I163265,I163268,I163274,I163259,I163271,I163262,I163283,I163286,I163280,I163332,I163335,I163338,I163341,I163344,I163347,I163350,I163353,I163356,I163359,I2224,I2231);
PAT_9 I_2281 (I163332,I163359,I163356,I163338,I163344,I163335,I163347,I163332,I163350,I163341,I163353,I163405,I163408,I163411,I163414,I163417,I163420,I163423,I163426,I163429,I2224,I2231);
PAT_0 I_2282 (I163414,I163426,I163405,I163408,I163411,I163405,I163420,I163423,I163417,I163429,I163408,I163475,I163478,I163481,I163484,I163487,I163490,I163493,I163496,I2224,I2231);
PAT_1 I_2283 (I163478,I163475,I163475,I163493,I163478,I163487,I163481,I163490,I163484,I163496,I163481,I163542,I163545,I163548,I163551,I163554,I163557,I163560,I163563,I163566,I2224,I2231);
PAT_10 I_2284 (I163557,I163554,I163545,I163542,I163545,I163560,I163548,I163563,I163566,I163551,I163542,I163612,I163615,I163618,I163621,I163624,I163627,I163630,I163633,I2224,I2231);
PAT_2 I_2285 (I163624,I163627,I163618,I163630,I163615,I163612,I163612,I163618,I163633,I163621,I163615,I163679,I163682,I163685,I163688,I163691,I163694,I163697,I163700,I163703,I2224,I2231);
PAT_10 I_2286 (I163679,I163697,I163694,I163682,I163685,I163700,I163691,I163679,I163688,I163703,I163682,I163749,I163752,I163755,I163758,I163761,I163764,I163767,I163770,I2224,I2231);
PAT_5 I_2287 (I163770,I163749,I163758,I163752,I163767,I163764,I163755,I163755,I163749,I163752,I163761,I163816,I163819,I163822,I163825,I163828,I163831,I163834,I163837,I163840,I163843,I2224,I2231);
PAT_6 I_2288 (I163834,I163828,I163816,I163822,I163819,I163825,I163831,I163816,I163840,I163837,I163843,I163889,I163892,I163895,I163898,I163901,I163904,I163907,I163910,I163913,I163916,I2224,I2231);
PAT_10 I_2289 (I163889,I163904,I163907,I163898,I163889,I163913,I163916,I163892,I163901,I163895,I163910,I163962,I163965,I163968,I163971,I163974,I163977,I163980,I163983,I2224,I2231);
PAT_4 I_2290 (I163977,I163974,I163965,I163983,I163962,I163965,I163971,I163968,I163980,I163962,I163968,I164029,I164032,I164035,I164038,I164041,I164044,I164047,I164050,I164053,I2224,I2231);
PAT_11 I_2291 (I164041,I164050,I164032,I164044,I164029,I164032,I164029,I164038,I164053,I164047,I164035,I164099,I164102,I164105,I164108,I164111,I164114,I164117,I164120,I164123,I164126,I2224,I2231);
PAT_4 I_2292 (I164105,I164126,I164099,I164117,I164108,I164099,I164120,I164102,I164111,I164123,I164114,I164172,I164175,I164178,I164181,I164184,I164187,I164190,I164193,I164196,I2224,I2231);
PAT_0 I_2293 (I164178,I164196,I164172,I164172,I164187,I164193,I164184,I164190,I164181,I164175,I164175,I164242,I164245,I164248,I164251,I164254,I164257,I164260,I164263,I2224,I2231);
PAT_13 I_2294 (I164251,I164260,I164242,I164245,I164245,I164248,I164254,I164248,I164242,I164257,I164263,I164309,I164312,I164315,I164318,I164321,I164324,I164327,I164330,I164333,I2224,I2231);
PAT_10 I_2295 (I164330,I164324,I164318,I164312,I164333,I164312,I164321,I164309,I164309,I164327,I164315,I164379,I164382,I164385,I164388,I164391,I164394,I164397,I164400,I2224,I2231);
PAT_13 I_2296 (I164385,I164391,I164385,I164382,I164397,I164400,I164379,I164379,I164394,I164382,I164388,I164446,I164449,I164452,I164455,I164458,I164461,I164464,I164467,I164470,I2224,I2231);
PAT_4 I_2297 (I164455,I164458,I164470,I164452,I164467,I164464,I164449,I164461,I164449,I164446,I164446,I164516,I164519,I164522,I164525,I164528,I164531,I164534,I164537,I164540,I2224,I2231);
PAT_17 I_2298 (I164528,I164525,I164537,I164531,I164516,I164534,I164540,I164519,I164522,I164519,I164516,I164586,I164589,I164592,I164595,I164598,I164601,I164604,I164607,I164610,I164613,I2224,I2231);
PAT_10 I_2299 (I164586,I164592,I164613,I164595,I164610,I164589,I164604,I164598,I164607,I164601,I164586,I164659,I164662,I164665,I164668,I164671,I164674,I164677,I164680,I2224,I2231);
PAT_7 I_2300 (I164680,I164677,I164674,I164659,I164662,I164665,I164662,I164671,I164659,I164665,I164668,I164726,I164729,I164732,I164735,I164738,I164741,I164744,I164747,I164750,I2224,I2231);
PAT_13 I_2301 (I164732,I164750,I164741,I164726,I164738,I164726,I164747,I164729,I164735,I164729,I164744,I164796,I164799,I164802,I164805,I164808,I164811,I164814,I164817,I164820,I2224,I2231);
PAT_12 I_2302 (I164805,I164796,I164796,I164820,I164817,I164799,I164814,I164808,I164799,I164802,I164811,I164866,I164869,I164872,I164875,I164878,I164881,I164884,I164887,I2224,I2231);
PAT_11 I_2303 (I164872,I164875,I164872,I164884,I164887,I164881,I164869,I164878,I164866,I164869,I164866,I164933,I164936,I164939,I164942,I164945,I164948,I164951,I164954,I164957,I164960,I2224,I2231);
PAT_9 I_2304 (I164939,I164951,I164942,I164954,I164933,I164936,I164945,I164933,I164948,I164957,I164960,I165006,I165009,I165012,I165015,I165018,I165021,I165024,I165027,I165030,I2224,I2231);
PAT_5 I_2305 (I165027,I165006,I165021,I165006,I165012,I165015,I165009,I165009,I165024,I165018,I165030,I165076,I165079,I165082,I165085,I165088,I165091,I165094,I165097,I165100,I165103,I2224,I2231);
PAT_0 I_2306 (I165097,I165076,I165103,I165100,I165076,I165094,I165088,I165079,I165085,I165091,I165082,I165149,I165152,I165155,I165158,I165161,I165164,I165167,I165170,I2224,I2231);
PAT_9 I_2307 (I165155,I165167,I165152,I165161,I165164,I165152,I165149,I165158,I165170,I165155,I165149,I165216,I165219,I165222,I165225,I165228,I165231,I165234,I165237,I165240,I2224,I2231);
PAT_17 I_2308 (I165219,I165225,I165240,I165231,I165234,I165222,I165216,I165228,I165216,I165219,I165237,I165286,I165289,I165292,I165295,I165298,I165301,I165304,I165307,I165310,I165313,I2224,I2231);
PAT_5 I_2309 (I165298,I165292,I165289,I165310,I165295,I165301,I165304,I165286,I165286,I165307,I165313,I165359,I165362,I165365,I165368,I165371,I165374,I165377,I165380,I165383,I165386,I2224,I2231);
PAT_6 I_2310 (I165377,I165371,I165359,I165365,I165362,I165368,I165374,I165359,I165383,I165380,I165386,I165432,I165435,I165438,I165441,I165444,I165447,I165450,I165453,I165456,I165459,I2224,I2231);
PAT_9 I_2311 (I165432,I165459,I165456,I165438,I165444,I165435,I165447,I165432,I165450,I165441,I165453,I165505,I165508,I165511,I165514,I165517,I165520,I165523,I165526,I165529,I2224,I2231);
PAT_2 I_2312 (I165520,I165523,I165514,I165529,I165505,I165508,I165511,I165508,I165526,I165517,I165505,I165575,I165578,I165581,I165584,I165587,I165590,I165593,I165596,I165599,I2224,I2231);
PAT_11 I_2313 (I165578,I165590,I165575,I165587,I165584,I165596,I165593,I165578,I165599,I165581,I165575,I165645,I165648,I165651,I165654,I165657,I165660,I165663,I165666,I165669,I165672,I2224,I2231);
PAT_13 I_2314 (I165645,I165648,I165657,I165669,I165672,I165660,I165666,I165654,I165663,I165651,I165645,I165718,I165721,I165724,I165727,I165730,I165733,I165736,I165739,I165742,I2224,I2231);
PAT_4 I_2315 (I165727,I165730,I165742,I165724,I165739,I165736,I165721,I165733,I165721,I165718,I165718,I165788,I165791,I165794,I165797,I165800,I165803,I165806,I165809,I165812,I2224,I2231);
PAT_12 I_2316 (I165788,I165791,I165809,I165812,I165803,I165794,I165800,I165797,I165788,I165806,I165791,I165858,I165861,I165864,I165867,I165870,I165873,I165876,I165879,I2224,I2231);
PAT_17 I_2317 (I165873,I165867,I165861,I165858,I165858,I165864,I165864,I165876,I165879,I165861,I165870,I165925,I165928,I165931,I165934,I165937,I165940,I165943,I165946,I165949,I165952,I2224,I2231);
PAT_5 I_2318 (I165937,I165931,I165928,I165949,I165934,I165940,I165943,I165925,I165925,I165946,I165952,I165998,I166001,I166004,I166007,I166010,I166013,I166016,I166019,I166022,I166025,I2224,I2231);
PAT_9 I_2319 (I166013,I166010,I166019,I166016,I166007,I165998,I166004,I166025,I166001,I166022,I165998,I166071,I166074,I166077,I166080,I166083,I166086,I166089,I166092,I166095,I2224,I2231);
PAT_13 I_2320 (I166071,I166092,I166074,I166089,I166083,I166080,I166095,I166071,I166077,I166086,I166074,I166141,I166144,I166147,I166150,I166153,I166156,I166159,I166162,I166165,I2224,I2231);
PAT_4 I_2321 (I166150,I166153,I166165,I166147,I166162,I166159,I166144,I166156,I166144,I166141,I166141,I166211,I166214,I166217,I166220,I166223,I166226,I166229,I166232,I166235,I2224,I2231);
PAT_8 I_2322 (I166223,I166211,I166232,I166217,I166214,I166235,I166220,I166229,I166214,I166211,I166226,I166281,I166284,I166287,I166290,I166293,I166296,I166299,I166302,I166305,I2224,I2231);
PAT_6 I_2323 (I166284,I166281,I166287,I166299,I166296,I166290,I166293,I166281,I166302,I166284,I166305,I166351,I166354,I166357,I166360,I166363,I166366,I166369,I166372,I166375,I166378,I2224,I2231);
PAT_9 I_2324 (I166351,I166378,I166375,I166357,I166363,I166354,I166366,I166351,I166369,I166360,I166372,I166424,I166427,I166430,I166433,I166436,I166439,I166442,I166445,I166448,I2224,I2231);
PAT_2 I_2325 (I166439,I166442,I166433,I166448,I166424,I166427,I166430,I166427,I166445,I166436,I166424,I166494,I166497,I166500,I166503,I166506,I166509,I166512,I166515,I166518,I2224,I2231);
PAT_11 I_2326 (I166497,I166509,I166494,I166506,I166503,I166515,I166512,I166497,I166518,I166500,I166494,I166564,I166567,I166570,I166573,I166576,I166579,I166582,I166585,I166588,I166591,I2224,I2231);
PAT_2 I_2327 (I166564,I166588,I166576,I166570,I166579,I166582,I166567,I166591,I166585,I166573,I166564,I166637,I166640,I166643,I166646,I166649,I166652,I166655,I166658,I166661,I2224,I2231);
PAT_9 I_2328 (I166652,I166661,I166637,I166643,I166646,I166655,I166640,I166649,I166658,I166640,I166637,I166707,I166710,I166713,I166716,I166719,I166722,I166725,I166728,I166731,I2224,I2231);
PAT_2 I_2329 (I166722,I166725,I166716,I166731,I166707,I166710,I166713,I166710,I166728,I166719,I166707,I166777,I166780,I166783,I166786,I166789,I166792,I166795,I166798,I166801,I2224,I2231);
PAT_4 I_2330 (I166777,I166783,I166801,I166795,I166792,I166789,I166780,I166798,I166777,I166780,I166786,I166847,I166850,I166853,I166856,I166859,I166862,I166865,I166868,I166871,I2224,I2231);
PAT_8 I_2331 (I166859,I166847,I166868,I166853,I166850,I166871,I166856,I166865,I166850,I166847,I166862,I166917,I166920,I166923,I166926,I166929,I166932,I166935,I166938,I166941,I2224,I2231);
PAT_4 I_2332 (I166935,I166920,I166926,I166917,I166917,I166929,I166920,I166938,I166941,I166923,I166932,I166987,I166990,I166993,I166996,I166999,I167002,I167005,I167008,I167011,I2224,I2231);
PAT_13 I_2333 (I167002,I166996,I167008,I166993,I166999,I166987,I167011,I167005,I166990,I166987,I166990,I167057,I167060,I167063,I167066,I167069,I167072,I167075,I167078,I167081,I2224,I2231);
PAT_2 I_2334 (I167075,I167069,I167066,I167072,I167057,I167081,I167060,I167078,I167057,I167063,I167060,I167127,I167130,I167133,I167136,I167139,I167142,I167145,I167148,I167151,I2224,I2231);
PAT_9 I_2335 (I167142,I167151,I167127,I167133,I167136,I167145,I167130,I167139,I167148,I167130,I167127,I167197,I167200,I167203,I167206,I167209,I167212,I167215,I167218,I167221,I2224,I2231);
PAT_14 I_2336 (I167206,I167197,I167221,I167203,I167200,I167197,I167212,I167218,I167209,I167200,I167215,I167267,I167270,I167273,I167276,I167279,I167282,I167285,I167288,I167291,I2224,I2231);
PAT_4 I_2337 (I167276,I167282,I167273,I167267,I167291,I167279,I167267,I167270,I167288,I167270,I167285,I167337,I167340,I167343,I167346,I167349,I167352,I167355,I167358,I167361,I2224,I2231);
PAT_11 I_2338 (I167349,I167358,I167340,I167352,I167337,I167340,I167337,I167346,I167361,I167355,I167343,I167407,I167410,I167413,I167416,I167419,I167422,I167425,I167428,I167431,I167434,I2224,I2231);
PAT_5 I_2339 (I167428,I167407,I167434,I167422,I167419,I167431,I167413,I167407,I167425,I167410,I167416,I167480,I167483,I167486,I167489,I167492,I167495,I167498,I167501,I167504,I167507,I2224,I2231);
PAT_17 I_2340 (I167507,I167483,I167486,I167489,I167480,I167492,I167480,I167504,I167498,I167495,I167501,I167553,I167556,I167559,I167562,I167565,I167568,I167571,I167574,I167577,I167580,I2224,I2231);
PAT_5 I_2341 (I167565,I167559,I167556,I167577,I167562,I167568,I167571,I167553,I167553,I167574,I167580,I167626,I167629,I167632,I167635,I167638,I167641,I167644,I167647,I167650,I167653,I2224,I2231);
PAT_6 I_2342 (I167644,I167638,I167626,I167632,I167629,I167635,I167641,I167626,I167650,I167647,I167653,I167699,I167702,I167705,I167708,I167711,I167714,I167717,I167720,I167723,I167726,I2224,I2231);
PAT_5 I_2343 (I167720,I167699,I167705,I167708,I167714,I167717,I167699,I167723,I167702,I167711,I167726,I167772,I167775,I167778,I167781,I167784,I167787,I167790,I167793,I167796,I167799,I2224,I2231);
PAT_0 I_2344 (I167793,I167772,I167799,I167796,I167772,I167790,I167784,I167775,I167781,I167787,I167778,I167845,I167848,I167851,I167854,I167857,I167860,I167863,I167866,I2224,I2231);
PAT_12 I_2345 (I167857,I167866,I167848,I167848,I167845,I167845,I167854,I167851,I167860,I167863,I167851,I167912,I167915,I167918,I167921,I167924,I167927,I167930,I167933,I2224,I2231);
PAT_4 I_2346 (I167918,I167915,I167930,I167933,I167927,I167921,I167912,I167912,I167918,I167924,I167915,I167979,I167982,I167985,I167988,I167991,I167994,I167997,I168000,I168003,I2224,I2231);
PAT_9 I_2347 (I168000,I167982,I167985,I167994,I167997,I167979,I167988,I167982,I168003,I167979,I167991,I168049,I168052,I168055,I168058,I168061,I168064,I168067,I168070,I168073,I2224,I2231);
PAT_8 I_2348 (I168070,I168058,I168067,I168049,I168052,I168064,I168073,I168052,I168055,I168061,I168049,I168119,I168122,I168125,I168128,I168131,I168134,I168137,I168140,I168143,I2224,I2231);
PAT_11 I_2349 (I168140,I168131,I168119,I168122,I168137,I168125,I168128,I168119,I168143,I168134,I168122,I168189,I168192,I168195,I168198,I168201,I168204,I168207,I168210,I168213,I168216,I2224,I2231);
PAT_0 I_2350 (I168189,I168198,I168192,I168189,I168207,I168213,I168195,I168216,I168204,I168210,I168201,I168262,I168265,I168268,I168271,I168274,I168277,I168280,I168283,I2224,I2231);
PAT_2 I_2351 (I168268,I168271,I168280,I168265,I168268,I168265,I168274,I168262,I168262,I168277,I168283,I168329,I168332,I168335,I168338,I168341,I168344,I168347,I168350,I168353,I2224,I2231);
PAT_6 I_2352 (I168353,I168329,I168344,I168341,I168347,I168338,I168332,I168350,I168329,I168335,I168332,I168399,I168402,I168405,I168408,I168411,I168414,I168417,I168420,I168423,I168426,I2224,I2231);
PAT_13 I_2353 (I168423,I168405,I168420,I168399,I168402,I168408,I168426,I168411,I168417,I168399,I168414,I168472,I168475,I168478,I168481,I168484,I168487,I168490,I168493,I168496,I2224,I2231);
PAT_4 I_2354 (I168481,I168484,I168496,I168478,I168493,I168490,I168475,I168487,I168475,I168472,I168472,I168542,I168545,I168548,I168551,I168554,I168557,I168560,I168563,I168566,I2224,I2231);
PAT_11 I_2355 (I168554,I168563,I168545,I168557,I168542,I168545,I168542,I168551,I168566,I168560,I168548,I168612,I168615,I168618,I168621,I168624,I168627,I168630,I168633,I168636,I168639,I2224,I2231);
PAT_4 I_2356 (I168618,I168639,I168612,I168630,I168621,I168612,I168633,I168615,I168624,I168636,I168627,I168685,I168688,I168691,I168694,I168697,I168700,I168703,I168706,I168709,I2224,I2231);
PAT_10 I_2357 (I168685,I168685,I168709,I168688,I168694,I168703,I168700,I168688,I168706,I168691,I168697,I168755,I168758,I168761,I168764,I168767,I168770,I168773,I168776,I2224,I2231);
PAT_5 I_2358 (I168776,I168755,I168764,I168758,I168773,I168770,I168761,I168761,I168755,I168758,I168767,I168822,I168825,I168828,I168831,I168834,I168837,I168840,I168843,I168846,I168849,I2224,I2231);
PAT_2 I_2359 (I168837,I168822,I168834,I168828,I168843,I168825,I168840,I168831,I168846,I168849,I168822,I168895,I168898,I168901,I168904,I168907,I168910,I168913,I168916,I168919,I2224,I2231);
PAT_12 I_2360 (I168904,I168901,I168895,I168898,I168919,I168913,I168916,I168898,I168910,I168895,I168907,I168965,I168968,I168971,I168974,I168977,I168980,I168983,I168986,I2224,I2231);
PAT_13 I_2361 (I168977,I168980,I168971,I168986,I168983,I168965,I168968,I168974,I168971,I168968,I168965,I169032,I169035,I169038,I169041,I169044,I169047,I169050,I169053,I169056,I2224,I2231);
PAT_10 I_2362 (I169053,I169047,I169041,I169035,I169056,I169035,I169044,I169032,I169032,I169050,I169038,I169102,I169105,I169108,I169111,I169114,I169117,I169120,I169123,I2224,I2231);
PAT_2 I_2363 (I169114,I169117,I169108,I169120,I169105,I169102,I169102,I169108,I169123,I169111,I169105,I169169,I169172,I169175,I169178,I169181,I169184,I169187,I169190,I169193,I2224,I2231);
PAT_9 I_2364 (I169184,I169193,I169169,I169175,I169178,I169187,I169172,I169181,I169190,I169172,I169169,I169239,I169242,I169245,I169248,I169251,I169254,I169257,I169260,I169263,I2224,I2231);
PAT_4 I_2365 (I169239,I169263,I169257,I169245,I169242,I169260,I169242,I169239,I169254,I169248,I169251,I169309,I169312,I169315,I169318,I169321,I169324,I169327,I169330,I169333,I2224,I2231);
PAT_13 I_2366 (I169324,I169318,I169330,I169315,I169321,I169309,I169333,I169327,I169312,I169309,I169312,I169379,I169382,I169385,I169388,I169391,I169394,I169397,I169400,I169403,I2224,I2231);
PAT_6 I_2367 (I169379,I169391,I169388,I169400,I169397,I169403,I169379,I169394,I169382,I169382,I169385,I169449,I169452,I169455,I169458,I169461,I169464,I169467,I169470,I169473,I169476,I2224,I2231);
PAT_13 I_2368 (I169473,I169455,I169470,I169449,I169452,I169458,I169476,I169461,I169467,I169449,I169464,I169522,I169525,I169528,I169531,I169534,I169537,I169540,I169543,I169546,I2224,I2231);
PAT_17 I_2369 (I169546,I169534,I169543,I169540,I169531,I169522,I169525,I169528,I169522,I169537,I169525,I169592,I169595,I169598,I169601,I169604,I169607,I169610,I169613,I169616,I169619,I2224,I2231);
PAT_10 I_2370 (I169592,I169598,I169619,I169601,I169616,I169595,I169610,I169604,I169613,I169607,I169592,I169665,I169668,I169671,I169674,I169677,I169680,I169683,I169686,I2224,I2231);
PAT_7 I_2371 (I169686,I169683,I169680,I169665,I169668,I169671,I169668,I169677,I169665,I169671,I169674,I169732,I169735,I169738,I169741,I169744,I169747,I169750,I169753,I169756,I2224,I2231);
PAT_15 I_2372 (I169750,I169735,I169735,I169747,I169732,I169756,I169738,I169744,I169753,I169732,I169741,I169802,I169805,I169808,I169811,I169814,I169817,I169820,I169823,I169826,I2224,I2231);
PAT_17 I_2373 (I169802,I169802,I169814,I169805,I169808,I169826,I169823,I169817,I169805,I169811,I169820,I169872,I169875,I169878,I169881,I169884,I169887,I169890,I169893,I169896,I169899,I2224,I2231);
PAT_4 I_2374 (I169881,I169872,I169890,I169887,I169899,I169896,I169875,I169872,I169878,I169884,I169893,I169945,I169948,I169951,I169954,I169957,I169960,I169963,I169966,I169969,I2224,I2231);
PAT_6 I_2375 (I169945,I169951,I169948,I169960,I169963,I169957,I169969,I169966,I169945,I169954,I169948,I170015,I170018,I170021,I170024,I170027,I170030,I170033,I170036,I170039,I170042,I2224,I2231);
PAT_5 I_2376 (I170036,I170015,I170021,I170024,I170030,I170033,I170015,I170039,I170018,I170027,I170042,I170088,I170091,I170094,I170097,I170100,I170103,I170106,I170109,I170112,I170115,I2224,I2231);
PAT_6 I_2377 (I170106,I170100,I170088,I170094,I170091,I170097,I170103,I170088,I170112,I170109,I170115,I170161,I170164,I170167,I170170,I170173,I170176,I170179,I170182,I170185,I170188,I2224,I2231);
PAT_13 I_2378 (I170185,I170167,I170182,I170161,I170164,I170170,I170188,I170173,I170179,I170161,I170176,I170234,I170237,I170240,I170243,I170246,I170249,I170252,I170255,I170258,I2224,I2231);
PAT_5 I_2379 (I170246,I170237,I170243,I170255,I170237,I170258,I170240,I170249,I170234,I170234,I170252,I170304,I170307,I170310,I170313,I170316,I170319,I170322,I170325,I170328,I170331,I2224,I2231);
PAT_17 I_2380 (I170331,I170307,I170310,I170313,I170304,I170316,I170304,I170328,I170322,I170319,I170325,I170377,I170380,I170383,I170386,I170389,I170392,I170395,I170398,I170401,I170404,I2224,I2231);
PAT_15 I_2381 (I170404,I170398,I170395,I170377,I170386,I170383,I170389,I170380,I170377,I170401,I170392,I170450,I170453,I170456,I170459,I170462,I170465,I170468,I170471,I170474,I2224,I2231);
PAT_2 I_2382 (I170453,I170453,I170456,I170462,I170450,I170450,I170459,I170474,I170468,I170471,I170465,I170520,I170523,I170526,I170529,I170532,I170535,I170538,I170541,I170544,I2224,I2231);
PAT_15 I_2383 (I170523,I170535,I170541,I170544,I170526,I170538,I170520,I170529,I170520,I170532,I170523,I170590,I170593,I170596,I170599,I170602,I170605,I170608,I170611,I170614,I2224,I2231);
PAT_5 I_2384 (I170593,I170590,I170596,I170614,I170611,I170599,I170608,I170602,I170593,I170605,I170590,I170660,I170663,I170666,I170669,I170672,I170675,I170678,I170681,I170684,I170687,I2224,I2231);
PAT_14 I_2385 (I170681,I170666,I170660,I170684,I170687,I170660,I170678,I170663,I170669,I170672,I170675,I170733,I170736,I170739,I170742,I170745,I170748,I170751,I170754,I170757,I2224,I2231);
PAT_13 I_2386 (I170742,I170757,I170736,I170745,I170733,I170736,I170751,I170739,I170733,I170754,I170748,I170803,I170806,I170809,I170812,I170815,I170818,I170821,I170824,I170827,I2224,I2231);
PAT_10 I_2387 (I170824,I170818,I170812,I170806,I170827,I170806,I170815,I170803,I170803,I170821,I170809,I170873,I170876,I170879,I170882,I170885,I170888,I170891,I170894,I2224,I2231);
PAT_14 I_2388 (I170873,I170894,I170879,I170888,I170885,I170891,I170882,I170876,I170876,I170879,I170873,I170940,I170943,I170946,I170949,I170952,I170955,I170958,I170961,I170964,I2224,I2231);
PAT_10 I_2389 (I170943,I170940,I170946,I170964,I170961,I170955,I170943,I170958,I170940,I170952,I170949,I171010,I171013,I171016,I171019,I171022,I171025,I171028,I171031,I2224,I2231);
PAT_5 I_2390 (I171031,I171010,I171019,I171013,I171028,I171025,I171016,I171016,I171010,I171013,I171022,I171077,I171080,I171083,I171086,I171089,I171092,I171095,I171098,I171101,I171104,I2224,I2231);
PAT_11 I_2391 (I171089,I171086,I171080,I171098,I171101,I171077,I171095,I171092,I171104,I171083,I171077,I171150,I171153,I171156,I171159,I171162,I171165,I171168,I171171,I171174,I171177,I2224,I2231);
PAT_17 I_2392 (I171162,I171153,I171177,I171150,I171159,I171171,I171168,I171165,I171150,I171174,I171156,I171223,I171226,I171229,I171232,I171235,I171238,I171241,I171244,I171247,I171250,I2224,I2231);
PAT_5 I_2393 (I171235,I171229,I171226,I171247,I171232,I171238,I171241,I171223,I171223,I171244,I171250,I171296,I171299,I171302,I171305,I171308,I171311,I171314,I171317,I171320,I171323,I2224,I2231);
PAT_17 I_2394 (I171323,I171299,I171302,I171305,I171296,I171308,I171296,I171320,I171314,I171311,I171317,I171369,I171372,I171375,I171378,I171381,I171384,I171387,I171390,I171393,I171396,I2224,I2231);
PAT_9 I_2395 (I171390,I171372,I171378,I171393,I171375,I171387,I171369,I171381,I171369,I171396,I171384,I171442,I171445,I171448,I171451,I171454,I171457,I171460,I171463,I171466,I2224,I2231);
PAT_5 I_2396 (I171463,I171442,I171457,I171442,I171448,I171451,I171445,I171445,I171460,I171454,I171466,I171512,I171515,I171518,I171521,I171524,I171527,I171530,I171533,I171536,I171539,I2224,I2231);
PAT_7 I_2397 (I171530,I171533,I171539,I171536,I171521,I171518,I171512,I171524,I171512,I171515,I171527,I171585,I171588,I171591,I171594,I171597,I171600,I171603,I171606,I171609,I2224,I2231);
PAT_13 I_2398 (I171591,I171609,I171600,I171585,I171597,I171585,I171606,I171588,I171594,I171588,I171603,I171655,I171658,I171661,I171664,I171667,I171670,I171673,I171676,I171679,I2224,I2231);
PAT_4 I_2399 (I171664,I171667,I171679,I171661,I171676,I171673,I171658,I171670,I171658,I171655,I171655,I171725,I171728,I171731,I171734,I171737,I171740,I171743,I171746,I171749,I2224,I2231);
PAT_9 I_2400 (I171746,I171728,I171731,I171740,I171743,I171725,I171734,I171728,I171749,I171725,I171737,I171795,I171798,I171801,I171804,I171807,I171810,I171813,I171816,I171819,I2224,I2231);
PAT_11 I_2401 (I171807,I171813,I171819,I171816,I171804,I171798,I171798,I171795,I171810,I171795,I171801,I171865,I171868,I171871,I171874,I171877,I171880,I171883,I171886,I171889,I171892,I2224,I2231);
PAT_5 I_2402 (I171886,I171865,I171892,I171880,I171877,I171889,I171871,I171865,I171883,I171868,I171874,I171938,I171941,I171944,I171947,I171950,I171953,I171956,I171959,I171962,I171965,I2224,I2231);
PAT_2 I_2403 (I171953,I171938,I171950,I171944,I171959,I171941,I171956,I171947,I171962,I171965,I171938,I172011,I172014,I172017,I172020,I172023,I172026,I172029,I172032,I172035,I2224,I2231);
PAT_12 I_2404 (I172020,I172017,I172011,I172014,I172035,I172029,I172032,I172014,I172026,I172011,I172023,I172081,I172084,I172087,I172090,I172093,I172096,I172099,I172102,I2224,I2231);
PAT_6 I_2405 (I172090,I172084,I172102,I172087,I172084,I172087,I172096,I172081,I172099,I172081,I172093,I172148,I172151,I172154,I172157,I172160,I172163,I172166,I172169,I172172,I172175,I2224,I2231);
PAT_5 I_2406 (I172169,I172148,I172154,I172157,I172163,I172166,I172148,I172172,I172151,I172160,I172175,I172221,I172224,I172227,I172230,I172233,I172236,I172239,I172242,I172245,I172248,I2224,I2231);
PAT_6 I_2407 (I172239,I172233,I172221,I172227,I172224,I172230,I172236,I172221,I172245,I172242,I172248,I172294,I172297,I172300,I172303,I172306,I172309,I172312,I172315,I172318,I172321,I2224,I2231);
PAT_9 I_2408 (I172294,I172321,I172318,I172300,I172306,I172297,I172309,I172294,I172312,I172303,I172315,I172367,I172370,I172373,I172376,I172379,I172382,I172385,I172388,I172391,I2224,I2231);
PAT_6 I_2409 (I172385,I172367,I172379,I172388,I172367,I172376,I172373,I172391,I172382,I172370,I172370,I172437,I172440,I172443,I172446,I172449,I172452,I172455,I172458,I172461,I172464,I2224,I2231);
PAT_12 I_2410 (I172437,I172464,I172443,I172446,I172440,I172437,I172458,I172452,I172455,I172449,I172461,I172510,I172513,I172516,I172519,I172522,I172525,I172528,I172531,I2224,I2231);
PAT_4 I_2411 (I172516,I172513,I172528,I172531,I172525,I172519,I172510,I172510,I172516,I172522,I172513,I172577,I172580,I172583,I172586,I172589,I172592,I172595,I172598,I172601,I2224,I2231);
PAT_2 I_2412 (I172586,I172580,I172580,I172601,I172577,I172595,I172592,I172583,I172577,I172589,I172598,I172647,I172650,I172653,I172656,I172659,I172662,I172665,I172668,I172671,I2224,I2231);
PAT_8 I_2413 (I172659,I172650,I172656,I172647,I172653,I172668,I172665,I172647,I172662,I172650,I172671,I172717,I172720,I172723,I172726,I172729,I172732,I172735,I172738,I172741,I2224,I2231);
PAT_5 I_2414 (I172723,I172741,I172717,I172738,I172726,I172729,I172720,I172717,I172720,I172732,I172735,I172787,I172790,I172793,I172796,I172799,I172802,I172805,I172808,I172811,I172814,I2224,I2231);
PAT_9 I_2415 (I172802,I172799,I172808,I172805,I172796,I172787,I172793,I172814,I172790,I172811,I172787,I172860,I172863,I172866,I172869,I172872,I172875,I172878,I172881,I172884,I2224,I2231);
PAT_14 I_2416 (I172869,I172860,I172884,I172866,I172863,I172860,I172875,I172881,I172872,I172863,I172878,I172930,I172933,I172936,I172939,I172942,I172945,I172948,I172951,I172954,I2224,I2231);
PAT_8 I_2417 (I172936,I172939,I172933,I172945,I172954,I172933,I172930,I172951,I172930,I172942,I172948,I173000,I173003,I173006,I173009,I173012,I173015,I173018,I173021,I173024,I2224,I2231);
PAT_16 I_2418 (I173021,I173000,I173000,I173009,I173006,I173018,I173003,I173012,I173015,I173024,I173003,I173070,I173073,I173076,I173079,I173082,I173085,I173088,I173091,I173094,I173097,I2224,I2231);
PAT_1 I_2419 (I173073,I173076,I173097,I173079,I173082,I173088,I173070,I173085,I173091,I173094,I173070,I173143,I173146,I173149,I173152,I173155,I173158,I173161,I173164,I173167,I2224,I2231);
PAT_13 I_2420 (I173152,I173161,I173167,I173143,I173158,I173155,I173164,I173149,I173146,I173143,I173146,I173213,I173216,I173219,I173222,I173225,I173228,I173231,I173234,I173237,I2224,I2231);
PAT_12 I_2421 (I173222,I173213,I173213,I173237,I173234,I173216,I173231,I173225,I173216,I173219,I173228,I173283,I173286,I173289,I173292,I173295,I173298,I173301,I173304,I2224,I2231);
PAT_17 I_2422 (I173298,I173292,I173286,I173283,I173283,I173289,I173289,I173301,I173304,I173286,I173295,I173350,I173353,I173356,I173359,I173362,I173365,I173368,I173371,I173374,I173377,I2224,I2231);
PAT_1 I_2423 (I173374,I173377,I173356,I173365,I173350,I173371,I173362,I173353,I173359,I173350,I173368,I173423,I173426,I173429,I173432,I173435,I173438,I173441,I173444,I173447,I2224,I2231);
PAT_9 I_2424 (I173438,I173444,I173429,I173447,I173426,I173441,I173426,I173432,I173423,I173435,I173423,I173493,I173496,I173499,I173502,I173505,I173508,I173511,I173514,I173517,I2224,I2231);
PAT_5 I_2425 (I173514,I173493,I173508,I173493,I173499,I173502,I173496,I173496,I173511,I173505,I173517,I173563,I173566,I173569,I173572,I173575,I173578,I173581,I173584,I173587,I173590,I2224,I2231);
PAT_2 I_2426 (I173578,I173563,I173575,I173569,I173584,I173566,I173581,I173572,I173587,I173590,I173563,I173636,I173639,I173642,I173645,I173648,I173651,I173654,I173657,I173660,I2224,I2231);
PAT_11 I_2427 (I173639,I173651,I173636,I173648,I173645,I173657,I173654,I173639,I173660,I173642,I173636,I173706,I173709,I173712,I173715,I173718,I173721,I173724,I173727,I173730,I173733,I2224,I2231);
PAT_10 I_2428 (I173721,I173727,I173718,I173712,I173730,I173715,I173733,I173724,I173706,I173709,I173706,I173779,I173782,I173785,I173788,I173791,I173794,I173797,I173800,I2224,I2231);
PAT_17 I_2429 (I173791,I173800,I173794,I173779,I173785,I173797,I173782,I173782,I173779,I173785,I173788,I173846,I173849,I173852,I173855,I173858,I173861,I173864,I173867,I173870,I173873,I2224,I2231);
PAT_5 I_2430 (I173858,I173852,I173849,I173870,I173855,I173861,I173864,I173846,I173846,I173867,I173873,I173919,I173922,I173925,I173928,I173931,I173934,I173937,I173940,I173943,I173946,I2224,I2231);
PAT_9 I_2431 (I173934,I173931,I173940,I173937,I173928,I173919,I173925,I173946,I173922,I173943,I173919,I173992,I173995,I173998,I174001,I174004,I174007,I174010,I174013,I174016,I2224,I2231);
PAT_12 I_2432 (I174013,I174010,I174004,I173992,I174001,I173992,I173995,I173998,I174016,I174007,I173995,I174062,I174065,I174068,I174071,I174074,I174077,I174080,I174083,I2224,I2231);
PAT_10 I_2433 (I174062,I174083,I174074,I174077,I174068,I174065,I174062,I174080,I174068,I174071,I174065,I174129,I174132,I174135,I174138,I174141,I174144,I174147,I174150,I2224,I2231);
PAT_6 I_2434 (I174150,I174144,I174138,I174132,I174129,I174135,I174129,I174135,I174132,I174141,I174147,I174196,I174199,I174202,I174205,I174208,I174211,I174214,I174217,I174220,I174223,I2224,I2231);
PAT_1 I_2435 (I174223,I174214,I174202,I174205,I174217,I174208,I174211,I174196,I174199,I174196,I174220,I174269,I174272,I174275,I174278,I174281,I174284,I174287,I174290,I174293,I2224,I2231);
PAT_11 I_2436 (I174272,I174287,I174284,I174290,I174293,I174272,I174278,I174281,I174269,I174275,I174269,I174339,I174342,I174345,I174348,I174351,I174354,I174357,I174360,I174363,I174366,I2224,I2231);
PAT_4 I_2437 (I174345,I174366,I174339,I174357,I174348,I174339,I174360,I174342,I174351,I174363,I174354,I174412,I174415,I174418,I174421,I174424,I174427,I174430,I174433,I174436,I2224,I2231);
PAT_10 I_2438 (I174412,I174412,I174436,I174415,I174421,I174430,I174427,I174415,I174433,I174418,I174424,I174482,I174485,I174488,I174491,I174494,I174497,I174500,I174503,I2224,I2231);
PAT_7 I_2439 (I174503,I174500,I174497,I174482,I174485,I174488,I174485,I174494,I174482,I174488,I174491,I174549,I174552,I174555,I174558,I174561,I174564,I174567,I174570,I174573,I2224,I2231);
PAT_15 I_2440 (I174567,I174552,I174552,I174564,I174549,I174573,I174555,I174561,I174570,I174549,I174558,I174619,I174622,I174625,I174628,I174631,I174634,I174637,I174640,I174643,I2224,I2231);
PAT_5 I_2441 (I174622,I174619,I174625,I174643,I174640,I174628,I174637,I174631,I174622,I174634,I174619,I174689,I174692,I174695,I174698,I174701,I174704,I174707,I174710,I174713,I174716,I2224,I2231);
PAT_17 I_2442 (I174716,I174692,I174695,I174698,I174689,I174701,I174689,I174713,I174707,I174704,I174710,I174762,I174765,I174768,I174771,I174774,I174777,I174780,I174783,I174786,I174789,I2224,I2231);
PAT_5 I_2443 (I174774,I174768,I174765,I174786,I174771,I174777,I174780,I174762,I174762,I174783,I174789,I174835,I174838,I174841,I174844,I174847,I174850,I174853,I174856,I174859,I174862,I2224,I2231);
PAT_4 I_2444 (I174853,I174859,I174862,I174841,I174844,I174856,I174838,I174835,I174847,I174850,I174835,I174908,I174911,I174914,I174917,I174920,I174923,I174926,I174929,I174932,I2224,I2231);
PAT_2 I_2445 (I174917,I174911,I174911,I174932,I174908,I174926,I174923,I174914,I174908,I174920,I174929,I174978,I174981,I174984,I174987,I174990,I174993,I174996,I174999,I175002,I2224,I2231);
PAT_9 I_2446 (I174993,I175002,I174978,I174984,I174987,I174996,I174981,I174990,I174999,I174981,I174978,I175048,I175051,I175054,I175057,I175060,I175063,I175066,I175069,I175072,I2224,I2231);
PAT_4 I_2447 (I175048,I175072,I175066,I175054,I175051,I175069,I175051,I175048,I175063,I175057,I175060,I175118,I175121,I175124,I175127,I175130,I175133,I175136,I175139,I175142,I2224,I2231);
PAT_12 I_2448 (I175118,I175121,I175139,I175142,I175133,I175124,I175130,I175127,I175118,I175136,I175121,I175188,I175191,I175194,I175197,I175200,I175203,I175206,I175209,I2224,I2231);
PAT_8 I_2449 (I175188,I175197,I175194,I175191,I175203,I175188,I175191,I175194,I175206,I175200,I175209,I175255,I175258,I175261,I175264,I175267,I175270,I175273,I175276,I175279,I2224,I2231);
PAT_4 I_2450 (I175273,I175258,I175264,I175255,I175255,I175267,I175258,I175276,I175279,I175261,I175270,I175325,I175328,I175331,I175334,I175337,I175340,I175343,I175346,I175349,I2224,I2231);
PAT_11 I_2451 (I175337,I175346,I175328,I175340,I175325,I175328,I175325,I175334,I175349,I175343,I175331,I175395,I175398,I175401,I175404,I175407,I175410,I175413,I175416,I175419,I175422,I2224,I2231);
PAT_9 I_2452 (I175401,I175413,I175404,I175416,I175395,I175398,I175407,I175395,I175410,I175419,I175422,I175468,I175471,I175474,I175477,I175480,I175483,I175486,I175489,I175492,I2224,I2231);
PAT_11 I_2453 (I175480,I175486,I175492,I175489,I175477,I175471,I175471,I175468,I175483,I175468,I175474,I175538,I175541,I175544,I175547,I175550,I175553,I175556,I175559,I175562,I175565,I2224,I2231);
PAT_5 I_2454 (I175559,I175538,I175565,I175553,I175550,I175562,I175544,I175538,I175556,I175541,I175547,I175611,I175614,I175617,I175620,I175623,I175626,I175629,I175632,I175635,I175638,I2224,I2231);
PAT_8 I_2455 (I175611,I175638,I175629,I175626,I175620,I175611,I175623,I175635,I175614,I175632,I175617,I175684,I175687,I175690,I175693,I175696,I175699,I175702,I175705,I175708,I2224,I2231);
PAT_13 I_2456 (I175696,I175705,I175687,I175708,I175690,I175684,I175684,I175693,I175702,I175699,I175687,I175754,I175757,I175760,I175763,I175766,I175769,I175772,I175775,I175778,I2224,I2231);
PAT_4 I_2457 (I175763,I175766,I175778,I175760,I175775,I175772,I175757,I175769,I175757,I175754,I175754,I175824,I175827,I175830,I175833,I175836,I175839,I175842,I175845,I175848,I2224,I2231);
PAT_12 I_2458 (I175824,I175827,I175845,I175848,I175839,I175830,I175836,I175833,I175824,I175842,I175827,I175894,I175897,I175900,I175903,I175906,I175909,I175912,I175915,I2224,I2231);
PAT_17 I_2459 (I175909,I175903,I175897,I175894,I175894,I175900,I175900,I175912,I175915,I175897,I175906,I175961,I175964,I175967,I175970,I175973,I175976,I175979,I175982,I175985,I175988,I2224,I2231);
PAT_11 I_2460 (I175973,I175982,I175988,I175964,I175961,I175979,I175970,I175976,I175967,I175985,I175961,I176034,I176037,I176040,I176043,I176046,I176049,I176052,I176055,I176058,I176061,I2224,I2231);
PAT_5 I_2461 (I176055,I176034,I176061,I176049,I176046,I176058,I176040,I176034,I176052,I176037,I176043,I176107,I176110,I176113,I176116,I176119,I176122,I176125,I176128,I176131,I176134,I2224,I2231);
PAT_6 I_2462 (I176125,I176119,I176107,I176113,I176110,I176116,I176122,I176107,I176131,I176128,I176134,I176180,I176183,I176186,I176189,I176192,I176195,I176198,I176201,I176204,I176207,I2224,I2231);
PAT_12 I_2463 (I176180,I176207,I176186,I176189,I176183,I176180,I176201,I176195,I176198,I176192,I176204,I176253,I176256,I176259,I176262,I176265,I176268,I176271,I176274,I2224,I2231);
PAT_8 I_2464 (I176253,I176262,I176259,I176256,I176268,I176253,I176256,I176259,I176271,I176265,I176274,I176320,I176323,I176326,I176329,I176332,I176335,I176338,I176341,I176344,I2224,I2231);
PAT_17 I_2465 (I176344,I176332,I176329,I176323,I176326,I176338,I176320,I176323,I176320,I176335,I176341,I176390,I176393,I176396,I176399,I176402,I176405,I176408,I176411,I176414,I176417,I2224,I2231);
PAT_1 I_2466 (I176414,I176417,I176396,I176405,I176390,I176411,I176402,I176393,I176399,I176390,I176408,I176463,I176466,I176469,I176472,I176475,I176478,I176481,I176484,I176487,I2224,I2231);
PAT_9 I_2467 (I176478,I176484,I176469,I176487,I176466,I176481,I176466,I176472,I176463,I176475,I176463,I176533,I176536,I176539,I176542,I176545,I176548,I176551,I176554,I176557,I2224,I2231);
PAT_4 I_2468 (I176533,I176557,I176551,I176539,I176536,I176554,I176536,I176533,I176548,I176542,I176545,I176603,I176606,I176609,I176612,I176615,I176618,I176621,I176624,I176627,I2224,I2231);
PAT_9 I_2469 (I176624,I176606,I176609,I176618,I176621,I176603,I176612,I176606,I176627,I176603,I176615,I176673,I176676,I176679,I176682,I176685,I176688,I176691,I176694,I176697,I2224,I2231);
PAT_6 I_2470 (I176691,I176673,I176685,I176694,I176673,I176682,I176679,I176697,I176688,I176676,I176676,I176743,I176746,I176749,I176752,I176755,I176758,I176761,I176764,I176767,I176770,I2224,I2231);
PAT_5 I_2471 (I176764,I176743,I176749,I176752,I176758,I176761,I176743,I176767,I176746,I176755,I176770,I176816,I176819,I176822,I176825,I176828,I176831,I176834,I176837,I176840,I176843,I2224,I2231);
PAT_13 I_2472 (I176822,I176831,I176816,I176819,I176840,I176825,I176837,I176816,I176834,I176843,I176828,I176889,I176892,I176895,I176898,I176901,I176904,I176907,I176910,I176913,I2224,I2231);
PAT_3 I_2473 (I176913,I176892,I176907,I176895,I176901,I176910,I176889,I176898,I176889,I176892,I176904,I176959,I176962,I176965,I176968,I176971,I176974,I176977,I176980,I176983,I176986,I2224,I2231);
PAT_12 I_2474 (I176974,I176980,I176959,I176986,I176977,I176968,I176971,I176962,I176959,I176965,I176983,I177032,I177035,I177038,I177041,I177044,I177047,I177050,I177053,I2224,I2231);
PAT_4 I_2475 (I177038,I177035,I177050,I177053,I177047,I177041,I177032,I177032,I177038,I177044,I177035,I177099,I177102,I177105,I177108,I177111,I177114,I177117,I177120,I177123,I2224,I2231);
PAT_13 I_2476 (I177114,I177108,I177120,I177105,I177111,I177099,I177123,I177117,I177102,I177099,I177102,I177169,I177172,I177175,I177178,I177181,I177184,I177187,I177190,I177193,I2224,I2231);
PAT_10 I_2477 (I177190,I177184,I177178,I177172,I177193,I177172,I177181,I177169,I177169,I177187,I177175,I177239,I177242,I177245,I177248,I177251,I177254,I177257,I177260,I2224,I2231);
PAT_0 I_2478 (I177242,I177245,I177254,I177242,I177260,I177257,I177251,I177239,I177245,I177248,I177239,I177306,I177309,I177312,I177315,I177318,I177321,I177324,I177327,I2224,I2231);
PAT_11 I_2479 (I177312,I177321,I177327,I177306,I177324,I177312,I177309,I177315,I177318,I177306,I177309,I177373,I177376,I177379,I177382,I177385,I177388,I177391,I177394,I177397,I177400,I2224,I2231);
PAT_1 I_2480 (I177388,I177379,I177382,I177373,I177394,I177391,I177376,I177373,I177400,I177397,I177385,I177446,I177449,I177452,I177455,I177458,I177461,I177464,I177467,I177470,I2224,I2231);
PAT_9 I_2481 (I177461,I177467,I177452,I177470,I177449,I177464,I177449,I177455,I177446,I177458,I177446,I177516,I177519,I177522,I177525,I177528,I177531,I177534,I177537,I177540,I2224,I2231);
PAT_1 I_2482 (I177516,I177534,I177516,I177528,I177519,I177525,I177531,I177537,I177540,I177522,I177519,I177586,I177589,I177592,I177595,I177598,I177601,I177604,I177607,I177610,I2224,I2231);
PAT_4 I_2483 (I177598,I177604,I177586,I177589,I177592,I177595,I177607,I177589,I177601,I177586,I177610,I177656,I177659,I177662,I177665,I177668,I177671,I177674,I177677,I177680,I2224,I2231);
PAT_1 I_2484 (I177656,I177677,I177674,I177659,I177671,I177656,I177659,I177680,I177665,I177662,I177668,I177726,I177729,I177732,I177735,I177738,I177741,I177744,I177747,I177750,I2224,I2231);
PAT_13 I_2485 (I177735,I177744,I177750,I177726,I177741,I177738,I177747,I177732,I177729,I177726,I177729,I177796,I177799,I177802,I177805,I177808,I177811,I177814,I177817,I177820,I2224,I2231);
PAT_9 I_2486 (I177817,I177799,I177799,I177796,I177820,I177802,I177805,I177796,I177808,I177814,I177811,I177866,I177869,I177872,I177875,I177878,I177881,I177884,I177887,I177890,I2224,I2231);
PAT_17 I_2487 (I177869,I177875,I177890,I177881,I177884,I177872,I177866,I177878,I177866,I177869,I177887,I177936,I177939,I177942,I177945,I177948,I177951,I177954,I177957,I177960,I177963,I2224,I2231);
PAT_9 I_2488 (I177957,I177939,I177945,I177960,I177942,I177954,I177936,I177948,I177936,I177963,I177951,I178009,I178012,I178015,I178018,I178021,I178024,I178027,I178030,I178033,I2224,I2231);
PAT_13 I_2489 (I178009,I178030,I178012,I178027,I178021,I178018,I178033,I178009,I178015,I178024,I178012,I178079,I178082,I178085,I178088,I178091,I178094,I178097,I178100,I178103,I2224,I2231);
PAT_7 I_2490 (I178088,I178091,I178079,I178094,I178100,I178085,I178082,I178103,I178082,I178079,I178097,I178149,I178152,I178155,I178158,I178161,I178164,I178167,I178170,I178173,I2224,I2231);
PAT_13 I_2491 (I178155,I178173,I178164,I178149,I178161,I178149,I178170,I178152,I178158,I178152,I178167,I178219,I178222,I178225,I178228,I178231,I178234,I178237,I178240,I178243,I2224,I2231);
PAT_14 I_2492 (I178222,I178237,I178225,I178234,I178228,I178219,I178231,I178240,I178219,I178243,I178222,I178289,I178292,I178295,I178298,I178301,I178304,I178307,I178310,I178313,I2224,I2231);
PAT_17 I_2493 (I178304,I178292,I178313,I178289,I178310,I178298,I178295,I178307,I178301,I178292,I178289,I178359,I178362,I178365,I178368,I178371,I178374,I178377,I178380,I178383,I178386,I2224,I2231);
PAT_9 I_2494 (I178380,I178362,I178368,I178383,I178365,I178377,I178359,I178371,I178359,I178386,I178374,I178432,I178435,I178438,I178441,I178444,I178447,I178450,I178453,I178456,I2224,I2231);
PAT_4 I_2495 (I178432,I178456,I178450,I178438,I178435,I178453,I178435,I178432,I178447,I178441,I178444,I178502,I178505,I178508,I178511,I178514,I178517,I178520,I178523,I178526,I2224,I2231);
PAT_9 I_2496 (I178523,I178505,I178508,I178517,I178520,I178502,I178511,I178505,I178526,I178502,I178514,I178572,I178575,I178578,I178581,I178584,I178587,I178590,I178593,I178596,I2224,I2231);
PAT_5 I_2497 (I178593,I178572,I178587,I178572,I178578,I178581,I178575,I178575,I178590,I178584,I178596,I178642,I178645,I178648,I178651,I178654,I178657,I178660,I178663,I178666,I178669,I2224,I2231);
PAT_4 I_2498 (I178660,I178666,I178669,I178648,I178651,I178663,I178645,I178642,I178654,I178657,I178642,I178715,I178718,I178721,I178724,I178727,I178730,I178733,I178736,I178739,I2224,I2231);
PAT_10 I_2499 (I178715,I178715,I178739,I178718,I178724,I178733,I178730,I178718,I178736,I178721,I178727,I178785,I178788,I178791,I178794,I178797,I178800,I178803,I178806,I2224,I2231);
PAT_9 I_2500 (I178797,I178785,I178788,I178791,I178785,I178791,I178794,I178788,I178806,I178800,I178803,I178852,I178855,I178858,I178861,I178864,I178867,I178870,I178873,I178876,I2224,I2231);
PAT_10 I_2501 (I178873,I178870,I178858,I178855,I178876,I178861,I178867,I178855,I178852,I178852,I178864,I178922,I178925,I178928,I178931,I178934,I178937,I178940,I178943,I2224,I2231);
PAT_6 I_2502 (I178943,I178937,I178931,I178925,I178922,I178928,I178922,I178928,I178925,I178934,I178940,I178989,I178992,I178995,I178998,I179001,I179004,I179007,I179010,I179013,I179016,I2224,I2231);
PAT_8 I_2503 (I178998,I179004,I178995,I179007,I178989,I178992,I179010,I178989,I179016,I179013,I179001,I179062,I179065,I179068,I179071,I179074,I179077,I179080,I179083,I179086,I2224,I2231);
PAT_17 I_2504 (I179086,I179074,I179071,I179065,I179068,I179080,I179062,I179065,I179062,I179077,I179083,I179132,I179135,I179138,I179141,I179144,I179147,I179150,I179153,I179156,I179159,I2224,I2231);
PAT_11 I_2505 (I179144,I179153,I179159,I179135,I179132,I179150,I179141,I179147,I179138,I179156,I179132,I179205,I179208,I179211,I179214,I179217,I179220,I179223,I179226,I179229,I179232,I2224,I2231);
PAT_10 I_2506 (I179220,I179226,I179217,I179211,I179229,I179214,I179232,I179223,I179205,I179208,I179205,I179278,I179281,I179284,I179287,I179290,I179293,I179296,I179299,I2224,I2231);
PAT_11 I_2507 (I179287,I179290,I179299,I179293,I179296,I179278,I179278,I179284,I179281,I179281,I179284,I179345,I179348,I179351,I179354,I179357,I179360,I179363,I179366,I179369,I179372,I2224,I2231);
PAT_9 I_2508 (I179351,I179363,I179354,I179366,I179345,I179348,I179357,I179345,I179360,I179369,I179372,I179418,I179421,I179424,I179427,I179430,I179433,I179436,I179439,I179442,I2224,I2231);
PAT_6 I_2509 (I179436,I179418,I179430,I179439,I179418,I179427,I179424,I179442,I179433,I179421,I179421,I179488,I179491,I179494,I179497,I179500,I179503,I179506,I179509,I179512,I179515,I2224,I2231);
PAT_9 I_2510 (I179488,I179515,I179512,I179494,I179500,I179491,I179503,I179488,I179506,I179497,I179509,I179561,I179564,I179567,I179570,I179573,I179576,I179579,I179582,I179585,I2224,I2231);
PAT_6 I_2511 (I1585,I1705,I1553,I2017,I2185,I1913,I1961,I2089,I2065,I1545,I1641,I179631,I179634,I179637,I179640,I179643,I179646,I179649,I179652,I179655,I179658,I2224,I2231);
PAT_7 I_2512 (I179637,I179646,I179649,I179631,I179640,I179634,I179643,I179658,I179652,I179655,I179631,I179704,I179707,I179710,I179713,I179716,I179719,I179722,I179725,I179728,I2224,I2231);
PAT_10 I_2513 (I179704,I179707,I179704,I179725,I179713,I179716,I179707,I179728,I179719,I179710,I179722,I179774,I179777,I179780,I179783,I179786,I179789,I179792,I179795,I2224,I2231);
PAT_9 I_2514 (I179786,I179774,I179777,I179780,I179774,I179780,I179783,I179777,I179795,I179789,I179792,I179841,I179844,I179847,I179850,I179853,I179856,I179859,I179862,I179865,I2224,I2231);
PAT_6 I_2515 (I179859,I179841,I179853,I179862,I179841,I179850,I179847,I179865,I179856,I179844,I179844,I179911,I179914,I179917,I179920,I179923,I179926,I179929,I179932,I179935,I179938,I2224,I2231);
PAT_5 I_2516 (I179932,I179911,I179917,I179920,I179926,I179929,I179911,I179935,I179914,I179923,I179938,I179984,I179987,I179990,I179993,I179996,I179999,I180002,I180005,I180008,I180011,I2224,I2231);
PAT_2 I_2517 (I179999,I179984,I179996,I179990,I180005,I179987,I180002,I179993,I180008,I180011,I179984,I180057,I180060,I180063,I180066,I180069,I180072,I180075,I180078,I180081,I2224,I2231);
PAT_9 I_2518 (I180072,I180081,I180057,I180063,I180066,I180075,I180060,I180069,I180078,I180060,I180057,I180127,I180130,I180133,I180136,I180139,I180142,I180145,I180148,I180151,I2224,I2231);
PAT_6 I_2519 (I180145,I180127,I180139,I180148,I180127,I180136,I180133,I180151,I180142,I180130,I180130,I180197,I180200,I180203,I180206,I180209,I180212,I180215,I180218,I180221,I180224,I2224,I2231);
PAT_9 I_2520 (I180197,I180224,I180221,I180203,I180209,I180200,I180212,I180197,I180215,I180206,I180218,I180270,I180273,I180276,I180279,I180282,I180285,I180288,I180291,I180294,I2224,I2231);
PAT_13 I_2521 (I180270,I180291,I180273,I180288,I180282,I180279,I180294,I180270,I180276,I180285,I180273,I180340,I180343,I180346,I180349,I180352,I180355,I180358,I180361,I180364,I2224,I2231);
PAT_5 I_2522 (I180352,I180343,I180349,I180361,I180343,I180364,I180346,I180355,I180340,I180340,I180358,I180410,I180413,I180416,I180419,I180422,I180425,I180428,I180431,I180434,I180437,I2224,I2231);
PAT_4 I_2523 (I180428,I180434,I180437,I180416,I180419,I180431,I180413,I180410,I180422,I180425,I180410,I180483,I180486,I180489,I180492,I180495,I180498,I180501,I180504,I180507,I2224,I2231);
PAT_10 I_2524 (I180483,I180483,I180507,I180486,I180492,I180501,I180498,I180486,I180504,I180489,I180495,I180553,I180556,I180559,I180562,I180565,I180568,I180571,I180574,I2224,I2231);
PAT_11 I_2525 (I180562,I180565,I180574,I180568,I180571,I180553,I180553,I180559,I180556,I180556,I180559,I180620,I180623,I180626,I180629,I180632,I180635,I180638,I180641,I180644,I180647,I2224,I2231);
PAT_8 I_2526 (I180629,I180635,I180638,I180644,I180641,I180632,I180620,I180620,I180647,I180623,I180626,I180693,I180696,I180699,I180702,I180705,I180708,I180711,I180714,I180717,I2224,I2231);
PAT_11 I_2527 (I180714,I180705,I180693,I180696,I180711,I180699,I180702,I180693,I180717,I180708,I180696,I180763,I180766,I180769,I180772,I180775,I180778,I180781,I180784,I180787,I180790,I2224,I2231);
PAT_9 I_2528 (I180769,I180781,I180772,I180784,I180763,I180766,I180775,I180763,I180778,I180787,I180790,I180836,I180839,I180842,I180845,I180848,I180851,I180854,I180857,I180860,I2224,I2231);
PAT_2 I_2529 (I180851,I180854,I180845,I180860,I180836,I180839,I180842,I180839,I180857,I180848,I180836,I180906,I180909,I180912,I180915,I180918,I180921,I180924,I180927,I180930,I2224,I2231);
PAT_15 I_2530 (I180909,I180921,I180927,I180930,I180912,I180924,I180906,I180915,I180906,I180918,I180909,I180976,I180979,I180982,I180985,I180988,I180991,I180994,I180997,I181000,I2224,I2231);
PAT_4 I_2531 (I180988,I180994,I180976,I180979,I180982,I180976,I181000,I180997,I180985,I180991,I180979,I181046,I181049,I181052,I181055,I181058,I181061,I181064,I181067,I181070,I2224,I2231);
PAT_6 I_2532 (I181046,I181052,I181049,I181061,I181064,I181058,I181070,I181067,I181046,I181055,I181049,I181116,I181119,I181122,I181125,I181128,I181131,I181134,I181137,I181140,I181143,I2224,I2231);
PAT_12 I_2533 (I181116,I181143,I181122,I181125,I181119,I181116,I181137,I181131,I181134,I181128,I181140,I181189,I181192,I181195,I181198,I181201,I181204,I181207,I181210,I2224,I2231);
PAT_4 I_2534 (I181195,I181192,I181207,I181210,I181204,I181198,I181189,I181189,I181195,I181201,I181192,I181256,I181259,I181262,I181265,I181268,I181271,I181274,I181277,I181280,I2224,I2231);
PAT_5 I_2535 (I181277,I181259,I181259,I181271,I181274,I181268,I181265,I181256,I181262,I181256,I181280,I181326,I181329,I181332,I181335,I181338,I181341,I181344,I181347,I181350,I181353,I2224,I2231);
PAT_9 I_2536 (I181341,I181338,I181347,I181344,I181335,I181326,I181332,I181353,I181329,I181350,I181326,I181399,I181402,I181405,I181408,I181411,I181414,I181417,I181420,I181423,I2224,I2231);
PAT_13 I_2537 (I181399,I181420,I181402,I181417,I181411,I181408,I181423,I181399,I181405,I181414,I181402,I181469,I181472,I181475,I181478,I181481,I181484,I181487,I181490,I181493,I2224,I2231);
PAT_11 I_2538 (I181469,I181481,I181484,I181475,I181472,I181493,I181472,I181490,I181478,I181469,I181487,I181539,I181542,I181545,I181548,I181551,I181554,I181557,I181560,I181563,I181566,I2224,I2231);
PAT_5 I_2539 (I181560,I181539,I181566,I181554,I181551,I181563,I181545,I181539,I181557,I181542,I181548,I181612,I181615,I181618,I181621,I181624,I181627,I181630,I181633,I181636,I181639,I2224,I2231);
PAT_14 I_2540 (I181633,I181618,I181612,I181636,I181639,I181612,I181630,I181615,I181621,I181624,I181627,I181685,I181688,I181691,I181694,I181697,I181700,I181703,I181706,I181709,I2224,I2231);
PAT_10 I_2541 (I181688,I181685,I181691,I181709,I181706,I181700,I181688,I181703,I181685,I181697,I181694,I181755,I181758,I181761,I181764,I181767,I181770,I181773,I181776,I2224,I2231);
PAT_13 I_2542 (I181761,I181767,I181761,I181758,I181773,I181776,I181755,I181755,I181770,I181758,I181764,I181822,I181825,I181828,I181831,I181834,I181837,I181840,I181843,I181846,I2224,I2231);
PAT_5 I_2543 (I181834,I181825,I181831,I181843,I181825,I181846,I181828,I181837,I181822,I181822,I181840,I181892,I181895,I181898,I181901,I181904,I181907,I181910,I181913,I181916,I181919,I2224,I2231);
PAT_11 I_2544 (I181904,I181901,I181895,I181913,I181916,I181892,I181910,I181907,I181919,I181898,I181892,I181965,I181968,I181971,I181974,I181977,I181980,I181983,I181986,I181989,I181992,I2224,I2231);
PAT_4 I_2545 (I181971,I181992,I181965,I181983,I181974,I181965,I181986,I181968,I181977,I181989,I181980,I182038,I182041,I182044,I182047,I182050,I182053,I182056,I182059,I182062,I2224,I2231);
PAT_16 I_2546 (I182044,I182056,I182038,I182041,I182053,I182047,I182041,I182059,I182050,I182038,I182062,I182108,I182111,I182114,I182117,I182120,I182123,I182126,I182129,I182132,I182135,I2224,I2231);
PAT_14 I_2547 (I182114,I182123,I182108,I182108,I182111,I182129,I182126,I182117,I182132,I182135,I182120,I182181,I182184,I182187,I182190,I182193,I182196,I182199,I182202,I182205,I2224,I2231);
PAT_9 I_2548 (I182190,I182202,I182181,I182199,I182184,I182187,I182205,I182184,I182193,I182181,I182196,I182251,I182254,I182257,I182260,I182263,I182266,I182269,I182272,I182275,I2224,I2231);
PAT_11 I_2549 (I182263,I182269,I182275,I182272,I182260,I182254,I182254,I182251,I182266,I182251,I182257,I182321,I182324,I182327,I182330,I182333,I182336,I182339,I182342,I182345,I182348,I2224,I2231);
PAT_13 I_2550 (I182321,I182324,I182333,I182345,I182348,I182336,I182342,I182330,I182339,I182327,I182321,I182394,I182397,I182400,I182403,I182406,I182409,I182412,I182415,I182418,I2224,I2231);
PAT_6 I_2551 (I182394,I182406,I182403,I182415,I182412,I182418,I182394,I182409,I182397,I182397,I182400,I182464,I182467,I182470,I182473,I182476,I182479,I182482,I182485,I182488,I182491,I2224,I2231);
PAT_11 I_2552 (I182464,I182479,I182464,I182476,I182473,I182491,I182488,I182485,I182482,I182467,I182470,I182537,I182540,I182543,I182546,I182549,I182552,I182555,I182558,I182561,I182564,I2224,I2231);
PAT_10 I_2553 (I182552,I182558,I182549,I182543,I182561,I182546,I182564,I182555,I182537,I182540,I182537,I182610,I182613,I182616,I182619,I182622,I182625,I182628,I182631,I2224,I2231);
PAT_12 I_2554 (I182616,I182610,I182610,I182622,I182625,I182613,I182613,I182628,I182631,I182616,I182619,I182677,I182680,I182683,I182686,I182689,I182692,I182695,I182698,I2224,I2231);
PAT_9 I_2555 (I182686,I182692,I182677,I182683,I182689,I182680,I182677,I182680,I182698,I182683,I182695,I182744,I182747,I182750,I182753,I182756,I182759,I182762,I182765,I182768,I2224,I2231);
PAT_7 I_2556 (I182750,I182759,I182744,I182765,I182756,I182744,I182747,I182768,I182762,I182747,I182753,I182814,I182817,I182820,I182823,I182826,I182829,I182832,I182835,I182838,I2224,I2231);
PAT_11 I_2557 (I182826,I182820,I182814,I182835,I182838,I182823,I182817,I182832,I182814,I182829,I182817,I182884,I182887,I182890,I182893,I182896,I182899,I182902,I182905,I182908,I182911,I2224,I2231);
PAT_9 I_2558 (I182890,I182902,I182893,I182905,I182884,I182887,I182896,I182884,I182899,I182908,I182911,I182957,I182960,I182963,I182966,I182969,I182972,I182975,I182978,I182981,I2224,I2231);
PAT_2 I_2559 (I182972,I182975,I182966,I182981,I182957,I182960,I182963,I182960,I182978,I182969,I182957,I183027,I183030,I183033,I183036,I183039,I183042,I183045,I183048,I183051,I2224,I2231);
PAT_17 I_2560 (I183027,I183027,I183039,I183030,I183033,I183045,I183042,I183051,I183030,I183036,I183048,I183097,I183100,I183103,I183106,I183109,I183112,I183115,I183118,I183121,I183124,I2224,I2231);
PAT_5 I_2561 (I183109,I183103,I183100,I183121,I183106,I183112,I183115,I183097,I183097,I183118,I183124,I183170,I183173,I183176,I183179,I183182,I183185,I183188,I183191,I183194,I183197,I2224,I2231);
PAT_13 I_2562 (I183176,I183185,I183170,I183173,I183194,I183179,I183191,I183170,I183188,I183197,I183182,I183243,I183246,I183249,I183252,I183255,I183258,I183261,I183264,I183267,I2224,I2231);
PAT_17 I_2563 (I183267,I183255,I183264,I183261,I183252,I183243,I183246,I183249,I183243,I183258,I183246,I183313,I183316,I183319,I183322,I183325,I183328,I183331,I183334,I183337,I183340,I2224,I2231);
PAT_4 I_2564 (I183322,I183313,I183331,I183328,I183340,I183337,I183316,I183313,I183319,I183325,I183334,I183386,I183389,I183392,I183395,I183398,I183401,I183404,I183407,I183410,I2224,I2231);
PAT_16 I_2565 (I183392,I183404,I183386,I183389,I183401,I183395,I183389,I183407,I183398,I183386,I183410,I183456,I183459,I183462,I183465,I183468,I183471,I183474,I183477,I183480,I183483,I2224,I2231);
PAT_10 I_2566 (I183456,I183468,I183483,I183471,I183477,I183480,I183465,I183456,I183474,I183462,I183459,I183529,I183532,I183535,I183538,I183541,I183544,I183547,I183550,I2224,I2231);
PAT_11 I_2567 (I183538,I183541,I183550,I183544,I183547,I183529,I183529,I183535,I183532,I183532,I183535,I183596,I183599,I183602,I183605,I183608,I183611,I183614,I183617,I183620,I183623,I2224,I2231);
PAT_5 I_2568 (I183617,I183596,I183623,I183611,I183608,I183620,I183602,I183596,I183614,I183599,I183605,I183669,I183672,I183675,I183678,I183681,I183684,I183687,I183690,I183693,I183696,I2224,I2231);
PAT_3 I_2569 (I183681,I183669,I183696,I183690,I183693,I183669,I183684,I183672,I183675,I183678,I183687,I183742,I183745,I183748,I183751,I183754,I183757,I183760,I183763,I183766,I183769,I2224,I2231);
PAT_13 I_2570 (I183763,I183751,I183769,I183748,I183754,I183757,I183745,I183760,I183742,I183742,I183766,I183815,I183818,I183821,I183824,I183827,I183830,I183833,I183836,I183839,I2224,I2231);
PAT_1 I_2571 (I183815,I183824,I183818,I183836,I183830,I183821,I183833,I183827,I183818,I183839,I183815,I183885,I183888,I183891,I183894,I183897,I183900,I183903,I183906,I183909,I2224,I2231);
PAT_15 I_2572 (I183888,I183897,I183885,I183900,I183894,I183888,I183909,I183906,I183903,I183891,I183885,I183955,I183958,I183961,I183964,I183967,I183970,I183973,I183976,I183979,I2224,I2231);
PAT_13 I_2573 (I183964,I183955,I183973,I183958,I183958,I183976,I183967,I183955,I183970,I183979,I183961,I184025,I184028,I184031,I184034,I184037,I184040,I184043,I184046,I184049,I2224,I2231);
PAT_17 I_2574 (I184049,I184037,I184046,I184043,I184034,I184025,I184028,I184031,I184025,I184040,I184028,I184095,I184098,I184101,I184104,I184107,I184110,I184113,I184116,I184119,I184122,I2224,I2231);
PAT_12 I_2575 (I184119,I184101,I184095,I184113,I184107,I184116,I184098,I184122,I184095,I184104,I184110,I184168,I184171,I184174,I184177,I184180,I184183,I184186,I184189,I2224,I2231);
PAT_13 I_2576 (I184180,I184183,I184174,I184189,I184186,I184168,I184171,I184177,I184174,I184171,I184168,I184235,I184238,I184241,I184244,I184247,I184250,I184253,I184256,I184259,I2224,I2231);
PAT_14 I_2577 (I184238,I184253,I184241,I184250,I184244,I184235,I184247,I184256,I184235,I184259,I184238,I184305,I184308,I184311,I184314,I184317,I184320,I184323,I184326,I184329,I2224,I2231);
PAT_9 I_2578 (I184314,I184326,I184305,I184323,I184308,I184311,I184329,I184308,I184317,I184305,I184320,I184375,I184378,I184381,I184384,I184387,I184390,I184393,I184396,I184399,I2224,I2231);
PAT_1 I_2579 (I184375,I184393,I184375,I184387,I184378,I184384,I184390,I184396,I184399,I184381,I184378,I184445,I184448,I184451,I184454,I184457,I184460,I184463,I184466,I184469,I2224,I2231);
PAT_5 I_2580 (I184463,I184466,I184448,I184457,I184454,I184451,I184460,I184469,I184448,I184445,I184445,I184515,I184518,I184521,I184524,I184527,I184530,I184533,I184536,I184539,I184542,I2224,I2231);
PAT_10 I_2581 (I184539,I184542,I184521,I184527,I184530,I184536,I184518,I184515,I184515,I184524,I184533,I184588,I184591,I184594,I184597,I184600,I184603,I184606,I184609,I2224,I2231);
PAT_12 I_2582 (I184594,I184588,I184588,I184600,I184603,I184591,I184591,I184606,I184609,I184594,I184597,I184655,I184658,I184661,I184664,I184667,I184670,I184673,I184676,I2224,I2231);
PAT_10 I_2583 (I184655,I184676,I184667,I184670,I184661,I184658,I184655,I184673,I184661,I184664,I184658,I184722,I184725,I184728,I184731,I184734,I184737,I184740,I184743,I2224,I2231);
PAT_13 I_2584 (I184728,I184734,I184728,I184725,I184740,I184743,I184722,I184722,I184737,I184725,I184731,I184789,I184792,I184795,I184798,I184801,I184804,I184807,I184810,I184813,I2224,I2231);
PAT_14 I_2585 (I184792,I184807,I184795,I184804,I184798,I184789,I184801,I184810,I184789,I184813,I184792,I184859,I184862,I184865,I184868,I184871,I184874,I184877,I184880,I184883,I2224,I2231);
PAT_9 I_2586 (I184868,I184880,I184859,I184877,I184862,I184865,I184883,I184862,I184871,I184859,I184874,I184929,I184932,I184935,I184938,I184941,I184944,I184947,I184950,I184953,I2224,I2231);
PAT_4 I_2587 (I184929,I184953,I184947,I184935,I184932,I184950,I184932,I184929,I184944,I184938,I184941,I184999,I185002,I185005,I185008,I185011,I185014,I185017,I185020,I185023,I2224,I2231);
PAT_14 I_2588 (I185002,I185017,I185014,I184999,I185011,I185002,I184999,I185005,I185020,I185008,I185023,I185069,I185072,I185075,I185078,I185081,I185084,I185087,I185090,I185093,I2224,I2231);
PAT_10 I_2589 (I185072,I185069,I185075,I185093,I185090,I185084,I185072,I185087,I185069,I185081,I185078,I185139,I185142,I185145,I185148,I185151,I185154,I185157,I185160,I2224,I2231);
PAT_2 I_2590 (I185151,I185154,I185145,I185157,I185142,I185139,I185139,I185145,I185160,I185148,I185142,I185206,I185209,I185212,I185215,I185218,I185221,I185224,I185227,I185230,I2224,I2231);
PAT_5 I_2591 (I185227,I185206,I185206,I185218,I185215,I185224,I185212,I185221,I185230,I185209,I185209,I185276,I185279,I185282,I185285,I185288,I185291,I185294,I185297,I185300,I185303,I2224,I2231);
PAT_13 I_2592 (I185282,I185291,I185276,I185279,I185300,I185285,I185297,I185276,I185294,I185303,I185288,I185349,I185352,I185355,I185358,I185361,I185364,I185367,I185370,I185373,I2224,I2231);
PAT_1 I_2593 (I185349,I185358,I185352,I185370,I185364,I185355,I185367,I185361,I185352,I185373,I185349,I185419,I185422,I185425,I185428,I185431,I185434,I185437,I185440,I185443,I2224,I2231);
PAT_10 I_2594 (I185434,I185431,I185422,I185419,I185422,I185437,I185425,I185440,I185443,I185428,I185419,I185489,I185492,I185495,I185498,I185501,I185504,I185507,I185510,I2224,I2231);
PAT_15 I_2595 (I185504,I185507,I185495,I185501,I185489,I185489,I185495,I185510,I185498,I185492,I185492,I185556,I185559,I185562,I185565,I185568,I185571,I185574,I185577,I185580,I2224,I2231);
PAT_13 I_2596 (I185565,I185556,I185574,I185559,I185559,I185577,I185568,I185556,I185571,I185580,I185562,I185626,I185629,I185632,I185635,I185638,I185641,I185644,I185647,I185650,I2224,I2231);
PAT_8 I_2597 (I185635,I185647,I185638,I185641,I185650,I185629,I185644,I185626,I185629,I185632,I185626,I185696,I185699,I185702,I185705,I185708,I185711,I185714,I185717,I185720,I2224,I2231);
PAT_17 I_2598 (I185720,I185708,I185705,I185699,I185702,I185714,I185696,I185699,I185696,I185711,I185717,I185766,I185769,I185772,I185775,I185778,I185781,I185784,I185787,I185790,I185793,I2224,I2231);
PAT_4 I_2599 (I185775,I185766,I185784,I185781,I185793,I185790,I185769,I185766,I185772,I185778,I185787,I185839,I185842,I185845,I185848,I185851,I185854,I185857,I185860,I185863,I2224,I2231);
PAT_9 I_2600 (I185860,I185842,I185845,I185854,I185857,I185839,I185848,I185842,I185863,I185839,I185851,I185909,I185912,I185915,I185918,I185921,I185924,I185927,I185930,I185933,I2224,I2231);
PAT_11 I_2601 (I185921,I185927,I185933,I185930,I185918,I185912,I185912,I185909,I185924,I185909,I185915,I185979,I185982,I185985,I185988,I185991,I185994,I185997,I186000,I186003,I186006,I2224,I2231);
PAT_10 I_2602 (I185994,I186000,I185991,I185985,I186003,I185988,I186006,I185997,I185979,I185982,I185979,I186052,I186055,I186058,I186061,I186064,I186067,I186070,I186073,I2224,I2231);
PAT_11 I_2603 (I186061,I186064,I186073,I186067,I186070,I186052,I186052,I186058,I186055,I186055,I186058,I186119,I186122,I186125,I186128,I186131,I186134,I186137,I186140,I186143,I186146,I2224,I2231);
PAT_8 I_2604 (I186128,I186134,I186137,I186143,I186140,I186131,I186119,I186119,I186146,I186122,I186125,I186192,I186195,I186198,I186201,I186204,I186207,I186210,I186213,I186216,I2224,I2231);
PAT_11 I_2605 (I186213,I186204,I186192,I186195,I186210,I186198,I186201,I186192,I186216,I186207,I186195,I186262,I186265,I186268,I186271,I186274,I186277,I186280,I186283,I186286,I186289,I2224,I2231);
PAT_2 I_2606 (I186262,I186286,I186274,I186268,I186277,I186280,I186265,I186289,I186283,I186271,I186262,I186335,I186338,I186341,I186344,I186347,I186350,I186353,I186356,I186359,I2224,I2231);
PAT_9 I_2607 (I186350,I186359,I186335,I186341,I186344,I186353,I186338,I186347,I186356,I186338,I186335,I186405,I186408,I186411,I186414,I186417,I186420,I186423,I186426,I186429,I2224,I2231);
PAT_13 I_2608 (I186405,I186426,I186408,I186423,I186417,I186414,I186429,I186405,I186411,I186420,I186408,I186475,I186478,I186481,I186484,I186487,I186490,I186493,I186496,I186499,I2224,I2231);
PAT_12 I_2609 (I186484,I186475,I186475,I186499,I186496,I186478,I186493,I186487,I186478,I186481,I186490,I186545,I186548,I186551,I186554,I186557,I186560,I186563,I186566,I2224,I2231);
PAT_6 I_2610 (I186554,I186548,I186566,I186551,I186548,I186551,I186560,I186545,I186563,I186545,I186557,I186612,I186615,I186618,I186621,I186624,I186627,I186630,I186633,I186636,I186639,I2224,I2231);
PAT_9 I_2611 (I186612,I186639,I186636,I186618,I186624,I186615,I186627,I186612,I186630,I186621,I186633,I186685,I186688,I186691,I186694,I186697,I186700,I186703,I186706,I186709,I2224,I2231);
PAT_4 I_2612 (I186685,I186709,I186703,I186691,I186688,I186706,I186688,I186685,I186700,I186694,I186697,I186755,I186758,I186761,I186764,I186767,I186770,I186773,I186776,I186779,I2224,I2231);
PAT_9 I_2613 (I186776,I186758,I186761,I186770,I186773,I186755,I186764,I186758,I186779,I186755,I186767,I186825,I186828,I186831,I186834,I186837,I186840,I186843,I186846,I186849,I2224,I2231);
PAT_4 I_2614 (I186825,I186849,I186843,I186831,I186828,I186846,I186828,I186825,I186840,I186834,I186837,I186895,I186898,I186901,I186904,I186907,I186910,I186913,I186916,I186919,I2224,I2231);
PAT_13 I_2615 (I186910,I186904,I186916,I186901,I186907,I186895,I186919,I186913,I186898,I186895,I186898,I186965,I186968,I186971,I186974,I186977,I186980,I186983,I186986,I186989,I2224,I2231);
PAT_11 I_2616 (I186965,I186977,I186980,I186971,I186968,I186989,I186968,I186986,I186974,I186965,I186983,I187035,I187038,I187041,I187044,I187047,I187050,I187053,I187056,I187059,I187062,I2224,I2231);
PAT_8 I_2617 (I187044,I187050,I187053,I187059,I187056,I187047,I187035,I187035,I187062,I187038,I187041,I187108,I187111,I187114,I187117,I187120,I187123,I187126,I187129,I187132,I2224,I2231);
PAT_13 I_2618 (I187120,I187129,I187111,I187132,I187114,I187108,I187108,I187117,I187126,I187123,I187111,I187178,I187181,I187184,I187187,I187190,I187193,I187196,I187199,I187202,I2224,I2231);
PAT_16 I_2619 (I187184,I187187,I187196,I187190,I187202,I187178,I187199,I187193,I187181,I187181,I187178,I187248,I187251,I187254,I187257,I187260,I187263,I187266,I187269,I187272,I187275,I2224,I2231);
PAT_13 I_2620 (I187260,I187251,I187248,I187254,I187263,I187272,I187269,I187266,I187257,I187248,I187275,I187321,I187324,I187327,I187330,I187333,I187336,I187339,I187342,I187345,I2224,I2231);
PAT_11 I_2621 (I187321,I187333,I187336,I187327,I187324,I187345,I187324,I187342,I187330,I187321,I187339,I187391,I187394,I187397,I187400,I187403,I187406,I187409,I187412,I187415,I187418,I2224,I2231);
PAT_5 I_2622 (I187412,I187391,I187418,I187406,I187403,I187415,I187397,I187391,I187409,I187394,I187400,I187464,I187467,I187470,I187473,I187476,I187479,I187482,I187485,I187488,I187491,I2224,I2231);
PAT_13 I_2623 (I187470,I187479,I187464,I187467,I187488,I187473,I187485,I187464,I187482,I187491,I187476,I187537,I187540,I187543,I187546,I187549,I187552,I187555,I187558,I187561,I2224,I2231);
PAT_14 I_2624 (I187540,I187555,I187543,I187552,I187546,I187537,I187549,I187558,I187537,I187561,I187540,I187607,I187610,I187613,I187616,I187619,I187622,I187625,I187628,I187631,I2224,I2231);
PAT_17 I_2625 (I187622,I187610,I187631,I187607,I187628,I187616,I187613,I187625,I187619,I187610,I187607,I187677,I187680,I187683,I187686,I187689,I187692,I187695,I187698,I187701,I187704,I2224,I2231);
PAT_13 I_2626 (I187695,I187698,I187683,I187677,I187689,I187701,I187680,I187692,I187677,I187704,I187686,I187750,I187753,I187756,I187759,I187762,I187765,I187768,I187771,I187774,I2224,I2231);
PAT_4 I_2627 (I187759,I187762,I187774,I187756,I187771,I187768,I187753,I187765,I187753,I187750,I187750,I187820,I187823,I187826,I187829,I187832,I187835,I187838,I187841,I187844,I2224,I2231);
PAT_17 I_2628 (I187832,I187829,I187841,I187835,I187820,I187838,I187844,I187823,I187826,I187823,I187820,I187890,I187893,I187896,I187899,I187902,I187905,I187908,I187911,I187914,I187917,I2224,I2231);
PAT_4 I_2629 (I187899,I187890,I187908,I187905,I187917,I187914,I187893,I187890,I187896,I187902,I187911,I187963,I187966,I187969,I187972,I187975,I187978,I187981,I187984,I187987,I2224,I2231);
PAT_9 I_2630 (I187984,I187966,I187969,I187978,I187981,I187963,I187972,I187966,I187987,I187963,I187975,I188033,I188036,I188039,I188042,I188045,I188048,I188051,I188054,I188057,I2224,I2231);
PAT_15 I_2631 (I188045,I188054,I188057,I188036,I188051,I188039,I188042,I188033,I188048,I188033,I188036,I188103,I188106,I188109,I188112,I188115,I188118,I188121,I188124,I188127,I2224,I2231);
PAT_14 I_2632 (I188106,I188106,I188127,I188103,I188109,I188103,I188118,I188115,I188124,I188112,I188121,I188173,I188176,I188179,I188182,I188185,I188188,I188191,I188194,I188197,I2224,I2231);
PAT_9 I_2633 (I188182,I188194,I188173,I188191,I188176,I188179,I188197,I188176,I188185,I188173,I188188,I188243,I188246,I188249,I188252,I188255,I188258,I188261,I188264,I188267,I2224,I2231);
PAT_14 I_2634 (I188252,I188243,I188267,I188249,I188246,I188243,I188258,I188264,I188255,I188246,I188261,I188313,I188316,I188319,I188322,I188325,I188328,I188331,I188334,I188337,I2224,I2231);
PAT_12 I_2635 (I188322,I188328,I188313,I188337,I188316,I188316,I188331,I188313,I188334,I188325,I188319,I188383,I188386,I188389,I188392,I188395,I188398,I188401,I188404,I2224,I2231);
PAT_15 I_2636 (I188404,I188386,I188383,I188383,I188398,I188401,I188395,I188386,I188389,I188392,I188389,I188450,I188453,I188456,I188459,I188462,I188465,I188468,I188471,I188474,I2224,I2231);
PAT_11 I_2637 (I188471,I188453,I188450,I188465,I188456,I188450,I188468,I188474,I188462,I188453,I188459,I188520,I188523,I188526,I188529,I188532,I188535,I188538,I188541,I188544,I188547,I2224,I2231);
PAT_8 I_2638 (I188529,I188535,I188538,I188544,I188541,I188532,I188520,I188520,I188547,I188523,I188526,I188593,I188596,I188599,I188602,I188605,I188608,I188611,I188614,I188617,I2224,I2231);
PAT_9 I_2639 (I188596,I188605,I188596,I188593,I188608,I188599,I188614,I188602,I188611,I188593,I188617,I188663,I188666,I188669,I188672,I188675,I188678,I188681,I188684,I188687,I2224,I2231);
PAT_4 I_2640 (I188663,I188687,I188681,I188669,I188666,I188684,I188666,I188663,I188678,I188672,I188675,I188733,I188736,I188739,I188742,I188745,I188748,I188751,I188754,I188757,I2224,I2231);
PAT_17 I_2641 (I188745,I188742,I188754,I188748,I188733,I188751,I188757,I188736,I188739,I188736,I188733,I188803,I188806,I188809,I188812,I188815,I188818,I188821,I188824,I188827,I188830,I2224,I2231);
PAT_14 I_2642 (I188806,I188821,I188803,I188827,I188812,I188818,I188803,I188824,I188809,I188830,I188815,I188876,I188879,I188882,I188885,I188888,I188891,I188894,I188897,I188900,I2224,I2231);
PAT_10 I_2643 (I188879,I188876,I188882,I188900,I188897,I188891,I188879,I188894,I188876,I188888,I188885,I188946,I188949,I188952,I188955,I188958,I188961,I188964,I188967,I2224,I2231);
PAT_11 I_2644 (I188955,I188958,I188967,I188961,I188964,I188946,I188946,I188952,I188949,I188949,I188952,I189013,I189016,I189019,I189022,I189025,I189028,I189031,I189034,I189037,I189040,I2224,I2231);
PAT_6 I_2645 (I189013,I189040,I189028,I189037,I189031,I189025,I189016,I189034,I189022,I189019,I189013,I189086,I189089,I189092,I189095,I189098,I189101,I189104,I189107,I189110,I189113,I2224,I2231);
PAT_8 I_2646 (I189095,I189101,I189092,I189104,I189086,I189089,I189107,I189086,I189113,I189110,I189098,I189159,I189162,I189165,I189168,I189171,I189174,I189177,I189180,I189183,I2224,I2231);
PAT_2 I_2647 (I189162,I189177,I189183,I189159,I189171,I189174,I189162,I189180,I189165,I189168,I189159,I189229,I189232,I189235,I189238,I189241,I189244,I189247,I189250,I189253,I2224,I2231);
PAT_14 I_2648 (I189235,I189238,I189253,I189244,I189229,I189232,I189247,I189241,I189229,I189250,I189232,I189299,I189302,I189305,I189308,I189311,I189314,I189317,I189320,I189323,I2224,I2231);
PAT_17 I_2649 (I189314,I189302,I189323,I189299,I189320,I189308,I189305,I189317,I189311,I189302,I189299,I189369,I189372,I189375,I189378,I189381,I189384,I189387,I189390,I189393,I189396,I2224,I2231);
PAT_4 I_2650 (I189378,I189369,I189387,I189384,I189396,I189393,I189372,I189369,I189375,I189381,I189390,I189442,I189445,I189448,I189451,I189454,I189457,I189460,I189463,I189466,I2224,I2231);
PAT_10 I_2651 (I189442,I189442,I189466,I189445,I189451,I189460,I189457,I189445,I189463,I189448,I189454,I189512,I189515,I189518,I189521,I189524,I189527,I189530,I189533,I2224,I2231);
PAT_4 I_2652 (I189527,I189524,I189515,I189533,I189512,I189515,I189521,I189518,I189530,I189512,I189518,I189579,I189582,I189585,I189588,I189591,I189594,I189597,I189600,I189603,I2224,I2231);
PAT_11 I_2653 (I189591,I189600,I189582,I189594,I189579,I189582,I189579,I189588,I189603,I189597,I189585,I189649,I189652,I189655,I189658,I189661,I189664,I189667,I189670,I189673,I189676,I2224,I2231);
PAT_10 I_2654 (I189664,I189670,I189661,I189655,I189673,I189658,I189676,I189667,I189649,I189652,I189649,I189722,I189725,I189728,I189731,I189734,I189737,I189740,I189743,I2224,I2231);
PAT_2 I_2655 (I189734,I189737,I189728,I189740,I189725,I189722,I189722,I189728,I189743,I189731,I189725,I189789,I189792,I189795,I189798,I189801,I189804,I189807,I189810,I189813,I2224,I2231);
PAT_5 I_2656 (I189810,I189789,I189789,I189801,I189798,I189807,I189795,I189804,I189813,I189792,I189792,I189859,I189862,I189865,I189868,I189871,I189874,I189877,I189880,I189883,I189886,I2224,I2231);
PAT_2 I_2657 (I189874,I189859,I189871,I189865,I189880,I189862,I189877,I189868,I189883,I189886,I189859,I189932,I189935,I189938,I189941,I189944,I189947,I189950,I189953,I189956,I2224,I2231);
PAT_9 I_2658 (I189947,I189956,I189932,I189938,I189941,I189950,I189935,I189944,I189953,I189935,I189932,I190002,I190005,I190008,I190011,I190014,I190017,I190020,I190023,I190026,I2224,I2231);
PAT_6 I_2659 (I190020,I190002,I190014,I190023,I190002,I190011,I190008,I190026,I190017,I190005,I190005,I190072,I190075,I190078,I190081,I190084,I190087,I190090,I190093,I190096,I190099,I2224,I2231);
PAT_4 I_2660 (I190072,I190087,I190075,I190078,I190081,I190072,I190099,I190090,I190093,I190084,I190096,I190145,I190148,I190151,I190154,I190157,I190160,I190163,I190166,I190169,I2224,I2231);
PAT_6 I_2661 (I190145,I190151,I190148,I190160,I190163,I190157,I190169,I190166,I190145,I190154,I190148,I190215,I190218,I190221,I190224,I190227,I190230,I190233,I190236,I190239,I190242,I2224,I2231);
PAT_5 I_2662 (I190236,I190215,I190221,I190224,I190230,I190233,I190215,I190239,I190218,I190227,I190242,I190288,I190291,I190294,I190297,I190300,I190303,I190306,I190309,I190312,I190315,I2224,I2231);
PAT_4 I_2663 (I190306,I190312,I190315,I190294,I190297,I190309,I190291,I190288,I190300,I190303,I190288,I190361,I190364,I190367,I190370,I190373,I190376,I190379,I190382,I190385,I2224,I2231);
PAT_7 I_2664 (I190376,I190370,I190367,I190361,I190373,I190379,I190364,I190364,I190382,I190385,I190361,I190431,I190434,I190437,I190440,I190443,I190446,I190449,I190452,I190455,I2224,I2231);
PAT_2 I_2665 (I190452,I190446,I190437,I190431,I190440,I190434,I190443,I190455,I190449,I190434,I190431,I190501,I190504,I190507,I190510,I190513,I190516,I190519,I190522,I190525,I2224,I2231);
PAT_1 I_2666 (I190513,I190501,I190507,I190510,I190501,I190516,I190525,I190504,I190519,I190504,I190522,I190571,I190574,I190577,I190580,I190583,I190586,I190589,I190592,I190595,I2224,I2231);
PAT_8 I_2667 (I190592,I190574,I190580,I190571,I190589,I190583,I190586,I190571,I190595,I190577,I190574,I190641,I190644,I190647,I190650,I190653,I190656,I190659,I190662,I190665,I2224,I2231);
PAT_5 I_2668 (I190647,I190665,I190641,I190662,I190650,I190653,I190644,I190641,I190644,I190656,I190659,I190711,I190714,I190717,I190720,I190723,I190726,I190729,I190732,I190735,I190738,I2224,I2231);
PAT_7 I_2669 (I190729,I190732,I190738,I190735,I190720,I190717,I190711,I190723,I190711,I190714,I190726,I190784,I190787,I190790,I190793,I190796,I190799,I190802,I190805,I190808,I2224,I2231);
PAT_6 I_2670 (I190784,I190802,I190784,I190793,I190799,I190787,I190805,I190790,I190808,I190787,I190796,I190854,I190857,I190860,I190863,I190866,I190869,I190872,I190875,I190878,I190881,I2224,I2231);
PAT_10 I_2671 (I190854,I190869,I190872,I190863,I190854,I190878,I190881,I190857,I190866,I190860,I190875,I190927,I190930,I190933,I190936,I190939,I190942,I190945,I190948,I2224,I2231);
PAT_12 I_2672 (I190933,I190927,I190927,I190939,I190942,I190930,I190930,I190945,I190948,I190933,I190936,I190994,I190997,I191000,I191003,I191006,I191009,I191012,I191015,I2224,I2231);
PAT_5 I_2673 (I191003,I191009,I191015,I191000,I191000,I190994,I191012,I190994,I190997,I190997,I191006,I191061,I191064,I191067,I191070,I191073,I191076,I191079,I191082,I191085,I191088,I2224,I2231);
PAT_2 I_2674 (I191076,I191061,I191073,I191067,I191082,I191064,I191079,I191070,I191085,I191088,I191061,I191134,I191137,I191140,I191143,I191146,I191149,I191152,I191155,I191158,I2224,I2231);
PAT_13 I_2675 (I191143,I191137,I191134,I191155,I191146,I191149,I191137,I191140,I191152,I191158,I191134,I191204,I191207,I191210,I191213,I191216,I191219,I191222,I191225,I191228,I2224,I2231);
PAT_4 I_2676 (I191213,I191216,I191228,I191210,I191225,I191222,I191207,I191219,I191207,I191204,I191204,I191274,I191277,I191280,I191283,I191286,I191289,I191292,I191295,I191298,I2224,I2231);
PAT_10 I_2677 (I191274,I191274,I191298,I191277,I191283,I191292,I191289,I191277,I191295,I191280,I191286,I191344,I191347,I191350,I191353,I191356,I191359,I191362,I191365,I2224,I2231);
PAT_9 I_2678 (I191356,I191344,I191347,I191350,I191344,I191350,I191353,I191347,I191365,I191359,I191362,I191411,I191414,I191417,I191420,I191423,I191426,I191429,I191432,I191435,I2224,I2231);
PAT_2 I_2679 (I191426,I191429,I191420,I191435,I191411,I191414,I191417,I191414,I191432,I191423,I191411,I191481,I191484,I191487,I191490,I191493,I191496,I191499,I191502,I191505,I2224,I2231);
PAT_11 I_2680 (I191484,I191496,I191481,I191493,I191490,I191502,I191499,I191484,I191505,I191487,I191481,I191551,I191554,I191557,I191560,I191563,I191566,I191569,I191572,I191575,I191578,I2224,I2231);
PAT_13 I_2681 (I191551,I191554,I191563,I191575,I191578,I191566,I191572,I191560,I191569,I191557,I191551,I191624,I191627,I191630,I191633,I191636,I191639,I191642,I191645,I191648,I2224,I2231);
PAT_5 I_2682 (I191636,I191627,I191633,I191645,I191627,I191648,I191630,I191639,I191624,I191624,I191642,I191694,I191697,I191700,I191703,I191706,I191709,I191712,I191715,I191718,I191721,I2224,I2231);
PAT_8 I_2683 (I191694,I191721,I191712,I191709,I191703,I191694,I191706,I191718,I191697,I191715,I191700,I191767,I191770,I191773,I191776,I191779,I191782,I191785,I191788,I191791,I2224,I2231);
PAT_2 I_2684 (I191770,I191785,I191791,I191767,I191779,I191782,I191770,I191788,I191773,I191776,I191767,I191837,I191840,I191843,I191846,I191849,I191852,I191855,I191858,I191861,I2224,I2231);
PAT_1 I_2685 (I191849,I191837,I191843,I191846,I191837,I191852,I191861,I191840,I191855,I191840,I191858,I191907,I191910,I191913,I191916,I191919,I191922,I191925,I191928,I191931,I2224,I2231);
PAT_2 I_2686 (I191907,I191913,I191907,I191922,I191910,I191910,I191916,I191919,I191925,I191931,I191928,I191977,I191980,I191983,I191986,I191989,I191992,I191995,I191998,I192001,I2224,I2231);
PAT_11 I_2687 (I191980,I191992,I191977,I191989,I191986,I191998,I191995,I191980,I192001,I191983,I191977,I192047,I192050,I192053,I192056,I192059,I192062,I192065,I192068,I192071,I192074,I2224,I2231);
PAT_13 I_2688 (I192047,I192050,I192059,I192071,I192074,I192062,I192068,I192056,I192065,I192053,I192047,I192120,I192123,I192126,I192129,I192132,I192135,I192138,I192141,I192144,I2224,I2231);
PAT_12 I_2689 (I192129,I192120,I192120,I192144,I192141,I192123,I192138,I192132,I192123,I192126,I192135,I192190,I192193,I192196,I192199,I192202,I192205,I192208,I192211,I2224,I2231);
PAT_10 I_2690 (I192190,I192211,I192202,I192205,I192196,I192193,I192190,I192208,I192196,I192199,I192193,I192257,I192260,I192263,I192266,I192269,I192272,I192275,I192278,I2224,I2231);
PAT_17 I_2691 (I192269,I192278,I192272,I192257,I192263,I192275,I192260,I192260,I192257,I192263,I192266,I192324,I192327,I192330,I192333,I192336,I192339,I192342,I192345,I192348,I192351,I2224,I2231);
PAT_4 I_2692 (I192333,I192324,I192342,I192339,I192351,I192348,I192327,I192324,I192330,I192336,I192345,I192397,I192400,I192403,I192406,I192409,I192412,I192415,I192418,I192421,I2224,I2231);
PAT_9 I_2693 (I192418,I192400,I192403,I192412,I192415,I192397,I192406,I192400,I192421,I192397,I192409,I192467,I192470,I192473,I192476,I192479,I192482,I192485,I192488,I192491,I2224,I2231);
PAT_17 I_2694 (I192470,I192476,I192491,I192482,I192485,I192473,I192467,I192479,I192467,I192470,I192488,I192537,I192540,I192543,I192546,I192549,I192552,I192555,I192558,I192561,I192564,I2224,I2231);
PAT_11 I_2695 (I192549,I192558,I192564,I192540,I192537,I192555,I192546,I192552,I192543,I192561,I192537,I192610,I192613,I192616,I192619,I192622,I192625,I192628,I192631,I192634,I192637,I2224,I2231);
PAT_12 I_2696 (I192619,I192634,I192616,I192613,I192622,I192625,I192631,I192610,I192628,I192637,I192610,I192683,I192686,I192689,I192692,I192695,I192698,I192701,I192704,I2224,I2231);
PAT_11 I_2697 (I192689,I192692,I192689,I192701,I192704,I192698,I192686,I192695,I192683,I192686,I192683,I192750,I192753,I192756,I192759,I192762,I192765,I192768,I192771,I192774,I192777,I2224,I2231);
PAT_13 I_2698 (I192750,I192753,I192762,I192774,I192777,I192765,I192771,I192759,I192768,I192756,I192750,I192823,I192826,I192829,I192832,I192835,I192838,I192841,I192844,I192847,I2224,I2231);
PAT_7 I_2699 (I192832,I192835,I192823,I192838,I192844,I192829,I192826,I192847,I192826,I192823,I192841,I192893,I192896,I192899,I192902,I192905,I192908,I192911,I192914,I192917,I2224,I2231);
PAT_9 I_2700 (I192914,I192902,I192911,I192917,I192899,I192905,I192896,I192908,I192893,I192893,I192896,I192963,I192966,I192969,I192972,I192975,I192978,I192981,I192984,I192987,I2224,I2231);
PAT_6 I_2701 (I192981,I192963,I192975,I192984,I192963,I192972,I192969,I192987,I192978,I192966,I192966,I193033,I193036,I193039,I193042,I193045,I193048,I193051,I193054,I193057,I193060,I2224,I2231);
PAT_1 I_2702 (I193060,I193051,I193039,I193042,I193054,I193045,I193048,I193033,I193036,I193033,I193057,I193106,I193109,I193112,I193115,I193118,I193121,I193124,I193127,I193130,I2224,I2231);
PAT_13 I_2703 (I193115,I193124,I193130,I193106,I193121,I193118,I193127,I193112,I193109,I193106,I193109,I193176,I193179,I193182,I193185,I193188,I193191,I193194,I193197,I193200,I2224,I2231);
PAT_2 I_2704 (I193194,I193188,I193185,I193191,I193176,I193200,I193179,I193197,I193176,I193182,I193179,I193246,I193249,I193252,I193255,I193258,I193261,I193264,I193267,I193270,I2224,I2231);
PAT_12 I_2705 (I193255,I193252,I193246,I193249,I193270,I193264,I193267,I193249,I193261,I193246,I193258,I193316,I193319,I193322,I193325,I193328,I193331,I193334,I193337,I2224,I2231);
PAT_5 I_2706 (I193325,I193331,I193337,I193322,I193322,I193316,I193334,I193316,I193319,I193319,I193328,I193383,I193386,I193389,I193392,I193395,I193398,I193401,I193404,I193407,I193410,I2224,I2231);
PAT_2 I_2707 (I193398,I193383,I193395,I193389,I193404,I193386,I193401,I193392,I193407,I193410,I193383,I193456,I193459,I193462,I193465,I193468,I193471,I193474,I193477,I193480,I2224,I2231);
PAT_14 I_2708 (I193462,I193465,I193480,I193471,I193456,I193459,I193474,I193468,I193456,I193477,I193459,I193526,I193529,I193532,I193535,I193538,I193541,I193544,I193547,I193550,I2224,I2231);
PAT_13 I_2709 (I193535,I193550,I193529,I193538,I193526,I193529,I193544,I193532,I193526,I193547,I193541,I193596,I193599,I193602,I193605,I193608,I193611,I193614,I193617,I193620,I2224,I2231);
PAT_9 I_2710 (I193617,I193599,I193599,I193596,I193620,I193602,I193605,I193596,I193608,I193614,I193611,I193666,I193669,I193672,I193675,I193678,I193681,I193684,I193687,I193690,I2224,I2231);
PAT_4 I_2711 (I193666,I193690,I193684,I193672,I193669,I193687,I193669,I193666,I193681,I193675,I193678,I193736,I193739,I193742,I193745,I193748,I193751,I193754,I193757,I193760,I2224,I2231);
PAT_10 I_2712 (I193736,I193736,I193760,I193739,I193745,I193754,I193751,I193739,I193757,I193742,I193748,I193806,I193809,I193812,I193815,I193818,I193821,I193824,I193827,I2224,I2231);
PAT_15 I_2713 (I193821,I193824,I193812,I193818,I193806,I193806,I193812,I193827,I193815,I193809,I193809,I193873,I193876,I193879,I193882,I193885,I193888,I193891,I193894,I193897,I2224,I2231);
PAT_9 I_2714 (I193873,I193894,I193882,I193876,I193888,I193876,I193891,I193897,I193879,I193873,I193885,I193943,I193946,I193949,I193952,I193955,I193958,I193961,I193964,I193967,I2224,I2231);
PAT_7 I_2715 (I193949,I193958,I193943,I193964,I193955,I193943,I193946,I193967,I193961,I193946,I193952,I194013,I194016,I194019,I194022,I194025,I194028,I194031,I194034,I194037,I2224,I2231);
PAT_6 I_2716 (I194013,I194031,I194013,I194022,I194028,I194016,I194034,I194019,I194037,I194016,I194025,I194083,I194086,I194089,I194092,I194095,I194098,I194101,I194104,I194107,I194110,I2224,I2231);
PAT_10 I_2717 (I194083,I194098,I194101,I194092,I194083,I194107,I194110,I194086,I194095,I194089,I194104,I194156,I194159,I194162,I194165,I194168,I194171,I194174,I194177,I2224,I2231);
PAT_6 I_2718 (I194177,I194171,I194165,I194159,I194156,I194162,I194156,I194162,I194159,I194168,I194174,I194223,I194226,I194229,I194232,I194235,I194238,I194241,I194244,I194247,I194250,I2224,I2231);
PAT_2 I_2719 (I194244,I194250,I194232,I194238,I194223,I194229,I194223,I194235,I194226,I194241,I194247,I194296,I194299,I194302,I194305,I194308,I194311,I194314,I194317,I194320,I2224,I2231);
PAT_12 I_2720 (I194305,I194302,I194296,I194299,I194320,I194314,I194317,I194299,I194311,I194296,I194308,I194366,I194369,I194372,I194375,I194378,I194381,I194384,I194387,I2224,I2231);
PAT_6 I_2721 (I194375,I194369,I194387,I194372,I194369,I194372,I194381,I194366,I194384,I194366,I194378,I194433,I194436,I194439,I194442,I194445,I194448,I194451,I194454,I194457,I194460,I2224,I2231);
PAT_8 I_2722 (I194442,I194448,I194439,I194451,I194433,I194436,I194454,I194433,I194460,I194457,I194445,I194506,I194509,I194512,I194515,I194518,I194521,I194524,I194527,I194530,I2224,I2231);
PAT_9 I_2723 (I194509,I194518,I194509,I194506,I194521,I194512,I194527,I194515,I194524,I194506,I194530,I194576,I194579,I194582,I194585,I194588,I194591,I194594,I194597,I194600,I2224,I2231);
PAT_10 I_2724 (I194597,I194594,I194582,I194579,I194600,I194585,I194591,I194579,I194576,I194576,I194588,I194646,I194649,I194652,I194655,I194658,I194661,I194664,I194667,I2224,I2231);
PAT_11 I_2725 (I194655,I194658,I194667,I194661,I194664,I194646,I194646,I194652,I194649,I194649,I194652,I194713,I194716,I194719,I194722,I194725,I194728,I194731,I194734,I194737,I194740,I2224,I2231);
PAT_9 I_2726 (I194719,I194731,I194722,I194734,I194713,I194716,I194725,I194713,I194728,I194737,I194740,I194786,I194789,I194792,I194795,I194798,I194801,I194804,I194807,I194810,I2224,I2231);
PAT_13 I_2727 (I194786,I194807,I194789,I194804,I194798,I194795,I194810,I194786,I194792,I194801,I194789,I194856,I194859,I194862,I194865,I194868,I194871,I194874,I194877,I194880,I2224,I2231);
PAT_11 I_2728 (I194856,I194868,I194871,I194862,I194859,I194880,I194859,I194877,I194865,I194856,I194874,I194926,I194929,I194932,I194935,I194938,I194941,I194944,I194947,I194950,I194953,I2224,I2231);
PAT_13 I_2729 (I194926,I194929,I194938,I194950,I194953,I194941,I194947,I194935,I194944,I194932,I194926,I194999,I195002,I195005,I195008,I195011,I195014,I195017,I195020,I195023,I2224,I2231);
PAT_9 I_2730 (I195020,I195002,I195002,I194999,I195023,I195005,I195008,I194999,I195011,I195017,I195014,I195069,I195072,I195075,I195078,I195081,I195084,I195087,I195090,I195093,I2224,I2231);
PAT_2 I_2731 (I195084,I195087,I195078,I195093,I195069,I195072,I195075,I195072,I195090,I195081,I195069,I195139,I195142,I195145,I195148,I195151,I195154,I195157,I195160,I195163,I2224,I2231);
PAT_10 I_2732 (I195139,I195157,I195154,I195142,I195145,I195160,I195151,I195139,I195148,I195163,I195142,I195209,I195212,I195215,I195218,I195221,I195224,I195227,I195230,I2224,I2231);
PAT_9 I_2733 (I195221,I195209,I195212,I195215,I195209,I195215,I195218,I195212,I195230,I195224,I195227,I195276,I195279,I195282,I195285,I195288,I195291,I195294,I195297,I195300,I2224,I2231);
PAT_4 I_2734 (I195276,I195300,I195294,I195282,I195279,I195297,I195279,I195276,I195291,I195285,I195288,I195346,I195349,I195352,I195355,I195358,I195361,I195364,I195367,I195370,I2224,I2231);
PAT_9 I_2735 (I195367,I195349,I195352,I195361,I195364,I195346,I195355,I195349,I195370,I195346,I195358,I195416,I195419,I195422,I195425,I195428,I195431,I195434,I195437,I195440,I2224,I2231);
PAT_5 I_2736 (I195437,I195416,I195431,I195416,I195422,I195425,I195419,I195419,I195434,I195428,I195440,I195486,I195489,I195492,I195495,I195498,I195501,I195504,I195507,I195510,I195513,I2224,I2231);
PAT_4 I_2737 (I195504,I195510,I195513,I195492,I195495,I195507,I195489,I195486,I195498,I195501,I195486,I195559,I195562,I195565,I195568,I195571,I195574,I195577,I195580,I195583,I2224,I2231);
PAT_9 I_2738 (I195580,I195562,I195565,I195574,I195577,I195559,I195568,I195562,I195583,I195559,I195571,I195629,I195632,I195635,I195638,I195641,I195644,I195647,I195650,I195653,I2224,I2231);
PAT_7 I_2739 (I195635,I195644,I195629,I195650,I195641,I195629,I195632,I195653,I195647,I195632,I195638,I195699,I195702,I195705,I195708,I195711,I195714,I195717,I195720,I195723,I2224,I2231);
PAT_2 I_2740 (I195720,I195714,I195705,I195699,I195708,I195702,I195711,I195723,I195717,I195702,I195699,I195769,I195772,I195775,I195778,I195781,I195784,I195787,I195790,I195793,I2224,I2231);
PAT_15 I_2741 (I195772,I195784,I195790,I195793,I195775,I195787,I195769,I195778,I195769,I195781,I195772,I195839,I195842,I195845,I195848,I195851,I195854,I195857,I195860,I195863,I2224,I2231);
PAT_8 I_2742 (I195860,I195839,I195839,I195848,I195845,I195842,I195857,I195854,I195842,I195863,I195851,I195909,I195912,I195915,I195918,I195921,I195924,I195927,I195930,I195933,I2224,I2231);
PAT_13 I_2743 (I195921,I195930,I195912,I195933,I195915,I195909,I195909,I195918,I195927,I195924,I195912,I195979,I195982,I195985,I195988,I195991,I195994,I195997,I196000,I196003,I2224,I2231);
PAT_17 I_2744 (I196003,I195991,I196000,I195997,I195988,I195979,I195982,I195985,I195979,I195994,I195982,I196049,I196052,I196055,I196058,I196061,I196064,I196067,I196070,I196073,I196076,I2224,I2231);
PAT_5 I_2745 (I196061,I196055,I196052,I196073,I196058,I196064,I196067,I196049,I196049,I196070,I196076,I196122,I196125,I196128,I196131,I196134,I196137,I196140,I196143,I196146,I196149,I2224,I2231);
PAT_1 I_2746 (I196137,I196125,I196143,I196122,I196128,I196122,I196131,I196146,I196140,I196149,I196134,I196195,I196198,I196201,I196204,I196207,I196210,I196213,I196216,I196219,I2224,I2231);
PAT_9 I_2747 (I196210,I196216,I196201,I196219,I196198,I196213,I196198,I196204,I196195,I196207,I196195,I196265,I196268,I196271,I196274,I196277,I196280,I196283,I196286,I196289,I2224,I2231);
PAT_3 I_2748 (I196289,I196268,I196271,I196283,I196274,I196268,I196277,I196265,I196286,I196265,I196280,I196335,I196338,I196341,I196344,I196347,I196350,I196353,I196356,I196359,I196362,I2224,I2231);
PAT_6 I_2749 (I196362,I196350,I196344,I196335,I196335,I196353,I196341,I196356,I196359,I196347,I196338,I196408,I196411,I196414,I196417,I196420,I196423,I196426,I196429,I196432,I196435,I2224,I2231);
PAT_17 I_2750 (I196420,I196423,I196429,I196417,I196411,I196432,I196426,I196408,I196435,I196414,I196408,I196481,I196484,I196487,I196490,I196493,I196496,I196499,I196502,I196505,I196508,I2224,I2231);
PAT_6 I_2751 (I196481,I196499,I196487,I196490,I196496,I196481,I196493,I196484,I196505,I196508,I196502,I196554,I196557,I196560,I196563,I196566,I196569,I196572,I196575,I196578,I196581,I2224,I2231);
PAT_1 I_2752 (I196581,I196572,I196560,I196563,I196575,I196566,I196569,I196554,I196557,I196554,I196578,I196627,I196630,I196633,I196636,I196639,I196642,I196645,I196648,I196651,I2224,I2231);
PAT_2 I_2753 (I196627,I196633,I196627,I196642,I196630,I196630,I196636,I196639,I196645,I196651,I196648,I196697,I196700,I196703,I196706,I196709,I196712,I196715,I196718,I196721,I2224,I2231);
PAT_13 I_2754 (I196706,I196700,I196697,I196718,I196709,I196712,I196700,I196703,I196715,I196721,I196697,I196767,I196770,I196773,I196776,I196779,I196782,I196785,I196788,I196791,I2224,I2231);
PAT_2 I_2755 (I196785,I196779,I196776,I196782,I196767,I196791,I196770,I196788,I196767,I196773,I196770,I196837,I196840,I196843,I196846,I196849,I196852,I196855,I196858,I196861,I2224,I2231);
PAT_11 I_2756 (I196840,I196852,I196837,I196849,I196846,I196858,I196855,I196840,I196861,I196843,I196837,I196907,I196910,I196913,I196916,I196919,I196922,I196925,I196928,I196931,I196934,I2224,I2231);
PAT_14 I_2757 (I196928,I196916,I196910,I196931,I196922,I196925,I196913,I196934,I196919,I196907,I196907,I196980,I196983,I196986,I196989,I196992,I196995,I196998,I197001,I197004,I2224,I2231);
PAT_13 I_2758 (I196989,I197004,I196983,I196992,I196980,I196983,I196998,I196986,I196980,I197001,I196995,I197050,I197053,I197056,I197059,I197062,I197065,I197068,I197071,I197074,I2224,I2231);
PAT_5 I_2759 (I197062,I197053,I197059,I197071,I197053,I197074,I197056,I197065,I197050,I197050,I197068,I197120,I197123,I197126,I197129,I197132,I197135,I197138,I197141,I197144,I197147,I2224,I2231);
PAT_17 I_2760 (I197147,I197123,I197126,I197129,I197120,I197132,I197120,I197144,I197138,I197135,I197141,I197193,I197196,I197199,I197202,I197205,I197208,I197211,I197214,I197217,I197220,I2224,I2231);
PAT_5 I_2761 (I197205,I197199,I197196,I197217,I197202,I197208,I197211,I197193,I197193,I197214,I197220,I197266,I197269,I197272,I197275,I197278,I197281,I197284,I197287,I197290,I197293,I2224,I2231);
PAT_13 I_2762 (I197272,I197281,I197266,I197269,I197290,I197275,I197287,I197266,I197284,I197293,I197278,I197339,I197342,I197345,I197348,I197351,I197354,I197357,I197360,I197363,I2224,I2231);
PAT_12 I_2763 (I197348,I197339,I197339,I197363,I197360,I197342,I197357,I197351,I197342,I197345,I197354,I197409,I197412,I197415,I197418,I197421,I197424,I197427,I197430,I2224,I2231);
PAT_11 I_2764 (I197415,I197418,I197415,I197427,I197430,I197424,I197412,I197421,I197409,I197412,I197409,I197476,I197479,I197482,I197485,I197488,I197491,I197494,I197497,I197500,I197503,I2224,I2231);
PAT_1 I_2765 (I197491,I197482,I197485,I197476,I197497,I197494,I197479,I197476,I197503,I197500,I197488,I197549,I197552,I197555,I197558,I197561,I197564,I197567,I197570,I197573,I2224,I2231);
PAT_3 I_2766 (I197558,I197552,I197552,I197555,I197567,I197570,I197573,I197561,I197549,I197549,I197564,I197619,I197622,I197625,I197628,I197631,I197634,I197637,I197640,I197643,I197646,I2224,I2231);
PAT_13 I_2767 (I197640,I197628,I197646,I197625,I197631,I197634,I197622,I197637,I197619,I197619,I197643,I197692,I197695,I197698,I197701,I197704,I197707,I197710,I197713,I197716,I2224,I2231);
PAT_4 I_2768 (I197701,I197704,I197716,I197698,I197713,I197710,I197695,I197707,I197695,I197692,I197692,I197762,I197765,I197768,I197771,I197774,I197777,I197780,I197783,I197786,I2224,I2231);
PAT_14 I_2769 (I197765,I197780,I197777,I197762,I197774,I197765,I197762,I197768,I197783,I197771,I197786,I197832,I197835,I197838,I197841,I197844,I197847,I197850,I197853,I197856,I2224,I2231);
PAT_7 I_2770 (I197832,I197841,I197838,I197844,I197835,I197856,I197835,I197853,I197850,I197847,I197832,I197902,I197905,I197908,I197911,I197914,I197917,I197920,I197923,I197926,I2224,I2231);
PAT_9 I_2771 (I197923,I197911,I197920,I197926,I197908,I197914,I197905,I197917,I197902,I197902,I197905,I197972,I197975,I197978,I197981,I197984,I197987,I197990,I197993,I197996,I2224,I2231);
PAT_10 I_2772 (I197993,I197990,I197978,I197975,I197996,I197981,I197987,I197975,I197972,I197972,I197984,I198042,I198045,I198048,I198051,I198054,I198057,I198060,I198063,I2224,I2231);
PAT_5 I_2773 (I198063,I198042,I198051,I198045,I198060,I198057,I198048,I198048,I198042,I198045,I198054,I198109,I198112,I198115,I198118,I198121,I198124,I198127,I198130,I198133,I198136,I2224,I2231);
PAT_11 I_2774 (I198121,I198118,I198112,I198130,I198133,I198109,I198127,I198124,I198136,I198115,I198109,I198182,I198185,I198188,I198191,I198194,I198197,I198200,I198203,I198206,I198209,I2224,I2231);
PAT_4 I_2775 (I198188,I198209,I198182,I198200,I198191,I198182,I198203,I198185,I198194,I198206,I198197,I198255,I198258,I198261,I198264,I198267,I198270,I198273,I198276,I198279,I2224,I2231);
PAT_9 I_2776 (I198276,I198258,I198261,I198270,I198273,I198255,I198264,I198258,I198279,I198255,I198267,I198325,I198328,I198331,I198334,I198337,I198340,I198343,I198346,I198349,I2224,I2231);
PAT_15 I_2777 (I198337,I198346,I198349,I198328,I198343,I198331,I198334,I198325,I198340,I198325,I198328,I198395,I198398,I198401,I198404,I198407,I198410,I198413,I198416,I198419,I2224,I2231);
PAT_2 I_2778 (I198398,I198398,I198401,I198407,I198395,I198395,I198404,I198419,I198413,I198416,I198410,I198465,I198468,I198471,I198474,I198477,I198480,I198483,I198486,I198489,I2224,I2231);
PAT_5 I_2779 (I198486,I198465,I198465,I198477,I198474,I198483,I198471,I198480,I198489,I198468,I198468,I198535,I198538,I198541,I198544,I198547,I198550,I198553,I198556,I198559,I198562,I2224,I2231);
PAT_8 I_2780 (I198535,I198562,I198553,I198550,I198544,I198535,I198547,I198559,I198538,I198556,I198541,I198608,I198611,I198614,I198617,I198620,I198623,I198626,I198629,I198632,I2224,I2231);
PAT_3 I_2781 (I198629,I198620,I198611,I198617,I198614,I198626,I198611,I198632,I198608,I198623,I198608,I198678,I198681,I198684,I198687,I198690,I198693,I198696,I198699,I198702,I198705,I2224,I2231);
PAT_10 I_2782 (I198687,I198690,I198681,I198705,I198678,I198693,I198699,I198678,I198696,I198702,I198684,I198751,I198754,I198757,I198760,I198763,I198766,I198769,I198772,I2224,I2231);
PAT_13 I_2783 (I198757,I198763,I198757,I198754,I198769,I198772,I198751,I198751,I198766,I198754,I198760,I198818,I198821,I198824,I198827,I198830,I198833,I198836,I198839,I198842,I2224,I2231);
PAT_5 I_2784 (I198830,I198821,I198827,I198839,I198821,I198842,I198824,I198833,I198818,I198818,I198836,I198888,I198891,I198894,I198897,I198900,I198903,I198906,I198909,I198912,I198915,I2224,I2231);
PAT_10 I_2785 (I198912,I198915,I198894,I198900,I198903,I198909,I198891,I198888,I198888,I198897,I198906,I198961,I198964,I198967,I198970,I198973,I198976,I198979,I198982,I2224,I2231);
PAT_2 I_2786 (I198973,I198976,I198967,I198979,I198964,I198961,I198961,I198967,I198982,I198970,I198964,I199028,I199031,I199034,I199037,I199040,I199043,I199046,I199049,I199052,I2224,I2231);
PAT_17 I_2787 (I199028,I199028,I199040,I199031,I199034,I199046,I199043,I199052,I199031,I199037,I199049,I199098,I199101,I199104,I199107,I199110,I199113,I199116,I199119,I199122,I199125,I2224,I2231);
PAT_8 I_2788 (I199107,I199119,I199125,I199116,I199101,I199110,I199113,I199122,I199104,I199098,I199098,I199171,I199174,I199177,I199180,I199183,I199186,I199189,I199192,I199195,I2224,I2231);
PAT_6 I_2789 (I199174,I199171,I199177,I199189,I199186,I199180,I199183,I199171,I199192,I199174,I199195,I199241,I199244,I199247,I199250,I199253,I199256,I199259,I199262,I199265,I199268,I2224,I2231);
endmodule


