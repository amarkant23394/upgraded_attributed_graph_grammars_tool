module test_I16551(I13162,I1477,I14503,I1470,I16551);
input I13162,I1477,I14503,I1470;
output I16551;
wire I14667,I13189,I14901,I14537,I14808,I14344,I14520,I16534,I16240,I14370,I13174,I14650,I14335,I14715;
and I_0(I14667,I14650,I13189);
DFFARX1 I_1(I1470,,,I13189,);
DFFARX1 I_2(I14808,I1470,I14370,,,I14901,);
DFFARX1 I_3(I14520,I1470,I14370,,,I14537,);
DFFARX1 I_4(I13162,I1470,I14370,,,I14808,);
nand I_5(I14344,I14537,I14715);
and I_6(I14520,I14503,I13174);
DFFARX1 I_7(I14335,I1470,I16240,,,I16534,);
not I_8(I16240,I1477);
not I_9(I14370,I1477);
DFFARX1 I_10(I1470,,,I13174,);
DFFARX1 I_11(I1470,I14370,,,I14650,);
and I_12(I16551,I16534,I14344);
and I_13(I14335,I14808,I14901);
not I_14(I14715,I14667);
endmodule


