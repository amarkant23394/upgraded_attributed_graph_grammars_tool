module test_I11947(I10154,I10038,I1477,I1470,I11947);
input I10154,I10038,I1477,I1470;
output I11947;
wire I10219,I12425,I10020,I12106,I12524,I12442,I10052,I11973,I10287;
nand I_0(I11947,I12106,I12524);
DFFARX1 I_1(I1470,I10052,,,I10219,);
DFFARX1 I_2(I10038,I1470,I11973,,,I12425,);
DFFARX1 I_3(I10287,I1470,I10052,,,I10020,);
not I_4(I12106,I10020);
not I_5(I12524,I12442);
not I_6(I12442,I12425);
not I_7(I10052,I1477);
not I_8(I11973,I1477);
and I_9(I10287,I10219,I10154);
endmodule


