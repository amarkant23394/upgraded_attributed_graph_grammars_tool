module test_final(IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2,n4_7_l_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
nor I_0(N1371_0_r_2,n32_2,n35_2);
nor I_1(N1508_0_r_2,n32_2,n55_2);
not I_2(N1372_1_r_2,n54_2);
nor I_3(N1508_1_r_2,n59_2,n54_2);
nor I_4(N6147_2_r_2,n42_2,n43_2);
nor I_5(N1507_6_r_2,n40_2,n53_2);
nor I_6(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_7(n4_7_r_2,blif_clk_net_8_r_10,n11_10,G42_7_r_2,);
nor I_8(n_572_7_r_2,n36_2,n37_2);
or I_9(n_573_7_r_2,n34_2,n35_2);
nor I_10(n_549_7_r_2,n40_2,n41_2);
nand I_11(n_569_7_r_2,n38_2,n39_2);
nor I_12(n_452_7_r_2,n59_2,n35_2);
nor I_13(n4_7_l_2,G18_7_l_2,IN_1_7_l_2);
DFFARX1 I_14(n4_7_l_2,blif_clk_net_8_r_10,n11_10,n59_2,);
not I_15(n33_2,n59_2);
and I_16(N3_8_l_2,IN_6_8_l_2,n49_2);
DFFARX1 I_17(N3_8_l_2,blif_clk_net_8_r_10,n11_10,n32_internal_2,);
not I_18(n32_2,n32_internal_2);
nor I_19(n4_7_r_2,n59_2,n36_2);
not I_20(n34_2,n39_2);
nor I_21(n35_2,IN_1_8_l_2,IN_3_8_l_2);
nor I_22(n36_2,G18_7_l_2,IN_5_7_l_2);
or I_23(n37_2,IN_9_7_l_2,IN_10_7_l_2);
not I_24(n38_2,n40_2);
nand I_25(n39_2,n45_2,n57_2);
nor I_26(n40_2,IN_3_1_l_2,n47_2);
nor I_27(n41_2,n32_2,n36_2);
not I_28(n42_2,n53_2);
nand I_29(n43_2,n44_2,n45_2);
nand I_30(n44_2,n38_2,n46_2);
not I_31(n45_2,IN_10_7_l_2);
nand I_32(n46_2,n47_2,n48_2);
nand I_33(n47_2,IN_1_1_l_2,IN_2_1_l_2);
or I_34(n48_2,G15_7_l_2,IN_7_7_l_2);
nand I_35(n49_2,IN_2_8_l_2,IN_3_8_l_2);
nand I_36(n50_2,n51_2,n52_2);
not I_37(n51_2,n47_2);
nand I_38(n52_2,n38_2,n53_2);
nor I_39(n53_2,IN_5_7_l_2,IN_9_7_l_2);
nand I_40(n54_2,n42_2,n56_2);
nor I_41(n55_2,n34_2,n56_2);
nor I_42(n56_2,G15_7_l_2,IN_7_7_l_2);
nand I_43(n57_2,IN_4_7_l_2,n58_2);
not I_44(n58_2,G15_7_l_2);
nor I_45(N1371_0_r_10,n37_10,n38_10);
nor I_46(N1508_0_r_10,n37_10,n58_10);
nand I_47(N6147_2_r_10,n39_10,n40_10);
not I_48(N6147_3_r_10,n39_10);
nor I_49(N1372_4_r_10,n46_10,n49_10);
nor I_50(N1508_4_r_10,n51_10,n52_10);
nor I_51(N1507_6_r_10,n49_10,n60_10);
nor I_52(N1508_6_r_10,n49_10,n50_10);
nor I_53(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_54(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_55(N6147_9_r_10,n36_10,n37_10);
nor I_56(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_57(I_BUFF_1_9_r_10,n48_10);
nor I_58(N3_8_r_10,n44_10,n47_10);
not I_59(n11_10,blif_reset_net_8_r_10);
not I_60(n35_10,n49_10);
nor I_61(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_62(n37_10,N1372_1_r_2);
not I_63(n38_10,n46_10);
nand I_64(n39_10,n43_10,n44_10);
nand I_65(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_66(n41_10,n42_10,N1372_1_r_2);
not I_67(n42_10,n44_10);
nor I_68(n43_10,n45_10,N1372_1_r_2);
nand I_69(n44_10,n54_10,n_573_7_r_2);
nor I_70(n45_10,n59_10,N6147_2_r_2);
nand I_71(n46_10,n61_10,N1508_1_r_2);
nor I_72(n47_10,n46_10,n48_10);
nand I_73(n48_10,n62_10,n63_10);
nand I_74(n49_10,n56_10,N1507_6_r_2);
not I_75(n50_10,n45_10);
nor I_76(n51_10,n42_10,n53_10);
not I_77(n52_10,N1372_4_r_10);
nor I_78(n53_10,n48_10,n50_10);
and I_79(n54_10,n55_10,n_452_7_r_2);
nand I_80(n55_10,n56_10,n57_10);
nand I_81(n56_10,N1371_0_r_2,n_569_7_r_2);
not I_82(n57_10,N1507_6_r_2);
nor I_83(n58_10,n35_10,n45_10);
nor I_84(n59_10,n_572_7_r_2,N1371_0_r_2);
nor I_85(n60_10,n37_10,n46_10);
or I_86(n61_10,n_572_7_r_2,N1371_0_r_2);
nor I_87(n62_10,G42_7_r_2,n_549_7_r_2);
or I_88(n63_10,n64_10,N1508_0_r_2);
nor I_89(n64_10,N1508_0_r_2,N1508_6_r_2);
endmodule


