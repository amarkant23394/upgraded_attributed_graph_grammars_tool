module test_I4000(I1415,I1351,I1447,I1477,I3028,I1470,I1407,I4000);
input I1415,I1351,I1447,I1477,I3028,I1470,I1407;
output I4000;
wire I2721,I2878,I2759,I3045,I3155,I3076,I2861,I2724,I2980,I2776;
nand I_0(I2721,I2980,I2878);
not I_1(I2878,I2861);
not I_2(I2759,I1477);
and I_3(I3045,I2861,I3028);
or I_4(I3155,I3076,I3045);
nand I_5(I4000,I2721,I2724);
DFFARX1 I_6(I1447,I1470,I2759,,,I3076,);
not I_7(I2861,I1351);
DFFARX1 I_8(I3155,I1470,I2759,,,I2724,);
nand I_9(I2980,I2776,I1415);
not I_10(I2776,I1407);
endmodule


