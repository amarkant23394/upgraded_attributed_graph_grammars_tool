module Benchmark_testing25000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2595,I2602,I17674,I17665,I17662,I17668,I17656,I17650,I17671,I17659,I17653,I58627,I58603,I58615,I58609,I58624,I58618,I58612,I58606,I58621,I62197,I62173,I62185,I62179,I62194,I62188,I62182,I62176,I62191,I90107,I90131,I90113,I90116,I90104,I90122,I90125,I90110,I90119,I90128,I108025,I108049,I108031,I108034,I108022,I108040,I108043,I108028,I108037,I108046,I154099,I154096,I154081,I154093,I154087,I154075,I154084,I154090,I154078,I244618,I244621,I244612,I244603,I244606,I244615,I244600,I244609,I251996,I251999,I251990,I251981,I251984,I251993,I251978,I251987,I266738,I266741,I266717,I266729,I266744,I266732,I266726,I266720,I266723,I266735,I289348,I289330,I289333,I289342,I289345,I289339,I289327,I289336,I319483,I319471,I319492,I319468,I319489,I319480,I319486,I319477,I319474,I347542,I347521,I347524,I347539,I347536,I347533,I347530,I347518,I347527,I350806,I350785,I350788,I350803,I350800,I350797,I350794,I350782,I350791,I370047,I370050,I370035,I370038,I370032,I370029,I370053,I370044,I370026,I370041);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2595,I2602;
output I17674,I17665,I17662,I17668,I17656,I17650,I17671,I17659,I17653,I58627,I58603,I58615,I58609,I58624,I58618,I58612,I58606,I58621,I62197,I62173,I62185,I62179,I62194,I62188,I62182,I62176,I62191,I90107,I90131,I90113,I90116,I90104,I90122,I90125,I90110,I90119,I90128,I108025,I108049,I108031,I108034,I108022,I108040,I108043,I108028,I108037,I108046,I154099,I154096,I154081,I154093,I154087,I154075,I154084,I154090,I154078,I244618,I244621,I244612,I244603,I244606,I244615,I244600,I244609,I251996,I251999,I251990,I251981,I251984,I251993,I251978,I251987,I266738,I266741,I266717,I266729,I266744,I266732,I266726,I266720,I266723,I266735,I289348,I289330,I289333,I289342,I289345,I289339,I289327,I289336,I319483,I319471,I319492,I319468,I319489,I319480,I319486,I319477,I319474,I347542,I347521,I347524,I347539,I347536,I347533,I347530,I347518,I347527,I350806,I350785,I350788,I350803,I350800,I350797,I350794,I350782,I350791,I370047,I370050,I370035,I370038,I370032,I370029,I370053,I370044,I370026,I370041;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2595,I2602,I2634,I185940,I2660,I2668,I185919,I2685,I2626,I185928,I2725,I2733,I2750,I185934,I2767,I185931,I2784,I2801,I2605,I2832,I2849,I2866,I185922,I185916,I2608,I2897,I2914,I185937,I2931,I2948,I2965,I2982,I2617,I3013,I185925,I3030,I3047,I2623,I3078,I2620,I3109,I3135,I3143,I3160,I2614,I2611,I3229,I339701,I3255,I3263,I3280,I3221,I339716,I3320,I3328,I3345,I339713,I3362,I339722,I3379,I3396,I3200,I3427,I3444,I3461,I339710,I339719,I3203,I3492,I3509,I339707,I3526,I339698,I3543,I3560,I3577,I3212,I3608,I339704,I3625,I3642,I3218,I3673,I3215,I3704,I3730,I3738,I3755,I3209,I3206,I3824,I346454,I3850,I3858,I346442,I3875,I3816,I346430,I3915,I3923,I3940,I3957,I346436,I3974,I3991,I3795,I4022,I4039,I4056,I346433,I346448,I3798,I4087,I4104,I346439,I4121,I346451,I4138,I4155,I4172,I3807,I4203,I346445,I4220,I4237,I3813,I4268,I3810,I4299,I4325,I4333,I4350,I3804,I3801,I4419,I100659,I4445,I4453,I100650,I4470,I4411,I100653,I4510,I4518,I4535,I100647,I4552,I100656,I4569,I4586,I4390,I4617,I4634,I4651,I100644,I100662,I4393,I4682,I4699,I4716,I100668,I4733,I4750,I4767,I4402,I4798,I100665,I4815,I4832,I4408,I4863,I4405,I4894,I100671,I4920,I4928,I4945,I4399,I4396,I5014,I82741,I5040,I5048,I82732,I5065,I5006,I82735,I5105,I5113,I5130,I82729,I5147,I82738,I5164,I5181,I4985,I5212,I5229,I5246,I82726,I82744,I4988,I5277,I5294,I5311,I82750,I5328,I5345,I5362,I4997,I5393,I82747,I5410,I5427,I5003,I5458,I5000,I5489,I82753,I5515,I5523,I5540,I4994,I4991,I5609,I335655,I5635,I5643,I5660,I5601,I335670,I5700,I5708,I5725,I335667,I5742,I335676,I5759,I5776,I5580,I5807,I5824,I5841,I335664,I335673,I5583,I5872,I5889,I335661,I5906,I335652,I5923,I5940,I5957,I5592,I5988,I335658,I6005,I6022,I5598,I6053,I5595,I6084,I6110,I6118,I6135,I5589,I5586,I6204,I154670,I6230,I6238,I154691,I6255,I6196,I154688,I6295,I6303,I6320,I6337,I154682,I6354,I6371,I6175,I6402,I6419,I6436,I154685,I154694,I6178,I6467,I6484,I154673,I6501,I154676,I6518,I6535,I6552,I6187,I6583,I6600,I6617,I6193,I6648,I6190,I6679,I154679,I6705,I6713,I6730,I6184,I6181,I6799,I360237,I6825,I6833,I360243,I6850,I6791,I360246,I6890,I6898,I6915,I360234,I6932,I360252,I6949,I6966,I6770,I6997,I7014,I7031,I360249,I360258,I6773,I7062,I7079,I7096,I360255,I7113,I7130,I7147,I6782,I7178,I360240,I7195,I7212,I6788,I7243,I6785,I7274,I7300,I7308,I7325,I6779,I6776,I7394,I342591,I7420,I7428,I7445,I7386,I342606,I7485,I7493,I7510,I342603,I7527,I342612,I7544,I7561,I7365,I7592,I7609,I7626,I342600,I342609,I7368,I7657,I7674,I342597,I7691,I342588,I7708,I7725,I7742,I7377,I7773,I342594,I7790,I7807,I7383,I7838,I7380,I7869,I7895,I7903,I7920,I7374,I7371,I7989,I277720,I8015,I8023,I277711,I8040,I7981,I277714,I8080,I8088,I8105,I277726,I8122,I277705,I8139,I8156,I7960,I8187,I8204,I8221,I277717,I277723,I7963,I8252,I8269,I277708,I8286,I277699,I8303,I8320,I8337,I7972,I8368,I8385,I8402,I7978,I8433,I7975,I8464,I277702,I8490,I8498,I8515,I7969,I7966,I8584,I217730,I8610,I8618,I217709,I8635,I8576,I217718,I8675,I8683,I8700,I217724,I8717,I217721,I8734,I8751,I8555,I8782,I8799,I8816,I217712,I217706,I8558,I8847,I8864,I217727,I8881,I8898,I8915,I8932,I8567,I8963,I217715,I8980,I8997,I8573,I9028,I8570,I9059,I9085,I9093,I9110,I8564,I8561,I9179,I32945,I9205,I9213,I32936,I9230,I9171,I32957,I9270,I9278,I9295,I32933,I9312,I9329,I9346,I9150,I9377,I9394,I9411,I32942,I9153,I9442,I9459,I32954,I9476,I32951,I9493,I9510,I9527,I9162,I9558,I32948,I9575,I9592,I9168,I9623,I9165,I9654,I32939,I9680,I9688,I9705,I9159,I9156,I9777,I201528,I9803,I9820,I9828,I9845,I201543,I201546,I9862,I201525,I9888,I9769,I9760,I201531,I9933,I9941,I201537,I9958,I9757,I9998,I10006,I9763,I9751,I10051,I201540,I201522,I10068,I201534,I10094,I10102,I9745,I10133,I10150,I10167,I10184,I10201,I9766,I10232,I9754,I9748,I10304,I289894,I10330,I10347,I10355,I10372,I289888,I289909,I10389,I10415,I10296,I10287,I289891,I10460,I10468,I289900,I10485,I10284,I10525,I10533,I10290,I10278,I10578,I289906,I10595,I289897,I10621,I10629,I10272,I10660,I10677,I289903,I10694,I10711,I10728,I10293,I10759,I10281,I10275,I10831,I268679,I10857,I10874,I10882,I10899,I268655,I268682,I10916,I268667,I10942,I10823,I10814,I268673,I10987,I10995,I268658,I11012,I10811,I268676,I11052,I11060,I10817,I10805,I11105,I268661,I268664,I11122,I11148,I11156,I10799,I11187,I11204,I268670,I11221,I11238,I11255,I10820,I11286,I10808,I10802,I11358,I31882,I11384,I11401,I11409,I11426,I31897,I11443,I31900,I11469,I11350,I11341,I31894,I11514,I11522,I31903,I11539,I11338,I31879,I11579,I11587,I11344,I11332,I11632,I31885,I11649,I31888,I11675,I11683,I11326,I11714,I11731,I31891,I11748,I11765,I11782,I11347,I11813,I11335,I11329,I11885,I225226,I11911,I11928,I11936,I11953,I225241,I225244,I11970,I225223,I11996,I11877,I11868,I225229,I12041,I12049,I225235,I12066,I11865,I12106,I12114,I11871,I11859,I12159,I225238,I225220,I12176,I225232,I12202,I12210,I11853,I12241,I12258,I12275,I12292,I12309,I11874,I12340,I11862,I11856,I12412,I194014,I12438,I12455,I12463,I12480,I194029,I194032,I12497,I194011,I12523,I12404,I12395,I194017,I12568,I12576,I194023,I12593,I12392,I12633,I12641,I12398,I12386,I12686,I194026,I194008,I12703,I194020,I12729,I12737,I12380,I12768,I12785,I12802,I12819,I12836,I12401,I12867,I12389,I12383,I12939,I74674,I12965,I12982,I12990,I13007,I74692,I74677,I13024,I74680,I13050,I12931,I12922,I74668,I13095,I13103,I74671,I13120,I12919,I74683,I13160,I13168,I12925,I12913,I13213,I74689,I74686,I13230,I13256,I13264,I12907,I13295,I13312,I13329,I13346,I13363,I12928,I13394,I12916,I12910,I13466,I309666,I13492,I13509,I13517,I13534,I309654,I309645,I13551,I309642,I13577,I13458,I13449,I309648,I13622,I13630,I309660,I13647,I13446,I309657,I13687,I13695,I13452,I13440,I13740,I309651,I13757,I309663,I13783,I13791,I13434,I13822,I13839,I13856,I13873,I13890,I13455,I13921,I13443,I13437,I13993,I189390,I14019,I14036,I14044,I14061,I189405,I189408,I14078,I189387,I14104,I13985,I13976,I189393,I14149,I14157,I189399,I14174,I13973,I14214,I14222,I13979,I13967,I14267,I189402,I189384,I14284,I189396,I14310,I14318,I13961,I14349,I14366,I14383,I14400,I14417,I13982,I14448,I13970,I13964,I14520,I14546,I14563,I14571,I14588,I14605,I14631,I14512,I14503,I14676,I14684,I14701,I14500,I14741,I14749,I14506,I14494,I14794,I14811,I14837,I14845,I14488,I14876,I14893,I14910,I14927,I14944,I14509,I14975,I14497,I14491,I15047,I15073,I15090,I15098,I15115,I15132,I15158,I15039,I15030,I15203,I15211,I15228,I15027,I15268,I15276,I15033,I15021,I15321,I15338,I15364,I15372,I15015,I15403,I15420,I15437,I15454,I15471,I15036,I15502,I15024,I15018,I15574,I327006,I15600,I15617,I15625,I15642,I326994,I326985,I15659,I326982,I15685,I15566,I15557,I326988,I15730,I15738,I327000,I15755,I15554,I326997,I15795,I15803,I15560,I15548,I15848,I326991,I15865,I327003,I15891,I15899,I15542,I15930,I15947,I15964,I15981,I15998,I15563,I16029,I15551,I15545,I16101,I30828,I16127,I16144,I16152,I16169,I30843,I16186,I30846,I16212,I16093,I16084,I30840,I16257,I16265,I30849,I16282,I16081,I30825,I16322,I16330,I16087,I16075,I16375,I30831,I16392,I30834,I16418,I16426,I16069,I16457,I16474,I30837,I16491,I16508,I16525,I16090,I16556,I16078,I16072,I16628,I99617,I16654,I16671,I16679,I16696,I99614,I99608,I16713,I99602,I16739,I16620,I16611,I99590,I16784,I16792,I99599,I16809,I16608,I99596,I16849,I16857,I16614,I16602,I16902,I99593,I99611,I16919,I16945,I16953,I16596,I16984,I17001,I99605,I17018,I17035,I17052,I16617,I17083,I16605,I16599,I17155,I280307,I17181,I17198,I17206,I17223,I280283,I280310,I17240,I280295,I17266,I17147,I17138,I280301,I17311,I17319,I280286,I17336,I17135,I280304,I17376,I17384,I17141,I17129,I17429,I280289,I280292,I17446,I17472,I17480,I17123,I17511,I17528,I280298,I17545,I17562,I17579,I17144,I17610,I17132,I17126,I17682,I165123,I17708,I17725,I17733,I17750,I165108,I165126,I17767,I165120,I17793,I165117,I17838,I17846,I17863,I165111,I17903,I17911,I17956,I165132,I165114,I17973,I165129,I17999,I18007,I18038,I18055,I18072,I18089,I18106,I18137,I18209,I127929,I18235,I18252,I18260,I18277,I127932,I18294,I127953,I18320,I18201,I18192,I127941,I18365,I18373,I127944,I18390,I18189,I127950,I18430,I18438,I18195,I18183,I18483,I127947,I127935,I18500,I127938,I18526,I18534,I18177,I18565,I18582,I127956,I18599,I18616,I18633,I18198,I18664,I18186,I18180,I18736,I160499,I18762,I18779,I18787,I18804,I160484,I160502,I18821,I160496,I18847,I18728,I18719,I160493,I18892,I18900,I18917,I18716,I160487,I18957,I18965,I18722,I18710,I19010,I160508,I160490,I19027,I160505,I19053,I19061,I18704,I19092,I19109,I19126,I19143,I19160,I18725,I19191,I18713,I18707,I19263,I390783,I19289,I19306,I19314,I19331,I390786,I390792,I19348,I390801,I19374,I19255,I19246,I390804,I19419,I19427,I390795,I19444,I19243,I19484,I19492,I19249,I19237,I19537,I390810,I390789,I19554,I390798,I19580,I19588,I19231,I19619,I19636,I390807,I19653,I19670,I19687,I19252,I19718,I19240,I19234,I19790,I291577,I19816,I19833,I19841,I19858,I291571,I291592,I19875,I19901,I19782,I19773,I291574,I19946,I19954,I291583,I19971,I19770,I20011,I20019,I19776,I19764,I20064,I291589,I20081,I291580,I20107,I20115,I19758,I20146,I20163,I291586,I20180,I20197,I20214,I19779,I20245,I19767,I19761,I20317,I359671,I20343,I20360,I20368,I20385,I359674,I359668,I20402,I359677,I20428,I20309,I20300,I359665,I20473,I20481,I359680,I20498,I20297,I359656,I20538,I20546,I20303,I20291,I20591,I359659,I20608,I20634,I20642,I20285,I20673,I20690,I359662,I20707,I20724,I20741,I20306,I20772,I20294,I20288,I20844,I288059,I20870,I20887,I20895,I20912,I288035,I288062,I20929,I288047,I20955,I20836,I20827,I288053,I21000,I21008,I288038,I21025,I20824,I288056,I21065,I21073,I20830,I20818,I21118,I288041,I288044,I21135,I21161,I21169,I20812,I21200,I21217,I288050,I21234,I21251,I21268,I20833,I21299,I20821,I20815,I21371,I35044,I21397,I21414,I21422,I21439,I35059,I21456,I35062,I21482,I21363,I21354,I35056,I21527,I21535,I35065,I21552,I21351,I35041,I21592,I21600,I21357,I21345,I21645,I35047,I21662,I35050,I21688,I21696,I21339,I21727,I21744,I35053,I21761,I21778,I21795,I21360,I21826,I21348,I21342,I21898,I108576,I21924,I21941,I21949,I21966,I108573,I108567,I21983,I108561,I22009,I21890,I21881,I108549,I22054,I22062,I108558,I22079,I21878,I108555,I22119,I22127,I21884,I21872,I22172,I108552,I108570,I22189,I22215,I22223,I21866,I22254,I22271,I108564,I22288,I22305,I22322,I21887,I22353,I21875,I21869,I22425,I293260,I22451,I22468,I22476,I22493,I293254,I293275,I22510,I22536,I22417,I22408,I293257,I22581,I22589,I293266,I22606,I22405,I22646,I22654,I22411,I22399,I22699,I293272,I22716,I293263,I22742,I22750,I22393,I22781,I22798,I293269,I22815,I22832,I22849,I22414,I22880,I22402,I22396,I22952,I368928,I22978,I22995,I23003,I23020,I368919,I368925,I23037,I368904,I23063,I22944,I22935,I368922,I23108,I23116,I23133,I22932,I368916,I23173,I23181,I22938,I22926,I23226,I368910,I368931,I23243,I368913,I23269,I23277,I22920,I23308,I23325,I368907,I23342,I23359,I23376,I22941,I23407,I22929,I22923,I23479,I138827,I23505,I23513,I23530,I138821,I138812,I23547,I138833,I23573,I138815,I23590,I23598,I138809,I23615,I23447,I23646,I23663,I23459,I23703,I23468,I23725,I138836,I138818,I23742,I138824,I23768,I23785,I23471,I23807,I23456,I23838,I138830,I23855,I23872,I23889,I23465,I23920,I23453,I23462,I23450,I24006,I273832,I24032,I24040,I24057,I273850,I273844,I24074,I273823,I24100,I273841,I24117,I24125,I273826,I24142,I23974,I24173,I24190,I23986,I273838,I24230,I23995,I24252,I273847,I273835,I24269,I273829,I24295,I24312,I23998,I24334,I23983,I24365,I24382,I24399,I24416,I23992,I24447,I23980,I23989,I23977,I24533,I178411,I24559,I24567,I24584,I178423,I178408,I24601,I178402,I24627,I178417,I24644,I24652,I178405,I24669,I24501,I24700,I24717,I24513,I178414,I24757,I24522,I24779,I178420,I178426,I24796,I24822,I24839,I24525,I24861,I24510,I24892,I24909,I24926,I24943,I24519,I24974,I24507,I24516,I24504,I25060,I113319,I25086,I25094,I25111,I113301,I113316,I25128,I113292,I25154,I113295,I25171,I25179,I113310,I25196,I25028,I25227,I25244,I25040,I113313,I25284,I25049,I25306,I113304,I25323,I113298,I25349,I25366,I25052,I25388,I25037,I25419,I113307,I25436,I25453,I25470,I25046,I25501,I25034,I25043,I25031,I25587,I99090,I25613,I25621,I25638,I99072,I99087,I25655,I99063,I25681,I99066,I25698,I25706,I99081,I25723,I25555,I25754,I25771,I25567,I99084,I25811,I25576,I25833,I99075,I25850,I99069,I25876,I25893,I25579,I25915,I25564,I25946,I99078,I25963,I25980,I25997,I25573,I26028,I25561,I25570,I25558,I26114,I56830,I26140,I26148,I26165,I56824,I56818,I26182,I56839,I26208,I56836,I26225,I26233,I56833,I26250,I26082,I26281,I26298,I26094,I26338,I26103,I26360,I56821,I26377,I56842,I26403,I26420,I26106,I26442,I26091,I26473,I56827,I26490,I26507,I26524,I26100,I26555,I26088,I26097,I26085,I26641,I83807,I26667,I26675,I26692,I83789,I83804,I26709,I83780,I26735,I83783,I26752,I26760,I83798,I26777,I26609,I26808,I26825,I26621,I83801,I26865,I26630,I26887,I83792,I26904,I83786,I26930,I26947,I26633,I26969,I26618,I27000,I83795,I27017,I27034,I27051,I26627,I27082,I26615,I26624,I26612,I27168,I222342,I27194,I27202,I27219,I222333,I222351,I27236,I222330,I27262,I27279,I27287,I222336,I27304,I27136,I27335,I27352,I27148,I27392,I27157,I27414,I222348,I222339,I27431,I222354,I27457,I27474,I27160,I27496,I27145,I27527,I222345,I27544,I27561,I27578,I27154,I27609,I27142,I27151,I27139,I27695,I49690,I27721,I27729,I27746,I49684,I49678,I27763,I49699,I27789,I49696,I27806,I27814,I49693,I27831,I27663,I27862,I27879,I27675,I27919,I27684,I27941,I49681,I27958,I49702,I27984,I28001,I27687,I28023,I27672,I28054,I49687,I28071,I28088,I28105,I27681,I28136,I27669,I27678,I27666,I28222,I385440,I28248,I28256,I28273,I385434,I385455,I28290,I385431,I28316,I385452,I28333,I28341,I385449,I28358,I28190,I28389,I28406,I28202,I385437,I28446,I28211,I28468,I385446,I385443,I28485,I385428,I28511,I28528,I28214,I28550,I28199,I28581,I28598,I28615,I28632,I28208,I28663,I28196,I28205,I28193,I28749,I199222,I28775,I28783,I28800,I199213,I199231,I28817,I199210,I28843,I28860,I28868,I199216,I28885,I28717,I28916,I28933,I28729,I28973,I28738,I28995,I199228,I199219,I29012,I199234,I29038,I29055,I28741,I29077,I28726,I29108,I199225,I29125,I29142,I29159,I28735,I29190,I28723,I28732,I28720,I29276,I276416,I29302,I29310,I29327,I276434,I276428,I29344,I276407,I29370,I276425,I29387,I29395,I276410,I29412,I29244,I29443,I29460,I29256,I276422,I29500,I29265,I29522,I276431,I276419,I29539,I276413,I29565,I29582,I29268,I29604,I29253,I29635,I29652,I29669,I29686,I29262,I29717,I29250,I29259,I29247,I29803,I60400,I29829,I29837,I29854,I60394,I60388,I29871,I60409,I29897,I60406,I29914,I29922,I60403,I29939,I29771,I29970,I29987,I29783,I30027,I29792,I30049,I60391,I30066,I60412,I30092,I30109,I29795,I30131,I29780,I30162,I60397,I30179,I30196,I30213,I29789,I30244,I29777,I29786,I29774,I30330,I299989,I30356,I30364,I30381,I299986,I299992,I30398,I30424,I30441,I30449,I30466,I30298,I30497,I30514,I30310,I299995,I30554,I30319,I30576,I299998,I300007,I30593,I300001,I30619,I30636,I30322,I30658,I30307,I30689,I300004,I30706,I30723,I30740,I30316,I30771,I30304,I30313,I30301,I30857,I326410,I30883,I30891,I30908,I326425,I326404,I30925,I326407,I30951,I326428,I30968,I30976,I30993,I31024,I31041,I31081,I31103,I326416,I326413,I31120,I326419,I31146,I31163,I31185,I31216,I326422,I31233,I31250,I31267,I31298,I31384,I131211,I31410,I31418,I31435,I131205,I131196,I31452,I131217,I31478,I131199,I31495,I31503,I131193,I31520,I31352,I31551,I31568,I31364,I31608,I31373,I31630,I131220,I131202,I31647,I131208,I31673,I31690,I31376,I31712,I31361,I31743,I131214,I31760,I31777,I31794,I31370,I31825,I31358,I31367,I31355,I31911,I88023,I31937,I31945,I31962,I88005,I88020,I31979,I87996,I32005,I87999,I32022,I32030,I88014,I32047,I32078,I32095,I88017,I32135,I32157,I88008,I32174,I88002,I32200,I32217,I32239,I32270,I88011,I32287,I32304,I32321,I32352,I32438,I302794,I32464,I32472,I32489,I302791,I302797,I32506,I32532,I32549,I32557,I32574,I32406,I32605,I32622,I32418,I302800,I32662,I32427,I32684,I302803,I302812,I32701,I302806,I32727,I32744,I32430,I32766,I32415,I32797,I302809,I32814,I32831,I32848,I32424,I32879,I32412,I32421,I32409,I32965,I94347,I32991,I32999,I33016,I94329,I94344,I33033,I94320,I33059,I94323,I33076,I33084,I94338,I33101,I33132,I33149,I94341,I33189,I33211,I94332,I33228,I94326,I33254,I33271,I33293,I33324,I94335,I33341,I33358,I33375,I33406,I33492,I236704,I33518,I33526,I33543,I236701,I236716,I33560,I236698,I33586,I236695,I33603,I33611,I33628,I33460,I33659,I33676,I33472,I33716,I33481,I33738,I236710,I33755,I236713,I33781,I33798,I33484,I33820,I33469,I33851,I236707,I33868,I33885,I33902,I33478,I33933,I33466,I33475,I33463,I34019,I372945,I34045,I34053,I34070,I372939,I372960,I34087,I372936,I34113,I372957,I34130,I34138,I372954,I34155,I33987,I34186,I34203,I33999,I372942,I34243,I34008,I34265,I372951,I372948,I34282,I372933,I34308,I34325,I34011,I34347,I33996,I34378,I34395,I34412,I34429,I34005,I34460,I33993,I34002,I33990,I34546,I133931,I34572,I34580,I34597,I133925,I133916,I34614,I133937,I34640,I133919,I34657,I34665,I133913,I34682,I34514,I34713,I34730,I34526,I34770,I34535,I34792,I133940,I133922,I34809,I133928,I34835,I34852,I34538,I34874,I34523,I34905,I133934,I34922,I34939,I34956,I34532,I34987,I34520,I34529,I34517,I35073,I325832,I35099,I35107,I35124,I325847,I325826,I35141,I325829,I35167,I325850,I35184,I35192,I35209,I35240,I35257,I35297,I35319,I325838,I325835,I35336,I325841,I35362,I35379,I35401,I35432,I325844,I35449,I35466,I35483,I35514,I35600,I369465,I35626,I35634,I35651,I369471,I369489,I35668,I369486,I35694,I369483,I35711,I35719,I369477,I35736,I35568,I35767,I35784,I35580,I35824,I35589,I35846,I369480,I369468,I35863,I369492,I35889,I35906,I35592,I35928,I35577,I35959,I369474,I35976,I35993,I36010,I35586,I36041,I35574,I35583,I35571,I36127,I299428,I36153,I36161,I36178,I299425,I299431,I36195,I36221,I36238,I36246,I36263,I36095,I36294,I36311,I36107,I299434,I36351,I36116,I36373,I299437,I299446,I36390,I299440,I36416,I36433,I36119,I36455,I36104,I36486,I299443,I36503,I36520,I36537,I36113,I36568,I36101,I36110,I36098,I36654,I159337,I36680,I36688,I36705,I159349,I159334,I36722,I159328,I36748,I159343,I36765,I36773,I159331,I36790,I36622,I36821,I36838,I36634,I159340,I36878,I36643,I36900,I159346,I159352,I36917,I36943,I36960,I36646,I36982,I36631,I37013,I37030,I37047,I37064,I36640,I37095,I36628,I36637,I36625,I37181,I126315,I37207,I37215,I37232,I126309,I126300,I37249,I126321,I37275,I126303,I37292,I37300,I126297,I37317,I37149,I37348,I37365,I37161,I37405,I37170,I37427,I126324,I126306,I37444,I126312,I37470,I37487,I37173,I37509,I37158,I37540,I126318,I37557,I37574,I37591,I37167,I37622,I37155,I37164,I37152,I37708,I356228,I37734,I37742,I37759,I356222,I356243,I37776,I356234,I37802,I356225,I37819,I37827,I356237,I37844,I37676,I37875,I37892,I37688,I37932,I37697,I37954,I356246,I356231,I37971,I37997,I38014,I37700,I38036,I37685,I38067,I356240,I38084,I38101,I38118,I37694,I38149,I37682,I37691,I37679,I38235,I346980,I38261,I38269,I38286,I346974,I346995,I38303,I346986,I38329,I346977,I38346,I38354,I346989,I38371,I38203,I38402,I38419,I38215,I38459,I38224,I38481,I346998,I346983,I38498,I38524,I38541,I38227,I38563,I38212,I38594,I346992,I38611,I38628,I38645,I38221,I38676,I38209,I38218,I38206,I38762,I233542,I38788,I38796,I38813,I233539,I233554,I38830,I233536,I38856,I233533,I38873,I38881,I38898,I38730,I38929,I38946,I38742,I38986,I38751,I39008,I233548,I39025,I233551,I39051,I39068,I38754,I39090,I38739,I39121,I233545,I39138,I39155,I39172,I38748,I39203,I38736,I38745,I38733,I39289,I129035,I39315,I39323,I39340,I129029,I129020,I39357,I129041,I39383,I129023,I39400,I39408,I129017,I39425,I39257,I39456,I39473,I39269,I39513,I39278,I39535,I129044,I129026,I39552,I129032,I39578,I39595,I39281,I39617,I39266,I39648,I129038,I39665,I39682,I39699,I39275,I39730,I39263,I39272,I39260,I39816,I78845,I39842,I39850,I39867,I78839,I78833,I39884,I78854,I39910,I78851,I39927,I39935,I78848,I39952,I39784,I39983,I40000,I39796,I40040,I39805,I40062,I78836,I40079,I78857,I40105,I40122,I39808,I40144,I39793,I40175,I78842,I40192,I40209,I40226,I39802,I40257,I39790,I39799,I39787,I40343,I344804,I40369,I40377,I40394,I344798,I344819,I40411,I344810,I40437,I344801,I40454,I40462,I344813,I40479,I40311,I40510,I40527,I40323,I40567,I40332,I40589,I344822,I344807,I40606,I40632,I40649,I40335,I40671,I40320,I40702,I344816,I40719,I40736,I40753,I40329,I40784,I40317,I40326,I40314,I40870,I355140,I40896,I40904,I40921,I355134,I355155,I40938,I355146,I40964,I355137,I40981,I40989,I355149,I41006,I40838,I41037,I41054,I40850,I41094,I40859,I41116,I355158,I355143,I41133,I41159,I41176,I40862,I41198,I40847,I41229,I355152,I41246,I41263,I41280,I40856,I41311,I40844,I40853,I40841,I41397,I331034,I41423,I41431,I41448,I331049,I331028,I41465,I331031,I41491,I331052,I41508,I41516,I41533,I41365,I41564,I41581,I41377,I41621,I41386,I41643,I331040,I331037,I41660,I331043,I41686,I41703,I41389,I41725,I41374,I41756,I331046,I41773,I41790,I41807,I41383,I41838,I41371,I41380,I41368,I41924,I41950,I41958,I41975,I41992,I42018,I42035,I42043,I42060,I41892,I42091,I42108,I41904,I42148,I41913,I42170,I42187,I42213,I42230,I41916,I42252,I41901,I42283,I42300,I42317,I42334,I41910,I42365,I41898,I41907,I41895,I42451,I341438,I42477,I42485,I42502,I341453,I341432,I42519,I341435,I42545,I341456,I42562,I42570,I42587,I42419,I42618,I42635,I42431,I42675,I42440,I42697,I341444,I341441,I42714,I341447,I42740,I42757,I42443,I42779,I42428,I42810,I341450,I42827,I42844,I42861,I42437,I42892,I42425,I42434,I42422,I42978,I303916,I43004,I43012,I43029,I303913,I303919,I43046,I43072,I43089,I43097,I43114,I42946,I43145,I43162,I42958,I303922,I43202,I42967,I43224,I303925,I303934,I43241,I303928,I43267,I43284,I42970,I43306,I42955,I43337,I303931,I43354,I43371,I43388,I42964,I43419,I42952,I42961,I42949,I43505,I285460,I43531,I43539,I43556,I285478,I285472,I43573,I285451,I43599,I285469,I43616,I43624,I285454,I43641,I43473,I43672,I43689,I43485,I285466,I43729,I43494,I43751,I285475,I285463,I43768,I285457,I43794,I43811,I43497,I43833,I43482,I43864,I43881,I43898,I43915,I43491,I43946,I43479,I43488,I43476,I44032,I195754,I44058,I44066,I44083,I195745,I195763,I44100,I195742,I44126,I44143,I44151,I195748,I44168,I44000,I44199,I44216,I44012,I44256,I44021,I44278,I195760,I195751,I44295,I195766,I44321,I44338,I44024,I44360,I44009,I44391,I195757,I44408,I44425,I44442,I44018,I44473,I44006,I44015,I44003,I44559,I44585,I44593,I44610,I44627,I44653,I44670,I44678,I44695,I44527,I44726,I44743,I44539,I44783,I44548,I44805,I44822,I44848,I44865,I44551,I44887,I44536,I44918,I44935,I44952,I44969,I44545,I45000,I44533,I44542,I44530,I45086,I45112,I45120,I45137,I45154,I45180,I45197,I45205,I45222,I45054,I45253,I45270,I45066,I45310,I45075,I45332,I45349,I45375,I45392,I45078,I45414,I45063,I45445,I45462,I45479,I45496,I45072,I45527,I45060,I45069,I45057,I45613,I318318,I45639,I45647,I45664,I318333,I318312,I45681,I318315,I45707,I318336,I45724,I45732,I45749,I45581,I45780,I45797,I45593,I45837,I45602,I45859,I318324,I318321,I45876,I318327,I45902,I45919,I45605,I45941,I45590,I45972,I318330,I45989,I46006,I46023,I45599,I46054,I45587,I45596,I45584,I46143,I298873,I46169,I46177,I298867,I46203,I46211,I46228,I298885,I46245,I46120,I46276,I298870,I46114,I46307,I298876,I46324,I46341,I298864,I298882,I46358,I46375,I46392,I46129,I46126,I46132,I46451,I46468,I46485,I46511,I46111,I46542,I46550,I298879,I46135,I46581,I46598,I46615,I46117,I46646,I46663,I46108,I46123,I46738,I222908,I46764,I46772,I222929,I46798,I46806,I46823,I222920,I46840,I46715,I46871,I222917,I46709,I46902,I222926,I46919,I46936,I222911,I46953,I46970,I46987,I46724,I46721,I46727,I47046,I47063,I47080,I222932,I222914,I47106,I46706,I47137,I47145,I222923,I46730,I47176,I47193,I47210,I46712,I47241,I47258,I46703,I46718,I47333,I75287,I47359,I47367,I75281,I47393,I47401,I75266,I47418,I75275,I47435,I47310,I47466,I75263,I47304,I47497,I75269,I47514,I47531,I75272,I75284,I47548,I47565,I47582,I47319,I47316,I47322,I47641,I47658,I47675,I75278,I47701,I47301,I47732,I47740,I47325,I47771,I47788,I47805,I47307,I47836,I47853,I47298,I47313,I47928,I132849,I47954,I47962,I132843,I47988,I47996,I132840,I48013,I132831,I48030,I47905,I48061,I132834,I47899,I48092,I132837,I48109,I48126,I132825,I132852,I48143,I48160,I48177,I47914,I47911,I47917,I48236,I48253,I48270,I132828,I48296,I47896,I48327,I48335,I132846,I47920,I48366,I48383,I48400,I47902,I48431,I48448,I47893,I47908,I48520,I295501,I48546,I48563,I48512,I48585,I295510,I48611,I48619,I48636,I295504,I48653,I295498,I48670,I48687,I295513,I48704,I48721,I295507,I48738,I48488,I48769,I48786,I48803,I48820,I48500,I48494,I48865,I48509,I48503,I48910,I48927,I295519,I48944,I295516,I48961,I48987,I48995,I48497,I48491,I49049,I49057,I48506,I49115,I315422,I49141,I49158,I49107,I49180,I49206,I49214,I49231,I315425,I49248,I315437,I49265,I49282,I315443,I49299,I315434,I49316,I315440,I49333,I49083,I49364,I49381,I49398,I49415,I49095,I49089,I49460,I315431,I49104,I49098,I49505,I49522,I315428,I49539,I315446,I49556,I49582,I49590,I49092,I49086,I49644,I49652,I49101,I49710,I176105,I49736,I49753,I49775,I176096,I49801,I49809,I49826,I176114,I49843,I176111,I49860,I49877,I176090,I49894,I176093,I49911,I176102,I49928,I49959,I49976,I49993,I50010,I50055,I176108,I50100,I50117,I50134,I176099,I50151,I50177,I50185,I50239,I50247,I50305,I218874,I50331,I50348,I50297,I50370,I218871,I50396,I50404,I50421,I218877,I50438,I218862,I50455,I50472,I218865,I50489,I218886,I50506,I218883,I50523,I50273,I50554,I50571,I50588,I50605,I50285,I50279,I50650,I50294,I50288,I50695,I50712,I218868,I50729,I218880,I50746,I50772,I50780,I50282,I50276,I50834,I50842,I50291,I50900,I181304,I50926,I50943,I50892,I50965,I181301,I50991,I50999,I51016,I181307,I51033,I181292,I51050,I51067,I181295,I51084,I181316,I51101,I181313,I51118,I50868,I51149,I51166,I51183,I51200,I50880,I50874,I51245,I50889,I50883,I51290,I51307,I181298,I51324,I181310,I51341,I51367,I51375,I50877,I50871,I51429,I51437,I50886,I51495,I179573,I51521,I51538,I51487,I51560,I179564,I51586,I51594,I51611,I179582,I51628,I179579,I51645,I51662,I179558,I51679,I179561,I51696,I179570,I51713,I51463,I51744,I51761,I51778,I51795,I51475,I51469,I51840,I179576,I51484,I51478,I51885,I51902,I51919,I179567,I51936,I51962,I51970,I51472,I51466,I52024,I52032,I51481,I52090,I211938,I52116,I52133,I52082,I52155,I211935,I52181,I52189,I52206,I211941,I52223,I211926,I52240,I52257,I211929,I52274,I211950,I52291,I211947,I52308,I52058,I52339,I52356,I52373,I52390,I52070,I52064,I52435,I52079,I52073,I52480,I52497,I211932,I52514,I211944,I52531,I52557,I52565,I52067,I52061,I52619,I52627,I52076,I52685,I200378,I52711,I52728,I52677,I52750,I200375,I52776,I52784,I52801,I200381,I52818,I200366,I52835,I52852,I200369,I52869,I200390,I52886,I200387,I52903,I52653,I52934,I52951,I52968,I52985,I52665,I52659,I53030,I52674,I52668,I53075,I53092,I200372,I53109,I200384,I53126,I53152,I53160,I52662,I52656,I53214,I53222,I52671,I53280,I312532,I53306,I53323,I53272,I53345,I53371,I53379,I53396,I312535,I53413,I312547,I53430,I53447,I312553,I53464,I312544,I53481,I312550,I53498,I53248,I53529,I53546,I53563,I53580,I53260,I53254,I53625,I312541,I53269,I53263,I53670,I53687,I312538,I53704,I312556,I53721,I53747,I53755,I53257,I53251,I53809,I53817,I53266,I53875,I101698,I53901,I53918,I53867,I53940,I101713,I53966,I53974,I53991,I101710,I54008,I54025,I54042,I101707,I54059,I101722,I54076,I101719,I54093,I53843,I54124,I54141,I54158,I54175,I53855,I53849,I54220,I101716,I53864,I53858,I54265,I54282,I101704,I54299,I101725,I54316,I101701,I54342,I54350,I53852,I53846,I54404,I54412,I53861,I54470,I241971,I54496,I54513,I54462,I54535,I241965,I54561,I54569,I54586,I241983,I54603,I54620,I54637,I54654,I241977,I54671,I241968,I54688,I54438,I54719,I54736,I54753,I54770,I54450,I54444,I54815,I241980,I54459,I54453,I54860,I54877,I241986,I54894,I54911,I241974,I54937,I54945,I54447,I54441,I54999,I55007,I54456,I55065,I239863,I55091,I55108,I55057,I55130,I239857,I55156,I55164,I55181,I239875,I55198,I55215,I55232,I55249,I239869,I55266,I239860,I55283,I55033,I55314,I55331,I55348,I55365,I55045,I55039,I55410,I239872,I55054,I55048,I55455,I55472,I239878,I55489,I55506,I239866,I55532,I55540,I55042,I55036,I55594,I55602,I55051,I55660,I151112,I55686,I55703,I55652,I55725,I151106,I55751,I55759,I55776,I151121,I55793,I151118,I55810,I55827,I151109,I55844,I151100,I55861,I151103,I55878,I55628,I55909,I55926,I55943,I55960,I55640,I55634,I56005,I151124,I55649,I55643,I56050,I56067,I151115,I56084,I56101,I56127,I56135,I55637,I55631,I56189,I56197,I55646,I56255,I56281,I56298,I56247,I56320,I56346,I56354,I56371,I56388,I56405,I56422,I56439,I56456,I56473,I56223,I56504,I56521,I56538,I56555,I56235,I56229,I56600,I56244,I56238,I56645,I56662,I56679,I56696,I56722,I56730,I56232,I56226,I56784,I56792,I56241,I56850,I177839,I56876,I56893,I56915,I177830,I56941,I56949,I56966,I177848,I56983,I177845,I57000,I57017,I177824,I57034,I177827,I57051,I177836,I57068,I57099,I57116,I57133,I57150,I57195,I177842,I57240,I57257,I57274,I177833,I57291,I57317,I57325,I57379,I57387,I57445,I208470,I57471,I57488,I57437,I57510,I208467,I57536,I57544,I57561,I208473,I57578,I208458,I57595,I57612,I208461,I57629,I208482,I57646,I208479,I57663,I57413,I57694,I57711,I57728,I57745,I57425,I57419,I57790,I57434,I57428,I57835,I57852,I208464,I57869,I208476,I57886,I57912,I57920,I57422,I57416,I57974,I57982,I57431,I58040,I122513,I58066,I58083,I58032,I58105,I122501,I58131,I58139,I58156,I122510,I58173,I122507,I58190,I58207,I122498,I58224,I122504,I58241,I122489,I58258,I58008,I58289,I58306,I58323,I58340,I58020,I58014,I58385,I58029,I58023,I58430,I58447,I122495,I58464,I122492,I58481,I122516,I58507,I58515,I58017,I58011,I58569,I58577,I58026,I58635,I111711,I58661,I58678,I58700,I111726,I58726,I58734,I58751,I111723,I58768,I58785,I58802,I111720,I58819,I111735,I58836,I111732,I58853,I58884,I58901,I58918,I58935,I58980,I111729,I59025,I59042,I111717,I59059,I111738,I59076,I111714,I59102,I59110,I59164,I59172,I59230,I357347,I59256,I59273,I59222,I59295,I357359,I59321,I59329,I59346,I357353,I59363,I357365,I59380,I59397,I357350,I59414,I357362,I59431,I357344,I59448,I59198,I59479,I59496,I59513,I59530,I59210,I59204,I59575,I357356,I59219,I59213,I59620,I59637,I59654,I59671,I357368,I59697,I59705,I59207,I59201,I59759,I59767,I59216,I59825,I305596,I59851,I59868,I59817,I59890,I59916,I59924,I59941,I305599,I59958,I305611,I59975,I59992,I305617,I60009,I305608,I60026,I305614,I60043,I59793,I60074,I60091,I60108,I60125,I59805,I59799,I60170,I305605,I59814,I59808,I60215,I60232,I305602,I60249,I305620,I60266,I60292,I60300,I59802,I59796,I60354,I60362,I59811,I60420,I365439,I60446,I60463,I60485,I365451,I60511,I60519,I60536,I365445,I60553,I365457,I60570,I60587,I365442,I60604,I365454,I60621,I365436,I60638,I60669,I60686,I60703,I60720,I60765,I365448,I60810,I60827,I60844,I60861,I365460,I60887,I60895,I60949,I60957,I61015,I114346,I61041,I61058,I61007,I61080,I114361,I61106,I61114,I61131,I114358,I61148,I61165,I61182,I114355,I61199,I114370,I61216,I114367,I61233,I60983,I61264,I61281,I61298,I61315,I60995,I60989,I61360,I114364,I61004,I60998,I61405,I61422,I114352,I61439,I114373,I61456,I114349,I61482,I61490,I60992,I60986,I61544,I61552,I61001,I61610,I282882,I61636,I61653,I61602,I61675,I282891,I61701,I61709,I61726,I282879,I61743,I282870,I61760,I61777,I282876,I61794,I282894,I61811,I282867,I61828,I61578,I61859,I61876,I61893,I61910,I61590,I61584,I61955,I282873,I61599,I61593,I62000,I62017,I282885,I62034,I62051,I282888,I62077,I62085,I61587,I61581,I62139,I62147,I61596,I62205,I106968,I62231,I62248,I62270,I106983,I62296,I62304,I62321,I106980,I62338,I62355,I62372,I106977,I62389,I106992,I62406,I106989,I62423,I62454,I62471,I62488,I62505,I62550,I106986,I62595,I62612,I106974,I62629,I106995,I62646,I106971,I62672,I62680,I62734,I62742,I62800,I155277,I62826,I62843,I62792,I62865,I155271,I62891,I62899,I62916,I155286,I62933,I155283,I62950,I62967,I155274,I62984,I155265,I63001,I155268,I63018,I62768,I63049,I63066,I63083,I63100,I62780,I62774,I63145,I155289,I62789,I62783,I63190,I63207,I155280,I63224,I63241,I63267,I63275,I62777,I62771,I63329,I63337,I62786,I63395,I63421,I63438,I63387,I63460,I63486,I63494,I63511,I63528,I63545,I63562,I63579,I63596,I63613,I63363,I63644,I63661,I63678,I63695,I63375,I63369,I63740,I63384,I63378,I63785,I63802,I63819,I63836,I63862,I63870,I63372,I63366,I63924,I63932,I63381,I63990,I345360,I64016,I64033,I63982,I64055,I345345,I64081,I64089,I64106,I345363,I64123,I64140,I64157,I345366,I64174,I345357,I64191,I345354,I64208,I63958,I64239,I64256,I64273,I64290,I63970,I63964,I64335,I345351,I63979,I63973,I64380,I64397,I345342,I64414,I345348,I64431,I64457,I64465,I63967,I63961,I64519,I64527,I63976,I64585,I306752,I64611,I64628,I64577,I64650,I64676,I64684,I64701,I306755,I64718,I306767,I64735,I64752,I306773,I64769,I306764,I64786,I306770,I64803,I64553,I64834,I64851,I64868,I64885,I64565,I64559,I64930,I306761,I64574,I64568,I64975,I64992,I306758,I65009,I306776,I65026,I65052,I65060,I64562,I64556,I65114,I65122,I64571,I65180,I193442,I65206,I65223,I65172,I65245,I193439,I65271,I65279,I65296,I193445,I65313,I193430,I65330,I65347,I193433,I65364,I193454,I65381,I193451,I65398,I65148,I65429,I65446,I65463,I65480,I65160,I65154,I65525,I65169,I65163,I65570,I65587,I193436,I65604,I193448,I65621,I65647,I65655,I65157,I65151,I65709,I65717,I65166,I65775,I255750,I65801,I65818,I65767,I65840,I255759,I65866,I65874,I65891,I255747,I65908,I255738,I65925,I65942,I255744,I65959,I255762,I65976,I255735,I65993,I65743,I66024,I66041,I66058,I66075,I65755,I65749,I66120,I255741,I65764,I65758,I66165,I66182,I255753,I66199,I66216,I255756,I66242,I66250,I65752,I65746,I66304,I66312,I65761,I66370,I149922,I66396,I66413,I66362,I66435,I149916,I66461,I66469,I66486,I149931,I66503,I149928,I66520,I66537,I149919,I66554,I149910,I66571,I149913,I66588,I66338,I66619,I66636,I66653,I66670,I66350,I66344,I66715,I149934,I66359,I66353,I66760,I66777,I149925,I66794,I66811,I66837,I66845,I66347,I66341,I66899,I66907,I66356,I66965,I127409,I66991,I67008,I66957,I67030,I127397,I67056,I67064,I67081,I127406,I67098,I127403,I67115,I67132,I127394,I67149,I127400,I67166,I127385,I67183,I66933,I67214,I67231,I67248,I67265,I66945,I66939,I67310,I66954,I66948,I67355,I67372,I127391,I67389,I127388,I67406,I127412,I67432,I67440,I66942,I66936,I67494,I67502,I66951,I67560,I237755,I67586,I67603,I67552,I67625,I237749,I67651,I67659,I67676,I237767,I67693,I67710,I67727,I67744,I237761,I67761,I237752,I67778,I67528,I67809,I67826,I67843,I67860,I67540,I67534,I67905,I237764,I67549,I67543,I67950,I67967,I237770,I67984,I68001,I237758,I68027,I68035,I67537,I67531,I68089,I68097,I67546,I68155,I248822,I68181,I68198,I68147,I68220,I248816,I68246,I68254,I68271,I248834,I68288,I68305,I68322,I68339,I248828,I68356,I248819,I68373,I68123,I68404,I68421,I68438,I68455,I68135,I68129,I68500,I248831,I68144,I68138,I68545,I68562,I248837,I68579,I68596,I248825,I68622,I68630,I68132,I68126,I68684,I68692,I68141,I68750,I306174,I68776,I68793,I68742,I68815,I68841,I68849,I68866,I306177,I68883,I306189,I68900,I68917,I306195,I68934,I306186,I68951,I306192,I68968,I68718,I68999,I69016,I69033,I69050,I68730,I68724,I69095,I306183,I68739,I68733,I69140,I69157,I306180,I69174,I306198,I69191,I69217,I69225,I68727,I68721,I69279,I69287,I68736,I69345,I316578,I69371,I69388,I69337,I69410,I69436,I69444,I69461,I316581,I69478,I316593,I69495,I69512,I316599,I69529,I316590,I69546,I316596,I69563,I69313,I69594,I69611,I69628,I69645,I69325,I69319,I69690,I316587,I69334,I69328,I69735,I69752,I316584,I69769,I316602,I69786,I69812,I69820,I69322,I69316,I69874,I69882,I69331,I69940,I121969,I69966,I69983,I69932,I70005,I121957,I70031,I70039,I70056,I121966,I70073,I121963,I70090,I70107,I121954,I70124,I121960,I70141,I121945,I70158,I69908,I70189,I70206,I70223,I70240,I69920,I69914,I70285,I69929,I69923,I70330,I70347,I121951,I70364,I121948,I70381,I121972,I70407,I70415,I69917,I69911,I70469,I70477,I69926,I70535,I70561,I70578,I70527,I70600,I70626,I70634,I70651,I70668,I70685,I70702,I70719,I70736,I70753,I70503,I70784,I70801,I70818,I70835,I70515,I70509,I70880,I70524,I70518,I70925,I70942,I70959,I70976,I71002,I71010,I70512,I70506,I71064,I71072,I70521,I71130,I344272,I71156,I71173,I71122,I71195,I344257,I71221,I71229,I71246,I344275,I71263,I71280,I71297,I344278,I71314,I344269,I71331,I344266,I71348,I71098,I71379,I71396,I71413,I71430,I71110,I71104,I71475,I344263,I71119,I71113,I71520,I71537,I344254,I71554,I344260,I71571,I71597,I71605,I71107,I71101,I71659,I71667,I71116,I71725,I226388,I71751,I71768,I71717,I71790,I226385,I71816,I71824,I71841,I226391,I71858,I226376,I71875,I71892,I226379,I71909,I226400,I71926,I226397,I71943,I71693,I71974,I71991,I72008,I72025,I71705,I71699,I72070,I71714,I71708,I72115,I72132,I226382,I72149,I226394,I72166,I72192,I72200,I71702,I71696,I72254,I72262,I71711,I72320,I202690,I72346,I72363,I72312,I72385,I202687,I72411,I72419,I72436,I202693,I72453,I202678,I72470,I72487,I202681,I72504,I202702,I72521,I202699,I72538,I72288,I72569,I72586,I72603,I72620,I72300,I72294,I72665,I72309,I72303,I72710,I72727,I202684,I72744,I202696,I72761,I72787,I72795,I72297,I72291,I72849,I72857,I72306,I72915,I126865,I72941,I72958,I72907,I72980,I126853,I73006,I73014,I73031,I126862,I73048,I126859,I73065,I73082,I126850,I73099,I126856,I73116,I126841,I73133,I72883,I73164,I73181,I73198,I73215,I72895,I72889,I73260,I72904,I72898,I73305,I73322,I126847,I73339,I126844,I73356,I126868,I73382,I73390,I72892,I72886,I73444,I73452,I72901,I73510,I73536,I73553,I73502,I73575,I73601,I73609,I73626,I73643,I73660,I73677,I73694,I73711,I73728,I73478,I73759,I73776,I73793,I73810,I73490,I73484,I73855,I73499,I73493,I73900,I73917,I73934,I73951,I73977,I73985,I73487,I73481,I74039,I74047,I73496,I74105,I138289,I74131,I74148,I74097,I74170,I138277,I74196,I74204,I74221,I138286,I74238,I138283,I74255,I74272,I138274,I74289,I138280,I74306,I138265,I74323,I74073,I74354,I74371,I74388,I74405,I74085,I74079,I74450,I74094,I74088,I74495,I74512,I138271,I74529,I138268,I74546,I138292,I74572,I74580,I74082,I74076,I74634,I74642,I74091,I74700,I183038,I74726,I74743,I74765,I183035,I74791,I74799,I74816,I183041,I74833,I183026,I74850,I74867,I183029,I74884,I183050,I74901,I183047,I74918,I74949,I74966,I74983,I75000,I75045,I75090,I75107,I183032,I75124,I183044,I75141,I75167,I75175,I75229,I75237,I75295,I75321,I75338,I75360,I75386,I75394,I75411,I75428,I75445,I75462,I75479,I75496,I75513,I75544,I75561,I75578,I75595,I75640,I75685,I75702,I75719,I75736,I75762,I75770,I75824,I75832,I75890,I116529,I75916,I75933,I75882,I75955,I116517,I75981,I75989,I76006,I116526,I76023,I116523,I76040,I76057,I116514,I76074,I116520,I76091,I116505,I76108,I75858,I76139,I76156,I76173,I76190,I75870,I75864,I76235,I75879,I75873,I76280,I76297,I116511,I76314,I116508,I76331,I116532,I76357,I76365,I75867,I75861,I76419,I76427,I75876,I76485,I158765,I76511,I76528,I76477,I76550,I158756,I76576,I76584,I76601,I158774,I76618,I158771,I76635,I76652,I158750,I76669,I158753,I76686,I158762,I76703,I76453,I76734,I76751,I76768,I76785,I76465,I76459,I76830,I158768,I76474,I76468,I76875,I76892,I76909,I158759,I76926,I76952,I76960,I76462,I76456,I77014,I77022,I76471,I77080,I221764,I77106,I77123,I77072,I77145,I221761,I77171,I77179,I77196,I221767,I77213,I221752,I77230,I77247,I221755,I77264,I221776,I77281,I221773,I77298,I77048,I77329,I77346,I77363,I77380,I77060,I77054,I77425,I77069,I77063,I77470,I77487,I221758,I77504,I221770,I77521,I77547,I77555,I77057,I77051,I77609,I77617,I77066,I77675,I115441,I77701,I77718,I77667,I77740,I115429,I77766,I77774,I77791,I115438,I77808,I115435,I77825,I77842,I115426,I77859,I115432,I77876,I115417,I77893,I77643,I77924,I77941,I77958,I77975,I77655,I77649,I78020,I77664,I77658,I78065,I78082,I115423,I78099,I115420,I78116,I115444,I78142,I78150,I77652,I77646,I78204,I78212,I77661,I78270,I308486,I78296,I78313,I78262,I78335,I78361,I78369,I78386,I308489,I78403,I308501,I78420,I78437,I308507,I78454,I308498,I78471,I308504,I78488,I78238,I78519,I78536,I78553,I78570,I78250,I78244,I78615,I308495,I78259,I78253,I78660,I78677,I308492,I78694,I308510,I78711,I78737,I78745,I78247,I78241,I78799,I78807,I78256,I78865,I215406,I78891,I78908,I78930,I215403,I78956,I78964,I78981,I215409,I78998,I215394,I79015,I79032,I215397,I79049,I215418,I79066,I215415,I79083,I79114,I79131,I79148,I79165,I79210,I79255,I79272,I215400,I79289,I215412,I79306,I79332,I79340,I79394,I79402,I79460,I240917,I79486,I79503,I79452,I79525,I240911,I79551,I79559,I79576,I240929,I79593,I79610,I79627,I79644,I240923,I79661,I240914,I79678,I79428,I79709,I79726,I79743,I79760,I79440,I79434,I79805,I240926,I79449,I79443,I79850,I79867,I240932,I79884,I79901,I240920,I79927,I79935,I79437,I79431,I79989,I79997,I79446,I80055,I270608,I80081,I80098,I80047,I80120,I270617,I80146,I80154,I80171,I270605,I80188,I270596,I80205,I80222,I270602,I80239,I270620,I80256,I270593,I80273,I80023,I80304,I80321,I80338,I80355,I80035,I80029,I80400,I270599,I80044,I80038,I80445,I80462,I270611,I80479,I80496,I270614,I80522,I80530,I80032,I80026,I80584,I80592,I80041,I80653,I131749,I80679,I80687,I131761,I131740,I80704,I131764,I80730,I80621,I80752,I131755,I80778,I80786,I131737,I80803,I80829,I80645,I80851,I80627,I131752,I80891,I80908,I80916,I80933,I80630,I80964,I131743,I80981,I131746,I81007,I81015,I80618,I80636,I81060,I131758,I81077,I80639,I80624,I80633,I80642,I81180,I81206,I81214,I81231,I81257,I81148,I81279,I81305,I81313,I81330,I81356,I81172,I81378,I81154,I81418,I81435,I81443,I81460,I81157,I81491,I81508,I81534,I81542,I81145,I81163,I81587,I81604,I81166,I81151,I81160,I81169,I81707,I307330,I81733,I81741,I307345,I81758,I307348,I81784,I81675,I81806,I307354,I81832,I81840,I307336,I81857,I81883,I81699,I81905,I81681,I307333,I81945,I81962,I81970,I81987,I81684,I82018,I307339,I82035,I307351,I82061,I82069,I81672,I81690,I82114,I307342,I82131,I81693,I81678,I81687,I81696,I82234,I328716,I82260,I82268,I328731,I82285,I328734,I82311,I82202,I82333,I328740,I82359,I82367,I328722,I82384,I82410,I82226,I82432,I82208,I328719,I82472,I82489,I82497,I82514,I82211,I82545,I328725,I82562,I328737,I82588,I82596,I82199,I82217,I82641,I328728,I82658,I82220,I82205,I82214,I82223,I82761,I82787,I82795,I82812,I82838,I82860,I82886,I82894,I82911,I82937,I82959,I82999,I83016,I83024,I83041,I83072,I83089,I83115,I83123,I83168,I83185,I83288,I240387,I83314,I83322,I240390,I240384,I83339,I240396,I83365,I83256,I83387,I240399,I83413,I83421,I83438,I83464,I83280,I83486,I83262,I240402,I83526,I83543,I83551,I83568,I83265,I83599,I240393,I83616,I83642,I83650,I83253,I83271,I83695,I240405,I83712,I83274,I83259,I83268,I83277,I83815,I291013,I83841,I83849,I291010,I83866,I291022,I83892,I83914,I83940,I83948,I291028,I83965,I83991,I84013,I291016,I84053,I84070,I84078,I84095,I84126,I291025,I291031,I84143,I84169,I84177,I84222,I291019,I84239,I84342,I320046,I84368,I84376,I320061,I84393,I320064,I84419,I84310,I84441,I320070,I84467,I84475,I320052,I84492,I84518,I84334,I84540,I84316,I320049,I84580,I84597,I84605,I84622,I84319,I84653,I320055,I84670,I320067,I84696,I84704,I84307,I84325,I84749,I320058,I84766,I84328,I84313,I84322,I84331,I84869,I249873,I84895,I84903,I249876,I249870,I84920,I249882,I84946,I84837,I84968,I249885,I84994,I85002,I85019,I85045,I84861,I85067,I84843,I249888,I85107,I85124,I85132,I85149,I84846,I85180,I249879,I85197,I85223,I85231,I84834,I84852,I85276,I249891,I85293,I84855,I84840,I84849,I84858,I85396,I210204,I85422,I85430,I210195,I210210,I85447,I210216,I85473,I85364,I85495,I210201,I85521,I85529,I85546,I85572,I85388,I85594,I85370,I210198,I85634,I85651,I85659,I85676,I85373,I85707,I210192,I210207,I85724,I85750,I85758,I85361,I85379,I85803,I210213,I85820,I85382,I85367,I85376,I85385,I85923,I85949,I85957,I85974,I86000,I85891,I86022,I86048,I86056,I86073,I86099,I85915,I86121,I85897,I86161,I86178,I86186,I86203,I85900,I86234,I86251,I86277,I86285,I85888,I85906,I86330,I86347,I85909,I85894,I85903,I85912,I86450,I203268,I86476,I86484,I203259,I203274,I86501,I203280,I86527,I86418,I86549,I203265,I86575,I86583,I86600,I86626,I86442,I86648,I86424,I203262,I86688,I86705,I86713,I86730,I86427,I86761,I203256,I203271,I86778,I86804,I86812,I86415,I86433,I86857,I203277,I86874,I86436,I86421,I86430,I86439,I86977,I87003,I87011,I87028,I87054,I86945,I87076,I87102,I87110,I87127,I87153,I86969,I87175,I86951,I87215,I87232,I87240,I87257,I86954,I87288,I87305,I87331,I87339,I86942,I86960,I87384,I87401,I86963,I86948,I86957,I86966,I87504,I381284,I87530,I87538,I381263,I87555,I381290,I87581,I87472,I87603,I381278,I87629,I87637,I381281,I87654,I87680,I87496,I87702,I87478,I381272,I87742,I87759,I87767,I87784,I87481,I87815,I381269,I381266,I87832,I381287,I87858,I87866,I87469,I87487,I87911,I381275,I87928,I87490,I87475,I87484,I87493,I88031,I149318,I88057,I88065,I149330,I88082,I149315,I88108,I88130,I149339,I88156,I88164,I149336,I88181,I88207,I88229,I149327,I88269,I88286,I88294,I88311,I88342,I149324,I88359,I149333,I88385,I88393,I88438,I149321,I88455,I88558,I88584,I88592,I88609,I88635,I88526,I88657,I88683,I88691,I88708,I88734,I88550,I88756,I88532,I88796,I88813,I88821,I88838,I88535,I88869,I88886,I88912,I88920,I88523,I88541,I88965,I88982,I88544,I88529,I88538,I88547,I89085,I322936,I89111,I89119,I322951,I89136,I322954,I89162,I89053,I89184,I322960,I89210,I89218,I322942,I89235,I89261,I89077,I89283,I89059,I322939,I89323,I89340,I89348,I89365,I89062,I89396,I322945,I89413,I322957,I89439,I89447,I89050,I89068,I89492,I322948,I89509,I89071,I89056,I89065,I89074,I89612,I89638,I89646,I89663,I89689,I89580,I89711,I89737,I89745,I89762,I89788,I89604,I89810,I89586,I89850,I89867,I89875,I89892,I89589,I89923,I89940,I89966,I89974,I89577,I89595,I90019,I90036,I89598,I89583,I89592,I89601,I90139,I320624,I90165,I90173,I320639,I90190,I320642,I90216,I90238,I320648,I90264,I90272,I320630,I90289,I90315,I90337,I320627,I90377,I90394,I90402,I90419,I90450,I320633,I90467,I320645,I90493,I90501,I90546,I320636,I90563,I90666,I249346,I90692,I90700,I249349,I249343,I90717,I249355,I90743,I90634,I90765,I249358,I90791,I90799,I90816,I90842,I90658,I90864,I90640,I249361,I90904,I90921,I90929,I90946,I90643,I90977,I249352,I90994,I91020,I91028,I90631,I90649,I91073,I249364,I91090,I90652,I90637,I90646,I90655,I91193,I139909,I91219,I91227,I139921,I139900,I91244,I139924,I91270,I91161,I91292,I139915,I91318,I91326,I139897,I91343,I91369,I91185,I91391,I91167,I139912,I91431,I91448,I91456,I91473,I91170,I91504,I139903,I91521,I139906,I91547,I91555,I91158,I91176,I91600,I139918,I91617,I91179,I91164,I91173,I91182,I91720,I262844,I91746,I91754,I262841,I262859,I91771,I262850,I91797,I91688,I91819,I262865,I91845,I91853,I262847,I91870,I91896,I91712,I91918,I91694,I262853,I91958,I91975,I91983,I92000,I91697,I92031,I262868,I92048,I262856,I92074,I92082,I91685,I91703,I92127,I262862,I92144,I91706,I91691,I91700,I91709,I92247,I234590,I92273,I92281,I234593,I234587,I92298,I234599,I92324,I92215,I92346,I234602,I92372,I92380,I92397,I92423,I92239,I92445,I92221,I234605,I92485,I92502,I92510,I92527,I92224,I92558,I234596,I92575,I92601,I92609,I92212,I92230,I92654,I234608,I92671,I92233,I92218,I92227,I92236,I92774,I206736,I92800,I92808,I206727,I206742,I92825,I206748,I92851,I92742,I92873,I206733,I92899,I92907,I92924,I92950,I92766,I92972,I92748,I206730,I93012,I93029,I93037,I93054,I92751,I93085,I206724,I206739,I93102,I93128,I93136,I92739,I92757,I93181,I206745,I93198,I92760,I92745,I92754,I92763,I93301,I209626,I93327,I93335,I209617,I209632,I93352,I209638,I93378,I93269,I93400,I209623,I93426,I93434,I93451,I93477,I93293,I93499,I93275,I209620,I93539,I93556,I93564,I93581,I93278,I93612,I209614,I209629,I93629,I93655,I93663,I93266,I93284,I93708,I209635,I93725,I93287,I93272,I93281,I93290,I93828,I204424,I93854,I93862,I204415,I204430,I93879,I204436,I93905,I93796,I93927,I204421,I93953,I93961,I93978,I94004,I93820,I94026,I93802,I204418,I94066,I94083,I94091,I94108,I93805,I94139,I204412,I204427,I94156,I94182,I94190,I93793,I93811,I94235,I204433,I94252,I93814,I93799,I93808,I93817,I94355,I387234,I94381,I94389,I387213,I94406,I387240,I94432,I94454,I387228,I94480,I94488,I387231,I94505,I94531,I94553,I387222,I94593,I94610,I94618,I94635,I94666,I387219,I387216,I94683,I387237,I94709,I94717,I94762,I387225,I94779,I94882,I242495,I94908,I94916,I242498,I242492,I94933,I242504,I94959,I94850,I94981,I242507,I95007,I95015,I95032,I95058,I94874,I95080,I94856,I242510,I95120,I95137,I95145,I95162,I94859,I95193,I242501,I95210,I95236,I95244,I94847,I94865,I95289,I242513,I95306,I94868,I94853,I94862,I94871,I95409,I95435,I95443,I95460,I95486,I95377,I95508,I95534,I95542,I95559,I95585,I95401,I95607,I95383,I95647,I95664,I95672,I95689,I95386,I95720,I95737,I95763,I95771,I95374,I95392,I95816,I95833,I95395,I95380,I95389,I95398,I95936,I115973,I95962,I95970,I115985,I115964,I95987,I115988,I96013,I95904,I96035,I115979,I96061,I96069,I115961,I96086,I96112,I95928,I96134,I95910,I115976,I96174,I96191,I96199,I96216,I95913,I96247,I115967,I96264,I115970,I96290,I96298,I95901,I95919,I96343,I115982,I96360,I95922,I95907,I95916,I95925,I96463,I207892,I96489,I96497,I207883,I207898,I96514,I207904,I96540,I96431,I96562,I207889,I96588,I96596,I96613,I96639,I96455,I96661,I96437,I207886,I96701,I96718,I96726,I96743,I96440,I96774,I207880,I207895,I96791,I96817,I96825,I96428,I96446,I96870,I207901,I96887,I96449,I96434,I96443,I96452,I96990,I275764,I97016,I97024,I275761,I275779,I97041,I275770,I97067,I96958,I97089,I275785,I97115,I97123,I275767,I97140,I97166,I96982,I97188,I96964,I275773,I97228,I97245,I97253,I97270,I96967,I97301,I275788,I97318,I275776,I97344,I97352,I96955,I96973,I97397,I275782,I97414,I96976,I96961,I96970,I96979,I97517,I328138,I97543,I97551,I328153,I97568,I328156,I97594,I97485,I97616,I328162,I97642,I97650,I328144,I97667,I97693,I97509,I97715,I97491,I328141,I97755,I97772,I97780,I97797,I97494,I97828,I328147,I97845,I328159,I97871,I97879,I97482,I97500,I97924,I328150,I97941,I97503,I97488,I97497,I97506,I98044,I378309,I98070,I98078,I378288,I98095,I378315,I98121,I98012,I98143,I378303,I98169,I98177,I378306,I98194,I98220,I98036,I98242,I98018,I378297,I98282,I98299,I98307,I98324,I98021,I98355,I378294,I378291,I98372,I378312,I98398,I98406,I98009,I98027,I98451,I378300,I98468,I98030,I98015,I98024,I98033,I98571,I210782,I98597,I98605,I210773,I210788,I98622,I210794,I98648,I98539,I98670,I210779,I98696,I98704,I98721,I98747,I98563,I98769,I98545,I210776,I98809,I98826,I98834,I98851,I98548,I98882,I210770,I210785,I98899,I98925,I98933,I98536,I98554,I98978,I210791,I98995,I98557,I98542,I98551,I98560,I99098,I99124,I99132,I99149,I99175,I99197,I99223,I99231,I99248,I99274,I99296,I99336,I99353,I99361,I99378,I99409,I99426,I99452,I99460,I99505,I99522,I99625,I99651,I99659,I99676,I99702,I99724,I99750,I99758,I99775,I99801,I99823,I99863,I99880,I99888,I99905,I99936,I99953,I99979,I99987,I100032,I100049,I100152,I162233,I100178,I100186,I162218,I162221,I100203,I162236,I100229,I100120,I100251,I162230,I100277,I100285,I100302,I100328,I100144,I100350,I100126,I162227,I100390,I100407,I100415,I100432,I100129,I100463,I162242,I100480,I162239,I100506,I100514,I100117,I100135,I100559,I162224,I100576,I100138,I100123,I100132,I100141,I100679,I245130,I100705,I100713,I245133,I245127,I100730,I245139,I100756,I100778,I245142,I100804,I100812,I100829,I100855,I100877,I245145,I100917,I100934,I100942,I100959,I100990,I245136,I101007,I101033,I101041,I101086,I245148,I101103,I101206,I101232,I101240,I101257,I101283,I101174,I101305,I101331,I101339,I101356,I101382,I101198,I101404,I101180,I101444,I101461,I101469,I101486,I101183,I101517,I101534,I101560,I101568,I101171,I101189,I101613,I101630,I101192,I101177,I101186,I101195,I101733,I133381,I101759,I101767,I133393,I133372,I101784,I133396,I101810,I101832,I133387,I101858,I101866,I133369,I101883,I101909,I101931,I133384,I101971,I101988,I101996,I102013,I102044,I133375,I102061,I133378,I102087,I102095,I102140,I133390,I102157,I102260,I180729,I102286,I102294,I180714,I180717,I102311,I180732,I102337,I102228,I102359,I180726,I102385,I102393,I102410,I102436,I102252,I102458,I102234,I180723,I102498,I102515,I102523,I102540,I102237,I102571,I180738,I102588,I180735,I102614,I102622,I102225,I102243,I102667,I180720,I102684,I102246,I102231,I102240,I102249,I102787,I386639,I102813,I102821,I386618,I102838,I386645,I102864,I102755,I102886,I386633,I102912,I102920,I386636,I102937,I102963,I102779,I102985,I102761,I386627,I103025,I103042,I103050,I103067,I102764,I103098,I386624,I386621,I103115,I386642,I103141,I103149,I102752,I102770,I103194,I386630,I103211,I102773,I102758,I102767,I102776,I103314,I103340,I103348,I103365,I103391,I103282,I103413,I103439,I103447,I103464,I103490,I103306,I103512,I103288,I103552,I103569,I103577,I103594,I103291,I103625,I103642,I103668,I103676,I103279,I103297,I103721,I103738,I103300,I103285,I103294,I103303,I103841,I202112,I103867,I103875,I202103,I202118,I103892,I202124,I103918,I103809,I103940,I202109,I103966,I103974,I103991,I104017,I103833,I104039,I103815,I202106,I104079,I104096,I104104,I104121,I103818,I104152,I202100,I202115,I104169,I104195,I104203,I103806,I103824,I104248,I202121,I104265,I103827,I103812,I103821,I103830,I104368,I343728,I104394,I104402,I343710,I343734,I104419,I343725,I104445,I104336,I104467,I343731,I104493,I104501,I343719,I104518,I104544,I104360,I104566,I104342,I104606,I104623,I104631,I104648,I104345,I104679,I343716,I343713,I104696,I343722,I104722,I104730,I104333,I104351,I104775,I104792,I104354,I104339,I104348,I104357,I104895,I104921,I104929,I104946,I104972,I104863,I104994,I105020,I105028,I105045,I105071,I104887,I105093,I104869,I105133,I105150,I105158,I105175,I104872,I105206,I105223,I105249,I105257,I104860,I104878,I105302,I105319,I104881,I104866,I104875,I104884,I105422,I134469,I105448,I105456,I134481,I134460,I105473,I134484,I105499,I105390,I105521,I134475,I105547,I105555,I134457,I105572,I105598,I105414,I105620,I105396,I134472,I105660,I105677,I105685,I105702,I105399,I105733,I134463,I105750,I134466,I105776,I105784,I105387,I105405,I105829,I134478,I105846,I105408,I105393,I105402,I105411,I105949,I200956,I105975,I105983,I200947,I200962,I106000,I200968,I106026,I105917,I106048,I200953,I106074,I106082,I106099,I106125,I105941,I106147,I105923,I200950,I106187,I106204,I106212,I106229,I105926,I106260,I200944,I200959,I106277,I106303,I106311,I105914,I105932,I106356,I200965,I106373,I105935,I105920,I105929,I105938,I106476,I321780,I106502,I106510,I321795,I106527,I321798,I106553,I106444,I106575,I321804,I106601,I106609,I321786,I106626,I106652,I106468,I106674,I106450,I321783,I106714,I106731,I106739,I106756,I106453,I106787,I321789,I106804,I321801,I106830,I106838,I106441,I106459,I106883,I321792,I106900,I106462,I106447,I106456,I106465,I107003,I170325,I107029,I107037,I170310,I170313,I107054,I170328,I107080,I107102,I170322,I107128,I107136,I107153,I107179,I107201,I170319,I107241,I107258,I107266,I107283,I107314,I170334,I107331,I170331,I107357,I107365,I107410,I170316,I107427,I107530,I321202,I107556,I107564,I321217,I107581,I321220,I107607,I107498,I107629,I321226,I107655,I107663,I321208,I107680,I107706,I107522,I107728,I107504,I321205,I107768,I107785,I107793,I107810,I107507,I107841,I321211,I107858,I321223,I107884,I107892,I107495,I107513,I107937,I321214,I107954,I107516,I107501,I107510,I107519,I108057,I108083,I108091,I108108,I108134,I108156,I108182,I108190,I108207,I108233,I108255,I108295,I108312,I108320,I108337,I108368,I108385,I108411,I108419,I108464,I108481,I108584,I108610,I108618,I108635,I108661,I108683,I108709,I108717,I108734,I108760,I108782,I108822,I108839,I108847,I108864,I108895,I108912,I108938,I108946,I108991,I109008,I109111,I109137,I109145,I109162,I109188,I109079,I109210,I109236,I109244,I109261,I109287,I109103,I109309,I109085,I109349,I109366,I109374,I109391,I109088,I109422,I109439,I109465,I109473,I109076,I109094,I109518,I109535,I109097,I109082,I109091,I109100,I109638,I109664,I109672,I109689,I109715,I109606,I109737,I109763,I109771,I109788,I109814,I109630,I109836,I109612,I109876,I109893,I109901,I109918,I109615,I109949,I109966,I109992,I110000,I109603,I109621,I110045,I110062,I109624,I109609,I109618,I109627,I110165,I110191,I110199,I110216,I110242,I110133,I110264,I110290,I110298,I110315,I110341,I110157,I110363,I110139,I110403,I110420,I110428,I110445,I110142,I110476,I110493,I110519,I110527,I110130,I110148,I110572,I110589,I110151,I110136,I110145,I110154,I110692,I283516,I110718,I110726,I283513,I283531,I110743,I283522,I110769,I110660,I110791,I283537,I110817,I110825,I283519,I110842,I110868,I110684,I110890,I110666,I283525,I110930,I110947,I110955,I110972,I110669,I111003,I283540,I111020,I283528,I111046,I111054,I110657,I110675,I111099,I283534,I111116,I110678,I110663,I110672,I110681,I111219,I212516,I111245,I111253,I212507,I212522,I111270,I212528,I111296,I111187,I111318,I212513,I111344,I111352,I111369,I111395,I111211,I111417,I111193,I212510,I111457,I111474,I111482,I111499,I111196,I111530,I212504,I212519,I111547,I111573,I111581,I111184,I111202,I111626,I212525,I111643,I111205,I111190,I111199,I111208,I111746,I333340,I111772,I111780,I333355,I111797,I333358,I111823,I111845,I333364,I111871,I111879,I333346,I111896,I111922,I111944,I333343,I111984,I112001,I112009,I112026,I112057,I333349,I112074,I333361,I112100,I112108,I112153,I333352,I112170,I112273,I145748,I112299,I112307,I145760,I112324,I145745,I112350,I112241,I112372,I145769,I112398,I112406,I145766,I112423,I112449,I112265,I112471,I112247,I145757,I112511,I112528,I112536,I112553,I112250,I112584,I145754,I112601,I145763,I112627,I112635,I112238,I112256,I112680,I145751,I112697,I112259,I112244,I112253,I112262,I112800,I188240,I112826,I112834,I188231,I188246,I112851,I188252,I112877,I112768,I112899,I188237,I112925,I112933,I112950,I112976,I112792,I112998,I112774,I188234,I113038,I113055,I113063,I113080,I112777,I113111,I188228,I188243,I113128,I113154,I113162,I112765,I112783,I113207,I188249,I113224,I112786,I112771,I112780,I112789,I113327,I272534,I113353,I113361,I272531,I272549,I113378,I272540,I113404,I113426,I272555,I113452,I113460,I272537,I113477,I113503,I113525,I272543,I113565,I113582,I113590,I113607,I113638,I272558,I113655,I272546,I113681,I113689,I113734,I272552,I113751,I113854,I195176,I113880,I113888,I195167,I195182,I113905,I195188,I113931,I113822,I113953,I195173,I113979,I113987,I114004,I114030,I113846,I114052,I113828,I195170,I114092,I114109,I114117,I114134,I113831,I114165,I195164,I195179,I114182,I114208,I114216,I113819,I113837,I114261,I195185,I114278,I113840,I113825,I113834,I113843,I114381,I119781,I114407,I114415,I119793,I119772,I114432,I119796,I114458,I114480,I119787,I114506,I114514,I119769,I114531,I114557,I114579,I119784,I114619,I114636,I114644,I114661,I114692,I119775,I114709,I119778,I114735,I114743,I114788,I119790,I114805,I114908,I282227,I114934,I114951,I114900,I114973,I114990,I282242,I282230,I115007,I282221,I115033,I115041,I282233,I115067,I115075,I282224,I115092,I114879,I282239,I115132,I115140,I114873,I114888,I115185,I282248,I282236,I115202,I282245,I115228,I114876,I115250,I115267,I115284,I114891,I115315,I115332,I114882,I115363,I114885,I114897,I114894,I115452,I155863,I115478,I115495,I115517,I115534,I155860,I155881,I115551,I155884,I115577,I115585,I155869,I115611,I115619,I155872,I115636,I155875,I115676,I115684,I115729,I155866,I115746,I155878,I115772,I115794,I115811,I115828,I115859,I115876,I115907,I115996,I116022,I116039,I116061,I116078,I116095,I116121,I116129,I116155,I116163,I116180,I116220,I116228,I116273,I116290,I116316,I116338,I116355,I116372,I116403,I116420,I116451,I116540,I377125,I116566,I116583,I116605,I116622,I377101,I377122,I116639,I377119,I116665,I116673,I377098,I116699,I116707,I377110,I116724,I377113,I116764,I116772,I116817,I377116,I377104,I116834,I377107,I116860,I116882,I116899,I116916,I116947,I116964,I116995,I117084,I325251,I117110,I117127,I117076,I117149,I117166,I325263,I117183,I325254,I117209,I117217,I325272,I117243,I117251,I325248,I117268,I117055,I325266,I117308,I117316,I117049,I117064,I117361,I325260,I325257,I117378,I325269,I117404,I117052,I117426,I117443,I117460,I117067,I117491,I117508,I117058,I117539,I117061,I117073,I117070,I117628,I361408,I117654,I117671,I117620,I117693,I117710,I361405,I361402,I117727,I361390,I117753,I117761,I361414,I117787,I117795,I361399,I117812,I117599,I361393,I117852,I117860,I117593,I117608,I117905,I361396,I117922,I361411,I117948,I117596,I117970,I117987,I118004,I117611,I118035,I118052,I117602,I118083,I117605,I117617,I117614,I118172,I250409,I118198,I118215,I118164,I118237,I118254,I250403,I250400,I118271,I250415,I118297,I118305,I118331,I118339,I250397,I118356,I118143,I118396,I118404,I118137,I118152,I118449,I250412,I250406,I118466,I118492,I118140,I118514,I118531,I118548,I118155,I118579,I118596,I250418,I118146,I118627,I118149,I118161,I118158,I118716,I224067,I118742,I118759,I118708,I118781,I118798,I224088,I224079,I118815,I118841,I118849,I224073,I118875,I118883,I224070,I118900,I118687,I224064,I118940,I118948,I118681,I118696,I118993,I224076,I119010,I224085,I119036,I118684,I119058,I119075,I119092,I118699,I119123,I119140,I224082,I118690,I119171,I118693,I118705,I118702,I119260,I181873,I119286,I119303,I119252,I119325,I119342,I181894,I181885,I119359,I119385,I119393,I181879,I119419,I119427,I181876,I119444,I119231,I181870,I119484,I119492,I119225,I119240,I119537,I181882,I119554,I181891,I119580,I119228,I119602,I119619,I119636,I119243,I119667,I119684,I181888,I119234,I119715,I119237,I119249,I119246,I119804,I245666,I119830,I119847,I119869,I119886,I245660,I245657,I119903,I245672,I119929,I119937,I119963,I119971,I245654,I119988,I120028,I120036,I120081,I245669,I245663,I120098,I120124,I120146,I120163,I120180,I120211,I120228,I245675,I120259,I120348,I355681,I120374,I120391,I120340,I120413,I120430,I355693,I355696,I120447,I355699,I120473,I120481,I355684,I120507,I120515,I355690,I120532,I120319,I355678,I120572,I120580,I120313,I120328,I120625,I355702,I120642,I355687,I120668,I120316,I120690,I120707,I120724,I120331,I120755,I120772,I120322,I120803,I120325,I120337,I120334,I120892,I225801,I120918,I120935,I120884,I120957,I120974,I225822,I225813,I120991,I121017,I121025,I225807,I121051,I121059,I225804,I121076,I120863,I225798,I121116,I121124,I120857,I120872,I121169,I225810,I121186,I225819,I121212,I120860,I121234,I121251,I121268,I120875,I121299,I121316,I225816,I120866,I121347,I120869,I120881,I120878,I121436,I362564,I121462,I121479,I121428,I121501,I121518,I362561,I362558,I121535,I362546,I121561,I121569,I362570,I121595,I121603,I362555,I121620,I121407,I362549,I121660,I121668,I121401,I121416,I121713,I362552,I121730,I362567,I121756,I121404,I121778,I121795,I121812,I121419,I121843,I121860,I121410,I121891,I121413,I121425,I121422,I121980,I348609,I122006,I122023,I122045,I122062,I348621,I348624,I122079,I348627,I122105,I122113,I348612,I122139,I122147,I348618,I122164,I348606,I122204,I122212,I122257,I348630,I122274,I348615,I122300,I122322,I122339,I122356,I122387,I122404,I122435,I122524,I122550,I122567,I122589,I122606,I122623,I122649,I122657,I122683,I122691,I122708,I122748,I122756,I122801,I122818,I122844,I122866,I122883,I122900,I122931,I122948,I122979,I123068,I297742,I123094,I123111,I123060,I123133,I123150,I297760,I123167,I297754,I123193,I123201,I297748,I123227,I123235,I297757,I123252,I123039,I297745,I123292,I123300,I123033,I123048,I123345,I297763,I123362,I123388,I123036,I123410,I123427,I123444,I123051,I123475,I123492,I297751,I123042,I123523,I123045,I123057,I123054,I123612,I168001,I123638,I123655,I123604,I123677,I123694,I167998,I168019,I123711,I168022,I123737,I123745,I168007,I123771,I123779,I168010,I123796,I123583,I168013,I123836,I123844,I123577,I123592,I123889,I168004,I123906,I168016,I123932,I123580,I123954,I123971,I123988,I123595,I124019,I124036,I123586,I124067,I123589,I123601,I123598,I124156,I152888,I124182,I124199,I124148,I124221,I124238,I152891,I152909,I124255,I152897,I124281,I124289,I124315,I124323,I152906,I124340,I124127,I152900,I124380,I124388,I124121,I124136,I124433,I152903,I152885,I124450,I152894,I124476,I124124,I124498,I124515,I124532,I124139,I124563,I124580,I124130,I124611,I124133,I124145,I124142,I124700,I331609,I124726,I124743,I124692,I124765,I124782,I331621,I124799,I331612,I124825,I124833,I331630,I124859,I124867,I331606,I124884,I124671,I331624,I124924,I124932,I124665,I124680,I124977,I331618,I331615,I124994,I331627,I125020,I124668,I125042,I125059,I125076,I124683,I125107,I125124,I124674,I125155,I124677,I124689,I124686,I125244,I142178,I125270,I125287,I125236,I125309,I125326,I142181,I142199,I125343,I142187,I125369,I125377,I125403,I125411,I142196,I125428,I125215,I142190,I125468,I125476,I125209,I125224,I125521,I142193,I142175,I125538,I142184,I125564,I125212,I125586,I125603,I125620,I125227,I125651,I125668,I125218,I125699,I125221,I125233,I125230,I125788,I382480,I125814,I125831,I125780,I125853,I125870,I382456,I382477,I125887,I382474,I125913,I125921,I382453,I125947,I125955,I382465,I125972,I125759,I382468,I126012,I126020,I125753,I125768,I126065,I382471,I382459,I126082,I382462,I126108,I125756,I126130,I126147,I126164,I125771,I126195,I126212,I125762,I126243,I125765,I125777,I125774,I126332,I126358,I126375,I126397,I126414,I126431,I126457,I126465,I126491,I126499,I126516,I126556,I126564,I126609,I126626,I126652,I126674,I126691,I126708,I126739,I126756,I126787,I126876,I171469,I126902,I126919,I126941,I126958,I171466,I171487,I126975,I171490,I127001,I127009,I171475,I127035,I127043,I171478,I127060,I171481,I127100,I127108,I127153,I171472,I127170,I171484,I127196,I127218,I127235,I127252,I127283,I127300,I127331,I127420,I127446,I127463,I127485,I127502,I127519,I127545,I127553,I127579,I127587,I127604,I127644,I127652,I127697,I127714,I127740,I127762,I127779,I127796,I127827,I127844,I127875,I127964,I127990,I128007,I128029,I128046,I128063,I128089,I128097,I128123,I128131,I128148,I128188,I128196,I128241,I128258,I128284,I128306,I128323,I128340,I128371,I128388,I128419,I128508,I128534,I128551,I128500,I128573,I128590,I128607,I128633,I128641,I128667,I128675,I128692,I128479,I128732,I128740,I128473,I128488,I128785,I128802,I128828,I128476,I128850,I128867,I128884,I128491,I128915,I128932,I128482,I128963,I128485,I128497,I128494,I129052,I197479,I129078,I129095,I129117,I129134,I197500,I197491,I129151,I129177,I129185,I197485,I129211,I129219,I197482,I129236,I197476,I129276,I129284,I129329,I197488,I129346,I197497,I129372,I129394,I129411,I129428,I129459,I129476,I197494,I129507,I129596,I129622,I129639,I129588,I129661,I129678,I129695,I129721,I129729,I129755,I129763,I129780,I129567,I129820,I129828,I129561,I129576,I129873,I129890,I129916,I129564,I129938,I129955,I129972,I129579,I130003,I130020,I129570,I130051,I129573,I129585,I129582,I130140,I130166,I130183,I130132,I130205,I130222,I130239,I130265,I130273,I130299,I130307,I130324,I130111,I130364,I130372,I130105,I130120,I130417,I130434,I130460,I130108,I130482,I130499,I130516,I130123,I130547,I130564,I130114,I130595,I130117,I130129,I130126,I130684,I235126,I130710,I130727,I130676,I130749,I130766,I235120,I235117,I130783,I235132,I130809,I130817,I130843,I130851,I235114,I130868,I130655,I130908,I130916,I130649,I130664,I130961,I235129,I235123,I130978,I131004,I130652,I131026,I131043,I131060,I130667,I131091,I131108,I235135,I130658,I131139,I130661,I130673,I130670,I131228,I131254,I131271,I131293,I131310,I131327,I131353,I131361,I131387,I131395,I131412,I131452,I131460,I131505,I131522,I131548,I131570,I131587,I131604,I131635,I131652,I131683,I131772,I237234,I131798,I131815,I131837,I131854,I237228,I237225,I131871,I237240,I131897,I131905,I131931,I131939,I237222,I131956,I131996,I132004,I132049,I237237,I237231,I132066,I132092,I132114,I132131,I132148,I132179,I132196,I237243,I132227,I132316,I132342,I132359,I132308,I132381,I132398,I132415,I132441,I132449,I132475,I132483,I132500,I132287,I132540,I132548,I132281,I132296,I132593,I132610,I132636,I132284,I132658,I132675,I132692,I132299,I132723,I132740,I132290,I132771,I132293,I132305,I132302,I132860,I368344,I132886,I132903,I132925,I132942,I368341,I368338,I132959,I368326,I132985,I132993,I368350,I133019,I133027,I368335,I133044,I368329,I133084,I133092,I133137,I368332,I133154,I368347,I133180,I133202,I133219,I133236,I133267,I133284,I133315,I133404,I367188,I133430,I133447,I133469,I133486,I367185,I367182,I133503,I367170,I133529,I133537,I367194,I133563,I133571,I367179,I133588,I367173,I133628,I133636,I133681,I367176,I133698,I367191,I133724,I133746,I133763,I133780,I133811,I133828,I133859,I133948,I216553,I133974,I133991,I134013,I134030,I216574,I216565,I134047,I134073,I134081,I216559,I134107,I134115,I216556,I134132,I216550,I134172,I134180,I134225,I216562,I134242,I216571,I134268,I134290,I134307,I134324,I134355,I134372,I216568,I134403,I134492,I209039,I134518,I134535,I134557,I134574,I209060,I209051,I134591,I134617,I134625,I209045,I134651,I134659,I209042,I134676,I209036,I134716,I134724,I134769,I209048,I134786,I209057,I134812,I134834,I134851,I134868,I134899,I134916,I209054,I134947,I135036,I174937,I135062,I135079,I135028,I135101,I135118,I174934,I174955,I135135,I174958,I135161,I135169,I174943,I135195,I135203,I174946,I135220,I135007,I174949,I135260,I135268,I135001,I135016,I135313,I174940,I135330,I174952,I135356,I135004,I135378,I135395,I135412,I135019,I135443,I135460,I135010,I135491,I135013,I135025,I135022,I135580,I135606,I135623,I135572,I135645,I135662,I135679,I135705,I135713,I135739,I135747,I135764,I135551,I135804,I135812,I135545,I135560,I135857,I135874,I135900,I135548,I135922,I135939,I135956,I135563,I135987,I136004,I135554,I136035,I135557,I135569,I135566,I136124,I173781,I136150,I136167,I136116,I136189,I136206,I173778,I173799,I136223,I173802,I136249,I136257,I173787,I136283,I136291,I173790,I136308,I136095,I173793,I136348,I136356,I136089,I136104,I136401,I173784,I136418,I173796,I136444,I136092,I136466,I136483,I136500,I136107,I136531,I136548,I136098,I136579,I136101,I136113,I136110,I136668,I233018,I136694,I136711,I136660,I136733,I136750,I233012,I233009,I136767,I233024,I136793,I136801,I136827,I136835,I233006,I136852,I136639,I136892,I136900,I136633,I136648,I136945,I233021,I233015,I136962,I136988,I136636,I137010,I137027,I137044,I136651,I137075,I137092,I233027,I136642,I137123,I136645,I136657,I136654,I137212,I137238,I137255,I137204,I137277,I137294,I137311,I137337,I137345,I137371,I137379,I137396,I137183,I137436,I137444,I137177,I137192,I137489,I137506,I137532,I137180,I137554,I137571,I137588,I137195,I137619,I137636,I137186,I137667,I137189,I137201,I137198,I137756,I307911,I137782,I137799,I137748,I137821,I137838,I307923,I137855,I307914,I137881,I137889,I307932,I137915,I137923,I307908,I137940,I137727,I307926,I137980,I137988,I137721,I137736,I138033,I307920,I307917,I138050,I307929,I138076,I137724,I138098,I138115,I138132,I137739,I138163,I138180,I137730,I138211,I137733,I137745,I137742,I138300,I138326,I138343,I138365,I138382,I138399,I138425,I138433,I138459,I138467,I138484,I138524,I138532,I138577,I138594,I138620,I138642,I138659,I138676,I138707,I138724,I138755,I138844,I247774,I138870,I138887,I138909,I138926,I247768,I247765,I138943,I247780,I138969,I138977,I139003,I139011,I247762,I139028,I139068,I139076,I139121,I247777,I247771,I139138,I139164,I139186,I139203,I139220,I139251,I139268,I247783,I139299,I139388,I139414,I139431,I139380,I139453,I139470,I139487,I139513,I139521,I139547,I139555,I139572,I139359,I139612,I139620,I139353,I139368,I139665,I139682,I139708,I139356,I139730,I139747,I139764,I139371,I139795,I139812,I139362,I139843,I139365,I139377,I139374,I139932,I211351,I139958,I139975,I139997,I140014,I211372,I211363,I140031,I140057,I140065,I211357,I140091,I140099,I211354,I140116,I211348,I140156,I140164,I140209,I211360,I140226,I211369,I140252,I140274,I140291,I140308,I140339,I140356,I211366,I140387,I140476,I178983,I140502,I140519,I140468,I140541,I140558,I178980,I179001,I140575,I179004,I140601,I140609,I178989,I140635,I140643,I178992,I140660,I140447,I178995,I140700,I140708,I140441,I140456,I140753,I178986,I140770,I178998,I140796,I140444,I140818,I140835,I140852,I140459,I140883,I140900,I140450,I140931,I140453,I140465,I140462,I141017,I141043,I141060,I141009,I141091,I141099,I141116,I141133,I141150,I141167,I141184,I141201,I141006,I141232,I141249,I141266,I140991,I141003,I141311,I141328,I140997,I141359,I141376,I140985,I141407,I141424,I141441,I141467,I141475,I140994,I141506,I141523,I141000,I141554,I140988,I141612,I141638,I141655,I141604,I141686,I141694,I141711,I141728,I141745,I141762,I141779,I141796,I141601,I141827,I141844,I141861,I141586,I141598,I141906,I141923,I141592,I141954,I141971,I141580,I142002,I142019,I142036,I142062,I142070,I141589,I142101,I142118,I141595,I142149,I141583,I142207,I142233,I142250,I142281,I142289,I142306,I142323,I142340,I142357,I142374,I142391,I142422,I142439,I142456,I142501,I142518,I142549,I142566,I142597,I142614,I142631,I142657,I142665,I142696,I142713,I142744,I142802,I204999,I142828,I142845,I142794,I204993,I142876,I142884,I204990,I142901,I142918,I205002,I142935,I205005,I142952,I142969,I142986,I142791,I143017,I205014,I143034,I205008,I143051,I142776,I142788,I143096,I143113,I142782,I143144,I204996,I143161,I142770,I143192,I205011,I143209,I143226,I143252,I143260,I142779,I143291,I143308,I142785,I143339,I142773,I143397,I271254,I143423,I143440,I143389,I271242,I143471,I143479,I271239,I143496,I143513,I271251,I143530,I271248,I143547,I143564,I143581,I143386,I143612,I271257,I143629,I271260,I143646,I143371,I143383,I143691,I143708,I143377,I143739,I271263,I143756,I143365,I143787,I271266,I143804,I271245,I143821,I143847,I143855,I143374,I143886,I143903,I143380,I143934,I143368,I143992,I144018,I144035,I143984,I144066,I144074,I144091,I144108,I144125,I144142,I144159,I144176,I143981,I144207,I144224,I144241,I143966,I143978,I144286,I144303,I143972,I144334,I144351,I143960,I144382,I144399,I144416,I144442,I144450,I143969,I144481,I144498,I143975,I144529,I143963,I144587,I267378,I144613,I144630,I144579,I267366,I144661,I144669,I267363,I144686,I144703,I267375,I144720,I267372,I144737,I144754,I144771,I144576,I144802,I267381,I144819,I267384,I144836,I144561,I144573,I144881,I144898,I144567,I144929,I267387,I144946,I144555,I144977,I267390,I144994,I267369,I145011,I145037,I145045,I144564,I145076,I145093,I144570,I145124,I144558,I145182,I145208,I145225,I145174,I145256,I145264,I145281,I145298,I145315,I145332,I145349,I145366,I145171,I145397,I145414,I145431,I145156,I145168,I145476,I145493,I145162,I145524,I145541,I145150,I145572,I145589,I145606,I145632,I145640,I145159,I145671,I145688,I145165,I145719,I145153,I145777,I293815,I145803,I145820,I293818,I145851,I145859,I293821,I145876,I145893,I293833,I145910,I293824,I145927,I145944,I145961,I145992,I293830,I146009,I146026,I146071,I146088,I146119,I146136,I146167,I293827,I146184,I146201,I293836,I146227,I146235,I146266,I146283,I146314,I146372,I383643,I146398,I146415,I146364,I383649,I146446,I146454,I383664,I146471,I146488,I383655,I146505,I383652,I146522,I146539,I146556,I146361,I146587,I146604,I383667,I146621,I146346,I146358,I146666,I146683,I146352,I146714,I383661,I146731,I146340,I146762,I383646,I146779,I383658,I146796,I383670,I146822,I146830,I146349,I146861,I146878,I146355,I146909,I146343,I146967,I239339,I146993,I147010,I146959,I239336,I147041,I147049,I147066,I147083,I239333,I147100,I239348,I147117,I147134,I147151,I146956,I147182,I239342,I147199,I239330,I147216,I146941,I146953,I147261,I147278,I146947,I147309,I239351,I147326,I146935,I147357,I147374,I239345,I147391,I147417,I147425,I146944,I147456,I147473,I146950,I147504,I146938,I147562,I248298,I147588,I147605,I147554,I248295,I147636,I147644,I147661,I147678,I248292,I147695,I248307,I147712,I147729,I147746,I147551,I147777,I248301,I147794,I248289,I147811,I147536,I147548,I147856,I147873,I147542,I147904,I248310,I147921,I147530,I147952,I147969,I248304,I147986,I148012,I148020,I147539,I148051,I148068,I147545,I148099,I147533,I148157,I354590,I148183,I148200,I148149,I354605,I148231,I148239,I354614,I148256,I148273,I354593,I148290,I354599,I148307,I148324,I148341,I148146,I148372,I354611,I148389,I354608,I148406,I148131,I148143,I148451,I148468,I148137,I148499,I148516,I148125,I148547,I354602,I148564,I354596,I148581,I148607,I148615,I148134,I148646,I148663,I148140,I148694,I148128,I148752,I265440,I148778,I148795,I148744,I265428,I148826,I148834,I265425,I148851,I148868,I265437,I148885,I265434,I148902,I148919,I148936,I148741,I148967,I265443,I148984,I265446,I149001,I148726,I148738,I149046,I149063,I148732,I149094,I265449,I149111,I148720,I149142,I265452,I149159,I265431,I149176,I149202,I149210,I148729,I149241,I149258,I148735,I149289,I148723,I149347,I236177,I149373,I149390,I236174,I149421,I149429,I149446,I149463,I236171,I149480,I236186,I149497,I149514,I149531,I149562,I236180,I149579,I236168,I149596,I149641,I149658,I149689,I236189,I149706,I149737,I149754,I236183,I149771,I149797,I149805,I149836,I149853,I149884,I149942,I340872,I149968,I149985,I340854,I150016,I150024,I340860,I150041,I150058,I340875,I150075,I340866,I150092,I150109,I150126,I150157,I340878,I150174,I340857,I150191,I150236,I150253,I150284,I340863,I150301,I150332,I340869,I150349,I150366,I150392,I150400,I150431,I150448,I150479,I150537,I343166,I150563,I150580,I150529,I343181,I150611,I150619,I343190,I150636,I150653,I343169,I150670,I343175,I150687,I150704,I150721,I150526,I150752,I343187,I150769,I343184,I150786,I150511,I150523,I150831,I150848,I150517,I150879,I150896,I150505,I150927,I343178,I150944,I343172,I150961,I150987,I150995,I150514,I151026,I151043,I150520,I151074,I150508,I151132,I196329,I151158,I151175,I196323,I151206,I151214,I196320,I151231,I151248,I196332,I151265,I196335,I151282,I151299,I151316,I151347,I196344,I151364,I196338,I151381,I151426,I151443,I151474,I196326,I151491,I151522,I196341,I151539,I151556,I151582,I151590,I151621,I151638,I151669,I151727,I230907,I151753,I151770,I151719,I230904,I151801,I151809,I151826,I151843,I230901,I151860,I230916,I151877,I151894,I151911,I151716,I151942,I230910,I151959,I230898,I151976,I151701,I151713,I152021,I152038,I151707,I152069,I230919,I152086,I151695,I152117,I152134,I230913,I152151,I152177,I152185,I151704,I152216,I152233,I151710,I152264,I151698,I152322,I175515,I152348,I152365,I152314,I175527,I152396,I152404,I175512,I152421,I152438,I175530,I152455,I175521,I152472,I152489,I152506,I152311,I152537,I175533,I152554,I175536,I152571,I152296,I152308,I152616,I152633,I152302,I152664,I152681,I152290,I152712,I175524,I152729,I175518,I152746,I152772,I152780,I152299,I152811,I152828,I152305,I152859,I152293,I152917,I152943,I152960,I152991,I152999,I153016,I153033,I153050,I153067,I153084,I153101,I153132,I153149,I153166,I153211,I153228,I153259,I153276,I153307,I153324,I153341,I153367,I153375,I153406,I153423,I153454,I153512,I389593,I153538,I153555,I153504,I389599,I153586,I153594,I389614,I153611,I153628,I389605,I153645,I389602,I153662,I153679,I153696,I153501,I153727,I153744,I389617,I153761,I153486,I153498,I153806,I153823,I153492,I153854,I389611,I153871,I153480,I153902,I389596,I153919,I389608,I153936,I389620,I153962,I153970,I153489,I154001,I154018,I153495,I154049,I153483,I154107,I154133,I154150,I154181,I154189,I154206,I154223,I154240,I154257,I154274,I154291,I154322,I154339,I154356,I154401,I154418,I154449,I154466,I154497,I154514,I154531,I154557,I154565,I154596,I154613,I154644,I154702,I154728,I154745,I154776,I154784,I154801,I154818,I154835,I154852,I154869,I154886,I154917,I154934,I154951,I154996,I155013,I155044,I155061,I155092,I155109,I155126,I155152,I155160,I155191,I155208,I155239,I155297,I217137,I155323,I155340,I217131,I155371,I155379,I217128,I155396,I155413,I217140,I155430,I217143,I155447,I155464,I155481,I155512,I217152,I155529,I217146,I155546,I155591,I155608,I155639,I217134,I155656,I155687,I217149,I155704,I155721,I155747,I155755,I155786,I155803,I155834,I155892,I336230,I155918,I155926,I336236,I155952,I155960,I155977,I336233,I155994,I156011,I336251,I156028,I156059,I156076,I156093,I336254,I156110,I156155,I156200,I336239,I156217,I156234,I156265,I336245,I156282,I336242,I156299,I336248,I156325,I156333,I156378,I156395,I156412,I156470,I351888,I156496,I156504,I351882,I156530,I156538,I351891,I156555,I351870,I156572,I156589,I351879,I156606,I156456,I156637,I156654,I156671,I351894,I156688,I351873,I156453,I156444,I156733,I156447,I156441,I156778,I351876,I156795,I156812,I156450,I156843,I351885,I156860,I156877,I156903,I156911,I156438,I156462,I156956,I156973,I156990,I156459,I157048,I157074,I157082,I157108,I157116,I157133,I157150,I157167,I157184,I157034,I157215,I157232,I157249,I157266,I157031,I157022,I157311,I157025,I157019,I157356,I157373,I157390,I157028,I157421,I157438,I157455,I157481,I157489,I157016,I157040,I157534,I157551,I157568,I157037,I157626,I391973,I157652,I157660,I157686,I157694,I391997,I157711,I391979,I157728,I157745,I391994,I157762,I157612,I157793,I157810,I157827,I391976,I157844,I391985,I157609,I157600,I157889,I157603,I157597,I157934,I391982,I157951,I157968,I157606,I157999,I391991,I158016,I392000,I158033,I391988,I158059,I158067,I157594,I157618,I158112,I158129,I158146,I157615,I158204,I158230,I158238,I158264,I158272,I158289,I158306,I158323,I158340,I158190,I158371,I158388,I158405,I158422,I158187,I158178,I158467,I158181,I158175,I158512,I158529,I158546,I158184,I158577,I158594,I158611,I158637,I158645,I158172,I158196,I158690,I158707,I158724,I158193,I158782,I246714,I158808,I158816,I158842,I158850,I246711,I158867,I246726,I158884,I158901,I246720,I158918,I158949,I158966,I158983,I246717,I159000,I246708,I159045,I159090,I246729,I159107,I159124,I159155,I159172,I159189,I246723,I159215,I159223,I159268,I159285,I159302,I159360,I318890,I159386,I159394,I318896,I159420,I159428,I159445,I318893,I159462,I159479,I318911,I159496,I159527,I159544,I159561,I318914,I159578,I159623,I159668,I318899,I159685,I159702,I159733,I318905,I159750,I318902,I159767,I318908,I159793,I159801,I159846,I159863,I159880,I159938,I372338,I159964,I159972,I159998,I160006,I372362,I160023,I372344,I160040,I160057,I372359,I160074,I159924,I160105,I160122,I160139,I372341,I160156,I372350,I159921,I159912,I160201,I159915,I159909,I160246,I372347,I160263,I160280,I159918,I160311,I372356,I160328,I372365,I160345,I372353,I160371,I160379,I159906,I159930,I160424,I160441,I160458,I159927,I160516,I160542,I160550,I160576,I160584,I160601,I160618,I160635,I160652,I160683,I160700,I160717,I160734,I160779,I160824,I160841,I160858,I160889,I160906,I160923,I160949,I160957,I161002,I161019,I161036,I161094,I187650,I161120,I161128,I187662,I161154,I161162,I187653,I161179,I187656,I161196,I161213,I187659,I161230,I161080,I161261,I161278,I161295,I161312,I187665,I161077,I161068,I161357,I161071,I161065,I161402,I187671,I161419,I161436,I161074,I161467,I161484,I187668,I161501,I187674,I161527,I161535,I161062,I161086,I161580,I161597,I161614,I161083,I161672,I384238,I161698,I161706,I161732,I161740,I384262,I161757,I384244,I161774,I161791,I384259,I161808,I161658,I161839,I161856,I161873,I384241,I161890,I384250,I161655,I161646,I161935,I161649,I161643,I161980,I384247,I161997,I162014,I161652,I162045,I384256,I162062,I384265,I162079,I384253,I162105,I162113,I161640,I161664,I162158,I162175,I162192,I161661,I162250,I162276,I162284,I162310,I162318,I162335,I162352,I162369,I162386,I162417,I162434,I162451,I162468,I162513,I162558,I162575,I162592,I162623,I162640,I162657,I162683,I162691,I162736,I162753,I162770,I162828,I379478,I162854,I162862,I162888,I162896,I379502,I162913,I379484,I162930,I162947,I379499,I162964,I162814,I162995,I163012,I163029,I379481,I163046,I379490,I162811,I162802,I163091,I162805,I162799,I163136,I379487,I163153,I163170,I162808,I163201,I379496,I163218,I379505,I163235,I379493,I163261,I163269,I162796,I162820,I163314,I163331,I163348,I162817,I163406,I163432,I163440,I163466,I163474,I163491,I163508,I163525,I163542,I163392,I163573,I163590,I163607,I163624,I163389,I163380,I163669,I163383,I163377,I163714,I163731,I163748,I163386,I163779,I163796,I163813,I163839,I163847,I163374,I163398,I163892,I163909,I163926,I163395,I163984,I164010,I164018,I164044,I164052,I164069,I164086,I164103,I164120,I163970,I164151,I164168,I164185,I164202,I163967,I163958,I164247,I163961,I163955,I164292,I164309,I164326,I163964,I164357,I164374,I164391,I164417,I164425,I163952,I163976,I164470,I164487,I164504,I163973,I164562,I164588,I164596,I164622,I164630,I164647,I164664,I164681,I164698,I164548,I164729,I164746,I164763,I164780,I164545,I164536,I164825,I164539,I164533,I164870,I164887,I164904,I164542,I164935,I164952,I164969,I164995,I165003,I164530,I164554,I165048,I165065,I165082,I164551,I165140,I165166,I165174,I165200,I165208,I165225,I165242,I165259,I165276,I165307,I165324,I165341,I165358,I165403,I165448,I165465,I165482,I165513,I165530,I165547,I165573,I165581,I165626,I165643,I165660,I165718,I165744,I165752,I165778,I165786,I165803,I165820,I165837,I165854,I165704,I165885,I165902,I165919,I165936,I165701,I165692,I165981,I165695,I165689,I166026,I166043,I166060,I165698,I166091,I166108,I166125,I166151,I166159,I165686,I165710,I166204,I166221,I166238,I165707,I166296,I364870,I166322,I166330,I364882,I166356,I166364,I364873,I166381,I364861,I166398,I166415,I364858,I166432,I166282,I166463,I166480,I166497,I364864,I166514,I166279,I166270,I166559,I166273,I166267,I166604,I364879,I166621,I166638,I166276,I166669,I364867,I166686,I166703,I364876,I166729,I166737,I166264,I166288,I166782,I166799,I166816,I166285,I166874,I166900,I166908,I166934,I166942,I166959,I166976,I166993,I167010,I166860,I167041,I167058,I167075,I167092,I166857,I166848,I167137,I166851,I166845,I167182,I167199,I167216,I166854,I167247,I167264,I167281,I167307,I167315,I166842,I166866,I167360,I167377,I167394,I166863,I167452,I268015,I167478,I167486,I268012,I167512,I167520,I268009,I167537,I268036,I167554,I167571,I268024,I167588,I167438,I167619,I167636,I167653,I268030,I167670,I268021,I167435,I167426,I167715,I167429,I167423,I167760,I268018,I167777,I167794,I167432,I167825,I268033,I167842,I268027,I167859,I167885,I167893,I167420,I167444,I167938,I167955,I167972,I167441,I168030,I287395,I168056,I168064,I287392,I168090,I168098,I287389,I168115,I287416,I168132,I168149,I287404,I168166,I168197,I168214,I168231,I287410,I168248,I287401,I168293,I168338,I287398,I168355,I168372,I168403,I287413,I168420,I287407,I168437,I168463,I168471,I168516,I168533,I168550,I168608,I205568,I168634,I168642,I205580,I168668,I168676,I205571,I168693,I205574,I168710,I168727,I205577,I168744,I168594,I168775,I168792,I168809,I168826,I205583,I168591,I168582,I168871,I168585,I168579,I168916,I205589,I168933,I168950,I168588,I168981,I168998,I205586,I169015,I205592,I169041,I169049,I168576,I168600,I169094,I169111,I169128,I168597,I169186,I366604,I169212,I169220,I366616,I169246,I169254,I366607,I169271,I366595,I169288,I169305,I366592,I169322,I169172,I169353,I169370,I169387,I366598,I169404,I169169,I169160,I169449,I169163,I169157,I169494,I366613,I169511,I169528,I169166,I169559,I366601,I169576,I169593,I366610,I169619,I169627,I169154,I169178,I169672,I169689,I169706,I169175,I169764,I169790,I169798,I169824,I169832,I169849,I169866,I169883,I169900,I169750,I169931,I169948,I169965,I169982,I169747,I169738,I170027,I169741,I169735,I170072,I170089,I170106,I169744,I170137,I170154,I170171,I170197,I170205,I169732,I169756,I170250,I170267,I170284,I169753,I170342,I170368,I170376,I170402,I170410,I170427,I170444,I170461,I170478,I170509,I170526,I170543,I170560,I170605,I170650,I170667,I170684,I170715,I170732,I170749,I170775,I170783,I170828,I170845,I170862,I170920,I170946,I170954,I170980,I170988,I171005,I171022,I171039,I171056,I170906,I171087,I171104,I171121,I171138,I170903,I170894,I171183,I170897,I170891,I171228,I171245,I171262,I170900,I171293,I171310,I171327,I171353,I171361,I170888,I170912,I171406,I171423,I171440,I170909,I171498,I171524,I171532,I171558,I171566,I171583,I171600,I171617,I171634,I171665,I171682,I171699,I171716,I171761,I171806,I171823,I171840,I171871,I171888,I171905,I171931,I171939,I171984,I172001,I172018,I172076,I329872,I172102,I172110,I329878,I172136,I172144,I172161,I329875,I172178,I172195,I329893,I172212,I172062,I172243,I172260,I172277,I329896,I172294,I172059,I172050,I172339,I172053,I172047,I172384,I329881,I172401,I172418,I172056,I172449,I329887,I172466,I329884,I172483,I329890,I172509,I172517,I172044,I172068,I172562,I172579,I172596,I172065,I172654,I250930,I172680,I172688,I172714,I172722,I250927,I172739,I250942,I172756,I172773,I250936,I172790,I172640,I172821,I172838,I172855,I250933,I172872,I250924,I172637,I172628,I172917,I172631,I172625,I172962,I250945,I172979,I172996,I172634,I173027,I173044,I173061,I250939,I173087,I173095,I172622,I172646,I173140,I173157,I173174,I172643,I173232,I339120,I173258,I173266,I339126,I173292,I173300,I173317,I339123,I173334,I173351,I339141,I173368,I173218,I173399,I173416,I173433,I339144,I173450,I173215,I173206,I173495,I173209,I173203,I173540,I339129,I173557,I173574,I173212,I173605,I339135,I173622,I339132,I173639,I339138,I173665,I173673,I173200,I173224,I173718,I173735,I173752,I173221,I173810,I353520,I173836,I173844,I353514,I173870,I173878,I353523,I173895,I353502,I173912,I173929,I353511,I173946,I173977,I173994,I174011,I353526,I174028,I353505,I174073,I174118,I353508,I174135,I174152,I174183,I353517,I174200,I174217,I174243,I174251,I174296,I174313,I174330,I174388,I214238,I174414,I174422,I214250,I174448,I174456,I214241,I174473,I214244,I174490,I174507,I214247,I174524,I174374,I174555,I174572,I174589,I174606,I214253,I174371,I174362,I174651,I174365,I174359,I174696,I214259,I174713,I174730,I174368,I174761,I174778,I214256,I174795,I214262,I174821,I174829,I174356,I174380,I174874,I174891,I174908,I174377,I174966,I174992,I175000,I175026,I175034,I175051,I175068,I175085,I175102,I175133,I175150,I175167,I175184,I175229,I175274,I175291,I175308,I175339,I175356,I175373,I175399,I175407,I175452,I175469,I175486,I175544,I175570,I175578,I175604,I175612,I175629,I175646,I175663,I175680,I175711,I175728,I175745,I175762,I175807,I175852,I175869,I175886,I175917,I175934,I175951,I175977,I175985,I176030,I176047,I176064,I176122,I220596,I176148,I176156,I220608,I176182,I176190,I220599,I176207,I220602,I176224,I176241,I220605,I176258,I176289,I176306,I176323,I176340,I220611,I176385,I176430,I220617,I176447,I176464,I176495,I176512,I220614,I176529,I220620,I176555,I176563,I176608,I176625,I176642,I176700,I277059,I176726,I176734,I277056,I176760,I176768,I277053,I176785,I277080,I176802,I176819,I277068,I176836,I176686,I176867,I176884,I176901,I277074,I176918,I277065,I176683,I176674,I176963,I176677,I176671,I177008,I277062,I177025,I177042,I176680,I177073,I277077,I177090,I277071,I177107,I177133,I177141,I176668,I176692,I177186,I177203,I177220,I176689,I177278,I177304,I177312,I177338,I177346,I177363,I177380,I177397,I177414,I177264,I177445,I177462,I177479,I177496,I177261,I177252,I177541,I177255,I177249,I177586,I177603,I177620,I177258,I177651,I177668,I177685,I177711,I177719,I177246,I177270,I177764,I177781,I177798,I177267,I177856,I177882,I177890,I177916,I177924,I177941,I177958,I177975,I177992,I178023,I178040,I178057,I178074,I178119,I178164,I178181,I178198,I178229,I178246,I178263,I178289,I178297,I178342,I178359,I178376,I178434,I178460,I178468,I178494,I178502,I178519,I178536,I178553,I178570,I178601,I178618,I178635,I178652,I178697,I178742,I178759,I178776,I178807,I178824,I178841,I178867,I178875,I178920,I178937,I178954,I179012,I354064,I179038,I179046,I354058,I179072,I179080,I354067,I179097,I354046,I179114,I179131,I354055,I179148,I179179,I179196,I179213,I354070,I179230,I354049,I179275,I179320,I354052,I179337,I179354,I179385,I354061,I179402,I179419,I179445,I179453,I179498,I179515,I179532,I179590,I179616,I179624,I179650,I179658,I179675,I179692,I179709,I179726,I179757,I179774,I179791,I179808,I179853,I179898,I179915,I179932,I179963,I179980,I179997,I180023,I180031,I180076,I180093,I180110,I180168,I241444,I180194,I180202,I180228,I180236,I241441,I180253,I241456,I180270,I180287,I241450,I180304,I180154,I180335,I180352,I180369,I241447,I180386,I241438,I180151,I180142,I180431,I180145,I180139,I180476,I241459,I180493,I180510,I180148,I180541,I180558,I180575,I241453,I180601,I180609,I180136,I180160,I180654,I180671,I180688,I180157,I180746,I180772,I180780,I180806,I180814,I180831,I180848,I180865,I180882,I180913,I180930,I180947,I180964,I181009,I181054,I181071,I181088,I181119,I181136,I181153,I181179,I181187,I181232,I181249,I181266,I181324,I181350,I181358,I181375,I181392,I181418,I181426,I181452,I181460,I181477,I181494,I181511,I181551,I181559,I181576,I181593,I181610,I181641,I181658,I181684,I181692,I181723,I181754,I181771,I181802,I181902,I181928,I181936,I181953,I181970,I181996,I182004,I182030,I182038,I182055,I182072,I182089,I182129,I182137,I182154,I182171,I182188,I182219,I182236,I182262,I182270,I182301,I182332,I182349,I182380,I182480,I182506,I182514,I182531,I182548,I182574,I182582,I182608,I182616,I182633,I182650,I182667,I182463,I182707,I182715,I182732,I182749,I182766,I182466,I182797,I182814,I182840,I182848,I182448,I182879,I182457,I182910,I182927,I182469,I182958,I182460,I182451,I182454,I182472,I183058,I183084,I183092,I183109,I183126,I183152,I183160,I183186,I183194,I183211,I183228,I183245,I183285,I183293,I183310,I183327,I183344,I183375,I183392,I183418,I183426,I183457,I183488,I183505,I183536,I183636,I183662,I183670,I183687,I183704,I183730,I183738,I183764,I183772,I183789,I183806,I183823,I183619,I183863,I183871,I183888,I183905,I183922,I183622,I183953,I183970,I183996,I184004,I183604,I184035,I183613,I184066,I184083,I183625,I184114,I183616,I183607,I183610,I183628,I184214,I184240,I184248,I184265,I184282,I184308,I184316,I184342,I184350,I184367,I184384,I184401,I184197,I184441,I184449,I184466,I184483,I184500,I184200,I184531,I184548,I184574,I184582,I184182,I184613,I184191,I184644,I184661,I184203,I184692,I184194,I184185,I184188,I184206,I184792,I184818,I184826,I184843,I184860,I184886,I184894,I184920,I184928,I184945,I184962,I184979,I184775,I185019,I185027,I185044,I185061,I185078,I184778,I185109,I185126,I185152,I185160,I184760,I185191,I184769,I185222,I185239,I184781,I185270,I184772,I184763,I184766,I184784,I185370,I185396,I185404,I185421,I185438,I185464,I185472,I185498,I185506,I185523,I185540,I185557,I185353,I185597,I185605,I185622,I185639,I185656,I185356,I185687,I185704,I185730,I185738,I185338,I185769,I185347,I185800,I185817,I185359,I185848,I185350,I185341,I185344,I185362,I185948,I298309,I185974,I185982,I185999,I298306,I298324,I186016,I298321,I186042,I186050,I298303,I186076,I186084,I186101,I186118,I186135,I298315,I186175,I186183,I186200,I186217,I186234,I186265,I298318,I186282,I186308,I186316,I186347,I186378,I186395,I186426,I298312,I186526,I374150,I186552,I186560,I186577,I374135,I374123,I186594,I374138,I186620,I186628,I374141,I186654,I186662,I186679,I186696,I186713,I186509,I374129,I186753,I186761,I186778,I186795,I186812,I186512,I186843,I374126,I374132,I186860,I374147,I186886,I186894,I186494,I186925,I186503,I186956,I186973,I186515,I187004,I374144,I186506,I186497,I186500,I186518,I187104,I381885,I187130,I187138,I187155,I381870,I381858,I187172,I381873,I187198,I187206,I381876,I187232,I187240,I187257,I187274,I187291,I187087,I381864,I187331,I187339,I187356,I187373,I187390,I187090,I187421,I381861,I381867,I187438,I381882,I187464,I187472,I187072,I187503,I187081,I187534,I187551,I187093,I187582,I381879,I187084,I187075,I187078,I187096,I187682,I187708,I187716,I187733,I187750,I187776,I187784,I187810,I187818,I187835,I187852,I187869,I187909,I187917,I187934,I187951,I187968,I187999,I188016,I188042,I188050,I188081,I188112,I188129,I188160,I188260,I255113,I188286,I188294,I188311,I255089,I255104,I188328,I255116,I188354,I188362,I255101,I255092,I188388,I188396,I188413,I188430,I188447,I188487,I188495,I188512,I188529,I188546,I188577,I255107,I255098,I188594,I255110,I188620,I188628,I188659,I188690,I188707,I188738,I255095,I188838,I231967,I188864,I188872,I188889,I231955,I231973,I188906,I231970,I188932,I188940,I231961,I231958,I188966,I188974,I188991,I189008,I189025,I188821,I231952,I189065,I189073,I189090,I189107,I189124,I188824,I189155,I189172,I189198,I189206,I188806,I189237,I188815,I189268,I189285,I188827,I189316,I231964,I188818,I188809,I188812,I188830,I189416,I189442,I189450,I189467,I189484,I189510,I189518,I189544,I189552,I189569,I189586,I189603,I189643,I189651,I189668,I189685,I189702,I189733,I189750,I189776,I189784,I189815,I189846,I189863,I189894,I189994,I190020,I190028,I190045,I190062,I190088,I190096,I190122,I190130,I190147,I190164,I190181,I189977,I190221,I190229,I190246,I190263,I190280,I189980,I190311,I190328,I190354,I190362,I189962,I190393,I189971,I190424,I190441,I189983,I190472,I189974,I189965,I189968,I189986,I190572,I190598,I190606,I190623,I190640,I190666,I190674,I190700,I190708,I190725,I190742,I190759,I190555,I190799,I190807,I190824,I190841,I190858,I190558,I190889,I190906,I190932,I190940,I190540,I190971,I190549,I191002,I191019,I190561,I191050,I190552,I190543,I190546,I190564,I191150,I257697,I191176,I191184,I191201,I257673,I257688,I191218,I257700,I191244,I191252,I257685,I257676,I191278,I191286,I191303,I191320,I191337,I191133,I191377,I191385,I191402,I191419,I191436,I191136,I191467,I257691,I257682,I191484,I257694,I191510,I191518,I191118,I191549,I191127,I191580,I191597,I191139,I191628,I257679,I191130,I191121,I191124,I191142,I191728,I191754,I191762,I191779,I191796,I191822,I191830,I191856,I191864,I191881,I191898,I191915,I191711,I191955,I191963,I191980,I191997,I192014,I191714,I192045,I192062,I192088,I192096,I191696,I192127,I191705,I192158,I192175,I191717,I192206,I191708,I191699,I191702,I191720,I192306,I192332,I192340,I192357,I192374,I192400,I192408,I192434,I192442,I192459,I192476,I192493,I192289,I192533,I192541,I192558,I192575,I192592,I192292,I192623,I192640,I192666,I192674,I192274,I192705,I192283,I192736,I192753,I192295,I192784,I192286,I192277,I192280,I192298,I192884,I192910,I192918,I192935,I192952,I192978,I192986,I193012,I193020,I193037,I193054,I193071,I192867,I193111,I193119,I193136,I193153,I193170,I192870,I193201,I193218,I193244,I193252,I192852,I193283,I192861,I193314,I193331,I192873,I193362,I192864,I192855,I192858,I192876,I193462,I309082,I193488,I193496,I193513,I309064,I309076,I193530,I309079,I193556,I193564,I309073,I309070,I193590,I193598,I193615,I193632,I193649,I309088,I193689,I193697,I193714,I193731,I193748,I193779,I309067,I193796,I193822,I193830,I193861,I193892,I193909,I193940,I309085,I194040,I324688,I194066,I194074,I194091,I324670,I324682,I194108,I324685,I194134,I194142,I324679,I324676,I194168,I194176,I194193,I194210,I194227,I324694,I194267,I194275,I194292,I194309,I194326,I194357,I324673,I194374,I194400,I194408,I194439,I194470,I194487,I194518,I324691,I194618,I373555,I194644,I194652,I194669,I373540,I373528,I194686,I373543,I194712,I194720,I373546,I194746,I194754,I194771,I194788,I194805,I194601,I373534,I194845,I194853,I194870,I194887,I194904,I194604,I194935,I373531,I373537,I194952,I373552,I194978,I194986,I194586,I195017,I194595,I195048,I195065,I194607,I195096,I373549,I194598,I194589,I194592,I194610,I195196,I350238,I195222,I195230,I195247,I350241,I350250,I195264,I350253,I195290,I195298,I350262,I350244,I195324,I195332,I195349,I195366,I195383,I195423,I195431,I195448,I195465,I195482,I195513,I350259,I195530,I350256,I195556,I195564,I195595,I195626,I195643,I195674,I350247,I195774,I195800,I195808,I195825,I195842,I195868,I195876,I195902,I195910,I195927,I195944,I195961,I196001,I196009,I196026,I196043,I196060,I196091,I196108,I196134,I196142,I196173,I196204,I196221,I196252,I196352,I313706,I196378,I196386,I196403,I313688,I313700,I196420,I313703,I196446,I196454,I313697,I313694,I196480,I196488,I196505,I196522,I196539,I313712,I196579,I196587,I196604,I196621,I196638,I196669,I313691,I196686,I196712,I196720,I196751,I196782,I196799,I196830,I313709,I196930,I323532,I196956,I196964,I196981,I323514,I323526,I196998,I323529,I197024,I197032,I323523,I323520,I197058,I197066,I197083,I197100,I197117,I196913,I323538,I197157,I197165,I197182,I197199,I197216,I196916,I197247,I323517,I197264,I197290,I197298,I196898,I197329,I196907,I197360,I197377,I196919,I197408,I323535,I196910,I196901,I196904,I196922,I197508,I197534,I197542,I197559,I197576,I197602,I197610,I197636,I197644,I197661,I197678,I197695,I197735,I197743,I197760,I197777,I197794,I197825,I197842,I197868,I197876,I197907,I197938,I197955,I197986,I198086,I364280,I198112,I198120,I198137,I364304,I364286,I198154,I364292,I198180,I198188,I364298,I364283,I198214,I198222,I198239,I198256,I198273,I198069,I364295,I198313,I198321,I198338,I198355,I198372,I198072,I198403,I364301,I364289,I198420,I198446,I198454,I198054,I198485,I198063,I198516,I198533,I198075,I198564,I198066,I198057,I198060,I198078,I198664,I260281,I198690,I198698,I198715,I260257,I260272,I198732,I260284,I198758,I198766,I260269,I260260,I198792,I198800,I198817,I198834,I198851,I198647,I198891,I198899,I198916,I198933,I198950,I198650,I198981,I260275,I260266,I198998,I260278,I199024,I199032,I198632,I199063,I198641,I199094,I199111,I198653,I199142,I260263,I198644,I198635,I198638,I198656,I199242,I199268,I199276,I199293,I199310,I199336,I199344,I199370,I199378,I199395,I199412,I199429,I199469,I199477,I199494,I199511,I199528,I199559,I199576,I199602,I199610,I199641,I199672,I199689,I199720,I199820,I199846,I199854,I199871,I199888,I199914,I199922,I199948,I199956,I199973,I199990,I200007,I199803,I200047,I200055,I200072,I200089,I200106,I199806,I200137,I200154,I200180,I200188,I199788,I200219,I199797,I200250,I200267,I199809,I200298,I199800,I199791,I199794,I199812,I200398,I200424,I200432,I200449,I200466,I200492,I200500,I200526,I200534,I200551,I200568,I200585,I200625,I200633,I200650,I200667,I200684,I200715,I200732,I200758,I200766,I200797,I200828,I200845,I200876,I200976,I201002,I201010,I201027,I201044,I201070,I201078,I201104,I201112,I201129,I201146,I201163,I201203,I201211,I201228,I201245,I201262,I201293,I201310,I201336,I201344,I201375,I201406,I201423,I201454,I201554,I201580,I201588,I201605,I201622,I201648,I201656,I201682,I201690,I201707,I201724,I201741,I201781,I201789,I201806,I201823,I201840,I201871,I201888,I201914,I201922,I201953,I201984,I202001,I202032,I202132,I202158,I202166,I202183,I202200,I202226,I202234,I202260,I202268,I202285,I202302,I202319,I202359,I202367,I202384,I202401,I202418,I202449,I202466,I202492,I202500,I202531,I202562,I202579,I202610,I202710,I202736,I202744,I202761,I202778,I202804,I202812,I202838,I202846,I202863,I202880,I202897,I202937,I202945,I202962,I202979,I202996,I203027,I203044,I203070,I203078,I203109,I203140,I203157,I203188,I203288,I203314,I203322,I203339,I203356,I203382,I203390,I203416,I203424,I203441,I203458,I203475,I203515,I203523,I203540,I203557,I203574,I203605,I203622,I203648,I203656,I203687,I203718,I203735,I203766,I203866,I203892,I203900,I203917,I203934,I203960,I203968,I203994,I204002,I204019,I204036,I204053,I203849,I204093,I204101,I204118,I204135,I204152,I203852,I204183,I204200,I204226,I204234,I203834,I204265,I203843,I204296,I204313,I203855,I204344,I203846,I203837,I203840,I203858,I204444,I204470,I204478,I204495,I204512,I204538,I204546,I204572,I204580,I204597,I204614,I204631,I204671,I204679,I204696,I204713,I204730,I204761,I204778,I204804,I204812,I204843,I204874,I204891,I204922,I205022,I286767,I205048,I205056,I205073,I286743,I286758,I205090,I286770,I205116,I205124,I286755,I286746,I205150,I205158,I205175,I205192,I205209,I205249,I205257,I205274,I205291,I205308,I205339,I286761,I286752,I205356,I286764,I205382,I205390,I205421,I205452,I205469,I205500,I286749,I205600,I264803,I205626,I205634,I205651,I264779,I264794,I205668,I264806,I205694,I205702,I264791,I264782,I205728,I205736,I205753,I205770,I205787,I205827,I205835,I205852,I205869,I205886,I205917,I264797,I264788,I205934,I264800,I205960,I205968,I205999,I206030,I206047,I206078,I264785,I206178,I206204,I206212,I206229,I206246,I206272,I206280,I206306,I206314,I206331,I206348,I206365,I206161,I206405,I206413,I206430,I206447,I206464,I206164,I206495,I206512,I206538,I206546,I206146,I206577,I206155,I206608,I206625,I206167,I206656,I206158,I206149,I206152,I206170,I206756,I258989,I206782,I206790,I206807,I258965,I258980,I206824,I258992,I206850,I206858,I258977,I258968,I206884,I206892,I206909,I206926,I206943,I206983,I206991,I207008,I207025,I207042,I207073,I258983,I258974,I207090,I258986,I207116,I207124,I207155,I207186,I207203,I207234,I258971,I207334,I333936,I207360,I207368,I207385,I333918,I333930,I207402,I333933,I207428,I207436,I333927,I333924,I207462,I207470,I207487,I207504,I207521,I207317,I333942,I207561,I207569,I207586,I207603,I207620,I207320,I207651,I333921,I207668,I207694,I207702,I207302,I207733,I207311,I207764,I207781,I207323,I207812,I333939,I207314,I207305,I207308,I207326,I207912,I279661,I207938,I207946,I207963,I279637,I279652,I207980,I279664,I208006,I208014,I279649,I279640,I208040,I208048,I208065,I208082,I208099,I208139,I208147,I208164,I208181,I208198,I208229,I279655,I279646,I208246,I279658,I208272,I208280,I208311,I208342,I208359,I208390,I279643,I208490,I342028,I208516,I208524,I208541,I342010,I342022,I208558,I342025,I208584,I208592,I342019,I342016,I208618,I208626,I208643,I208660,I208677,I342034,I208717,I208725,I208742,I208759,I208776,I208807,I342013,I208824,I208850,I208858,I208889,I208920,I208937,I208968,I342031,I209068,I209094,I209102,I209119,I209136,I209162,I209170,I209196,I209204,I209221,I209238,I209255,I209295,I209303,I209320,I209337,I209354,I209385,I209402,I209428,I209436,I209467,I209498,I209515,I209546,I209646,I317174,I209672,I209680,I209697,I317156,I317168,I209714,I317171,I209740,I209748,I317165,I317162,I209774,I209782,I209799,I209816,I209833,I317180,I209873,I209881,I209898,I209915,I209932,I209963,I317159,I209980,I210006,I210014,I210045,I210076,I210093,I210124,I317177,I210224,I210250,I210258,I210275,I210292,I210318,I210326,I210352,I210360,I210377,I210394,I210411,I210451,I210459,I210476,I210493,I210510,I210541,I210558,I210584,I210592,I210623,I210654,I210671,I210702,I210802,I275139,I210828,I210836,I210853,I275115,I275130,I210870,I275142,I210896,I210904,I275127,I275118,I210930,I210938,I210955,I210972,I210989,I211029,I211037,I211054,I211071,I211088,I211119,I275133,I275124,I211136,I275136,I211162,I211170,I211201,I211232,I211249,I211280,I275121,I211380,I211406,I211414,I211431,I211448,I211474,I211482,I211508,I211516,I211533,I211550,I211567,I211607,I211615,I211632,I211649,I211666,I211697,I211714,I211740,I211748,I211779,I211810,I211827,I211858,I211958,I211984,I211992,I212009,I212026,I212052,I212060,I212086,I212094,I212111,I212128,I212145,I212185,I212193,I212210,I212227,I212244,I212275,I212292,I212318,I212326,I212357,I212388,I212405,I212436,I212536,I247250,I212562,I212570,I212587,I247238,I247256,I212604,I247253,I212630,I212638,I247244,I247241,I212664,I212672,I212689,I212706,I212723,I247235,I212763,I212771,I212788,I212805,I212822,I212853,I212870,I212896,I212904,I212935,I212966,I212983,I213014,I247247,I213114,I259635,I213140,I213148,I213165,I259611,I259626,I213182,I259638,I213208,I213216,I259623,I259614,I213242,I213250,I213267,I213284,I213301,I213097,I213341,I213349,I213366,I213383,I213400,I213100,I213431,I259629,I259620,I213448,I259632,I213474,I213482,I213082,I213513,I213091,I213544,I213561,I213103,I213592,I259617,I213094,I213085,I213088,I213106,I213692,I213718,I213726,I213743,I213760,I213786,I213794,I213820,I213828,I213845,I213862,I213879,I213675,I213919,I213927,I213944,I213961,I213978,I213678,I214009,I214026,I214052,I214060,I213660,I214091,I213669,I214122,I214139,I213681,I214170,I213672,I213663,I213666,I213684,I214270,I214296,I214304,I214321,I214338,I214364,I214372,I214398,I214406,I214423,I214440,I214457,I214497,I214505,I214522,I214539,I214556,I214587,I214604,I214630,I214638,I214669,I214700,I214717,I214748,I214848,I380100,I214874,I214882,I214899,I380085,I380073,I214916,I380088,I214942,I214950,I380091,I214976,I214984,I215001,I215018,I215035,I214831,I380079,I215075,I215083,I215100,I215117,I215134,I214834,I215165,I380076,I380082,I215182,I380097,I215208,I215216,I214816,I215247,I214825,I215278,I215295,I214837,I215326,I380094,I214828,I214819,I214822,I214840,I215426,I215452,I215460,I215477,I215494,I215520,I215528,I215554,I215562,I215579,I215596,I215613,I215653,I215661,I215678,I215695,I215712,I215743,I215760,I215786,I215794,I215825,I215856,I215873,I215904,I216004,I216030,I216038,I216055,I216072,I216098,I216106,I216132,I216140,I216157,I216174,I216191,I215987,I216231,I216239,I216256,I216273,I216290,I215990,I216321,I216338,I216364,I216372,I215972,I216403,I215981,I216434,I216451,I215993,I216482,I215984,I215975,I215978,I215996,I216582,I216608,I216616,I216633,I216650,I216676,I216684,I216710,I216718,I216735,I216752,I216769,I216809,I216817,I216834,I216851,I216868,I216899,I216916,I216942,I216950,I216981,I217012,I217029,I217060,I217160,I253175,I217186,I217194,I217211,I253151,I253166,I217228,I253178,I217254,I217262,I253163,I253154,I217288,I217296,I217313,I217330,I217347,I217387,I217395,I217412,I217429,I217446,I217477,I253169,I253160,I217494,I253172,I217520,I217528,I217559,I217590,I217607,I217638,I253157,I217738,I377720,I217764,I217772,I217789,I377705,I377693,I217806,I377708,I217832,I217840,I377711,I217866,I217874,I217891,I217908,I217925,I377699,I217965,I217973,I217990,I218007,I218024,I218055,I377696,I377702,I218072,I377717,I218098,I218106,I218137,I218168,I218185,I218216,I377714,I218316,I370602,I218342,I218350,I218367,I370590,I370608,I218384,I370599,I218410,I218418,I370614,I370611,I218444,I218452,I218469,I218486,I218503,I218299,I370593,I218543,I218551,I218568,I218585,I218602,I218302,I218633,I370587,I218650,I370596,I218676,I218684,I218284,I218715,I218293,I218746,I218763,I218305,I218794,I370605,I218296,I218287,I218290,I218308,I218894,I335092,I218920,I218928,I218945,I335074,I335086,I218962,I335089,I218988,I218996,I335083,I335080,I219022,I219030,I219047,I219064,I219081,I335098,I219121,I219129,I219146,I219163,I219180,I219211,I335077,I219228,I219254,I219262,I219293,I219324,I219341,I219372,I335095,I219472,I219498,I219506,I219523,I219540,I219566,I219574,I219600,I219608,I219625,I219642,I219659,I219455,I219699,I219707,I219724,I219741,I219758,I219458,I219789,I219806,I219832,I219840,I219440,I219871,I219449,I219902,I219919,I219461,I219950,I219452,I219443,I219446,I219464,I220050,I220076,I220084,I220101,I220118,I220144,I220152,I220178,I220186,I220203,I220220,I220237,I220033,I220277,I220285,I220302,I220319,I220336,I220036,I220367,I220384,I220410,I220418,I220018,I220449,I220027,I220480,I220497,I220039,I220528,I220030,I220021,I220024,I220042,I220628,I220654,I220662,I220679,I220696,I220722,I220730,I220756,I220764,I220781,I220798,I220815,I220855,I220863,I220880,I220897,I220914,I220945,I220962,I220988,I220996,I221027,I221058,I221075,I221106,I221206,I384860,I221232,I221240,I221257,I384845,I384833,I221274,I384848,I221300,I221308,I384851,I221334,I221342,I221359,I221376,I221393,I221189,I384839,I221433,I221441,I221458,I221475,I221492,I221192,I221523,I384836,I384842,I221540,I384857,I221566,I221574,I221174,I221605,I221183,I221636,I221653,I221195,I221684,I384854,I221186,I221177,I221180,I221198,I221784,I221810,I221818,I221835,I221852,I221878,I221886,I221912,I221920,I221937,I221954,I221971,I222011,I222019,I222036,I222053,I222070,I222101,I222118,I222144,I222152,I222183,I222214,I222231,I222262,I222362,I222388,I222396,I222413,I222430,I222456,I222464,I222490,I222498,I222515,I222532,I222549,I222589,I222597,I222614,I222631,I222648,I222679,I222696,I222722,I222730,I222761,I222792,I222809,I222840,I222940,I222966,I222974,I222991,I223008,I223034,I223042,I223068,I223076,I223093,I223110,I223127,I223167,I223175,I223192,I223209,I223226,I223257,I223274,I223300,I223308,I223339,I223370,I223387,I223418,I223518,I223544,I223552,I223569,I223586,I223612,I223620,I223646,I223654,I223671,I223688,I223705,I223501,I223745,I223753,I223770,I223787,I223804,I223504,I223835,I223852,I223878,I223886,I223486,I223917,I223495,I223948,I223965,I223507,I223996,I223498,I223489,I223492,I223510,I224096,I224122,I224130,I224147,I224164,I224190,I224198,I224224,I224232,I224249,I224266,I224283,I224323,I224331,I224348,I224365,I224382,I224413,I224430,I224456,I224464,I224495,I224526,I224543,I224574,I224674,I352414,I224700,I224708,I224725,I352417,I352426,I224742,I352429,I224768,I224776,I352438,I352420,I224802,I224810,I224827,I224844,I224861,I224657,I224901,I224909,I224926,I224943,I224960,I224660,I224991,I352435,I225008,I352432,I225034,I225042,I224642,I225073,I224651,I225104,I225121,I224663,I225152,I352423,I224654,I224645,I224648,I224666,I225252,I371770,I225278,I225286,I225303,I371755,I371743,I225320,I371758,I225346,I225354,I371761,I225380,I225388,I225405,I225422,I225439,I371749,I225479,I225487,I225504,I225521,I225538,I225569,I371746,I371752,I225586,I371767,I225612,I225620,I225651,I225682,I225699,I225730,I371764,I225830,I225856,I225864,I225881,I225898,I225924,I225932,I225958,I225966,I225983,I226000,I226017,I226057,I226065,I226082,I226099,I226116,I226147,I226164,I226190,I226198,I226229,I226260,I226277,I226308,I226408,I226434,I226442,I226459,I226476,I226502,I226510,I226536,I226544,I226561,I226578,I226595,I226635,I226643,I226660,I226677,I226694,I226725,I226742,I226768,I226776,I226807,I226838,I226855,I226886,I226986,I284183,I227012,I227020,I227037,I284159,I284174,I227054,I284186,I227080,I227088,I284171,I284162,I227114,I227122,I227139,I227156,I227173,I226969,I227213,I227221,I227238,I227255,I227272,I226972,I227303,I284177,I284168,I227320,I284180,I227346,I227354,I226954,I227385,I226963,I227416,I227433,I226975,I227464,I284165,I226966,I226957,I226960,I226978,I227564,I340294,I227590,I227598,I227615,I340276,I340288,I227632,I340291,I227658,I227666,I340285,I340282,I227692,I227700,I227717,I227734,I227751,I227547,I340300,I227791,I227799,I227816,I227833,I227850,I227550,I227881,I340279,I227898,I227924,I227932,I227532,I227963,I227541,I227994,I228011,I227553,I228042,I340297,I227544,I227535,I227538,I227556,I228142,I279015,I228168,I228176,I228193,I278991,I279006,I228210,I279018,I228236,I228244,I279003,I278994,I228270,I228278,I228295,I228312,I228329,I228125,I228369,I228377,I228394,I228411,I228428,I228128,I228459,I279009,I279000,I228476,I279012,I228502,I228510,I228110,I228541,I228119,I228572,I228589,I228131,I228620,I278997,I228122,I228113,I228116,I228134,I228720,I228746,I228754,I228771,I228788,I228814,I228822,I228848,I228856,I228873,I228890,I228907,I228703,I228947,I228955,I228972,I228989,I229006,I228706,I229037,I229054,I229080,I229088,I228688,I229119,I228697,I229150,I229167,I228709,I229198,I228700,I228691,I228694,I228712,I229298,I317752,I229324,I229332,I229349,I317734,I317746,I229366,I317749,I229392,I229400,I317743,I317740,I229426,I229434,I229451,I229468,I229485,I229281,I317758,I229525,I229533,I229550,I229567,I229584,I229284,I229615,I317737,I229632,I229658,I229666,I229266,I229697,I229275,I229728,I229745,I229287,I229776,I317755,I229278,I229269,I229272,I229290,I229873,I257030,I229899,I229907,I229924,I257045,I257027,I229941,I229967,I229862,I257036,I229998,I230006,I257054,I230023,I230049,I230057,I229865,I257051,I230097,I229856,I229847,I230133,I257048,I257039,I230150,I257033,I230176,I230184,I230201,I229850,I230232,I257042,I230249,I230266,I229859,I230297,I229844,I230328,I230345,I229853,I230400,I230426,I230434,I230451,I230468,I230494,I230389,I230525,I230533,I230550,I230576,I230584,I230392,I230624,I230383,I230374,I230660,I230677,I230703,I230711,I230728,I230377,I230759,I230776,I230793,I230386,I230824,I230371,I230855,I230872,I230380,I230927,I230953,I230961,I230978,I230995,I231021,I231052,I231060,I231077,I231103,I231111,I231151,I231187,I231204,I231230,I231238,I231255,I231286,I231303,I231320,I231351,I231382,I231399,I231454,I302239,I231480,I231488,I231505,I302248,I302236,I231522,I302233,I231548,I231443,I231579,I231587,I302230,I231604,I231630,I231638,I231446,I231678,I231437,I231428,I231714,I302251,I302242,I231731,I302245,I231757,I231765,I231782,I231431,I231813,I231830,I231847,I231440,I231878,I231425,I231909,I231926,I231434,I231981,I232007,I232015,I232032,I232049,I232075,I232106,I232114,I232131,I232157,I232165,I232205,I232241,I232258,I232284,I232292,I232309,I232340,I232357,I232374,I232405,I232436,I232453,I232508,I232534,I232542,I232559,I232576,I232602,I232497,I232633,I232641,I232658,I232684,I232692,I232500,I232732,I232491,I232482,I232768,I232785,I232811,I232819,I232836,I232485,I232867,I232884,I232901,I232494,I232932,I232479,I232963,I232980,I232488,I233035,I338560,I233061,I233069,I233086,I338542,I233103,I338548,I233129,I338545,I233160,I233168,I338554,I233185,I233211,I233219,I338566,I233259,I233295,I338557,I338551,I233312,I233338,I233346,I233363,I233394,I338563,I233411,I233428,I233459,I233490,I233507,I233562,I260906,I233588,I233596,I233613,I260921,I260903,I233630,I233656,I260912,I233687,I233695,I260930,I233712,I233738,I233746,I260927,I233786,I233822,I260924,I260915,I233839,I260909,I233865,I233873,I233890,I233921,I260918,I233938,I233955,I233986,I234017,I234034,I234089,I234115,I234123,I234140,I234157,I234183,I234078,I234214,I234222,I234239,I234265,I234273,I234081,I234313,I234072,I234063,I234349,I234366,I234392,I234400,I234417,I234066,I234448,I234465,I234482,I234075,I234513,I234060,I234544,I234561,I234069,I234616,I391393,I234642,I234650,I234667,I391390,I391399,I234684,I391378,I234710,I391381,I234741,I234749,I391396,I234766,I234792,I234800,I391402,I234840,I234876,I391384,I391405,I234893,I391387,I234919,I234927,I234944,I234975,I234992,I235009,I235040,I235071,I235088,I235143,I235169,I235177,I235194,I235211,I235237,I235268,I235276,I235293,I235319,I235327,I235367,I235403,I235420,I235446,I235454,I235471,I235502,I235519,I235536,I235567,I235598,I235615,I235670,I235696,I235704,I235721,I235738,I235764,I235659,I235795,I235803,I235820,I235846,I235854,I235662,I235894,I235653,I235644,I235930,I235947,I235973,I235981,I235998,I235647,I236029,I236046,I236063,I235656,I236094,I235641,I236125,I236142,I235650,I236197,I236223,I236231,I236248,I236265,I236291,I236322,I236330,I236347,I236373,I236381,I236421,I236457,I236474,I236500,I236508,I236525,I236556,I236573,I236590,I236621,I236652,I236669,I236724,I236750,I236758,I236775,I236792,I236818,I236849,I236857,I236874,I236900,I236908,I236948,I236984,I237001,I237027,I237035,I237052,I237083,I237100,I237117,I237148,I237179,I237196,I237251,I237277,I237285,I237302,I237319,I237345,I237376,I237384,I237401,I237427,I237435,I237475,I237511,I237528,I237554,I237562,I237579,I237610,I237627,I237644,I237675,I237706,I237723,I237778,I261552,I237804,I237812,I237829,I261567,I261549,I237846,I237872,I261558,I237903,I237911,I261576,I237928,I237954,I237962,I261573,I238002,I238038,I261570,I261561,I238055,I261555,I238081,I238089,I238106,I238137,I261564,I238154,I238171,I238202,I238233,I238250,I238305,I238331,I238339,I238356,I238373,I238399,I238294,I238430,I238438,I238455,I238481,I238489,I238297,I238529,I238288,I238279,I238565,I238582,I238608,I238616,I238633,I238282,I238664,I238681,I238698,I238291,I238729,I238276,I238760,I238777,I238285,I238832,I296629,I238858,I238866,I238883,I296638,I296626,I238900,I296623,I238926,I238821,I238957,I238965,I296620,I238982,I239008,I239016,I238824,I239056,I238815,I238806,I239092,I296641,I296632,I239109,I296635,I239135,I239143,I239160,I238809,I239191,I239208,I239225,I238818,I239256,I238803,I239287,I239304,I238812,I239359,I239385,I239393,I239410,I239427,I239453,I239484,I239492,I239509,I239535,I239543,I239583,I239619,I239636,I239662,I239670,I239687,I239718,I239735,I239752,I239783,I239814,I239831,I239886,I239912,I239920,I239937,I239954,I239980,I240011,I240019,I240036,I240062,I240070,I240110,I240146,I240163,I240189,I240197,I240214,I240245,I240262,I240279,I240310,I240341,I240358,I240413,I322376,I240439,I240447,I240464,I322358,I240481,I322364,I240507,I322361,I240538,I240546,I322370,I240563,I240589,I240597,I322382,I240637,I240673,I322373,I322367,I240690,I240716,I240724,I240741,I240772,I322379,I240789,I240806,I240837,I240868,I240885,I240940,I240966,I240974,I240991,I241008,I241034,I241065,I241073,I241090,I241116,I241124,I241164,I241200,I241217,I241243,I241251,I241268,I241299,I241316,I241333,I241364,I241395,I241412,I241467,I313128,I241493,I241501,I241518,I313110,I241535,I313116,I241561,I313113,I241592,I241600,I313122,I241617,I241643,I241651,I313134,I241691,I241727,I313125,I313119,I241744,I241770,I241778,I241795,I241826,I313131,I241843,I241860,I241891,I241922,I241939,I241994,I374733,I242020,I242028,I242045,I374730,I374739,I242062,I374718,I242088,I374721,I242119,I242127,I374736,I242144,I242170,I242178,I374742,I242218,I242254,I374724,I374745,I242271,I374727,I242297,I242305,I242322,I242353,I242370,I242387,I242418,I242449,I242466,I242521,I242547,I242555,I242572,I242589,I242615,I242646,I242654,I242671,I242697,I242705,I242745,I242781,I242798,I242824,I242832,I242849,I242880,I242897,I242914,I242945,I242976,I242993,I243048,I376518,I243074,I243082,I243099,I376515,I376524,I243116,I376503,I243142,I243037,I376506,I243173,I243181,I376521,I243198,I243224,I243232,I243040,I376527,I243272,I243031,I243022,I243308,I376509,I376530,I243325,I376512,I243351,I243359,I243376,I243025,I243407,I243424,I243441,I243034,I243472,I243019,I243503,I243520,I243028,I243575,I243601,I243609,I243626,I243643,I243669,I243564,I243700,I243708,I243725,I243751,I243759,I243567,I243799,I243558,I243549,I243835,I243852,I243878,I243886,I243903,I243552,I243934,I243951,I243968,I243561,I243999,I243546,I244030,I244047,I243555,I244102,I301117,I244128,I244136,I244153,I301126,I301114,I244170,I301111,I244196,I244091,I244227,I244235,I301108,I244252,I244278,I244286,I244094,I244326,I244085,I244076,I244362,I301129,I301120,I244379,I301123,I244405,I244413,I244430,I244079,I244461,I244478,I244495,I244088,I244526,I244073,I244557,I244574,I244082,I244629,I244655,I244663,I244680,I244697,I244723,I244754,I244762,I244779,I244805,I244813,I244853,I244889,I244906,I244932,I244940,I244957,I244988,I245005,I245022,I245053,I245084,I245101,I245156,I245182,I245190,I245207,I245224,I245250,I245281,I245289,I245306,I245332,I245340,I245380,I245416,I245433,I245459,I245467,I245484,I245515,I245532,I245549,I245580,I245611,I245628,I245683,I314284,I245709,I245717,I245734,I314266,I245751,I314272,I245777,I314269,I245808,I245816,I314278,I245833,I245859,I245867,I314290,I245907,I245943,I314281,I314275,I245960,I245986,I245994,I246011,I246042,I314287,I246059,I246076,I246107,I246138,I246155,I246210,I330468,I246236,I246244,I246261,I330450,I246278,I330456,I246304,I246199,I330453,I246335,I246343,I330462,I246360,I246386,I246394,I246202,I330474,I246434,I246193,I246184,I246470,I330465,I330459,I246487,I246513,I246521,I246538,I246187,I246569,I330471,I246586,I246603,I246196,I246634,I246181,I246665,I246682,I246190,I246737,I264136,I246763,I246771,I246788,I264151,I264133,I246805,I246831,I264142,I246862,I246870,I264160,I246887,I246913,I246921,I264157,I246961,I246997,I264154,I264145,I247014,I264139,I247040,I247048,I247065,I247096,I264148,I247113,I247130,I247161,I247192,I247209,I247264,I247290,I247298,I247315,I247332,I247358,I247389,I247397,I247414,I247440,I247448,I247488,I247524,I247541,I247567,I247575,I247592,I247623,I247640,I247657,I247688,I247719,I247736,I247791,I375923,I247817,I247825,I247842,I375920,I375929,I247859,I375908,I247885,I375911,I247916,I247924,I375926,I247941,I247967,I247975,I375932,I248015,I248051,I375914,I375935,I248068,I375917,I248094,I248102,I248119,I248150,I248167,I248184,I248215,I248246,I248263,I248318,I348074,I248344,I248352,I248369,I348080,I348062,I248386,I348071,I248412,I348077,I248443,I248451,I348065,I248468,I248494,I248502,I348083,I248542,I248578,I348068,I248595,I348086,I248621,I248629,I248646,I248677,I248694,I248711,I248742,I248773,I248790,I248845,I300556,I248871,I248879,I248896,I300565,I300553,I248913,I300550,I248939,I248970,I248978,I300547,I248995,I249021,I249029,I249069,I249105,I300568,I300559,I249122,I300562,I249148,I249156,I249173,I249204,I249221,I249238,I249269,I249300,I249317,I249372,I249398,I249406,I249423,I249440,I249466,I249497,I249505,I249522,I249548,I249556,I249596,I249632,I249649,I249675,I249683,I249700,I249731,I249748,I249765,I249796,I249827,I249844,I249899,I249925,I249933,I249950,I249967,I249993,I250024,I250032,I250049,I250075,I250083,I250123,I250159,I250176,I250202,I250210,I250227,I250258,I250275,I250292,I250323,I250354,I250371,I250426,I352970,I250452,I250460,I250477,I352976,I352958,I250494,I352967,I250520,I352973,I250551,I250559,I352961,I250576,I250602,I250610,I352979,I250650,I250686,I352964,I250703,I352982,I250729,I250737,I250754,I250785,I250802,I250819,I250850,I250881,I250898,I250953,I250979,I250987,I251004,I251021,I251047,I251078,I251086,I251103,I251129,I251137,I251177,I251213,I251230,I251256,I251264,I251281,I251312,I251329,I251346,I251377,I251408,I251425,I251480,I269304,I251506,I251514,I251531,I269319,I269301,I251548,I251574,I251469,I269310,I251605,I251613,I269328,I251630,I251656,I251664,I251472,I269325,I251704,I251463,I251454,I251740,I269322,I269313,I251757,I269307,I251783,I251791,I251808,I251457,I251839,I269316,I251856,I251873,I251466,I251904,I251451,I251935,I251952,I251460,I252007,I252033,I252041,I252058,I252075,I252101,I252132,I252140,I252157,I252183,I252191,I252231,I252267,I252284,I252310,I252318,I252335,I252366,I252383,I252400,I252431,I252462,I252479,I252540,I252566,I252583,I252591,I252608,I252625,I252642,I252659,I252676,I252526,I252707,I252724,I252529,I252755,I252772,I252789,I252505,I252820,I252517,I252860,I252868,I252885,I252902,I252919,I252532,I252950,I252967,I252984,I253010,I252520,I253032,I253049,I252514,I253080,I252508,I252511,I253125,I252523,I253186,I253212,I253229,I253237,I253254,I253271,I253288,I253305,I253322,I253353,I253370,I253401,I253418,I253435,I253466,I253506,I253514,I253531,I253548,I253565,I253596,I253613,I253630,I253656,I253678,I253695,I253726,I253771,I253832,I303352,I253858,I303355,I253875,I253883,I253900,I253917,I303364,I253934,I303373,I253951,I303361,I253968,I253818,I253999,I254016,I253821,I254047,I254064,I303367,I254081,I253797,I254112,I253809,I254152,I254160,I254177,I254194,I303358,I254211,I253824,I254242,I303370,I254259,I254276,I254302,I253812,I254324,I254341,I253806,I254372,I253800,I253803,I254417,I253815,I254478,I254504,I254521,I254529,I254546,I254563,I254580,I254597,I254614,I254464,I254645,I254662,I254467,I254693,I254710,I254727,I254443,I254758,I254455,I254798,I254806,I254823,I254840,I254857,I254470,I254888,I254905,I254922,I254948,I254458,I254970,I254987,I254452,I255018,I254446,I254449,I255063,I254461,I255124,I255150,I255167,I255175,I255192,I255209,I255226,I255243,I255260,I255291,I255308,I255339,I255356,I255373,I255404,I255444,I255452,I255469,I255486,I255503,I255534,I255551,I255568,I255594,I255616,I255633,I255664,I255709,I255770,I255796,I255813,I255821,I255838,I255855,I255872,I255889,I255906,I255937,I255954,I255985,I256002,I256019,I256050,I256090,I256098,I256115,I256132,I256149,I256180,I256197,I256214,I256240,I256262,I256279,I256310,I256355,I256416,I256442,I256459,I256467,I256484,I256501,I256518,I256535,I256552,I256402,I256583,I256600,I256405,I256631,I256648,I256665,I256381,I256696,I256393,I256736,I256744,I256761,I256778,I256795,I256408,I256826,I256843,I256860,I256886,I256396,I256908,I256925,I256390,I256956,I256384,I256387,I257001,I256399,I257062,I257088,I257105,I257113,I257130,I257147,I257164,I257181,I257198,I257229,I257246,I257277,I257294,I257311,I257342,I257382,I257390,I257407,I257424,I257441,I257472,I257489,I257506,I257532,I257554,I257571,I257602,I257647,I257708,I257734,I257751,I257759,I257776,I257793,I257810,I257827,I257844,I257875,I257892,I257923,I257940,I257957,I257988,I258028,I258036,I258053,I258070,I258087,I258118,I258135,I258152,I258178,I258200,I258217,I258248,I258293,I258354,I258380,I258397,I258405,I258422,I258439,I258456,I258473,I258490,I258340,I258521,I258538,I258343,I258569,I258586,I258603,I258319,I258634,I258331,I258674,I258682,I258699,I258716,I258733,I258346,I258764,I258781,I258798,I258824,I258334,I258846,I258863,I258328,I258894,I258322,I258325,I258939,I258337,I259000,I259026,I259043,I259051,I259068,I259085,I259102,I259119,I259136,I259167,I259184,I259215,I259232,I259249,I259280,I259320,I259328,I259345,I259362,I259379,I259410,I259427,I259444,I259470,I259492,I259509,I259540,I259585,I259646,I390188,I259672,I390212,I259689,I259697,I259714,I390194,I259731,I390203,I259748,I259765,I390209,I259782,I259813,I259830,I259861,I259878,I390206,I259895,I259926,I259966,I259974,I259991,I260008,I390200,I260025,I260056,I390191,I260073,I390215,I260090,I390197,I260116,I260138,I260155,I260186,I260231,I260292,I260318,I260335,I260343,I260360,I260377,I260394,I260411,I260428,I260459,I260476,I260507,I260524,I260541,I260572,I260612,I260620,I260637,I260654,I260671,I260702,I260719,I260736,I260762,I260784,I260801,I260832,I260877,I260938,I260964,I260981,I260989,I261006,I261023,I261040,I261057,I261074,I261105,I261122,I261153,I261170,I261187,I261218,I261258,I261266,I261283,I261300,I261317,I261348,I261365,I261382,I261408,I261430,I261447,I261478,I261523,I261584,I261610,I261627,I261635,I261652,I261669,I261686,I261703,I261720,I261751,I261768,I261799,I261816,I261833,I261864,I261904,I261912,I261929,I261946,I261963,I261994,I262011,I262028,I262054,I262076,I262093,I262124,I262169,I262230,I294376,I262256,I294379,I262273,I262281,I262298,I262315,I294388,I262332,I294397,I262349,I294385,I262366,I262216,I262397,I262414,I262219,I262445,I262462,I294391,I262479,I262195,I262510,I262207,I262550,I262558,I262575,I262592,I294382,I262609,I262222,I262640,I294394,I262657,I262674,I262700,I262210,I262722,I262739,I262204,I262770,I262198,I262201,I262815,I262213,I262876,I332780,I262902,I332762,I262919,I262927,I262944,I332771,I262961,I332783,I262978,I332765,I262995,I332774,I263012,I263043,I263060,I263091,I263108,I332786,I263125,I263156,I263196,I263204,I263221,I263238,I263255,I263286,I332768,I263303,I332777,I263320,I263346,I263368,I263385,I263416,I263461,I263522,I263548,I263565,I263573,I263590,I263607,I263624,I263641,I263658,I263508,I263689,I263706,I263511,I263737,I263754,I263771,I263487,I263802,I263499,I263842,I263850,I263867,I263884,I263901,I263514,I263932,I263949,I263966,I263992,I263502,I264014,I264031,I263496,I264062,I263490,I263493,I264107,I263505,I264168,I264194,I264211,I264219,I264236,I264253,I264270,I264287,I264304,I264335,I264352,I264383,I264400,I264417,I264448,I264488,I264496,I264513,I264530,I264547,I264578,I264595,I264612,I264638,I264660,I264677,I264708,I264753,I264814,I264840,I264857,I264865,I264882,I264899,I264916,I264933,I264950,I264981,I264998,I265029,I265046,I265063,I265094,I265134,I265142,I265159,I265176,I265193,I265224,I265241,I265258,I265284,I265306,I265323,I265354,I265399,I265460,I265486,I265503,I265511,I265528,I265545,I265562,I265579,I265596,I265627,I265644,I265675,I265692,I265709,I265740,I265780,I265788,I265805,I265822,I265839,I265870,I265887,I265904,I265930,I265952,I265969,I266000,I266045,I266106,I266132,I266149,I266157,I266174,I266191,I266208,I266225,I266242,I266092,I266273,I266290,I266095,I266321,I266338,I266355,I266071,I266386,I266083,I266426,I266434,I266451,I266468,I266485,I266098,I266516,I266533,I266550,I266576,I266086,I266598,I266615,I266080,I266646,I266074,I266077,I266691,I266089,I266752,I304474,I266778,I304477,I266795,I266803,I266820,I266837,I304486,I266854,I304495,I266871,I304483,I266888,I266919,I266936,I266967,I266984,I304489,I267001,I267032,I267072,I267080,I267097,I267114,I304480,I267131,I267162,I304492,I267179,I267196,I267222,I267244,I267261,I267292,I267337,I267398,I267424,I267441,I267449,I267466,I267483,I267500,I267517,I267534,I267565,I267582,I267613,I267630,I267647,I267678,I267718,I267726,I267743,I267760,I267777,I267808,I267825,I267842,I267868,I267890,I267907,I267938,I267983,I268044,I268070,I268087,I268095,I268112,I268129,I268146,I268163,I268180,I268211,I268228,I268259,I268276,I268293,I268324,I268364,I268372,I268389,I268406,I268423,I268454,I268471,I268488,I268514,I268536,I268553,I268584,I268629,I268690,I268716,I268733,I268741,I268758,I268775,I268792,I268809,I268826,I268857,I268874,I268905,I268922,I268939,I268970,I269010,I269018,I269035,I269052,I269069,I269100,I269117,I269134,I269160,I269182,I269199,I269230,I269275,I269336,I269362,I269379,I269387,I269404,I269421,I269438,I269455,I269472,I269503,I269520,I269551,I269568,I269585,I269616,I269656,I269664,I269681,I269698,I269715,I269746,I269763,I269780,I269806,I269828,I269845,I269876,I269921,I269982,I270008,I270025,I270033,I270050,I270067,I270084,I270101,I270118,I269968,I270149,I270166,I269971,I270197,I270214,I270231,I269947,I270262,I269959,I270302,I270310,I270327,I270344,I270361,I269974,I270392,I270409,I270426,I270452,I269962,I270474,I270491,I269956,I270522,I269950,I269953,I270567,I269965,I270628,I311972,I270654,I311954,I270671,I270679,I270696,I311963,I270713,I311975,I270730,I311957,I270747,I311966,I270764,I270795,I270812,I270843,I270860,I311978,I270877,I270908,I270948,I270956,I270973,I270990,I271007,I271038,I311960,I271055,I311969,I271072,I271098,I271120,I271137,I271168,I271213,I271274,I392568,I271300,I392592,I271317,I271325,I271342,I392574,I271359,I392583,I271376,I271393,I392589,I271410,I271441,I271458,I271489,I271506,I392586,I271523,I271554,I271594,I271602,I271619,I271636,I392580,I271653,I271684,I392571,I271701,I392595,I271718,I392577,I271744,I271766,I271783,I271814,I271859,I271920,I271946,I271963,I271971,I271988,I272005,I272022,I272039,I272056,I271906,I272087,I272104,I271909,I272135,I272152,I272169,I271885,I272200,I271897,I272240,I272248,I272265,I272282,I272299,I271912,I272330,I272347,I272364,I272390,I271900,I272412,I272429,I271894,I272460,I271888,I271891,I272505,I271903,I272566,I272592,I272609,I272617,I272634,I272651,I272668,I272685,I272702,I272733,I272750,I272781,I272798,I272815,I272846,I272886,I272894,I272911,I272928,I272945,I272976,I272993,I273010,I273036,I273058,I273075,I273106,I273151,I273212,I387808,I273238,I387832,I273255,I273263,I273280,I387814,I273297,I387823,I273314,I273331,I387829,I273348,I273198,I273379,I273396,I273201,I273427,I273444,I387826,I273461,I273177,I273492,I273189,I273532,I273540,I273557,I273574,I387820,I273591,I273204,I273622,I387811,I273639,I387835,I273656,I387817,I273682,I273192,I273704,I273721,I273186,I273752,I273180,I273183,I273797,I273195,I273858,I363711,I273884,I363705,I273901,I273909,I273926,I363714,I273943,I363726,I273960,I363708,I273977,I273994,I274025,I274042,I274073,I274090,I363702,I274107,I274138,I274178,I274186,I274203,I274220,I363723,I274237,I274268,I363717,I274285,I274302,I363720,I274328,I274350,I274367,I274398,I274443,I274504,I274530,I274547,I274555,I274572,I274589,I274606,I274623,I274640,I274490,I274671,I274688,I274493,I274719,I274736,I274753,I274469,I274784,I274481,I274824,I274832,I274849,I274866,I274883,I274496,I274914,I274931,I274948,I274974,I274484,I274996,I275013,I274478,I275044,I274472,I274475,I275089,I274487,I275150,I275176,I275193,I275201,I275218,I275235,I275252,I275269,I275286,I275317,I275334,I275365,I275382,I275399,I275430,I275470,I275478,I275495,I275512,I275529,I275560,I275577,I275594,I275620,I275642,I275659,I275690,I275735,I275796,I336826,I275822,I336808,I275839,I275847,I275864,I336817,I275881,I336829,I275898,I336811,I275915,I336820,I275932,I275963,I275980,I276011,I276028,I336832,I276045,I276076,I276116,I276124,I276141,I276158,I276175,I276206,I336814,I276223,I336823,I276240,I276266,I276288,I276305,I276336,I276381,I276442,I276468,I276485,I276493,I276510,I276527,I276544,I276561,I276578,I276609,I276626,I276657,I276674,I276691,I276722,I276762,I276770,I276787,I276804,I276821,I276852,I276869,I276886,I276912,I276934,I276951,I276982,I277027,I277088,I277114,I277131,I277139,I277156,I277173,I277190,I277207,I277224,I277255,I277272,I277303,I277320,I277337,I277368,I277408,I277416,I277433,I277450,I277467,I277498,I277515,I277532,I277558,I277580,I277597,I277628,I277673,I277734,I277760,I277777,I277785,I277802,I277819,I277836,I277853,I277870,I277901,I277918,I277949,I277966,I277983,I278014,I278054,I278062,I278079,I278096,I278113,I278144,I278161,I278178,I278204,I278226,I278243,I278274,I278319,I278380,I290449,I278406,I290452,I278423,I278431,I278448,I278465,I290461,I278482,I290470,I278499,I290458,I278516,I278366,I278547,I278564,I278369,I278595,I278612,I290464,I278629,I278345,I278660,I278357,I278700,I278708,I278725,I278742,I290455,I278759,I278372,I278790,I290467,I278807,I278824,I278850,I278360,I278872,I278889,I278354,I278920,I278348,I278351,I278965,I278363,I279026,I279052,I279069,I279077,I279094,I279111,I279128,I279145,I279162,I279193,I279210,I279241,I279258,I279275,I279306,I279346,I279354,I279371,I279388,I279405,I279436,I279453,I279470,I279496,I279518,I279535,I279566,I279611,I279672,I345904,I279698,I345910,I279715,I279723,I279740,I345907,I279757,I345886,I279774,I345889,I279791,I345895,I279808,I279839,I279856,I279887,I279904,I279921,I279952,I279992,I280000,I280017,I280034,I345898,I280051,I280082,I280099,I345892,I280116,I345901,I280142,I280164,I280181,I280212,I280257,I280318,I280344,I280361,I280369,I280386,I280403,I280420,I280437,I280454,I280485,I280502,I280533,I280550,I280567,I280598,I280638,I280646,I280663,I280680,I280697,I280728,I280745,I280762,I280788,I280810,I280827,I280858,I280903,I280964,I280990,I281007,I281015,I281032,I281049,I281066,I281083,I281100,I280950,I281131,I281148,I280953,I281179,I281196,I281213,I280929,I281244,I280941,I281284,I281292,I281309,I281326,I281343,I280956,I281374,I281391,I281408,I281434,I280944,I281456,I281473,I280938,I281504,I280932,I280935,I281549,I280947,I281610,I281636,I281653,I281661,I281678,I281695,I281712,I281729,I281746,I281596,I281777,I281794,I281599,I281825,I281842,I281859,I281575,I281890,I281587,I281930,I281938,I281955,I281972,I281989,I281602,I282020,I282037,I282054,I282080,I281590,I282102,I282119,I281584,I282150,I281578,I281581,I282195,I281593,I282256,I349168,I282282,I349174,I282299,I282307,I282324,I349171,I282341,I349150,I282358,I349153,I282375,I349159,I282392,I282423,I282440,I282471,I282488,I282505,I282536,I282576,I282584,I282601,I282618,I349162,I282635,I282666,I282683,I349156,I282700,I349165,I282726,I282748,I282765,I282796,I282841,I282902,I314862,I282928,I314844,I282945,I282953,I282970,I314853,I282987,I314865,I283004,I314847,I283021,I314856,I283038,I283069,I283086,I283117,I283134,I314868,I283151,I283182,I283222,I283230,I283247,I283264,I283281,I283312,I314850,I283329,I314859,I283346,I283372,I283394,I283411,I283442,I283487,I283548,I283574,I283591,I283599,I283616,I283633,I283650,I283667,I283684,I283715,I283732,I283763,I283780,I283797,I283828,I283868,I283876,I283893,I283910,I283927,I283958,I283975,I283992,I284018,I284040,I284057,I284088,I284133,I284194,I284220,I284237,I284245,I284262,I284279,I284296,I284313,I284330,I284361,I284378,I284409,I284426,I284443,I284474,I284514,I284522,I284539,I284556,I284573,I284604,I284621,I284638,I284664,I284686,I284703,I284734,I284779,I284840,I284866,I284883,I284891,I284908,I284925,I284942,I284959,I284976,I284826,I285007,I285024,I284829,I285055,I285072,I285089,I284805,I285120,I284817,I285160,I285168,I285185,I285202,I285219,I284832,I285250,I285267,I285284,I285310,I284820,I285332,I285349,I284814,I285380,I284808,I284811,I285425,I284823,I285486,I285512,I285529,I285537,I285554,I285571,I285588,I285605,I285622,I285653,I285670,I285701,I285718,I285735,I285766,I285806,I285814,I285831,I285848,I285865,I285896,I285913,I285930,I285956,I285978,I285995,I286026,I286071,I286132,I292693,I286158,I292696,I286175,I286183,I286200,I286217,I292705,I286234,I292714,I286251,I292702,I286268,I286118,I286299,I286316,I286121,I286347,I286364,I292708,I286381,I286097,I286412,I286109,I286452,I286460,I286477,I286494,I292699,I286511,I286124,I286542,I292711,I286559,I286576,I286602,I286112,I286624,I286641,I286106,I286672,I286100,I286103,I286717,I286115,I286778,I388403,I286804,I388427,I286821,I286829,I286846,I388409,I286863,I388418,I286880,I286897,I388424,I286914,I286945,I286962,I286993,I287010,I388421,I287027,I287058,I287098,I287106,I287123,I287140,I388415,I287157,I287188,I388406,I287205,I388430,I287222,I388412,I287248,I287270,I287287,I287318,I287363,I287424,I358509,I287450,I358503,I287467,I287475,I287492,I358512,I287509,I358524,I287526,I358506,I287543,I287560,I287591,I287608,I287639,I287656,I358500,I287673,I287704,I287744,I287752,I287769,I287786,I358521,I287803,I287834,I358515,I287851,I287868,I358518,I287894,I287916,I287933,I287964,I288009,I288070,I288096,I288113,I288121,I288138,I288155,I288172,I288189,I288206,I288237,I288254,I288285,I288302,I288319,I288350,I288390,I288398,I288415,I288432,I288449,I288480,I288497,I288514,I288540,I288562,I288579,I288610,I288655,I288716,I288742,I288759,I288767,I288784,I288801,I288818,I288835,I288852,I288702,I288883,I288900,I288705,I288931,I288948,I288965,I288681,I288996,I288693,I289036,I289044,I289061,I289078,I289095,I288708,I289126,I289143,I289160,I289186,I288696,I289208,I289225,I288690,I289256,I288684,I288687,I289301,I288699,I289356,I289382,I289399,I289421,I289447,I289455,I289472,I289489,I289506,I289523,I289540,I289557,I289588,I289619,I289636,I289653,I289670,I289701,I289746,I289763,I289780,I289806,I289814,I289845,I289862,I289917,I289943,I289960,I289982,I290008,I290016,I290033,I290050,I290067,I290084,I290101,I290118,I290149,I290180,I290197,I290214,I290231,I290262,I290307,I290324,I290341,I290367,I290375,I290406,I290423,I290478,I290504,I290521,I290543,I290569,I290577,I290594,I290611,I290628,I290645,I290662,I290679,I290710,I290741,I290758,I290775,I290792,I290823,I290868,I290885,I290902,I290928,I290936,I290967,I290984,I291039,I291065,I291082,I291104,I291130,I291138,I291155,I291172,I291189,I291206,I291223,I291240,I291271,I291302,I291319,I291336,I291353,I291384,I291429,I291446,I291463,I291489,I291497,I291528,I291545,I291600,I351332,I291626,I291643,I291665,I351338,I291691,I291699,I351347,I291716,I291733,I351326,I291750,I351329,I291767,I291784,I351341,I291801,I291832,I291863,I351335,I291880,I291897,I291914,I291945,I291990,I351350,I292007,I292024,I351344,I292050,I292058,I292089,I292106,I292161,I292187,I292204,I292153,I292226,I292252,I292260,I292277,I292294,I292311,I292328,I292345,I292362,I292135,I292393,I292138,I292424,I292441,I292458,I292475,I292147,I292506,I292150,I292144,I292551,I292568,I292585,I292611,I292619,I292132,I292650,I292667,I292141,I292722,I366017,I292748,I292765,I292787,I366014,I292813,I292821,I366020,I292838,I292855,I366029,I292872,I366023,I292889,I292906,I366035,I292923,I292954,I292985,I366032,I293002,I293019,I293036,I293067,I293112,I366026,I293129,I366038,I293146,I293172,I293180,I293211,I293228,I293283,I293309,I293326,I293348,I293374,I293382,I293399,I293416,I293433,I293450,I293467,I293484,I293515,I293546,I293563,I293580,I293597,I293628,I293673,I293690,I293707,I293733,I293741,I293772,I293789,I293844,I293870,I293887,I293909,I293935,I293943,I293960,I293977,I293994,I294011,I294028,I294045,I294076,I294107,I294124,I294141,I294158,I294189,I294234,I294251,I294268,I294294,I294302,I294333,I294350,I294405,I294431,I294448,I294470,I294496,I294504,I294521,I294538,I294555,I294572,I294589,I294606,I294637,I294668,I294685,I294702,I294719,I294750,I294795,I294812,I294829,I294855,I294863,I294894,I294911,I294966,I329309,I294992,I295009,I294958,I295031,I329300,I295057,I295065,I329297,I295082,I295099,I329306,I295116,I329315,I295133,I295150,I329294,I295167,I294940,I295198,I294943,I295229,I329303,I295246,I295263,I295280,I294952,I295311,I294955,I294949,I295356,I329318,I295373,I295390,I329312,I295416,I295424,I294937,I295455,I295472,I294946,I295527,I383063,I295553,I295570,I295592,I383057,I295618,I295626,I383048,I295643,I295660,I383075,I295677,I383060,I383069,I295694,I295711,I383054,I295728,I295759,I295790,I383072,I295807,I295824,I295841,I295872,I295917,I383066,I295934,I295951,I383051,I295977,I295985,I296016,I296033,I296088,I296114,I296131,I296080,I296153,I296179,I296187,I296204,I296221,I296238,I296255,I296272,I296289,I296062,I296320,I296065,I296351,I296368,I296385,I296402,I296074,I296433,I296077,I296071,I296478,I296495,I296512,I296538,I296546,I296059,I296577,I296594,I296068,I296649,I296675,I296692,I296714,I296740,I296748,I296765,I296782,I296799,I296816,I296833,I296850,I296881,I296912,I296929,I296946,I296963,I296994,I297039,I297056,I297073,I297099,I297107,I297138,I297155,I297210,I357925,I297236,I297253,I297202,I297275,I357922,I297301,I297309,I357928,I297326,I297343,I357937,I297360,I357931,I297377,I297394,I357943,I297411,I297184,I297442,I297187,I297473,I357940,I297490,I297507,I297524,I297196,I297555,I297199,I297193,I297600,I357934,I297617,I357946,I297634,I297660,I297668,I297181,I297699,I297716,I297190,I297771,I297797,I297814,I297836,I297862,I297870,I297887,I297904,I297921,I297938,I297955,I297972,I298003,I298034,I298051,I298068,I298085,I298116,I298161,I298178,I298195,I298221,I298229,I298260,I298277,I298332,I298358,I298375,I298397,I298423,I298431,I298448,I298465,I298482,I298499,I298516,I298533,I298564,I298595,I298612,I298629,I298646,I298677,I298722,I298739,I298756,I298782,I298790,I298821,I298838,I298893,I298919,I298936,I298958,I298984,I298992,I299009,I299026,I299043,I299060,I299077,I299094,I299125,I299156,I299173,I299190,I299207,I299238,I299283,I299300,I299317,I299343,I299351,I299382,I299399,I299454,I299480,I299497,I299519,I299545,I299553,I299570,I299587,I299604,I299621,I299638,I299655,I299686,I299717,I299734,I299751,I299768,I299799,I299844,I299861,I299878,I299904,I299912,I299943,I299960,I300015,I300041,I300058,I300080,I300106,I300114,I300131,I300148,I300165,I300182,I300199,I300216,I300247,I300278,I300295,I300312,I300329,I300360,I300405,I300422,I300439,I300465,I300473,I300504,I300521,I300576,I300602,I300619,I300641,I300667,I300675,I300692,I300709,I300726,I300743,I300760,I300777,I300808,I300839,I300856,I300873,I300890,I300921,I300966,I300983,I301000,I301026,I301034,I301065,I301082,I301137,I301163,I301180,I301202,I301228,I301236,I301253,I301270,I301287,I301304,I301321,I301338,I301369,I301400,I301417,I301434,I301451,I301482,I301527,I301544,I301561,I301587,I301595,I301626,I301643,I301698,I301724,I301741,I301690,I301763,I301789,I301797,I301814,I301831,I301848,I301865,I301882,I301899,I301672,I301930,I301675,I301961,I301978,I301995,I302012,I301684,I302043,I301687,I301681,I302088,I302105,I302122,I302148,I302156,I301669,I302187,I302204,I301678,I302259,I302285,I302302,I302324,I302350,I302358,I302375,I302392,I302409,I302426,I302443,I302460,I302491,I302522,I302539,I302556,I302573,I302604,I302649,I302666,I302683,I302709,I302717,I302748,I302765,I302820,I310235,I302846,I302863,I302885,I310226,I302911,I302919,I310223,I302936,I302953,I310232,I302970,I310241,I302987,I303004,I310220,I303021,I303052,I303083,I310229,I303100,I303117,I303134,I303165,I303210,I310244,I303227,I303244,I310238,I303270,I303278,I303309,I303326,I303381,I303407,I303424,I303446,I303472,I303480,I303497,I303514,I303531,I303548,I303565,I303582,I303613,I303644,I303661,I303678,I303695,I303726,I303771,I303788,I303805,I303831,I303839,I303870,I303887,I303942,I386038,I303968,I303985,I304007,I386032,I304033,I304041,I386023,I304058,I304075,I386050,I304092,I386035,I386044,I304109,I304126,I386029,I304143,I304174,I304205,I386047,I304222,I304239,I304256,I304287,I304332,I386041,I304349,I304366,I386026,I304392,I304400,I304431,I304448,I304503,I389013,I304529,I304546,I304568,I389007,I304594,I304602,I388998,I304619,I304636,I389025,I304653,I389010,I389019,I304670,I304687,I389004,I304704,I304735,I304766,I389022,I304783,I304800,I304817,I304848,I304893,I389016,I304910,I304927,I389001,I304953,I304961,I304992,I305009,I305064,I305090,I305107,I305056,I305129,I305155,I305163,I305180,I305197,I305214,I305231,I305248,I305265,I305038,I305296,I305041,I305327,I305344,I305361,I305378,I305050,I305409,I305053,I305047,I305454,I305471,I305488,I305514,I305522,I305035,I305553,I305570,I305044,I305628,I305654,I305662,I305702,I305710,I305727,I305744,I305784,I305806,I305823,I305849,I305857,I305874,I305891,I305908,I305925,I305970,I306001,I306018,I306044,I306052,I306083,I306100,I306117,I306134,I306206,I306232,I306240,I306280,I306288,I306305,I306322,I306362,I306384,I306401,I306427,I306435,I306452,I306469,I306486,I306503,I306548,I306579,I306596,I306622,I306630,I306661,I306678,I306695,I306712,I306784,I306810,I306818,I306858,I306866,I306883,I306900,I306940,I306962,I306979,I307005,I307013,I307030,I307047,I307064,I307081,I307126,I307157,I307174,I307200,I307208,I307239,I307256,I307273,I307290,I307362,I307388,I307396,I307436,I307444,I307461,I307478,I307518,I307540,I307557,I307583,I307591,I307608,I307625,I307642,I307659,I307704,I307735,I307752,I307778,I307786,I307817,I307834,I307851,I307868,I307940,I307966,I307974,I308014,I308022,I308039,I308056,I308096,I308118,I308135,I308161,I308169,I308186,I308203,I308220,I308237,I308282,I308313,I308330,I308356,I308364,I308395,I308412,I308429,I308446,I308518,I380695,I308544,I308552,I380677,I380668,I308592,I308600,I380683,I308617,I380671,I308634,I308674,I308696,I380680,I308713,I308739,I308747,I308764,I380689,I308781,I308798,I308815,I308860,I380692,I308891,I308908,I380686,I380674,I308934,I308942,I308973,I308990,I309007,I309024,I309096,I309122,I309130,I309170,I309178,I309195,I309212,I309252,I309274,I309291,I309317,I309325,I309342,I309359,I309376,I309393,I309438,I309469,I309486,I309512,I309520,I309551,I309568,I309585,I309602,I309674,I309700,I309708,I309748,I309756,I309773,I309790,I309830,I309852,I309869,I309895,I309903,I309920,I309937,I309954,I309971,I310016,I310047,I310064,I310090,I310098,I310129,I310146,I310163,I310180,I310252,I310278,I310286,I310326,I310334,I310351,I310368,I310408,I310430,I310447,I310473,I310481,I310498,I310515,I310532,I310549,I310594,I310625,I310642,I310668,I310676,I310707,I310724,I310741,I310758,I310830,I310856,I310864,I310813,I310904,I310912,I310929,I310946,I310801,I310986,I310822,I311008,I311025,I311051,I311059,I311076,I311093,I311110,I311127,I310798,I310819,I311172,I310810,I311203,I311220,I311246,I311254,I310816,I311285,I311302,I311319,I311336,I310807,I310804,I311408,I311434,I311442,I311391,I311482,I311490,I311507,I311524,I311379,I311564,I311400,I311586,I311603,I311629,I311637,I311654,I311671,I311688,I311705,I311376,I311397,I311750,I311388,I311781,I311798,I311824,I311832,I311394,I311863,I311880,I311897,I311914,I311385,I311382,I311986,I312012,I312020,I312060,I312068,I312085,I312102,I312142,I312164,I312181,I312207,I312215,I312232,I312249,I312266,I312283,I312328,I312359,I312376,I312402,I312410,I312441,I312458,I312475,I312492,I312564,I312590,I312598,I312638,I312646,I312663,I312680,I312720,I312742,I312759,I312785,I312793,I312810,I312827,I312844,I312861,I312906,I312937,I312954,I312980,I312988,I313019,I313036,I313053,I313070,I313142,I313168,I313176,I313216,I313224,I313241,I313258,I313298,I313320,I313337,I313363,I313371,I313388,I313405,I313422,I313439,I313484,I313515,I313532,I313558,I313566,I313597,I313614,I313631,I313648,I313720,I313746,I313754,I313794,I313802,I313819,I313836,I313876,I313898,I313915,I313941,I313949,I313966,I313983,I314000,I314017,I314062,I314093,I314110,I314136,I314144,I314175,I314192,I314209,I314226,I314298,I314324,I314332,I314372,I314380,I314397,I314414,I314454,I314476,I314493,I314519,I314527,I314544,I314561,I314578,I314595,I314640,I314671,I314688,I314714,I314722,I314753,I314770,I314787,I314804,I314876,I314902,I314910,I314950,I314958,I314975,I314992,I315032,I315054,I315071,I315097,I315105,I315122,I315139,I315156,I315173,I315218,I315249,I315266,I315292,I315300,I315331,I315348,I315365,I315382,I315454,I315480,I315488,I315528,I315536,I315553,I315570,I315610,I315632,I315649,I315675,I315683,I315700,I315717,I315734,I315751,I315796,I315827,I315844,I315870,I315878,I315909,I315926,I315943,I315960,I316032,I316058,I316066,I316015,I316106,I316114,I316131,I316148,I316003,I316188,I316024,I316210,I316227,I316253,I316261,I316278,I316295,I316312,I316329,I316000,I316021,I316374,I316012,I316405,I316422,I316448,I316456,I316018,I316487,I316504,I316521,I316538,I316009,I316006,I316610,I375340,I316636,I316644,I375322,I375313,I316684,I316692,I375328,I316709,I375316,I316726,I316766,I316788,I375325,I316805,I316831,I316839,I316856,I375334,I316873,I316890,I316907,I316952,I375337,I316983,I317000,I375331,I375319,I317026,I317034,I317065,I317082,I317099,I317116,I317188,I317214,I317222,I317262,I317270,I317287,I317304,I317344,I317366,I317383,I317409,I317417,I317434,I317451,I317468,I317485,I317530,I317561,I317578,I317604,I317612,I317643,I317660,I317677,I317694,I317766,I317792,I317800,I317840,I317848,I317865,I317882,I317922,I317944,I317961,I317987,I317995,I318012,I318029,I318046,I318063,I318108,I318139,I318156,I318182,I318190,I318221,I318238,I318255,I318272,I318344,I318370,I318378,I318418,I318426,I318443,I318460,I318500,I318522,I318539,I318565,I318573,I318590,I318607,I318624,I318641,I318686,I318717,I318734,I318760,I318768,I318799,I318816,I318833,I318850,I318922,I318948,I318956,I318996,I319004,I319021,I319038,I319078,I319100,I319117,I319143,I319151,I319168,I319185,I319202,I319219,I319264,I319295,I319312,I319338,I319346,I319377,I319394,I319411,I319428,I319500,I319526,I319534,I319574,I319582,I319599,I319616,I319656,I319678,I319695,I319721,I319729,I319746,I319763,I319780,I319797,I319842,I319873,I319890,I319916,I319924,I319955,I319972,I319989,I320006,I320078,I320104,I320112,I320152,I320160,I320177,I320194,I320234,I320256,I320273,I320299,I320307,I320324,I320341,I320358,I320375,I320420,I320451,I320468,I320494,I320502,I320533,I320550,I320567,I320584,I320656,I320682,I320690,I320730,I320738,I320755,I320772,I320812,I320834,I320851,I320877,I320885,I320902,I320919,I320936,I320953,I320998,I321029,I321046,I321072,I321080,I321111,I321128,I321145,I321162,I321234,I321260,I321268,I321308,I321316,I321333,I321350,I321390,I321412,I321429,I321455,I321463,I321480,I321497,I321514,I321531,I321576,I321607,I321624,I321650,I321658,I321689,I321706,I321723,I321740,I321812,I321838,I321846,I321886,I321894,I321911,I321928,I321968,I321990,I322007,I322033,I322041,I322058,I322075,I322092,I322109,I322154,I322185,I322202,I322228,I322236,I322267,I322284,I322301,I322318,I322390,I322416,I322424,I322464,I322472,I322489,I322506,I322546,I322568,I322585,I322611,I322619,I322636,I322653,I322670,I322687,I322732,I322763,I322780,I322806,I322814,I322845,I322862,I322879,I322896,I322968,I322994,I323002,I323042,I323050,I323067,I323084,I323124,I323146,I323163,I323189,I323197,I323214,I323231,I323248,I323265,I323310,I323341,I323358,I323384,I323392,I323423,I323440,I323457,I323474,I323546,I323572,I323580,I323620,I323628,I323645,I323662,I323702,I323724,I323741,I323767,I323775,I323792,I323809,I323826,I323843,I323888,I323919,I323936,I323962,I323970,I324001,I324018,I324035,I324052,I324124,I324150,I324158,I324107,I324198,I324206,I324223,I324240,I324095,I324280,I324116,I324302,I324319,I324345,I324353,I324370,I324387,I324404,I324421,I324092,I324113,I324466,I324104,I324497,I324514,I324540,I324548,I324110,I324579,I324596,I324613,I324630,I324101,I324098,I324702,I324728,I324736,I324776,I324784,I324801,I324818,I324858,I324880,I324897,I324923,I324931,I324948,I324965,I324982,I324999,I325044,I325075,I325092,I325118,I325126,I325157,I325174,I325191,I325208,I325280,I325306,I325314,I325354,I325362,I325379,I325396,I325436,I325458,I325475,I325501,I325509,I325526,I325543,I325560,I325577,I325622,I325653,I325670,I325696,I325704,I325735,I325752,I325769,I325786,I325858,I325884,I325892,I325932,I325940,I325957,I325974,I326014,I326036,I326053,I326079,I326087,I326104,I326121,I326138,I326155,I326200,I326231,I326248,I326274,I326282,I326313,I326330,I326347,I326364,I326436,I359102,I326462,I326470,I359084,I359093,I326510,I326518,I359078,I326535,I359090,I326552,I326592,I326614,I359081,I326631,I326657,I326665,I326682,I326699,I326716,I326733,I326778,I359099,I326809,I326826,I359087,I359096,I326852,I326860,I326891,I326908,I326925,I326942,I327014,I327040,I327048,I327088,I327096,I327113,I327130,I327170,I327192,I327209,I327235,I327243,I327260,I327277,I327294,I327311,I327356,I327387,I327404,I327430,I327438,I327469,I327486,I327503,I327520,I327592,I327618,I327626,I327575,I327666,I327674,I327691,I327708,I327563,I327748,I327584,I327770,I327787,I327813,I327821,I327838,I327855,I327872,I327889,I327560,I327581,I327934,I327572,I327965,I327982,I328008,I328016,I327578,I328047,I328064,I328081,I328098,I327569,I327566,I328170,I328196,I328204,I328244,I328252,I328269,I328286,I328326,I328348,I328365,I328391,I328399,I328416,I328433,I328450,I328467,I328512,I328543,I328560,I328586,I328594,I328625,I328642,I328659,I328676,I328748,I328774,I328782,I328822,I328830,I328847,I328864,I328904,I328926,I328943,I328969,I328977,I328994,I329011,I329028,I329045,I329090,I329121,I329138,I329164,I329172,I329203,I329220,I329237,I329254,I329326,I329352,I329360,I329400,I329408,I329425,I329442,I329482,I329504,I329521,I329547,I329555,I329572,I329589,I329606,I329623,I329668,I329699,I329716,I329742,I329750,I329781,I329798,I329815,I329832,I329904,I329930,I329938,I329978,I329986,I330003,I330020,I330060,I330082,I330099,I330125,I330133,I330150,I330167,I330184,I330201,I330246,I330277,I330294,I330320,I330328,I330359,I330376,I330393,I330410,I330482,I371175,I330508,I330516,I371157,I371148,I330556,I330564,I371163,I330581,I371151,I330598,I330638,I330660,I371160,I330677,I330703,I330711,I330728,I371169,I330745,I330762,I330779,I330824,I371172,I330855,I330872,I371166,I371154,I330898,I330906,I330937,I330954,I330971,I330988,I331060,I331086,I331094,I331134,I331142,I331159,I331176,I331216,I331238,I331255,I331281,I331289,I331306,I331323,I331340,I331357,I331402,I331433,I331450,I331476,I331484,I331515,I331532,I331549,I331566,I331638,I331664,I331672,I331712,I331720,I331737,I331754,I331794,I331816,I331833,I331859,I331867,I331884,I331901,I331918,I331935,I331980,I332011,I332028,I332054,I332062,I332093,I332110,I332127,I332144,I332216,I332242,I332250,I332199,I332290,I332298,I332315,I332332,I332187,I332372,I332208,I332394,I332411,I332437,I332445,I332462,I332479,I332496,I332513,I332184,I332205,I332558,I332196,I332589,I332606,I332632,I332640,I332202,I332671,I332688,I332705,I332722,I332193,I332190,I332794,I332820,I332828,I332868,I332876,I332893,I332910,I332950,I332972,I332989,I333015,I333023,I333040,I333057,I333074,I333091,I333136,I333167,I333184,I333210,I333218,I333249,I333266,I333283,I333300,I333372,I333398,I333406,I333446,I333454,I333471,I333488,I333528,I333550,I333567,I333593,I333601,I333618,I333635,I333652,I333669,I333714,I333745,I333762,I333788,I333796,I333827,I333844,I333861,I333878,I333950,I333976,I333984,I334024,I334032,I334049,I334066,I334106,I334128,I334145,I334171,I334179,I334196,I334213,I334230,I334247,I334292,I334323,I334340,I334366,I334374,I334405,I334422,I334439,I334456,I334528,I334554,I334562,I334511,I334602,I334610,I334627,I334644,I334499,I334684,I334520,I334706,I334723,I334749,I334757,I334774,I334791,I334808,I334825,I334496,I334517,I334870,I334508,I334901,I334918,I334944,I334952,I334514,I334983,I335000,I335017,I335034,I334505,I334502,I335106,I335132,I335140,I335180,I335188,I335205,I335222,I335262,I335284,I335301,I335327,I335335,I335352,I335369,I335386,I335403,I335448,I335479,I335496,I335522,I335530,I335561,I335578,I335595,I335612,I335684,I335710,I335718,I335758,I335766,I335783,I335800,I335840,I335862,I335879,I335905,I335913,I335930,I335947,I335964,I335981,I336026,I336057,I336074,I336100,I336108,I336139,I336156,I336173,I336190,I336262,I336288,I336296,I336336,I336344,I336361,I336378,I336418,I336440,I336457,I336483,I336491,I336508,I336525,I336542,I336559,I336604,I336635,I336652,I336678,I336686,I336717,I336734,I336751,I336768,I336840,I336866,I336874,I336914,I336922,I336939,I336956,I336996,I337018,I337035,I337061,I337069,I337086,I337103,I337120,I337137,I337182,I337213,I337230,I337256,I337264,I337295,I337312,I337329,I337346,I337418,I337444,I337452,I337401,I337492,I337500,I337517,I337534,I337389,I337574,I337410,I337596,I337613,I337639,I337647,I337664,I337681,I337698,I337715,I337386,I337407,I337760,I337398,I337791,I337808,I337834,I337842,I337404,I337873,I337890,I337907,I337924,I337395,I337392,I337996,I338022,I338030,I337979,I338070,I338078,I338095,I338112,I337967,I338152,I337988,I338174,I338191,I338217,I338225,I338242,I338259,I338276,I338293,I337964,I337985,I338338,I337976,I338369,I338386,I338412,I338420,I337982,I338451,I338468,I338485,I338502,I337973,I337970,I338574,I338600,I338608,I338648,I338656,I338673,I338690,I338730,I338752,I338769,I338795,I338803,I338820,I338837,I338854,I338871,I338916,I338947,I338964,I338990,I338998,I339029,I339046,I339063,I339080,I339152,I339178,I339186,I339226,I339234,I339251,I339268,I339308,I339330,I339347,I339373,I339381,I339398,I339415,I339432,I339449,I339494,I339525,I339542,I339568,I339576,I339607,I339624,I339641,I339658,I339730,I339756,I339764,I339804,I339812,I339829,I339846,I339886,I339908,I339925,I339951,I339959,I339976,I339993,I340010,I340027,I340072,I340103,I340120,I340146,I340154,I340185,I340202,I340219,I340236,I340308,I378910,I340334,I340342,I378892,I378883,I340382,I340390,I378898,I340407,I378886,I340424,I340464,I340486,I378895,I340503,I340529,I340537,I340554,I378904,I340571,I340588,I340605,I340650,I378907,I340681,I340698,I378901,I378889,I340724,I340732,I340763,I340780,I340797,I340814,I340886,I340912,I340920,I340960,I340968,I340985,I341002,I341042,I341064,I341081,I341107,I341115,I341132,I341149,I341166,I341183,I341228,I341259,I341276,I341302,I341310,I341341,I341358,I341375,I341392,I341464,I341490,I341498,I341538,I341546,I341563,I341580,I341620,I341642,I341659,I341685,I341693,I341710,I341727,I341744,I341761,I341806,I341837,I341854,I341880,I341888,I341919,I341936,I341953,I341970,I342042,I342068,I342076,I342116,I342124,I342141,I342158,I342198,I342220,I342237,I342263,I342271,I342288,I342305,I342322,I342339,I342384,I342415,I342432,I342458,I342466,I342497,I342514,I342531,I342548,I342620,I342646,I342654,I342694,I342702,I342719,I342736,I342776,I342798,I342815,I342841,I342849,I342866,I342883,I342900,I342917,I342962,I342993,I343010,I343036,I343044,I343075,I343092,I343109,I343126,I343198,I343224,I343232,I343258,I343275,I343297,I343314,I343331,I343348,I343365,I343396,I343413,I343430,I343447,I343492,I343509,I343526,I343585,I343611,I343619,I343636,I343653,I343684,I343742,I343768,I343776,I343802,I343819,I343841,I343858,I343875,I343892,I343909,I343940,I343957,I343974,I343991,I344036,I344053,I344070,I344129,I344155,I344163,I344180,I344197,I344228,I344286,I344312,I344320,I344346,I344363,I344385,I344402,I344419,I344436,I344453,I344484,I344501,I344518,I344535,I344580,I344597,I344614,I344673,I344699,I344707,I344724,I344741,I344772,I344830,I344856,I344864,I344890,I344907,I344929,I344946,I344963,I344980,I344997,I345028,I345045,I345062,I345079,I345124,I345141,I345158,I345217,I345243,I345251,I345268,I345285,I345316,I345374,I345400,I345408,I345434,I345451,I345473,I345490,I345507,I345524,I345541,I345572,I345589,I345606,I345623,I345668,I345685,I345702,I345761,I345787,I345795,I345812,I345829,I345860,I345918,I345944,I345952,I345978,I345995,I346017,I346034,I346051,I346068,I346085,I346116,I346133,I346150,I346167,I346212,I346229,I346246,I346305,I346331,I346339,I346356,I346373,I346404,I346462,I346488,I346496,I346522,I346539,I346561,I346578,I346595,I346612,I346629,I346660,I346677,I346694,I346711,I346756,I346773,I346790,I346849,I346875,I346883,I346900,I346917,I346948,I347006,I347032,I347040,I347066,I347083,I347105,I347122,I347139,I347156,I347173,I347204,I347221,I347238,I347255,I347300,I347317,I347334,I347393,I347419,I347427,I347444,I347461,I347492,I347550,I347576,I347584,I347610,I347627,I347649,I347666,I347683,I347700,I347717,I347748,I347765,I347782,I347799,I347844,I347861,I347878,I347937,I347963,I347971,I347988,I348005,I348036,I348094,I348120,I348128,I348154,I348171,I348193,I348210,I348227,I348244,I348261,I348292,I348309,I348326,I348343,I348388,I348405,I348422,I348481,I348507,I348515,I348532,I348549,I348580,I348638,I348664,I348672,I348698,I348715,I348737,I348754,I348771,I348788,I348805,I348836,I348853,I348870,I348887,I348932,I348949,I348966,I349025,I349051,I349059,I349076,I349093,I349124,I349182,I349208,I349216,I349242,I349259,I349281,I349298,I349315,I349332,I349349,I349380,I349397,I349414,I349431,I349476,I349493,I349510,I349569,I349595,I349603,I349620,I349637,I349668,I349726,I349752,I349760,I349786,I349803,I349718,I349825,I349842,I349859,I349876,I349893,I349697,I349924,I349941,I349958,I349975,I349700,I349715,I350020,I350037,I350054,I349712,I349709,I349706,I350113,I350139,I350147,I350164,I350181,I349694,I350212,I349703,I350270,I356775,I350296,I350304,I356784,I356787,I350330,I350347,I350369,I356781,I350386,I356778,I350403,I356772,I350420,I350437,I350468,I356769,I350485,I356766,I350502,I350519,I350564,I350581,I350598,I350657,I356790,I350683,I350691,I350708,I350725,I350756,I350814,I350840,I350848,I350874,I350891,I350913,I350930,I350947,I350964,I350981,I351012,I351029,I351046,I351063,I351108,I351125,I351142,I351201,I351227,I351235,I351252,I351269,I351300,I351358,I351384,I351392,I351418,I351435,I351457,I351474,I351491,I351508,I351525,I351556,I351573,I351590,I351607,I351652,I351669,I351686,I351745,I351771,I351779,I351796,I351813,I351844,I351902,I351928,I351936,I351962,I351979,I352001,I352018,I352035,I352052,I352069,I352100,I352117,I352134,I352151,I352196,I352213,I352230,I352289,I352315,I352323,I352340,I352357,I352388,I352446,I363133,I352472,I352480,I363142,I363145,I352506,I352523,I352545,I363139,I352562,I363136,I352579,I363130,I352596,I352613,I352644,I363127,I352661,I363124,I352678,I352695,I352740,I352757,I352774,I352833,I363148,I352859,I352867,I352884,I352901,I352932,I352990,I353016,I353024,I353050,I353067,I353089,I353106,I353123,I353140,I353157,I353188,I353205,I353222,I353239,I353284,I353301,I353318,I353377,I353403,I353411,I353428,I353445,I353476,I353534,I353560,I353568,I353594,I353611,I353633,I353650,I353667,I353684,I353701,I353732,I353749,I353766,I353783,I353828,I353845,I353862,I353921,I353947,I353955,I353972,I353989,I354020,I354078,I354104,I354112,I354138,I354155,I354177,I354194,I354211,I354228,I354245,I354276,I354293,I354310,I354327,I354372,I354389,I354406,I354465,I354491,I354499,I354516,I354533,I354564,I354622,I354648,I354656,I354682,I354699,I354721,I354738,I354755,I354772,I354789,I354820,I354837,I354854,I354871,I354916,I354933,I354950,I355009,I355035,I355043,I355060,I355077,I355108,I355166,I355192,I355200,I355226,I355243,I355265,I355282,I355299,I355316,I355333,I355364,I355381,I355398,I355415,I355460,I355477,I355494,I355553,I355579,I355587,I355604,I355621,I355652,I355710,I355736,I355744,I355770,I355787,I355809,I355826,I355843,I355860,I355877,I355908,I355925,I355942,I355959,I356004,I356021,I356038,I356097,I356123,I356131,I356148,I356165,I356196,I356254,I356280,I356288,I356314,I356331,I356353,I356370,I356387,I356404,I356421,I356452,I356469,I356486,I356503,I356548,I356565,I356582,I356641,I356667,I356675,I356692,I356709,I356740,I356798,I356824,I356832,I356849,I356875,I356883,I356900,I356917,I356934,I356951,I356982,I356999,I357016,I357047,I357064,I357104,I357112,I357143,I357160,I357177,I357194,I357225,I357256,I357282,I357304,I357376,I357402,I357410,I357427,I357453,I357461,I357478,I357495,I357512,I357529,I357560,I357577,I357594,I357625,I357642,I357682,I357690,I357721,I357738,I357755,I357772,I357803,I357834,I357860,I357882,I357954,I357980,I357988,I358005,I358031,I358039,I358056,I358073,I358090,I358107,I358138,I358155,I358172,I358203,I358220,I358260,I358268,I358299,I358316,I358333,I358350,I358381,I358412,I358438,I358460,I358532,I358558,I358566,I358583,I358609,I358617,I358634,I358651,I358668,I358685,I358716,I358733,I358750,I358781,I358798,I358838,I358846,I358877,I358894,I358911,I358928,I358959,I358990,I359016,I359038,I359110,I359136,I359144,I359161,I359187,I359195,I359212,I359229,I359246,I359263,I359294,I359311,I359328,I359359,I359376,I359416,I359424,I359455,I359472,I359489,I359506,I359537,I359568,I359594,I359616,I359688,I359714,I359722,I359739,I359765,I359773,I359790,I359807,I359824,I359841,I359872,I359889,I359906,I359937,I359954,I359994,I360002,I360033,I360050,I360067,I360084,I360115,I360146,I360172,I360194,I360266,I360292,I360300,I360317,I360343,I360351,I360368,I360385,I360402,I360419,I360450,I360467,I360484,I360515,I360532,I360572,I360580,I360611,I360628,I360645,I360662,I360693,I360724,I360750,I360772,I360844,I360870,I360878,I360895,I360921,I360929,I360946,I360963,I360980,I360997,I360836,I361028,I361045,I361062,I360815,I361093,I361110,I360821,I361150,I361158,I360830,I361189,I361206,I361223,I361240,I360833,I361271,I360812,I361302,I361328,I360827,I361350,I360824,I360818,I361422,I361448,I361456,I361473,I361499,I361507,I361524,I361541,I361558,I361575,I361606,I361623,I361640,I361671,I361688,I361728,I361736,I361767,I361784,I361801,I361818,I361849,I361880,I361906,I361928,I362000,I362026,I362034,I362051,I362077,I362085,I362102,I362119,I362136,I362153,I361992,I362184,I362201,I362218,I361971,I362249,I362266,I361977,I362306,I362314,I361986,I362345,I362362,I362379,I362396,I361989,I362427,I361968,I362458,I362484,I361983,I362506,I361980,I361974,I362578,I362604,I362612,I362629,I362655,I362663,I362680,I362697,I362714,I362731,I362762,I362779,I362796,I362827,I362844,I362884,I362892,I362923,I362940,I362957,I362974,I363005,I363036,I363062,I363084,I363156,I363182,I363190,I363207,I363233,I363241,I363258,I363275,I363292,I363309,I363340,I363357,I363374,I363405,I363422,I363462,I363470,I363501,I363518,I363535,I363552,I363583,I363614,I363640,I363662,I363734,I363760,I363768,I363785,I363811,I363819,I363836,I363853,I363870,I363887,I363918,I363935,I363952,I363983,I364000,I364040,I364048,I364079,I364096,I364113,I364130,I364161,I364192,I364218,I364240,I364312,I364338,I364346,I364363,I364389,I364397,I364414,I364431,I364448,I364465,I364496,I364513,I364530,I364561,I364578,I364618,I364626,I364657,I364674,I364691,I364708,I364739,I364770,I364796,I364818,I364890,I364916,I364924,I364941,I364967,I364975,I364992,I365009,I365026,I365043,I365074,I365091,I365108,I365139,I365156,I365196,I365204,I365235,I365252,I365269,I365286,I365317,I365348,I365374,I365396,I365468,I365494,I365502,I365519,I365545,I365553,I365570,I365587,I365604,I365621,I365652,I365669,I365686,I365717,I365734,I365774,I365782,I365813,I365830,I365847,I365864,I365895,I365926,I365952,I365974,I366046,I366072,I366080,I366097,I366123,I366131,I366148,I366165,I366182,I366199,I366230,I366247,I366264,I366295,I366312,I366352,I366360,I366391,I366408,I366425,I366442,I366473,I366504,I366530,I366552,I366624,I366650,I366658,I366675,I366701,I366709,I366726,I366743,I366760,I366777,I366808,I366825,I366842,I366873,I366890,I366930,I366938,I366969,I366986,I367003,I367020,I367051,I367082,I367108,I367130,I367202,I367228,I367236,I367253,I367279,I367287,I367304,I367321,I367338,I367355,I367386,I367403,I367420,I367451,I367468,I367508,I367516,I367547,I367564,I367581,I367598,I367629,I367660,I367686,I367708,I367780,I367806,I367814,I367831,I367857,I367865,I367882,I367899,I367916,I367933,I367772,I367964,I367981,I367998,I367751,I368029,I368046,I367757,I368086,I368094,I367766,I368125,I368142,I368159,I368176,I367769,I368207,I367748,I368238,I368264,I367763,I368286,I367760,I367754,I368358,I368384,I368392,I368409,I368435,I368443,I368460,I368477,I368494,I368511,I368542,I368559,I368576,I368607,I368624,I368664,I368672,I368703,I368720,I368737,I368754,I368785,I368816,I368842,I368864,I368939,I368965,I368973,I368990,I369016,I369024,I369041,I369058,I369089,I369120,I369137,I369154,I369171,I369188,I369219,I369278,I369295,I369321,I369343,I369369,I369377,I369394,I369425,I369500,I369526,I369534,I369551,I369577,I369585,I369602,I369619,I369650,I369681,I369698,I369715,I369732,I369749,I369780,I369839,I369856,I369882,I369904,I369930,I369938,I369955,I369986,I370061,I370087,I370095,I370112,I370138,I370146,I370163,I370180,I370211,I370242,I370259,I370276,I370293,I370310,I370341,I370400,I370417,I370443,I370465,I370491,I370499,I370516,I370547,I370622,I370648,I370656,I370673,I370699,I370707,I370724,I370741,I370772,I370803,I370820,I370837,I370854,I370871,I370902,I370961,I370978,I371004,I371026,I371052,I371060,I371077,I371108,I371183,I371209,I371226,I371234,I371279,I371296,I371313,I371330,I371347,I371364,I371381,I371412,I371429,I371474,I371491,I371508,I371539,I371565,I371573,I371604,I371621,I371638,I371664,I371672,I371689,I371778,I371804,I371821,I371829,I371874,I371891,I371908,I371925,I371942,I371959,I371976,I372007,I372024,I372069,I372086,I372103,I372134,I372160,I372168,I372199,I372216,I372233,I372259,I372267,I372284,I372373,I372399,I372416,I372424,I372469,I372486,I372503,I372520,I372537,I372554,I372571,I372602,I372619,I372664,I372681,I372698,I372729,I372755,I372763,I372794,I372811,I372828,I372854,I372862,I372879,I372968,I372994,I373011,I373019,I373064,I373081,I373098,I373115,I373132,I373149,I373166,I373197,I373214,I373259,I373276,I373293,I373324,I373350,I373358,I373389,I373406,I373423,I373449,I373457,I373474,I373563,I373589,I373606,I373614,I373659,I373676,I373693,I373710,I373727,I373744,I373761,I373792,I373809,I373854,I373871,I373888,I373919,I373945,I373953,I373984,I374001,I374018,I374044,I374052,I374069,I374158,I374184,I374201,I374209,I374254,I374271,I374288,I374305,I374322,I374339,I374356,I374387,I374404,I374449,I374466,I374483,I374514,I374540,I374548,I374579,I374596,I374613,I374639,I374647,I374664,I374753,I374779,I374796,I374804,I374849,I374866,I374883,I374900,I374917,I374934,I374951,I374982,I374999,I375044,I375061,I375078,I375109,I375135,I375143,I375174,I375191,I375208,I375234,I375242,I375259,I375348,I375374,I375391,I375399,I375444,I375461,I375478,I375495,I375512,I375529,I375546,I375577,I375594,I375639,I375656,I375673,I375704,I375730,I375738,I375769,I375786,I375803,I375829,I375837,I375854,I375943,I375969,I375986,I375994,I376039,I376056,I376073,I376090,I376107,I376124,I376141,I376172,I376189,I376234,I376251,I376268,I376299,I376325,I376333,I376364,I376381,I376398,I376424,I376432,I376449,I376538,I376564,I376581,I376589,I376634,I376651,I376668,I376685,I376702,I376719,I376736,I376767,I376784,I376829,I376846,I376863,I376894,I376920,I376928,I376959,I376976,I376993,I377019,I377027,I377044,I377133,I377159,I377176,I377184,I377229,I377246,I377263,I377280,I377297,I377314,I377331,I377362,I377379,I377424,I377441,I377458,I377489,I377515,I377523,I377554,I377571,I377588,I377614,I377622,I377639,I377728,I377754,I377771,I377779,I377824,I377841,I377858,I377875,I377892,I377909,I377926,I377957,I377974,I378019,I378036,I378053,I378084,I378110,I378118,I378149,I378166,I378183,I378209,I378217,I378234,I378323,I378349,I378366,I378374,I378419,I378436,I378453,I378470,I378487,I378504,I378521,I378552,I378569,I378614,I378631,I378648,I378679,I378705,I378713,I378744,I378761,I378778,I378804,I378812,I378829,I378918,I378944,I378961,I378969,I379014,I379031,I379048,I379065,I379082,I379099,I379116,I379147,I379164,I379209,I379226,I379243,I379274,I379300,I379308,I379339,I379356,I379373,I379399,I379407,I379424,I379513,I379539,I379556,I379564,I379609,I379626,I379643,I379660,I379677,I379694,I379711,I379742,I379759,I379804,I379821,I379838,I379869,I379895,I379903,I379934,I379951,I379968,I379994,I380002,I380019,I380108,I380134,I380151,I380159,I380204,I380221,I380238,I380255,I380272,I380289,I380306,I380337,I380354,I380399,I380416,I380433,I380464,I380490,I380498,I380529,I380546,I380563,I380589,I380597,I380614,I380703,I380729,I380746,I380754,I380799,I380816,I380833,I380850,I380867,I380884,I380901,I380932,I380949,I380994,I381011,I381028,I381059,I381085,I381093,I381124,I381141,I381158,I381184,I381192,I381209,I381298,I381324,I381341,I381349,I381394,I381411,I381428,I381445,I381462,I381479,I381496,I381527,I381544,I381589,I381606,I381623,I381654,I381680,I381688,I381719,I381736,I381753,I381779,I381787,I381804,I381893,I381919,I381936,I381944,I381989,I382006,I382023,I382040,I382057,I382074,I382091,I382122,I382139,I382184,I382201,I382218,I382249,I382275,I382283,I382314,I382331,I382348,I382374,I382382,I382399,I382488,I382514,I382531,I382539,I382584,I382601,I382618,I382635,I382652,I382669,I382686,I382717,I382734,I382779,I382796,I382813,I382844,I382870,I382878,I382909,I382926,I382943,I382969,I382977,I382994,I383083,I383109,I383126,I383134,I383179,I383196,I383213,I383230,I383247,I383264,I383281,I383312,I383329,I383374,I383391,I383408,I383439,I383465,I383473,I383504,I383521,I383538,I383564,I383572,I383589,I383678,I383704,I383721,I383729,I383774,I383791,I383808,I383825,I383842,I383859,I383876,I383907,I383924,I383969,I383986,I384003,I384034,I384060,I384068,I384099,I384116,I384133,I384159,I384167,I384184,I384273,I384299,I384316,I384324,I384369,I384386,I384403,I384420,I384437,I384454,I384471,I384502,I384519,I384564,I384581,I384598,I384629,I384655,I384663,I384694,I384711,I384728,I384754,I384762,I384779,I384868,I384894,I384911,I384919,I384964,I384981,I384998,I385015,I385032,I385049,I385066,I385097,I385114,I385159,I385176,I385193,I385224,I385250,I385258,I385289,I385306,I385323,I385349,I385357,I385374,I385463,I385489,I385506,I385514,I385559,I385576,I385593,I385610,I385627,I385644,I385661,I385692,I385709,I385754,I385771,I385788,I385819,I385845,I385853,I385884,I385901,I385918,I385944,I385952,I385969,I386058,I386084,I386101,I386109,I386154,I386171,I386188,I386205,I386222,I386239,I386256,I386287,I386304,I386349,I386366,I386383,I386414,I386440,I386448,I386479,I386496,I386513,I386539,I386547,I386564,I386653,I386679,I386696,I386704,I386749,I386766,I386783,I386800,I386817,I386834,I386851,I386882,I386899,I386944,I386961,I386978,I387009,I387035,I387043,I387074,I387091,I387108,I387134,I387142,I387159,I387248,I387274,I387291,I387299,I387344,I387361,I387378,I387395,I387412,I387429,I387446,I387477,I387494,I387539,I387556,I387573,I387604,I387630,I387638,I387669,I387686,I387703,I387729,I387737,I387754,I387843,I387869,I387886,I387894,I387939,I387956,I387973,I387990,I388007,I388024,I388041,I388072,I388089,I388134,I388151,I388168,I388199,I388225,I388233,I388264,I388281,I388298,I388324,I388332,I388349,I388438,I388464,I388481,I388489,I388534,I388551,I388568,I388585,I388602,I388619,I388636,I388667,I388684,I388729,I388746,I388763,I388794,I388820,I388828,I388859,I388876,I388893,I388919,I388927,I388944,I389033,I389059,I389076,I389084,I389129,I389146,I389163,I389180,I389197,I389214,I389231,I389262,I389279,I389324,I389341,I389358,I389389,I389415,I389423,I389454,I389471,I389488,I389514,I389522,I389539,I389628,I389654,I389671,I389679,I389724,I389741,I389758,I389775,I389792,I389809,I389826,I389857,I389874,I389919,I389936,I389953,I389984,I390010,I390018,I390049,I390066,I390083,I390109,I390117,I390134,I390223,I390249,I390266,I390274,I390319,I390336,I390353,I390370,I390387,I390404,I390421,I390452,I390469,I390514,I390531,I390548,I390579,I390605,I390613,I390644,I390661,I390678,I390704,I390712,I390729,I390818,I390844,I390861,I390869,I390914,I390931,I390948,I390965,I390982,I390999,I391016,I391047,I391064,I391109,I391126,I391143,I391174,I391200,I391208,I391239,I391256,I391273,I391299,I391307,I391324,I391413,I391439,I391456,I391464,I391509,I391526,I391543,I391560,I391577,I391594,I391611,I391642,I391659,I391704,I391721,I391738,I391769,I391795,I391803,I391834,I391851,I391868,I391894,I391902,I391919,I392008,I392034,I392051,I392059,I392104,I392121,I392138,I392155,I392172,I392189,I392206,I392237,I392254,I392299,I392316,I392333,I392364,I392390,I392398,I392429,I392446,I392463,I392489,I392497,I392514,I392603,I392629,I392646,I392654,I392699,I392716,I392733,I392750,I392767,I392784,I392801,I392832,I392849,I392894,I392911,I392928,I392959,I392985,I392993,I393024,I393041,I393058,I393084,I393092,I393109;
not I_0 (I2634,I2602);
DFFARX1 I_1 (I185940,I2595,I2634,I2660,);
nand I_2 (I2668,I2660,I185919);
not I_3 (I2685,I2668);
DFFARX1 I_4 (I2685,I2595,I2634,I2626,);
DFFARX1 I_5 (I185928,I2595,I2634,I2725,);
not I_6 (I2733,I2725);
not I_7 (I2750,I185934);
not I_8 (I2767,I185931);
nand I_9 (I2784,I2733,I2767);
nor I_10 (I2801,I2784,I185934);
DFFARX1 I_11 (I2801,I2595,I2634,I2605,);
nor I_12 (I2832,I185931,I185934);
nand I_13 (I2849,I2725,I2832);
nor I_14 (I2866,I185922,I185916);
nor I_15 (I2608,I2784,I185922);
not I_16 (I2897,I185922);
not I_17 (I2914,I185937);
nand I_18 (I2931,I2914,I185919);
nand I_19 (I2948,I2750,I2931);
not I_20 (I2965,I2948);
nor I_21 (I2982,I185937,I185916);
nor I_22 (I2617,I2965,I2982);
nor I_23 (I3013,I185925,I185937);
and I_24 (I3030,I3013,I2866);
nor I_25 (I3047,I2948,I3030);
DFFARX1 I_26 (I3047,I2595,I2634,I2623,);
nor I_27 (I3078,I2668,I3030);
DFFARX1 I_28 (I3078,I2595,I2634,I2620,);
nor I_29 (I3109,I185925,I185916);
DFFARX1 I_30 (I3109,I2595,I2634,I3135,);
nor I_31 (I3143,I3135,I185931);
nand I_32 (I3160,I3143,I2750);
nand I_33 (I2614,I3160,I2849);
nand I_34 (I2611,I3143,I2897);
not I_35 (I3229,I2602);
DFFARX1 I_36 (I339701,I2595,I3229,I3255,);
nand I_37 (I3263,I3255,I339701);
not I_38 (I3280,I3263);
DFFARX1 I_39 (I3280,I2595,I3229,I3221,);
DFFARX1 I_40 (I339716,I2595,I3229,I3320,);
not I_41 (I3328,I3320);
not I_42 (I3345,I339713);
not I_43 (I3362,I339722);
nand I_44 (I3379,I3328,I3362);
nor I_45 (I3396,I3379,I339713);
DFFARX1 I_46 (I3396,I2595,I3229,I3200,);
nor I_47 (I3427,I339722,I339713);
nand I_48 (I3444,I3320,I3427);
nor I_49 (I3461,I339710,I339719);
nor I_50 (I3203,I3379,I339710);
not I_51 (I3492,I339710);
not I_52 (I3509,I339707);
nand I_53 (I3526,I3509,I339698);
nand I_54 (I3543,I3345,I3526);
not I_55 (I3560,I3543);
nor I_56 (I3577,I339707,I339719);
nor I_57 (I3212,I3560,I3577);
nor I_58 (I3608,I339704,I339707);
and I_59 (I3625,I3608,I3461);
nor I_60 (I3642,I3543,I3625);
DFFARX1 I_61 (I3642,I2595,I3229,I3218,);
nor I_62 (I3673,I3263,I3625);
DFFARX1 I_63 (I3673,I2595,I3229,I3215,);
nor I_64 (I3704,I339704,I339698);
DFFARX1 I_65 (I3704,I2595,I3229,I3730,);
nor I_66 (I3738,I3730,I339722);
nand I_67 (I3755,I3738,I3345);
nand I_68 (I3209,I3755,I3444);
nand I_69 (I3206,I3738,I3492);
not I_70 (I3824,I2602);
DFFARX1 I_71 (I346454,I2595,I3824,I3850,);
nand I_72 (I3858,I3850,I346442);
not I_73 (I3875,I3858);
DFFARX1 I_74 (I3875,I2595,I3824,I3816,);
DFFARX1 I_75 (I346430,I2595,I3824,I3915,);
not I_76 (I3923,I3915);
not I_77 (I3940,I346430);
not I_78 (I3957,I346436);
nand I_79 (I3974,I3923,I3957);
nor I_80 (I3991,I3974,I346430);
DFFARX1 I_81 (I3991,I2595,I3824,I3795,);
nor I_82 (I4022,I346436,I346430);
nand I_83 (I4039,I3915,I4022);
nor I_84 (I4056,I346433,I346448);
nor I_85 (I3798,I3974,I346433);
not I_86 (I4087,I346433);
not I_87 (I4104,I346439);
nand I_88 (I4121,I4104,I346451);
nand I_89 (I4138,I3940,I4121);
not I_90 (I4155,I4138);
nor I_91 (I4172,I346439,I346448);
nor I_92 (I3807,I4155,I4172);
nor I_93 (I4203,I346445,I346439);
and I_94 (I4220,I4203,I4056);
nor I_95 (I4237,I4138,I4220);
DFFARX1 I_96 (I4237,I2595,I3824,I3813,);
nor I_97 (I4268,I3858,I4220);
DFFARX1 I_98 (I4268,I2595,I3824,I3810,);
nor I_99 (I4299,I346445,I346433);
DFFARX1 I_100 (I4299,I2595,I3824,I4325,);
nor I_101 (I4333,I4325,I346436);
nand I_102 (I4350,I4333,I3940);
nand I_103 (I3804,I4350,I4039);
nand I_104 (I3801,I4333,I4087);
not I_105 (I4419,I2602);
DFFARX1 I_106 (I100659,I2595,I4419,I4445,);
nand I_107 (I4453,I4445,I100650);
not I_108 (I4470,I4453);
DFFARX1 I_109 (I4470,I2595,I4419,I4411,);
DFFARX1 I_110 (I100653,I2595,I4419,I4510,);
not I_111 (I4518,I4510);
not I_112 (I4535,I100647);
not I_113 (I4552,I100656);
nand I_114 (I4569,I4518,I4552);
nor I_115 (I4586,I4569,I100647);
DFFARX1 I_116 (I4586,I2595,I4419,I4390,);
nor I_117 (I4617,I100656,I100647);
nand I_118 (I4634,I4510,I4617);
nor I_119 (I4651,I100644,I100662);
nor I_120 (I4393,I4569,I100644);
not I_121 (I4682,I100644);
not I_122 (I4699,I100644);
nand I_123 (I4716,I4699,I100668);
nand I_124 (I4733,I4535,I4716);
not I_125 (I4750,I4733);
nor I_126 (I4767,I100644,I100662);
nor I_127 (I4402,I4750,I4767);
nor I_128 (I4798,I100665,I100644);
and I_129 (I4815,I4798,I4651);
nor I_130 (I4832,I4733,I4815);
DFFARX1 I_131 (I4832,I2595,I4419,I4408,);
nor I_132 (I4863,I4453,I4815);
DFFARX1 I_133 (I4863,I2595,I4419,I4405,);
nor I_134 (I4894,I100665,I100671);
DFFARX1 I_135 (I4894,I2595,I4419,I4920,);
nor I_136 (I4928,I4920,I100656);
nand I_137 (I4945,I4928,I4535);
nand I_138 (I4399,I4945,I4634);
nand I_139 (I4396,I4928,I4682);
not I_140 (I5014,I2602);
DFFARX1 I_141 (I82741,I2595,I5014,I5040,);
nand I_142 (I5048,I5040,I82732);
not I_143 (I5065,I5048);
DFFARX1 I_144 (I5065,I2595,I5014,I5006,);
DFFARX1 I_145 (I82735,I2595,I5014,I5105,);
not I_146 (I5113,I5105);
not I_147 (I5130,I82729);
not I_148 (I5147,I82738);
nand I_149 (I5164,I5113,I5147);
nor I_150 (I5181,I5164,I82729);
DFFARX1 I_151 (I5181,I2595,I5014,I4985,);
nor I_152 (I5212,I82738,I82729);
nand I_153 (I5229,I5105,I5212);
nor I_154 (I5246,I82726,I82744);
nor I_155 (I4988,I5164,I82726);
not I_156 (I5277,I82726);
not I_157 (I5294,I82726);
nand I_158 (I5311,I5294,I82750);
nand I_159 (I5328,I5130,I5311);
not I_160 (I5345,I5328);
nor I_161 (I5362,I82726,I82744);
nor I_162 (I4997,I5345,I5362);
nor I_163 (I5393,I82747,I82726);
and I_164 (I5410,I5393,I5246);
nor I_165 (I5427,I5328,I5410);
DFFARX1 I_166 (I5427,I2595,I5014,I5003,);
nor I_167 (I5458,I5048,I5410);
DFFARX1 I_168 (I5458,I2595,I5014,I5000,);
nor I_169 (I5489,I82747,I82753);
DFFARX1 I_170 (I5489,I2595,I5014,I5515,);
nor I_171 (I5523,I5515,I82738);
nand I_172 (I5540,I5523,I5130);
nand I_173 (I4994,I5540,I5229);
nand I_174 (I4991,I5523,I5277);
not I_175 (I5609,I2602);
DFFARX1 I_176 (I335655,I2595,I5609,I5635,);
nand I_177 (I5643,I5635,I335655);
not I_178 (I5660,I5643);
DFFARX1 I_179 (I5660,I2595,I5609,I5601,);
DFFARX1 I_180 (I335670,I2595,I5609,I5700,);
not I_181 (I5708,I5700);
not I_182 (I5725,I335667);
not I_183 (I5742,I335676);
nand I_184 (I5759,I5708,I5742);
nor I_185 (I5776,I5759,I335667);
DFFARX1 I_186 (I5776,I2595,I5609,I5580,);
nor I_187 (I5807,I335676,I335667);
nand I_188 (I5824,I5700,I5807);
nor I_189 (I5841,I335664,I335673);
nor I_190 (I5583,I5759,I335664);
not I_191 (I5872,I335664);
not I_192 (I5889,I335661);
nand I_193 (I5906,I5889,I335652);
nand I_194 (I5923,I5725,I5906);
not I_195 (I5940,I5923);
nor I_196 (I5957,I335661,I335673);
nor I_197 (I5592,I5940,I5957);
nor I_198 (I5988,I335658,I335661);
and I_199 (I6005,I5988,I5841);
nor I_200 (I6022,I5923,I6005);
DFFARX1 I_201 (I6022,I2595,I5609,I5598,);
nor I_202 (I6053,I5643,I6005);
DFFARX1 I_203 (I6053,I2595,I5609,I5595,);
nor I_204 (I6084,I335658,I335652);
DFFARX1 I_205 (I6084,I2595,I5609,I6110,);
nor I_206 (I6118,I6110,I335676);
nand I_207 (I6135,I6118,I5725);
nand I_208 (I5589,I6135,I5824);
nand I_209 (I5586,I6118,I5872);
not I_210 (I6204,I2602);
DFFARX1 I_211 (I154670,I2595,I6204,I6230,);
nand I_212 (I6238,I6230,I154691);
not I_213 (I6255,I6238);
DFFARX1 I_214 (I6255,I2595,I6204,I6196,);
DFFARX1 I_215 (I154688,I2595,I6204,I6295,);
not I_216 (I6303,I6295);
not I_217 (I6320,I154670);
not I_218 (I6337,I154682);
nand I_219 (I6354,I6303,I6337);
nor I_220 (I6371,I6354,I154670);
DFFARX1 I_221 (I6371,I2595,I6204,I6175,);
nor I_222 (I6402,I154682,I154670);
nand I_223 (I6419,I6295,I6402);
nor I_224 (I6436,I154685,I154694);
nor I_225 (I6178,I6354,I154685);
not I_226 (I6467,I154685);
not I_227 (I6484,I154673);
nand I_228 (I6501,I6484,I154676);
nand I_229 (I6518,I6320,I6501);
not I_230 (I6535,I6518);
nor I_231 (I6552,I154673,I154694);
nor I_232 (I6187,I6535,I6552);
nor I_233 (I6583,I154673,I154673);
and I_234 (I6600,I6583,I6436);
nor I_235 (I6617,I6518,I6600);
DFFARX1 I_236 (I6617,I2595,I6204,I6193,);
nor I_237 (I6648,I6238,I6600);
DFFARX1 I_238 (I6648,I2595,I6204,I6190,);
nor I_239 (I6679,I154673,I154679);
DFFARX1 I_240 (I6679,I2595,I6204,I6705,);
nor I_241 (I6713,I6705,I154682);
nand I_242 (I6730,I6713,I6320);
nand I_243 (I6184,I6730,I6419);
nand I_244 (I6181,I6713,I6467);
not I_245 (I6799,I2602);
DFFARX1 I_246 (I360237,I2595,I6799,I6825,);
nand I_247 (I6833,I6825,I360243);
not I_248 (I6850,I6833);
DFFARX1 I_249 (I6850,I2595,I6799,I6791,);
DFFARX1 I_250 (I360246,I2595,I6799,I6890,);
not I_251 (I6898,I6890);
not I_252 (I6915,I360234);
not I_253 (I6932,I360252);
nand I_254 (I6949,I6898,I6932);
nor I_255 (I6966,I6949,I360234);
DFFARX1 I_256 (I6966,I2595,I6799,I6770,);
nor I_257 (I6997,I360252,I360234);
nand I_258 (I7014,I6890,I6997);
nor I_259 (I7031,I360249,I360258);
nor I_260 (I6773,I6949,I360249);
not I_261 (I7062,I360249);
not I_262 (I7079,I360237);
nand I_263 (I7096,I7079,I360255);
nand I_264 (I7113,I6915,I7096);
not I_265 (I7130,I7113);
nor I_266 (I7147,I360237,I360258);
nor I_267 (I6782,I7130,I7147);
nor I_268 (I7178,I360240,I360237);
and I_269 (I7195,I7178,I7031);
nor I_270 (I7212,I7113,I7195);
DFFARX1 I_271 (I7212,I2595,I6799,I6788,);
nor I_272 (I7243,I6833,I7195);
DFFARX1 I_273 (I7243,I2595,I6799,I6785,);
nor I_274 (I7274,I360240,I360234);
DFFARX1 I_275 (I7274,I2595,I6799,I7300,);
nor I_276 (I7308,I7300,I360252);
nand I_277 (I7325,I7308,I6915);
nand I_278 (I6779,I7325,I7014);
nand I_279 (I6776,I7308,I7062);
not I_280 (I7394,I2602);
DFFARX1 I_281 (I342591,I2595,I7394,I7420,);
nand I_282 (I7428,I7420,I342591);
not I_283 (I7445,I7428);
DFFARX1 I_284 (I7445,I2595,I7394,I7386,);
DFFARX1 I_285 (I342606,I2595,I7394,I7485,);
not I_286 (I7493,I7485);
not I_287 (I7510,I342603);
not I_288 (I7527,I342612);
nand I_289 (I7544,I7493,I7527);
nor I_290 (I7561,I7544,I342603);
DFFARX1 I_291 (I7561,I2595,I7394,I7365,);
nor I_292 (I7592,I342612,I342603);
nand I_293 (I7609,I7485,I7592);
nor I_294 (I7626,I342600,I342609);
nor I_295 (I7368,I7544,I342600);
not I_296 (I7657,I342600);
not I_297 (I7674,I342597);
nand I_298 (I7691,I7674,I342588);
nand I_299 (I7708,I7510,I7691);
not I_300 (I7725,I7708);
nor I_301 (I7742,I342597,I342609);
nor I_302 (I7377,I7725,I7742);
nor I_303 (I7773,I342594,I342597);
and I_304 (I7790,I7773,I7626);
nor I_305 (I7807,I7708,I7790);
DFFARX1 I_306 (I7807,I2595,I7394,I7383,);
nor I_307 (I7838,I7428,I7790);
DFFARX1 I_308 (I7838,I2595,I7394,I7380,);
nor I_309 (I7869,I342594,I342588);
DFFARX1 I_310 (I7869,I2595,I7394,I7895,);
nor I_311 (I7903,I7895,I342612);
nand I_312 (I7920,I7903,I7510);
nand I_313 (I7374,I7920,I7609);
nand I_314 (I7371,I7903,I7657);
not I_315 (I7989,I2602);
DFFARX1 I_316 (I277720,I2595,I7989,I8015,);
nand I_317 (I8023,I8015,I277711);
not I_318 (I8040,I8023);
DFFARX1 I_319 (I8040,I2595,I7989,I7981,);
DFFARX1 I_320 (I277714,I2595,I7989,I8080,);
not I_321 (I8088,I8080);
not I_322 (I8105,I277726);
not I_323 (I8122,I277705);
nand I_324 (I8139,I8088,I8122);
nor I_325 (I8156,I8139,I277726);
DFFARX1 I_326 (I8156,I2595,I7989,I7960,);
nor I_327 (I8187,I277705,I277726);
nand I_328 (I8204,I8080,I8187);
nor I_329 (I8221,I277717,I277723);
nor I_330 (I7963,I8139,I277717);
not I_331 (I8252,I277717);
not I_332 (I8269,I277708);
nand I_333 (I8286,I8269,I277699);
nand I_334 (I8303,I8105,I8286);
not I_335 (I8320,I8303);
nor I_336 (I8337,I277708,I277723);
nor I_337 (I7972,I8320,I8337);
nor I_338 (I8368,I277699,I277708);
and I_339 (I8385,I8368,I8221);
nor I_340 (I8402,I8303,I8385);
DFFARX1 I_341 (I8402,I2595,I7989,I7978,);
nor I_342 (I8433,I8023,I8385);
DFFARX1 I_343 (I8433,I2595,I7989,I7975,);
nor I_344 (I8464,I277699,I277702);
DFFARX1 I_345 (I8464,I2595,I7989,I8490,);
nor I_346 (I8498,I8490,I277705);
nand I_347 (I8515,I8498,I8105);
nand I_348 (I7969,I8515,I8204);
nand I_349 (I7966,I8498,I8252);
not I_350 (I8584,I2602);
DFFARX1 I_351 (I217730,I2595,I8584,I8610,);
nand I_352 (I8618,I8610,I217709);
not I_353 (I8635,I8618);
DFFARX1 I_354 (I8635,I2595,I8584,I8576,);
DFFARX1 I_355 (I217718,I2595,I8584,I8675,);
not I_356 (I8683,I8675);
not I_357 (I8700,I217724);
not I_358 (I8717,I217721);
nand I_359 (I8734,I8683,I8717);
nor I_360 (I8751,I8734,I217724);
DFFARX1 I_361 (I8751,I2595,I8584,I8555,);
nor I_362 (I8782,I217721,I217724);
nand I_363 (I8799,I8675,I8782);
nor I_364 (I8816,I217712,I217706);
nor I_365 (I8558,I8734,I217712);
not I_366 (I8847,I217712);
not I_367 (I8864,I217727);
nand I_368 (I8881,I8864,I217709);
nand I_369 (I8898,I8700,I8881);
not I_370 (I8915,I8898);
nor I_371 (I8932,I217727,I217706);
nor I_372 (I8567,I8915,I8932);
nor I_373 (I8963,I217715,I217727);
and I_374 (I8980,I8963,I8816);
nor I_375 (I8997,I8898,I8980);
DFFARX1 I_376 (I8997,I2595,I8584,I8573,);
nor I_377 (I9028,I8618,I8980);
DFFARX1 I_378 (I9028,I2595,I8584,I8570,);
nor I_379 (I9059,I217715,I217706);
DFFARX1 I_380 (I9059,I2595,I8584,I9085,);
nor I_381 (I9093,I9085,I217721);
nand I_382 (I9110,I9093,I8700);
nand I_383 (I8564,I9110,I8799);
nand I_384 (I8561,I9093,I8847);
not I_385 (I9179,I2602);
DFFARX1 I_386 (I32945,I2595,I9179,I9205,);
nand I_387 (I9213,I9205,I32936);
not I_388 (I9230,I9213);
DFFARX1 I_389 (I9230,I2595,I9179,I9171,);
DFFARX1 I_390 (I32957,I2595,I9179,I9270,);
not I_391 (I9278,I9270);
not I_392 (I9295,I32933);
not I_393 (I9312,I32933);
nand I_394 (I9329,I9278,I9312);
nor I_395 (I9346,I9329,I32933);
DFFARX1 I_396 (I9346,I2595,I9179,I9150,);
nor I_397 (I9377,I32933,I32933);
nand I_398 (I9394,I9270,I9377);
nor I_399 (I9411,I32942,I32936);
nor I_400 (I9153,I9329,I32942);
not I_401 (I9442,I32942);
not I_402 (I9459,I32954);
nand I_403 (I9476,I9459,I32951);
nand I_404 (I9493,I9295,I9476);
not I_405 (I9510,I9493);
nor I_406 (I9527,I32954,I32936);
nor I_407 (I9162,I9510,I9527);
nor I_408 (I9558,I32948,I32954);
and I_409 (I9575,I9558,I9411);
nor I_410 (I9592,I9493,I9575);
DFFARX1 I_411 (I9592,I2595,I9179,I9168,);
nor I_412 (I9623,I9213,I9575);
DFFARX1 I_413 (I9623,I2595,I9179,I9165,);
nor I_414 (I9654,I32948,I32939);
DFFARX1 I_415 (I9654,I2595,I9179,I9680,);
nor I_416 (I9688,I9680,I32933);
nand I_417 (I9705,I9688,I9295);
nand I_418 (I9159,I9705,I9394);
nand I_419 (I9156,I9688,I9442);
not I_420 (I9777,I2602);
DFFARX1 I_421 (I201528,I2595,I9777,I9803,);
DFFARX1 I_422 (I9803,I2595,I9777,I9820,);
not I_423 (I9828,I9820);
nand I_424 (I9845,I201543,I201546);
and I_425 (I9862,I9845,I201525);
DFFARX1 I_426 (I9862,I2595,I9777,I9888,);
DFFARX1 I_427 (I9888,I2595,I9777,I9769,);
DFFARX1 I_428 (I9888,I2595,I9777,I9760,);
DFFARX1 I_429 (I201531,I2595,I9777,I9933,);
nand I_430 (I9941,I9933,I201537);
not I_431 (I9958,I9941);
nor I_432 (I9757,I9803,I9958);
DFFARX1 I_433 (I201525,I2595,I9777,I9998,);
not I_434 (I10006,I9998);
nor I_435 (I9763,I10006,I9828);
nand I_436 (I9751,I10006,I9941);
nand I_437 (I10051,I201540,I201522);
and I_438 (I10068,I10051,I201534);
DFFARX1 I_439 (I10068,I2595,I9777,I10094,);
nor I_440 (I10102,I10094,I9803);
DFFARX1 I_441 (I10102,I2595,I9777,I9745,);
not I_442 (I10133,I10094);
nor I_443 (I10150,I201522,I201522);
not I_444 (I10167,I10150);
nor I_445 (I10184,I9941,I10167);
nor I_446 (I10201,I10133,I10184);
DFFARX1 I_447 (I10201,I2595,I9777,I9766,);
nor I_448 (I10232,I10094,I10167);
nor I_449 (I9754,I9958,I10232);
nor I_450 (I9748,I10094,I10150);
not I_451 (I10304,I2602);
DFFARX1 I_452 (I289894,I2595,I10304,I10330,);
DFFARX1 I_453 (I10330,I2595,I10304,I10347,);
not I_454 (I10355,I10347);
nand I_455 (I10372,I289888,I289909);
and I_456 (I10389,I10372,I289894);
DFFARX1 I_457 (I10389,I2595,I10304,I10415,);
DFFARX1 I_458 (I10415,I2595,I10304,I10296,);
DFFARX1 I_459 (I10415,I2595,I10304,I10287,);
DFFARX1 I_460 (I289891,I2595,I10304,I10460,);
nand I_461 (I10468,I10460,I289900);
not I_462 (I10485,I10468);
nor I_463 (I10284,I10330,I10485);
DFFARX1 I_464 (I289888,I2595,I10304,I10525,);
not I_465 (I10533,I10525);
nor I_466 (I10290,I10533,I10355);
nand I_467 (I10278,I10533,I10468);
nand I_468 (I10578,I289891,I289906);
and I_469 (I10595,I10578,I289897);
DFFARX1 I_470 (I10595,I2595,I10304,I10621,);
nor I_471 (I10629,I10621,I10330);
DFFARX1 I_472 (I10629,I2595,I10304,I10272,);
not I_473 (I10660,I10621);
nor I_474 (I10677,I289903,I289906);
not I_475 (I10694,I10677);
nor I_476 (I10711,I10468,I10694);
nor I_477 (I10728,I10660,I10711);
DFFARX1 I_478 (I10728,I2595,I10304,I10293,);
nor I_479 (I10759,I10621,I10694);
nor I_480 (I10281,I10485,I10759);
nor I_481 (I10275,I10621,I10677);
not I_482 (I10831,I2602);
DFFARX1 I_483 (I268679,I2595,I10831,I10857,);
DFFARX1 I_484 (I10857,I2595,I10831,I10874,);
not I_485 (I10882,I10874);
nand I_486 (I10899,I268655,I268682);
and I_487 (I10916,I10899,I268667);
DFFARX1 I_488 (I10916,I2595,I10831,I10942,);
DFFARX1 I_489 (I10942,I2595,I10831,I10823,);
DFFARX1 I_490 (I10942,I2595,I10831,I10814,);
DFFARX1 I_491 (I268673,I2595,I10831,I10987,);
nand I_492 (I10995,I10987,I268658);
not I_493 (I11012,I10995);
nor I_494 (I10811,I10857,I11012);
DFFARX1 I_495 (I268676,I2595,I10831,I11052,);
not I_496 (I11060,I11052);
nor I_497 (I10817,I11060,I10882);
nand I_498 (I10805,I11060,I10995);
nand I_499 (I11105,I268661,I268664);
and I_500 (I11122,I11105,I268655);
DFFARX1 I_501 (I11122,I2595,I10831,I11148,);
nor I_502 (I11156,I11148,I10857);
DFFARX1 I_503 (I11156,I2595,I10831,I10799,);
not I_504 (I11187,I11148);
nor I_505 (I11204,I268670,I268664);
not I_506 (I11221,I11204);
nor I_507 (I11238,I10995,I11221);
nor I_508 (I11255,I11187,I11238);
DFFARX1 I_509 (I11255,I2595,I10831,I10820,);
nor I_510 (I11286,I11148,I11221);
nor I_511 (I10808,I11012,I11286);
nor I_512 (I10802,I11148,I11204);
not I_513 (I11358,I2602);
DFFARX1 I_514 (I31882,I2595,I11358,I11384,);
DFFARX1 I_515 (I11384,I2595,I11358,I11401,);
not I_516 (I11409,I11401);
nand I_517 (I11426,I31882,I31897);
and I_518 (I11443,I11426,I31900);
DFFARX1 I_519 (I11443,I2595,I11358,I11469,);
DFFARX1 I_520 (I11469,I2595,I11358,I11350,);
DFFARX1 I_521 (I11469,I2595,I11358,I11341,);
DFFARX1 I_522 (I31894,I2595,I11358,I11514,);
nand I_523 (I11522,I11514,I31903);
not I_524 (I11539,I11522);
nor I_525 (I11338,I11384,I11539);
DFFARX1 I_526 (I31879,I2595,I11358,I11579,);
not I_527 (I11587,I11579);
nor I_528 (I11344,I11587,I11409);
nand I_529 (I11332,I11587,I11522);
nand I_530 (I11632,I31879,I31885);
and I_531 (I11649,I11632,I31888);
DFFARX1 I_532 (I11649,I2595,I11358,I11675,);
nor I_533 (I11683,I11675,I11384);
DFFARX1 I_534 (I11683,I2595,I11358,I11326,);
not I_535 (I11714,I11675);
nor I_536 (I11731,I31891,I31885);
not I_537 (I11748,I11731);
nor I_538 (I11765,I11522,I11748);
nor I_539 (I11782,I11714,I11765);
DFFARX1 I_540 (I11782,I2595,I11358,I11347,);
nor I_541 (I11813,I11675,I11748);
nor I_542 (I11335,I11539,I11813);
nor I_543 (I11329,I11675,I11731);
not I_544 (I11885,I2602);
DFFARX1 I_545 (I225226,I2595,I11885,I11911,);
DFFARX1 I_546 (I11911,I2595,I11885,I11928,);
not I_547 (I11936,I11928);
nand I_548 (I11953,I225241,I225244);
and I_549 (I11970,I11953,I225223);
DFFARX1 I_550 (I11970,I2595,I11885,I11996,);
DFFARX1 I_551 (I11996,I2595,I11885,I11877,);
DFFARX1 I_552 (I11996,I2595,I11885,I11868,);
DFFARX1 I_553 (I225229,I2595,I11885,I12041,);
nand I_554 (I12049,I12041,I225235);
not I_555 (I12066,I12049);
nor I_556 (I11865,I11911,I12066);
DFFARX1 I_557 (I225223,I2595,I11885,I12106,);
not I_558 (I12114,I12106);
nor I_559 (I11871,I12114,I11936);
nand I_560 (I11859,I12114,I12049);
nand I_561 (I12159,I225238,I225220);
and I_562 (I12176,I12159,I225232);
DFFARX1 I_563 (I12176,I2595,I11885,I12202,);
nor I_564 (I12210,I12202,I11911);
DFFARX1 I_565 (I12210,I2595,I11885,I11853,);
not I_566 (I12241,I12202);
nor I_567 (I12258,I225220,I225220);
not I_568 (I12275,I12258);
nor I_569 (I12292,I12049,I12275);
nor I_570 (I12309,I12241,I12292);
DFFARX1 I_571 (I12309,I2595,I11885,I11874,);
nor I_572 (I12340,I12202,I12275);
nor I_573 (I11862,I12066,I12340);
nor I_574 (I11856,I12202,I12258);
not I_575 (I12412,I2602);
DFFARX1 I_576 (I194014,I2595,I12412,I12438,);
DFFARX1 I_577 (I12438,I2595,I12412,I12455,);
not I_578 (I12463,I12455);
nand I_579 (I12480,I194029,I194032);
and I_580 (I12497,I12480,I194011);
DFFARX1 I_581 (I12497,I2595,I12412,I12523,);
DFFARX1 I_582 (I12523,I2595,I12412,I12404,);
DFFARX1 I_583 (I12523,I2595,I12412,I12395,);
DFFARX1 I_584 (I194017,I2595,I12412,I12568,);
nand I_585 (I12576,I12568,I194023);
not I_586 (I12593,I12576);
nor I_587 (I12392,I12438,I12593);
DFFARX1 I_588 (I194011,I2595,I12412,I12633,);
not I_589 (I12641,I12633);
nor I_590 (I12398,I12641,I12463);
nand I_591 (I12386,I12641,I12576);
nand I_592 (I12686,I194026,I194008);
and I_593 (I12703,I12686,I194020);
DFFARX1 I_594 (I12703,I2595,I12412,I12729,);
nor I_595 (I12737,I12729,I12438);
DFFARX1 I_596 (I12737,I2595,I12412,I12380,);
not I_597 (I12768,I12729);
nor I_598 (I12785,I194008,I194008);
not I_599 (I12802,I12785);
nor I_600 (I12819,I12576,I12802);
nor I_601 (I12836,I12768,I12819);
DFFARX1 I_602 (I12836,I2595,I12412,I12401,);
nor I_603 (I12867,I12729,I12802);
nor I_604 (I12389,I12593,I12867);
nor I_605 (I12383,I12729,I12785);
not I_606 (I12939,I2602);
DFFARX1 I_607 (I74674,I2595,I12939,I12965,);
DFFARX1 I_608 (I12965,I2595,I12939,I12982,);
not I_609 (I12990,I12982);
nand I_610 (I13007,I74692,I74677);
and I_611 (I13024,I13007,I74680);
DFFARX1 I_612 (I13024,I2595,I12939,I13050,);
DFFARX1 I_613 (I13050,I2595,I12939,I12931,);
DFFARX1 I_614 (I13050,I2595,I12939,I12922,);
DFFARX1 I_615 (I74668,I2595,I12939,I13095,);
nand I_616 (I13103,I13095,I74671);
not I_617 (I13120,I13103);
nor I_618 (I12919,I12965,I13120);
DFFARX1 I_619 (I74683,I2595,I12939,I13160,);
not I_620 (I13168,I13160);
nor I_621 (I12925,I13168,I12990);
nand I_622 (I12913,I13168,I13103);
nand I_623 (I13213,I74689,I74686);
and I_624 (I13230,I13213,I74671);
DFFARX1 I_625 (I13230,I2595,I12939,I13256,);
nor I_626 (I13264,I13256,I12965);
DFFARX1 I_627 (I13264,I2595,I12939,I12907,);
not I_628 (I13295,I13256);
nor I_629 (I13312,I74668,I74686);
not I_630 (I13329,I13312);
nor I_631 (I13346,I13103,I13329);
nor I_632 (I13363,I13295,I13346);
DFFARX1 I_633 (I13363,I2595,I12939,I12928,);
nor I_634 (I13394,I13256,I13329);
nor I_635 (I12916,I13120,I13394);
nor I_636 (I12910,I13256,I13312);
not I_637 (I13466,I2602);
DFFARX1 I_638 (I309666,I2595,I13466,I13492,);
DFFARX1 I_639 (I13492,I2595,I13466,I13509,);
not I_640 (I13517,I13509);
nand I_641 (I13534,I309654,I309645);
and I_642 (I13551,I13534,I309642);
DFFARX1 I_643 (I13551,I2595,I13466,I13577,);
DFFARX1 I_644 (I13577,I2595,I13466,I13458,);
DFFARX1 I_645 (I13577,I2595,I13466,I13449,);
DFFARX1 I_646 (I309648,I2595,I13466,I13622,);
nand I_647 (I13630,I13622,I309660);
not I_648 (I13647,I13630);
nor I_649 (I13446,I13492,I13647);
DFFARX1 I_650 (I309657,I2595,I13466,I13687,);
not I_651 (I13695,I13687);
nor I_652 (I13452,I13695,I13517);
nand I_653 (I13440,I13695,I13630);
nand I_654 (I13740,I309651,I309645);
and I_655 (I13757,I13740,I309663);
DFFARX1 I_656 (I13757,I2595,I13466,I13783,);
nor I_657 (I13791,I13783,I13492);
DFFARX1 I_658 (I13791,I2595,I13466,I13434,);
not I_659 (I13822,I13783);
nor I_660 (I13839,I309642,I309645);
not I_661 (I13856,I13839);
nor I_662 (I13873,I13630,I13856);
nor I_663 (I13890,I13822,I13873);
DFFARX1 I_664 (I13890,I2595,I13466,I13455,);
nor I_665 (I13921,I13783,I13856);
nor I_666 (I13443,I13647,I13921);
nor I_667 (I13437,I13783,I13839);
not I_668 (I13993,I2602);
DFFARX1 I_669 (I189390,I2595,I13993,I14019,);
DFFARX1 I_670 (I14019,I2595,I13993,I14036,);
not I_671 (I14044,I14036);
nand I_672 (I14061,I189405,I189408);
and I_673 (I14078,I14061,I189387);
DFFARX1 I_674 (I14078,I2595,I13993,I14104,);
DFFARX1 I_675 (I14104,I2595,I13993,I13985,);
DFFARX1 I_676 (I14104,I2595,I13993,I13976,);
DFFARX1 I_677 (I189393,I2595,I13993,I14149,);
nand I_678 (I14157,I14149,I189399);
not I_679 (I14174,I14157);
nor I_680 (I13973,I14019,I14174);
DFFARX1 I_681 (I189387,I2595,I13993,I14214,);
not I_682 (I14222,I14214);
nor I_683 (I13979,I14222,I14044);
nand I_684 (I13967,I14222,I14157);
nand I_685 (I14267,I189402,I189384);
and I_686 (I14284,I14267,I189396);
DFFARX1 I_687 (I14284,I2595,I13993,I14310,);
nor I_688 (I14318,I14310,I14019);
DFFARX1 I_689 (I14318,I2595,I13993,I13961,);
not I_690 (I14349,I14310);
nor I_691 (I14366,I189384,I189384);
not I_692 (I14383,I14366);
nor I_693 (I14400,I14157,I14383);
nor I_694 (I14417,I14349,I14400);
DFFARX1 I_695 (I14417,I2595,I13993,I13982,);
nor I_696 (I14448,I14310,I14383);
nor I_697 (I13970,I14174,I14448);
nor I_698 (I13964,I14310,I14366);
not I_699 (I14520,I2602);
DFFARX1 I_700 (I1916,I2595,I14520,I14546,);
DFFARX1 I_701 (I14546,I2595,I14520,I14563,);
not I_702 (I14571,I14563);
nand I_703 (I14588,I1588,I1764);
and I_704 (I14605,I14588,I2188);
DFFARX1 I_705 (I14605,I2595,I14520,I14631,);
DFFARX1 I_706 (I14631,I2595,I14520,I14512,);
DFFARX1 I_707 (I14631,I2595,I14520,I14503,);
DFFARX1 I_708 (I2420,I2595,I14520,I14676,);
nand I_709 (I14684,I14676,I1812);
not I_710 (I14701,I14684);
nor I_711 (I14500,I14546,I14701);
DFFARX1 I_712 (I2564,I2595,I14520,I14741,);
not I_713 (I14749,I14741);
nor I_714 (I14506,I14749,I14571);
nand I_715 (I14494,I14749,I14684);
nand I_716 (I14794,I1708,I2484);
and I_717 (I14811,I14794,I1404);
DFFARX1 I_718 (I14811,I2595,I14520,I14837,);
nor I_719 (I14845,I14837,I14546);
DFFARX1 I_720 (I14845,I2595,I14520,I14488,);
not I_721 (I14876,I14837);
nor I_722 (I14893,I2212,I2484);
not I_723 (I14910,I14893);
nor I_724 (I14927,I14684,I14910);
nor I_725 (I14944,I14876,I14927);
DFFARX1 I_726 (I14944,I2595,I14520,I14509,);
nor I_727 (I14975,I14837,I14910);
nor I_728 (I14497,I14701,I14975);
nor I_729 (I14491,I14837,I14893);
not I_730 (I15047,I2602);
DFFARX1 I_731 (I1660,I2595,I15047,I15073,);
DFFARX1 I_732 (I15073,I2595,I15047,I15090,);
not I_733 (I15098,I15090);
nand I_734 (I15115,I1500,I2196);
and I_735 (I15132,I15115,I2252);
DFFARX1 I_736 (I15132,I2595,I15047,I15158,);
DFFARX1 I_737 (I15158,I2595,I15047,I15039,);
DFFARX1 I_738 (I15158,I2595,I15047,I15030,);
DFFARX1 I_739 (I1444,I2595,I15047,I15203,);
nand I_740 (I15211,I15203,I1428);
not I_741 (I15228,I15211);
nor I_742 (I15027,I15073,I15228);
DFFARX1 I_743 (I1612,I2595,I15047,I15268,);
not I_744 (I15276,I15268);
nor I_745 (I15033,I15276,I15098);
nand I_746 (I15021,I15276,I15211);
nand I_747 (I15321,I1844,I1876);
and I_748 (I15338,I15321,I1476);
DFFARX1 I_749 (I15338,I2595,I15047,I15364,);
nor I_750 (I15372,I15364,I15073);
DFFARX1 I_751 (I15372,I2595,I15047,I15015,);
not I_752 (I15403,I15364);
nor I_753 (I15420,I2060,I1876);
not I_754 (I15437,I15420);
nor I_755 (I15454,I15211,I15437);
nor I_756 (I15471,I15403,I15454);
DFFARX1 I_757 (I15471,I2595,I15047,I15036,);
nor I_758 (I15502,I15364,I15437);
nor I_759 (I15024,I15228,I15502);
nor I_760 (I15018,I15364,I15420);
not I_761 (I15574,I2602);
DFFARX1 I_762 (I327006,I2595,I15574,I15600,);
DFFARX1 I_763 (I15600,I2595,I15574,I15617,);
not I_764 (I15625,I15617);
nand I_765 (I15642,I326994,I326985);
and I_766 (I15659,I15642,I326982);
DFFARX1 I_767 (I15659,I2595,I15574,I15685,);
DFFARX1 I_768 (I15685,I2595,I15574,I15566,);
DFFARX1 I_769 (I15685,I2595,I15574,I15557,);
DFFARX1 I_770 (I326988,I2595,I15574,I15730,);
nand I_771 (I15738,I15730,I327000);
not I_772 (I15755,I15738);
nor I_773 (I15554,I15600,I15755);
DFFARX1 I_774 (I326997,I2595,I15574,I15795,);
not I_775 (I15803,I15795);
nor I_776 (I15560,I15803,I15625);
nand I_777 (I15548,I15803,I15738);
nand I_778 (I15848,I326991,I326985);
and I_779 (I15865,I15848,I327003);
DFFARX1 I_780 (I15865,I2595,I15574,I15891,);
nor I_781 (I15899,I15891,I15600);
DFFARX1 I_782 (I15899,I2595,I15574,I15542,);
not I_783 (I15930,I15891);
nor I_784 (I15947,I326982,I326985);
not I_785 (I15964,I15947);
nor I_786 (I15981,I15738,I15964);
nor I_787 (I15998,I15930,I15981);
DFFARX1 I_788 (I15998,I2595,I15574,I15563,);
nor I_789 (I16029,I15891,I15964);
nor I_790 (I15551,I15755,I16029);
nor I_791 (I15545,I15891,I15947);
not I_792 (I16101,I2602);
DFFARX1 I_793 (I30828,I2595,I16101,I16127,);
DFFARX1 I_794 (I16127,I2595,I16101,I16144,);
not I_795 (I16152,I16144);
nand I_796 (I16169,I30828,I30843);
and I_797 (I16186,I16169,I30846);
DFFARX1 I_798 (I16186,I2595,I16101,I16212,);
DFFARX1 I_799 (I16212,I2595,I16101,I16093,);
DFFARX1 I_800 (I16212,I2595,I16101,I16084,);
DFFARX1 I_801 (I30840,I2595,I16101,I16257,);
nand I_802 (I16265,I16257,I30849);
not I_803 (I16282,I16265);
nor I_804 (I16081,I16127,I16282);
DFFARX1 I_805 (I30825,I2595,I16101,I16322,);
not I_806 (I16330,I16322);
nor I_807 (I16087,I16330,I16152);
nand I_808 (I16075,I16330,I16265);
nand I_809 (I16375,I30825,I30831);
and I_810 (I16392,I16375,I30834);
DFFARX1 I_811 (I16392,I2595,I16101,I16418,);
nor I_812 (I16426,I16418,I16127);
DFFARX1 I_813 (I16426,I2595,I16101,I16069,);
not I_814 (I16457,I16418);
nor I_815 (I16474,I30837,I30831);
not I_816 (I16491,I16474);
nor I_817 (I16508,I16265,I16491);
nor I_818 (I16525,I16457,I16508);
DFFARX1 I_819 (I16525,I2595,I16101,I16090,);
nor I_820 (I16556,I16418,I16491);
nor I_821 (I16078,I16282,I16556);
nor I_822 (I16072,I16418,I16474);
not I_823 (I16628,I2602);
DFFARX1 I_824 (I99617,I2595,I16628,I16654,);
DFFARX1 I_825 (I16654,I2595,I16628,I16671,);
not I_826 (I16679,I16671);
nand I_827 (I16696,I99614,I99608);
and I_828 (I16713,I16696,I99602);
DFFARX1 I_829 (I16713,I2595,I16628,I16739,);
DFFARX1 I_830 (I16739,I2595,I16628,I16620,);
DFFARX1 I_831 (I16739,I2595,I16628,I16611,);
DFFARX1 I_832 (I99590,I2595,I16628,I16784,);
nand I_833 (I16792,I16784,I99599);
not I_834 (I16809,I16792);
nor I_835 (I16608,I16654,I16809);
DFFARX1 I_836 (I99596,I2595,I16628,I16849,);
not I_837 (I16857,I16849);
nor I_838 (I16614,I16857,I16679);
nand I_839 (I16602,I16857,I16792);
nand I_840 (I16902,I99593,I99611);
and I_841 (I16919,I16902,I99590);
DFFARX1 I_842 (I16919,I2595,I16628,I16945,);
nor I_843 (I16953,I16945,I16654);
DFFARX1 I_844 (I16953,I2595,I16628,I16596,);
not I_845 (I16984,I16945);
nor I_846 (I17001,I99605,I99611);
not I_847 (I17018,I17001);
nor I_848 (I17035,I16792,I17018);
nor I_849 (I17052,I16984,I17035);
DFFARX1 I_850 (I17052,I2595,I16628,I16617,);
nor I_851 (I17083,I16945,I17018);
nor I_852 (I16605,I16809,I17083);
nor I_853 (I16599,I16945,I17001);
not I_854 (I17155,I2602);
DFFARX1 I_855 (I280307,I2595,I17155,I17181,);
DFFARX1 I_856 (I17181,I2595,I17155,I17198,);
not I_857 (I17206,I17198);
nand I_858 (I17223,I280283,I280310);
and I_859 (I17240,I17223,I280295);
DFFARX1 I_860 (I17240,I2595,I17155,I17266,);
DFFARX1 I_861 (I17266,I2595,I17155,I17147,);
DFFARX1 I_862 (I17266,I2595,I17155,I17138,);
DFFARX1 I_863 (I280301,I2595,I17155,I17311,);
nand I_864 (I17319,I17311,I280286);
not I_865 (I17336,I17319);
nor I_866 (I17135,I17181,I17336);
DFFARX1 I_867 (I280304,I2595,I17155,I17376,);
not I_868 (I17384,I17376);
nor I_869 (I17141,I17384,I17206);
nand I_870 (I17129,I17384,I17319);
nand I_871 (I17429,I280289,I280292);
and I_872 (I17446,I17429,I280283);
DFFARX1 I_873 (I17446,I2595,I17155,I17472,);
nor I_874 (I17480,I17472,I17181);
DFFARX1 I_875 (I17480,I2595,I17155,I17123,);
not I_876 (I17511,I17472);
nor I_877 (I17528,I280298,I280292);
not I_878 (I17545,I17528);
nor I_879 (I17562,I17319,I17545);
nor I_880 (I17579,I17511,I17562);
DFFARX1 I_881 (I17579,I2595,I17155,I17144,);
nor I_882 (I17610,I17472,I17545);
nor I_883 (I17132,I17336,I17610);
nor I_884 (I17126,I17472,I17528);
not I_885 (I17682,I2602);
DFFARX1 I_886 (I165123,I2595,I17682,I17708,);
DFFARX1 I_887 (I17708,I2595,I17682,I17725,);
not I_888 (I17733,I17725);
nand I_889 (I17750,I165108,I165126);
and I_890 (I17767,I17750,I165120);
DFFARX1 I_891 (I17767,I2595,I17682,I17793,);
DFFARX1 I_892 (I17793,I2595,I17682,I17674,);
DFFARX1 I_893 (I17793,I2595,I17682,I17665,);
DFFARX1 I_894 (I165117,I2595,I17682,I17838,);
nand I_895 (I17846,I17838,I165108);
not I_896 (I17863,I17846);
nor I_897 (I17662,I17708,I17863);
DFFARX1 I_898 (I165111,I2595,I17682,I17903,);
not I_899 (I17911,I17903);
nor I_900 (I17668,I17911,I17733);
nand I_901 (I17656,I17911,I17846);
nand I_902 (I17956,I165132,I165114);
and I_903 (I17973,I17956,I165129);
DFFARX1 I_904 (I17973,I2595,I17682,I17999,);
nor I_905 (I18007,I17999,I17708);
DFFARX1 I_906 (I18007,I2595,I17682,I17650,);
not I_907 (I18038,I17999);
nor I_908 (I18055,I165111,I165114);
not I_909 (I18072,I18055);
nor I_910 (I18089,I17846,I18072);
nor I_911 (I18106,I18038,I18089);
DFFARX1 I_912 (I18106,I2595,I17682,I17671,);
nor I_913 (I18137,I17999,I18072);
nor I_914 (I17659,I17863,I18137);
nor I_915 (I17653,I17999,I18055);
not I_916 (I18209,I2602);
DFFARX1 I_917 (I127929,I2595,I18209,I18235,);
DFFARX1 I_918 (I18235,I2595,I18209,I18252,);
not I_919 (I18260,I18252);
nand I_920 (I18277,I127929,I127932);
and I_921 (I18294,I18277,I127953);
DFFARX1 I_922 (I18294,I2595,I18209,I18320,);
DFFARX1 I_923 (I18320,I2595,I18209,I18201,);
DFFARX1 I_924 (I18320,I2595,I18209,I18192,);
DFFARX1 I_925 (I127941,I2595,I18209,I18365,);
nand I_926 (I18373,I18365,I127944);
not I_927 (I18390,I18373);
nor I_928 (I18189,I18235,I18390);
DFFARX1 I_929 (I127950,I2595,I18209,I18430,);
not I_930 (I18438,I18430);
nor I_931 (I18195,I18438,I18260);
nand I_932 (I18183,I18438,I18373);
nand I_933 (I18483,I127947,I127935);
and I_934 (I18500,I18483,I127938);
DFFARX1 I_935 (I18500,I2595,I18209,I18526,);
nor I_936 (I18534,I18526,I18235);
DFFARX1 I_937 (I18534,I2595,I18209,I18177,);
not I_938 (I18565,I18526);
nor I_939 (I18582,I127956,I127935);
not I_940 (I18599,I18582);
nor I_941 (I18616,I18373,I18599);
nor I_942 (I18633,I18565,I18616);
DFFARX1 I_943 (I18633,I2595,I18209,I18198,);
nor I_944 (I18664,I18526,I18599);
nor I_945 (I18186,I18390,I18664);
nor I_946 (I18180,I18526,I18582);
not I_947 (I18736,I2602);
DFFARX1 I_948 (I160499,I2595,I18736,I18762,);
DFFARX1 I_949 (I18762,I2595,I18736,I18779,);
not I_950 (I18787,I18779);
nand I_951 (I18804,I160484,I160502);
and I_952 (I18821,I18804,I160496);
DFFARX1 I_953 (I18821,I2595,I18736,I18847,);
DFFARX1 I_954 (I18847,I2595,I18736,I18728,);
DFFARX1 I_955 (I18847,I2595,I18736,I18719,);
DFFARX1 I_956 (I160493,I2595,I18736,I18892,);
nand I_957 (I18900,I18892,I160484);
not I_958 (I18917,I18900);
nor I_959 (I18716,I18762,I18917);
DFFARX1 I_960 (I160487,I2595,I18736,I18957,);
not I_961 (I18965,I18957);
nor I_962 (I18722,I18965,I18787);
nand I_963 (I18710,I18965,I18900);
nand I_964 (I19010,I160508,I160490);
and I_965 (I19027,I19010,I160505);
DFFARX1 I_966 (I19027,I2595,I18736,I19053,);
nor I_967 (I19061,I19053,I18762);
DFFARX1 I_968 (I19061,I2595,I18736,I18704,);
not I_969 (I19092,I19053);
nor I_970 (I19109,I160487,I160490);
not I_971 (I19126,I19109);
nor I_972 (I19143,I18900,I19126);
nor I_973 (I19160,I19092,I19143);
DFFARX1 I_974 (I19160,I2595,I18736,I18725,);
nor I_975 (I19191,I19053,I19126);
nor I_976 (I18713,I18917,I19191);
nor I_977 (I18707,I19053,I19109);
not I_978 (I19263,I2602);
DFFARX1 I_979 (I390783,I2595,I19263,I19289,);
DFFARX1 I_980 (I19289,I2595,I19263,I19306,);
not I_981 (I19314,I19306);
nand I_982 (I19331,I390786,I390792);
and I_983 (I19348,I19331,I390801);
DFFARX1 I_984 (I19348,I2595,I19263,I19374,);
DFFARX1 I_985 (I19374,I2595,I19263,I19255,);
DFFARX1 I_986 (I19374,I2595,I19263,I19246,);
DFFARX1 I_987 (I390804,I2595,I19263,I19419,);
nand I_988 (I19427,I19419,I390795);
not I_989 (I19444,I19427);
nor I_990 (I19243,I19289,I19444);
DFFARX1 I_991 (I390783,I2595,I19263,I19484,);
not I_992 (I19492,I19484);
nor I_993 (I19249,I19492,I19314);
nand I_994 (I19237,I19492,I19427);
nand I_995 (I19537,I390810,I390789);
and I_996 (I19554,I19537,I390798);
DFFARX1 I_997 (I19554,I2595,I19263,I19580,);
nor I_998 (I19588,I19580,I19289);
DFFARX1 I_999 (I19588,I2595,I19263,I19231,);
not I_1000 (I19619,I19580);
nor I_1001 (I19636,I390807,I390789);
not I_1002 (I19653,I19636);
nor I_1003 (I19670,I19427,I19653);
nor I_1004 (I19687,I19619,I19670);
DFFARX1 I_1005 (I19687,I2595,I19263,I19252,);
nor I_1006 (I19718,I19580,I19653);
nor I_1007 (I19240,I19444,I19718);
nor I_1008 (I19234,I19580,I19636);
not I_1009 (I19790,I2602);
DFFARX1 I_1010 (I291577,I2595,I19790,I19816,);
DFFARX1 I_1011 (I19816,I2595,I19790,I19833,);
not I_1012 (I19841,I19833);
nand I_1013 (I19858,I291571,I291592);
and I_1014 (I19875,I19858,I291577);
DFFARX1 I_1015 (I19875,I2595,I19790,I19901,);
DFFARX1 I_1016 (I19901,I2595,I19790,I19782,);
DFFARX1 I_1017 (I19901,I2595,I19790,I19773,);
DFFARX1 I_1018 (I291574,I2595,I19790,I19946,);
nand I_1019 (I19954,I19946,I291583);
not I_1020 (I19971,I19954);
nor I_1021 (I19770,I19816,I19971);
DFFARX1 I_1022 (I291571,I2595,I19790,I20011,);
not I_1023 (I20019,I20011);
nor I_1024 (I19776,I20019,I19841);
nand I_1025 (I19764,I20019,I19954);
nand I_1026 (I20064,I291574,I291589);
and I_1027 (I20081,I20064,I291580);
DFFARX1 I_1028 (I20081,I2595,I19790,I20107,);
nor I_1029 (I20115,I20107,I19816);
DFFARX1 I_1030 (I20115,I2595,I19790,I19758,);
not I_1031 (I20146,I20107);
nor I_1032 (I20163,I291586,I291589);
not I_1033 (I20180,I20163);
nor I_1034 (I20197,I19954,I20180);
nor I_1035 (I20214,I20146,I20197);
DFFARX1 I_1036 (I20214,I2595,I19790,I19779,);
nor I_1037 (I20245,I20107,I20180);
nor I_1038 (I19767,I19971,I20245);
nor I_1039 (I19761,I20107,I20163);
not I_1040 (I20317,I2602);
DFFARX1 I_1041 (I359671,I2595,I20317,I20343,);
DFFARX1 I_1042 (I20343,I2595,I20317,I20360,);
not I_1043 (I20368,I20360);
nand I_1044 (I20385,I359674,I359668);
and I_1045 (I20402,I20385,I359677);
DFFARX1 I_1046 (I20402,I2595,I20317,I20428,);
DFFARX1 I_1047 (I20428,I2595,I20317,I20309,);
DFFARX1 I_1048 (I20428,I2595,I20317,I20300,);
DFFARX1 I_1049 (I359665,I2595,I20317,I20473,);
nand I_1050 (I20481,I20473,I359680);
not I_1051 (I20498,I20481);
nor I_1052 (I20297,I20343,I20498);
DFFARX1 I_1053 (I359656,I2595,I20317,I20538,);
not I_1054 (I20546,I20538);
nor I_1055 (I20303,I20546,I20368);
nand I_1056 (I20291,I20546,I20481);
nand I_1057 (I20591,I359659,I359659);
and I_1058 (I20608,I20591,I359656);
DFFARX1 I_1059 (I20608,I2595,I20317,I20634,);
nor I_1060 (I20642,I20634,I20343);
DFFARX1 I_1061 (I20642,I2595,I20317,I20285,);
not I_1062 (I20673,I20634);
nor I_1063 (I20690,I359662,I359659);
not I_1064 (I20707,I20690);
nor I_1065 (I20724,I20481,I20707);
nor I_1066 (I20741,I20673,I20724);
DFFARX1 I_1067 (I20741,I2595,I20317,I20306,);
nor I_1068 (I20772,I20634,I20707);
nor I_1069 (I20294,I20498,I20772);
nor I_1070 (I20288,I20634,I20690);
not I_1071 (I20844,I2602);
DFFARX1 I_1072 (I288059,I2595,I20844,I20870,);
DFFARX1 I_1073 (I20870,I2595,I20844,I20887,);
not I_1074 (I20895,I20887);
nand I_1075 (I20912,I288035,I288062);
and I_1076 (I20929,I20912,I288047);
DFFARX1 I_1077 (I20929,I2595,I20844,I20955,);
DFFARX1 I_1078 (I20955,I2595,I20844,I20836,);
DFFARX1 I_1079 (I20955,I2595,I20844,I20827,);
DFFARX1 I_1080 (I288053,I2595,I20844,I21000,);
nand I_1081 (I21008,I21000,I288038);
not I_1082 (I21025,I21008);
nor I_1083 (I20824,I20870,I21025);
DFFARX1 I_1084 (I288056,I2595,I20844,I21065,);
not I_1085 (I21073,I21065);
nor I_1086 (I20830,I21073,I20895);
nand I_1087 (I20818,I21073,I21008);
nand I_1088 (I21118,I288041,I288044);
and I_1089 (I21135,I21118,I288035);
DFFARX1 I_1090 (I21135,I2595,I20844,I21161,);
nor I_1091 (I21169,I21161,I20870);
DFFARX1 I_1092 (I21169,I2595,I20844,I20812,);
not I_1093 (I21200,I21161);
nor I_1094 (I21217,I288050,I288044);
not I_1095 (I21234,I21217);
nor I_1096 (I21251,I21008,I21234);
nor I_1097 (I21268,I21200,I21251);
DFFARX1 I_1098 (I21268,I2595,I20844,I20833,);
nor I_1099 (I21299,I21161,I21234);
nor I_1100 (I20821,I21025,I21299);
nor I_1101 (I20815,I21161,I21217);
not I_1102 (I21371,I2602);
DFFARX1 I_1103 (I35044,I2595,I21371,I21397,);
DFFARX1 I_1104 (I21397,I2595,I21371,I21414,);
not I_1105 (I21422,I21414);
nand I_1106 (I21439,I35044,I35059);
and I_1107 (I21456,I21439,I35062);
DFFARX1 I_1108 (I21456,I2595,I21371,I21482,);
DFFARX1 I_1109 (I21482,I2595,I21371,I21363,);
DFFARX1 I_1110 (I21482,I2595,I21371,I21354,);
DFFARX1 I_1111 (I35056,I2595,I21371,I21527,);
nand I_1112 (I21535,I21527,I35065);
not I_1113 (I21552,I21535);
nor I_1114 (I21351,I21397,I21552);
DFFARX1 I_1115 (I35041,I2595,I21371,I21592,);
not I_1116 (I21600,I21592);
nor I_1117 (I21357,I21600,I21422);
nand I_1118 (I21345,I21600,I21535);
nand I_1119 (I21645,I35041,I35047);
and I_1120 (I21662,I21645,I35050);
DFFARX1 I_1121 (I21662,I2595,I21371,I21688,);
nor I_1122 (I21696,I21688,I21397);
DFFARX1 I_1123 (I21696,I2595,I21371,I21339,);
not I_1124 (I21727,I21688);
nor I_1125 (I21744,I35053,I35047);
not I_1126 (I21761,I21744);
nor I_1127 (I21778,I21535,I21761);
nor I_1128 (I21795,I21727,I21778);
DFFARX1 I_1129 (I21795,I2595,I21371,I21360,);
nor I_1130 (I21826,I21688,I21761);
nor I_1131 (I21348,I21552,I21826);
nor I_1132 (I21342,I21688,I21744);
not I_1133 (I21898,I2602);
DFFARX1 I_1134 (I108576,I2595,I21898,I21924,);
DFFARX1 I_1135 (I21924,I2595,I21898,I21941,);
not I_1136 (I21949,I21941);
nand I_1137 (I21966,I108573,I108567);
and I_1138 (I21983,I21966,I108561);
DFFARX1 I_1139 (I21983,I2595,I21898,I22009,);
DFFARX1 I_1140 (I22009,I2595,I21898,I21890,);
DFFARX1 I_1141 (I22009,I2595,I21898,I21881,);
DFFARX1 I_1142 (I108549,I2595,I21898,I22054,);
nand I_1143 (I22062,I22054,I108558);
not I_1144 (I22079,I22062);
nor I_1145 (I21878,I21924,I22079);
DFFARX1 I_1146 (I108555,I2595,I21898,I22119,);
not I_1147 (I22127,I22119);
nor I_1148 (I21884,I22127,I21949);
nand I_1149 (I21872,I22127,I22062);
nand I_1150 (I22172,I108552,I108570);
and I_1151 (I22189,I22172,I108549);
DFFARX1 I_1152 (I22189,I2595,I21898,I22215,);
nor I_1153 (I22223,I22215,I21924);
DFFARX1 I_1154 (I22223,I2595,I21898,I21866,);
not I_1155 (I22254,I22215);
nor I_1156 (I22271,I108564,I108570);
not I_1157 (I22288,I22271);
nor I_1158 (I22305,I22062,I22288);
nor I_1159 (I22322,I22254,I22305);
DFFARX1 I_1160 (I22322,I2595,I21898,I21887,);
nor I_1161 (I22353,I22215,I22288);
nor I_1162 (I21875,I22079,I22353);
nor I_1163 (I21869,I22215,I22271);
not I_1164 (I22425,I2602);
DFFARX1 I_1165 (I293260,I2595,I22425,I22451,);
DFFARX1 I_1166 (I22451,I2595,I22425,I22468,);
not I_1167 (I22476,I22468);
nand I_1168 (I22493,I293254,I293275);
and I_1169 (I22510,I22493,I293260);
DFFARX1 I_1170 (I22510,I2595,I22425,I22536,);
DFFARX1 I_1171 (I22536,I2595,I22425,I22417,);
DFFARX1 I_1172 (I22536,I2595,I22425,I22408,);
DFFARX1 I_1173 (I293257,I2595,I22425,I22581,);
nand I_1174 (I22589,I22581,I293266);
not I_1175 (I22606,I22589);
nor I_1176 (I22405,I22451,I22606);
DFFARX1 I_1177 (I293254,I2595,I22425,I22646,);
not I_1178 (I22654,I22646);
nor I_1179 (I22411,I22654,I22476);
nand I_1180 (I22399,I22654,I22589);
nand I_1181 (I22699,I293257,I293272);
and I_1182 (I22716,I22699,I293263);
DFFARX1 I_1183 (I22716,I2595,I22425,I22742,);
nor I_1184 (I22750,I22742,I22451);
DFFARX1 I_1185 (I22750,I2595,I22425,I22393,);
not I_1186 (I22781,I22742);
nor I_1187 (I22798,I293269,I293272);
not I_1188 (I22815,I22798);
nor I_1189 (I22832,I22589,I22815);
nor I_1190 (I22849,I22781,I22832);
DFFARX1 I_1191 (I22849,I2595,I22425,I22414,);
nor I_1192 (I22880,I22742,I22815);
nor I_1193 (I22402,I22606,I22880);
nor I_1194 (I22396,I22742,I22798);
not I_1195 (I22952,I2602);
DFFARX1 I_1196 (I368928,I2595,I22952,I22978,);
DFFARX1 I_1197 (I22978,I2595,I22952,I22995,);
not I_1198 (I23003,I22995);
nand I_1199 (I23020,I368919,I368925);
and I_1200 (I23037,I23020,I368904);
DFFARX1 I_1201 (I23037,I2595,I22952,I23063,);
DFFARX1 I_1202 (I23063,I2595,I22952,I22944,);
DFFARX1 I_1203 (I23063,I2595,I22952,I22935,);
DFFARX1 I_1204 (I368922,I2595,I22952,I23108,);
nand I_1205 (I23116,I23108,I368904);
not I_1206 (I23133,I23116);
nor I_1207 (I22932,I22978,I23133);
DFFARX1 I_1208 (I368916,I2595,I22952,I23173,);
not I_1209 (I23181,I23173);
nor I_1210 (I22938,I23181,I23003);
nand I_1211 (I22926,I23181,I23116);
nand I_1212 (I23226,I368910,I368931);
and I_1213 (I23243,I23226,I368913);
DFFARX1 I_1214 (I23243,I2595,I22952,I23269,);
nor I_1215 (I23277,I23269,I22978);
DFFARX1 I_1216 (I23277,I2595,I22952,I22920,);
not I_1217 (I23308,I23269);
nor I_1218 (I23325,I368907,I368931);
not I_1219 (I23342,I23325);
nor I_1220 (I23359,I23116,I23342);
nor I_1221 (I23376,I23308,I23359);
DFFARX1 I_1222 (I23376,I2595,I22952,I22941,);
nor I_1223 (I23407,I23269,I23342);
nor I_1224 (I22929,I23133,I23407);
nor I_1225 (I22923,I23269,I23325);
not I_1226 (I23479,I2602);
DFFARX1 I_1227 (I138827,I2595,I23479,I23505,);
not I_1228 (I23513,I23505);
nand I_1229 (I23530,I138821,I138812);
and I_1230 (I23547,I23530,I138833);
DFFARX1 I_1231 (I23547,I2595,I23479,I23573,);
DFFARX1 I_1232 (I138815,I2595,I23479,I23590,);
and I_1233 (I23598,I23590,I138809);
nor I_1234 (I23615,I23573,I23598);
DFFARX1 I_1235 (I23615,I2595,I23479,I23447,);
nand I_1236 (I23646,I23590,I138809);
nand I_1237 (I23663,I23513,I23646);
not I_1238 (I23459,I23663);
DFFARX1 I_1239 (I138809,I2595,I23479,I23703,);
DFFARX1 I_1240 (I23703,I2595,I23479,I23468,);
nand I_1241 (I23725,I138836,I138818);
and I_1242 (I23742,I23725,I138824);
DFFARX1 I_1243 (I23742,I2595,I23479,I23768,);
DFFARX1 I_1244 (I23768,I2595,I23479,I23785,);
not I_1245 (I23471,I23785);
not I_1246 (I23807,I23768);
nand I_1247 (I23456,I23807,I23646);
nor I_1248 (I23838,I138830,I138818);
not I_1249 (I23855,I23838);
nor I_1250 (I23872,I23807,I23855);
nor I_1251 (I23889,I23513,I23872);
DFFARX1 I_1252 (I23889,I2595,I23479,I23465,);
nor I_1253 (I23920,I23573,I23855);
nor I_1254 (I23453,I23768,I23920);
nor I_1255 (I23462,I23703,I23838);
nor I_1256 (I23450,I23573,I23838);
not I_1257 (I24006,I2602);
DFFARX1 I_1258 (I273832,I2595,I24006,I24032,);
not I_1259 (I24040,I24032);
nand I_1260 (I24057,I273850,I273844);
and I_1261 (I24074,I24057,I273823);
DFFARX1 I_1262 (I24074,I2595,I24006,I24100,);
DFFARX1 I_1263 (I273841,I2595,I24006,I24117,);
and I_1264 (I24125,I24117,I273826);
nor I_1265 (I24142,I24100,I24125);
DFFARX1 I_1266 (I24142,I2595,I24006,I23974,);
nand I_1267 (I24173,I24117,I273826);
nand I_1268 (I24190,I24040,I24173);
not I_1269 (I23986,I24190);
DFFARX1 I_1270 (I273838,I2595,I24006,I24230,);
DFFARX1 I_1271 (I24230,I2595,I24006,I23995,);
nand I_1272 (I24252,I273847,I273835);
and I_1273 (I24269,I24252,I273829);
DFFARX1 I_1274 (I24269,I2595,I24006,I24295,);
DFFARX1 I_1275 (I24295,I2595,I24006,I24312,);
not I_1276 (I23998,I24312);
not I_1277 (I24334,I24295);
nand I_1278 (I23983,I24334,I24173);
nor I_1279 (I24365,I273823,I273835);
not I_1280 (I24382,I24365);
nor I_1281 (I24399,I24334,I24382);
nor I_1282 (I24416,I24040,I24399);
DFFARX1 I_1283 (I24416,I2595,I24006,I23992,);
nor I_1284 (I24447,I24100,I24382);
nor I_1285 (I23980,I24295,I24447);
nor I_1286 (I23989,I24230,I24365);
nor I_1287 (I23977,I24100,I24365);
not I_1288 (I24533,I2602);
DFFARX1 I_1289 (I178411,I2595,I24533,I24559,);
not I_1290 (I24567,I24559);
nand I_1291 (I24584,I178423,I178408);
and I_1292 (I24601,I24584,I178402);
DFFARX1 I_1293 (I24601,I2595,I24533,I24627,);
DFFARX1 I_1294 (I178417,I2595,I24533,I24644,);
and I_1295 (I24652,I24644,I178405);
nor I_1296 (I24669,I24627,I24652);
DFFARX1 I_1297 (I24669,I2595,I24533,I24501,);
nand I_1298 (I24700,I24644,I178405);
nand I_1299 (I24717,I24567,I24700);
not I_1300 (I24513,I24717);
DFFARX1 I_1301 (I178414,I2595,I24533,I24757,);
DFFARX1 I_1302 (I24757,I2595,I24533,I24522,);
nand I_1303 (I24779,I178420,I178426);
and I_1304 (I24796,I24779,I178402);
DFFARX1 I_1305 (I24796,I2595,I24533,I24822,);
DFFARX1 I_1306 (I24822,I2595,I24533,I24839,);
not I_1307 (I24525,I24839);
not I_1308 (I24861,I24822);
nand I_1309 (I24510,I24861,I24700);
nor I_1310 (I24892,I178405,I178426);
not I_1311 (I24909,I24892);
nor I_1312 (I24926,I24861,I24909);
nor I_1313 (I24943,I24567,I24926);
DFFARX1 I_1314 (I24943,I2595,I24533,I24519,);
nor I_1315 (I24974,I24627,I24909);
nor I_1316 (I24507,I24822,I24974);
nor I_1317 (I24516,I24757,I24892);
nor I_1318 (I24504,I24627,I24892);
not I_1319 (I25060,I2602);
DFFARX1 I_1320 (I113319,I2595,I25060,I25086,);
not I_1321 (I25094,I25086);
nand I_1322 (I25111,I113301,I113316);
and I_1323 (I25128,I25111,I113292);
DFFARX1 I_1324 (I25128,I2595,I25060,I25154,);
DFFARX1 I_1325 (I113295,I2595,I25060,I25171,);
and I_1326 (I25179,I25171,I113310);
nor I_1327 (I25196,I25154,I25179);
DFFARX1 I_1328 (I25196,I2595,I25060,I25028,);
nand I_1329 (I25227,I25171,I113310);
nand I_1330 (I25244,I25094,I25227);
not I_1331 (I25040,I25244);
DFFARX1 I_1332 (I113313,I2595,I25060,I25284,);
DFFARX1 I_1333 (I25284,I2595,I25060,I25049,);
nand I_1334 (I25306,I113292,I113304);
and I_1335 (I25323,I25306,I113298);
DFFARX1 I_1336 (I25323,I2595,I25060,I25349,);
DFFARX1 I_1337 (I25349,I2595,I25060,I25366,);
not I_1338 (I25052,I25366);
not I_1339 (I25388,I25349);
nand I_1340 (I25037,I25388,I25227);
nor I_1341 (I25419,I113307,I113304);
not I_1342 (I25436,I25419);
nor I_1343 (I25453,I25388,I25436);
nor I_1344 (I25470,I25094,I25453);
DFFARX1 I_1345 (I25470,I2595,I25060,I25046,);
nor I_1346 (I25501,I25154,I25436);
nor I_1347 (I25034,I25349,I25501);
nor I_1348 (I25043,I25284,I25419);
nor I_1349 (I25031,I25154,I25419);
not I_1350 (I25587,I2602);
DFFARX1 I_1351 (I99090,I2595,I25587,I25613,);
not I_1352 (I25621,I25613);
nand I_1353 (I25638,I99072,I99087);
and I_1354 (I25655,I25638,I99063);
DFFARX1 I_1355 (I25655,I2595,I25587,I25681,);
DFFARX1 I_1356 (I99066,I2595,I25587,I25698,);
and I_1357 (I25706,I25698,I99081);
nor I_1358 (I25723,I25681,I25706);
DFFARX1 I_1359 (I25723,I2595,I25587,I25555,);
nand I_1360 (I25754,I25698,I99081);
nand I_1361 (I25771,I25621,I25754);
not I_1362 (I25567,I25771);
DFFARX1 I_1363 (I99084,I2595,I25587,I25811,);
DFFARX1 I_1364 (I25811,I2595,I25587,I25576,);
nand I_1365 (I25833,I99063,I99075);
and I_1366 (I25850,I25833,I99069);
DFFARX1 I_1367 (I25850,I2595,I25587,I25876,);
DFFARX1 I_1368 (I25876,I2595,I25587,I25893,);
not I_1369 (I25579,I25893);
not I_1370 (I25915,I25876);
nand I_1371 (I25564,I25915,I25754);
nor I_1372 (I25946,I99078,I99075);
not I_1373 (I25963,I25946);
nor I_1374 (I25980,I25915,I25963);
nor I_1375 (I25997,I25621,I25980);
DFFARX1 I_1376 (I25997,I2595,I25587,I25573,);
nor I_1377 (I26028,I25681,I25963);
nor I_1378 (I25561,I25876,I26028);
nor I_1379 (I25570,I25811,I25946);
nor I_1380 (I25558,I25681,I25946);
not I_1381 (I26114,I2602);
DFFARX1 I_1382 (I56830,I2595,I26114,I26140,);
not I_1383 (I26148,I26140);
nand I_1384 (I26165,I56824,I56818);
and I_1385 (I26182,I26165,I56839);
DFFARX1 I_1386 (I26182,I2595,I26114,I26208,);
DFFARX1 I_1387 (I56836,I2595,I26114,I26225,);
and I_1388 (I26233,I26225,I56833);
nor I_1389 (I26250,I26208,I26233);
DFFARX1 I_1390 (I26250,I2595,I26114,I26082,);
nand I_1391 (I26281,I26225,I56833);
nand I_1392 (I26298,I26148,I26281);
not I_1393 (I26094,I26298);
DFFARX1 I_1394 (I56818,I2595,I26114,I26338,);
DFFARX1 I_1395 (I26338,I2595,I26114,I26103,);
nand I_1396 (I26360,I56821,I56821);
and I_1397 (I26377,I26360,I56842);
DFFARX1 I_1398 (I26377,I2595,I26114,I26403,);
DFFARX1 I_1399 (I26403,I2595,I26114,I26420,);
not I_1400 (I26106,I26420);
not I_1401 (I26442,I26403);
nand I_1402 (I26091,I26442,I26281);
nor I_1403 (I26473,I56827,I56821);
not I_1404 (I26490,I26473);
nor I_1405 (I26507,I26442,I26490);
nor I_1406 (I26524,I26148,I26507);
DFFARX1 I_1407 (I26524,I2595,I26114,I26100,);
nor I_1408 (I26555,I26208,I26490);
nor I_1409 (I26088,I26403,I26555);
nor I_1410 (I26097,I26338,I26473);
nor I_1411 (I26085,I26208,I26473);
not I_1412 (I26641,I2602);
DFFARX1 I_1413 (I83807,I2595,I26641,I26667,);
not I_1414 (I26675,I26667);
nand I_1415 (I26692,I83789,I83804);
and I_1416 (I26709,I26692,I83780);
DFFARX1 I_1417 (I26709,I2595,I26641,I26735,);
DFFARX1 I_1418 (I83783,I2595,I26641,I26752,);
and I_1419 (I26760,I26752,I83798);
nor I_1420 (I26777,I26735,I26760);
DFFARX1 I_1421 (I26777,I2595,I26641,I26609,);
nand I_1422 (I26808,I26752,I83798);
nand I_1423 (I26825,I26675,I26808);
not I_1424 (I26621,I26825);
DFFARX1 I_1425 (I83801,I2595,I26641,I26865,);
DFFARX1 I_1426 (I26865,I2595,I26641,I26630,);
nand I_1427 (I26887,I83780,I83792);
and I_1428 (I26904,I26887,I83786);
DFFARX1 I_1429 (I26904,I2595,I26641,I26930,);
DFFARX1 I_1430 (I26930,I2595,I26641,I26947,);
not I_1431 (I26633,I26947);
not I_1432 (I26969,I26930);
nand I_1433 (I26618,I26969,I26808);
nor I_1434 (I27000,I83795,I83792);
not I_1435 (I27017,I27000);
nor I_1436 (I27034,I26969,I27017);
nor I_1437 (I27051,I26675,I27034);
DFFARX1 I_1438 (I27051,I2595,I26641,I26627,);
nor I_1439 (I27082,I26735,I27017);
nor I_1440 (I26615,I26930,I27082);
nor I_1441 (I26624,I26865,I27000);
nor I_1442 (I26612,I26735,I27000);
not I_1443 (I27168,I2602);
DFFARX1 I_1444 (I222342,I2595,I27168,I27194,);
not I_1445 (I27202,I27194);
nand I_1446 (I27219,I222333,I222351);
and I_1447 (I27236,I27219,I222330);
DFFARX1 I_1448 (I27236,I2595,I27168,I27262,);
DFFARX1 I_1449 (I222333,I2595,I27168,I27279,);
and I_1450 (I27287,I27279,I222336);
nor I_1451 (I27304,I27262,I27287);
DFFARX1 I_1452 (I27304,I2595,I27168,I27136,);
nand I_1453 (I27335,I27279,I222336);
nand I_1454 (I27352,I27202,I27335);
not I_1455 (I27148,I27352);
DFFARX1 I_1456 (I222330,I2595,I27168,I27392,);
DFFARX1 I_1457 (I27392,I2595,I27168,I27157,);
nand I_1458 (I27414,I222348,I222339);
and I_1459 (I27431,I27414,I222354);
DFFARX1 I_1460 (I27431,I2595,I27168,I27457,);
DFFARX1 I_1461 (I27457,I2595,I27168,I27474,);
not I_1462 (I27160,I27474);
not I_1463 (I27496,I27457);
nand I_1464 (I27145,I27496,I27335);
nor I_1465 (I27527,I222345,I222339);
not I_1466 (I27544,I27527);
nor I_1467 (I27561,I27496,I27544);
nor I_1468 (I27578,I27202,I27561);
DFFARX1 I_1469 (I27578,I2595,I27168,I27154,);
nor I_1470 (I27609,I27262,I27544);
nor I_1471 (I27142,I27457,I27609);
nor I_1472 (I27151,I27392,I27527);
nor I_1473 (I27139,I27262,I27527);
not I_1474 (I27695,I2602);
DFFARX1 I_1475 (I49690,I2595,I27695,I27721,);
not I_1476 (I27729,I27721);
nand I_1477 (I27746,I49684,I49678);
and I_1478 (I27763,I27746,I49699);
DFFARX1 I_1479 (I27763,I2595,I27695,I27789,);
DFFARX1 I_1480 (I49696,I2595,I27695,I27806,);
and I_1481 (I27814,I27806,I49693);
nor I_1482 (I27831,I27789,I27814);
DFFARX1 I_1483 (I27831,I2595,I27695,I27663,);
nand I_1484 (I27862,I27806,I49693);
nand I_1485 (I27879,I27729,I27862);
not I_1486 (I27675,I27879);
DFFARX1 I_1487 (I49678,I2595,I27695,I27919,);
DFFARX1 I_1488 (I27919,I2595,I27695,I27684,);
nand I_1489 (I27941,I49681,I49681);
and I_1490 (I27958,I27941,I49702);
DFFARX1 I_1491 (I27958,I2595,I27695,I27984,);
DFFARX1 I_1492 (I27984,I2595,I27695,I28001,);
not I_1493 (I27687,I28001);
not I_1494 (I28023,I27984);
nand I_1495 (I27672,I28023,I27862);
nor I_1496 (I28054,I49687,I49681);
not I_1497 (I28071,I28054);
nor I_1498 (I28088,I28023,I28071);
nor I_1499 (I28105,I27729,I28088);
DFFARX1 I_1500 (I28105,I2595,I27695,I27681,);
nor I_1501 (I28136,I27789,I28071);
nor I_1502 (I27669,I27984,I28136);
nor I_1503 (I27678,I27919,I28054);
nor I_1504 (I27666,I27789,I28054);
not I_1505 (I28222,I2602);
DFFARX1 I_1506 (I385440,I2595,I28222,I28248,);
not I_1507 (I28256,I28248);
nand I_1508 (I28273,I385434,I385455);
and I_1509 (I28290,I28273,I385431);
DFFARX1 I_1510 (I28290,I2595,I28222,I28316,);
DFFARX1 I_1511 (I385452,I2595,I28222,I28333,);
and I_1512 (I28341,I28333,I385449);
nor I_1513 (I28358,I28316,I28341);
DFFARX1 I_1514 (I28358,I2595,I28222,I28190,);
nand I_1515 (I28389,I28333,I385449);
nand I_1516 (I28406,I28256,I28389);
not I_1517 (I28202,I28406);
DFFARX1 I_1518 (I385437,I2595,I28222,I28446,);
DFFARX1 I_1519 (I28446,I2595,I28222,I28211,);
nand I_1520 (I28468,I385446,I385443);
and I_1521 (I28485,I28468,I385428);
DFFARX1 I_1522 (I28485,I2595,I28222,I28511,);
DFFARX1 I_1523 (I28511,I2595,I28222,I28528,);
not I_1524 (I28214,I28528);
not I_1525 (I28550,I28511);
nand I_1526 (I28199,I28550,I28389);
nor I_1527 (I28581,I385428,I385443);
not I_1528 (I28598,I28581);
nor I_1529 (I28615,I28550,I28598);
nor I_1530 (I28632,I28256,I28615);
DFFARX1 I_1531 (I28632,I2595,I28222,I28208,);
nor I_1532 (I28663,I28316,I28598);
nor I_1533 (I28196,I28511,I28663);
nor I_1534 (I28205,I28446,I28581);
nor I_1535 (I28193,I28316,I28581);
not I_1536 (I28749,I2602);
DFFARX1 I_1537 (I199222,I2595,I28749,I28775,);
not I_1538 (I28783,I28775);
nand I_1539 (I28800,I199213,I199231);
and I_1540 (I28817,I28800,I199210);
DFFARX1 I_1541 (I28817,I2595,I28749,I28843,);
DFFARX1 I_1542 (I199213,I2595,I28749,I28860,);
and I_1543 (I28868,I28860,I199216);
nor I_1544 (I28885,I28843,I28868);
DFFARX1 I_1545 (I28885,I2595,I28749,I28717,);
nand I_1546 (I28916,I28860,I199216);
nand I_1547 (I28933,I28783,I28916);
not I_1548 (I28729,I28933);
DFFARX1 I_1549 (I199210,I2595,I28749,I28973,);
DFFARX1 I_1550 (I28973,I2595,I28749,I28738,);
nand I_1551 (I28995,I199228,I199219);
and I_1552 (I29012,I28995,I199234);
DFFARX1 I_1553 (I29012,I2595,I28749,I29038,);
DFFARX1 I_1554 (I29038,I2595,I28749,I29055,);
not I_1555 (I28741,I29055);
not I_1556 (I29077,I29038);
nand I_1557 (I28726,I29077,I28916);
nor I_1558 (I29108,I199225,I199219);
not I_1559 (I29125,I29108);
nor I_1560 (I29142,I29077,I29125);
nor I_1561 (I29159,I28783,I29142);
DFFARX1 I_1562 (I29159,I2595,I28749,I28735,);
nor I_1563 (I29190,I28843,I29125);
nor I_1564 (I28723,I29038,I29190);
nor I_1565 (I28732,I28973,I29108);
nor I_1566 (I28720,I28843,I29108);
not I_1567 (I29276,I2602);
DFFARX1 I_1568 (I276416,I2595,I29276,I29302,);
not I_1569 (I29310,I29302);
nand I_1570 (I29327,I276434,I276428);
and I_1571 (I29344,I29327,I276407);
DFFARX1 I_1572 (I29344,I2595,I29276,I29370,);
DFFARX1 I_1573 (I276425,I2595,I29276,I29387,);
and I_1574 (I29395,I29387,I276410);
nor I_1575 (I29412,I29370,I29395);
DFFARX1 I_1576 (I29412,I2595,I29276,I29244,);
nand I_1577 (I29443,I29387,I276410);
nand I_1578 (I29460,I29310,I29443);
not I_1579 (I29256,I29460);
DFFARX1 I_1580 (I276422,I2595,I29276,I29500,);
DFFARX1 I_1581 (I29500,I2595,I29276,I29265,);
nand I_1582 (I29522,I276431,I276419);
and I_1583 (I29539,I29522,I276413);
DFFARX1 I_1584 (I29539,I2595,I29276,I29565,);
DFFARX1 I_1585 (I29565,I2595,I29276,I29582,);
not I_1586 (I29268,I29582);
not I_1587 (I29604,I29565);
nand I_1588 (I29253,I29604,I29443);
nor I_1589 (I29635,I276407,I276419);
not I_1590 (I29652,I29635);
nor I_1591 (I29669,I29604,I29652);
nor I_1592 (I29686,I29310,I29669);
DFFARX1 I_1593 (I29686,I2595,I29276,I29262,);
nor I_1594 (I29717,I29370,I29652);
nor I_1595 (I29250,I29565,I29717);
nor I_1596 (I29259,I29500,I29635);
nor I_1597 (I29247,I29370,I29635);
not I_1598 (I29803,I2602);
DFFARX1 I_1599 (I60400,I2595,I29803,I29829,);
not I_1600 (I29837,I29829);
nand I_1601 (I29854,I60394,I60388);
and I_1602 (I29871,I29854,I60409);
DFFARX1 I_1603 (I29871,I2595,I29803,I29897,);
DFFARX1 I_1604 (I60406,I2595,I29803,I29914,);
and I_1605 (I29922,I29914,I60403);
nor I_1606 (I29939,I29897,I29922);
DFFARX1 I_1607 (I29939,I2595,I29803,I29771,);
nand I_1608 (I29970,I29914,I60403);
nand I_1609 (I29987,I29837,I29970);
not I_1610 (I29783,I29987);
DFFARX1 I_1611 (I60388,I2595,I29803,I30027,);
DFFARX1 I_1612 (I30027,I2595,I29803,I29792,);
nand I_1613 (I30049,I60391,I60391);
and I_1614 (I30066,I30049,I60412);
DFFARX1 I_1615 (I30066,I2595,I29803,I30092,);
DFFARX1 I_1616 (I30092,I2595,I29803,I30109,);
not I_1617 (I29795,I30109);
not I_1618 (I30131,I30092);
nand I_1619 (I29780,I30131,I29970);
nor I_1620 (I30162,I60397,I60391);
not I_1621 (I30179,I30162);
nor I_1622 (I30196,I30131,I30179);
nor I_1623 (I30213,I29837,I30196);
DFFARX1 I_1624 (I30213,I2595,I29803,I29789,);
nor I_1625 (I30244,I29897,I30179);
nor I_1626 (I29777,I30092,I30244);
nor I_1627 (I29786,I30027,I30162);
nor I_1628 (I29774,I29897,I30162);
not I_1629 (I30330,I2602);
DFFARX1 I_1630 (I299989,I2595,I30330,I30356,);
not I_1631 (I30364,I30356);
nand I_1632 (I30381,I299986,I299992);
and I_1633 (I30398,I30381,I299989);
DFFARX1 I_1634 (I30398,I2595,I30330,I30424,);
DFFARX1 I_1635 (I299992,I2595,I30330,I30441,);
and I_1636 (I30449,I30441,I299986);
nor I_1637 (I30466,I30424,I30449);
DFFARX1 I_1638 (I30466,I2595,I30330,I30298,);
nand I_1639 (I30497,I30441,I299986);
nand I_1640 (I30514,I30364,I30497);
not I_1641 (I30310,I30514);
DFFARX1 I_1642 (I299995,I2595,I30330,I30554,);
DFFARX1 I_1643 (I30554,I2595,I30330,I30319,);
nand I_1644 (I30576,I299998,I300007);
and I_1645 (I30593,I30576,I300001);
DFFARX1 I_1646 (I30593,I2595,I30330,I30619,);
DFFARX1 I_1647 (I30619,I2595,I30330,I30636,);
not I_1648 (I30322,I30636);
not I_1649 (I30658,I30619);
nand I_1650 (I30307,I30658,I30497);
nor I_1651 (I30689,I300004,I300007);
not I_1652 (I30706,I30689);
nor I_1653 (I30723,I30658,I30706);
nor I_1654 (I30740,I30364,I30723);
DFFARX1 I_1655 (I30740,I2595,I30330,I30316,);
nor I_1656 (I30771,I30424,I30706);
nor I_1657 (I30304,I30619,I30771);
nor I_1658 (I30313,I30554,I30689);
nor I_1659 (I30301,I30424,I30689);
not I_1660 (I30857,I2602);
DFFARX1 I_1661 (I326410,I2595,I30857,I30883,);
not I_1662 (I30891,I30883);
nand I_1663 (I30908,I326425,I326404);
and I_1664 (I30925,I30908,I326407);
DFFARX1 I_1665 (I30925,I2595,I30857,I30951,);
DFFARX1 I_1666 (I326428,I2595,I30857,I30968,);
and I_1667 (I30976,I30968,I326407);
nor I_1668 (I30993,I30951,I30976);
DFFARX1 I_1669 (I30993,I2595,I30857,I30825,);
nand I_1670 (I31024,I30968,I326407);
nand I_1671 (I31041,I30891,I31024);
not I_1672 (I30837,I31041);
DFFARX1 I_1673 (I326404,I2595,I30857,I31081,);
DFFARX1 I_1674 (I31081,I2595,I30857,I30846,);
nand I_1675 (I31103,I326416,I326413);
and I_1676 (I31120,I31103,I326419);
DFFARX1 I_1677 (I31120,I2595,I30857,I31146,);
DFFARX1 I_1678 (I31146,I2595,I30857,I31163,);
not I_1679 (I30849,I31163);
not I_1680 (I31185,I31146);
nand I_1681 (I30834,I31185,I31024);
nor I_1682 (I31216,I326422,I326413);
not I_1683 (I31233,I31216);
nor I_1684 (I31250,I31185,I31233);
nor I_1685 (I31267,I30891,I31250);
DFFARX1 I_1686 (I31267,I2595,I30857,I30843,);
nor I_1687 (I31298,I30951,I31233);
nor I_1688 (I30831,I31146,I31298);
nor I_1689 (I30840,I31081,I31216);
nor I_1690 (I30828,I30951,I31216);
not I_1691 (I31384,I2602);
DFFARX1 I_1692 (I131211,I2595,I31384,I31410,);
not I_1693 (I31418,I31410);
nand I_1694 (I31435,I131205,I131196);
and I_1695 (I31452,I31435,I131217);
DFFARX1 I_1696 (I31452,I2595,I31384,I31478,);
DFFARX1 I_1697 (I131199,I2595,I31384,I31495,);
and I_1698 (I31503,I31495,I131193);
nor I_1699 (I31520,I31478,I31503);
DFFARX1 I_1700 (I31520,I2595,I31384,I31352,);
nand I_1701 (I31551,I31495,I131193);
nand I_1702 (I31568,I31418,I31551);
not I_1703 (I31364,I31568);
DFFARX1 I_1704 (I131193,I2595,I31384,I31608,);
DFFARX1 I_1705 (I31608,I2595,I31384,I31373,);
nand I_1706 (I31630,I131220,I131202);
and I_1707 (I31647,I31630,I131208);
DFFARX1 I_1708 (I31647,I2595,I31384,I31673,);
DFFARX1 I_1709 (I31673,I2595,I31384,I31690,);
not I_1710 (I31376,I31690);
not I_1711 (I31712,I31673);
nand I_1712 (I31361,I31712,I31551);
nor I_1713 (I31743,I131214,I131202);
not I_1714 (I31760,I31743);
nor I_1715 (I31777,I31712,I31760);
nor I_1716 (I31794,I31418,I31777);
DFFARX1 I_1717 (I31794,I2595,I31384,I31370,);
nor I_1718 (I31825,I31478,I31760);
nor I_1719 (I31358,I31673,I31825);
nor I_1720 (I31367,I31608,I31743);
nor I_1721 (I31355,I31478,I31743);
not I_1722 (I31911,I2602);
DFFARX1 I_1723 (I88023,I2595,I31911,I31937,);
not I_1724 (I31945,I31937);
nand I_1725 (I31962,I88005,I88020);
and I_1726 (I31979,I31962,I87996);
DFFARX1 I_1727 (I31979,I2595,I31911,I32005,);
DFFARX1 I_1728 (I87999,I2595,I31911,I32022,);
and I_1729 (I32030,I32022,I88014);
nor I_1730 (I32047,I32005,I32030);
DFFARX1 I_1731 (I32047,I2595,I31911,I31879,);
nand I_1732 (I32078,I32022,I88014);
nand I_1733 (I32095,I31945,I32078);
not I_1734 (I31891,I32095);
DFFARX1 I_1735 (I88017,I2595,I31911,I32135,);
DFFARX1 I_1736 (I32135,I2595,I31911,I31900,);
nand I_1737 (I32157,I87996,I88008);
and I_1738 (I32174,I32157,I88002);
DFFARX1 I_1739 (I32174,I2595,I31911,I32200,);
DFFARX1 I_1740 (I32200,I2595,I31911,I32217,);
not I_1741 (I31903,I32217);
not I_1742 (I32239,I32200);
nand I_1743 (I31888,I32239,I32078);
nor I_1744 (I32270,I88011,I88008);
not I_1745 (I32287,I32270);
nor I_1746 (I32304,I32239,I32287);
nor I_1747 (I32321,I31945,I32304);
DFFARX1 I_1748 (I32321,I2595,I31911,I31897,);
nor I_1749 (I32352,I32005,I32287);
nor I_1750 (I31885,I32200,I32352);
nor I_1751 (I31894,I32135,I32270);
nor I_1752 (I31882,I32005,I32270);
not I_1753 (I32438,I2602);
DFFARX1 I_1754 (I302794,I2595,I32438,I32464,);
not I_1755 (I32472,I32464);
nand I_1756 (I32489,I302791,I302797);
and I_1757 (I32506,I32489,I302794);
DFFARX1 I_1758 (I32506,I2595,I32438,I32532,);
DFFARX1 I_1759 (I302797,I2595,I32438,I32549,);
and I_1760 (I32557,I32549,I302791);
nor I_1761 (I32574,I32532,I32557);
DFFARX1 I_1762 (I32574,I2595,I32438,I32406,);
nand I_1763 (I32605,I32549,I302791);
nand I_1764 (I32622,I32472,I32605);
not I_1765 (I32418,I32622);
DFFARX1 I_1766 (I302800,I2595,I32438,I32662,);
DFFARX1 I_1767 (I32662,I2595,I32438,I32427,);
nand I_1768 (I32684,I302803,I302812);
and I_1769 (I32701,I32684,I302806);
DFFARX1 I_1770 (I32701,I2595,I32438,I32727,);
DFFARX1 I_1771 (I32727,I2595,I32438,I32744,);
not I_1772 (I32430,I32744);
not I_1773 (I32766,I32727);
nand I_1774 (I32415,I32766,I32605);
nor I_1775 (I32797,I302809,I302812);
not I_1776 (I32814,I32797);
nor I_1777 (I32831,I32766,I32814);
nor I_1778 (I32848,I32472,I32831);
DFFARX1 I_1779 (I32848,I2595,I32438,I32424,);
nor I_1780 (I32879,I32532,I32814);
nor I_1781 (I32412,I32727,I32879);
nor I_1782 (I32421,I32662,I32797);
nor I_1783 (I32409,I32532,I32797);
not I_1784 (I32965,I2602);
DFFARX1 I_1785 (I94347,I2595,I32965,I32991,);
not I_1786 (I32999,I32991);
nand I_1787 (I33016,I94329,I94344);
and I_1788 (I33033,I33016,I94320);
DFFARX1 I_1789 (I33033,I2595,I32965,I33059,);
DFFARX1 I_1790 (I94323,I2595,I32965,I33076,);
and I_1791 (I33084,I33076,I94338);
nor I_1792 (I33101,I33059,I33084);
DFFARX1 I_1793 (I33101,I2595,I32965,I32933,);
nand I_1794 (I33132,I33076,I94338);
nand I_1795 (I33149,I32999,I33132);
not I_1796 (I32945,I33149);
DFFARX1 I_1797 (I94341,I2595,I32965,I33189,);
DFFARX1 I_1798 (I33189,I2595,I32965,I32954,);
nand I_1799 (I33211,I94320,I94332);
and I_1800 (I33228,I33211,I94326);
DFFARX1 I_1801 (I33228,I2595,I32965,I33254,);
DFFARX1 I_1802 (I33254,I2595,I32965,I33271,);
not I_1803 (I32957,I33271);
not I_1804 (I33293,I33254);
nand I_1805 (I32942,I33293,I33132);
nor I_1806 (I33324,I94335,I94332);
not I_1807 (I33341,I33324);
nor I_1808 (I33358,I33293,I33341);
nor I_1809 (I33375,I32999,I33358);
DFFARX1 I_1810 (I33375,I2595,I32965,I32951,);
nor I_1811 (I33406,I33059,I33341);
nor I_1812 (I32939,I33254,I33406);
nor I_1813 (I32948,I33189,I33324);
nor I_1814 (I32936,I33059,I33324);
not I_1815 (I33492,I2602);
DFFARX1 I_1816 (I236704,I2595,I33492,I33518,);
not I_1817 (I33526,I33518);
nand I_1818 (I33543,I236701,I236716);
and I_1819 (I33560,I33543,I236698);
DFFARX1 I_1820 (I33560,I2595,I33492,I33586,);
DFFARX1 I_1821 (I236695,I2595,I33492,I33603,);
and I_1822 (I33611,I33603,I236695);
nor I_1823 (I33628,I33586,I33611);
DFFARX1 I_1824 (I33628,I2595,I33492,I33460,);
nand I_1825 (I33659,I33603,I236695);
nand I_1826 (I33676,I33526,I33659);
not I_1827 (I33472,I33676);
DFFARX1 I_1828 (I236698,I2595,I33492,I33716,);
DFFARX1 I_1829 (I33716,I2595,I33492,I33481,);
nand I_1830 (I33738,I236710,I236701);
and I_1831 (I33755,I33738,I236713);
DFFARX1 I_1832 (I33755,I2595,I33492,I33781,);
DFFARX1 I_1833 (I33781,I2595,I33492,I33798,);
not I_1834 (I33484,I33798);
not I_1835 (I33820,I33781);
nand I_1836 (I33469,I33820,I33659);
nor I_1837 (I33851,I236707,I236701);
not I_1838 (I33868,I33851);
nor I_1839 (I33885,I33820,I33868);
nor I_1840 (I33902,I33526,I33885);
DFFARX1 I_1841 (I33902,I2595,I33492,I33478,);
nor I_1842 (I33933,I33586,I33868);
nor I_1843 (I33466,I33781,I33933);
nor I_1844 (I33475,I33716,I33851);
nor I_1845 (I33463,I33586,I33851);
not I_1846 (I34019,I2602);
DFFARX1 I_1847 (I372945,I2595,I34019,I34045,);
not I_1848 (I34053,I34045);
nand I_1849 (I34070,I372939,I372960);
and I_1850 (I34087,I34070,I372936);
DFFARX1 I_1851 (I34087,I2595,I34019,I34113,);
DFFARX1 I_1852 (I372957,I2595,I34019,I34130,);
and I_1853 (I34138,I34130,I372954);
nor I_1854 (I34155,I34113,I34138);
DFFARX1 I_1855 (I34155,I2595,I34019,I33987,);
nand I_1856 (I34186,I34130,I372954);
nand I_1857 (I34203,I34053,I34186);
not I_1858 (I33999,I34203);
DFFARX1 I_1859 (I372942,I2595,I34019,I34243,);
DFFARX1 I_1860 (I34243,I2595,I34019,I34008,);
nand I_1861 (I34265,I372951,I372948);
and I_1862 (I34282,I34265,I372933);
DFFARX1 I_1863 (I34282,I2595,I34019,I34308,);
DFFARX1 I_1864 (I34308,I2595,I34019,I34325,);
not I_1865 (I34011,I34325);
not I_1866 (I34347,I34308);
nand I_1867 (I33996,I34347,I34186);
nor I_1868 (I34378,I372933,I372948);
not I_1869 (I34395,I34378);
nor I_1870 (I34412,I34347,I34395);
nor I_1871 (I34429,I34053,I34412);
DFFARX1 I_1872 (I34429,I2595,I34019,I34005,);
nor I_1873 (I34460,I34113,I34395);
nor I_1874 (I33993,I34308,I34460);
nor I_1875 (I34002,I34243,I34378);
nor I_1876 (I33990,I34113,I34378);
not I_1877 (I34546,I2602);
DFFARX1 I_1878 (I133931,I2595,I34546,I34572,);
not I_1879 (I34580,I34572);
nand I_1880 (I34597,I133925,I133916);
and I_1881 (I34614,I34597,I133937);
DFFARX1 I_1882 (I34614,I2595,I34546,I34640,);
DFFARX1 I_1883 (I133919,I2595,I34546,I34657,);
and I_1884 (I34665,I34657,I133913);
nor I_1885 (I34682,I34640,I34665);
DFFARX1 I_1886 (I34682,I2595,I34546,I34514,);
nand I_1887 (I34713,I34657,I133913);
nand I_1888 (I34730,I34580,I34713);
not I_1889 (I34526,I34730);
DFFARX1 I_1890 (I133913,I2595,I34546,I34770,);
DFFARX1 I_1891 (I34770,I2595,I34546,I34535,);
nand I_1892 (I34792,I133940,I133922);
and I_1893 (I34809,I34792,I133928);
DFFARX1 I_1894 (I34809,I2595,I34546,I34835,);
DFFARX1 I_1895 (I34835,I2595,I34546,I34852,);
not I_1896 (I34538,I34852);
not I_1897 (I34874,I34835);
nand I_1898 (I34523,I34874,I34713);
nor I_1899 (I34905,I133934,I133922);
not I_1900 (I34922,I34905);
nor I_1901 (I34939,I34874,I34922);
nor I_1902 (I34956,I34580,I34939);
DFFARX1 I_1903 (I34956,I2595,I34546,I34532,);
nor I_1904 (I34987,I34640,I34922);
nor I_1905 (I34520,I34835,I34987);
nor I_1906 (I34529,I34770,I34905);
nor I_1907 (I34517,I34640,I34905);
not I_1908 (I35073,I2602);
DFFARX1 I_1909 (I325832,I2595,I35073,I35099,);
not I_1910 (I35107,I35099);
nand I_1911 (I35124,I325847,I325826);
and I_1912 (I35141,I35124,I325829);
DFFARX1 I_1913 (I35141,I2595,I35073,I35167,);
DFFARX1 I_1914 (I325850,I2595,I35073,I35184,);
and I_1915 (I35192,I35184,I325829);
nor I_1916 (I35209,I35167,I35192);
DFFARX1 I_1917 (I35209,I2595,I35073,I35041,);
nand I_1918 (I35240,I35184,I325829);
nand I_1919 (I35257,I35107,I35240);
not I_1920 (I35053,I35257);
DFFARX1 I_1921 (I325826,I2595,I35073,I35297,);
DFFARX1 I_1922 (I35297,I2595,I35073,I35062,);
nand I_1923 (I35319,I325838,I325835);
and I_1924 (I35336,I35319,I325841);
DFFARX1 I_1925 (I35336,I2595,I35073,I35362,);
DFFARX1 I_1926 (I35362,I2595,I35073,I35379,);
not I_1927 (I35065,I35379);
not I_1928 (I35401,I35362);
nand I_1929 (I35050,I35401,I35240);
nor I_1930 (I35432,I325844,I325835);
not I_1931 (I35449,I35432);
nor I_1932 (I35466,I35401,I35449);
nor I_1933 (I35483,I35107,I35466);
DFFARX1 I_1934 (I35483,I2595,I35073,I35059,);
nor I_1935 (I35514,I35167,I35449);
nor I_1936 (I35047,I35362,I35514);
nor I_1937 (I35056,I35297,I35432);
nor I_1938 (I35044,I35167,I35432);
not I_1939 (I35600,I2602);
DFFARX1 I_1940 (I369465,I2595,I35600,I35626,);
not I_1941 (I35634,I35626);
nand I_1942 (I35651,I369471,I369489);
and I_1943 (I35668,I35651,I369486);
DFFARX1 I_1944 (I35668,I2595,I35600,I35694,);
DFFARX1 I_1945 (I369483,I2595,I35600,I35711,);
and I_1946 (I35719,I35711,I369477);
nor I_1947 (I35736,I35694,I35719);
DFFARX1 I_1948 (I35736,I2595,I35600,I35568,);
nand I_1949 (I35767,I35711,I369477);
nand I_1950 (I35784,I35634,I35767);
not I_1951 (I35580,I35784);
DFFARX1 I_1952 (I369465,I2595,I35600,I35824,);
DFFARX1 I_1953 (I35824,I2595,I35600,I35589,);
nand I_1954 (I35846,I369480,I369468);
and I_1955 (I35863,I35846,I369492);
DFFARX1 I_1956 (I35863,I2595,I35600,I35889,);
DFFARX1 I_1957 (I35889,I2595,I35600,I35906,);
not I_1958 (I35592,I35906);
not I_1959 (I35928,I35889);
nand I_1960 (I35577,I35928,I35767);
nor I_1961 (I35959,I369474,I369468);
not I_1962 (I35976,I35959);
nor I_1963 (I35993,I35928,I35976);
nor I_1964 (I36010,I35634,I35993);
DFFARX1 I_1965 (I36010,I2595,I35600,I35586,);
nor I_1966 (I36041,I35694,I35976);
nor I_1967 (I35574,I35889,I36041);
nor I_1968 (I35583,I35824,I35959);
nor I_1969 (I35571,I35694,I35959);
not I_1970 (I36127,I2602);
DFFARX1 I_1971 (I299428,I2595,I36127,I36153,);
not I_1972 (I36161,I36153);
nand I_1973 (I36178,I299425,I299431);
and I_1974 (I36195,I36178,I299428);
DFFARX1 I_1975 (I36195,I2595,I36127,I36221,);
DFFARX1 I_1976 (I299431,I2595,I36127,I36238,);
and I_1977 (I36246,I36238,I299425);
nor I_1978 (I36263,I36221,I36246);
DFFARX1 I_1979 (I36263,I2595,I36127,I36095,);
nand I_1980 (I36294,I36238,I299425);
nand I_1981 (I36311,I36161,I36294);
not I_1982 (I36107,I36311);
DFFARX1 I_1983 (I299434,I2595,I36127,I36351,);
DFFARX1 I_1984 (I36351,I2595,I36127,I36116,);
nand I_1985 (I36373,I299437,I299446);
and I_1986 (I36390,I36373,I299440);
DFFARX1 I_1987 (I36390,I2595,I36127,I36416,);
DFFARX1 I_1988 (I36416,I2595,I36127,I36433,);
not I_1989 (I36119,I36433);
not I_1990 (I36455,I36416);
nand I_1991 (I36104,I36455,I36294);
nor I_1992 (I36486,I299443,I299446);
not I_1993 (I36503,I36486);
nor I_1994 (I36520,I36455,I36503);
nor I_1995 (I36537,I36161,I36520);
DFFARX1 I_1996 (I36537,I2595,I36127,I36113,);
nor I_1997 (I36568,I36221,I36503);
nor I_1998 (I36101,I36416,I36568);
nor I_1999 (I36110,I36351,I36486);
nor I_2000 (I36098,I36221,I36486);
not I_2001 (I36654,I2602);
DFFARX1 I_2002 (I159337,I2595,I36654,I36680,);
not I_2003 (I36688,I36680);
nand I_2004 (I36705,I159349,I159334);
and I_2005 (I36722,I36705,I159328);
DFFARX1 I_2006 (I36722,I2595,I36654,I36748,);
DFFARX1 I_2007 (I159343,I2595,I36654,I36765,);
and I_2008 (I36773,I36765,I159331);
nor I_2009 (I36790,I36748,I36773);
DFFARX1 I_2010 (I36790,I2595,I36654,I36622,);
nand I_2011 (I36821,I36765,I159331);
nand I_2012 (I36838,I36688,I36821);
not I_2013 (I36634,I36838);
DFFARX1 I_2014 (I159340,I2595,I36654,I36878,);
DFFARX1 I_2015 (I36878,I2595,I36654,I36643,);
nand I_2016 (I36900,I159346,I159352);
and I_2017 (I36917,I36900,I159328);
DFFARX1 I_2018 (I36917,I2595,I36654,I36943,);
DFFARX1 I_2019 (I36943,I2595,I36654,I36960,);
not I_2020 (I36646,I36960);
not I_2021 (I36982,I36943);
nand I_2022 (I36631,I36982,I36821);
nor I_2023 (I37013,I159331,I159352);
not I_2024 (I37030,I37013);
nor I_2025 (I37047,I36982,I37030);
nor I_2026 (I37064,I36688,I37047);
DFFARX1 I_2027 (I37064,I2595,I36654,I36640,);
nor I_2028 (I37095,I36748,I37030);
nor I_2029 (I36628,I36943,I37095);
nor I_2030 (I36637,I36878,I37013);
nor I_2031 (I36625,I36748,I37013);
not I_2032 (I37181,I2602);
DFFARX1 I_2033 (I126315,I2595,I37181,I37207,);
not I_2034 (I37215,I37207);
nand I_2035 (I37232,I126309,I126300);
and I_2036 (I37249,I37232,I126321);
DFFARX1 I_2037 (I37249,I2595,I37181,I37275,);
DFFARX1 I_2038 (I126303,I2595,I37181,I37292,);
and I_2039 (I37300,I37292,I126297);
nor I_2040 (I37317,I37275,I37300);
DFFARX1 I_2041 (I37317,I2595,I37181,I37149,);
nand I_2042 (I37348,I37292,I126297);
nand I_2043 (I37365,I37215,I37348);
not I_2044 (I37161,I37365);
DFFARX1 I_2045 (I126297,I2595,I37181,I37405,);
DFFARX1 I_2046 (I37405,I2595,I37181,I37170,);
nand I_2047 (I37427,I126324,I126306);
and I_2048 (I37444,I37427,I126312);
DFFARX1 I_2049 (I37444,I2595,I37181,I37470,);
DFFARX1 I_2050 (I37470,I2595,I37181,I37487,);
not I_2051 (I37173,I37487);
not I_2052 (I37509,I37470);
nand I_2053 (I37158,I37509,I37348);
nor I_2054 (I37540,I126318,I126306);
not I_2055 (I37557,I37540);
nor I_2056 (I37574,I37509,I37557);
nor I_2057 (I37591,I37215,I37574);
DFFARX1 I_2058 (I37591,I2595,I37181,I37167,);
nor I_2059 (I37622,I37275,I37557);
nor I_2060 (I37155,I37470,I37622);
nor I_2061 (I37164,I37405,I37540);
nor I_2062 (I37152,I37275,I37540);
not I_2063 (I37708,I2602);
DFFARX1 I_2064 (I356228,I2595,I37708,I37734,);
not I_2065 (I37742,I37734);
nand I_2066 (I37759,I356222,I356243);
and I_2067 (I37776,I37759,I356234);
DFFARX1 I_2068 (I37776,I2595,I37708,I37802,);
DFFARX1 I_2069 (I356225,I2595,I37708,I37819,);
and I_2070 (I37827,I37819,I356237);
nor I_2071 (I37844,I37802,I37827);
DFFARX1 I_2072 (I37844,I2595,I37708,I37676,);
nand I_2073 (I37875,I37819,I356237);
nand I_2074 (I37892,I37742,I37875);
not I_2075 (I37688,I37892);
DFFARX1 I_2076 (I356225,I2595,I37708,I37932,);
DFFARX1 I_2077 (I37932,I2595,I37708,I37697,);
nand I_2078 (I37954,I356246,I356231);
and I_2079 (I37971,I37954,I356222);
DFFARX1 I_2080 (I37971,I2595,I37708,I37997,);
DFFARX1 I_2081 (I37997,I2595,I37708,I38014,);
not I_2082 (I37700,I38014);
not I_2083 (I38036,I37997);
nand I_2084 (I37685,I38036,I37875);
nor I_2085 (I38067,I356240,I356231);
not I_2086 (I38084,I38067);
nor I_2087 (I38101,I38036,I38084);
nor I_2088 (I38118,I37742,I38101);
DFFARX1 I_2089 (I38118,I2595,I37708,I37694,);
nor I_2090 (I38149,I37802,I38084);
nor I_2091 (I37682,I37997,I38149);
nor I_2092 (I37691,I37932,I38067);
nor I_2093 (I37679,I37802,I38067);
not I_2094 (I38235,I2602);
DFFARX1 I_2095 (I346980,I2595,I38235,I38261,);
not I_2096 (I38269,I38261);
nand I_2097 (I38286,I346974,I346995);
and I_2098 (I38303,I38286,I346986);
DFFARX1 I_2099 (I38303,I2595,I38235,I38329,);
DFFARX1 I_2100 (I346977,I2595,I38235,I38346,);
and I_2101 (I38354,I38346,I346989);
nor I_2102 (I38371,I38329,I38354);
DFFARX1 I_2103 (I38371,I2595,I38235,I38203,);
nand I_2104 (I38402,I38346,I346989);
nand I_2105 (I38419,I38269,I38402);
not I_2106 (I38215,I38419);
DFFARX1 I_2107 (I346977,I2595,I38235,I38459,);
DFFARX1 I_2108 (I38459,I2595,I38235,I38224,);
nand I_2109 (I38481,I346998,I346983);
and I_2110 (I38498,I38481,I346974);
DFFARX1 I_2111 (I38498,I2595,I38235,I38524,);
DFFARX1 I_2112 (I38524,I2595,I38235,I38541,);
not I_2113 (I38227,I38541);
not I_2114 (I38563,I38524);
nand I_2115 (I38212,I38563,I38402);
nor I_2116 (I38594,I346992,I346983);
not I_2117 (I38611,I38594);
nor I_2118 (I38628,I38563,I38611);
nor I_2119 (I38645,I38269,I38628);
DFFARX1 I_2120 (I38645,I2595,I38235,I38221,);
nor I_2121 (I38676,I38329,I38611);
nor I_2122 (I38209,I38524,I38676);
nor I_2123 (I38218,I38459,I38594);
nor I_2124 (I38206,I38329,I38594);
not I_2125 (I38762,I2602);
DFFARX1 I_2126 (I233542,I2595,I38762,I38788,);
not I_2127 (I38796,I38788);
nand I_2128 (I38813,I233539,I233554);
and I_2129 (I38830,I38813,I233536);
DFFARX1 I_2130 (I38830,I2595,I38762,I38856,);
DFFARX1 I_2131 (I233533,I2595,I38762,I38873,);
and I_2132 (I38881,I38873,I233533);
nor I_2133 (I38898,I38856,I38881);
DFFARX1 I_2134 (I38898,I2595,I38762,I38730,);
nand I_2135 (I38929,I38873,I233533);
nand I_2136 (I38946,I38796,I38929);
not I_2137 (I38742,I38946);
DFFARX1 I_2138 (I233536,I2595,I38762,I38986,);
DFFARX1 I_2139 (I38986,I2595,I38762,I38751,);
nand I_2140 (I39008,I233548,I233539);
and I_2141 (I39025,I39008,I233551);
DFFARX1 I_2142 (I39025,I2595,I38762,I39051,);
DFFARX1 I_2143 (I39051,I2595,I38762,I39068,);
not I_2144 (I38754,I39068);
not I_2145 (I39090,I39051);
nand I_2146 (I38739,I39090,I38929);
nor I_2147 (I39121,I233545,I233539);
not I_2148 (I39138,I39121);
nor I_2149 (I39155,I39090,I39138);
nor I_2150 (I39172,I38796,I39155);
DFFARX1 I_2151 (I39172,I2595,I38762,I38748,);
nor I_2152 (I39203,I38856,I39138);
nor I_2153 (I38736,I39051,I39203);
nor I_2154 (I38745,I38986,I39121);
nor I_2155 (I38733,I38856,I39121);
not I_2156 (I39289,I2602);
DFFARX1 I_2157 (I129035,I2595,I39289,I39315,);
not I_2158 (I39323,I39315);
nand I_2159 (I39340,I129029,I129020);
and I_2160 (I39357,I39340,I129041);
DFFARX1 I_2161 (I39357,I2595,I39289,I39383,);
DFFARX1 I_2162 (I129023,I2595,I39289,I39400,);
and I_2163 (I39408,I39400,I129017);
nor I_2164 (I39425,I39383,I39408);
DFFARX1 I_2165 (I39425,I2595,I39289,I39257,);
nand I_2166 (I39456,I39400,I129017);
nand I_2167 (I39473,I39323,I39456);
not I_2168 (I39269,I39473);
DFFARX1 I_2169 (I129017,I2595,I39289,I39513,);
DFFARX1 I_2170 (I39513,I2595,I39289,I39278,);
nand I_2171 (I39535,I129044,I129026);
and I_2172 (I39552,I39535,I129032);
DFFARX1 I_2173 (I39552,I2595,I39289,I39578,);
DFFARX1 I_2174 (I39578,I2595,I39289,I39595,);
not I_2175 (I39281,I39595);
not I_2176 (I39617,I39578);
nand I_2177 (I39266,I39617,I39456);
nor I_2178 (I39648,I129038,I129026);
not I_2179 (I39665,I39648);
nor I_2180 (I39682,I39617,I39665);
nor I_2181 (I39699,I39323,I39682);
DFFARX1 I_2182 (I39699,I2595,I39289,I39275,);
nor I_2183 (I39730,I39383,I39665);
nor I_2184 (I39263,I39578,I39730);
nor I_2185 (I39272,I39513,I39648);
nor I_2186 (I39260,I39383,I39648);
not I_2187 (I39816,I2602);
DFFARX1 I_2188 (I78845,I2595,I39816,I39842,);
not I_2189 (I39850,I39842);
nand I_2190 (I39867,I78839,I78833);
and I_2191 (I39884,I39867,I78854);
DFFARX1 I_2192 (I39884,I2595,I39816,I39910,);
DFFARX1 I_2193 (I78851,I2595,I39816,I39927,);
and I_2194 (I39935,I39927,I78848);
nor I_2195 (I39952,I39910,I39935);
DFFARX1 I_2196 (I39952,I2595,I39816,I39784,);
nand I_2197 (I39983,I39927,I78848);
nand I_2198 (I40000,I39850,I39983);
not I_2199 (I39796,I40000);
DFFARX1 I_2200 (I78833,I2595,I39816,I40040,);
DFFARX1 I_2201 (I40040,I2595,I39816,I39805,);
nand I_2202 (I40062,I78836,I78836);
and I_2203 (I40079,I40062,I78857);
DFFARX1 I_2204 (I40079,I2595,I39816,I40105,);
DFFARX1 I_2205 (I40105,I2595,I39816,I40122,);
not I_2206 (I39808,I40122);
not I_2207 (I40144,I40105);
nand I_2208 (I39793,I40144,I39983);
nor I_2209 (I40175,I78842,I78836);
not I_2210 (I40192,I40175);
nor I_2211 (I40209,I40144,I40192);
nor I_2212 (I40226,I39850,I40209);
DFFARX1 I_2213 (I40226,I2595,I39816,I39802,);
nor I_2214 (I40257,I39910,I40192);
nor I_2215 (I39790,I40105,I40257);
nor I_2216 (I39799,I40040,I40175);
nor I_2217 (I39787,I39910,I40175);
not I_2218 (I40343,I2602);
DFFARX1 I_2219 (I344804,I2595,I40343,I40369,);
not I_2220 (I40377,I40369);
nand I_2221 (I40394,I344798,I344819);
and I_2222 (I40411,I40394,I344810);
DFFARX1 I_2223 (I40411,I2595,I40343,I40437,);
DFFARX1 I_2224 (I344801,I2595,I40343,I40454,);
and I_2225 (I40462,I40454,I344813);
nor I_2226 (I40479,I40437,I40462);
DFFARX1 I_2227 (I40479,I2595,I40343,I40311,);
nand I_2228 (I40510,I40454,I344813);
nand I_2229 (I40527,I40377,I40510);
not I_2230 (I40323,I40527);
DFFARX1 I_2231 (I344801,I2595,I40343,I40567,);
DFFARX1 I_2232 (I40567,I2595,I40343,I40332,);
nand I_2233 (I40589,I344822,I344807);
and I_2234 (I40606,I40589,I344798);
DFFARX1 I_2235 (I40606,I2595,I40343,I40632,);
DFFARX1 I_2236 (I40632,I2595,I40343,I40649,);
not I_2237 (I40335,I40649);
not I_2238 (I40671,I40632);
nand I_2239 (I40320,I40671,I40510);
nor I_2240 (I40702,I344816,I344807);
not I_2241 (I40719,I40702);
nor I_2242 (I40736,I40671,I40719);
nor I_2243 (I40753,I40377,I40736);
DFFARX1 I_2244 (I40753,I2595,I40343,I40329,);
nor I_2245 (I40784,I40437,I40719);
nor I_2246 (I40317,I40632,I40784);
nor I_2247 (I40326,I40567,I40702);
nor I_2248 (I40314,I40437,I40702);
not I_2249 (I40870,I2602);
DFFARX1 I_2250 (I355140,I2595,I40870,I40896,);
not I_2251 (I40904,I40896);
nand I_2252 (I40921,I355134,I355155);
and I_2253 (I40938,I40921,I355146);
DFFARX1 I_2254 (I40938,I2595,I40870,I40964,);
DFFARX1 I_2255 (I355137,I2595,I40870,I40981,);
and I_2256 (I40989,I40981,I355149);
nor I_2257 (I41006,I40964,I40989);
DFFARX1 I_2258 (I41006,I2595,I40870,I40838,);
nand I_2259 (I41037,I40981,I355149);
nand I_2260 (I41054,I40904,I41037);
not I_2261 (I40850,I41054);
DFFARX1 I_2262 (I355137,I2595,I40870,I41094,);
DFFARX1 I_2263 (I41094,I2595,I40870,I40859,);
nand I_2264 (I41116,I355158,I355143);
and I_2265 (I41133,I41116,I355134);
DFFARX1 I_2266 (I41133,I2595,I40870,I41159,);
DFFARX1 I_2267 (I41159,I2595,I40870,I41176,);
not I_2268 (I40862,I41176);
not I_2269 (I41198,I41159);
nand I_2270 (I40847,I41198,I41037);
nor I_2271 (I41229,I355152,I355143);
not I_2272 (I41246,I41229);
nor I_2273 (I41263,I41198,I41246);
nor I_2274 (I41280,I40904,I41263);
DFFARX1 I_2275 (I41280,I2595,I40870,I40856,);
nor I_2276 (I41311,I40964,I41246);
nor I_2277 (I40844,I41159,I41311);
nor I_2278 (I40853,I41094,I41229);
nor I_2279 (I40841,I40964,I41229);
not I_2280 (I41397,I2602);
DFFARX1 I_2281 (I331034,I2595,I41397,I41423,);
not I_2282 (I41431,I41423);
nand I_2283 (I41448,I331049,I331028);
and I_2284 (I41465,I41448,I331031);
DFFARX1 I_2285 (I41465,I2595,I41397,I41491,);
DFFARX1 I_2286 (I331052,I2595,I41397,I41508,);
and I_2287 (I41516,I41508,I331031);
nor I_2288 (I41533,I41491,I41516);
DFFARX1 I_2289 (I41533,I2595,I41397,I41365,);
nand I_2290 (I41564,I41508,I331031);
nand I_2291 (I41581,I41431,I41564);
not I_2292 (I41377,I41581);
DFFARX1 I_2293 (I331028,I2595,I41397,I41621,);
DFFARX1 I_2294 (I41621,I2595,I41397,I41386,);
nand I_2295 (I41643,I331040,I331037);
and I_2296 (I41660,I41643,I331043);
DFFARX1 I_2297 (I41660,I2595,I41397,I41686,);
DFFARX1 I_2298 (I41686,I2595,I41397,I41703,);
not I_2299 (I41389,I41703);
not I_2300 (I41725,I41686);
nand I_2301 (I41374,I41725,I41564);
nor I_2302 (I41756,I331046,I331037);
not I_2303 (I41773,I41756);
nor I_2304 (I41790,I41725,I41773);
nor I_2305 (I41807,I41431,I41790);
DFFARX1 I_2306 (I41807,I2595,I41397,I41383,);
nor I_2307 (I41838,I41491,I41773);
nor I_2308 (I41371,I41686,I41838);
nor I_2309 (I41380,I41621,I41756);
nor I_2310 (I41368,I41491,I41756);
not I_2311 (I41924,I2602);
DFFARX1 I_2312 (I22417,I2595,I41924,I41950,);
not I_2313 (I41958,I41950);
nand I_2314 (I41975,I22405,I22411);
and I_2315 (I41992,I41975,I22414);
DFFARX1 I_2316 (I41992,I2595,I41924,I42018,);
DFFARX1 I_2317 (I22396,I2595,I41924,I42035,);
and I_2318 (I42043,I42035,I22402);
nor I_2319 (I42060,I42018,I42043);
DFFARX1 I_2320 (I42060,I2595,I41924,I41892,);
nand I_2321 (I42091,I42035,I22402);
nand I_2322 (I42108,I41958,I42091);
not I_2323 (I41904,I42108);
DFFARX1 I_2324 (I22396,I2595,I41924,I42148,);
DFFARX1 I_2325 (I42148,I2595,I41924,I41913,);
nand I_2326 (I42170,I22399,I22393);
and I_2327 (I42187,I42170,I22408);
DFFARX1 I_2328 (I42187,I2595,I41924,I42213,);
DFFARX1 I_2329 (I42213,I2595,I41924,I42230,);
not I_2330 (I41916,I42230);
not I_2331 (I42252,I42213);
nand I_2332 (I41901,I42252,I42091);
nor I_2333 (I42283,I22393,I22393);
not I_2334 (I42300,I42283);
nor I_2335 (I42317,I42252,I42300);
nor I_2336 (I42334,I41958,I42317);
DFFARX1 I_2337 (I42334,I2595,I41924,I41910,);
nor I_2338 (I42365,I42018,I42300);
nor I_2339 (I41898,I42213,I42365);
nor I_2340 (I41907,I42148,I42283);
nor I_2341 (I41895,I42018,I42283);
not I_2342 (I42451,I2602);
DFFARX1 I_2343 (I341438,I2595,I42451,I42477,);
not I_2344 (I42485,I42477);
nand I_2345 (I42502,I341453,I341432);
and I_2346 (I42519,I42502,I341435);
DFFARX1 I_2347 (I42519,I2595,I42451,I42545,);
DFFARX1 I_2348 (I341456,I2595,I42451,I42562,);
and I_2349 (I42570,I42562,I341435);
nor I_2350 (I42587,I42545,I42570);
DFFARX1 I_2351 (I42587,I2595,I42451,I42419,);
nand I_2352 (I42618,I42562,I341435);
nand I_2353 (I42635,I42485,I42618);
not I_2354 (I42431,I42635);
DFFARX1 I_2355 (I341432,I2595,I42451,I42675,);
DFFARX1 I_2356 (I42675,I2595,I42451,I42440,);
nand I_2357 (I42697,I341444,I341441);
and I_2358 (I42714,I42697,I341447);
DFFARX1 I_2359 (I42714,I2595,I42451,I42740,);
DFFARX1 I_2360 (I42740,I2595,I42451,I42757,);
not I_2361 (I42443,I42757);
not I_2362 (I42779,I42740);
nand I_2363 (I42428,I42779,I42618);
nor I_2364 (I42810,I341450,I341441);
not I_2365 (I42827,I42810);
nor I_2366 (I42844,I42779,I42827);
nor I_2367 (I42861,I42485,I42844);
DFFARX1 I_2368 (I42861,I2595,I42451,I42437,);
nor I_2369 (I42892,I42545,I42827);
nor I_2370 (I42425,I42740,I42892);
nor I_2371 (I42434,I42675,I42810);
nor I_2372 (I42422,I42545,I42810);
not I_2373 (I42978,I2602);
DFFARX1 I_2374 (I303916,I2595,I42978,I43004,);
not I_2375 (I43012,I43004);
nand I_2376 (I43029,I303913,I303919);
and I_2377 (I43046,I43029,I303916);
DFFARX1 I_2378 (I43046,I2595,I42978,I43072,);
DFFARX1 I_2379 (I303919,I2595,I42978,I43089,);
and I_2380 (I43097,I43089,I303913);
nor I_2381 (I43114,I43072,I43097);
DFFARX1 I_2382 (I43114,I2595,I42978,I42946,);
nand I_2383 (I43145,I43089,I303913);
nand I_2384 (I43162,I43012,I43145);
not I_2385 (I42958,I43162);
DFFARX1 I_2386 (I303922,I2595,I42978,I43202,);
DFFARX1 I_2387 (I43202,I2595,I42978,I42967,);
nand I_2388 (I43224,I303925,I303934);
and I_2389 (I43241,I43224,I303928);
DFFARX1 I_2390 (I43241,I2595,I42978,I43267,);
DFFARX1 I_2391 (I43267,I2595,I42978,I43284,);
not I_2392 (I42970,I43284);
not I_2393 (I43306,I43267);
nand I_2394 (I42955,I43306,I43145);
nor I_2395 (I43337,I303931,I303934);
not I_2396 (I43354,I43337);
nor I_2397 (I43371,I43306,I43354);
nor I_2398 (I43388,I43012,I43371);
DFFARX1 I_2399 (I43388,I2595,I42978,I42964,);
nor I_2400 (I43419,I43072,I43354);
nor I_2401 (I42952,I43267,I43419);
nor I_2402 (I42961,I43202,I43337);
nor I_2403 (I42949,I43072,I43337);
not I_2404 (I43505,I2602);
DFFARX1 I_2405 (I285460,I2595,I43505,I43531,);
not I_2406 (I43539,I43531);
nand I_2407 (I43556,I285478,I285472);
and I_2408 (I43573,I43556,I285451);
DFFARX1 I_2409 (I43573,I2595,I43505,I43599,);
DFFARX1 I_2410 (I285469,I2595,I43505,I43616,);
and I_2411 (I43624,I43616,I285454);
nor I_2412 (I43641,I43599,I43624);
DFFARX1 I_2413 (I43641,I2595,I43505,I43473,);
nand I_2414 (I43672,I43616,I285454);
nand I_2415 (I43689,I43539,I43672);
not I_2416 (I43485,I43689);
DFFARX1 I_2417 (I285466,I2595,I43505,I43729,);
DFFARX1 I_2418 (I43729,I2595,I43505,I43494,);
nand I_2419 (I43751,I285475,I285463);
and I_2420 (I43768,I43751,I285457);
DFFARX1 I_2421 (I43768,I2595,I43505,I43794,);
DFFARX1 I_2422 (I43794,I2595,I43505,I43811,);
not I_2423 (I43497,I43811);
not I_2424 (I43833,I43794);
nand I_2425 (I43482,I43833,I43672);
nor I_2426 (I43864,I285451,I285463);
not I_2427 (I43881,I43864);
nor I_2428 (I43898,I43833,I43881);
nor I_2429 (I43915,I43539,I43898);
DFFARX1 I_2430 (I43915,I2595,I43505,I43491,);
nor I_2431 (I43946,I43599,I43881);
nor I_2432 (I43479,I43794,I43946);
nor I_2433 (I43488,I43729,I43864);
nor I_2434 (I43476,I43599,I43864);
not I_2435 (I44032,I2602);
DFFARX1 I_2436 (I195754,I2595,I44032,I44058,);
not I_2437 (I44066,I44058);
nand I_2438 (I44083,I195745,I195763);
and I_2439 (I44100,I44083,I195742);
DFFARX1 I_2440 (I44100,I2595,I44032,I44126,);
DFFARX1 I_2441 (I195745,I2595,I44032,I44143,);
and I_2442 (I44151,I44143,I195748);
nor I_2443 (I44168,I44126,I44151);
DFFARX1 I_2444 (I44168,I2595,I44032,I44000,);
nand I_2445 (I44199,I44143,I195748);
nand I_2446 (I44216,I44066,I44199);
not I_2447 (I44012,I44216);
DFFARX1 I_2448 (I195742,I2595,I44032,I44256,);
DFFARX1 I_2449 (I44256,I2595,I44032,I44021,);
nand I_2450 (I44278,I195760,I195751);
and I_2451 (I44295,I44278,I195766);
DFFARX1 I_2452 (I44295,I2595,I44032,I44321,);
DFFARX1 I_2453 (I44321,I2595,I44032,I44338,);
not I_2454 (I44024,I44338);
not I_2455 (I44360,I44321);
nand I_2456 (I44009,I44360,I44199);
nor I_2457 (I44391,I195757,I195751);
not I_2458 (I44408,I44391);
nor I_2459 (I44425,I44360,I44408);
nor I_2460 (I44442,I44066,I44425);
DFFARX1 I_2461 (I44442,I2595,I44032,I44018,);
nor I_2462 (I44473,I44126,I44408);
nor I_2463 (I44006,I44321,I44473);
nor I_2464 (I44015,I44256,I44391);
nor I_2465 (I44003,I44126,I44391);
not I_2466 (I44559,I2602);
DFFARX1 I_2467 (I12404,I2595,I44559,I44585,);
not I_2468 (I44593,I44585);
nand I_2469 (I44610,I12392,I12398);
and I_2470 (I44627,I44610,I12401);
DFFARX1 I_2471 (I44627,I2595,I44559,I44653,);
DFFARX1 I_2472 (I12383,I2595,I44559,I44670,);
and I_2473 (I44678,I44670,I12389);
nor I_2474 (I44695,I44653,I44678);
DFFARX1 I_2475 (I44695,I2595,I44559,I44527,);
nand I_2476 (I44726,I44670,I12389);
nand I_2477 (I44743,I44593,I44726);
not I_2478 (I44539,I44743);
DFFARX1 I_2479 (I12383,I2595,I44559,I44783,);
DFFARX1 I_2480 (I44783,I2595,I44559,I44548,);
nand I_2481 (I44805,I12386,I12380);
and I_2482 (I44822,I44805,I12395);
DFFARX1 I_2483 (I44822,I2595,I44559,I44848,);
DFFARX1 I_2484 (I44848,I2595,I44559,I44865,);
not I_2485 (I44551,I44865);
not I_2486 (I44887,I44848);
nand I_2487 (I44536,I44887,I44726);
nor I_2488 (I44918,I12380,I12380);
not I_2489 (I44935,I44918);
nor I_2490 (I44952,I44887,I44935);
nor I_2491 (I44969,I44593,I44952);
DFFARX1 I_2492 (I44969,I2595,I44559,I44545,);
nor I_2493 (I45000,I44653,I44935);
nor I_2494 (I44533,I44848,I45000);
nor I_2495 (I44542,I44783,I44918);
nor I_2496 (I44530,I44653,I44918);
not I_2497 (I45086,I2602);
DFFARX1 I_2498 (I16620,I2595,I45086,I45112,);
not I_2499 (I45120,I45112);
nand I_2500 (I45137,I16608,I16614);
and I_2501 (I45154,I45137,I16617);
DFFARX1 I_2502 (I45154,I2595,I45086,I45180,);
DFFARX1 I_2503 (I16599,I2595,I45086,I45197,);
and I_2504 (I45205,I45197,I16605);
nor I_2505 (I45222,I45180,I45205);
DFFARX1 I_2506 (I45222,I2595,I45086,I45054,);
nand I_2507 (I45253,I45197,I16605);
nand I_2508 (I45270,I45120,I45253);
not I_2509 (I45066,I45270);
DFFARX1 I_2510 (I16599,I2595,I45086,I45310,);
DFFARX1 I_2511 (I45310,I2595,I45086,I45075,);
nand I_2512 (I45332,I16602,I16596);
and I_2513 (I45349,I45332,I16611);
DFFARX1 I_2514 (I45349,I2595,I45086,I45375,);
DFFARX1 I_2515 (I45375,I2595,I45086,I45392,);
not I_2516 (I45078,I45392);
not I_2517 (I45414,I45375);
nand I_2518 (I45063,I45414,I45253);
nor I_2519 (I45445,I16596,I16596);
not I_2520 (I45462,I45445);
nor I_2521 (I45479,I45414,I45462);
nor I_2522 (I45496,I45120,I45479);
DFFARX1 I_2523 (I45496,I2595,I45086,I45072,);
nor I_2524 (I45527,I45180,I45462);
nor I_2525 (I45060,I45375,I45527);
nor I_2526 (I45069,I45310,I45445);
nor I_2527 (I45057,I45180,I45445);
not I_2528 (I45613,I2602);
DFFARX1 I_2529 (I318318,I2595,I45613,I45639,);
not I_2530 (I45647,I45639);
nand I_2531 (I45664,I318333,I318312);
and I_2532 (I45681,I45664,I318315);
DFFARX1 I_2533 (I45681,I2595,I45613,I45707,);
DFFARX1 I_2534 (I318336,I2595,I45613,I45724,);
and I_2535 (I45732,I45724,I318315);
nor I_2536 (I45749,I45707,I45732);
DFFARX1 I_2537 (I45749,I2595,I45613,I45581,);
nand I_2538 (I45780,I45724,I318315);
nand I_2539 (I45797,I45647,I45780);
not I_2540 (I45593,I45797);
DFFARX1 I_2541 (I318312,I2595,I45613,I45837,);
DFFARX1 I_2542 (I45837,I2595,I45613,I45602,);
nand I_2543 (I45859,I318324,I318321);
and I_2544 (I45876,I45859,I318327);
DFFARX1 I_2545 (I45876,I2595,I45613,I45902,);
DFFARX1 I_2546 (I45902,I2595,I45613,I45919,);
not I_2547 (I45605,I45919);
not I_2548 (I45941,I45902);
nand I_2549 (I45590,I45941,I45780);
nor I_2550 (I45972,I318330,I318321);
not I_2551 (I45989,I45972);
nor I_2552 (I46006,I45941,I45989);
nor I_2553 (I46023,I45647,I46006);
DFFARX1 I_2554 (I46023,I2595,I45613,I45599,);
nor I_2555 (I46054,I45707,I45989);
nor I_2556 (I45587,I45902,I46054);
nor I_2557 (I45596,I45837,I45972);
nor I_2558 (I45584,I45707,I45972);
not I_2559 (I46143,I2602);
DFFARX1 I_2560 (I298873,I2595,I46143,I46169,);
not I_2561 (I46177,I46169);
DFFARX1 I_2562 (I298867,I2595,I46143,I46203,);
not I_2563 (I46211,I298867);
or I_2564 (I46228,I298885,I298867);
nor I_2565 (I46245,I46203,I298885);
nand I_2566 (I46120,I46211,I46245);
nor I_2567 (I46276,I298870,I298885);
nand I_2568 (I46114,I46276,I46211);
not I_2569 (I46307,I298876);
nand I_2570 (I46324,I46211,I46307);
nor I_2571 (I46341,I298864,I298882);
not I_2572 (I46358,I46341);
nor I_2573 (I46375,I46358,I46324);
nor I_2574 (I46392,I46276,I46375);
DFFARX1 I_2575 (I46392,I2595,I46143,I46129,);
nor I_2576 (I46126,I46341,I46228);
DFFARX1 I_2577 (I46341,I2595,I46143,I46132,);
nor I_2578 (I46451,I46307,I298864);
nor I_2579 (I46468,I46451,I298867);
nor I_2580 (I46485,I298864,I298870);
DFFARX1 I_2581 (I46485,I2595,I46143,I46511,);
nor I_2582 (I46111,I46511,I46468);
DFFARX1 I_2583 (I46511,I2595,I46143,I46542,);
nand I_2584 (I46550,I46542,I298879);
nor I_2585 (I46135,I46177,I46550);
not I_2586 (I46581,I46511);
nand I_2587 (I46598,I46581,I298879);
nor I_2588 (I46615,I46177,I46598);
nor I_2589 (I46117,I46203,I46615);
nor I_2590 (I46646,I298864,I298870);
nor I_2591 (I46663,I46203,I46646);
DFFARX1 I_2592 (I46663,I2595,I46143,I46108,);
and I_2593 (I46123,I46276,I298864);
not I_2594 (I46738,I2602);
DFFARX1 I_2595 (I222908,I2595,I46738,I46764,);
not I_2596 (I46772,I46764);
DFFARX1 I_2597 (I222929,I2595,I46738,I46798,);
not I_2598 (I46806,I222908);
or I_2599 (I46823,I222920,I222908);
nor I_2600 (I46840,I46798,I222920);
nand I_2601 (I46715,I46806,I46840);
nor I_2602 (I46871,I222917,I222920);
nand I_2603 (I46709,I46871,I46806);
not I_2604 (I46902,I222926);
nand I_2605 (I46919,I46806,I46902);
nor I_2606 (I46936,I222911,I222911);
not I_2607 (I46953,I46936);
nor I_2608 (I46970,I46953,I46919);
nor I_2609 (I46987,I46871,I46970);
DFFARX1 I_2610 (I46987,I2595,I46738,I46724,);
nor I_2611 (I46721,I46936,I46823);
DFFARX1 I_2612 (I46936,I2595,I46738,I46727,);
nor I_2613 (I47046,I46902,I222911);
nor I_2614 (I47063,I47046,I222908);
nor I_2615 (I47080,I222932,I222914);
DFFARX1 I_2616 (I47080,I2595,I46738,I47106,);
nor I_2617 (I46706,I47106,I47063);
DFFARX1 I_2618 (I47106,I2595,I46738,I47137,);
nand I_2619 (I47145,I47137,I222923);
nor I_2620 (I46730,I46772,I47145);
not I_2621 (I47176,I47106);
nand I_2622 (I47193,I47176,I222923);
nor I_2623 (I47210,I46772,I47193);
nor I_2624 (I46712,I46798,I47210);
nor I_2625 (I47241,I222932,I222917);
nor I_2626 (I47258,I46798,I47241);
DFFARX1 I_2627 (I47258,I2595,I46738,I46703,);
and I_2628 (I46718,I46871,I222932);
not I_2629 (I47333,I2602);
DFFARX1 I_2630 (I75287,I2595,I47333,I47359,);
not I_2631 (I47367,I47359);
DFFARX1 I_2632 (I75281,I2595,I47333,I47393,);
not I_2633 (I47401,I75266);
or I_2634 (I47418,I75275,I75266);
nor I_2635 (I47435,I47393,I75275);
nand I_2636 (I47310,I47401,I47435);
nor I_2637 (I47466,I75263,I75275);
nand I_2638 (I47304,I47466,I47401);
not I_2639 (I47497,I75269);
nand I_2640 (I47514,I47401,I47497);
nor I_2641 (I47531,I75272,I75284);
not I_2642 (I47548,I47531);
nor I_2643 (I47565,I47548,I47514);
nor I_2644 (I47582,I47466,I47565);
DFFARX1 I_2645 (I47582,I2595,I47333,I47319,);
nor I_2646 (I47316,I47531,I47418);
DFFARX1 I_2647 (I47531,I2595,I47333,I47322,);
nor I_2648 (I47641,I47497,I75272);
nor I_2649 (I47658,I47641,I75266);
nor I_2650 (I47675,I75278,I75266);
DFFARX1 I_2651 (I47675,I2595,I47333,I47701,);
nor I_2652 (I47301,I47701,I47658);
DFFARX1 I_2653 (I47701,I2595,I47333,I47732,);
nand I_2654 (I47740,I47732,I75263);
nor I_2655 (I47325,I47367,I47740);
not I_2656 (I47771,I47701);
nand I_2657 (I47788,I47771,I75263);
nor I_2658 (I47805,I47367,I47788);
nor I_2659 (I47307,I47393,I47805);
nor I_2660 (I47836,I75278,I75263);
nor I_2661 (I47853,I47393,I47836);
DFFARX1 I_2662 (I47853,I2595,I47333,I47298,);
and I_2663 (I47313,I47466,I75278);
not I_2664 (I47928,I2602);
DFFARX1 I_2665 (I132849,I2595,I47928,I47954,);
not I_2666 (I47962,I47954);
DFFARX1 I_2667 (I132843,I2595,I47928,I47988,);
not I_2668 (I47996,I132840);
or I_2669 (I48013,I132831,I132840);
nor I_2670 (I48030,I47988,I132831);
nand I_2671 (I47905,I47996,I48030);
nor I_2672 (I48061,I132834,I132831);
nand I_2673 (I47899,I48061,I47996);
not I_2674 (I48092,I132837);
nand I_2675 (I48109,I47996,I48092);
nor I_2676 (I48126,I132825,I132852);
not I_2677 (I48143,I48126);
nor I_2678 (I48160,I48143,I48109);
nor I_2679 (I48177,I48061,I48160);
DFFARX1 I_2680 (I48177,I2595,I47928,I47914,);
nor I_2681 (I47911,I48126,I48013);
DFFARX1 I_2682 (I48126,I2595,I47928,I47917,);
nor I_2683 (I48236,I48092,I132825);
nor I_2684 (I48253,I48236,I132840);
nor I_2685 (I48270,I132828,I132825);
DFFARX1 I_2686 (I48270,I2595,I47928,I48296,);
nor I_2687 (I47896,I48296,I48253);
DFFARX1 I_2688 (I48296,I2595,I47928,I48327,);
nand I_2689 (I48335,I48327,I132846);
nor I_2690 (I47920,I47962,I48335);
not I_2691 (I48366,I48296);
nand I_2692 (I48383,I48366,I132846);
nor I_2693 (I48400,I47962,I48383);
nor I_2694 (I47902,I47988,I48400);
nor I_2695 (I48431,I132828,I132834);
nor I_2696 (I48448,I47988,I48431);
DFFARX1 I_2697 (I48448,I2595,I47928,I47893,);
and I_2698 (I47908,I48061,I132828);
not I_2699 (I48520,I2602);
DFFARX1 I_2700 (I295501,I2595,I48520,I48546,);
DFFARX1 I_2701 (I48546,I2595,I48520,I48563,);
not I_2702 (I48512,I48563);
not I_2703 (I48585,I48546);
DFFARX1 I_2704 (I295510,I2595,I48520,I48611,);
not I_2705 (I48619,I48611);
and I_2706 (I48636,I48585,I295504);
not I_2707 (I48653,I295498);
nand I_2708 (I48670,I48653,I295504);
not I_2709 (I48687,I295513);
nor I_2710 (I48704,I48687,I295501);
nand I_2711 (I48721,I48704,I295507);
nor I_2712 (I48738,I48721,I48670);
DFFARX1 I_2713 (I48738,I2595,I48520,I48488,);
not I_2714 (I48769,I48721);
not I_2715 (I48786,I295501);
nand I_2716 (I48803,I48786,I295504);
nor I_2717 (I48820,I295501,I295498);
nand I_2718 (I48500,I48636,I48820);
nand I_2719 (I48494,I48585,I295501);
nand I_2720 (I48865,I48687,I295504);
DFFARX1 I_2721 (I48865,I2595,I48520,I48509,);
DFFARX1 I_2722 (I48865,I2595,I48520,I48503,);
not I_2723 (I48910,I295504);
nor I_2724 (I48927,I48910,I295519);
and I_2725 (I48944,I48927,I295516);
or I_2726 (I48961,I48944,I295498);
DFFARX1 I_2727 (I48961,I2595,I48520,I48987,);
nand I_2728 (I48995,I48987,I48653);
nor I_2729 (I48497,I48995,I48803);
nor I_2730 (I48491,I48987,I48619);
DFFARX1 I_2731 (I48987,I2595,I48520,I49049,);
not I_2732 (I49057,I49049);
nor I_2733 (I48506,I49057,I48769);
not I_2734 (I49115,I2602);
DFFARX1 I_2735 (I315422,I2595,I49115,I49141,);
DFFARX1 I_2736 (I49141,I2595,I49115,I49158,);
not I_2737 (I49107,I49158);
not I_2738 (I49180,I49141);
DFFARX1 I_2739 (I315422,I2595,I49115,I49206,);
not I_2740 (I49214,I49206);
and I_2741 (I49231,I49180,I315425);
not I_2742 (I49248,I315437);
nand I_2743 (I49265,I49248,I315425);
not I_2744 (I49282,I315443);
nor I_2745 (I49299,I49282,I315434);
nand I_2746 (I49316,I49299,I315440);
nor I_2747 (I49333,I49316,I49265);
DFFARX1 I_2748 (I49333,I2595,I49115,I49083,);
not I_2749 (I49364,I49316);
not I_2750 (I49381,I315434);
nand I_2751 (I49398,I49381,I315425);
nor I_2752 (I49415,I315434,I315437);
nand I_2753 (I49095,I49231,I49415);
nand I_2754 (I49089,I49180,I315434);
nand I_2755 (I49460,I49282,I315431);
DFFARX1 I_2756 (I49460,I2595,I49115,I49104,);
DFFARX1 I_2757 (I49460,I2595,I49115,I49098,);
not I_2758 (I49505,I315431);
nor I_2759 (I49522,I49505,I315428);
and I_2760 (I49539,I49522,I315446);
or I_2761 (I49556,I49539,I315425);
DFFARX1 I_2762 (I49556,I2595,I49115,I49582,);
nand I_2763 (I49590,I49582,I49248);
nor I_2764 (I49092,I49590,I49398);
nor I_2765 (I49086,I49582,I49214);
DFFARX1 I_2766 (I49582,I2595,I49115,I49644,);
not I_2767 (I49652,I49644);
nor I_2768 (I49101,I49652,I49364);
not I_2769 (I49710,I2602);
DFFARX1 I_2770 (I176105,I2595,I49710,I49736,);
DFFARX1 I_2771 (I49736,I2595,I49710,I49753,);
not I_2772 (I49702,I49753);
not I_2773 (I49775,I49736);
DFFARX1 I_2774 (I176096,I2595,I49710,I49801,);
not I_2775 (I49809,I49801);
and I_2776 (I49826,I49775,I176114);
not I_2777 (I49843,I176111);
nand I_2778 (I49860,I49843,I176114);
not I_2779 (I49877,I176090);
nor I_2780 (I49894,I49877,I176093);
nand I_2781 (I49911,I49894,I176102);
nor I_2782 (I49928,I49911,I49860);
DFFARX1 I_2783 (I49928,I2595,I49710,I49678,);
not I_2784 (I49959,I49911);
not I_2785 (I49976,I176093);
nand I_2786 (I49993,I49976,I176114);
nor I_2787 (I50010,I176093,I176111);
nand I_2788 (I49690,I49826,I50010);
nand I_2789 (I49684,I49775,I176093);
nand I_2790 (I50055,I49877,I176108);
DFFARX1 I_2791 (I50055,I2595,I49710,I49699,);
DFFARX1 I_2792 (I50055,I2595,I49710,I49693,);
not I_2793 (I50100,I176108);
nor I_2794 (I50117,I50100,I176090);
and I_2795 (I50134,I50117,I176099);
or I_2796 (I50151,I50134,I176093);
DFFARX1 I_2797 (I50151,I2595,I49710,I50177,);
nand I_2798 (I50185,I50177,I49843);
nor I_2799 (I49687,I50185,I49993);
nor I_2800 (I49681,I50177,I49809);
DFFARX1 I_2801 (I50177,I2595,I49710,I50239,);
not I_2802 (I50247,I50239);
nor I_2803 (I49696,I50247,I49959);
not I_2804 (I50305,I2602);
DFFARX1 I_2805 (I218874,I2595,I50305,I50331,);
DFFARX1 I_2806 (I50331,I2595,I50305,I50348,);
not I_2807 (I50297,I50348);
not I_2808 (I50370,I50331);
DFFARX1 I_2809 (I218871,I2595,I50305,I50396,);
not I_2810 (I50404,I50396);
and I_2811 (I50421,I50370,I218877);
not I_2812 (I50438,I218862);
nand I_2813 (I50455,I50438,I218877);
not I_2814 (I50472,I218865);
nor I_2815 (I50489,I50472,I218886);
nand I_2816 (I50506,I50489,I218883);
nor I_2817 (I50523,I50506,I50455);
DFFARX1 I_2818 (I50523,I2595,I50305,I50273,);
not I_2819 (I50554,I50506);
not I_2820 (I50571,I218886);
nand I_2821 (I50588,I50571,I218877);
nor I_2822 (I50605,I218886,I218862);
nand I_2823 (I50285,I50421,I50605);
nand I_2824 (I50279,I50370,I218886);
nand I_2825 (I50650,I50472,I218862);
DFFARX1 I_2826 (I50650,I2595,I50305,I50294,);
DFFARX1 I_2827 (I50650,I2595,I50305,I50288,);
not I_2828 (I50695,I218862);
nor I_2829 (I50712,I50695,I218868);
and I_2830 (I50729,I50712,I218880);
or I_2831 (I50746,I50729,I218865);
DFFARX1 I_2832 (I50746,I2595,I50305,I50772,);
nand I_2833 (I50780,I50772,I50438);
nor I_2834 (I50282,I50780,I50588);
nor I_2835 (I50276,I50772,I50404);
DFFARX1 I_2836 (I50772,I2595,I50305,I50834,);
not I_2837 (I50842,I50834);
nor I_2838 (I50291,I50842,I50554);
not I_2839 (I50900,I2602);
DFFARX1 I_2840 (I181304,I2595,I50900,I50926,);
DFFARX1 I_2841 (I50926,I2595,I50900,I50943,);
not I_2842 (I50892,I50943);
not I_2843 (I50965,I50926);
DFFARX1 I_2844 (I181301,I2595,I50900,I50991,);
not I_2845 (I50999,I50991);
and I_2846 (I51016,I50965,I181307);
not I_2847 (I51033,I181292);
nand I_2848 (I51050,I51033,I181307);
not I_2849 (I51067,I181295);
nor I_2850 (I51084,I51067,I181316);
nand I_2851 (I51101,I51084,I181313);
nor I_2852 (I51118,I51101,I51050);
DFFARX1 I_2853 (I51118,I2595,I50900,I50868,);
not I_2854 (I51149,I51101);
not I_2855 (I51166,I181316);
nand I_2856 (I51183,I51166,I181307);
nor I_2857 (I51200,I181316,I181292);
nand I_2858 (I50880,I51016,I51200);
nand I_2859 (I50874,I50965,I181316);
nand I_2860 (I51245,I51067,I181292);
DFFARX1 I_2861 (I51245,I2595,I50900,I50889,);
DFFARX1 I_2862 (I51245,I2595,I50900,I50883,);
not I_2863 (I51290,I181292);
nor I_2864 (I51307,I51290,I181298);
and I_2865 (I51324,I51307,I181310);
or I_2866 (I51341,I51324,I181295);
DFFARX1 I_2867 (I51341,I2595,I50900,I51367,);
nand I_2868 (I51375,I51367,I51033);
nor I_2869 (I50877,I51375,I51183);
nor I_2870 (I50871,I51367,I50999);
DFFARX1 I_2871 (I51367,I2595,I50900,I51429,);
not I_2872 (I51437,I51429);
nor I_2873 (I50886,I51437,I51149);
not I_2874 (I51495,I2602);
DFFARX1 I_2875 (I179573,I2595,I51495,I51521,);
DFFARX1 I_2876 (I51521,I2595,I51495,I51538,);
not I_2877 (I51487,I51538);
not I_2878 (I51560,I51521);
DFFARX1 I_2879 (I179564,I2595,I51495,I51586,);
not I_2880 (I51594,I51586);
and I_2881 (I51611,I51560,I179582);
not I_2882 (I51628,I179579);
nand I_2883 (I51645,I51628,I179582);
not I_2884 (I51662,I179558);
nor I_2885 (I51679,I51662,I179561);
nand I_2886 (I51696,I51679,I179570);
nor I_2887 (I51713,I51696,I51645);
DFFARX1 I_2888 (I51713,I2595,I51495,I51463,);
not I_2889 (I51744,I51696);
not I_2890 (I51761,I179561);
nand I_2891 (I51778,I51761,I179582);
nor I_2892 (I51795,I179561,I179579);
nand I_2893 (I51475,I51611,I51795);
nand I_2894 (I51469,I51560,I179561);
nand I_2895 (I51840,I51662,I179576);
DFFARX1 I_2896 (I51840,I2595,I51495,I51484,);
DFFARX1 I_2897 (I51840,I2595,I51495,I51478,);
not I_2898 (I51885,I179576);
nor I_2899 (I51902,I51885,I179558);
and I_2900 (I51919,I51902,I179567);
or I_2901 (I51936,I51919,I179561);
DFFARX1 I_2902 (I51936,I2595,I51495,I51962,);
nand I_2903 (I51970,I51962,I51628);
nor I_2904 (I51472,I51970,I51778);
nor I_2905 (I51466,I51962,I51594);
DFFARX1 I_2906 (I51962,I2595,I51495,I52024,);
not I_2907 (I52032,I52024);
nor I_2908 (I51481,I52032,I51744);
not I_2909 (I52090,I2602);
DFFARX1 I_2910 (I211938,I2595,I52090,I52116,);
DFFARX1 I_2911 (I52116,I2595,I52090,I52133,);
not I_2912 (I52082,I52133);
not I_2913 (I52155,I52116);
DFFARX1 I_2914 (I211935,I2595,I52090,I52181,);
not I_2915 (I52189,I52181);
and I_2916 (I52206,I52155,I211941);
not I_2917 (I52223,I211926);
nand I_2918 (I52240,I52223,I211941);
not I_2919 (I52257,I211929);
nor I_2920 (I52274,I52257,I211950);
nand I_2921 (I52291,I52274,I211947);
nor I_2922 (I52308,I52291,I52240);
DFFARX1 I_2923 (I52308,I2595,I52090,I52058,);
not I_2924 (I52339,I52291);
not I_2925 (I52356,I211950);
nand I_2926 (I52373,I52356,I211941);
nor I_2927 (I52390,I211950,I211926);
nand I_2928 (I52070,I52206,I52390);
nand I_2929 (I52064,I52155,I211950);
nand I_2930 (I52435,I52257,I211926);
DFFARX1 I_2931 (I52435,I2595,I52090,I52079,);
DFFARX1 I_2932 (I52435,I2595,I52090,I52073,);
not I_2933 (I52480,I211926);
nor I_2934 (I52497,I52480,I211932);
and I_2935 (I52514,I52497,I211944);
or I_2936 (I52531,I52514,I211929);
DFFARX1 I_2937 (I52531,I2595,I52090,I52557,);
nand I_2938 (I52565,I52557,I52223);
nor I_2939 (I52067,I52565,I52373);
nor I_2940 (I52061,I52557,I52189);
DFFARX1 I_2941 (I52557,I2595,I52090,I52619,);
not I_2942 (I52627,I52619);
nor I_2943 (I52076,I52627,I52339);
not I_2944 (I52685,I2602);
DFFARX1 I_2945 (I200378,I2595,I52685,I52711,);
DFFARX1 I_2946 (I52711,I2595,I52685,I52728,);
not I_2947 (I52677,I52728);
not I_2948 (I52750,I52711);
DFFARX1 I_2949 (I200375,I2595,I52685,I52776,);
not I_2950 (I52784,I52776);
and I_2951 (I52801,I52750,I200381);
not I_2952 (I52818,I200366);
nand I_2953 (I52835,I52818,I200381);
not I_2954 (I52852,I200369);
nor I_2955 (I52869,I52852,I200390);
nand I_2956 (I52886,I52869,I200387);
nor I_2957 (I52903,I52886,I52835);
DFFARX1 I_2958 (I52903,I2595,I52685,I52653,);
not I_2959 (I52934,I52886);
not I_2960 (I52951,I200390);
nand I_2961 (I52968,I52951,I200381);
nor I_2962 (I52985,I200390,I200366);
nand I_2963 (I52665,I52801,I52985);
nand I_2964 (I52659,I52750,I200390);
nand I_2965 (I53030,I52852,I200366);
DFFARX1 I_2966 (I53030,I2595,I52685,I52674,);
DFFARX1 I_2967 (I53030,I2595,I52685,I52668,);
not I_2968 (I53075,I200366);
nor I_2969 (I53092,I53075,I200372);
and I_2970 (I53109,I53092,I200384);
or I_2971 (I53126,I53109,I200369);
DFFARX1 I_2972 (I53126,I2595,I52685,I53152,);
nand I_2973 (I53160,I53152,I52818);
nor I_2974 (I52662,I53160,I52968);
nor I_2975 (I52656,I53152,I52784);
DFFARX1 I_2976 (I53152,I2595,I52685,I53214,);
not I_2977 (I53222,I53214);
nor I_2978 (I52671,I53222,I52934);
not I_2979 (I53280,I2602);
DFFARX1 I_2980 (I312532,I2595,I53280,I53306,);
DFFARX1 I_2981 (I53306,I2595,I53280,I53323,);
not I_2982 (I53272,I53323);
not I_2983 (I53345,I53306);
DFFARX1 I_2984 (I312532,I2595,I53280,I53371,);
not I_2985 (I53379,I53371);
and I_2986 (I53396,I53345,I312535);
not I_2987 (I53413,I312547);
nand I_2988 (I53430,I53413,I312535);
not I_2989 (I53447,I312553);
nor I_2990 (I53464,I53447,I312544);
nand I_2991 (I53481,I53464,I312550);
nor I_2992 (I53498,I53481,I53430);
DFFARX1 I_2993 (I53498,I2595,I53280,I53248,);
not I_2994 (I53529,I53481);
not I_2995 (I53546,I312544);
nand I_2996 (I53563,I53546,I312535);
nor I_2997 (I53580,I312544,I312547);
nand I_2998 (I53260,I53396,I53580);
nand I_2999 (I53254,I53345,I312544);
nand I_3000 (I53625,I53447,I312541);
DFFARX1 I_3001 (I53625,I2595,I53280,I53269,);
DFFARX1 I_3002 (I53625,I2595,I53280,I53263,);
not I_3003 (I53670,I312541);
nor I_3004 (I53687,I53670,I312538);
and I_3005 (I53704,I53687,I312556);
or I_3006 (I53721,I53704,I312535);
DFFARX1 I_3007 (I53721,I2595,I53280,I53747,);
nand I_3008 (I53755,I53747,I53413);
nor I_3009 (I53257,I53755,I53563);
nor I_3010 (I53251,I53747,I53379);
DFFARX1 I_3011 (I53747,I2595,I53280,I53809,);
not I_3012 (I53817,I53809);
nor I_3013 (I53266,I53817,I53529);
not I_3014 (I53875,I2602);
DFFARX1 I_3015 (I101698,I2595,I53875,I53901,);
DFFARX1 I_3016 (I53901,I2595,I53875,I53918,);
not I_3017 (I53867,I53918);
not I_3018 (I53940,I53901);
DFFARX1 I_3019 (I101713,I2595,I53875,I53966,);
not I_3020 (I53974,I53966);
and I_3021 (I53991,I53940,I101710);
not I_3022 (I54008,I101698);
nand I_3023 (I54025,I54008,I101710);
not I_3024 (I54042,I101707);
nor I_3025 (I54059,I54042,I101722);
nand I_3026 (I54076,I54059,I101719);
nor I_3027 (I54093,I54076,I54025);
DFFARX1 I_3028 (I54093,I2595,I53875,I53843,);
not I_3029 (I54124,I54076);
not I_3030 (I54141,I101722);
nand I_3031 (I54158,I54141,I101710);
nor I_3032 (I54175,I101722,I101698);
nand I_3033 (I53855,I53991,I54175);
nand I_3034 (I53849,I53940,I101722);
nand I_3035 (I54220,I54042,I101716);
DFFARX1 I_3036 (I54220,I2595,I53875,I53864,);
DFFARX1 I_3037 (I54220,I2595,I53875,I53858,);
not I_3038 (I54265,I101716);
nor I_3039 (I54282,I54265,I101704);
and I_3040 (I54299,I54282,I101725);
or I_3041 (I54316,I54299,I101701);
DFFARX1 I_3042 (I54316,I2595,I53875,I54342,);
nand I_3043 (I54350,I54342,I54008);
nor I_3044 (I53852,I54350,I54158);
nor I_3045 (I53846,I54342,I53974);
DFFARX1 I_3046 (I54342,I2595,I53875,I54404,);
not I_3047 (I54412,I54404);
nor I_3048 (I53861,I54412,I54124);
not I_3049 (I54470,I2602);
DFFARX1 I_3050 (I241971,I2595,I54470,I54496,);
DFFARX1 I_3051 (I54496,I2595,I54470,I54513,);
not I_3052 (I54462,I54513);
not I_3053 (I54535,I54496);
DFFARX1 I_3054 (I241965,I2595,I54470,I54561,);
not I_3055 (I54569,I54561);
and I_3056 (I54586,I54535,I241983);
not I_3057 (I54603,I241971);
nand I_3058 (I54620,I54603,I241983);
not I_3059 (I54637,I241965);
nor I_3060 (I54654,I54637,I241977);
nand I_3061 (I54671,I54654,I241968);
nor I_3062 (I54688,I54671,I54620);
DFFARX1 I_3063 (I54688,I2595,I54470,I54438,);
not I_3064 (I54719,I54671);
not I_3065 (I54736,I241977);
nand I_3066 (I54753,I54736,I241983);
nor I_3067 (I54770,I241977,I241971);
nand I_3068 (I54450,I54586,I54770);
nand I_3069 (I54444,I54535,I241977);
nand I_3070 (I54815,I54637,I241980);
DFFARX1 I_3071 (I54815,I2595,I54470,I54459,);
DFFARX1 I_3072 (I54815,I2595,I54470,I54453,);
not I_3073 (I54860,I241980);
nor I_3074 (I54877,I54860,I241986);
and I_3075 (I54894,I54877,I241968);
or I_3076 (I54911,I54894,I241974);
DFFARX1 I_3077 (I54911,I2595,I54470,I54937,);
nand I_3078 (I54945,I54937,I54603);
nor I_3079 (I54447,I54945,I54753);
nor I_3080 (I54441,I54937,I54569);
DFFARX1 I_3081 (I54937,I2595,I54470,I54999,);
not I_3082 (I55007,I54999);
nor I_3083 (I54456,I55007,I54719);
not I_3084 (I55065,I2602);
DFFARX1 I_3085 (I239863,I2595,I55065,I55091,);
DFFARX1 I_3086 (I55091,I2595,I55065,I55108,);
not I_3087 (I55057,I55108);
not I_3088 (I55130,I55091);
DFFARX1 I_3089 (I239857,I2595,I55065,I55156,);
not I_3090 (I55164,I55156);
and I_3091 (I55181,I55130,I239875);
not I_3092 (I55198,I239863);
nand I_3093 (I55215,I55198,I239875);
not I_3094 (I55232,I239857);
nor I_3095 (I55249,I55232,I239869);
nand I_3096 (I55266,I55249,I239860);
nor I_3097 (I55283,I55266,I55215);
DFFARX1 I_3098 (I55283,I2595,I55065,I55033,);
not I_3099 (I55314,I55266);
not I_3100 (I55331,I239869);
nand I_3101 (I55348,I55331,I239875);
nor I_3102 (I55365,I239869,I239863);
nand I_3103 (I55045,I55181,I55365);
nand I_3104 (I55039,I55130,I239869);
nand I_3105 (I55410,I55232,I239872);
DFFARX1 I_3106 (I55410,I2595,I55065,I55054,);
DFFARX1 I_3107 (I55410,I2595,I55065,I55048,);
not I_3108 (I55455,I239872);
nor I_3109 (I55472,I55455,I239878);
and I_3110 (I55489,I55472,I239860);
or I_3111 (I55506,I55489,I239866);
DFFARX1 I_3112 (I55506,I2595,I55065,I55532,);
nand I_3113 (I55540,I55532,I55198);
nor I_3114 (I55042,I55540,I55348);
nor I_3115 (I55036,I55532,I55164);
DFFARX1 I_3116 (I55532,I2595,I55065,I55594,);
not I_3117 (I55602,I55594);
nor I_3118 (I55051,I55602,I55314);
not I_3119 (I55660,I2602);
DFFARX1 I_3120 (I151112,I2595,I55660,I55686,);
DFFARX1 I_3121 (I55686,I2595,I55660,I55703,);
not I_3122 (I55652,I55703);
not I_3123 (I55725,I55686);
DFFARX1 I_3124 (I151106,I2595,I55660,I55751,);
not I_3125 (I55759,I55751);
and I_3126 (I55776,I55725,I151121);
not I_3127 (I55793,I151118);
nand I_3128 (I55810,I55793,I151121);
not I_3129 (I55827,I151109);
nor I_3130 (I55844,I55827,I151100);
nand I_3131 (I55861,I55844,I151103);
nor I_3132 (I55878,I55861,I55810);
DFFARX1 I_3133 (I55878,I2595,I55660,I55628,);
not I_3134 (I55909,I55861);
not I_3135 (I55926,I151100);
nand I_3136 (I55943,I55926,I151121);
nor I_3137 (I55960,I151100,I151118);
nand I_3138 (I55640,I55776,I55960);
nand I_3139 (I55634,I55725,I151100);
nand I_3140 (I56005,I55827,I151124);
DFFARX1 I_3141 (I56005,I2595,I55660,I55649,);
DFFARX1 I_3142 (I56005,I2595,I55660,I55643,);
not I_3143 (I56050,I151124);
nor I_3144 (I56067,I56050,I151115);
and I_3145 (I56084,I56067,I151100);
or I_3146 (I56101,I56084,I151103);
DFFARX1 I_3147 (I56101,I2595,I55660,I56127,);
nand I_3148 (I56135,I56127,I55793);
nor I_3149 (I55637,I56135,I55943);
nor I_3150 (I55631,I56127,I55759);
DFFARX1 I_3151 (I56127,I2595,I55660,I56189,);
not I_3152 (I56197,I56189);
nor I_3153 (I55646,I56197,I55909);
not I_3154 (I56255,I2602);
DFFARX1 I_3155 (I18201,I2595,I56255,I56281,);
DFFARX1 I_3156 (I56281,I2595,I56255,I56298,);
not I_3157 (I56247,I56298);
not I_3158 (I56320,I56281);
DFFARX1 I_3159 (I18177,I2595,I56255,I56346,);
not I_3160 (I56354,I56346);
and I_3161 (I56371,I56320,I18192);
not I_3162 (I56388,I18180);
nand I_3163 (I56405,I56388,I18192);
not I_3164 (I56422,I18183);
nor I_3165 (I56439,I56422,I18195);
nand I_3166 (I56456,I56439,I18186);
nor I_3167 (I56473,I56456,I56405);
DFFARX1 I_3168 (I56473,I2595,I56255,I56223,);
not I_3169 (I56504,I56456);
not I_3170 (I56521,I18195);
nand I_3171 (I56538,I56521,I18192);
nor I_3172 (I56555,I18195,I18180);
nand I_3173 (I56235,I56371,I56555);
nand I_3174 (I56229,I56320,I18195);
nand I_3175 (I56600,I56422,I18189);
DFFARX1 I_3176 (I56600,I2595,I56255,I56244,);
DFFARX1 I_3177 (I56600,I2595,I56255,I56238,);
not I_3178 (I56645,I18189);
nor I_3179 (I56662,I56645,I18180);
and I_3180 (I56679,I56662,I18177);
or I_3181 (I56696,I56679,I18198);
DFFARX1 I_3182 (I56696,I2595,I56255,I56722,);
nand I_3183 (I56730,I56722,I56388);
nor I_3184 (I56232,I56730,I56538);
nor I_3185 (I56226,I56722,I56354);
DFFARX1 I_3186 (I56722,I2595,I56255,I56784,);
not I_3187 (I56792,I56784);
nor I_3188 (I56241,I56792,I56504);
not I_3189 (I56850,I2602);
DFFARX1 I_3190 (I177839,I2595,I56850,I56876,);
DFFARX1 I_3191 (I56876,I2595,I56850,I56893,);
not I_3192 (I56842,I56893);
not I_3193 (I56915,I56876);
DFFARX1 I_3194 (I177830,I2595,I56850,I56941,);
not I_3195 (I56949,I56941);
and I_3196 (I56966,I56915,I177848);
not I_3197 (I56983,I177845);
nand I_3198 (I57000,I56983,I177848);
not I_3199 (I57017,I177824);
nor I_3200 (I57034,I57017,I177827);
nand I_3201 (I57051,I57034,I177836);
nor I_3202 (I57068,I57051,I57000);
DFFARX1 I_3203 (I57068,I2595,I56850,I56818,);
not I_3204 (I57099,I57051);
not I_3205 (I57116,I177827);
nand I_3206 (I57133,I57116,I177848);
nor I_3207 (I57150,I177827,I177845);
nand I_3208 (I56830,I56966,I57150);
nand I_3209 (I56824,I56915,I177827);
nand I_3210 (I57195,I57017,I177842);
DFFARX1 I_3211 (I57195,I2595,I56850,I56839,);
DFFARX1 I_3212 (I57195,I2595,I56850,I56833,);
not I_3213 (I57240,I177842);
nor I_3214 (I57257,I57240,I177824);
and I_3215 (I57274,I57257,I177833);
or I_3216 (I57291,I57274,I177827);
DFFARX1 I_3217 (I57291,I2595,I56850,I57317,);
nand I_3218 (I57325,I57317,I56983);
nor I_3219 (I56827,I57325,I57133);
nor I_3220 (I56821,I57317,I56949);
DFFARX1 I_3221 (I57317,I2595,I56850,I57379,);
not I_3222 (I57387,I57379);
nor I_3223 (I56836,I57387,I57099);
not I_3224 (I57445,I2602);
DFFARX1 I_3225 (I208470,I2595,I57445,I57471,);
DFFARX1 I_3226 (I57471,I2595,I57445,I57488,);
not I_3227 (I57437,I57488);
not I_3228 (I57510,I57471);
DFFARX1 I_3229 (I208467,I2595,I57445,I57536,);
not I_3230 (I57544,I57536);
and I_3231 (I57561,I57510,I208473);
not I_3232 (I57578,I208458);
nand I_3233 (I57595,I57578,I208473);
not I_3234 (I57612,I208461);
nor I_3235 (I57629,I57612,I208482);
nand I_3236 (I57646,I57629,I208479);
nor I_3237 (I57663,I57646,I57595);
DFFARX1 I_3238 (I57663,I2595,I57445,I57413,);
not I_3239 (I57694,I57646);
not I_3240 (I57711,I208482);
nand I_3241 (I57728,I57711,I208473);
nor I_3242 (I57745,I208482,I208458);
nand I_3243 (I57425,I57561,I57745);
nand I_3244 (I57419,I57510,I208482);
nand I_3245 (I57790,I57612,I208458);
DFFARX1 I_3246 (I57790,I2595,I57445,I57434,);
DFFARX1 I_3247 (I57790,I2595,I57445,I57428,);
not I_3248 (I57835,I208458);
nor I_3249 (I57852,I57835,I208464);
and I_3250 (I57869,I57852,I208476);
or I_3251 (I57886,I57869,I208461);
DFFARX1 I_3252 (I57886,I2595,I57445,I57912,);
nand I_3253 (I57920,I57912,I57578);
nor I_3254 (I57422,I57920,I57728);
nor I_3255 (I57416,I57912,I57544);
DFFARX1 I_3256 (I57912,I2595,I57445,I57974,);
not I_3257 (I57982,I57974);
nor I_3258 (I57431,I57982,I57694);
not I_3259 (I58040,I2602);
DFFARX1 I_3260 (I122513,I2595,I58040,I58066,);
DFFARX1 I_3261 (I58066,I2595,I58040,I58083,);
not I_3262 (I58032,I58083);
not I_3263 (I58105,I58066);
DFFARX1 I_3264 (I122501,I2595,I58040,I58131,);
not I_3265 (I58139,I58131);
and I_3266 (I58156,I58105,I122510);
not I_3267 (I58173,I122507);
nand I_3268 (I58190,I58173,I122510);
not I_3269 (I58207,I122498);
nor I_3270 (I58224,I58207,I122504);
nand I_3271 (I58241,I58224,I122489);
nor I_3272 (I58258,I58241,I58190);
DFFARX1 I_3273 (I58258,I2595,I58040,I58008,);
not I_3274 (I58289,I58241);
not I_3275 (I58306,I122504);
nand I_3276 (I58323,I58306,I122510);
nor I_3277 (I58340,I122504,I122507);
nand I_3278 (I58020,I58156,I58340);
nand I_3279 (I58014,I58105,I122504);
nand I_3280 (I58385,I58207,I122489);
DFFARX1 I_3281 (I58385,I2595,I58040,I58029,);
DFFARX1 I_3282 (I58385,I2595,I58040,I58023,);
not I_3283 (I58430,I122489);
nor I_3284 (I58447,I58430,I122495);
and I_3285 (I58464,I58447,I122492);
or I_3286 (I58481,I58464,I122516);
DFFARX1 I_3287 (I58481,I2595,I58040,I58507,);
nand I_3288 (I58515,I58507,I58173);
nor I_3289 (I58017,I58515,I58323);
nor I_3290 (I58011,I58507,I58139);
DFFARX1 I_3291 (I58507,I2595,I58040,I58569,);
not I_3292 (I58577,I58569);
nor I_3293 (I58026,I58577,I58289);
not I_3294 (I58635,I2602);
DFFARX1 I_3295 (I111711,I2595,I58635,I58661,);
DFFARX1 I_3296 (I58661,I2595,I58635,I58678,);
not I_3297 (I58627,I58678);
not I_3298 (I58700,I58661);
DFFARX1 I_3299 (I111726,I2595,I58635,I58726,);
not I_3300 (I58734,I58726);
and I_3301 (I58751,I58700,I111723);
not I_3302 (I58768,I111711);
nand I_3303 (I58785,I58768,I111723);
not I_3304 (I58802,I111720);
nor I_3305 (I58819,I58802,I111735);
nand I_3306 (I58836,I58819,I111732);
nor I_3307 (I58853,I58836,I58785);
DFFARX1 I_3308 (I58853,I2595,I58635,I58603,);
not I_3309 (I58884,I58836);
not I_3310 (I58901,I111735);
nand I_3311 (I58918,I58901,I111723);
nor I_3312 (I58935,I111735,I111711);
nand I_3313 (I58615,I58751,I58935);
nand I_3314 (I58609,I58700,I111735);
nand I_3315 (I58980,I58802,I111729);
DFFARX1 I_3316 (I58980,I2595,I58635,I58624,);
DFFARX1 I_3317 (I58980,I2595,I58635,I58618,);
not I_3318 (I59025,I111729);
nor I_3319 (I59042,I59025,I111717);
and I_3320 (I59059,I59042,I111738);
or I_3321 (I59076,I59059,I111714);
DFFARX1 I_3322 (I59076,I2595,I58635,I59102,);
nand I_3323 (I59110,I59102,I58768);
nor I_3324 (I58612,I59110,I58918);
nor I_3325 (I58606,I59102,I58734);
DFFARX1 I_3326 (I59102,I2595,I58635,I59164,);
not I_3327 (I59172,I59164);
nor I_3328 (I58621,I59172,I58884);
not I_3329 (I59230,I2602);
DFFARX1 I_3330 (I357347,I2595,I59230,I59256,);
DFFARX1 I_3331 (I59256,I2595,I59230,I59273,);
not I_3332 (I59222,I59273);
not I_3333 (I59295,I59256);
DFFARX1 I_3334 (I357359,I2595,I59230,I59321,);
not I_3335 (I59329,I59321);
and I_3336 (I59346,I59295,I357353);
not I_3337 (I59363,I357365);
nand I_3338 (I59380,I59363,I357353);
not I_3339 (I59397,I357350);
nor I_3340 (I59414,I59397,I357362);
nand I_3341 (I59431,I59414,I357344);
nor I_3342 (I59448,I59431,I59380);
DFFARX1 I_3343 (I59448,I2595,I59230,I59198,);
not I_3344 (I59479,I59431);
not I_3345 (I59496,I357362);
nand I_3346 (I59513,I59496,I357353);
nor I_3347 (I59530,I357362,I357365);
nand I_3348 (I59210,I59346,I59530);
nand I_3349 (I59204,I59295,I357362);
nand I_3350 (I59575,I59397,I357356);
DFFARX1 I_3351 (I59575,I2595,I59230,I59219,);
DFFARX1 I_3352 (I59575,I2595,I59230,I59213,);
not I_3353 (I59620,I357356);
nor I_3354 (I59637,I59620,I357347);
and I_3355 (I59654,I59637,I357344);
or I_3356 (I59671,I59654,I357368);
DFFARX1 I_3357 (I59671,I2595,I59230,I59697,);
nand I_3358 (I59705,I59697,I59363);
nor I_3359 (I59207,I59705,I59513);
nor I_3360 (I59201,I59697,I59329);
DFFARX1 I_3361 (I59697,I2595,I59230,I59759,);
not I_3362 (I59767,I59759);
nor I_3363 (I59216,I59767,I59479);
not I_3364 (I59825,I2602);
DFFARX1 I_3365 (I305596,I2595,I59825,I59851,);
DFFARX1 I_3366 (I59851,I2595,I59825,I59868,);
not I_3367 (I59817,I59868);
not I_3368 (I59890,I59851);
DFFARX1 I_3369 (I305596,I2595,I59825,I59916,);
not I_3370 (I59924,I59916);
and I_3371 (I59941,I59890,I305599);
not I_3372 (I59958,I305611);
nand I_3373 (I59975,I59958,I305599);
not I_3374 (I59992,I305617);
nor I_3375 (I60009,I59992,I305608);
nand I_3376 (I60026,I60009,I305614);
nor I_3377 (I60043,I60026,I59975);
DFFARX1 I_3378 (I60043,I2595,I59825,I59793,);
not I_3379 (I60074,I60026);
not I_3380 (I60091,I305608);
nand I_3381 (I60108,I60091,I305599);
nor I_3382 (I60125,I305608,I305611);
nand I_3383 (I59805,I59941,I60125);
nand I_3384 (I59799,I59890,I305608);
nand I_3385 (I60170,I59992,I305605);
DFFARX1 I_3386 (I60170,I2595,I59825,I59814,);
DFFARX1 I_3387 (I60170,I2595,I59825,I59808,);
not I_3388 (I60215,I305605);
nor I_3389 (I60232,I60215,I305602);
and I_3390 (I60249,I60232,I305620);
or I_3391 (I60266,I60249,I305599);
DFFARX1 I_3392 (I60266,I2595,I59825,I60292,);
nand I_3393 (I60300,I60292,I59958);
nor I_3394 (I59802,I60300,I60108);
nor I_3395 (I59796,I60292,I59924);
DFFARX1 I_3396 (I60292,I2595,I59825,I60354,);
not I_3397 (I60362,I60354);
nor I_3398 (I59811,I60362,I60074);
not I_3399 (I60420,I2602);
DFFARX1 I_3400 (I365439,I2595,I60420,I60446,);
DFFARX1 I_3401 (I60446,I2595,I60420,I60463,);
not I_3402 (I60412,I60463);
not I_3403 (I60485,I60446);
DFFARX1 I_3404 (I365451,I2595,I60420,I60511,);
not I_3405 (I60519,I60511);
and I_3406 (I60536,I60485,I365445);
not I_3407 (I60553,I365457);
nand I_3408 (I60570,I60553,I365445);
not I_3409 (I60587,I365442);
nor I_3410 (I60604,I60587,I365454);
nand I_3411 (I60621,I60604,I365436);
nor I_3412 (I60638,I60621,I60570);
DFFARX1 I_3413 (I60638,I2595,I60420,I60388,);
not I_3414 (I60669,I60621);
not I_3415 (I60686,I365454);
nand I_3416 (I60703,I60686,I365445);
nor I_3417 (I60720,I365454,I365457);
nand I_3418 (I60400,I60536,I60720);
nand I_3419 (I60394,I60485,I365454);
nand I_3420 (I60765,I60587,I365448);
DFFARX1 I_3421 (I60765,I2595,I60420,I60409,);
DFFARX1 I_3422 (I60765,I2595,I60420,I60403,);
not I_3423 (I60810,I365448);
nor I_3424 (I60827,I60810,I365439);
and I_3425 (I60844,I60827,I365436);
or I_3426 (I60861,I60844,I365460);
DFFARX1 I_3427 (I60861,I2595,I60420,I60887,);
nand I_3428 (I60895,I60887,I60553);
nor I_3429 (I60397,I60895,I60703);
nor I_3430 (I60391,I60887,I60519);
DFFARX1 I_3431 (I60887,I2595,I60420,I60949,);
not I_3432 (I60957,I60949);
nor I_3433 (I60406,I60957,I60669);
not I_3434 (I61015,I2602);
DFFARX1 I_3435 (I114346,I2595,I61015,I61041,);
DFFARX1 I_3436 (I61041,I2595,I61015,I61058,);
not I_3437 (I61007,I61058);
not I_3438 (I61080,I61041);
DFFARX1 I_3439 (I114361,I2595,I61015,I61106,);
not I_3440 (I61114,I61106);
and I_3441 (I61131,I61080,I114358);
not I_3442 (I61148,I114346);
nand I_3443 (I61165,I61148,I114358);
not I_3444 (I61182,I114355);
nor I_3445 (I61199,I61182,I114370);
nand I_3446 (I61216,I61199,I114367);
nor I_3447 (I61233,I61216,I61165);
DFFARX1 I_3448 (I61233,I2595,I61015,I60983,);
not I_3449 (I61264,I61216);
not I_3450 (I61281,I114370);
nand I_3451 (I61298,I61281,I114358);
nor I_3452 (I61315,I114370,I114346);
nand I_3453 (I60995,I61131,I61315);
nand I_3454 (I60989,I61080,I114370);
nand I_3455 (I61360,I61182,I114364);
DFFARX1 I_3456 (I61360,I2595,I61015,I61004,);
DFFARX1 I_3457 (I61360,I2595,I61015,I60998,);
not I_3458 (I61405,I114364);
nor I_3459 (I61422,I61405,I114352);
and I_3460 (I61439,I61422,I114373);
or I_3461 (I61456,I61439,I114349);
DFFARX1 I_3462 (I61456,I2595,I61015,I61482,);
nand I_3463 (I61490,I61482,I61148);
nor I_3464 (I60992,I61490,I61298);
nor I_3465 (I60986,I61482,I61114);
DFFARX1 I_3466 (I61482,I2595,I61015,I61544,);
not I_3467 (I61552,I61544);
nor I_3468 (I61001,I61552,I61264);
not I_3469 (I61610,I2602);
DFFARX1 I_3470 (I282882,I2595,I61610,I61636,);
DFFARX1 I_3471 (I61636,I2595,I61610,I61653,);
not I_3472 (I61602,I61653);
not I_3473 (I61675,I61636);
DFFARX1 I_3474 (I282891,I2595,I61610,I61701,);
not I_3475 (I61709,I61701);
and I_3476 (I61726,I61675,I282879);
not I_3477 (I61743,I282870);
nand I_3478 (I61760,I61743,I282879);
not I_3479 (I61777,I282876);
nor I_3480 (I61794,I61777,I282894);
nand I_3481 (I61811,I61794,I282867);
nor I_3482 (I61828,I61811,I61760);
DFFARX1 I_3483 (I61828,I2595,I61610,I61578,);
not I_3484 (I61859,I61811);
not I_3485 (I61876,I282894);
nand I_3486 (I61893,I61876,I282879);
nor I_3487 (I61910,I282894,I282870);
nand I_3488 (I61590,I61726,I61910);
nand I_3489 (I61584,I61675,I282894);
nand I_3490 (I61955,I61777,I282873);
DFFARX1 I_3491 (I61955,I2595,I61610,I61599,);
DFFARX1 I_3492 (I61955,I2595,I61610,I61593,);
not I_3493 (I62000,I282873);
nor I_3494 (I62017,I62000,I282885);
and I_3495 (I62034,I62017,I282867);
or I_3496 (I62051,I62034,I282888);
DFFARX1 I_3497 (I62051,I2595,I61610,I62077,);
nand I_3498 (I62085,I62077,I61743);
nor I_3499 (I61587,I62085,I61893);
nor I_3500 (I61581,I62077,I61709);
DFFARX1 I_3501 (I62077,I2595,I61610,I62139,);
not I_3502 (I62147,I62139);
nor I_3503 (I61596,I62147,I61859);
not I_3504 (I62205,I2602);
DFFARX1 I_3505 (I106968,I2595,I62205,I62231,);
DFFARX1 I_3506 (I62231,I2595,I62205,I62248,);
not I_3507 (I62197,I62248);
not I_3508 (I62270,I62231);
DFFARX1 I_3509 (I106983,I2595,I62205,I62296,);
not I_3510 (I62304,I62296);
and I_3511 (I62321,I62270,I106980);
not I_3512 (I62338,I106968);
nand I_3513 (I62355,I62338,I106980);
not I_3514 (I62372,I106977);
nor I_3515 (I62389,I62372,I106992);
nand I_3516 (I62406,I62389,I106989);
nor I_3517 (I62423,I62406,I62355);
DFFARX1 I_3518 (I62423,I2595,I62205,I62173,);
not I_3519 (I62454,I62406);
not I_3520 (I62471,I106992);
nand I_3521 (I62488,I62471,I106980);
nor I_3522 (I62505,I106992,I106968);
nand I_3523 (I62185,I62321,I62505);
nand I_3524 (I62179,I62270,I106992);
nand I_3525 (I62550,I62372,I106986);
DFFARX1 I_3526 (I62550,I2595,I62205,I62194,);
DFFARX1 I_3527 (I62550,I2595,I62205,I62188,);
not I_3528 (I62595,I106986);
nor I_3529 (I62612,I62595,I106974);
and I_3530 (I62629,I62612,I106995);
or I_3531 (I62646,I62629,I106971);
DFFARX1 I_3532 (I62646,I2595,I62205,I62672,);
nand I_3533 (I62680,I62672,I62338);
nor I_3534 (I62182,I62680,I62488);
nor I_3535 (I62176,I62672,I62304);
DFFARX1 I_3536 (I62672,I2595,I62205,I62734,);
not I_3537 (I62742,I62734);
nor I_3538 (I62191,I62742,I62454);
not I_3539 (I62800,I2602);
DFFARX1 I_3540 (I155277,I2595,I62800,I62826,);
DFFARX1 I_3541 (I62826,I2595,I62800,I62843,);
not I_3542 (I62792,I62843);
not I_3543 (I62865,I62826);
DFFARX1 I_3544 (I155271,I2595,I62800,I62891,);
not I_3545 (I62899,I62891);
and I_3546 (I62916,I62865,I155286);
not I_3547 (I62933,I155283);
nand I_3548 (I62950,I62933,I155286);
not I_3549 (I62967,I155274);
nor I_3550 (I62984,I62967,I155265);
nand I_3551 (I63001,I62984,I155268);
nor I_3552 (I63018,I63001,I62950);
DFFARX1 I_3553 (I63018,I2595,I62800,I62768,);
not I_3554 (I63049,I63001);
not I_3555 (I63066,I155265);
nand I_3556 (I63083,I63066,I155286);
nor I_3557 (I63100,I155265,I155283);
nand I_3558 (I62780,I62916,I63100);
nand I_3559 (I62774,I62865,I155265);
nand I_3560 (I63145,I62967,I155289);
DFFARX1 I_3561 (I63145,I2595,I62800,I62789,);
DFFARX1 I_3562 (I63145,I2595,I62800,I62783,);
not I_3563 (I63190,I155289);
nor I_3564 (I63207,I63190,I155280);
and I_3565 (I63224,I63207,I155265);
or I_3566 (I63241,I63224,I155268);
DFFARX1 I_3567 (I63241,I2595,I62800,I63267,);
nand I_3568 (I63275,I63267,I62933);
nor I_3569 (I62777,I63275,I63083);
nor I_3570 (I62771,I63267,I62899);
DFFARX1 I_3571 (I63267,I2595,I62800,I63329,);
not I_3572 (I63337,I63329);
nor I_3573 (I62786,I63337,I63049);
not I_3574 (I63395,I2602);
DFFARX1 I_3575 (I10823,I2595,I63395,I63421,);
DFFARX1 I_3576 (I63421,I2595,I63395,I63438,);
not I_3577 (I63387,I63438);
not I_3578 (I63460,I63421);
DFFARX1 I_3579 (I10799,I2595,I63395,I63486,);
not I_3580 (I63494,I63486);
and I_3581 (I63511,I63460,I10814);
not I_3582 (I63528,I10802);
nand I_3583 (I63545,I63528,I10814);
not I_3584 (I63562,I10805);
nor I_3585 (I63579,I63562,I10817);
nand I_3586 (I63596,I63579,I10808);
nor I_3587 (I63613,I63596,I63545);
DFFARX1 I_3588 (I63613,I2595,I63395,I63363,);
not I_3589 (I63644,I63596);
not I_3590 (I63661,I10817);
nand I_3591 (I63678,I63661,I10814);
nor I_3592 (I63695,I10817,I10802);
nand I_3593 (I63375,I63511,I63695);
nand I_3594 (I63369,I63460,I10817);
nand I_3595 (I63740,I63562,I10811);
DFFARX1 I_3596 (I63740,I2595,I63395,I63384,);
DFFARX1 I_3597 (I63740,I2595,I63395,I63378,);
not I_3598 (I63785,I10811);
nor I_3599 (I63802,I63785,I10802);
and I_3600 (I63819,I63802,I10799);
or I_3601 (I63836,I63819,I10820);
DFFARX1 I_3602 (I63836,I2595,I63395,I63862,);
nand I_3603 (I63870,I63862,I63528);
nor I_3604 (I63372,I63870,I63678);
nor I_3605 (I63366,I63862,I63494);
DFFARX1 I_3606 (I63862,I2595,I63395,I63924,);
not I_3607 (I63932,I63924);
nor I_3608 (I63381,I63932,I63644);
not I_3609 (I63990,I2602);
DFFARX1 I_3610 (I345360,I2595,I63990,I64016,);
DFFARX1 I_3611 (I64016,I2595,I63990,I64033,);
not I_3612 (I63982,I64033);
not I_3613 (I64055,I64016);
DFFARX1 I_3614 (I345345,I2595,I63990,I64081,);
not I_3615 (I64089,I64081);
and I_3616 (I64106,I64055,I345363);
not I_3617 (I64123,I345345);
nand I_3618 (I64140,I64123,I345363);
not I_3619 (I64157,I345366);
nor I_3620 (I64174,I64157,I345357);
nand I_3621 (I64191,I64174,I345354);
nor I_3622 (I64208,I64191,I64140);
DFFARX1 I_3623 (I64208,I2595,I63990,I63958,);
not I_3624 (I64239,I64191);
not I_3625 (I64256,I345357);
nand I_3626 (I64273,I64256,I345363);
nor I_3627 (I64290,I345357,I345345);
nand I_3628 (I63970,I64106,I64290);
nand I_3629 (I63964,I64055,I345357);
nand I_3630 (I64335,I64157,I345351);
DFFARX1 I_3631 (I64335,I2595,I63990,I63979,);
DFFARX1 I_3632 (I64335,I2595,I63990,I63973,);
not I_3633 (I64380,I345351);
nor I_3634 (I64397,I64380,I345342);
and I_3635 (I64414,I64397,I345348);
or I_3636 (I64431,I64414,I345342);
DFFARX1 I_3637 (I64431,I2595,I63990,I64457,);
nand I_3638 (I64465,I64457,I64123);
nor I_3639 (I63967,I64465,I64273);
nor I_3640 (I63961,I64457,I64089);
DFFARX1 I_3641 (I64457,I2595,I63990,I64519,);
not I_3642 (I64527,I64519);
nor I_3643 (I63976,I64527,I64239);
not I_3644 (I64585,I2602);
DFFARX1 I_3645 (I306752,I2595,I64585,I64611,);
DFFARX1 I_3646 (I64611,I2595,I64585,I64628,);
not I_3647 (I64577,I64628);
not I_3648 (I64650,I64611);
DFFARX1 I_3649 (I306752,I2595,I64585,I64676,);
not I_3650 (I64684,I64676);
and I_3651 (I64701,I64650,I306755);
not I_3652 (I64718,I306767);
nand I_3653 (I64735,I64718,I306755);
not I_3654 (I64752,I306773);
nor I_3655 (I64769,I64752,I306764);
nand I_3656 (I64786,I64769,I306770);
nor I_3657 (I64803,I64786,I64735);
DFFARX1 I_3658 (I64803,I2595,I64585,I64553,);
not I_3659 (I64834,I64786);
not I_3660 (I64851,I306764);
nand I_3661 (I64868,I64851,I306755);
nor I_3662 (I64885,I306764,I306767);
nand I_3663 (I64565,I64701,I64885);
nand I_3664 (I64559,I64650,I306764);
nand I_3665 (I64930,I64752,I306761);
DFFARX1 I_3666 (I64930,I2595,I64585,I64574,);
DFFARX1 I_3667 (I64930,I2595,I64585,I64568,);
not I_3668 (I64975,I306761);
nor I_3669 (I64992,I64975,I306758);
and I_3670 (I65009,I64992,I306776);
or I_3671 (I65026,I65009,I306755);
DFFARX1 I_3672 (I65026,I2595,I64585,I65052,);
nand I_3673 (I65060,I65052,I64718);
nor I_3674 (I64562,I65060,I64868);
nor I_3675 (I64556,I65052,I64684);
DFFARX1 I_3676 (I65052,I2595,I64585,I65114,);
not I_3677 (I65122,I65114);
nor I_3678 (I64571,I65122,I64834);
not I_3679 (I65180,I2602);
DFFARX1 I_3680 (I193442,I2595,I65180,I65206,);
DFFARX1 I_3681 (I65206,I2595,I65180,I65223,);
not I_3682 (I65172,I65223);
not I_3683 (I65245,I65206);
DFFARX1 I_3684 (I193439,I2595,I65180,I65271,);
not I_3685 (I65279,I65271);
and I_3686 (I65296,I65245,I193445);
not I_3687 (I65313,I193430);
nand I_3688 (I65330,I65313,I193445);
not I_3689 (I65347,I193433);
nor I_3690 (I65364,I65347,I193454);
nand I_3691 (I65381,I65364,I193451);
nor I_3692 (I65398,I65381,I65330);
DFFARX1 I_3693 (I65398,I2595,I65180,I65148,);
not I_3694 (I65429,I65381);
not I_3695 (I65446,I193454);
nand I_3696 (I65463,I65446,I193445);
nor I_3697 (I65480,I193454,I193430);
nand I_3698 (I65160,I65296,I65480);
nand I_3699 (I65154,I65245,I193454);
nand I_3700 (I65525,I65347,I193430);
DFFARX1 I_3701 (I65525,I2595,I65180,I65169,);
DFFARX1 I_3702 (I65525,I2595,I65180,I65163,);
not I_3703 (I65570,I193430);
nor I_3704 (I65587,I65570,I193436);
and I_3705 (I65604,I65587,I193448);
or I_3706 (I65621,I65604,I193433);
DFFARX1 I_3707 (I65621,I2595,I65180,I65647,);
nand I_3708 (I65655,I65647,I65313);
nor I_3709 (I65157,I65655,I65463);
nor I_3710 (I65151,I65647,I65279);
DFFARX1 I_3711 (I65647,I2595,I65180,I65709,);
not I_3712 (I65717,I65709);
nor I_3713 (I65166,I65717,I65429);
not I_3714 (I65775,I2602);
DFFARX1 I_3715 (I255750,I2595,I65775,I65801,);
DFFARX1 I_3716 (I65801,I2595,I65775,I65818,);
not I_3717 (I65767,I65818);
not I_3718 (I65840,I65801);
DFFARX1 I_3719 (I255759,I2595,I65775,I65866,);
not I_3720 (I65874,I65866);
and I_3721 (I65891,I65840,I255747);
not I_3722 (I65908,I255738);
nand I_3723 (I65925,I65908,I255747);
not I_3724 (I65942,I255744);
nor I_3725 (I65959,I65942,I255762);
nand I_3726 (I65976,I65959,I255735);
nor I_3727 (I65993,I65976,I65925);
DFFARX1 I_3728 (I65993,I2595,I65775,I65743,);
not I_3729 (I66024,I65976);
not I_3730 (I66041,I255762);
nand I_3731 (I66058,I66041,I255747);
nor I_3732 (I66075,I255762,I255738);
nand I_3733 (I65755,I65891,I66075);
nand I_3734 (I65749,I65840,I255762);
nand I_3735 (I66120,I65942,I255741);
DFFARX1 I_3736 (I66120,I2595,I65775,I65764,);
DFFARX1 I_3737 (I66120,I2595,I65775,I65758,);
not I_3738 (I66165,I255741);
nor I_3739 (I66182,I66165,I255753);
and I_3740 (I66199,I66182,I255735);
or I_3741 (I66216,I66199,I255756);
DFFARX1 I_3742 (I66216,I2595,I65775,I66242,);
nand I_3743 (I66250,I66242,I65908);
nor I_3744 (I65752,I66250,I66058);
nor I_3745 (I65746,I66242,I65874);
DFFARX1 I_3746 (I66242,I2595,I65775,I66304,);
not I_3747 (I66312,I66304);
nor I_3748 (I65761,I66312,I66024);
not I_3749 (I66370,I2602);
DFFARX1 I_3750 (I149922,I2595,I66370,I66396,);
DFFARX1 I_3751 (I66396,I2595,I66370,I66413,);
not I_3752 (I66362,I66413);
not I_3753 (I66435,I66396);
DFFARX1 I_3754 (I149916,I2595,I66370,I66461,);
not I_3755 (I66469,I66461);
and I_3756 (I66486,I66435,I149931);
not I_3757 (I66503,I149928);
nand I_3758 (I66520,I66503,I149931);
not I_3759 (I66537,I149919);
nor I_3760 (I66554,I66537,I149910);
nand I_3761 (I66571,I66554,I149913);
nor I_3762 (I66588,I66571,I66520);
DFFARX1 I_3763 (I66588,I2595,I66370,I66338,);
not I_3764 (I66619,I66571);
not I_3765 (I66636,I149910);
nand I_3766 (I66653,I66636,I149931);
nor I_3767 (I66670,I149910,I149928);
nand I_3768 (I66350,I66486,I66670);
nand I_3769 (I66344,I66435,I149910);
nand I_3770 (I66715,I66537,I149934);
DFFARX1 I_3771 (I66715,I2595,I66370,I66359,);
DFFARX1 I_3772 (I66715,I2595,I66370,I66353,);
not I_3773 (I66760,I149934);
nor I_3774 (I66777,I66760,I149925);
and I_3775 (I66794,I66777,I149910);
or I_3776 (I66811,I66794,I149913);
DFFARX1 I_3777 (I66811,I2595,I66370,I66837,);
nand I_3778 (I66845,I66837,I66503);
nor I_3779 (I66347,I66845,I66653);
nor I_3780 (I66341,I66837,I66469);
DFFARX1 I_3781 (I66837,I2595,I66370,I66899,);
not I_3782 (I66907,I66899);
nor I_3783 (I66356,I66907,I66619);
not I_3784 (I66965,I2602);
DFFARX1 I_3785 (I127409,I2595,I66965,I66991,);
DFFARX1 I_3786 (I66991,I2595,I66965,I67008,);
not I_3787 (I66957,I67008);
not I_3788 (I67030,I66991);
DFFARX1 I_3789 (I127397,I2595,I66965,I67056,);
not I_3790 (I67064,I67056);
and I_3791 (I67081,I67030,I127406);
not I_3792 (I67098,I127403);
nand I_3793 (I67115,I67098,I127406);
not I_3794 (I67132,I127394);
nor I_3795 (I67149,I67132,I127400);
nand I_3796 (I67166,I67149,I127385);
nor I_3797 (I67183,I67166,I67115);
DFFARX1 I_3798 (I67183,I2595,I66965,I66933,);
not I_3799 (I67214,I67166);
not I_3800 (I67231,I127400);
nand I_3801 (I67248,I67231,I127406);
nor I_3802 (I67265,I127400,I127403);
nand I_3803 (I66945,I67081,I67265);
nand I_3804 (I66939,I67030,I127400);
nand I_3805 (I67310,I67132,I127385);
DFFARX1 I_3806 (I67310,I2595,I66965,I66954,);
DFFARX1 I_3807 (I67310,I2595,I66965,I66948,);
not I_3808 (I67355,I127385);
nor I_3809 (I67372,I67355,I127391);
and I_3810 (I67389,I67372,I127388);
or I_3811 (I67406,I67389,I127412);
DFFARX1 I_3812 (I67406,I2595,I66965,I67432,);
nand I_3813 (I67440,I67432,I67098);
nor I_3814 (I66942,I67440,I67248);
nor I_3815 (I66936,I67432,I67064);
DFFARX1 I_3816 (I67432,I2595,I66965,I67494,);
not I_3817 (I67502,I67494);
nor I_3818 (I66951,I67502,I67214);
not I_3819 (I67560,I2602);
DFFARX1 I_3820 (I237755,I2595,I67560,I67586,);
DFFARX1 I_3821 (I67586,I2595,I67560,I67603,);
not I_3822 (I67552,I67603);
not I_3823 (I67625,I67586);
DFFARX1 I_3824 (I237749,I2595,I67560,I67651,);
not I_3825 (I67659,I67651);
and I_3826 (I67676,I67625,I237767);
not I_3827 (I67693,I237755);
nand I_3828 (I67710,I67693,I237767);
not I_3829 (I67727,I237749);
nor I_3830 (I67744,I67727,I237761);
nand I_3831 (I67761,I67744,I237752);
nor I_3832 (I67778,I67761,I67710);
DFFARX1 I_3833 (I67778,I2595,I67560,I67528,);
not I_3834 (I67809,I67761);
not I_3835 (I67826,I237761);
nand I_3836 (I67843,I67826,I237767);
nor I_3837 (I67860,I237761,I237755);
nand I_3838 (I67540,I67676,I67860);
nand I_3839 (I67534,I67625,I237761);
nand I_3840 (I67905,I67727,I237764);
DFFARX1 I_3841 (I67905,I2595,I67560,I67549,);
DFFARX1 I_3842 (I67905,I2595,I67560,I67543,);
not I_3843 (I67950,I237764);
nor I_3844 (I67967,I67950,I237770);
and I_3845 (I67984,I67967,I237752);
or I_3846 (I68001,I67984,I237758);
DFFARX1 I_3847 (I68001,I2595,I67560,I68027,);
nand I_3848 (I68035,I68027,I67693);
nor I_3849 (I67537,I68035,I67843);
nor I_3850 (I67531,I68027,I67659);
DFFARX1 I_3851 (I68027,I2595,I67560,I68089,);
not I_3852 (I68097,I68089);
nor I_3853 (I67546,I68097,I67809);
not I_3854 (I68155,I2602);
DFFARX1 I_3855 (I248822,I2595,I68155,I68181,);
DFFARX1 I_3856 (I68181,I2595,I68155,I68198,);
not I_3857 (I68147,I68198);
not I_3858 (I68220,I68181);
DFFARX1 I_3859 (I248816,I2595,I68155,I68246,);
not I_3860 (I68254,I68246);
and I_3861 (I68271,I68220,I248834);
not I_3862 (I68288,I248822);
nand I_3863 (I68305,I68288,I248834);
not I_3864 (I68322,I248816);
nor I_3865 (I68339,I68322,I248828);
nand I_3866 (I68356,I68339,I248819);
nor I_3867 (I68373,I68356,I68305);
DFFARX1 I_3868 (I68373,I2595,I68155,I68123,);
not I_3869 (I68404,I68356);
not I_3870 (I68421,I248828);
nand I_3871 (I68438,I68421,I248834);
nor I_3872 (I68455,I248828,I248822);
nand I_3873 (I68135,I68271,I68455);
nand I_3874 (I68129,I68220,I248828);
nand I_3875 (I68500,I68322,I248831);
DFFARX1 I_3876 (I68500,I2595,I68155,I68144,);
DFFARX1 I_3877 (I68500,I2595,I68155,I68138,);
not I_3878 (I68545,I248831);
nor I_3879 (I68562,I68545,I248837);
and I_3880 (I68579,I68562,I248819);
or I_3881 (I68596,I68579,I248825);
DFFARX1 I_3882 (I68596,I2595,I68155,I68622,);
nand I_3883 (I68630,I68622,I68288);
nor I_3884 (I68132,I68630,I68438);
nor I_3885 (I68126,I68622,I68254);
DFFARX1 I_3886 (I68622,I2595,I68155,I68684,);
not I_3887 (I68692,I68684);
nor I_3888 (I68141,I68692,I68404);
not I_3889 (I68750,I2602);
DFFARX1 I_3890 (I306174,I2595,I68750,I68776,);
DFFARX1 I_3891 (I68776,I2595,I68750,I68793,);
not I_3892 (I68742,I68793);
not I_3893 (I68815,I68776);
DFFARX1 I_3894 (I306174,I2595,I68750,I68841,);
not I_3895 (I68849,I68841);
and I_3896 (I68866,I68815,I306177);
not I_3897 (I68883,I306189);
nand I_3898 (I68900,I68883,I306177);
not I_3899 (I68917,I306195);
nor I_3900 (I68934,I68917,I306186);
nand I_3901 (I68951,I68934,I306192);
nor I_3902 (I68968,I68951,I68900);
DFFARX1 I_3903 (I68968,I2595,I68750,I68718,);
not I_3904 (I68999,I68951);
not I_3905 (I69016,I306186);
nand I_3906 (I69033,I69016,I306177);
nor I_3907 (I69050,I306186,I306189);
nand I_3908 (I68730,I68866,I69050);
nand I_3909 (I68724,I68815,I306186);
nand I_3910 (I69095,I68917,I306183);
DFFARX1 I_3911 (I69095,I2595,I68750,I68739,);
DFFARX1 I_3912 (I69095,I2595,I68750,I68733,);
not I_3913 (I69140,I306183);
nor I_3914 (I69157,I69140,I306180);
and I_3915 (I69174,I69157,I306198);
or I_3916 (I69191,I69174,I306177);
DFFARX1 I_3917 (I69191,I2595,I68750,I69217,);
nand I_3918 (I69225,I69217,I68883);
nor I_3919 (I68727,I69225,I69033);
nor I_3920 (I68721,I69217,I68849);
DFFARX1 I_3921 (I69217,I2595,I68750,I69279,);
not I_3922 (I69287,I69279);
nor I_3923 (I68736,I69287,I68999);
not I_3924 (I69345,I2602);
DFFARX1 I_3925 (I316578,I2595,I69345,I69371,);
DFFARX1 I_3926 (I69371,I2595,I69345,I69388,);
not I_3927 (I69337,I69388);
not I_3928 (I69410,I69371);
DFFARX1 I_3929 (I316578,I2595,I69345,I69436,);
not I_3930 (I69444,I69436);
and I_3931 (I69461,I69410,I316581);
not I_3932 (I69478,I316593);
nand I_3933 (I69495,I69478,I316581);
not I_3934 (I69512,I316599);
nor I_3935 (I69529,I69512,I316590);
nand I_3936 (I69546,I69529,I316596);
nor I_3937 (I69563,I69546,I69495);
DFFARX1 I_3938 (I69563,I2595,I69345,I69313,);
not I_3939 (I69594,I69546);
not I_3940 (I69611,I316590);
nand I_3941 (I69628,I69611,I316581);
nor I_3942 (I69645,I316590,I316593);
nand I_3943 (I69325,I69461,I69645);
nand I_3944 (I69319,I69410,I316590);
nand I_3945 (I69690,I69512,I316587);
DFFARX1 I_3946 (I69690,I2595,I69345,I69334,);
DFFARX1 I_3947 (I69690,I2595,I69345,I69328,);
not I_3948 (I69735,I316587);
nor I_3949 (I69752,I69735,I316584);
and I_3950 (I69769,I69752,I316602);
or I_3951 (I69786,I69769,I316581);
DFFARX1 I_3952 (I69786,I2595,I69345,I69812,);
nand I_3953 (I69820,I69812,I69478);
nor I_3954 (I69322,I69820,I69628);
nor I_3955 (I69316,I69812,I69444);
DFFARX1 I_3956 (I69812,I2595,I69345,I69874,);
not I_3957 (I69882,I69874);
nor I_3958 (I69331,I69882,I69594);
not I_3959 (I69940,I2602);
DFFARX1 I_3960 (I121969,I2595,I69940,I69966,);
DFFARX1 I_3961 (I69966,I2595,I69940,I69983,);
not I_3962 (I69932,I69983);
not I_3963 (I70005,I69966);
DFFARX1 I_3964 (I121957,I2595,I69940,I70031,);
not I_3965 (I70039,I70031);
and I_3966 (I70056,I70005,I121966);
not I_3967 (I70073,I121963);
nand I_3968 (I70090,I70073,I121966);
not I_3969 (I70107,I121954);
nor I_3970 (I70124,I70107,I121960);
nand I_3971 (I70141,I70124,I121945);
nor I_3972 (I70158,I70141,I70090);
DFFARX1 I_3973 (I70158,I2595,I69940,I69908,);
not I_3974 (I70189,I70141);
not I_3975 (I70206,I121960);
nand I_3976 (I70223,I70206,I121966);
nor I_3977 (I70240,I121960,I121963);
nand I_3978 (I69920,I70056,I70240);
nand I_3979 (I69914,I70005,I121960);
nand I_3980 (I70285,I70107,I121945);
DFFARX1 I_3981 (I70285,I2595,I69940,I69929,);
DFFARX1 I_3982 (I70285,I2595,I69940,I69923,);
not I_3983 (I70330,I121945);
nor I_3984 (I70347,I70330,I121951);
and I_3985 (I70364,I70347,I121948);
or I_3986 (I70381,I70364,I121972);
DFFARX1 I_3987 (I70381,I2595,I69940,I70407,);
nand I_3988 (I70415,I70407,I70073);
nor I_3989 (I69917,I70415,I70223);
nor I_3990 (I69911,I70407,I70039);
DFFARX1 I_3991 (I70407,I2595,I69940,I70469,);
not I_3992 (I70477,I70469);
nor I_3993 (I69926,I70477,I70189);
not I_3994 (I70535,I2602);
DFFARX1 I_3995 (I42955,I2595,I70535,I70561,);
DFFARX1 I_3996 (I70561,I2595,I70535,I70578,);
not I_3997 (I70527,I70578);
not I_3998 (I70600,I70561);
DFFARX1 I_3999 (I42949,I2595,I70535,I70626,);
not I_4000 (I70634,I70626);
and I_4001 (I70651,I70600,I42946);
not I_4002 (I70668,I42967);
nand I_4003 (I70685,I70668,I42946);
not I_4004 (I70702,I42961);
nor I_4005 (I70719,I70702,I42952);
nand I_4006 (I70736,I70719,I42958);
nor I_4007 (I70753,I70736,I70685);
DFFARX1 I_4008 (I70753,I2595,I70535,I70503,);
not I_4009 (I70784,I70736);
not I_4010 (I70801,I42952);
nand I_4011 (I70818,I70801,I42946);
nor I_4012 (I70835,I42952,I42967);
nand I_4013 (I70515,I70651,I70835);
nand I_4014 (I70509,I70600,I42952);
nand I_4015 (I70880,I70702,I42946);
DFFARX1 I_4016 (I70880,I2595,I70535,I70524,);
DFFARX1 I_4017 (I70880,I2595,I70535,I70518,);
not I_4018 (I70925,I42946);
nor I_4019 (I70942,I70925,I42964);
and I_4020 (I70959,I70942,I42970);
or I_4021 (I70976,I70959,I42949);
DFFARX1 I_4022 (I70976,I2595,I70535,I71002,);
nand I_4023 (I71010,I71002,I70668);
nor I_4024 (I70512,I71010,I70818);
nor I_4025 (I70506,I71002,I70634);
DFFARX1 I_4026 (I71002,I2595,I70535,I71064,);
not I_4027 (I71072,I71064);
nor I_4028 (I70521,I71072,I70784);
not I_4029 (I71130,I2602);
DFFARX1 I_4030 (I344272,I2595,I71130,I71156,);
DFFARX1 I_4031 (I71156,I2595,I71130,I71173,);
not I_4032 (I71122,I71173);
not I_4033 (I71195,I71156);
DFFARX1 I_4034 (I344257,I2595,I71130,I71221,);
not I_4035 (I71229,I71221);
and I_4036 (I71246,I71195,I344275);
not I_4037 (I71263,I344257);
nand I_4038 (I71280,I71263,I344275);
not I_4039 (I71297,I344278);
nor I_4040 (I71314,I71297,I344269);
nand I_4041 (I71331,I71314,I344266);
nor I_4042 (I71348,I71331,I71280);
DFFARX1 I_4043 (I71348,I2595,I71130,I71098,);
not I_4044 (I71379,I71331);
not I_4045 (I71396,I344269);
nand I_4046 (I71413,I71396,I344275);
nor I_4047 (I71430,I344269,I344257);
nand I_4048 (I71110,I71246,I71430);
nand I_4049 (I71104,I71195,I344269);
nand I_4050 (I71475,I71297,I344263);
DFFARX1 I_4051 (I71475,I2595,I71130,I71119,);
DFFARX1 I_4052 (I71475,I2595,I71130,I71113,);
not I_4053 (I71520,I344263);
nor I_4054 (I71537,I71520,I344254);
and I_4055 (I71554,I71537,I344260);
or I_4056 (I71571,I71554,I344254);
DFFARX1 I_4057 (I71571,I2595,I71130,I71597,);
nand I_4058 (I71605,I71597,I71263);
nor I_4059 (I71107,I71605,I71413);
nor I_4060 (I71101,I71597,I71229);
DFFARX1 I_4061 (I71597,I2595,I71130,I71659,);
not I_4062 (I71667,I71659);
nor I_4063 (I71116,I71667,I71379);
not I_4064 (I71725,I2602);
DFFARX1 I_4065 (I226388,I2595,I71725,I71751,);
DFFARX1 I_4066 (I71751,I2595,I71725,I71768,);
not I_4067 (I71717,I71768);
not I_4068 (I71790,I71751);
DFFARX1 I_4069 (I226385,I2595,I71725,I71816,);
not I_4070 (I71824,I71816);
and I_4071 (I71841,I71790,I226391);
not I_4072 (I71858,I226376);
nand I_4073 (I71875,I71858,I226391);
not I_4074 (I71892,I226379);
nor I_4075 (I71909,I71892,I226400);
nand I_4076 (I71926,I71909,I226397);
nor I_4077 (I71943,I71926,I71875);
DFFARX1 I_4078 (I71943,I2595,I71725,I71693,);
not I_4079 (I71974,I71926);
not I_4080 (I71991,I226400);
nand I_4081 (I72008,I71991,I226391);
nor I_4082 (I72025,I226400,I226376);
nand I_4083 (I71705,I71841,I72025);
nand I_4084 (I71699,I71790,I226400);
nand I_4085 (I72070,I71892,I226376);
DFFARX1 I_4086 (I72070,I2595,I71725,I71714,);
DFFARX1 I_4087 (I72070,I2595,I71725,I71708,);
not I_4088 (I72115,I226376);
nor I_4089 (I72132,I72115,I226382);
and I_4090 (I72149,I72132,I226394);
or I_4091 (I72166,I72149,I226379);
DFFARX1 I_4092 (I72166,I2595,I71725,I72192,);
nand I_4093 (I72200,I72192,I71858);
nor I_4094 (I71702,I72200,I72008);
nor I_4095 (I71696,I72192,I71824);
DFFARX1 I_4096 (I72192,I2595,I71725,I72254,);
not I_4097 (I72262,I72254);
nor I_4098 (I71711,I72262,I71974);
not I_4099 (I72320,I2602);
DFFARX1 I_4100 (I202690,I2595,I72320,I72346,);
DFFARX1 I_4101 (I72346,I2595,I72320,I72363,);
not I_4102 (I72312,I72363);
not I_4103 (I72385,I72346);
DFFARX1 I_4104 (I202687,I2595,I72320,I72411,);
not I_4105 (I72419,I72411);
and I_4106 (I72436,I72385,I202693);
not I_4107 (I72453,I202678);
nand I_4108 (I72470,I72453,I202693);
not I_4109 (I72487,I202681);
nor I_4110 (I72504,I72487,I202702);
nand I_4111 (I72521,I72504,I202699);
nor I_4112 (I72538,I72521,I72470);
DFFARX1 I_4113 (I72538,I2595,I72320,I72288,);
not I_4114 (I72569,I72521);
not I_4115 (I72586,I202702);
nand I_4116 (I72603,I72586,I202693);
nor I_4117 (I72620,I202702,I202678);
nand I_4118 (I72300,I72436,I72620);
nand I_4119 (I72294,I72385,I202702);
nand I_4120 (I72665,I72487,I202678);
DFFARX1 I_4121 (I72665,I2595,I72320,I72309,);
DFFARX1 I_4122 (I72665,I2595,I72320,I72303,);
not I_4123 (I72710,I202678);
nor I_4124 (I72727,I72710,I202684);
and I_4125 (I72744,I72727,I202696);
or I_4126 (I72761,I72744,I202681);
DFFARX1 I_4127 (I72761,I2595,I72320,I72787,);
nand I_4128 (I72795,I72787,I72453);
nor I_4129 (I72297,I72795,I72603);
nor I_4130 (I72291,I72787,I72419);
DFFARX1 I_4131 (I72787,I2595,I72320,I72849,);
not I_4132 (I72857,I72849);
nor I_4133 (I72306,I72857,I72569);
not I_4134 (I72915,I2602);
DFFARX1 I_4135 (I126865,I2595,I72915,I72941,);
DFFARX1 I_4136 (I72941,I2595,I72915,I72958,);
not I_4137 (I72907,I72958);
not I_4138 (I72980,I72941);
DFFARX1 I_4139 (I126853,I2595,I72915,I73006,);
not I_4140 (I73014,I73006);
and I_4141 (I73031,I72980,I126862);
not I_4142 (I73048,I126859);
nand I_4143 (I73065,I73048,I126862);
not I_4144 (I73082,I126850);
nor I_4145 (I73099,I73082,I126856);
nand I_4146 (I73116,I73099,I126841);
nor I_4147 (I73133,I73116,I73065);
DFFARX1 I_4148 (I73133,I2595,I72915,I72883,);
not I_4149 (I73164,I73116);
not I_4150 (I73181,I126856);
nand I_4151 (I73198,I73181,I126862);
nor I_4152 (I73215,I126856,I126859);
nand I_4153 (I72895,I73031,I73215);
nand I_4154 (I72889,I72980,I126856);
nand I_4155 (I73260,I73082,I126841);
DFFARX1 I_4156 (I73260,I2595,I72915,I72904,);
DFFARX1 I_4157 (I73260,I2595,I72915,I72898,);
not I_4158 (I73305,I126841);
nor I_4159 (I73322,I73305,I126847);
and I_4160 (I73339,I73322,I126844);
or I_4161 (I73356,I73339,I126868);
DFFARX1 I_4162 (I73356,I2595,I72915,I73382,);
nand I_4163 (I73390,I73382,I73048);
nor I_4164 (I72892,I73390,I73198);
nor I_4165 (I72886,I73382,I73014);
DFFARX1 I_4166 (I73382,I2595,I72915,I73444,);
not I_4167 (I73452,I73444);
nor I_4168 (I72901,I73452,I73164);
not I_4169 (I73510,I2602);
DFFARX1 I_4170 (I2623,I2595,I73510,I73536,);
DFFARX1 I_4171 (I73536,I2595,I73510,I73553,);
not I_4172 (I73502,I73553);
not I_4173 (I73575,I73536);
DFFARX1 I_4174 (I2620,I2595,I73510,I73601,);
not I_4175 (I73609,I73601);
and I_4176 (I73626,I73575,I2611);
not I_4177 (I73643,I2608);
nand I_4178 (I73660,I73643,I2611);
not I_4179 (I73677,I2608);
nor I_4180 (I73694,I73677,I2605);
nand I_4181 (I73711,I73694,I2617);
nor I_4182 (I73728,I73711,I73660);
DFFARX1 I_4183 (I73728,I2595,I73510,I73478,);
not I_4184 (I73759,I73711);
not I_4185 (I73776,I2605);
nand I_4186 (I73793,I73776,I2611);
nor I_4187 (I73810,I2605,I2608);
nand I_4188 (I73490,I73626,I73810);
nand I_4189 (I73484,I73575,I2605);
nand I_4190 (I73855,I73677,I2614);
DFFARX1 I_4191 (I73855,I2595,I73510,I73499,);
DFFARX1 I_4192 (I73855,I2595,I73510,I73493,);
not I_4193 (I73900,I2614);
nor I_4194 (I73917,I73900,I2626);
and I_4195 (I73934,I73917,I2611);
or I_4196 (I73951,I73934,I2605);
DFFARX1 I_4197 (I73951,I2595,I73510,I73977,);
nand I_4198 (I73985,I73977,I73643);
nor I_4199 (I73487,I73985,I73793);
nor I_4200 (I73481,I73977,I73609);
DFFARX1 I_4201 (I73977,I2595,I73510,I74039,);
not I_4202 (I74047,I74039);
nor I_4203 (I73496,I74047,I73759);
not I_4204 (I74105,I2602);
DFFARX1 I_4205 (I138289,I2595,I74105,I74131,);
DFFARX1 I_4206 (I74131,I2595,I74105,I74148,);
not I_4207 (I74097,I74148);
not I_4208 (I74170,I74131);
DFFARX1 I_4209 (I138277,I2595,I74105,I74196,);
not I_4210 (I74204,I74196);
and I_4211 (I74221,I74170,I138286);
not I_4212 (I74238,I138283);
nand I_4213 (I74255,I74238,I138286);
not I_4214 (I74272,I138274);
nor I_4215 (I74289,I74272,I138280);
nand I_4216 (I74306,I74289,I138265);
nor I_4217 (I74323,I74306,I74255);
DFFARX1 I_4218 (I74323,I2595,I74105,I74073,);
not I_4219 (I74354,I74306);
not I_4220 (I74371,I138280);
nand I_4221 (I74388,I74371,I138286);
nor I_4222 (I74405,I138280,I138283);
nand I_4223 (I74085,I74221,I74405);
nand I_4224 (I74079,I74170,I138280);
nand I_4225 (I74450,I74272,I138265);
DFFARX1 I_4226 (I74450,I2595,I74105,I74094,);
DFFARX1 I_4227 (I74450,I2595,I74105,I74088,);
not I_4228 (I74495,I138265);
nor I_4229 (I74512,I74495,I138271);
and I_4230 (I74529,I74512,I138268);
or I_4231 (I74546,I74529,I138292);
DFFARX1 I_4232 (I74546,I2595,I74105,I74572,);
nand I_4233 (I74580,I74572,I74238);
nor I_4234 (I74082,I74580,I74388);
nor I_4235 (I74076,I74572,I74204);
DFFARX1 I_4236 (I74572,I2595,I74105,I74634,);
not I_4237 (I74642,I74634);
nor I_4238 (I74091,I74642,I74354);
not I_4239 (I74700,I2602);
DFFARX1 I_4240 (I183038,I2595,I74700,I74726,);
DFFARX1 I_4241 (I74726,I2595,I74700,I74743,);
not I_4242 (I74692,I74743);
not I_4243 (I74765,I74726);
DFFARX1 I_4244 (I183035,I2595,I74700,I74791,);
not I_4245 (I74799,I74791);
and I_4246 (I74816,I74765,I183041);
not I_4247 (I74833,I183026);
nand I_4248 (I74850,I74833,I183041);
not I_4249 (I74867,I183029);
nor I_4250 (I74884,I74867,I183050);
nand I_4251 (I74901,I74884,I183047);
nor I_4252 (I74918,I74901,I74850);
DFFARX1 I_4253 (I74918,I2595,I74700,I74668,);
not I_4254 (I74949,I74901);
not I_4255 (I74966,I183050);
nand I_4256 (I74983,I74966,I183041);
nor I_4257 (I75000,I183050,I183026);
nand I_4258 (I74680,I74816,I75000);
nand I_4259 (I74674,I74765,I183050);
nand I_4260 (I75045,I74867,I183026);
DFFARX1 I_4261 (I75045,I2595,I74700,I74689,);
DFFARX1 I_4262 (I75045,I2595,I74700,I74683,);
not I_4263 (I75090,I183026);
nor I_4264 (I75107,I75090,I183032);
and I_4265 (I75124,I75107,I183044);
or I_4266 (I75141,I75124,I183029);
DFFARX1 I_4267 (I75141,I2595,I74700,I75167,);
nand I_4268 (I75175,I75167,I74833);
nor I_4269 (I74677,I75175,I74983);
nor I_4270 (I74671,I75167,I74799);
DFFARX1 I_4271 (I75167,I2595,I74700,I75229,);
not I_4272 (I75237,I75229);
nor I_4273 (I74686,I75237,I74949);
not I_4274 (I75295,I2602);
DFFARX1 I_4275 (I2476,I2595,I75295,I75321,);
DFFARX1 I_4276 (I75321,I2595,I75295,I75338,);
not I_4277 (I75287,I75338);
not I_4278 (I75360,I75321);
DFFARX1 I_4279 (I2452,I2595,I75295,I75386,);
not I_4280 (I75394,I75386);
and I_4281 (I75411,I75360,I2028);
not I_4282 (I75428,I1436);
nand I_4283 (I75445,I75428,I2028);
not I_4284 (I75462,I1948);
nor I_4285 (I75479,I75462,I1492);
nand I_4286 (I75496,I75479,I2204);
nor I_4287 (I75513,I75496,I75445);
DFFARX1 I_4288 (I75513,I2595,I75295,I75263,);
not I_4289 (I75544,I75496);
not I_4290 (I75561,I1492);
nand I_4291 (I75578,I75561,I2028);
nor I_4292 (I75595,I1492,I1436);
nand I_4293 (I75275,I75411,I75595);
nand I_4294 (I75269,I75360,I1492);
nand I_4295 (I75640,I75462,I1620);
DFFARX1 I_4296 (I75640,I2595,I75295,I75284,);
DFFARX1 I_4297 (I75640,I2595,I75295,I75278,);
not I_4298 (I75685,I1620);
nor I_4299 (I75702,I75685,I1860);
and I_4300 (I75719,I75702,I1828);
or I_4301 (I75736,I75719,I1396);
DFFARX1 I_4302 (I75736,I2595,I75295,I75762,);
nand I_4303 (I75770,I75762,I75428);
nor I_4304 (I75272,I75770,I75578);
nor I_4305 (I75266,I75762,I75394);
DFFARX1 I_4306 (I75762,I2595,I75295,I75824,);
not I_4307 (I75832,I75824);
nor I_4308 (I75281,I75832,I75544);
not I_4309 (I75890,I2602);
DFFARX1 I_4310 (I116529,I2595,I75890,I75916,);
DFFARX1 I_4311 (I75916,I2595,I75890,I75933,);
not I_4312 (I75882,I75933);
not I_4313 (I75955,I75916);
DFFARX1 I_4314 (I116517,I2595,I75890,I75981,);
not I_4315 (I75989,I75981);
and I_4316 (I76006,I75955,I116526);
not I_4317 (I76023,I116523);
nand I_4318 (I76040,I76023,I116526);
not I_4319 (I76057,I116514);
nor I_4320 (I76074,I76057,I116520);
nand I_4321 (I76091,I76074,I116505);
nor I_4322 (I76108,I76091,I76040);
DFFARX1 I_4323 (I76108,I2595,I75890,I75858,);
not I_4324 (I76139,I76091);
not I_4325 (I76156,I116520);
nand I_4326 (I76173,I76156,I116526);
nor I_4327 (I76190,I116520,I116523);
nand I_4328 (I75870,I76006,I76190);
nand I_4329 (I75864,I75955,I116520);
nand I_4330 (I76235,I76057,I116505);
DFFARX1 I_4331 (I76235,I2595,I75890,I75879,);
DFFARX1 I_4332 (I76235,I2595,I75890,I75873,);
not I_4333 (I76280,I116505);
nor I_4334 (I76297,I76280,I116511);
and I_4335 (I76314,I76297,I116508);
or I_4336 (I76331,I76314,I116532);
DFFARX1 I_4337 (I76331,I2595,I75890,I76357,);
nand I_4338 (I76365,I76357,I76023);
nor I_4339 (I75867,I76365,I76173);
nor I_4340 (I75861,I76357,I75989);
DFFARX1 I_4341 (I76357,I2595,I75890,I76419,);
not I_4342 (I76427,I76419);
nor I_4343 (I75876,I76427,I76139);
not I_4344 (I76485,I2602);
DFFARX1 I_4345 (I158765,I2595,I76485,I76511,);
DFFARX1 I_4346 (I76511,I2595,I76485,I76528,);
not I_4347 (I76477,I76528);
not I_4348 (I76550,I76511);
DFFARX1 I_4349 (I158756,I2595,I76485,I76576,);
not I_4350 (I76584,I76576);
and I_4351 (I76601,I76550,I158774);
not I_4352 (I76618,I158771);
nand I_4353 (I76635,I76618,I158774);
not I_4354 (I76652,I158750);
nor I_4355 (I76669,I76652,I158753);
nand I_4356 (I76686,I76669,I158762);
nor I_4357 (I76703,I76686,I76635);
DFFARX1 I_4358 (I76703,I2595,I76485,I76453,);
not I_4359 (I76734,I76686);
not I_4360 (I76751,I158753);
nand I_4361 (I76768,I76751,I158774);
nor I_4362 (I76785,I158753,I158771);
nand I_4363 (I76465,I76601,I76785);
nand I_4364 (I76459,I76550,I158753);
nand I_4365 (I76830,I76652,I158768);
DFFARX1 I_4366 (I76830,I2595,I76485,I76474,);
DFFARX1 I_4367 (I76830,I2595,I76485,I76468,);
not I_4368 (I76875,I158768);
nor I_4369 (I76892,I76875,I158750);
and I_4370 (I76909,I76892,I158759);
or I_4371 (I76926,I76909,I158753);
DFFARX1 I_4372 (I76926,I2595,I76485,I76952,);
nand I_4373 (I76960,I76952,I76618);
nor I_4374 (I76462,I76960,I76768);
nor I_4375 (I76456,I76952,I76584);
DFFARX1 I_4376 (I76952,I2595,I76485,I77014,);
not I_4377 (I77022,I77014);
nor I_4378 (I76471,I77022,I76734);
not I_4379 (I77080,I2602);
DFFARX1 I_4380 (I221764,I2595,I77080,I77106,);
DFFARX1 I_4381 (I77106,I2595,I77080,I77123,);
not I_4382 (I77072,I77123);
not I_4383 (I77145,I77106);
DFFARX1 I_4384 (I221761,I2595,I77080,I77171,);
not I_4385 (I77179,I77171);
and I_4386 (I77196,I77145,I221767);
not I_4387 (I77213,I221752);
nand I_4388 (I77230,I77213,I221767);
not I_4389 (I77247,I221755);
nor I_4390 (I77264,I77247,I221776);
nand I_4391 (I77281,I77264,I221773);
nor I_4392 (I77298,I77281,I77230);
DFFARX1 I_4393 (I77298,I2595,I77080,I77048,);
not I_4394 (I77329,I77281);
not I_4395 (I77346,I221776);
nand I_4396 (I77363,I77346,I221767);
nor I_4397 (I77380,I221776,I221752);
nand I_4398 (I77060,I77196,I77380);
nand I_4399 (I77054,I77145,I221776);
nand I_4400 (I77425,I77247,I221752);
DFFARX1 I_4401 (I77425,I2595,I77080,I77069,);
DFFARX1 I_4402 (I77425,I2595,I77080,I77063,);
not I_4403 (I77470,I221752);
nor I_4404 (I77487,I77470,I221758);
and I_4405 (I77504,I77487,I221770);
or I_4406 (I77521,I77504,I221755);
DFFARX1 I_4407 (I77521,I2595,I77080,I77547,);
nand I_4408 (I77555,I77547,I77213);
nor I_4409 (I77057,I77555,I77363);
nor I_4410 (I77051,I77547,I77179);
DFFARX1 I_4411 (I77547,I2595,I77080,I77609,);
not I_4412 (I77617,I77609);
nor I_4413 (I77066,I77617,I77329);
not I_4414 (I77675,I2602);
DFFARX1 I_4415 (I115441,I2595,I77675,I77701,);
DFFARX1 I_4416 (I77701,I2595,I77675,I77718,);
not I_4417 (I77667,I77718);
not I_4418 (I77740,I77701);
DFFARX1 I_4419 (I115429,I2595,I77675,I77766,);
not I_4420 (I77774,I77766);
and I_4421 (I77791,I77740,I115438);
not I_4422 (I77808,I115435);
nand I_4423 (I77825,I77808,I115438);
not I_4424 (I77842,I115426);
nor I_4425 (I77859,I77842,I115432);
nand I_4426 (I77876,I77859,I115417);
nor I_4427 (I77893,I77876,I77825);
DFFARX1 I_4428 (I77893,I2595,I77675,I77643,);
not I_4429 (I77924,I77876);
not I_4430 (I77941,I115432);
nand I_4431 (I77958,I77941,I115438);
nor I_4432 (I77975,I115432,I115435);
nand I_4433 (I77655,I77791,I77975);
nand I_4434 (I77649,I77740,I115432);
nand I_4435 (I78020,I77842,I115417);
DFFARX1 I_4436 (I78020,I2595,I77675,I77664,);
DFFARX1 I_4437 (I78020,I2595,I77675,I77658,);
not I_4438 (I78065,I115417);
nor I_4439 (I78082,I78065,I115423);
and I_4440 (I78099,I78082,I115420);
or I_4441 (I78116,I78099,I115444);
DFFARX1 I_4442 (I78116,I2595,I77675,I78142,);
nand I_4443 (I78150,I78142,I77808);
nor I_4444 (I77652,I78150,I77958);
nor I_4445 (I77646,I78142,I77774);
DFFARX1 I_4446 (I78142,I2595,I77675,I78204,);
not I_4447 (I78212,I78204);
nor I_4448 (I77661,I78212,I77924);
not I_4449 (I78270,I2602);
DFFARX1 I_4450 (I308486,I2595,I78270,I78296,);
DFFARX1 I_4451 (I78296,I2595,I78270,I78313,);
not I_4452 (I78262,I78313);
not I_4453 (I78335,I78296);
DFFARX1 I_4454 (I308486,I2595,I78270,I78361,);
not I_4455 (I78369,I78361);
and I_4456 (I78386,I78335,I308489);
not I_4457 (I78403,I308501);
nand I_4458 (I78420,I78403,I308489);
not I_4459 (I78437,I308507);
nor I_4460 (I78454,I78437,I308498);
nand I_4461 (I78471,I78454,I308504);
nor I_4462 (I78488,I78471,I78420);
DFFARX1 I_4463 (I78488,I2595,I78270,I78238,);
not I_4464 (I78519,I78471);
not I_4465 (I78536,I308498);
nand I_4466 (I78553,I78536,I308489);
nor I_4467 (I78570,I308498,I308501);
nand I_4468 (I78250,I78386,I78570);
nand I_4469 (I78244,I78335,I308498);
nand I_4470 (I78615,I78437,I308495);
DFFARX1 I_4471 (I78615,I2595,I78270,I78259,);
DFFARX1 I_4472 (I78615,I2595,I78270,I78253,);
not I_4473 (I78660,I308495);
nor I_4474 (I78677,I78660,I308492);
and I_4475 (I78694,I78677,I308510);
or I_4476 (I78711,I78694,I308489);
DFFARX1 I_4477 (I78711,I2595,I78270,I78737,);
nand I_4478 (I78745,I78737,I78403);
nor I_4479 (I78247,I78745,I78553);
nor I_4480 (I78241,I78737,I78369);
DFFARX1 I_4481 (I78737,I2595,I78270,I78799,);
not I_4482 (I78807,I78799);
nor I_4483 (I78256,I78807,I78519);
not I_4484 (I78865,I2602);
DFFARX1 I_4485 (I215406,I2595,I78865,I78891,);
DFFARX1 I_4486 (I78891,I2595,I78865,I78908,);
not I_4487 (I78857,I78908);
not I_4488 (I78930,I78891);
DFFARX1 I_4489 (I215403,I2595,I78865,I78956,);
not I_4490 (I78964,I78956);
and I_4491 (I78981,I78930,I215409);
not I_4492 (I78998,I215394);
nand I_4493 (I79015,I78998,I215409);
not I_4494 (I79032,I215397);
nor I_4495 (I79049,I79032,I215418);
nand I_4496 (I79066,I79049,I215415);
nor I_4497 (I79083,I79066,I79015);
DFFARX1 I_4498 (I79083,I2595,I78865,I78833,);
not I_4499 (I79114,I79066);
not I_4500 (I79131,I215418);
nand I_4501 (I79148,I79131,I215409);
nor I_4502 (I79165,I215418,I215394);
nand I_4503 (I78845,I78981,I79165);
nand I_4504 (I78839,I78930,I215418);
nand I_4505 (I79210,I79032,I215394);
DFFARX1 I_4506 (I79210,I2595,I78865,I78854,);
DFFARX1 I_4507 (I79210,I2595,I78865,I78848,);
not I_4508 (I79255,I215394);
nor I_4509 (I79272,I79255,I215400);
and I_4510 (I79289,I79272,I215412);
or I_4511 (I79306,I79289,I215397);
DFFARX1 I_4512 (I79306,I2595,I78865,I79332,);
nand I_4513 (I79340,I79332,I78998);
nor I_4514 (I78842,I79340,I79148);
nor I_4515 (I78836,I79332,I78964);
DFFARX1 I_4516 (I79332,I2595,I78865,I79394,);
not I_4517 (I79402,I79394);
nor I_4518 (I78851,I79402,I79114);
not I_4519 (I79460,I2602);
DFFARX1 I_4520 (I240917,I2595,I79460,I79486,);
DFFARX1 I_4521 (I79486,I2595,I79460,I79503,);
not I_4522 (I79452,I79503);
not I_4523 (I79525,I79486);
DFFARX1 I_4524 (I240911,I2595,I79460,I79551,);
not I_4525 (I79559,I79551);
and I_4526 (I79576,I79525,I240929);
not I_4527 (I79593,I240917);
nand I_4528 (I79610,I79593,I240929);
not I_4529 (I79627,I240911);
nor I_4530 (I79644,I79627,I240923);
nand I_4531 (I79661,I79644,I240914);
nor I_4532 (I79678,I79661,I79610);
DFFARX1 I_4533 (I79678,I2595,I79460,I79428,);
not I_4534 (I79709,I79661);
not I_4535 (I79726,I240923);
nand I_4536 (I79743,I79726,I240929);
nor I_4537 (I79760,I240923,I240917);
nand I_4538 (I79440,I79576,I79760);
nand I_4539 (I79434,I79525,I240923);
nand I_4540 (I79805,I79627,I240926);
DFFARX1 I_4541 (I79805,I2595,I79460,I79449,);
DFFARX1 I_4542 (I79805,I2595,I79460,I79443,);
not I_4543 (I79850,I240926);
nor I_4544 (I79867,I79850,I240932);
and I_4545 (I79884,I79867,I240914);
or I_4546 (I79901,I79884,I240920);
DFFARX1 I_4547 (I79901,I2595,I79460,I79927,);
nand I_4548 (I79935,I79927,I79593);
nor I_4549 (I79437,I79935,I79743);
nor I_4550 (I79431,I79927,I79559);
DFFARX1 I_4551 (I79927,I2595,I79460,I79989,);
not I_4552 (I79997,I79989);
nor I_4553 (I79446,I79997,I79709);
not I_4554 (I80055,I2602);
DFFARX1 I_4555 (I270608,I2595,I80055,I80081,);
DFFARX1 I_4556 (I80081,I2595,I80055,I80098,);
not I_4557 (I80047,I80098);
not I_4558 (I80120,I80081);
DFFARX1 I_4559 (I270617,I2595,I80055,I80146,);
not I_4560 (I80154,I80146);
and I_4561 (I80171,I80120,I270605);
not I_4562 (I80188,I270596);
nand I_4563 (I80205,I80188,I270605);
not I_4564 (I80222,I270602);
nor I_4565 (I80239,I80222,I270620);
nand I_4566 (I80256,I80239,I270593);
nor I_4567 (I80273,I80256,I80205);
DFFARX1 I_4568 (I80273,I2595,I80055,I80023,);
not I_4569 (I80304,I80256);
not I_4570 (I80321,I270620);
nand I_4571 (I80338,I80321,I270605);
nor I_4572 (I80355,I270620,I270596);
nand I_4573 (I80035,I80171,I80355);
nand I_4574 (I80029,I80120,I270620);
nand I_4575 (I80400,I80222,I270599);
DFFARX1 I_4576 (I80400,I2595,I80055,I80044,);
DFFARX1 I_4577 (I80400,I2595,I80055,I80038,);
not I_4578 (I80445,I270599);
nor I_4579 (I80462,I80445,I270611);
and I_4580 (I80479,I80462,I270593);
or I_4581 (I80496,I80479,I270614);
DFFARX1 I_4582 (I80496,I2595,I80055,I80522,);
nand I_4583 (I80530,I80522,I80188);
nor I_4584 (I80032,I80530,I80338);
nor I_4585 (I80026,I80522,I80154);
DFFARX1 I_4586 (I80522,I2595,I80055,I80584,);
not I_4587 (I80592,I80584);
nor I_4588 (I80041,I80592,I80304);
not I_4589 (I80653,I2602);
DFFARX1 I_4590 (I131749,I2595,I80653,I80679,);
nand I_4591 (I80687,I131761,I131740);
and I_4592 (I80704,I80687,I131764);
DFFARX1 I_4593 (I80704,I2595,I80653,I80730,);
nor I_4594 (I80621,I80730,I80679);
not I_4595 (I80752,I80730);
DFFARX1 I_4596 (I131755,I2595,I80653,I80778,);
nand I_4597 (I80786,I80778,I131737);
not I_4598 (I80803,I80786);
DFFARX1 I_4599 (I80803,I2595,I80653,I80829,);
not I_4600 (I80645,I80829);
nor I_4601 (I80851,I80679,I80786);
nor I_4602 (I80627,I80730,I80851);
DFFARX1 I_4603 (I131752,I2595,I80653,I80891,);
DFFARX1 I_4604 (I80891,I2595,I80653,I80908,);
not I_4605 (I80916,I80908);
not I_4606 (I80933,I80891);
nand I_4607 (I80630,I80933,I80752);
nand I_4608 (I80964,I131737,I131743);
and I_4609 (I80981,I80964,I131746);
DFFARX1 I_4610 (I80981,I2595,I80653,I81007,);
nor I_4611 (I81015,I81007,I80679);
DFFARX1 I_4612 (I81015,I2595,I80653,I80618,);
DFFARX1 I_4613 (I81007,I2595,I80653,I80636,);
nor I_4614 (I81060,I131758,I131743);
not I_4615 (I81077,I81060);
nor I_4616 (I80639,I80916,I81077);
nand I_4617 (I80624,I80933,I81077);
nor I_4618 (I80633,I80679,I81060);
DFFARX1 I_4619 (I81060,I2595,I80653,I80642,);
not I_4620 (I81180,I2602);
DFFARX1 I_4621 (I65743,I2595,I81180,I81206,);
nand I_4622 (I81214,I65743,I65749);
and I_4623 (I81231,I81214,I65767);
DFFARX1 I_4624 (I81231,I2595,I81180,I81257,);
nor I_4625 (I81148,I81257,I81206);
not I_4626 (I81279,I81257);
DFFARX1 I_4627 (I65755,I2595,I81180,I81305,);
nand I_4628 (I81313,I81305,I65752);
not I_4629 (I81330,I81313);
DFFARX1 I_4630 (I81330,I2595,I81180,I81356,);
not I_4631 (I81172,I81356);
nor I_4632 (I81378,I81206,I81313);
nor I_4633 (I81154,I81257,I81378);
DFFARX1 I_4634 (I65761,I2595,I81180,I81418,);
DFFARX1 I_4635 (I81418,I2595,I81180,I81435,);
not I_4636 (I81443,I81435);
not I_4637 (I81460,I81418);
nand I_4638 (I81157,I81460,I81279);
nand I_4639 (I81491,I65746,I65746);
and I_4640 (I81508,I81491,I65758);
DFFARX1 I_4641 (I81508,I2595,I81180,I81534,);
nor I_4642 (I81542,I81534,I81206);
DFFARX1 I_4643 (I81542,I2595,I81180,I81145,);
DFFARX1 I_4644 (I81534,I2595,I81180,I81163,);
nor I_4645 (I81587,I65764,I65746);
not I_4646 (I81604,I81587);
nor I_4647 (I81166,I81443,I81604);
nand I_4648 (I81151,I81460,I81604);
nor I_4649 (I81160,I81206,I81587);
DFFARX1 I_4650 (I81587,I2595,I81180,I81169,);
not I_4651 (I81707,I2602);
DFFARX1 I_4652 (I307330,I2595,I81707,I81733,);
nand I_4653 (I81741,I307345,I307330);
and I_4654 (I81758,I81741,I307348);
DFFARX1 I_4655 (I81758,I2595,I81707,I81784,);
nor I_4656 (I81675,I81784,I81733);
not I_4657 (I81806,I81784);
DFFARX1 I_4658 (I307354,I2595,I81707,I81832,);
nand I_4659 (I81840,I81832,I307336);
not I_4660 (I81857,I81840);
DFFARX1 I_4661 (I81857,I2595,I81707,I81883,);
not I_4662 (I81699,I81883);
nor I_4663 (I81905,I81733,I81840);
nor I_4664 (I81681,I81784,I81905);
DFFARX1 I_4665 (I307333,I2595,I81707,I81945,);
DFFARX1 I_4666 (I81945,I2595,I81707,I81962,);
not I_4667 (I81970,I81962);
not I_4668 (I81987,I81945);
nand I_4669 (I81684,I81987,I81806);
nand I_4670 (I82018,I307333,I307339);
and I_4671 (I82035,I82018,I307351);
DFFARX1 I_4672 (I82035,I2595,I81707,I82061,);
nor I_4673 (I82069,I82061,I81733);
DFFARX1 I_4674 (I82069,I2595,I81707,I81672,);
DFFARX1 I_4675 (I82061,I2595,I81707,I81690,);
nor I_4676 (I82114,I307342,I307339);
not I_4677 (I82131,I82114);
nor I_4678 (I81693,I81970,I82131);
nand I_4679 (I81678,I81987,I82131);
nor I_4680 (I81687,I81733,I82114);
DFFARX1 I_4681 (I82114,I2595,I81707,I81696,);
not I_4682 (I82234,I2602);
DFFARX1 I_4683 (I328716,I2595,I82234,I82260,);
nand I_4684 (I82268,I328731,I328716);
and I_4685 (I82285,I82268,I328734);
DFFARX1 I_4686 (I82285,I2595,I82234,I82311,);
nor I_4687 (I82202,I82311,I82260);
not I_4688 (I82333,I82311);
DFFARX1 I_4689 (I328740,I2595,I82234,I82359,);
nand I_4690 (I82367,I82359,I328722);
not I_4691 (I82384,I82367);
DFFARX1 I_4692 (I82384,I2595,I82234,I82410,);
not I_4693 (I82226,I82410);
nor I_4694 (I82432,I82260,I82367);
nor I_4695 (I82208,I82311,I82432);
DFFARX1 I_4696 (I328719,I2595,I82234,I82472,);
DFFARX1 I_4697 (I82472,I2595,I82234,I82489,);
not I_4698 (I82497,I82489);
not I_4699 (I82514,I82472);
nand I_4700 (I82211,I82514,I82333);
nand I_4701 (I82545,I328719,I328725);
and I_4702 (I82562,I82545,I328737);
DFFARX1 I_4703 (I82562,I2595,I82234,I82588,);
nor I_4704 (I82596,I82588,I82260);
DFFARX1 I_4705 (I82596,I2595,I82234,I82199,);
DFFARX1 I_4706 (I82588,I2595,I82234,I82217,);
nor I_4707 (I82641,I328728,I328725);
not I_4708 (I82658,I82641);
nor I_4709 (I82220,I82497,I82658);
nand I_4710 (I82205,I82514,I82658);
nor I_4711 (I82214,I82260,I82641);
DFFARX1 I_4712 (I82641,I2595,I82234,I82223,);
not I_4713 (I82761,I2602);
DFFARX1 I_4714 (I37152,I2595,I82761,I82787,);
nand I_4715 (I82795,I37164,I37173);
and I_4716 (I82812,I82795,I37152);
DFFARX1 I_4717 (I82812,I2595,I82761,I82838,);
nor I_4718 (I82729,I82838,I82787);
not I_4719 (I82860,I82838);
DFFARX1 I_4720 (I37167,I2595,I82761,I82886,);
nand I_4721 (I82894,I82886,I37155);
not I_4722 (I82911,I82894);
DFFARX1 I_4723 (I82911,I2595,I82761,I82937,);
not I_4724 (I82753,I82937);
nor I_4725 (I82959,I82787,I82894);
nor I_4726 (I82735,I82838,I82959);
DFFARX1 I_4727 (I37158,I2595,I82761,I82999,);
DFFARX1 I_4728 (I82999,I2595,I82761,I83016,);
not I_4729 (I83024,I83016);
not I_4730 (I83041,I82999);
nand I_4731 (I82738,I83041,I82860);
nand I_4732 (I83072,I37149,I37149);
and I_4733 (I83089,I83072,I37161);
DFFARX1 I_4734 (I83089,I2595,I82761,I83115,);
nor I_4735 (I83123,I83115,I82787);
DFFARX1 I_4736 (I83123,I2595,I82761,I82726,);
DFFARX1 I_4737 (I83115,I2595,I82761,I82744,);
nor I_4738 (I83168,I37170,I37149);
not I_4739 (I83185,I83168);
nor I_4740 (I82747,I83024,I83185);
nand I_4741 (I82732,I83041,I83185);
nor I_4742 (I82741,I82787,I83168);
DFFARX1 I_4743 (I83168,I2595,I82761,I82750,);
not I_4744 (I83288,I2602);
DFFARX1 I_4745 (I240387,I2595,I83288,I83314,);
nand I_4746 (I83322,I240390,I240384);
and I_4747 (I83339,I83322,I240396);
DFFARX1 I_4748 (I83339,I2595,I83288,I83365,);
nor I_4749 (I83256,I83365,I83314);
not I_4750 (I83387,I83365);
DFFARX1 I_4751 (I240399,I2595,I83288,I83413,);
nand I_4752 (I83421,I83413,I240390);
not I_4753 (I83438,I83421);
DFFARX1 I_4754 (I83438,I2595,I83288,I83464,);
not I_4755 (I83280,I83464);
nor I_4756 (I83486,I83314,I83421);
nor I_4757 (I83262,I83365,I83486);
DFFARX1 I_4758 (I240402,I2595,I83288,I83526,);
DFFARX1 I_4759 (I83526,I2595,I83288,I83543,);
not I_4760 (I83551,I83543);
not I_4761 (I83568,I83526);
nand I_4762 (I83265,I83568,I83387);
nand I_4763 (I83599,I240384,I240393);
and I_4764 (I83616,I83599,I240387);
DFFARX1 I_4765 (I83616,I2595,I83288,I83642,);
nor I_4766 (I83650,I83642,I83314);
DFFARX1 I_4767 (I83650,I2595,I83288,I83253,);
DFFARX1 I_4768 (I83642,I2595,I83288,I83271,);
nor I_4769 (I83695,I240405,I240393);
not I_4770 (I83712,I83695);
nor I_4771 (I83274,I83551,I83712);
nand I_4772 (I83259,I83568,I83712);
nor I_4773 (I83268,I83314,I83695);
DFFARX1 I_4774 (I83695,I2595,I83288,I83277,);
not I_4775 (I83815,I2602);
DFFARX1 I_4776 (I291013,I2595,I83815,I83841,);
nand I_4777 (I83849,I291010,I291013);
and I_4778 (I83866,I83849,I291022);
DFFARX1 I_4779 (I83866,I2595,I83815,I83892,);
nor I_4780 (I83783,I83892,I83841);
not I_4781 (I83914,I83892);
DFFARX1 I_4782 (I291010,I2595,I83815,I83940,);
nand I_4783 (I83948,I83940,I291028);
not I_4784 (I83965,I83948);
DFFARX1 I_4785 (I83965,I2595,I83815,I83991,);
not I_4786 (I83807,I83991);
nor I_4787 (I84013,I83841,I83948);
nor I_4788 (I83789,I83892,I84013);
DFFARX1 I_4789 (I291016,I2595,I83815,I84053,);
DFFARX1 I_4790 (I84053,I2595,I83815,I84070,);
not I_4791 (I84078,I84070);
not I_4792 (I84095,I84053);
nand I_4793 (I83792,I84095,I83914);
nand I_4794 (I84126,I291025,I291031);
and I_4795 (I84143,I84126,I291016);
DFFARX1 I_4796 (I84143,I2595,I83815,I84169,);
nor I_4797 (I84177,I84169,I83841);
DFFARX1 I_4798 (I84177,I2595,I83815,I83780,);
DFFARX1 I_4799 (I84169,I2595,I83815,I83798,);
nor I_4800 (I84222,I291019,I291031);
not I_4801 (I84239,I84222);
nor I_4802 (I83801,I84078,I84239);
nand I_4803 (I83786,I84095,I84239);
nor I_4804 (I83795,I83841,I84222);
DFFARX1 I_4805 (I84222,I2595,I83815,I83804,);
not I_4806 (I84342,I2602);
DFFARX1 I_4807 (I320046,I2595,I84342,I84368,);
nand I_4808 (I84376,I320061,I320046);
and I_4809 (I84393,I84376,I320064);
DFFARX1 I_4810 (I84393,I2595,I84342,I84419,);
nor I_4811 (I84310,I84419,I84368);
not I_4812 (I84441,I84419);
DFFARX1 I_4813 (I320070,I2595,I84342,I84467,);
nand I_4814 (I84475,I84467,I320052);
not I_4815 (I84492,I84475);
DFFARX1 I_4816 (I84492,I2595,I84342,I84518,);
not I_4817 (I84334,I84518);
nor I_4818 (I84540,I84368,I84475);
nor I_4819 (I84316,I84419,I84540);
DFFARX1 I_4820 (I320049,I2595,I84342,I84580,);
DFFARX1 I_4821 (I84580,I2595,I84342,I84597,);
not I_4822 (I84605,I84597);
not I_4823 (I84622,I84580);
nand I_4824 (I84319,I84622,I84441);
nand I_4825 (I84653,I320049,I320055);
and I_4826 (I84670,I84653,I320067);
DFFARX1 I_4827 (I84670,I2595,I84342,I84696,);
nor I_4828 (I84704,I84696,I84368);
DFFARX1 I_4829 (I84704,I2595,I84342,I84307,);
DFFARX1 I_4830 (I84696,I2595,I84342,I84325,);
nor I_4831 (I84749,I320058,I320055);
not I_4832 (I84766,I84749);
nor I_4833 (I84328,I84605,I84766);
nand I_4834 (I84313,I84622,I84766);
nor I_4835 (I84322,I84368,I84749);
DFFARX1 I_4836 (I84749,I2595,I84342,I84331,);
not I_4837 (I84869,I2602);
DFFARX1 I_4838 (I249873,I2595,I84869,I84895,);
nand I_4839 (I84903,I249876,I249870);
and I_4840 (I84920,I84903,I249882);
DFFARX1 I_4841 (I84920,I2595,I84869,I84946,);
nor I_4842 (I84837,I84946,I84895);
not I_4843 (I84968,I84946);
DFFARX1 I_4844 (I249885,I2595,I84869,I84994,);
nand I_4845 (I85002,I84994,I249876);
not I_4846 (I85019,I85002);
DFFARX1 I_4847 (I85019,I2595,I84869,I85045,);
not I_4848 (I84861,I85045);
nor I_4849 (I85067,I84895,I85002);
nor I_4850 (I84843,I84946,I85067);
DFFARX1 I_4851 (I249888,I2595,I84869,I85107,);
DFFARX1 I_4852 (I85107,I2595,I84869,I85124,);
not I_4853 (I85132,I85124);
not I_4854 (I85149,I85107);
nand I_4855 (I84846,I85149,I84968);
nand I_4856 (I85180,I249870,I249879);
and I_4857 (I85197,I85180,I249873);
DFFARX1 I_4858 (I85197,I2595,I84869,I85223,);
nor I_4859 (I85231,I85223,I84895);
DFFARX1 I_4860 (I85231,I2595,I84869,I84834,);
DFFARX1 I_4861 (I85223,I2595,I84869,I84852,);
nor I_4862 (I85276,I249891,I249879);
not I_4863 (I85293,I85276);
nor I_4864 (I84855,I85132,I85293);
nand I_4865 (I84840,I85149,I85293);
nor I_4866 (I84849,I84895,I85276);
DFFARX1 I_4867 (I85276,I2595,I84869,I84858,);
not I_4868 (I85396,I2602);
DFFARX1 I_4869 (I210204,I2595,I85396,I85422,);
nand I_4870 (I85430,I210195,I210210);
and I_4871 (I85447,I85430,I210216);
DFFARX1 I_4872 (I85447,I2595,I85396,I85473,);
nor I_4873 (I85364,I85473,I85422);
not I_4874 (I85495,I85473);
DFFARX1 I_4875 (I210201,I2595,I85396,I85521,);
nand I_4876 (I85529,I85521,I210195);
not I_4877 (I85546,I85529);
DFFARX1 I_4878 (I85546,I2595,I85396,I85572,);
not I_4879 (I85388,I85572);
nor I_4880 (I85594,I85422,I85529);
nor I_4881 (I85370,I85473,I85594);
DFFARX1 I_4882 (I210198,I2595,I85396,I85634,);
DFFARX1 I_4883 (I85634,I2595,I85396,I85651,);
not I_4884 (I85659,I85651);
not I_4885 (I85676,I85634);
nand I_4886 (I85373,I85676,I85495);
nand I_4887 (I85707,I210192,I210207);
and I_4888 (I85724,I85707,I210192);
DFFARX1 I_4889 (I85724,I2595,I85396,I85750,);
nor I_4890 (I85758,I85750,I85422);
DFFARX1 I_4891 (I85758,I2595,I85396,I85361,);
DFFARX1 I_4892 (I85750,I2595,I85396,I85379,);
nor I_4893 (I85803,I210213,I210207);
not I_4894 (I85820,I85803);
nor I_4895 (I85382,I85659,I85820);
nand I_4896 (I85367,I85676,I85820);
nor I_4897 (I85376,I85422,I85803);
DFFARX1 I_4898 (I85803,I2595,I85396,I85385,);
not I_4899 (I85923,I2602);
DFFARX1 I_4900 (I31355,I2595,I85923,I85949,);
nand I_4901 (I85957,I31367,I31376);
and I_4902 (I85974,I85957,I31355);
DFFARX1 I_4903 (I85974,I2595,I85923,I86000,);
nor I_4904 (I85891,I86000,I85949);
not I_4905 (I86022,I86000);
DFFARX1 I_4906 (I31370,I2595,I85923,I86048,);
nand I_4907 (I86056,I86048,I31358);
not I_4908 (I86073,I86056);
DFFARX1 I_4909 (I86073,I2595,I85923,I86099,);
not I_4910 (I85915,I86099);
nor I_4911 (I86121,I85949,I86056);
nor I_4912 (I85897,I86000,I86121);
DFFARX1 I_4913 (I31361,I2595,I85923,I86161,);
DFFARX1 I_4914 (I86161,I2595,I85923,I86178,);
not I_4915 (I86186,I86178);
not I_4916 (I86203,I86161);
nand I_4917 (I85900,I86203,I86022);
nand I_4918 (I86234,I31352,I31352);
and I_4919 (I86251,I86234,I31364);
DFFARX1 I_4920 (I86251,I2595,I85923,I86277,);
nor I_4921 (I86285,I86277,I85949);
DFFARX1 I_4922 (I86285,I2595,I85923,I85888,);
DFFARX1 I_4923 (I86277,I2595,I85923,I85906,);
nor I_4924 (I86330,I31373,I31352);
not I_4925 (I86347,I86330);
nor I_4926 (I85909,I86186,I86347);
nand I_4927 (I85894,I86203,I86347);
nor I_4928 (I85903,I85949,I86330);
DFFARX1 I_4929 (I86330,I2595,I85923,I85912,);
not I_4930 (I86450,I2602);
DFFARX1 I_4931 (I203268,I2595,I86450,I86476,);
nand I_4932 (I86484,I203259,I203274);
and I_4933 (I86501,I86484,I203280);
DFFARX1 I_4934 (I86501,I2595,I86450,I86527,);
nor I_4935 (I86418,I86527,I86476);
not I_4936 (I86549,I86527);
DFFARX1 I_4937 (I203265,I2595,I86450,I86575,);
nand I_4938 (I86583,I86575,I203259);
not I_4939 (I86600,I86583);
DFFARX1 I_4940 (I86600,I2595,I86450,I86626,);
not I_4941 (I86442,I86626);
nor I_4942 (I86648,I86476,I86583);
nor I_4943 (I86424,I86527,I86648);
DFFARX1 I_4944 (I203262,I2595,I86450,I86688,);
DFFARX1 I_4945 (I86688,I2595,I86450,I86705,);
not I_4946 (I86713,I86705);
not I_4947 (I86730,I86688);
nand I_4948 (I86427,I86730,I86549);
nand I_4949 (I86761,I203256,I203271);
and I_4950 (I86778,I86761,I203256);
DFFARX1 I_4951 (I86778,I2595,I86450,I86804,);
nor I_4952 (I86812,I86804,I86476);
DFFARX1 I_4953 (I86812,I2595,I86450,I86415,);
DFFARX1 I_4954 (I86804,I2595,I86450,I86433,);
nor I_4955 (I86857,I203277,I203271);
not I_4956 (I86874,I86857);
nor I_4957 (I86436,I86713,I86874);
nand I_4958 (I86421,I86730,I86874);
nor I_4959 (I86430,I86476,I86857);
DFFARX1 I_4960 (I86857,I2595,I86450,I86439,);
not I_4961 (I86977,I2602);
DFFARX1 I_4962 (I36625,I2595,I86977,I87003,);
nand I_4963 (I87011,I36637,I36646);
and I_4964 (I87028,I87011,I36625);
DFFARX1 I_4965 (I87028,I2595,I86977,I87054,);
nor I_4966 (I86945,I87054,I87003);
not I_4967 (I87076,I87054);
DFFARX1 I_4968 (I36640,I2595,I86977,I87102,);
nand I_4969 (I87110,I87102,I36628);
not I_4970 (I87127,I87110);
DFFARX1 I_4971 (I87127,I2595,I86977,I87153,);
not I_4972 (I86969,I87153);
nor I_4973 (I87175,I87003,I87110);
nor I_4974 (I86951,I87054,I87175);
DFFARX1 I_4975 (I36631,I2595,I86977,I87215,);
DFFARX1 I_4976 (I87215,I2595,I86977,I87232,);
not I_4977 (I87240,I87232);
not I_4978 (I87257,I87215);
nand I_4979 (I86954,I87257,I87076);
nand I_4980 (I87288,I36622,I36622);
and I_4981 (I87305,I87288,I36634);
DFFARX1 I_4982 (I87305,I2595,I86977,I87331,);
nor I_4983 (I87339,I87331,I87003);
DFFARX1 I_4984 (I87339,I2595,I86977,I86942,);
DFFARX1 I_4985 (I87331,I2595,I86977,I86960,);
nor I_4986 (I87384,I36643,I36622);
not I_4987 (I87401,I87384);
nor I_4988 (I86963,I87240,I87401);
nand I_4989 (I86948,I87257,I87401);
nor I_4990 (I86957,I87003,I87384);
DFFARX1 I_4991 (I87384,I2595,I86977,I86966,);
not I_4992 (I87504,I2602);
DFFARX1 I_4993 (I381284,I2595,I87504,I87530,);
nand I_4994 (I87538,I381263,I381263);
and I_4995 (I87555,I87538,I381290);
DFFARX1 I_4996 (I87555,I2595,I87504,I87581,);
nor I_4997 (I87472,I87581,I87530);
not I_4998 (I87603,I87581);
DFFARX1 I_4999 (I381278,I2595,I87504,I87629,);
nand I_5000 (I87637,I87629,I381281);
not I_5001 (I87654,I87637);
DFFARX1 I_5002 (I87654,I2595,I87504,I87680,);
not I_5003 (I87496,I87680);
nor I_5004 (I87702,I87530,I87637);
nor I_5005 (I87478,I87581,I87702);
DFFARX1 I_5006 (I381272,I2595,I87504,I87742,);
DFFARX1 I_5007 (I87742,I2595,I87504,I87759,);
not I_5008 (I87767,I87759);
not I_5009 (I87784,I87742);
nand I_5010 (I87481,I87784,I87603);
nand I_5011 (I87815,I381269,I381266);
and I_5012 (I87832,I87815,I381287);
DFFARX1 I_5013 (I87832,I2595,I87504,I87858,);
nor I_5014 (I87866,I87858,I87530);
DFFARX1 I_5015 (I87866,I2595,I87504,I87469,);
DFFARX1 I_5016 (I87858,I2595,I87504,I87487,);
nor I_5017 (I87911,I381275,I381266);
not I_5018 (I87928,I87911);
nor I_5019 (I87490,I87767,I87928);
nand I_5020 (I87475,I87784,I87928);
nor I_5021 (I87484,I87530,I87911);
DFFARX1 I_5022 (I87911,I2595,I87504,I87493,);
not I_5023 (I88031,I2602);
DFFARX1 I_5024 (I149318,I2595,I88031,I88057,);
nand I_5025 (I88065,I149318,I149330);
and I_5026 (I88082,I88065,I149315);
DFFARX1 I_5027 (I88082,I2595,I88031,I88108,);
nor I_5028 (I87999,I88108,I88057);
not I_5029 (I88130,I88108);
DFFARX1 I_5030 (I149339,I2595,I88031,I88156,);
nand I_5031 (I88164,I88156,I149336);
not I_5032 (I88181,I88164);
DFFARX1 I_5033 (I88181,I2595,I88031,I88207,);
not I_5034 (I88023,I88207);
nor I_5035 (I88229,I88057,I88164);
nor I_5036 (I88005,I88108,I88229);
DFFARX1 I_5037 (I149327,I2595,I88031,I88269,);
DFFARX1 I_5038 (I88269,I2595,I88031,I88286,);
not I_5039 (I88294,I88286);
not I_5040 (I88311,I88269);
nand I_5041 (I88008,I88311,I88130);
nand I_5042 (I88342,I149315,I149324);
and I_5043 (I88359,I88342,I149333);
DFFARX1 I_5044 (I88359,I2595,I88031,I88385,);
nor I_5045 (I88393,I88385,I88057);
DFFARX1 I_5046 (I88393,I2595,I88031,I87996,);
DFFARX1 I_5047 (I88385,I2595,I88031,I88014,);
nor I_5048 (I88438,I149321,I149324);
not I_5049 (I88455,I88438);
nor I_5050 (I88017,I88294,I88455);
nand I_5051 (I88002,I88311,I88455);
nor I_5052 (I88011,I88057,I88438);
DFFARX1 I_5053 (I88438,I2595,I88031,I88020,);
not I_5054 (I88558,I2602);
DFFARX1 I_5055 (I41895,I2595,I88558,I88584,);
nand I_5056 (I88592,I41907,I41916);
and I_5057 (I88609,I88592,I41895);
DFFARX1 I_5058 (I88609,I2595,I88558,I88635,);
nor I_5059 (I88526,I88635,I88584);
not I_5060 (I88657,I88635);
DFFARX1 I_5061 (I41910,I2595,I88558,I88683,);
nand I_5062 (I88691,I88683,I41898);
not I_5063 (I88708,I88691);
DFFARX1 I_5064 (I88708,I2595,I88558,I88734,);
not I_5065 (I88550,I88734);
nor I_5066 (I88756,I88584,I88691);
nor I_5067 (I88532,I88635,I88756);
DFFARX1 I_5068 (I41901,I2595,I88558,I88796,);
DFFARX1 I_5069 (I88796,I2595,I88558,I88813,);
not I_5070 (I88821,I88813);
not I_5071 (I88838,I88796);
nand I_5072 (I88535,I88838,I88657);
nand I_5073 (I88869,I41892,I41892);
and I_5074 (I88886,I88869,I41904);
DFFARX1 I_5075 (I88886,I2595,I88558,I88912,);
nor I_5076 (I88920,I88912,I88584);
DFFARX1 I_5077 (I88920,I2595,I88558,I88523,);
DFFARX1 I_5078 (I88912,I2595,I88558,I88541,);
nor I_5079 (I88965,I41913,I41892);
not I_5080 (I88982,I88965);
nor I_5081 (I88544,I88821,I88982);
nand I_5082 (I88529,I88838,I88982);
nor I_5083 (I88538,I88584,I88965);
DFFARX1 I_5084 (I88965,I2595,I88558,I88547,);
not I_5085 (I89085,I2602);
DFFARX1 I_5086 (I322936,I2595,I89085,I89111,);
nand I_5087 (I89119,I322951,I322936);
and I_5088 (I89136,I89119,I322954);
DFFARX1 I_5089 (I89136,I2595,I89085,I89162,);
nor I_5090 (I89053,I89162,I89111);
not I_5091 (I89184,I89162);
DFFARX1 I_5092 (I322960,I2595,I89085,I89210,);
nand I_5093 (I89218,I89210,I322942);
not I_5094 (I89235,I89218);
DFFARX1 I_5095 (I89235,I2595,I89085,I89261,);
not I_5096 (I89077,I89261);
nor I_5097 (I89283,I89111,I89218);
nor I_5098 (I89059,I89162,I89283);
DFFARX1 I_5099 (I322939,I2595,I89085,I89323,);
DFFARX1 I_5100 (I89323,I2595,I89085,I89340,);
not I_5101 (I89348,I89340);
not I_5102 (I89365,I89323);
nand I_5103 (I89062,I89365,I89184);
nand I_5104 (I89396,I322939,I322945);
and I_5105 (I89413,I89396,I322957);
DFFARX1 I_5106 (I89413,I2595,I89085,I89439,);
nor I_5107 (I89447,I89439,I89111);
DFFARX1 I_5108 (I89447,I2595,I89085,I89050,);
DFFARX1 I_5109 (I89439,I2595,I89085,I89068,);
nor I_5110 (I89492,I322948,I322945);
not I_5111 (I89509,I89492);
nor I_5112 (I89071,I89348,I89509);
nand I_5113 (I89056,I89365,I89509);
nor I_5114 (I89065,I89111,I89492);
DFFARX1 I_5115 (I89492,I2595,I89085,I89074,);
not I_5116 (I89612,I2602);
DFFARX1 I_5117 (I25558,I2595,I89612,I89638,);
nand I_5118 (I89646,I25570,I25579);
and I_5119 (I89663,I89646,I25558);
DFFARX1 I_5120 (I89663,I2595,I89612,I89689,);
nor I_5121 (I89580,I89689,I89638);
not I_5122 (I89711,I89689);
DFFARX1 I_5123 (I25573,I2595,I89612,I89737,);
nand I_5124 (I89745,I89737,I25561);
not I_5125 (I89762,I89745);
DFFARX1 I_5126 (I89762,I2595,I89612,I89788,);
not I_5127 (I89604,I89788);
nor I_5128 (I89810,I89638,I89745);
nor I_5129 (I89586,I89689,I89810);
DFFARX1 I_5130 (I25564,I2595,I89612,I89850,);
DFFARX1 I_5131 (I89850,I2595,I89612,I89867,);
not I_5132 (I89875,I89867);
not I_5133 (I89892,I89850);
nand I_5134 (I89589,I89892,I89711);
nand I_5135 (I89923,I25555,I25555);
and I_5136 (I89940,I89923,I25567);
DFFARX1 I_5137 (I89940,I2595,I89612,I89966,);
nor I_5138 (I89974,I89966,I89638);
DFFARX1 I_5139 (I89974,I2595,I89612,I89577,);
DFFARX1 I_5140 (I89966,I2595,I89612,I89595,);
nor I_5141 (I90019,I25576,I25555);
not I_5142 (I90036,I90019);
nor I_5143 (I89598,I89875,I90036);
nand I_5144 (I89583,I89892,I90036);
nor I_5145 (I89592,I89638,I90019);
DFFARX1 I_5146 (I90019,I2595,I89612,I89601,);
not I_5147 (I90139,I2602);
DFFARX1 I_5148 (I320624,I2595,I90139,I90165,);
nand I_5149 (I90173,I320639,I320624);
and I_5150 (I90190,I90173,I320642);
DFFARX1 I_5151 (I90190,I2595,I90139,I90216,);
nor I_5152 (I90107,I90216,I90165);
not I_5153 (I90238,I90216);
DFFARX1 I_5154 (I320648,I2595,I90139,I90264,);
nand I_5155 (I90272,I90264,I320630);
not I_5156 (I90289,I90272);
DFFARX1 I_5157 (I90289,I2595,I90139,I90315,);
not I_5158 (I90131,I90315);
nor I_5159 (I90337,I90165,I90272);
nor I_5160 (I90113,I90216,I90337);
DFFARX1 I_5161 (I320627,I2595,I90139,I90377,);
DFFARX1 I_5162 (I90377,I2595,I90139,I90394,);
not I_5163 (I90402,I90394);
not I_5164 (I90419,I90377);
nand I_5165 (I90116,I90419,I90238);
nand I_5166 (I90450,I320627,I320633);
and I_5167 (I90467,I90450,I320645);
DFFARX1 I_5168 (I90467,I2595,I90139,I90493,);
nor I_5169 (I90501,I90493,I90165);
DFFARX1 I_5170 (I90501,I2595,I90139,I90104,);
DFFARX1 I_5171 (I90493,I2595,I90139,I90122,);
nor I_5172 (I90546,I320636,I320633);
not I_5173 (I90563,I90546);
nor I_5174 (I90125,I90402,I90563);
nand I_5175 (I90110,I90419,I90563);
nor I_5176 (I90119,I90165,I90546);
DFFARX1 I_5177 (I90546,I2595,I90139,I90128,);
not I_5178 (I90666,I2602);
DFFARX1 I_5179 (I249346,I2595,I90666,I90692,);
nand I_5180 (I90700,I249349,I249343);
and I_5181 (I90717,I90700,I249355);
DFFARX1 I_5182 (I90717,I2595,I90666,I90743,);
nor I_5183 (I90634,I90743,I90692);
not I_5184 (I90765,I90743);
DFFARX1 I_5185 (I249358,I2595,I90666,I90791,);
nand I_5186 (I90799,I90791,I249349);
not I_5187 (I90816,I90799);
DFFARX1 I_5188 (I90816,I2595,I90666,I90842,);
not I_5189 (I90658,I90842);
nor I_5190 (I90864,I90692,I90799);
nor I_5191 (I90640,I90743,I90864);
DFFARX1 I_5192 (I249361,I2595,I90666,I90904,);
DFFARX1 I_5193 (I90904,I2595,I90666,I90921,);
not I_5194 (I90929,I90921);
not I_5195 (I90946,I90904);
nand I_5196 (I90643,I90946,I90765);
nand I_5197 (I90977,I249343,I249352);
and I_5198 (I90994,I90977,I249346);
DFFARX1 I_5199 (I90994,I2595,I90666,I91020,);
nor I_5200 (I91028,I91020,I90692);
DFFARX1 I_5201 (I91028,I2595,I90666,I90631,);
DFFARX1 I_5202 (I91020,I2595,I90666,I90649,);
nor I_5203 (I91073,I249364,I249352);
not I_5204 (I91090,I91073);
nor I_5205 (I90652,I90929,I91090);
nand I_5206 (I90637,I90946,I91090);
nor I_5207 (I90646,I90692,I91073);
DFFARX1 I_5208 (I91073,I2595,I90666,I90655,);
not I_5209 (I91193,I2602);
DFFARX1 I_5210 (I139909,I2595,I91193,I91219,);
nand I_5211 (I91227,I139921,I139900);
and I_5212 (I91244,I91227,I139924);
DFFARX1 I_5213 (I91244,I2595,I91193,I91270,);
nor I_5214 (I91161,I91270,I91219);
not I_5215 (I91292,I91270);
DFFARX1 I_5216 (I139915,I2595,I91193,I91318,);
nand I_5217 (I91326,I91318,I139897);
not I_5218 (I91343,I91326);
DFFARX1 I_5219 (I91343,I2595,I91193,I91369,);
not I_5220 (I91185,I91369);
nor I_5221 (I91391,I91219,I91326);
nor I_5222 (I91167,I91270,I91391);
DFFARX1 I_5223 (I139912,I2595,I91193,I91431,);
DFFARX1 I_5224 (I91431,I2595,I91193,I91448,);
not I_5225 (I91456,I91448);
not I_5226 (I91473,I91431);
nand I_5227 (I91170,I91473,I91292);
nand I_5228 (I91504,I139897,I139903);
and I_5229 (I91521,I91504,I139906);
DFFARX1 I_5230 (I91521,I2595,I91193,I91547,);
nor I_5231 (I91555,I91547,I91219);
DFFARX1 I_5232 (I91555,I2595,I91193,I91158,);
DFFARX1 I_5233 (I91547,I2595,I91193,I91176,);
nor I_5234 (I91600,I139918,I139903);
not I_5235 (I91617,I91600);
nor I_5236 (I91179,I91456,I91617);
nand I_5237 (I91164,I91473,I91617);
nor I_5238 (I91173,I91219,I91600);
DFFARX1 I_5239 (I91600,I2595,I91193,I91182,);
not I_5240 (I91720,I2602);
DFFARX1 I_5241 (I262844,I2595,I91720,I91746,);
nand I_5242 (I91754,I262841,I262859);
and I_5243 (I91771,I91754,I262850);
DFFARX1 I_5244 (I91771,I2595,I91720,I91797,);
nor I_5245 (I91688,I91797,I91746);
not I_5246 (I91819,I91797);
DFFARX1 I_5247 (I262865,I2595,I91720,I91845,);
nand I_5248 (I91853,I91845,I262847);
not I_5249 (I91870,I91853);
DFFARX1 I_5250 (I91870,I2595,I91720,I91896,);
not I_5251 (I91712,I91896);
nor I_5252 (I91918,I91746,I91853);
nor I_5253 (I91694,I91797,I91918);
DFFARX1 I_5254 (I262853,I2595,I91720,I91958,);
DFFARX1 I_5255 (I91958,I2595,I91720,I91975,);
not I_5256 (I91983,I91975);
not I_5257 (I92000,I91958);
nand I_5258 (I91697,I92000,I91819);
nand I_5259 (I92031,I262841,I262868);
and I_5260 (I92048,I92031,I262856);
DFFARX1 I_5261 (I92048,I2595,I91720,I92074,);
nor I_5262 (I92082,I92074,I91746);
DFFARX1 I_5263 (I92082,I2595,I91720,I91685,);
DFFARX1 I_5264 (I92074,I2595,I91720,I91703,);
nor I_5265 (I92127,I262862,I262868);
not I_5266 (I92144,I92127);
nor I_5267 (I91706,I91983,I92144);
nand I_5268 (I91691,I92000,I92144);
nor I_5269 (I91700,I91746,I92127);
DFFARX1 I_5270 (I92127,I2595,I91720,I91709,);
not I_5271 (I92247,I2602);
DFFARX1 I_5272 (I234590,I2595,I92247,I92273,);
nand I_5273 (I92281,I234593,I234587);
and I_5274 (I92298,I92281,I234599);
DFFARX1 I_5275 (I92298,I2595,I92247,I92324,);
nor I_5276 (I92215,I92324,I92273);
not I_5277 (I92346,I92324);
DFFARX1 I_5278 (I234602,I2595,I92247,I92372,);
nand I_5279 (I92380,I92372,I234593);
not I_5280 (I92397,I92380);
DFFARX1 I_5281 (I92397,I2595,I92247,I92423,);
not I_5282 (I92239,I92423);
nor I_5283 (I92445,I92273,I92380);
nor I_5284 (I92221,I92324,I92445);
DFFARX1 I_5285 (I234605,I2595,I92247,I92485,);
DFFARX1 I_5286 (I92485,I2595,I92247,I92502,);
not I_5287 (I92510,I92502);
not I_5288 (I92527,I92485);
nand I_5289 (I92224,I92527,I92346);
nand I_5290 (I92558,I234587,I234596);
and I_5291 (I92575,I92558,I234590);
DFFARX1 I_5292 (I92575,I2595,I92247,I92601,);
nor I_5293 (I92609,I92601,I92273);
DFFARX1 I_5294 (I92609,I2595,I92247,I92212,);
DFFARX1 I_5295 (I92601,I2595,I92247,I92230,);
nor I_5296 (I92654,I234608,I234596);
not I_5297 (I92671,I92654);
nor I_5298 (I92233,I92510,I92671);
nand I_5299 (I92218,I92527,I92671);
nor I_5300 (I92227,I92273,I92654);
DFFARX1 I_5301 (I92654,I2595,I92247,I92236,);
not I_5302 (I92774,I2602);
DFFARX1 I_5303 (I206736,I2595,I92774,I92800,);
nand I_5304 (I92808,I206727,I206742);
and I_5305 (I92825,I92808,I206748);
DFFARX1 I_5306 (I92825,I2595,I92774,I92851,);
nor I_5307 (I92742,I92851,I92800);
not I_5308 (I92873,I92851);
DFFARX1 I_5309 (I206733,I2595,I92774,I92899,);
nand I_5310 (I92907,I92899,I206727);
not I_5311 (I92924,I92907);
DFFARX1 I_5312 (I92924,I2595,I92774,I92950,);
not I_5313 (I92766,I92950);
nor I_5314 (I92972,I92800,I92907);
nor I_5315 (I92748,I92851,I92972);
DFFARX1 I_5316 (I206730,I2595,I92774,I93012,);
DFFARX1 I_5317 (I93012,I2595,I92774,I93029,);
not I_5318 (I93037,I93029);
not I_5319 (I93054,I93012);
nand I_5320 (I92751,I93054,I92873);
nand I_5321 (I93085,I206724,I206739);
and I_5322 (I93102,I93085,I206724);
DFFARX1 I_5323 (I93102,I2595,I92774,I93128,);
nor I_5324 (I93136,I93128,I92800);
DFFARX1 I_5325 (I93136,I2595,I92774,I92739,);
DFFARX1 I_5326 (I93128,I2595,I92774,I92757,);
nor I_5327 (I93181,I206745,I206739);
not I_5328 (I93198,I93181);
nor I_5329 (I92760,I93037,I93198);
nand I_5330 (I92745,I93054,I93198);
nor I_5331 (I92754,I92800,I93181);
DFFARX1 I_5332 (I93181,I2595,I92774,I92763,);
not I_5333 (I93301,I2602);
DFFARX1 I_5334 (I209626,I2595,I93301,I93327,);
nand I_5335 (I93335,I209617,I209632);
and I_5336 (I93352,I93335,I209638);
DFFARX1 I_5337 (I93352,I2595,I93301,I93378,);
nor I_5338 (I93269,I93378,I93327);
not I_5339 (I93400,I93378);
DFFARX1 I_5340 (I209623,I2595,I93301,I93426,);
nand I_5341 (I93434,I93426,I209617);
not I_5342 (I93451,I93434);
DFFARX1 I_5343 (I93451,I2595,I93301,I93477,);
not I_5344 (I93293,I93477);
nor I_5345 (I93499,I93327,I93434);
nor I_5346 (I93275,I93378,I93499);
DFFARX1 I_5347 (I209620,I2595,I93301,I93539,);
DFFARX1 I_5348 (I93539,I2595,I93301,I93556,);
not I_5349 (I93564,I93556);
not I_5350 (I93581,I93539);
nand I_5351 (I93278,I93581,I93400);
nand I_5352 (I93612,I209614,I209629);
and I_5353 (I93629,I93612,I209614);
DFFARX1 I_5354 (I93629,I2595,I93301,I93655,);
nor I_5355 (I93663,I93655,I93327);
DFFARX1 I_5356 (I93663,I2595,I93301,I93266,);
DFFARX1 I_5357 (I93655,I2595,I93301,I93284,);
nor I_5358 (I93708,I209635,I209629);
not I_5359 (I93725,I93708);
nor I_5360 (I93287,I93564,I93725);
nand I_5361 (I93272,I93581,I93725);
nor I_5362 (I93281,I93327,I93708);
DFFARX1 I_5363 (I93708,I2595,I93301,I93290,);
not I_5364 (I93828,I2602);
DFFARX1 I_5365 (I204424,I2595,I93828,I93854,);
nand I_5366 (I93862,I204415,I204430);
and I_5367 (I93879,I93862,I204436);
DFFARX1 I_5368 (I93879,I2595,I93828,I93905,);
nor I_5369 (I93796,I93905,I93854);
not I_5370 (I93927,I93905);
DFFARX1 I_5371 (I204421,I2595,I93828,I93953,);
nand I_5372 (I93961,I93953,I204415);
not I_5373 (I93978,I93961);
DFFARX1 I_5374 (I93978,I2595,I93828,I94004,);
not I_5375 (I93820,I94004);
nor I_5376 (I94026,I93854,I93961);
nor I_5377 (I93802,I93905,I94026);
DFFARX1 I_5378 (I204418,I2595,I93828,I94066,);
DFFARX1 I_5379 (I94066,I2595,I93828,I94083,);
not I_5380 (I94091,I94083);
not I_5381 (I94108,I94066);
nand I_5382 (I93805,I94108,I93927);
nand I_5383 (I94139,I204412,I204427);
and I_5384 (I94156,I94139,I204412);
DFFARX1 I_5385 (I94156,I2595,I93828,I94182,);
nor I_5386 (I94190,I94182,I93854);
DFFARX1 I_5387 (I94190,I2595,I93828,I93793,);
DFFARX1 I_5388 (I94182,I2595,I93828,I93811,);
nor I_5389 (I94235,I204433,I204427);
not I_5390 (I94252,I94235);
nor I_5391 (I93814,I94091,I94252);
nand I_5392 (I93799,I94108,I94252);
nor I_5393 (I93808,I93854,I94235);
DFFARX1 I_5394 (I94235,I2595,I93828,I93817,);
not I_5395 (I94355,I2602);
DFFARX1 I_5396 (I387234,I2595,I94355,I94381,);
nand I_5397 (I94389,I387213,I387213);
and I_5398 (I94406,I94389,I387240);
DFFARX1 I_5399 (I94406,I2595,I94355,I94432,);
nor I_5400 (I94323,I94432,I94381);
not I_5401 (I94454,I94432);
DFFARX1 I_5402 (I387228,I2595,I94355,I94480,);
nand I_5403 (I94488,I94480,I387231);
not I_5404 (I94505,I94488);
DFFARX1 I_5405 (I94505,I2595,I94355,I94531,);
not I_5406 (I94347,I94531);
nor I_5407 (I94553,I94381,I94488);
nor I_5408 (I94329,I94432,I94553);
DFFARX1 I_5409 (I387222,I2595,I94355,I94593,);
DFFARX1 I_5410 (I94593,I2595,I94355,I94610,);
not I_5411 (I94618,I94610);
not I_5412 (I94635,I94593);
nand I_5413 (I94332,I94635,I94454);
nand I_5414 (I94666,I387219,I387216);
and I_5415 (I94683,I94666,I387237);
DFFARX1 I_5416 (I94683,I2595,I94355,I94709,);
nor I_5417 (I94717,I94709,I94381);
DFFARX1 I_5418 (I94717,I2595,I94355,I94320,);
DFFARX1 I_5419 (I94709,I2595,I94355,I94338,);
nor I_5420 (I94762,I387225,I387216);
not I_5421 (I94779,I94762);
nor I_5422 (I94341,I94618,I94779);
nand I_5423 (I94326,I94635,I94779);
nor I_5424 (I94335,I94381,I94762);
DFFARX1 I_5425 (I94762,I2595,I94355,I94344,);
not I_5426 (I94882,I2602);
DFFARX1 I_5427 (I242495,I2595,I94882,I94908,);
nand I_5428 (I94916,I242498,I242492);
and I_5429 (I94933,I94916,I242504);
DFFARX1 I_5430 (I94933,I2595,I94882,I94959,);
nor I_5431 (I94850,I94959,I94908);
not I_5432 (I94981,I94959);
DFFARX1 I_5433 (I242507,I2595,I94882,I95007,);
nand I_5434 (I95015,I95007,I242498);
not I_5435 (I95032,I95015);
DFFARX1 I_5436 (I95032,I2595,I94882,I95058,);
not I_5437 (I94874,I95058);
nor I_5438 (I95080,I94908,I95015);
nor I_5439 (I94856,I94959,I95080);
DFFARX1 I_5440 (I242510,I2595,I94882,I95120,);
DFFARX1 I_5441 (I95120,I2595,I94882,I95137,);
not I_5442 (I95145,I95137);
not I_5443 (I95162,I95120);
nand I_5444 (I94859,I95162,I94981);
nand I_5445 (I95193,I242492,I242501);
and I_5446 (I95210,I95193,I242495);
DFFARX1 I_5447 (I95210,I2595,I94882,I95236,);
nor I_5448 (I95244,I95236,I94908);
DFFARX1 I_5449 (I95244,I2595,I94882,I94847,);
DFFARX1 I_5450 (I95236,I2595,I94882,I94865,);
nor I_5451 (I95289,I242513,I242501);
not I_5452 (I95306,I95289);
nor I_5453 (I94868,I95145,I95306);
nand I_5454 (I94853,I95162,I95306);
nor I_5455 (I94862,I94908,I95289);
DFFARX1 I_5456 (I95289,I2595,I94882,I94871,);
not I_5457 (I95409,I2602);
DFFARX1 I_5458 (I63363,I2595,I95409,I95435,);
nand I_5459 (I95443,I63363,I63369);
and I_5460 (I95460,I95443,I63387);
DFFARX1 I_5461 (I95460,I2595,I95409,I95486,);
nor I_5462 (I95377,I95486,I95435);
not I_5463 (I95508,I95486);
DFFARX1 I_5464 (I63375,I2595,I95409,I95534,);
nand I_5465 (I95542,I95534,I63372);
not I_5466 (I95559,I95542);
DFFARX1 I_5467 (I95559,I2595,I95409,I95585,);
not I_5468 (I95401,I95585);
nor I_5469 (I95607,I95435,I95542);
nor I_5470 (I95383,I95486,I95607);
DFFARX1 I_5471 (I63381,I2595,I95409,I95647,);
DFFARX1 I_5472 (I95647,I2595,I95409,I95664,);
not I_5473 (I95672,I95664);
not I_5474 (I95689,I95647);
nand I_5475 (I95386,I95689,I95508);
nand I_5476 (I95720,I63366,I63366);
and I_5477 (I95737,I95720,I63378);
DFFARX1 I_5478 (I95737,I2595,I95409,I95763,);
nor I_5479 (I95771,I95763,I95435);
DFFARX1 I_5480 (I95771,I2595,I95409,I95374,);
DFFARX1 I_5481 (I95763,I2595,I95409,I95392,);
nor I_5482 (I95816,I63384,I63366);
not I_5483 (I95833,I95816);
nor I_5484 (I95395,I95672,I95833);
nand I_5485 (I95380,I95689,I95833);
nor I_5486 (I95389,I95435,I95816);
DFFARX1 I_5487 (I95816,I2595,I95409,I95398,);
not I_5488 (I95936,I2602);
DFFARX1 I_5489 (I115973,I2595,I95936,I95962,);
nand I_5490 (I95970,I115985,I115964);
and I_5491 (I95987,I95970,I115988);
DFFARX1 I_5492 (I95987,I2595,I95936,I96013,);
nor I_5493 (I95904,I96013,I95962);
not I_5494 (I96035,I96013);
DFFARX1 I_5495 (I115979,I2595,I95936,I96061,);
nand I_5496 (I96069,I96061,I115961);
not I_5497 (I96086,I96069);
DFFARX1 I_5498 (I96086,I2595,I95936,I96112,);
not I_5499 (I95928,I96112);
nor I_5500 (I96134,I95962,I96069);
nor I_5501 (I95910,I96013,I96134);
DFFARX1 I_5502 (I115976,I2595,I95936,I96174,);
DFFARX1 I_5503 (I96174,I2595,I95936,I96191,);
not I_5504 (I96199,I96191);
not I_5505 (I96216,I96174);
nand I_5506 (I95913,I96216,I96035);
nand I_5507 (I96247,I115961,I115967);
and I_5508 (I96264,I96247,I115970);
DFFARX1 I_5509 (I96264,I2595,I95936,I96290,);
nor I_5510 (I96298,I96290,I95962);
DFFARX1 I_5511 (I96298,I2595,I95936,I95901,);
DFFARX1 I_5512 (I96290,I2595,I95936,I95919,);
nor I_5513 (I96343,I115982,I115967);
not I_5514 (I96360,I96343);
nor I_5515 (I95922,I96199,I96360);
nand I_5516 (I95907,I96216,I96360);
nor I_5517 (I95916,I95962,I96343);
DFFARX1 I_5518 (I96343,I2595,I95936,I95925,);
not I_5519 (I96463,I2602);
DFFARX1 I_5520 (I207892,I2595,I96463,I96489,);
nand I_5521 (I96497,I207883,I207898);
and I_5522 (I96514,I96497,I207904);
DFFARX1 I_5523 (I96514,I2595,I96463,I96540,);
nor I_5524 (I96431,I96540,I96489);
not I_5525 (I96562,I96540);
DFFARX1 I_5526 (I207889,I2595,I96463,I96588,);
nand I_5527 (I96596,I96588,I207883);
not I_5528 (I96613,I96596);
DFFARX1 I_5529 (I96613,I2595,I96463,I96639,);
not I_5530 (I96455,I96639);
nor I_5531 (I96661,I96489,I96596);
nor I_5532 (I96437,I96540,I96661);
DFFARX1 I_5533 (I207886,I2595,I96463,I96701,);
DFFARX1 I_5534 (I96701,I2595,I96463,I96718,);
not I_5535 (I96726,I96718);
not I_5536 (I96743,I96701);
nand I_5537 (I96440,I96743,I96562);
nand I_5538 (I96774,I207880,I207895);
and I_5539 (I96791,I96774,I207880);
DFFARX1 I_5540 (I96791,I2595,I96463,I96817,);
nor I_5541 (I96825,I96817,I96489);
DFFARX1 I_5542 (I96825,I2595,I96463,I96428,);
DFFARX1 I_5543 (I96817,I2595,I96463,I96446,);
nor I_5544 (I96870,I207901,I207895);
not I_5545 (I96887,I96870);
nor I_5546 (I96449,I96726,I96887);
nand I_5547 (I96434,I96743,I96887);
nor I_5548 (I96443,I96489,I96870);
DFFARX1 I_5549 (I96870,I2595,I96463,I96452,);
not I_5550 (I96990,I2602);
DFFARX1 I_5551 (I275764,I2595,I96990,I97016,);
nand I_5552 (I97024,I275761,I275779);
and I_5553 (I97041,I97024,I275770);
DFFARX1 I_5554 (I97041,I2595,I96990,I97067,);
nor I_5555 (I96958,I97067,I97016);
not I_5556 (I97089,I97067);
DFFARX1 I_5557 (I275785,I2595,I96990,I97115,);
nand I_5558 (I97123,I97115,I275767);
not I_5559 (I97140,I97123);
DFFARX1 I_5560 (I97140,I2595,I96990,I97166,);
not I_5561 (I96982,I97166);
nor I_5562 (I97188,I97016,I97123);
nor I_5563 (I96964,I97067,I97188);
DFFARX1 I_5564 (I275773,I2595,I96990,I97228,);
DFFARX1 I_5565 (I97228,I2595,I96990,I97245,);
not I_5566 (I97253,I97245);
not I_5567 (I97270,I97228);
nand I_5568 (I96967,I97270,I97089);
nand I_5569 (I97301,I275761,I275788);
and I_5570 (I97318,I97301,I275776);
DFFARX1 I_5571 (I97318,I2595,I96990,I97344,);
nor I_5572 (I97352,I97344,I97016);
DFFARX1 I_5573 (I97352,I2595,I96990,I96955,);
DFFARX1 I_5574 (I97344,I2595,I96990,I96973,);
nor I_5575 (I97397,I275782,I275788);
not I_5576 (I97414,I97397);
nor I_5577 (I96976,I97253,I97414);
nand I_5578 (I96961,I97270,I97414);
nor I_5579 (I96970,I97016,I97397);
DFFARX1 I_5580 (I97397,I2595,I96990,I96979,);
not I_5581 (I97517,I2602);
DFFARX1 I_5582 (I328138,I2595,I97517,I97543,);
nand I_5583 (I97551,I328153,I328138);
and I_5584 (I97568,I97551,I328156);
DFFARX1 I_5585 (I97568,I2595,I97517,I97594,);
nor I_5586 (I97485,I97594,I97543);
not I_5587 (I97616,I97594);
DFFARX1 I_5588 (I328162,I2595,I97517,I97642,);
nand I_5589 (I97650,I97642,I328144);
not I_5590 (I97667,I97650);
DFFARX1 I_5591 (I97667,I2595,I97517,I97693,);
not I_5592 (I97509,I97693);
nor I_5593 (I97715,I97543,I97650);
nor I_5594 (I97491,I97594,I97715);
DFFARX1 I_5595 (I328141,I2595,I97517,I97755,);
DFFARX1 I_5596 (I97755,I2595,I97517,I97772,);
not I_5597 (I97780,I97772);
not I_5598 (I97797,I97755);
nand I_5599 (I97494,I97797,I97616);
nand I_5600 (I97828,I328141,I328147);
and I_5601 (I97845,I97828,I328159);
DFFARX1 I_5602 (I97845,I2595,I97517,I97871,);
nor I_5603 (I97879,I97871,I97543);
DFFARX1 I_5604 (I97879,I2595,I97517,I97482,);
DFFARX1 I_5605 (I97871,I2595,I97517,I97500,);
nor I_5606 (I97924,I328150,I328147);
not I_5607 (I97941,I97924);
nor I_5608 (I97503,I97780,I97941);
nand I_5609 (I97488,I97797,I97941);
nor I_5610 (I97497,I97543,I97924);
DFFARX1 I_5611 (I97924,I2595,I97517,I97506,);
not I_5612 (I98044,I2602);
DFFARX1 I_5613 (I378309,I2595,I98044,I98070,);
nand I_5614 (I98078,I378288,I378288);
and I_5615 (I98095,I98078,I378315);
DFFARX1 I_5616 (I98095,I2595,I98044,I98121,);
nor I_5617 (I98012,I98121,I98070);
not I_5618 (I98143,I98121);
DFFARX1 I_5619 (I378303,I2595,I98044,I98169,);
nand I_5620 (I98177,I98169,I378306);
not I_5621 (I98194,I98177);
DFFARX1 I_5622 (I98194,I2595,I98044,I98220,);
not I_5623 (I98036,I98220);
nor I_5624 (I98242,I98070,I98177);
nor I_5625 (I98018,I98121,I98242);
DFFARX1 I_5626 (I378297,I2595,I98044,I98282,);
DFFARX1 I_5627 (I98282,I2595,I98044,I98299,);
not I_5628 (I98307,I98299);
not I_5629 (I98324,I98282);
nand I_5630 (I98021,I98324,I98143);
nand I_5631 (I98355,I378294,I378291);
and I_5632 (I98372,I98355,I378312);
DFFARX1 I_5633 (I98372,I2595,I98044,I98398,);
nor I_5634 (I98406,I98398,I98070);
DFFARX1 I_5635 (I98406,I2595,I98044,I98009,);
DFFARX1 I_5636 (I98398,I2595,I98044,I98027,);
nor I_5637 (I98451,I378300,I378291);
not I_5638 (I98468,I98451);
nor I_5639 (I98030,I98307,I98468);
nand I_5640 (I98015,I98324,I98468);
nor I_5641 (I98024,I98070,I98451);
DFFARX1 I_5642 (I98451,I2595,I98044,I98033,);
not I_5643 (I98571,I2602);
DFFARX1 I_5644 (I210782,I2595,I98571,I98597,);
nand I_5645 (I98605,I210773,I210788);
and I_5646 (I98622,I98605,I210794);
DFFARX1 I_5647 (I98622,I2595,I98571,I98648,);
nor I_5648 (I98539,I98648,I98597);
not I_5649 (I98670,I98648);
DFFARX1 I_5650 (I210779,I2595,I98571,I98696,);
nand I_5651 (I98704,I98696,I210773);
not I_5652 (I98721,I98704);
DFFARX1 I_5653 (I98721,I2595,I98571,I98747,);
not I_5654 (I98563,I98747);
nor I_5655 (I98769,I98597,I98704);
nor I_5656 (I98545,I98648,I98769);
DFFARX1 I_5657 (I210776,I2595,I98571,I98809,);
DFFARX1 I_5658 (I98809,I2595,I98571,I98826,);
not I_5659 (I98834,I98826);
not I_5660 (I98851,I98809);
nand I_5661 (I98548,I98851,I98670);
nand I_5662 (I98882,I210770,I210785);
and I_5663 (I98899,I98882,I210770);
DFFARX1 I_5664 (I98899,I2595,I98571,I98925,);
nor I_5665 (I98933,I98925,I98597);
DFFARX1 I_5666 (I98933,I2595,I98571,I98536,);
DFFARX1 I_5667 (I98925,I2595,I98571,I98554,);
nor I_5668 (I98978,I210791,I210785);
not I_5669 (I98995,I98978);
nor I_5670 (I98557,I98834,I98995);
nand I_5671 (I98542,I98851,I98995);
nor I_5672 (I98551,I98597,I98978);
DFFARX1 I_5673 (I98978,I2595,I98571,I98560,);
not I_5674 (I99098,I2602);
DFFARX1 I_5675 (I27666,I2595,I99098,I99124,);
nand I_5676 (I99132,I27678,I27687);
and I_5677 (I99149,I99132,I27666);
DFFARX1 I_5678 (I99149,I2595,I99098,I99175,);
nor I_5679 (I99066,I99175,I99124);
not I_5680 (I99197,I99175);
DFFARX1 I_5681 (I27681,I2595,I99098,I99223,);
nand I_5682 (I99231,I99223,I27669);
not I_5683 (I99248,I99231);
DFFARX1 I_5684 (I99248,I2595,I99098,I99274,);
not I_5685 (I99090,I99274);
nor I_5686 (I99296,I99124,I99231);
nor I_5687 (I99072,I99175,I99296);
DFFARX1 I_5688 (I27672,I2595,I99098,I99336,);
DFFARX1 I_5689 (I99336,I2595,I99098,I99353,);
not I_5690 (I99361,I99353);
not I_5691 (I99378,I99336);
nand I_5692 (I99075,I99378,I99197);
nand I_5693 (I99409,I27663,I27663);
and I_5694 (I99426,I99409,I27675);
DFFARX1 I_5695 (I99426,I2595,I99098,I99452,);
nor I_5696 (I99460,I99452,I99124);
DFFARX1 I_5697 (I99460,I2595,I99098,I99063,);
DFFARX1 I_5698 (I99452,I2595,I99098,I99081,);
nor I_5699 (I99505,I27684,I27663);
not I_5700 (I99522,I99505);
nor I_5701 (I99084,I99361,I99522);
nand I_5702 (I99069,I99378,I99522);
nor I_5703 (I99078,I99124,I99505);
DFFARX1 I_5704 (I99505,I2595,I99098,I99087,);
not I_5705 (I99625,I2602);
DFFARX1 I_5706 (I9165,I2595,I99625,I99651,);
nand I_5707 (I99659,I9156,I9159);
and I_5708 (I99676,I99659,I9150);
DFFARX1 I_5709 (I99676,I2595,I99625,I99702,);
nor I_5710 (I99593,I99702,I99651);
not I_5711 (I99724,I99702);
DFFARX1 I_5712 (I9156,I2595,I99625,I99750,);
nand I_5713 (I99758,I99750,I9162);
not I_5714 (I99775,I99758);
DFFARX1 I_5715 (I99775,I2595,I99625,I99801,);
not I_5716 (I99617,I99801);
nor I_5717 (I99823,I99651,I99758);
nor I_5718 (I99599,I99702,I99823);
DFFARX1 I_5719 (I9153,I2595,I99625,I99863,);
DFFARX1 I_5720 (I99863,I2595,I99625,I99880,);
not I_5721 (I99888,I99880);
not I_5722 (I99905,I99863);
nand I_5723 (I99602,I99905,I99724);
nand I_5724 (I99936,I9153,I9168);
and I_5725 (I99953,I99936,I9150);
DFFARX1 I_5726 (I99953,I2595,I99625,I99979,);
nor I_5727 (I99987,I99979,I99651);
DFFARX1 I_5728 (I99987,I2595,I99625,I99590,);
DFFARX1 I_5729 (I99979,I2595,I99625,I99608,);
nor I_5730 (I100032,I9171,I9168);
not I_5731 (I100049,I100032);
nor I_5732 (I99611,I99888,I100049);
nand I_5733 (I99596,I99905,I100049);
nor I_5734 (I99605,I99651,I100032);
DFFARX1 I_5735 (I100032,I2595,I99625,I99614,);
not I_5736 (I100152,I2602);
DFFARX1 I_5737 (I162233,I2595,I100152,I100178,);
nand I_5738 (I100186,I162218,I162221);
and I_5739 (I100203,I100186,I162236);
DFFARX1 I_5740 (I100203,I2595,I100152,I100229,);
nor I_5741 (I100120,I100229,I100178);
not I_5742 (I100251,I100229);
DFFARX1 I_5743 (I162230,I2595,I100152,I100277,);
nand I_5744 (I100285,I100277,I162221);
not I_5745 (I100302,I100285);
DFFARX1 I_5746 (I100302,I2595,I100152,I100328,);
not I_5747 (I100144,I100328);
nor I_5748 (I100350,I100178,I100285);
nor I_5749 (I100126,I100229,I100350);
DFFARX1 I_5750 (I162227,I2595,I100152,I100390,);
DFFARX1 I_5751 (I100390,I2595,I100152,I100407,);
not I_5752 (I100415,I100407);
not I_5753 (I100432,I100390);
nand I_5754 (I100129,I100432,I100251);
nand I_5755 (I100463,I162242,I162218);
and I_5756 (I100480,I100463,I162239);
DFFARX1 I_5757 (I100480,I2595,I100152,I100506,);
nor I_5758 (I100514,I100506,I100178);
DFFARX1 I_5759 (I100514,I2595,I100152,I100117,);
DFFARX1 I_5760 (I100506,I2595,I100152,I100135,);
nor I_5761 (I100559,I162224,I162218);
not I_5762 (I100576,I100559);
nor I_5763 (I100138,I100415,I100576);
nand I_5764 (I100123,I100432,I100576);
nor I_5765 (I100132,I100178,I100559);
DFFARX1 I_5766 (I100559,I2595,I100152,I100141,);
not I_5767 (I100679,I2602);
DFFARX1 I_5768 (I245130,I2595,I100679,I100705,);
nand I_5769 (I100713,I245133,I245127);
and I_5770 (I100730,I100713,I245139);
DFFARX1 I_5771 (I100730,I2595,I100679,I100756,);
nor I_5772 (I100647,I100756,I100705);
not I_5773 (I100778,I100756);
DFFARX1 I_5774 (I245142,I2595,I100679,I100804,);
nand I_5775 (I100812,I100804,I245133);
not I_5776 (I100829,I100812);
DFFARX1 I_5777 (I100829,I2595,I100679,I100855,);
not I_5778 (I100671,I100855);
nor I_5779 (I100877,I100705,I100812);
nor I_5780 (I100653,I100756,I100877);
DFFARX1 I_5781 (I245145,I2595,I100679,I100917,);
DFFARX1 I_5782 (I100917,I2595,I100679,I100934,);
not I_5783 (I100942,I100934);
not I_5784 (I100959,I100917);
nand I_5785 (I100656,I100959,I100778);
nand I_5786 (I100990,I245127,I245136);
and I_5787 (I101007,I100990,I245130);
DFFARX1 I_5788 (I101007,I2595,I100679,I101033,);
nor I_5789 (I101041,I101033,I100705);
DFFARX1 I_5790 (I101041,I2595,I100679,I100644,);
DFFARX1 I_5791 (I101033,I2595,I100679,I100662,);
nor I_5792 (I101086,I245148,I245136);
not I_5793 (I101103,I101086);
nor I_5794 (I100665,I100942,I101103);
nand I_5795 (I100650,I100959,I101103);
nor I_5796 (I100659,I100705,I101086);
DFFARX1 I_5797 (I101086,I2595,I100679,I100668,);
not I_5798 (I101206,I2602);
DFFARX1 I_5799 (I22920,I2595,I101206,I101232,);
nand I_5800 (I101240,I22944,I22923);
and I_5801 (I101257,I101240,I22920);
DFFARX1 I_5802 (I101257,I2595,I101206,I101283,);
nor I_5803 (I101174,I101283,I101232);
not I_5804 (I101305,I101283);
DFFARX1 I_5805 (I22926,I2595,I101206,I101331,);
nand I_5806 (I101339,I101331,I22935);
not I_5807 (I101356,I101339);
DFFARX1 I_5808 (I101356,I2595,I101206,I101382,);
not I_5809 (I101198,I101382);
nor I_5810 (I101404,I101232,I101339);
nor I_5811 (I101180,I101283,I101404);
DFFARX1 I_5812 (I22929,I2595,I101206,I101444,);
DFFARX1 I_5813 (I101444,I2595,I101206,I101461,);
not I_5814 (I101469,I101461);
not I_5815 (I101486,I101444);
nand I_5816 (I101183,I101486,I101305);
nand I_5817 (I101517,I22941,I22923);
and I_5818 (I101534,I101517,I22932);
DFFARX1 I_5819 (I101534,I2595,I101206,I101560,);
nor I_5820 (I101568,I101560,I101232);
DFFARX1 I_5821 (I101568,I2595,I101206,I101171,);
DFFARX1 I_5822 (I101560,I2595,I101206,I101189,);
nor I_5823 (I101613,I22938,I22923);
not I_5824 (I101630,I101613);
nor I_5825 (I101192,I101469,I101630);
nand I_5826 (I101177,I101486,I101630);
nor I_5827 (I101186,I101232,I101613);
DFFARX1 I_5828 (I101613,I2595,I101206,I101195,);
not I_5829 (I101733,I2602);
DFFARX1 I_5830 (I133381,I2595,I101733,I101759,);
nand I_5831 (I101767,I133393,I133372);
and I_5832 (I101784,I101767,I133396);
DFFARX1 I_5833 (I101784,I2595,I101733,I101810,);
nor I_5834 (I101701,I101810,I101759);
not I_5835 (I101832,I101810);
DFFARX1 I_5836 (I133387,I2595,I101733,I101858,);
nand I_5837 (I101866,I101858,I133369);
not I_5838 (I101883,I101866);
DFFARX1 I_5839 (I101883,I2595,I101733,I101909,);
not I_5840 (I101725,I101909);
nor I_5841 (I101931,I101759,I101866);
nor I_5842 (I101707,I101810,I101931);
DFFARX1 I_5843 (I133384,I2595,I101733,I101971,);
DFFARX1 I_5844 (I101971,I2595,I101733,I101988,);
not I_5845 (I101996,I101988);
not I_5846 (I102013,I101971);
nand I_5847 (I101710,I102013,I101832);
nand I_5848 (I102044,I133369,I133375);
and I_5849 (I102061,I102044,I133378);
DFFARX1 I_5850 (I102061,I2595,I101733,I102087,);
nor I_5851 (I102095,I102087,I101759);
DFFARX1 I_5852 (I102095,I2595,I101733,I101698,);
DFFARX1 I_5853 (I102087,I2595,I101733,I101716,);
nor I_5854 (I102140,I133390,I133375);
not I_5855 (I102157,I102140);
nor I_5856 (I101719,I101996,I102157);
nand I_5857 (I101704,I102013,I102157);
nor I_5858 (I101713,I101759,I102140);
DFFARX1 I_5859 (I102140,I2595,I101733,I101722,);
not I_5860 (I102260,I2602);
DFFARX1 I_5861 (I180729,I2595,I102260,I102286,);
nand I_5862 (I102294,I180714,I180717);
and I_5863 (I102311,I102294,I180732);
DFFARX1 I_5864 (I102311,I2595,I102260,I102337,);
nor I_5865 (I102228,I102337,I102286);
not I_5866 (I102359,I102337);
DFFARX1 I_5867 (I180726,I2595,I102260,I102385,);
nand I_5868 (I102393,I102385,I180717);
not I_5869 (I102410,I102393);
DFFARX1 I_5870 (I102410,I2595,I102260,I102436,);
not I_5871 (I102252,I102436);
nor I_5872 (I102458,I102286,I102393);
nor I_5873 (I102234,I102337,I102458);
DFFARX1 I_5874 (I180723,I2595,I102260,I102498,);
DFFARX1 I_5875 (I102498,I2595,I102260,I102515,);
not I_5876 (I102523,I102515);
not I_5877 (I102540,I102498);
nand I_5878 (I102237,I102540,I102359);
nand I_5879 (I102571,I180738,I180714);
and I_5880 (I102588,I102571,I180735);
DFFARX1 I_5881 (I102588,I2595,I102260,I102614,);
nor I_5882 (I102622,I102614,I102286);
DFFARX1 I_5883 (I102622,I2595,I102260,I102225,);
DFFARX1 I_5884 (I102614,I2595,I102260,I102243,);
nor I_5885 (I102667,I180720,I180714);
not I_5886 (I102684,I102667);
nor I_5887 (I102246,I102523,I102684);
nand I_5888 (I102231,I102540,I102684);
nor I_5889 (I102240,I102286,I102667);
DFFARX1 I_5890 (I102667,I2595,I102260,I102249,);
not I_5891 (I102787,I2602);
DFFARX1 I_5892 (I386639,I2595,I102787,I102813,);
nand I_5893 (I102821,I386618,I386618);
and I_5894 (I102838,I102821,I386645);
DFFARX1 I_5895 (I102838,I2595,I102787,I102864,);
nor I_5896 (I102755,I102864,I102813);
not I_5897 (I102886,I102864);
DFFARX1 I_5898 (I386633,I2595,I102787,I102912,);
nand I_5899 (I102920,I102912,I386636);
not I_5900 (I102937,I102920);
DFFARX1 I_5901 (I102937,I2595,I102787,I102963,);
not I_5902 (I102779,I102963);
nor I_5903 (I102985,I102813,I102920);
nor I_5904 (I102761,I102864,I102985);
DFFARX1 I_5905 (I386627,I2595,I102787,I103025,);
DFFARX1 I_5906 (I103025,I2595,I102787,I103042,);
not I_5907 (I103050,I103042);
not I_5908 (I103067,I103025);
nand I_5909 (I102764,I103067,I102886);
nand I_5910 (I103098,I386624,I386621);
and I_5911 (I103115,I103098,I386642);
DFFARX1 I_5912 (I103115,I2595,I102787,I103141,);
nor I_5913 (I103149,I103141,I102813);
DFFARX1 I_5914 (I103149,I2595,I102787,I102752,);
DFFARX1 I_5915 (I103141,I2595,I102787,I102770,);
nor I_5916 (I103194,I386630,I386621);
not I_5917 (I103211,I103194);
nor I_5918 (I102773,I103050,I103211);
nand I_5919 (I102758,I103067,I103211);
nor I_5920 (I102767,I102813,I103194);
DFFARX1 I_5921 (I103194,I2595,I102787,I102776,);
not I_5922 (I103314,I2602);
DFFARX1 I_5923 (I50273,I2595,I103314,I103340,);
nand I_5924 (I103348,I50273,I50279);
and I_5925 (I103365,I103348,I50297);
DFFARX1 I_5926 (I103365,I2595,I103314,I103391,);
nor I_5927 (I103282,I103391,I103340);
not I_5928 (I103413,I103391);
DFFARX1 I_5929 (I50285,I2595,I103314,I103439,);
nand I_5930 (I103447,I103439,I50282);
not I_5931 (I103464,I103447);
DFFARX1 I_5932 (I103464,I2595,I103314,I103490,);
not I_5933 (I103306,I103490);
nor I_5934 (I103512,I103340,I103447);
nor I_5935 (I103288,I103391,I103512);
DFFARX1 I_5936 (I50291,I2595,I103314,I103552,);
DFFARX1 I_5937 (I103552,I2595,I103314,I103569,);
not I_5938 (I103577,I103569);
not I_5939 (I103594,I103552);
nand I_5940 (I103291,I103594,I103413);
nand I_5941 (I103625,I50276,I50276);
and I_5942 (I103642,I103625,I50288);
DFFARX1 I_5943 (I103642,I2595,I103314,I103668,);
nor I_5944 (I103676,I103668,I103340);
DFFARX1 I_5945 (I103676,I2595,I103314,I103279,);
DFFARX1 I_5946 (I103668,I2595,I103314,I103297,);
nor I_5947 (I103721,I50294,I50276);
not I_5948 (I103738,I103721);
nor I_5949 (I103300,I103577,I103738);
nand I_5950 (I103285,I103594,I103738);
nor I_5951 (I103294,I103340,I103721);
DFFARX1 I_5952 (I103721,I2595,I103314,I103303,);
not I_5953 (I103841,I2602);
DFFARX1 I_5954 (I202112,I2595,I103841,I103867,);
nand I_5955 (I103875,I202103,I202118);
and I_5956 (I103892,I103875,I202124);
DFFARX1 I_5957 (I103892,I2595,I103841,I103918,);
nor I_5958 (I103809,I103918,I103867);
not I_5959 (I103940,I103918);
DFFARX1 I_5960 (I202109,I2595,I103841,I103966,);
nand I_5961 (I103974,I103966,I202103);
not I_5962 (I103991,I103974);
DFFARX1 I_5963 (I103991,I2595,I103841,I104017,);
not I_5964 (I103833,I104017);
nor I_5965 (I104039,I103867,I103974);
nor I_5966 (I103815,I103918,I104039);
DFFARX1 I_5967 (I202106,I2595,I103841,I104079,);
DFFARX1 I_5968 (I104079,I2595,I103841,I104096,);
not I_5969 (I104104,I104096);
not I_5970 (I104121,I104079);
nand I_5971 (I103818,I104121,I103940);
nand I_5972 (I104152,I202100,I202115);
and I_5973 (I104169,I104152,I202100);
DFFARX1 I_5974 (I104169,I2595,I103841,I104195,);
nor I_5975 (I104203,I104195,I103867);
DFFARX1 I_5976 (I104203,I2595,I103841,I103806,);
DFFARX1 I_5977 (I104195,I2595,I103841,I103824,);
nor I_5978 (I104248,I202121,I202115);
not I_5979 (I104265,I104248);
nor I_5980 (I103827,I104104,I104265);
nand I_5981 (I103812,I104121,I104265);
nor I_5982 (I103821,I103867,I104248);
DFFARX1 I_5983 (I104248,I2595,I103841,I103830,);
not I_5984 (I104368,I2602);
DFFARX1 I_5985 (I343728,I2595,I104368,I104394,);
nand I_5986 (I104402,I343710,I343734);
and I_5987 (I104419,I104402,I343725);
DFFARX1 I_5988 (I104419,I2595,I104368,I104445,);
nor I_5989 (I104336,I104445,I104394);
not I_5990 (I104467,I104445);
DFFARX1 I_5991 (I343731,I2595,I104368,I104493,);
nand I_5992 (I104501,I104493,I343719);
not I_5993 (I104518,I104501);
DFFARX1 I_5994 (I104518,I2595,I104368,I104544,);
not I_5995 (I104360,I104544);
nor I_5996 (I104566,I104394,I104501);
nor I_5997 (I104342,I104445,I104566);
DFFARX1 I_5998 (I343710,I2595,I104368,I104606,);
DFFARX1 I_5999 (I104606,I2595,I104368,I104623,);
not I_6000 (I104631,I104623);
not I_6001 (I104648,I104606);
nand I_6002 (I104345,I104648,I104467);
nand I_6003 (I104679,I343716,I343713);
and I_6004 (I104696,I104679,I343722);
DFFARX1 I_6005 (I104696,I2595,I104368,I104722,);
nor I_6006 (I104730,I104722,I104394);
DFFARX1 I_6007 (I104730,I2595,I104368,I104333,);
DFFARX1 I_6008 (I104722,I2595,I104368,I104351,);
nor I_6009 (I104775,I343713,I343713);
not I_6010 (I104792,I104775);
nor I_6011 (I104354,I104631,I104792);
nand I_6012 (I104339,I104648,I104792);
nor I_6013 (I104348,I104394,I104775);
DFFARX1 I_6014 (I104775,I2595,I104368,I104357,);
not I_6015 (I104895,I2602);
DFFARX1 I_6016 (I1604,I2595,I104895,I104921,);
nand I_6017 (I104929,I2052,I1964);
and I_6018 (I104946,I104929,I1884);
DFFARX1 I_6019 (I104946,I2595,I104895,I104972,);
nor I_6020 (I104863,I104972,I104921);
not I_6021 (I104994,I104972);
DFFARX1 I_6022 (I2556,I2595,I104895,I105020,);
nand I_6023 (I105028,I105020,I2148);
not I_6024 (I105045,I105028);
DFFARX1 I_6025 (I105045,I2595,I104895,I105071,);
not I_6026 (I104887,I105071);
nor I_6027 (I105093,I104921,I105028);
nor I_6028 (I104869,I104972,I105093);
DFFARX1 I_6029 (I2404,I2595,I104895,I105133,);
DFFARX1 I_6030 (I105133,I2595,I104895,I105150,);
not I_6031 (I105158,I105150);
not I_6032 (I105175,I105133);
nand I_6033 (I104872,I105175,I104994);
nand I_6034 (I105206,I1652,I1460);
and I_6035 (I105223,I105206,I2124);
DFFARX1 I_6036 (I105223,I2595,I104895,I105249,);
nor I_6037 (I105257,I105249,I104921);
DFFARX1 I_6038 (I105257,I2595,I104895,I104860,);
DFFARX1 I_6039 (I105249,I2595,I104895,I104878,);
nor I_6040 (I105302,I1932,I1460);
not I_6041 (I105319,I105302);
nor I_6042 (I104881,I105158,I105319);
nand I_6043 (I104866,I105175,I105319);
nor I_6044 (I104875,I104921,I105302);
DFFARX1 I_6045 (I105302,I2595,I104895,I104884,);
not I_6046 (I105422,I2602);
DFFARX1 I_6047 (I134469,I2595,I105422,I105448,);
nand I_6048 (I105456,I134481,I134460);
and I_6049 (I105473,I105456,I134484);
DFFARX1 I_6050 (I105473,I2595,I105422,I105499,);
nor I_6051 (I105390,I105499,I105448);
not I_6052 (I105521,I105499);
DFFARX1 I_6053 (I134475,I2595,I105422,I105547,);
nand I_6054 (I105555,I105547,I134457);
not I_6055 (I105572,I105555);
DFFARX1 I_6056 (I105572,I2595,I105422,I105598,);
not I_6057 (I105414,I105598);
nor I_6058 (I105620,I105448,I105555);
nor I_6059 (I105396,I105499,I105620);
DFFARX1 I_6060 (I134472,I2595,I105422,I105660,);
DFFARX1 I_6061 (I105660,I2595,I105422,I105677,);
not I_6062 (I105685,I105677);
not I_6063 (I105702,I105660);
nand I_6064 (I105399,I105702,I105521);
nand I_6065 (I105733,I134457,I134463);
and I_6066 (I105750,I105733,I134466);
DFFARX1 I_6067 (I105750,I2595,I105422,I105776,);
nor I_6068 (I105784,I105776,I105448);
DFFARX1 I_6069 (I105784,I2595,I105422,I105387,);
DFFARX1 I_6070 (I105776,I2595,I105422,I105405,);
nor I_6071 (I105829,I134478,I134463);
not I_6072 (I105846,I105829);
nor I_6073 (I105408,I105685,I105846);
nand I_6074 (I105393,I105702,I105846);
nor I_6075 (I105402,I105448,I105829);
DFFARX1 I_6076 (I105829,I2595,I105422,I105411,);
not I_6077 (I105949,I2602);
DFFARX1 I_6078 (I200956,I2595,I105949,I105975,);
nand I_6079 (I105983,I200947,I200962);
and I_6080 (I106000,I105983,I200968);
DFFARX1 I_6081 (I106000,I2595,I105949,I106026,);
nor I_6082 (I105917,I106026,I105975);
not I_6083 (I106048,I106026);
DFFARX1 I_6084 (I200953,I2595,I105949,I106074,);
nand I_6085 (I106082,I106074,I200947);
not I_6086 (I106099,I106082);
DFFARX1 I_6087 (I106099,I2595,I105949,I106125,);
not I_6088 (I105941,I106125);
nor I_6089 (I106147,I105975,I106082);
nor I_6090 (I105923,I106026,I106147);
DFFARX1 I_6091 (I200950,I2595,I105949,I106187,);
DFFARX1 I_6092 (I106187,I2595,I105949,I106204,);
not I_6093 (I106212,I106204);
not I_6094 (I106229,I106187);
nand I_6095 (I105926,I106229,I106048);
nand I_6096 (I106260,I200944,I200959);
and I_6097 (I106277,I106260,I200944);
DFFARX1 I_6098 (I106277,I2595,I105949,I106303,);
nor I_6099 (I106311,I106303,I105975);
DFFARX1 I_6100 (I106311,I2595,I105949,I105914,);
DFFARX1 I_6101 (I106303,I2595,I105949,I105932,);
nor I_6102 (I106356,I200965,I200959);
not I_6103 (I106373,I106356);
nor I_6104 (I105935,I106212,I106373);
nand I_6105 (I105920,I106229,I106373);
nor I_6106 (I105929,I105975,I106356);
DFFARX1 I_6107 (I106356,I2595,I105949,I105938,);
not I_6108 (I106476,I2602);
DFFARX1 I_6109 (I321780,I2595,I106476,I106502,);
nand I_6110 (I106510,I321795,I321780);
and I_6111 (I106527,I106510,I321798);
DFFARX1 I_6112 (I106527,I2595,I106476,I106553,);
nor I_6113 (I106444,I106553,I106502);
not I_6114 (I106575,I106553);
DFFARX1 I_6115 (I321804,I2595,I106476,I106601,);
nand I_6116 (I106609,I106601,I321786);
not I_6117 (I106626,I106609);
DFFARX1 I_6118 (I106626,I2595,I106476,I106652,);
not I_6119 (I106468,I106652);
nor I_6120 (I106674,I106502,I106609);
nor I_6121 (I106450,I106553,I106674);
DFFARX1 I_6122 (I321783,I2595,I106476,I106714,);
DFFARX1 I_6123 (I106714,I2595,I106476,I106731,);
not I_6124 (I106739,I106731);
not I_6125 (I106756,I106714);
nand I_6126 (I106453,I106756,I106575);
nand I_6127 (I106787,I321783,I321789);
and I_6128 (I106804,I106787,I321801);
DFFARX1 I_6129 (I106804,I2595,I106476,I106830,);
nor I_6130 (I106838,I106830,I106502);
DFFARX1 I_6131 (I106838,I2595,I106476,I106441,);
DFFARX1 I_6132 (I106830,I2595,I106476,I106459,);
nor I_6133 (I106883,I321792,I321789);
not I_6134 (I106900,I106883);
nor I_6135 (I106462,I106739,I106900);
nand I_6136 (I106447,I106756,I106900);
nor I_6137 (I106456,I106502,I106883);
DFFARX1 I_6138 (I106883,I2595,I106476,I106465,);
not I_6139 (I107003,I2602);
DFFARX1 I_6140 (I170325,I2595,I107003,I107029,);
nand I_6141 (I107037,I170310,I170313);
and I_6142 (I107054,I107037,I170328);
DFFARX1 I_6143 (I107054,I2595,I107003,I107080,);
nor I_6144 (I106971,I107080,I107029);
not I_6145 (I107102,I107080);
DFFARX1 I_6146 (I170322,I2595,I107003,I107128,);
nand I_6147 (I107136,I107128,I170313);
not I_6148 (I107153,I107136);
DFFARX1 I_6149 (I107153,I2595,I107003,I107179,);
not I_6150 (I106995,I107179);
nor I_6151 (I107201,I107029,I107136);
nor I_6152 (I106977,I107080,I107201);
DFFARX1 I_6153 (I170319,I2595,I107003,I107241,);
DFFARX1 I_6154 (I107241,I2595,I107003,I107258,);
not I_6155 (I107266,I107258);
not I_6156 (I107283,I107241);
nand I_6157 (I106980,I107283,I107102);
nand I_6158 (I107314,I170334,I170310);
and I_6159 (I107331,I107314,I170331);
DFFARX1 I_6160 (I107331,I2595,I107003,I107357,);
nor I_6161 (I107365,I107357,I107029);
DFFARX1 I_6162 (I107365,I2595,I107003,I106968,);
DFFARX1 I_6163 (I107357,I2595,I107003,I106986,);
nor I_6164 (I107410,I170316,I170310);
not I_6165 (I107427,I107410);
nor I_6166 (I106989,I107266,I107427);
nand I_6167 (I106974,I107283,I107427);
nor I_6168 (I106983,I107029,I107410);
DFFARX1 I_6169 (I107410,I2595,I107003,I106992,);
not I_6170 (I107530,I2602);
DFFARX1 I_6171 (I321202,I2595,I107530,I107556,);
nand I_6172 (I107564,I321217,I321202);
and I_6173 (I107581,I107564,I321220);
DFFARX1 I_6174 (I107581,I2595,I107530,I107607,);
nor I_6175 (I107498,I107607,I107556);
not I_6176 (I107629,I107607);
DFFARX1 I_6177 (I321226,I2595,I107530,I107655,);
nand I_6178 (I107663,I107655,I321208);
not I_6179 (I107680,I107663);
DFFARX1 I_6180 (I107680,I2595,I107530,I107706,);
not I_6181 (I107522,I107706);
nor I_6182 (I107728,I107556,I107663);
nor I_6183 (I107504,I107607,I107728);
DFFARX1 I_6184 (I321205,I2595,I107530,I107768,);
DFFARX1 I_6185 (I107768,I2595,I107530,I107785,);
not I_6186 (I107793,I107785);
not I_6187 (I107810,I107768);
nand I_6188 (I107507,I107810,I107629);
nand I_6189 (I107841,I321205,I321211);
and I_6190 (I107858,I107841,I321223);
DFFARX1 I_6191 (I107858,I2595,I107530,I107884,);
nor I_6192 (I107892,I107884,I107556);
DFFARX1 I_6193 (I107892,I2595,I107530,I107495,);
DFFARX1 I_6194 (I107884,I2595,I107530,I107513,);
nor I_6195 (I107937,I321214,I321211);
not I_6196 (I107954,I107937);
nor I_6197 (I107516,I107793,I107954);
nand I_6198 (I107501,I107810,I107954);
nor I_6199 (I107510,I107556,I107937);
DFFARX1 I_6200 (I107937,I2595,I107530,I107519,);
not I_6201 (I108057,I2602);
DFFARX1 I_6202 (I44530,I2595,I108057,I108083,);
nand I_6203 (I108091,I44542,I44551);
and I_6204 (I108108,I108091,I44530);
DFFARX1 I_6205 (I108108,I2595,I108057,I108134,);
nor I_6206 (I108025,I108134,I108083);
not I_6207 (I108156,I108134);
DFFARX1 I_6208 (I44545,I2595,I108057,I108182,);
nand I_6209 (I108190,I108182,I44533);
not I_6210 (I108207,I108190);
DFFARX1 I_6211 (I108207,I2595,I108057,I108233,);
not I_6212 (I108049,I108233);
nor I_6213 (I108255,I108083,I108190);
nor I_6214 (I108031,I108134,I108255);
DFFARX1 I_6215 (I44536,I2595,I108057,I108295,);
DFFARX1 I_6216 (I108295,I2595,I108057,I108312,);
not I_6217 (I108320,I108312);
not I_6218 (I108337,I108295);
nand I_6219 (I108034,I108337,I108156);
nand I_6220 (I108368,I44527,I44527);
and I_6221 (I108385,I108368,I44539);
DFFARX1 I_6222 (I108385,I2595,I108057,I108411,);
nor I_6223 (I108419,I108411,I108083);
DFFARX1 I_6224 (I108419,I2595,I108057,I108022,);
DFFARX1 I_6225 (I108411,I2595,I108057,I108040,);
nor I_6226 (I108464,I44548,I44527);
not I_6227 (I108481,I108464);
nor I_6228 (I108043,I108320,I108481);
nand I_6229 (I108028,I108337,I108481);
nor I_6230 (I108037,I108083,I108464);
DFFARX1 I_6231 (I108464,I2595,I108057,I108046,);
not I_6232 (I108584,I2602);
DFFARX1 I_6233 (I42422,I2595,I108584,I108610,);
nand I_6234 (I108618,I42434,I42443);
and I_6235 (I108635,I108618,I42422);
DFFARX1 I_6236 (I108635,I2595,I108584,I108661,);
nor I_6237 (I108552,I108661,I108610);
not I_6238 (I108683,I108661);
DFFARX1 I_6239 (I42437,I2595,I108584,I108709,);
nand I_6240 (I108717,I108709,I42425);
not I_6241 (I108734,I108717);
DFFARX1 I_6242 (I108734,I2595,I108584,I108760,);
not I_6243 (I108576,I108760);
nor I_6244 (I108782,I108610,I108717);
nor I_6245 (I108558,I108661,I108782);
DFFARX1 I_6246 (I42428,I2595,I108584,I108822,);
DFFARX1 I_6247 (I108822,I2595,I108584,I108839,);
not I_6248 (I108847,I108839);
not I_6249 (I108864,I108822);
nand I_6250 (I108561,I108864,I108683);
nand I_6251 (I108895,I42419,I42419);
and I_6252 (I108912,I108895,I42431);
DFFARX1 I_6253 (I108912,I2595,I108584,I108938,);
nor I_6254 (I108946,I108938,I108610);
DFFARX1 I_6255 (I108946,I2595,I108584,I108549,);
DFFARX1 I_6256 (I108938,I2595,I108584,I108567,);
nor I_6257 (I108991,I42440,I42419);
not I_6258 (I109008,I108991);
nor I_6259 (I108570,I108847,I109008);
nand I_6260 (I108555,I108864,I109008);
nor I_6261 (I108564,I108610,I108991);
DFFARX1 I_6262 (I108991,I2595,I108584,I108573,);
not I_6263 (I109111,I2602);
DFFARX1 I_6264 (I69313,I2595,I109111,I109137,);
nand I_6265 (I109145,I69313,I69319);
and I_6266 (I109162,I109145,I69337);
DFFARX1 I_6267 (I109162,I2595,I109111,I109188,);
nor I_6268 (I109079,I109188,I109137);
not I_6269 (I109210,I109188);
DFFARX1 I_6270 (I69325,I2595,I109111,I109236,);
nand I_6271 (I109244,I109236,I69322);
not I_6272 (I109261,I109244);
DFFARX1 I_6273 (I109261,I2595,I109111,I109287,);
not I_6274 (I109103,I109287);
nor I_6275 (I109309,I109137,I109244);
nor I_6276 (I109085,I109188,I109309);
DFFARX1 I_6277 (I69331,I2595,I109111,I109349,);
DFFARX1 I_6278 (I109349,I2595,I109111,I109366,);
not I_6279 (I109374,I109366);
not I_6280 (I109391,I109349);
nand I_6281 (I109088,I109391,I109210);
nand I_6282 (I109422,I69316,I69316);
and I_6283 (I109439,I109422,I69328);
DFFARX1 I_6284 (I109439,I2595,I109111,I109465,);
nor I_6285 (I109473,I109465,I109137);
DFFARX1 I_6286 (I109473,I2595,I109111,I109076,);
DFFARX1 I_6287 (I109465,I2595,I109111,I109094,);
nor I_6288 (I109518,I69334,I69316);
not I_6289 (I109535,I109518);
nor I_6290 (I109097,I109374,I109535);
nand I_6291 (I109082,I109391,I109535);
nor I_6292 (I109091,I109137,I109518);
DFFARX1 I_6293 (I109518,I2595,I109111,I109100,);
not I_6294 (I109638,I2602);
DFFARX1 I_6295 (I40314,I2595,I109638,I109664,);
nand I_6296 (I109672,I40326,I40335);
and I_6297 (I109689,I109672,I40314);
DFFARX1 I_6298 (I109689,I2595,I109638,I109715,);
nor I_6299 (I109606,I109715,I109664);
not I_6300 (I109737,I109715);
DFFARX1 I_6301 (I40329,I2595,I109638,I109763,);
nand I_6302 (I109771,I109763,I40317);
not I_6303 (I109788,I109771);
DFFARX1 I_6304 (I109788,I2595,I109638,I109814,);
not I_6305 (I109630,I109814);
nor I_6306 (I109836,I109664,I109771);
nor I_6307 (I109612,I109715,I109836);
DFFARX1 I_6308 (I40320,I2595,I109638,I109876,);
DFFARX1 I_6309 (I109876,I2595,I109638,I109893,);
not I_6310 (I109901,I109893);
not I_6311 (I109918,I109876);
nand I_6312 (I109615,I109918,I109737);
nand I_6313 (I109949,I40311,I40311);
and I_6314 (I109966,I109949,I40323);
DFFARX1 I_6315 (I109966,I2595,I109638,I109992,);
nor I_6316 (I110000,I109992,I109664);
DFFARX1 I_6317 (I110000,I2595,I109638,I109603,);
DFFARX1 I_6318 (I109992,I2595,I109638,I109621,);
nor I_6319 (I110045,I40332,I40311);
not I_6320 (I110062,I110045);
nor I_6321 (I109624,I109901,I110062);
nand I_6322 (I109609,I109918,I110062);
nor I_6323 (I109618,I109664,I110045);
DFFARX1 I_6324 (I110045,I2595,I109638,I109627,);
not I_6325 (I110165,I2602);
DFFARX1 I_6326 (I21866,I2595,I110165,I110191,);
nand I_6327 (I110199,I21890,I21869);
and I_6328 (I110216,I110199,I21866);
DFFARX1 I_6329 (I110216,I2595,I110165,I110242,);
nor I_6330 (I110133,I110242,I110191);
not I_6331 (I110264,I110242);
DFFARX1 I_6332 (I21872,I2595,I110165,I110290,);
nand I_6333 (I110298,I110290,I21881);
not I_6334 (I110315,I110298);
DFFARX1 I_6335 (I110315,I2595,I110165,I110341,);
not I_6336 (I110157,I110341);
nor I_6337 (I110363,I110191,I110298);
nor I_6338 (I110139,I110242,I110363);
DFFARX1 I_6339 (I21875,I2595,I110165,I110403,);
DFFARX1 I_6340 (I110403,I2595,I110165,I110420,);
not I_6341 (I110428,I110420);
not I_6342 (I110445,I110403);
nand I_6343 (I110142,I110445,I110264);
nand I_6344 (I110476,I21887,I21869);
and I_6345 (I110493,I110476,I21878);
DFFARX1 I_6346 (I110493,I2595,I110165,I110519,);
nor I_6347 (I110527,I110519,I110191);
DFFARX1 I_6348 (I110527,I2595,I110165,I110130,);
DFFARX1 I_6349 (I110519,I2595,I110165,I110148,);
nor I_6350 (I110572,I21884,I21869);
not I_6351 (I110589,I110572);
nor I_6352 (I110151,I110428,I110589);
nand I_6353 (I110136,I110445,I110589);
nor I_6354 (I110145,I110191,I110572);
DFFARX1 I_6355 (I110572,I2595,I110165,I110154,);
not I_6356 (I110692,I2602);
DFFARX1 I_6357 (I283516,I2595,I110692,I110718,);
nand I_6358 (I110726,I283513,I283531);
and I_6359 (I110743,I110726,I283522);
DFFARX1 I_6360 (I110743,I2595,I110692,I110769,);
nor I_6361 (I110660,I110769,I110718);
not I_6362 (I110791,I110769);
DFFARX1 I_6363 (I283537,I2595,I110692,I110817,);
nand I_6364 (I110825,I110817,I283519);
not I_6365 (I110842,I110825);
DFFARX1 I_6366 (I110842,I2595,I110692,I110868,);
not I_6367 (I110684,I110868);
nor I_6368 (I110890,I110718,I110825);
nor I_6369 (I110666,I110769,I110890);
DFFARX1 I_6370 (I283525,I2595,I110692,I110930,);
DFFARX1 I_6371 (I110930,I2595,I110692,I110947,);
not I_6372 (I110955,I110947);
not I_6373 (I110972,I110930);
nand I_6374 (I110669,I110972,I110791);
nand I_6375 (I111003,I283513,I283540);
and I_6376 (I111020,I111003,I283528);
DFFARX1 I_6377 (I111020,I2595,I110692,I111046,);
nor I_6378 (I111054,I111046,I110718);
DFFARX1 I_6379 (I111054,I2595,I110692,I110657,);
DFFARX1 I_6380 (I111046,I2595,I110692,I110675,);
nor I_6381 (I111099,I283534,I283540);
not I_6382 (I111116,I111099);
nor I_6383 (I110678,I110955,I111116);
nand I_6384 (I110663,I110972,I111116);
nor I_6385 (I110672,I110718,I111099);
DFFARX1 I_6386 (I111099,I2595,I110692,I110681,);
not I_6387 (I111219,I2602);
DFFARX1 I_6388 (I212516,I2595,I111219,I111245,);
nand I_6389 (I111253,I212507,I212522);
and I_6390 (I111270,I111253,I212528);
DFFARX1 I_6391 (I111270,I2595,I111219,I111296,);
nor I_6392 (I111187,I111296,I111245);
not I_6393 (I111318,I111296);
DFFARX1 I_6394 (I212513,I2595,I111219,I111344,);
nand I_6395 (I111352,I111344,I212507);
not I_6396 (I111369,I111352);
DFFARX1 I_6397 (I111369,I2595,I111219,I111395,);
not I_6398 (I111211,I111395);
nor I_6399 (I111417,I111245,I111352);
nor I_6400 (I111193,I111296,I111417);
DFFARX1 I_6401 (I212510,I2595,I111219,I111457,);
DFFARX1 I_6402 (I111457,I2595,I111219,I111474,);
not I_6403 (I111482,I111474);
not I_6404 (I111499,I111457);
nand I_6405 (I111196,I111499,I111318);
nand I_6406 (I111530,I212504,I212519);
and I_6407 (I111547,I111530,I212504);
DFFARX1 I_6408 (I111547,I2595,I111219,I111573,);
nor I_6409 (I111581,I111573,I111245);
DFFARX1 I_6410 (I111581,I2595,I111219,I111184,);
DFFARX1 I_6411 (I111573,I2595,I111219,I111202,);
nor I_6412 (I111626,I212525,I212519);
not I_6413 (I111643,I111626);
nor I_6414 (I111205,I111482,I111643);
nand I_6415 (I111190,I111499,I111643);
nor I_6416 (I111199,I111245,I111626);
DFFARX1 I_6417 (I111626,I2595,I111219,I111208,);
not I_6418 (I111746,I2602);
DFFARX1 I_6419 (I333340,I2595,I111746,I111772,);
nand I_6420 (I111780,I333355,I333340);
and I_6421 (I111797,I111780,I333358);
DFFARX1 I_6422 (I111797,I2595,I111746,I111823,);
nor I_6423 (I111714,I111823,I111772);
not I_6424 (I111845,I111823);
DFFARX1 I_6425 (I333364,I2595,I111746,I111871,);
nand I_6426 (I111879,I111871,I333346);
not I_6427 (I111896,I111879);
DFFARX1 I_6428 (I111896,I2595,I111746,I111922,);
not I_6429 (I111738,I111922);
nor I_6430 (I111944,I111772,I111879);
nor I_6431 (I111720,I111823,I111944);
DFFARX1 I_6432 (I333343,I2595,I111746,I111984,);
DFFARX1 I_6433 (I111984,I2595,I111746,I112001,);
not I_6434 (I112009,I112001);
not I_6435 (I112026,I111984);
nand I_6436 (I111723,I112026,I111845);
nand I_6437 (I112057,I333343,I333349);
and I_6438 (I112074,I112057,I333361);
DFFARX1 I_6439 (I112074,I2595,I111746,I112100,);
nor I_6440 (I112108,I112100,I111772);
DFFARX1 I_6441 (I112108,I2595,I111746,I111711,);
DFFARX1 I_6442 (I112100,I2595,I111746,I111729,);
nor I_6443 (I112153,I333352,I333349);
not I_6444 (I112170,I112153);
nor I_6445 (I111732,I112009,I112170);
nand I_6446 (I111717,I112026,I112170);
nor I_6447 (I111726,I111772,I112153);
DFFARX1 I_6448 (I112153,I2595,I111746,I111735,);
not I_6449 (I112273,I2602);
DFFARX1 I_6450 (I145748,I2595,I112273,I112299,);
nand I_6451 (I112307,I145748,I145760);
and I_6452 (I112324,I112307,I145745);
DFFARX1 I_6453 (I112324,I2595,I112273,I112350,);
nor I_6454 (I112241,I112350,I112299);
not I_6455 (I112372,I112350);
DFFARX1 I_6456 (I145769,I2595,I112273,I112398,);
nand I_6457 (I112406,I112398,I145766);
not I_6458 (I112423,I112406);
DFFARX1 I_6459 (I112423,I2595,I112273,I112449,);
not I_6460 (I112265,I112449);
nor I_6461 (I112471,I112299,I112406);
nor I_6462 (I112247,I112350,I112471);
DFFARX1 I_6463 (I145757,I2595,I112273,I112511,);
DFFARX1 I_6464 (I112511,I2595,I112273,I112528,);
not I_6465 (I112536,I112528);
not I_6466 (I112553,I112511);
nand I_6467 (I112250,I112553,I112372);
nand I_6468 (I112584,I145745,I145754);
and I_6469 (I112601,I112584,I145763);
DFFARX1 I_6470 (I112601,I2595,I112273,I112627,);
nor I_6471 (I112635,I112627,I112299);
DFFARX1 I_6472 (I112635,I2595,I112273,I112238,);
DFFARX1 I_6473 (I112627,I2595,I112273,I112256,);
nor I_6474 (I112680,I145751,I145754);
not I_6475 (I112697,I112680);
nor I_6476 (I112259,I112536,I112697);
nand I_6477 (I112244,I112553,I112697);
nor I_6478 (I112253,I112299,I112680);
DFFARX1 I_6479 (I112680,I2595,I112273,I112262,);
not I_6480 (I112800,I2602);
DFFARX1 I_6481 (I188240,I2595,I112800,I112826,);
nand I_6482 (I112834,I188231,I188246);
and I_6483 (I112851,I112834,I188252);
DFFARX1 I_6484 (I112851,I2595,I112800,I112877,);
nor I_6485 (I112768,I112877,I112826);
not I_6486 (I112899,I112877);
DFFARX1 I_6487 (I188237,I2595,I112800,I112925,);
nand I_6488 (I112933,I112925,I188231);
not I_6489 (I112950,I112933);
DFFARX1 I_6490 (I112950,I2595,I112800,I112976,);
not I_6491 (I112792,I112976);
nor I_6492 (I112998,I112826,I112933);
nor I_6493 (I112774,I112877,I112998);
DFFARX1 I_6494 (I188234,I2595,I112800,I113038,);
DFFARX1 I_6495 (I113038,I2595,I112800,I113055,);
not I_6496 (I113063,I113055);
not I_6497 (I113080,I113038);
nand I_6498 (I112777,I113080,I112899);
nand I_6499 (I113111,I188228,I188243);
and I_6500 (I113128,I113111,I188228);
DFFARX1 I_6501 (I113128,I2595,I112800,I113154,);
nor I_6502 (I113162,I113154,I112826);
DFFARX1 I_6503 (I113162,I2595,I112800,I112765,);
DFFARX1 I_6504 (I113154,I2595,I112800,I112783,);
nor I_6505 (I113207,I188249,I188243);
not I_6506 (I113224,I113207);
nor I_6507 (I112786,I113063,I113224);
nand I_6508 (I112771,I113080,I113224);
nor I_6509 (I112780,I112826,I113207);
DFFARX1 I_6510 (I113207,I2595,I112800,I112789,);
not I_6511 (I113327,I2602);
DFFARX1 I_6512 (I272534,I2595,I113327,I113353,);
nand I_6513 (I113361,I272531,I272549);
and I_6514 (I113378,I113361,I272540);
DFFARX1 I_6515 (I113378,I2595,I113327,I113404,);
nor I_6516 (I113295,I113404,I113353);
not I_6517 (I113426,I113404);
DFFARX1 I_6518 (I272555,I2595,I113327,I113452,);
nand I_6519 (I113460,I113452,I272537);
not I_6520 (I113477,I113460);
DFFARX1 I_6521 (I113477,I2595,I113327,I113503,);
not I_6522 (I113319,I113503);
nor I_6523 (I113525,I113353,I113460);
nor I_6524 (I113301,I113404,I113525);
DFFARX1 I_6525 (I272543,I2595,I113327,I113565,);
DFFARX1 I_6526 (I113565,I2595,I113327,I113582,);
not I_6527 (I113590,I113582);
not I_6528 (I113607,I113565);
nand I_6529 (I113304,I113607,I113426);
nand I_6530 (I113638,I272531,I272558);
and I_6531 (I113655,I113638,I272546);
DFFARX1 I_6532 (I113655,I2595,I113327,I113681,);
nor I_6533 (I113689,I113681,I113353);
DFFARX1 I_6534 (I113689,I2595,I113327,I113292,);
DFFARX1 I_6535 (I113681,I2595,I113327,I113310,);
nor I_6536 (I113734,I272552,I272558);
not I_6537 (I113751,I113734);
nor I_6538 (I113313,I113590,I113751);
nand I_6539 (I113298,I113607,I113751);
nor I_6540 (I113307,I113353,I113734);
DFFARX1 I_6541 (I113734,I2595,I113327,I113316,);
not I_6542 (I113854,I2602);
DFFARX1 I_6543 (I195176,I2595,I113854,I113880,);
nand I_6544 (I113888,I195167,I195182);
and I_6545 (I113905,I113888,I195188);
DFFARX1 I_6546 (I113905,I2595,I113854,I113931,);
nor I_6547 (I113822,I113931,I113880);
not I_6548 (I113953,I113931);
DFFARX1 I_6549 (I195173,I2595,I113854,I113979,);
nand I_6550 (I113987,I113979,I195167);
not I_6551 (I114004,I113987);
DFFARX1 I_6552 (I114004,I2595,I113854,I114030,);
not I_6553 (I113846,I114030);
nor I_6554 (I114052,I113880,I113987);
nor I_6555 (I113828,I113931,I114052);
DFFARX1 I_6556 (I195170,I2595,I113854,I114092,);
DFFARX1 I_6557 (I114092,I2595,I113854,I114109,);
not I_6558 (I114117,I114109);
not I_6559 (I114134,I114092);
nand I_6560 (I113831,I114134,I113953);
nand I_6561 (I114165,I195164,I195179);
and I_6562 (I114182,I114165,I195164);
DFFARX1 I_6563 (I114182,I2595,I113854,I114208,);
nor I_6564 (I114216,I114208,I113880);
DFFARX1 I_6565 (I114216,I2595,I113854,I113819,);
DFFARX1 I_6566 (I114208,I2595,I113854,I113837,);
nor I_6567 (I114261,I195185,I195179);
not I_6568 (I114278,I114261);
nor I_6569 (I113840,I114117,I114278);
nand I_6570 (I113825,I114134,I114278);
nor I_6571 (I113834,I113880,I114261);
DFFARX1 I_6572 (I114261,I2595,I113854,I113843,);
not I_6573 (I114381,I2602);
DFFARX1 I_6574 (I119781,I2595,I114381,I114407,);
nand I_6575 (I114415,I119793,I119772);
and I_6576 (I114432,I114415,I119796);
DFFARX1 I_6577 (I114432,I2595,I114381,I114458,);
nor I_6578 (I114349,I114458,I114407);
not I_6579 (I114480,I114458);
DFFARX1 I_6580 (I119787,I2595,I114381,I114506,);
nand I_6581 (I114514,I114506,I119769);
not I_6582 (I114531,I114514);
DFFARX1 I_6583 (I114531,I2595,I114381,I114557,);
not I_6584 (I114373,I114557);
nor I_6585 (I114579,I114407,I114514);
nor I_6586 (I114355,I114458,I114579);
DFFARX1 I_6587 (I119784,I2595,I114381,I114619,);
DFFARX1 I_6588 (I114619,I2595,I114381,I114636,);
not I_6589 (I114644,I114636);
not I_6590 (I114661,I114619);
nand I_6591 (I114358,I114661,I114480);
nand I_6592 (I114692,I119769,I119775);
and I_6593 (I114709,I114692,I119778);
DFFARX1 I_6594 (I114709,I2595,I114381,I114735,);
nor I_6595 (I114743,I114735,I114407);
DFFARX1 I_6596 (I114743,I2595,I114381,I114346,);
DFFARX1 I_6597 (I114735,I2595,I114381,I114364,);
nor I_6598 (I114788,I119790,I119775);
not I_6599 (I114805,I114788);
nor I_6600 (I114367,I114644,I114805);
nand I_6601 (I114352,I114661,I114805);
nor I_6602 (I114361,I114407,I114788);
DFFARX1 I_6603 (I114788,I2595,I114381,I114370,);
not I_6604 (I114908,I2602);
DFFARX1 I_6605 (I282227,I2595,I114908,I114934,);
DFFARX1 I_6606 (I114934,I2595,I114908,I114951,);
not I_6607 (I114900,I114951);
not I_6608 (I114973,I114934);
nand I_6609 (I114990,I282242,I282230);
and I_6610 (I115007,I114990,I282221);
DFFARX1 I_6611 (I115007,I2595,I114908,I115033,);
not I_6612 (I115041,I115033);
DFFARX1 I_6613 (I282233,I2595,I114908,I115067,);
and I_6614 (I115075,I115067,I282224);
nand I_6615 (I115092,I115067,I282224);
nand I_6616 (I114879,I115041,I115092);
DFFARX1 I_6617 (I282239,I2595,I114908,I115132,);
nor I_6618 (I115140,I115132,I115075);
DFFARX1 I_6619 (I115140,I2595,I114908,I114873,);
nor I_6620 (I114888,I115132,I115033);
nand I_6621 (I115185,I282248,I282236);
and I_6622 (I115202,I115185,I282245);
DFFARX1 I_6623 (I115202,I2595,I114908,I115228,);
nor I_6624 (I114876,I115228,I115132);
not I_6625 (I115250,I115228);
nor I_6626 (I115267,I115250,I115041);
nor I_6627 (I115284,I114973,I115267);
DFFARX1 I_6628 (I115284,I2595,I114908,I114891,);
nor I_6629 (I115315,I115250,I115132);
nor I_6630 (I115332,I282221,I282236);
nor I_6631 (I114882,I115332,I115315);
not I_6632 (I115363,I115332);
nand I_6633 (I114885,I115092,I115363);
DFFARX1 I_6634 (I115332,I2595,I114908,I114897,);
DFFARX1 I_6635 (I115332,I2595,I114908,I114894,);
not I_6636 (I115452,I2602);
DFFARX1 I_6637 (I155863,I2595,I115452,I115478,);
DFFARX1 I_6638 (I115478,I2595,I115452,I115495,);
not I_6639 (I115444,I115495);
not I_6640 (I115517,I115478);
nand I_6641 (I115534,I155860,I155881);
and I_6642 (I115551,I115534,I155884);
DFFARX1 I_6643 (I115551,I2595,I115452,I115577,);
not I_6644 (I115585,I115577);
DFFARX1 I_6645 (I155869,I2595,I115452,I115611,);
and I_6646 (I115619,I115611,I155872);
nand I_6647 (I115636,I115611,I155872);
nand I_6648 (I115423,I115585,I115636);
DFFARX1 I_6649 (I155875,I2595,I115452,I115676,);
nor I_6650 (I115684,I115676,I115619);
DFFARX1 I_6651 (I115684,I2595,I115452,I115417,);
nor I_6652 (I115432,I115676,I115577);
nand I_6653 (I115729,I155860,I155866);
and I_6654 (I115746,I115729,I155878);
DFFARX1 I_6655 (I115746,I2595,I115452,I115772,);
nor I_6656 (I115420,I115772,I115676);
not I_6657 (I115794,I115772);
nor I_6658 (I115811,I115794,I115585);
nor I_6659 (I115828,I115517,I115811);
DFFARX1 I_6660 (I115828,I2595,I115452,I115435,);
nor I_6661 (I115859,I115794,I115676);
nor I_6662 (I115876,I155863,I155866);
nor I_6663 (I115426,I115876,I115859);
not I_6664 (I115907,I115876);
nand I_6665 (I115429,I115636,I115907);
DFFARX1 I_6666 (I115876,I2595,I115452,I115441,);
DFFARX1 I_6667 (I115876,I2595,I115452,I115438,);
not I_6668 (I115996,I2602);
DFFARX1 I_6669 (I62777,I2595,I115996,I116022,);
DFFARX1 I_6670 (I116022,I2595,I115996,I116039,);
not I_6671 (I115988,I116039);
not I_6672 (I116061,I116022);
nand I_6673 (I116078,I62789,I62768);
and I_6674 (I116095,I116078,I62771);
DFFARX1 I_6675 (I116095,I2595,I115996,I116121,);
not I_6676 (I116129,I116121);
DFFARX1 I_6677 (I62780,I2595,I115996,I116155,);
and I_6678 (I116163,I116155,I62792);
nand I_6679 (I116180,I116155,I62792);
nand I_6680 (I115967,I116129,I116180);
DFFARX1 I_6681 (I62786,I2595,I115996,I116220,);
nor I_6682 (I116228,I116220,I116163);
DFFARX1 I_6683 (I116228,I2595,I115996,I115961,);
nor I_6684 (I115976,I116220,I116121);
nand I_6685 (I116273,I62774,I62771);
and I_6686 (I116290,I116273,I62783);
DFFARX1 I_6687 (I116290,I2595,I115996,I116316,);
nor I_6688 (I115964,I116316,I116220);
not I_6689 (I116338,I116316);
nor I_6690 (I116355,I116338,I116129);
nor I_6691 (I116372,I116061,I116355);
DFFARX1 I_6692 (I116372,I2595,I115996,I115979,);
nor I_6693 (I116403,I116338,I116220);
nor I_6694 (I116420,I62768,I62771);
nor I_6695 (I115970,I116420,I116403);
not I_6696 (I116451,I116420);
nand I_6697 (I115973,I116180,I116451);
DFFARX1 I_6698 (I116420,I2595,I115996,I115985,);
DFFARX1 I_6699 (I116420,I2595,I115996,I115982,);
not I_6700 (I116540,I2602);
DFFARX1 I_6701 (I377125,I2595,I116540,I116566,);
DFFARX1 I_6702 (I116566,I2595,I116540,I116583,);
not I_6703 (I116532,I116583);
not I_6704 (I116605,I116566);
nand I_6705 (I116622,I377101,I377122);
and I_6706 (I116639,I116622,I377119);
DFFARX1 I_6707 (I116639,I2595,I116540,I116665,);
not I_6708 (I116673,I116665);
DFFARX1 I_6709 (I377098,I2595,I116540,I116699,);
and I_6710 (I116707,I116699,I377110);
nand I_6711 (I116724,I116699,I377110);
nand I_6712 (I116511,I116673,I116724);
DFFARX1 I_6713 (I377113,I2595,I116540,I116764,);
nor I_6714 (I116772,I116764,I116707);
DFFARX1 I_6715 (I116772,I2595,I116540,I116505,);
nor I_6716 (I116520,I116764,I116665);
nand I_6717 (I116817,I377116,I377104);
and I_6718 (I116834,I116817,I377107);
DFFARX1 I_6719 (I116834,I2595,I116540,I116860,);
nor I_6720 (I116508,I116860,I116764);
not I_6721 (I116882,I116860);
nor I_6722 (I116899,I116882,I116673);
nor I_6723 (I116916,I116605,I116899);
DFFARX1 I_6724 (I116916,I2595,I116540,I116523,);
nor I_6725 (I116947,I116882,I116764);
nor I_6726 (I116964,I377098,I377104);
nor I_6727 (I116514,I116964,I116947);
not I_6728 (I116995,I116964);
nand I_6729 (I116517,I116724,I116995);
DFFARX1 I_6730 (I116964,I2595,I116540,I116529,);
DFFARX1 I_6731 (I116964,I2595,I116540,I116526,);
not I_6732 (I117084,I2602);
DFFARX1 I_6733 (I325251,I2595,I117084,I117110,);
DFFARX1 I_6734 (I117110,I2595,I117084,I117127,);
not I_6735 (I117076,I117127);
not I_6736 (I117149,I117110);
nand I_6737 (I117166,I325263,I325251);
and I_6738 (I117183,I117166,I325254);
DFFARX1 I_6739 (I117183,I2595,I117084,I117209,);
not I_6740 (I117217,I117209);
DFFARX1 I_6741 (I325272,I2595,I117084,I117243,);
and I_6742 (I117251,I117243,I325248);
nand I_6743 (I117268,I117243,I325248);
nand I_6744 (I117055,I117217,I117268);
DFFARX1 I_6745 (I325266,I2595,I117084,I117308,);
nor I_6746 (I117316,I117308,I117251);
DFFARX1 I_6747 (I117316,I2595,I117084,I117049,);
nor I_6748 (I117064,I117308,I117209);
nand I_6749 (I117361,I325260,I325257);
and I_6750 (I117378,I117361,I325269);
DFFARX1 I_6751 (I117378,I2595,I117084,I117404,);
nor I_6752 (I117052,I117404,I117308);
not I_6753 (I117426,I117404);
nor I_6754 (I117443,I117426,I117217);
nor I_6755 (I117460,I117149,I117443);
DFFARX1 I_6756 (I117460,I2595,I117084,I117067,);
nor I_6757 (I117491,I117426,I117308);
nor I_6758 (I117508,I325248,I325257);
nor I_6759 (I117058,I117508,I117491);
not I_6760 (I117539,I117508);
nand I_6761 (I117061,I117268,I117539);
DFFARX1 I_6762 (I117508,I2595,I117084,I117073,);
DFFARX1 I_6763 (I117508,I2595,I117084,I117070,);
not I_6764 (I117628,I2602);
DFFARX1 I_6765 (I361408,I2595,I117628,I117654,);
DFFARX1 I_6766 (I117654,I2595,I117628,I117671,);
not I_6767 (I117620,I117671);
not I_6768 (I117693,I117654);
nand I_6769 (I117710,I361405,I361402);
and I_6770 (I117727,I117710,I361390);
DFFARX1 I_6771 (I117727,I2595,I117628,I117753,);
not I_6772 (I117761,I117753);
DFFARX1 I_6773 (I361414,I2595,I117628,I117787,);
and I_6774 (I117795,I117787,I361399);
nand I_6775 (I117812,I117787,I361399);
nand I_6776 (I117599,I117761,I117812);
DFFARX1 I_6777 (I361393,I2595,I117628,I117852,);
nor I_6778 (I117860,I117852,I117795);
DFFARX1 I_6779 (I117860,I2595,I117628,I117593,);
nor I_6780 (I117608,I117852,I117753);
nand I_6781 (I117905,I361390,I361396);
and I_6782 (I117922,I117905,I361411);
DFFARX1 I_6783 (I117922,I2595,I117628,I117948,);
nor I_6784 (I117596,I117948,I117852);
not I_6785 (I117970,I117948);
nor I_6786 (I117987,I117970,I117761);
nor I_6787 (I118004,I117693,I117987);
DFFARX1 I_6788 (I118004,I2595,I117628,I117611,);
nor I_6789 (I118035,I117970,I117852);
nor I_6790 (I118052,I361393,I361396);
nor I_6791 (I117602,I118052,I118035);
not I_6792 (I118083,I118052);
nand I_6793 (I117605,I117812,I118083);
DFFARX1 I_6794 (I118052,I2595,I117628,I117617,);
DFFARX1 I_6795 (I118052,I2595,I117628,I117614,);
not I_6796 (I118172,I2602);
DFFARX1 I_6797 (I250409,I2595,I118172,I118198,);
DFFARX1 I_6798 (I118198,I2595,I118172,I118215,);
not I_6799 (I118164,I118215);
not I_6800 (I118237,I118198);
nand I_6801 (I118254,I250403,I250400);
and I_6802 (I118271,I118254,I250415);
DFFARX1 I_6803 (I118271,I2595,I118172,I118297,);
not I_6804 (I118305,I118297);
DFFARX1 I_6805 (I250403,I2595,I118172,I118331,);
and I_6806 (I118339,I118331,I250397);
nand I_6807 (I118356,I118331,I250397);
nand I_6808 (I118143,I118305,I118356);
DFFARX1 I_6809 (I250397,I2595,I118172,I118396,);
nor I_6810 (I118404,I118396,I118339);
DFFARX1 I_6811 (I118404,I2595,I118172,I118137,);
nor I_6812 (I118152,I118396,I118297);
nand I_6813 (I118449,I250412,I250406);
and I_6814 (I118466,I118449,I250400);
DFFARX1 I_6815 (I118466,I2595,I118172,I118492,);
nor I_6816 (I118140,I118492,I118396);
not I_6817 (I118514,I118492);
nor I_6818 (I118531,I118514,I118305);
nor I_6819 (I118548,I118237,I118531);
DFFARX1 I_6820 (I118548,I2595,I118172,I118155,);
nor I_6821 (I118579,I118514,I118396);
nor I_6822 (I118596,I250418,I250406);
nor I_6823 (I118146,I118596,I118579);
not I_6824 (I118627,I118596);
nand I_6825 (I118149,I118356,I118627);
DFFARX1 I_6826 (I118596,I2595,I118172,I118161,);
DFFARX1 I_6827 (I118596,I2595,I118172,I118158,);
not I_6828 (I118716,I2602);
DFFARX1 I_6829 (I224067,I2595,I118716,I118742,);
DFFARX1 I_6830 (I118742,I2595,I118716,I118759,);
not I_6831 (I118708,I118759);
not I_6832 (I118781,I118742);
nand I_6833 (I118798,I224088,I224079);
and I_6834 (I118815,I118798,I224067);
DFFARX1 I_6835 (I118815,I2595,I118716,I118841,);
not I_6836 (I118849,I118841);
DFFARX1 I_6837 (I224073,I2595,I118716,I118875,);
and I_6838 (I118883,I118875,I224070);
nand I_6839 (I118900,I118875,I224070);
nand I_6840 (I118687,I118849,I118900);
DFFARX1 I_6841 (I224064,I2595,I118716,I118940,);
nor I_6842 (I118948,I118940,I118883);
DFFARX1 I_6843 (I118948,I2595,I118716,I118681,);
nor I_6844 (I118696,I118940,I118841);
nand I_6845 (I118993,I224064,I224076);
and I_6846 (I119010,I118993,I224085);
DFFARX1 I_6847 (I119010,I2595,I118716,I119036,);
nor I_6848 (I118684,I119036,I118940);
not I_6849 (I119058,I119036);
nor I_6850 (I119075,I119058,I118849);
nor I_6851 (I119092,I118781,I119075);
DFFARX1 I_6852 (I119092,I2595,I118716,I118699,);
nor I_6853 (I119123,I119058,I118940);
nor I_6854 (I119140,I224082,I224076);
nor I_6855 (I118690,I119140,I119123);
not I_6856 (I119171,I119140);
nand I_6857 (I118693,I118900,I119171);
DFFARX1 I_6858 (I119140,I2595,I118716,I118705,);
DFFARX1 I_6859 (I119140,I2595,I118716,I118702,);
not I_6860 (I119260,I2602);
DFFARX1 I_6861 (I181873,I2595,I119260,I119286,);
DFFARX1 I_6862 (I119286,I2595,I119260,I119303,);
not I_6863 (I119252,I119303);
not I_6864 (I119325,I119286);
nand I_6865 (I119342,I181894,I181885);
and I_6866 (I119359,I119342,I181873);
DFFARX1 I_6867 (I119359,I2595,I119260,I119385,);
not I_6868 (I119393,I119385);
DFFARX1 I_6869 (I181879,I2595,I119260,I119419,);
and I_6870 (I119427,I119419,I181876);
nand I_6871 (I119444,I119419,I181876);
nand I_6872 (I119231,I119393,I119444);
DFFARX1 I_6873 (I181870,I2595,I119260,I119484,);
nor I_6874 (I119492,I119484,I119427);
DFFARX1 I_6875 (I119492,I2595,I119260,I119225,);
nor I_6876 (I119240,I119484,I119385);
nand I_6877 (I119537,I181870,I181882);
and I_6878 (I119554,I119537,I181891);
DFFARX1 I_6879 (I119554,I2595,I119260,I119580,);
nor I_6880 (I119228,I119580,I119484);
not I_6881 (I119602,I119580);
nor I_6882 (I119619,I119602,I119393);
nor I_6883 (I119636,I119325,I119619);
DFFARX1 I_6884 (I119636,I2595,I119260,I119243,);
nor I_6885 (I119667,I119602,I119484);
nor I_6886 (I119684,I181888,I181882);
nor I_6887 (I119234,I119684,I119667);
not I_6888 (I119715,I119684);
nand I_6889 (I119237,I119444,I119715);
DFFARX1 I_6890 (I119684,I2595,I119260,I119249,);
DFFARX1 I_6891 (I119684,I2595,I119260,I119246,);
not I_6892 (I119804,I2602);
DFFARX1 I_6893 (I245666,I2595,I119804,I119830,);
DFFARX1 I_6894 (I119830,I2595,I119804,I119847,);
not I_6895 (I119796,I119847);
not I_6896 (I119869,I119830);
nand I_6897 (I119886,I245660,I245657);
and I_6898 (I119903,I119886,I245672);
DFFARX1 I_6899 (I119903,I2595,I119804,I119929,);
not I_6900 (I119937,I119929);
DFFARX1 I_6901 (I245660,I2595,I119804,I119963,);
and I_6902 (I119971,I119963,I245654);
nand I_6903 (I119988,I119963,I245654);
nand I_6904 (I119775,I119937,I119988);
DFFARX1 I_6905 (I245654,I2595,I119804,I120028,);
nor I_6906 (I120036,I120028,I119971);
DFFARX1 I_6907 (I120036,I2595,I119804,I119769,);
nor I_6908 (I119784,I120028,I119929);
nand I_6909 (I120081,I245669,I245663);
and I_6910 (I120098,I120081,I245657);
DFFARX1 I_6911 (I120098,I2595,I119804,I120124,);
nor I_6912 (I119772,I120124,I120028);
not I_6913 (I120146,I120124);
nor I_6914 (I120163,I120146,I119937);
nor I_6915 (I120180,I119869,I120163);
DFFARX1 I_6916 (I120180,I2595,I119804,I119787,);
nor I_6917 (I120211,I120146,I120028);
nor I_6918 (I120228,I245675,I245663);
nor I_6919 (I119778,I120228,I120211);
not I_6920 (I120259,I120228);
nand I_6921 (I119781,I119988,I120259);
DFFARX1 I_6922 (I120228,I2595,I119804,I119793,);
DFFARX1 I_6923 (I120228,I2595,I119804,I119790,);
not I_6924 (I120348,I2602);
DFFARX1 I_6925 (I355681,I2595,I120348,I120374,);
DFFARX1 I_6926 (I120374,I2595,I120348,I120391,);
not I_6927 (I120340,I120391);
not I_6928 (I120413,I120374);
nand I_6929 (I120430,I355693,I355696);
and I_6930 (I120447,I120430,I355699);
DFFARX1 I_6931 (I120447,I2595,I120348,I120473,);
not I_6932 (I120481,I120473);
DFFARX1 I_6933 (I355684,I2595,I120348,I120507,);
and I_6934 (I120515,I120507,I355690);
nand I_6935 (I120532,I120507,I355690);
nand I_6936 (I120319,I120481,I120532);
DFFARX1 I_6937 (I355678,I2595,I120348,I120572,);
nor I_6938 (I120580,I120572,I120515);
DFFARX1 I_6939 (I120580,I2595,I120348,I120313,);
nor I_6940 (I120328,I120572,I120473);
nand I_6941 (I120625,I355681,I355702);
and I_6942 (I120642,I120625,I355687);
DFFARX1 I_6943 (I120642,I2595,I120348,I120668,);
nor I_6944 (I120316,I120668,I120572);
not I_6945 (I120690,I120668);
nor I_6946 (I120707,I120690,I120481);
nor I_6947 (I120724,I120413,I120707);
DFFARX1 I_6948 (I120724,I2595,I120348,I120331,);
nor I_6949 (I120755,I120690,I120572);
nor I_6950 (I120772,I355678,I355702);
nor I_6951 (I120322,I120772,I120755);
not I_6952 (I120803,I120772);
nand I_6953 (I120325,I120532,I120803);
DFFARX1 I_6954 (I120772,I2595,I120348,I120337,);
DFFARX1 I_6955 (I120772,I2595,I120348,I120334,);
not I_6956 (I120892,I2602);
DFFARX1 I_6957 (I225801,I2595,I120892,I120918,);
DFFARX1 I_6958 (I120918,I2595,I120892,I120935,);
not I_6959 (I120884,I120935);
not I_6960 (I120957,I120918);
nand I_6961 (I120974,I225822,I225813);
and I_6962 (I120991,I120974,I225801);
DFFARX1 I_6963 (I120991,I2595,I120892,I121017,);
not I_6964 (I121025,I121017);
DFFARX1 I_6965 (I225807,I2595,I120892,I121051,);
and I_6966 (I121059,I121051,I225804);
nand I_6967 (I121076,I121051,I225804);
nand I_6968 (I120863,I121025,I121076);
DFFARX1 I_6969 (I225798,I2595,I120892,I121116,);
nor I_6970 (I121124,I121116,I121059);
DFFARX1 I_6971 (I121124,I2595,I120892,I120857,);
nor I_6972 (I120872,I121116,I121017);
nand I_6973 (I121169,I225798,I225810);
and I_6974 (I121186,I121169,I225819);
DFFARX1 I_6975 (I121186,I2595,I120892,I121212,);
nor I_6976 (I120860,I121212,I121116);
not I_6977 (I121234,I121212);
nor I_6978 (I121251,I121234,I121025);
nor I_6979 (I121268,I120957,I121251);
DFFARX1 I_6980 (I121268,I2595,I120892,I120875,);
nor I_6981 (I121299,I121234,I121116);
nor I_6982 (I121316,I225816,I225810);
nor I_6983 (I120866,I121316,I121299);
not I_6984 (I121347,I121316);
nand I_6985 (I120869,I121076,I121347);
DFFARX1 I_6986 (I121316,I2595,I120892,I120881,);
DFFARX1 I_6987 (I121316,I2595,I120892,I120878,);
not I_6988 (I121436,I2602);
DFFARX1 I_6989 (I362564,I2595,I121436,I121462,);
DFFARX1 I_6990 (I121462,I2595,I121436,I121479,);
not I_6991 (I121428,I121479);
not I_6992 (I121501,I121462);
nand I_6993 (I121518,I362561,I362558);
and I_6994 (I121535,I121518,I362546);
DFFARX1 I_6995 (I121535,I2595,I121436,I121561,);
not I_6996 (I121569,I121561);
DFFARX1 I_6997 (I362570,I2595,I121436,I121595,);
and I_6998 (I121603,I121595,I362555);
nand I_6999 (I121620,I121595,I362555);
nand I_7000 (I121407,I121569,I121620);
DFFARX1 I_7001 (I362549,I2595,I121436,I121660,);
nor I_7002 (I121668,I121660,I121603);
DFFARX1 I_7003 (I121668,I2595,I121436,I121401,);
nor I_7004 (I121416,I121660,I121561);
nand I_7005 (I121713,I362546,I362552);
and I_7006 (I121730,I121713,I362567);
DFFARX1 I_7007 (I121730,I2595,I121436,I121756,);
nor I_7008 (I121404,I121756,I121660);
not I_7009 (I121778,I121756);
nor I_7010 (I121795,I121778,I121569);
nor I_7011 (I121812,I121501,I121795);
DFFARX1 I_7012 (I121812,I2595,I121436,I121419,);
nor I_7013 (I121843,I121778,I121660);
nor I_7014 (I121860,I362549,I362552);
nor I_7015 (I121410,I121860,I121843);
not I_7016 (I121891,I121860);
nand I_7017 (I121413,I121620,I121891);
DFFARX1 I_7018 (I121860,I2595,I121436,I121425,);
DFFARX1 I_7019 (I121860,I2595,I121436,I121422,);
not I_7020 (I121980,I2602);
DFFARX1 I_7021 (I348609,I2595,I121980,I122006,);
DFFARX1 I_7022 (I122006,I2595,I121980,I122023,);
not I_7023 (I121972,I122023);
not I_7024 (I122045,I122006);
nand I_7025 (I122062,I348621,I348624);
and I_7026 (I122079,I122062,I348627);
DFFARX1 I_7027 (I122079,I2595,I121980,I122105,);
not I_7028 (I122113,I122105);
DFFARX1 I_7029 (I348612,I2595,I121980,I122139,);
and I_7030 (I122147,I122139,I348618);
nand I_7031 (I122164,I122139,I348618);
nand I_7032 (I121951,I122113,I122164);
DFFARX1 I_7033 (I348606,I2595,I121980,I122204,);
nor I_7034 (I122212,I122204,I122147);
DFFARX1 I_7035 (I122212,I2595,I121980,I121945,);
nor I_7036 (I121960,I122204,I122105);
nand I_7037 (I122257,I348609,I348630);
and I_7038 (I122274,I122257,I348615);
DFFARX1 I_7039 (I122274,I2595,I121980,I122300,);
nor I_7040 (I121948,I122300,I122204);
not I_7041 (I122322,I122300);
nor I_7042 (I122339,I122322,I122113);
nor I_7043 (I122356,I122045,I122339);
DFFARX1 I_7044 (I122356,I2595,I121980,I121963,);
nor I_7045 (I122387,I122322,I122204);
nor I_7046 (I122404,I348606,I348630);
nor I_7047 (I121954,I122404,I122387);
not I_7048 (I122435,I122404);
nand I_7049 (I121957,I122164,I122435);
DFFARX1 I_7050 (I122404,I2595,I121980,I121969,);
DFFARX1 I_7051 (I122404,I2595,I121980,I121966,);
not I_7052 (I122524,I2602);
DFFARX1 I_7053 (I111205,I2595,I122524,I122550,);
DFFARX1 I_7054 (I122550,I2595,I122524,I122567,);
not I_7055 (I122516,I122567);
not I_7056 (I122589,I122550);
nand I_7057 (I122606,I111184,I111208);
and I_7058 (I122623,I122606,I111211);
DFFARX1 I_7059 (I122623,I2595,I122524,I122649,);
not I_7060 (I122657,I122649);
DFFARX1 I_7061 (I111193,I2595,I122524,I122683,);
and I_7062 (I122691,I122683,I111199);
nand I_7063 (I122708,I122683,I111199);
nand I_7064 (I122495,I122657,I122708);
DFFARX1 I_7065 (I111187,I2595,I122524,I122748,);
nor I_7066 (I122756,I122748,I122691);
DFFARX1 I_7067 (I122756,I2595,I122524,I122489,);
nor I_7068 (I122504,I122748,I122649);
nand I_7069 (I122801,I111196,I111184);
and I_7070 (I122818,I122801,I111190);
DFFARX1 I_7071 (I122818,I2595,I122524,I122844,);
nor I_7072 (I122492,I122844,I122748);
not I_7073 (I122866,I122844);
nor I_7074 (I122883,I122866,I122657);
nor I_7075 (I122900,I122589,I122883);
DFFARX1 I_7076 (I122900,I2595,I122524,I122507,);
nor I_7077 (I122931,I122866,I122748);
nor I_7078 (I122948,I111202,I111184);
nor I_7079 (I122498,I122948,I122931);
not I_7080 (I122979,I122948);
nand I_7081 (I122501,I122708,I122979);
DFFARX1 I_7082 (I122948,I2595,I122524,I122513,);
DFFARX1 I_7083 (I122948,I2595,I122524,I122510,);
not I_7084 (I123068,I2602);
DFFARX1 I_7085 (I297742,I2595,I123068,I123094,);
DFFARX1 I_7086 (I123094,I2595,I123068,I123111,);
not I_7087 (I123060,I123111);
not I_7088 (I123133,I123094);
nand I_7089 (I123150,I297742,I297760);
and I_7090 (I123167,I123150,I297754);
DFFARX1 I_7091 (I123167,I2595,I123068,I123193,);
not I_7092 (I123201,I123193);
DFFARX1 I_7093 (I297748,I2595,I123068,I123227,);
and I_7094 (I123235,I123227,I297757);
nand I_7095 (I123252,I123227,I297757);
nand I_7096 (I123039,I123201,I123252);
DFFARX1 I_7097 (I297745,I2595,I123068,I123292,);
nor I_7098 (I123300,I123292,I123235);
DFFARX1 I_7099 (I123300,I2595,I123068,I123033,);
nor I_7100 (I123048,I123292,I123193);
nand I_7101 (I123345,I297745,I297763);
and I_7102 (I123362,I123345,I297748);
DFFARX1 I_7103 (I123362,I2595,I123068,I123388,);
nor I_7104 (I123036,I123388,I123292);
not I_7105 (I123410,I123388);
nor I_7106 (I123427,I123410,I123201);
nor I_7107 (I123444,I123133,I123427);
DFFARX1 I_7108 (I123444,I2595,I123068,I123051,);
nor I_7109 (I123475,I123410,I123292);
nor I_7110 (I123492,I297751,I297763);
nor I_7111 (I123042,I123492,I123475);
not I_7112 (I123523,I123492);
nand I_7113 (I123045,I123252,I123523);
DFFARX1 I_7114 (I123492,I2595,I123068,I123057,);
DFFARX1 I_7115 (I123492,I2595,I123068,I123054,);
not I_7116 (I123612,I2602);
DFFARX1 I_7117 (I168001,I2595,I123612,I123638,);
DFFARX1 I_7118 (I123638,I2595,I123612,I123655,);
not I_7119 (I123604,I123655);
not I_7120 (I123677,I123638);
nand I_7121 (I123694,I167998,I168019);
and I_7122 (I123711,I123694,I168022);
DFFARX1 I_7123 (I123711,I2595,I123612,I123737,);
not I_7124 (I123745,I123737);
DFFARX1 I_7125 (I168007,I2595,I123612,I123771,);
and I_7126 (I123779,I123771,I168010);
nand I_7127 (I123796,I123771,I168010);
nand I_7128 (I123583,I123745,I123796);
DFFARX1 I_7129 (I168013,I2595,I123612,I123836,);
nor I_7130 (I123844,I123836,I123779);
DFFARX1 I_7131 (I123844,I2595,I123612,I123577,);
nor I_7132 (I123592,I123836,I123737);
nand I_7133 (I123889,I167998,I168004);
and I_7134 (I123906,I123889,I168016);
DFFARX1 I_7135 (I123906,I2595,I123612,I123932,);
nor I_7136 (I123580,I123932,I123836);
not I_7137 (I123954,I123932);
nor I_7138 (I123971,I123954,I123745);
nor I_7139 (I123988,I123677,I123971);
DFFARX1 I_7140 (I123988,I2595,I123612,I123595,);
nor I_7141 (I124019,I123954,I123836);
nor I_7142 (I124036,I168001,I168004);
nor I_7143 (I123586,I124036,I124019);
not I_7144 (I124067,I124036);
nand I_7145 (I123589,I123796,I124067);
DFFARX1 I_7146 (I124036,I2595,I123612,I123601,);
DFFARX1 I_7147 (I124036,I2595,I123612,I123598,);
not I_7148 (I124156,I2602);
DFFARX1 I_7149 (I152888,I2595,I124156,I124182,);
DFFARX1 I_7150 (I124182,I2595,I124156,I124199,);
not I_7151 (I124148,I124199);
not I_7152 (I124221,I124182);
nand I_7153 (I124238,I152891,I152909);
and I_7154 (I124255,I124238,I152897);
DFFARX1 I_7155 (I124255,I2595,I124156,I124281,);
not I_7156 (I124289,I124281);
DFFARX1 I_7157 (I152888,I2595,I124156,I124315,);
and I_7158 (I124323,I124315,I152906);
nand I_7159 (I124340,I124315,I152906);
nand I_7160 (I124127,I124289,I124340);
DFFARX1 I_7161 (I152900,I2595,I124156,I124380,);
nor I_7162 (I124388,I124380,I124323);
DFFARX1 I_7163 (I124388,I2595,I124156,I124121,);
nor I_7164 (I124136,I124380,I124281);
nand I_7165 (I124433,I152903,I152885);
and I_7166 (I124450,I124433,I152894);
DFFARX1 I_7167 (I124450,I2595,I124156,I124476,);
nor I_7168 (I124124,I124476,I124380);
not I_7169 (I124498,I124476);
nor I_7170 (I124515,I124498,I124289);
nor I_7171 (I124532,I124221,I124515);
DFFARX1 I_7172 (I124532,I2595,I124156,I124139,);
nor I_7173 (I124563,I124498,I124380);
nor I_7174 (I124580,I152885,I152885);
nor I_7175 (I124130,I124580,I124563);
not I_7176 (I124611,I124580);
nand I_7177 (I124133,I124340,I124611);
DFFARX1 I_7178 (I124580,I2595,I124156,I124145,);
DFFARX1 I_7179 (I124580,I2595,I124156,I124142,);
not I_7180 (I124700,I2602);
DFFARX1 I_7181 (I331609,I2595,I124700,I124726,);
DFFARX1 I_7182 (I124726,I2595,I124700,I124743,);
not I_7183 (I124692,I124743);
not I_7184 (I124765,I124726);
nand I_7185 (I124782,I331621,I331609);
and I_7186 (I124799,I124782,I331612);
DFFARX1 I_7187 (I124799,I2595,I124700,I124825,);
not I_7188 (I124833,I124825);
DFFARX1 I_7189 (I331630,I2595,I124700,I124859,);
and I_7190 (I124867,I124859,I331606);
nand I_7191 (I124884,I124859,I331606);
nand I_7192 (I124671,I124833,I124884);
DFFARX1 I_7193 (I331624,I2595,I124700,I124924,);
nor I_7194 (I124932,I124924,I124867);
DFFARX1 I_7195 (I124932,I2595,I124700,I124665,);
nor I_7196 (I124680,I124924,I124825);
nand I_7197 (I124977,I331618,I331615);
and I_7198 (I124994,I124977,I331627);
DFFARX1 I_7199 (I124994,I2595,I124700,I125020,);
nor I_7200 (I124668,I125020,I124924);
not I_7201 (I125042,I125020);
nor I_7202 (I125059,I125042,I124833);
nor I_7203 (I125076,I124765,I125059);
DFFARX1 I_7204 (I125076,I2595,I124700,I124683,);
nor I_7205 (I125107,I125042,I124924);
nor I_7206 (I125124,I331606,I331615);
nor I_7207 (I124674,I125124,I125107);
not I_7208 (I125155,I125124);
nand I_7209 (I124677,I124884,I125155);
DFFARX1 I_7210 (I125124,I2595,I124700,I124689,);
DFFARX1 I_7211 (I125124,I2595,I124700,I124686,);
not I_7212 (I125244,I2602);
DFFARX1 I_7213 (I142178,I2595,I125244,I125270,);
DFFARX1 I_7214 (I125270,I2595,I125244,I125287,);
not I_7215 (I125236,I125287);
not I_7216 (I125309,I125270);
nand I_7217 (I125326,I142181,I142199);
and I_7218 (I125343,I125326,I142187);
DFFARX1 I_7219 (I125343,I2595,I125244,I125369,);
not I_7220 (I125377,I125369);
DFFARX1 I_7221 (I142178,I2595,I125244,I125403,);
and I_7222 (I125411,I125403,I142196);
nand I_7223 (I125428,I125403,I142196);
nand I_7224 (I125215,I125377,I125428);
DFFARX1 I_7225 (I142190,I2595,I125244,I125468,);
nor I_7226 (I125476,I125468,I125411);
DFFARX1 I_7227 (I125476,I2595,I125244,I125209,);
nor I_7228 (I125224,I125468,I125369);
nand I_7229 (I125521,I142193,I142175);
and I_7230 (I125538,I125521,I142184);
DFFARX1 I_7231 (I125538,I2595,I125244,I125564,);
nor I_7232 (I125212,I125564,I125468);
not I_7233 (I125586,I125564);
nor I_7234 (I125603,I125586,I125377);
nor I_7235 (I125620,I125309,I125603);
DFFARX1 I_7236 (I125620,I2595,I125244,I125227,);
nor I_7237 (I125651,I125586,I125468);
nor I_7238 (I125668,I142175,I142175);
nor I_7239 (I125218,I125668,I125651);
not I_7240 (I125699,I125668);
nand I_7241 (I125221,I125428,I125699);
DFFARX1 I_7242 (I125668,I2595,I125244,I125233,);
DFFARX1 I_7243 (I125668,I2595,I125244,I125230,);
not I_7244 (I125788,I2602);
DFFARX1 I_7245 (I382480,I2595,I125788,I125814,);
DFFARX1 I_7246 (I125814,I2595,I125788,I125831,);
not I_7247 (I125780,I125831);
not I_7248 (I125853,I125814);
nand I_7249 (I125870,I382456,I382477);
and I_7250 (I125887,I125870,I382474);
DFFARX1 I_7251 (I125887,I2595,I125788,I125913,);
not I_7252 (I125921,I125913);
DFFARX1 I_7253 (I382453,I2595,I125788,I125947,);
and I_7254 (I125955,I125947,I382465);
nand I_7255 (I125972,I125947,I382465);
nand I_7256 (I125759,I125921,I125972);
DFFARX1 I_7257 (I382468,I2595,I125788,I126012,);
nor I_7258 (I126020,I126012,I125955);
DFFARX1 I_7259 (I126020,I2595,I125788,I125753,);
nor I_7260 (I125768,I126012,I125913);
nand I_7261 (I126065,I382471,I382459);
and I_7262 (I126082,I126065,I382462);
DFFARX1 I_7263 (I126082,I2595,I125788,I126108,);
nor I_7264 (I125756,I126108,I126012);
not I_7265 (I126130,I126108);
nor I_7266 (I126147,I126130,I125921);
nor I_7267 (I126164,I125853,I126147);
DFFARX1 I_7268 (I126164,I2595,I125788,I125771,);
nor I_7269 (I126195,I126130,I126012);
nor I_7270 (I126212,I382453,I382459);
nor I_7271 (I125762,I126212,I126195);
not I_7272 (I126243,I126212);
nand I_7273 (I125765,I125972,I126243);
DFFARX1 I_7274 (I126212,I2595,I125788,I125777,);
DFFARX1 I_7275 (I126212,I2595,I125788,I125774,);
not I_7276 (I126332,I2602);
DFFARX1 I_7277 (I91706,I2595,I126332,I126358,);
DFFARX1 I_7278 (I126358,I2595,I126332,I126375,);
not I_7279 (I126324,I126375);
not I_7280 (I126397,I126358);
nand I_7281 (I126414,I91685,I91709);
and I_7282 (I126431,I126414,I91712);
DFFARX1 I_7283 (I126431,I2595,I126332,I126457,);
not I_7284 (I126465,I126457);
DFFARX1 I_7285 (I91694,I2595,I126332,I126491,);
and I_7286 (I126499,I126491,I91700);
nand I_7287 (I126516,I126491,I91700);
nand I_7288 (I126303,I126465,I126516);
DFFARX1 I_7289 (I91688,I2595,I126332,I126556,);
nor I_7290 (I126564,I126556,I126499);
DFFARX1 I_7291 (I126564,I2595,I126332,I126297,);
nor I_7292 (I126312,I126556,I126457);
nand I_7293 (I126609,I91697,I91685);
and I_7294 (I126626,I126609,I91691);
DFFARX1 I_7295 (I126626,I2595,I126332,I126652,);
nor I_7296 (I126300,I126652,I126556);
not I_7297 (I126674,I126652);
nor I_7298 (I126691,I126674,I126465);
nor I_7299 (I126708,I126397,I126691);
DFFARX1 I_7300 (I126708,I2595,I126332,I126315,);
nor I_7301 (I126739,I126674,I126556);
nor I_7302 (I126756,I91703,I91685);
nor I_7303 (I126306,I126756,I126739);
not I_7304 (I126787,I126756);
nand I_7305 (I126309,I126516,I126787);
DFFARX1 I_7306 (I126756,I2595,I126332,I126321,);
DFFARX1 I_7307 (I126756,I2595,I126332,I126318,);
not I_7308 (I126876,I2602);
DFFARX1 I_7309 (I171469,I2595,I126876,I126902,);
DFFARX1 I_7310 (I126902,I2595,I126876,I126919,);
not I_7311 (I126868,I126919);
not I_7312 (I126941,I126902);
nand I_7313 (I126958,I171466,I171487);
and I_7314 (I126975,I126958,I171490);
DFFARX1 I_7315 (I126975,I2595,I126876,I127001,);
not I_7316 (I127009,I127001);
DFFARX1 I_7317 (I171475,I2595,I126876,I127035,);
and I_7318 (I127043,I127035,I171478);
nand I_7319 (I127060,I127035,I171478);
nand I_7320 (I126847,I127009,I127060);
DFFARX1 I_7321 (I171481,I2595,I126876,I127100,);
nor I_7322 (I127108,I127100,I127043);
DFFARX1 I_7323 (I127108,I2595,I126876,I126841,);
nor I_7324 (I126856,I127100,I127001);
nand I_7325 (I127153,I171466,I171472);
and I_7326 (I127170,I127153,I171484);
DFFARX1 I_7327 (I127170,I2595,I126876,I127196,);
nor I_7328 (I126844,I127196,I127100);
not I_7329 (I127218,I127196);
nor I_7330 (I127235,I127218,I127009);
nor I_7331 (I127252,I126941,I127235);
DFFARX1 I_7332 (I127252,I2595,I126876,I126859,);
nor I_7333 (I127283,I127218,I127100);
nor I_7334 (I127300,I171469,I171472);
nor I_7335 (I126850,I127300,I127283);
not I_7336 (I127331,I127300);
nand I_7337 (I126853,I127060,I127331);
DFFARX1 I_7338 (I127300,I2595,I126876,I126865,);
DFFARX1 I_7339 (I127300,I2595,I126876,I126862,);
not I_7340 (I127420,I2602);
DFFARX1 I_7341 (I102773,I2595,I127420,I127446,);
DFFARX1 I_7342 (I127446,I2595,I127420,I127463,);
not I_7343 (I127412,I127463);
not I_7344 (I127485,I127446);
nand I_7345 (I127502,I102752,I102776);
and I_7346 (I127519,I127502,I102779);
DFFARX1 I_7347 (I127519,I2595,I127420,I127545,);
not I_7348 (I127553,I127545);
DFFARX1 I_7349 (I102761,I2595,I127420,I127579,);
and I_7350 (I127587,I127579,I102767);
nand I_7351 (I127604,I127579,I102767);
nand I_7352 (I127391,I127553,I127604);
DFFARX1 I_7353 (I102755,I2595,I127420,I127644,);
nor I_7354 (I127652,I127644,I127587);
DFFARX1 I_7355 (I127652,I2595,I127420,I127385,);
nor I_7356 (I127400,I127644,I127545);
nand I_7357 (I127697,I102764,I102752);
and I_7358 (I127714,I127697,I102758);
DFFARX1 I_7359 (I127714,I2595,I127420,I127740,);
nor I_7360 (I127388,I127740,I127644);
not I_7361 (I127762,I127740);
nor I_7362 (I127779,I127762,I127553);
nor I_7363 (I127796,I127485,I127779);
DFFARX1 I_7364 (I127796,I2595,I127420,I127403,);
nor I_7365 (I127827,I127762,I127644);
nor I_7366 (I127844,I102770,I102752);
nor I_7367 (I127394,I127844,I127827);
not I_7368 (I127875,I127844);
nand I_7369 (I127397,I127604,I127875);
DFFARX1 I_7370 (I127844,I2595,I127420,I127409,);
DFFARX1 I_7371 (I127844,I2595,I127420,I127406,);
not I_7372 (I127964,I2602);
DFFARX1 I_7373 (I3813,I2595,I127964,I127990,);
DFFARX1 I_7374 (I127990,I2595,I127964,I128007,);
not I_7375 (I127956,I128007);
not I_7376 (I128029,I127990);
nand I_7377 (I128046,I3816,I3804);
and I_7378 (I128063,I128046,I3810);
DFFARX1 I_7379 (I128063,I2595,I127964,I128089,);
not I_7380 (I128097,I128089);
DFFARX1 I_7381 (I3798,I2595,I127964,I128123,);
and I_7382 (I128131,I128123,I3795);
nand I_7383 (I128148,I128123,I3795);
nand I_7384 (I127935,I128097,I128148);
DFFARX1 I_7385 (I3801,I2595,I127964,I128188,);
nor I_7386 (I128196,I128188,I128131);
DFFARX1 I_7387 (I128196,I2595,I127964,I127929,);
nor I_7388 (I127944,I128188,I128089);
nand I_7389 (I128241,I3801,I3798);
and I_7390 (I128258,I128241,I3795);
DFFARX1 I_7391 (I128258,I2595,I127964,I128284,);
nor I_7392 (I127932,I128284,I128188);
not I_7393 (I128306,I128284);
nor I_7394 (I128323,I128306,I128097);
nor I_7395 (I128340,I128029,I128323);
DFFARX1 I_7396 (I128340,I2595,I127964,I127947,);
nor I_7397 (I128371,I128306,I128188);
nor I_7398 (I128388,I3807,I3798);
nor I_7399 (I127938,I128388,I128371);
not I_7400 (I128419,I128388);
nand I_7401 (I127941,I128148,I128419);
DFFARX1 I_7402 (I128388,I2595,I127964,I127953,);
DFFARX1 I_7403 (I128388,I2595,I127964,I127950,);
not I_7404 (I128508,I2602);
DFFARX1 I_7405 (I71702,I2595,I128508,I128534,);
DFFARX1 I_7406 (I128534,I2595,I128508,I128551,);
not I_7407 (I128500,I128551);
not I_7408 (I128573,I128534);
nand I_7409 (I128590,I71714,I71693);
and I_7410 (I128607,I128590,I71696);
DFFARX1 I_7411 (I128607,I2595,I128508,I128633,);
not I_7412 (I128641,I128633);
DFFARX1 I_7413 (I71705,I2595,I128508,I128667,);
and I_7414 (I128675,I128667,I71717);
nand I_7415 (I128692,I128667,I71717);
nand I_7416 (I128479,I128641,I128692);
DFFARX1 I_7417 (I71711,I2595,I128508,I128732,);
nor I_7418 (I128740,I128732,I128675);
DFFARX1 I_7419 (I128740,I2595,I128508,I128473,);
nor I_7420 (I128488,I128732,I128633);
nand I_7421 (I128785,I71699,I71696);
and I_7422 (I128802,I128785,I71708);
DFFARX1 I_7423 (I128802,I2595,I128508,I128828,);
nor I_7424 (I128476,I128828,I128732);
not I_7425 (I128850,I128828);
nor I_7426 (I128867,I128850,I128641);
nor I_7427 (I128884,I128573,I128867);
DFFARX1 I_7428 (I128884,I2595,I128508,I128491,);
nor I_7429 (I128915,I128850,I128732);
nor I_7430 (I128932,I71693,I71696);
nor I_7431 (I128482,I128932,I128915);
not I_7432 (I128963,I128932);
nand I_7433 (I128485,I128692,I128963);
DFFARX1 I_7434 (I128932,I2595,I128508,I128497,);
DFFARX1 I_7435 (I128932,I2595,I128508,I128494,);
not I_7436 (I129052,I2602);
DFFARX1 I_7437 (I197479,I2595,I129052,I129078,);
DFFARX1 I_7438 (I129078,I2595,I129052,I129095,);
not I_7439 (I129044,I129095);
not I_7440 (I129117,I129078);
nand I_7441 (I129134,I197500,I197491);
and I_7442 (I129151,I129134,I197479);
DFFARX1 I_7443 (I129151,I2595,I129052,I129177,);
not I_7444 (I129185,I129177);
DFFARX1 I_7445 (I197485,I2595,I129052,I129211,);
and I_7446 (I129219,I129211,I197482);
nand I_7447 (I129236,I129211,I197482);
nand I_7448 (I129023,I129185,I129236);
DFFARX1 I_7449 (I197476,I2595,I129052,I129276,);
nor I_7450 (I129284,I129276,I129219);
DFFARX1 I_7451 (I129284,I2595,I129052,I129017,);
nor I_7452 (I129032,I129276,I129177);
nand I_7453 (I129329,I197476,I197488);
and I_7454 (I129346,I129329,I197497);
DFFARX1 I_7455 (I129346,I2595,I129052,I129372,);
nor I_7456 (I129020,I129372,I129276);
not I_7457 (I129394,I129372);
nor I_7458 (I129411,I129394,I129185);
nor I_7459 (I129428,I129117,I129411);
DFFARX1 I_7460 (I129428,I2595,I129052,I129035,);
nor I_7461 (I129459,I129394,I129276);
nor I_7462 (I129476,I197494,I197488);
nor I_7463 (I129026,I129476,I129459);
not I_7464 (I129507,I129476);
nand I_7465 (I129029,I129236,I129507);
DFFARX1 I_7466 (I129476,I2595,I129052,I129041,);
DFFARX1 I_7467 (I129476,I2595,I129052,I129038,);
not I_7468 (I129596,I2602);
DFFARX1 I_7469 (I85909,I2595,I129596,I129622,);
DFFARX1 I_7470 (I129622,I2595,I129596,I129639,);
not I_7471 (I129588,I129639);
not I_7472 (I129661,I129622);
nand I_7473 (I129678,I85888,I85912);
and I_7474 (I129695,I129678,I85915);
DFFARX1 I_7475 (I129695,I2595,I129596,I129721,);
not I_7476 (I129729,I129721);
DFFARX1 I_7477 (I85897,I2595,I129596,I129755,);
and I_7478 (I129763,I129755,I85903);
nand I_7479 (I129780,I129755,I85903);
nand I_7480 (I129567,I129729,I129780);
DFFARX1 I_7481 (I85891,I2595,I129596,I129820,);
nor I_7482 (I129828,I129820,I129763);
DFFARX1 I_7483 (I129828,I2595,I129596,I129561,);
nor I_7484 (I129576,I129820,I129721);
nand I_7485 (I129873,I85900,I85888);
and I_7486 (I129890,I129873,I85894);
DFFARX1 I_7487 (I129890,I2595,I129596,I129916,);
nor I_7488 (I129564,I129916,I129820);
not I_7489 (I129938,I129916);
nor I_7490 (I129955,I129938,I129729);
nor I_7491 (I129972,I129661,I129955);
DFFARX1 I_7492 (I129972,I2595,I129596,I129579,);
nor I_7493 (I130003,I129938,I129820);
nor I_7494 (I130020,I85906,I85888);
nor I_7495 (I129570,I130020,I130003);
not I_7496 (I130051,I130020);
nand I_7497 (I129573,I129780,I130051);
DFFARX1 I_7498 (I130020,I2595,I129596,I129585,);
DFFARX1 I_7499 (I130020,I2595,I129596,I129582,);
not I_7500 (I130140,I2602);
DFFARX1 I_7501 (I29250,I2595,I130140,I130166,);
DFFARX1 I_7502 (I130166,I2595,I130140,I130183,);
not I_7503 (I130132,I130183);
not I_7504 (I130205,I130166);
nand I_7505 (I130222,I29265,I29244);
and I_7506 (I130239,I130222,I29247);
DFFARX1 I_7507 (I130239,I2595,I130140,I130265,);
not I_7508 (I130273,I130265);
DFFARX1 I_7509 (I29253,I2595,I130140,I130299,);
and I_7510 (I130307,I130299,I29247);
nand I_7511 (I130324,I130299,I29247);
nand I_7512 (I130111,I130273,I130324);
DFFARX1 I_7513 (I29262,I2595,I130140,I130364,);
nor I_7514 (I130372,I130364,I130307);
DFFARX1 I_7515 (I130372,I2595,I130140,I130105,);
nor I_7516 (I130120,I130364,I130265);
nand I_7517 (I130417,I29244,I29259);
and I_7518 (I130434,I130417,I29256);
DFFARX1 I_7519 (I130434,I2595,I130140,I130460,);
nor I_7520 (I130108,I130460,I130364);
not I_7521 (I130482,I130460);
nor I_7522 (I130499,I130482,I130273);
nor I_7523 (I130516,I130205,I130499);
DFFARX1 I_7524 (I130516,I2595,I130140,I130123,);
nor I_7525 (I130547,I130482,I130364);
nor I_7526 (I130564,I29268,I29259);
nor I_7527 (I130114,I130564,I130547);
not I_7528 (I130595,I130564);
nand I_7529 (I130117,I130324,I130595);
DFFARX1 I_7530 (I130564,I2595,I130140,I130129,);
DFFARX1 I_7531 (I130564,I2595,I130140,I130126,);
not I_7532 (I130684,I2602);
DFFARX1 I_7533 (I235126,I2595,I130684,I130710,);
DFFARX1 I_7534 (I130710,I2595,I130684,I130727,);
not I_7535 (I130676,I130727);
not I_7536 (I130749,I130710);
nand I_7537 (I130766,I235120,I235117);
and I_7538 (I130783,I130766,I235132);
DFFARX1 I_7539 (I130783,I2595,I130684,I130809,);
not I_7540 (I130817,I130809);
DFFARX1 I_7541 (I235120,I2595,I130684,I130843,);
and I_7542 (I130851,I130843,I235114);
nand I_7543 (I130868,I130843,I235114);
nand I_7544 (I130655,I130817,I130868);
DFFARX1 I_7545 (I235114,I2595,I130684,I130908,);
nor I_7546 (I130916,I130908,I130851);
DFFARX1 I_7547 (I130916,I2595,I130684,I130649,);
nor I_7548 (I130664,I130908,I130809);
nand I_7549 (I130961,I235129,I235123);
and I_7550 (I130978,I130961,I235117);
DFFARX1 I_7551 (I130978,I2595,I130684,I131004,);
nor I_7552 (I130652,I131004,I130908);
not I_7553 (I131026,I131004);
nor I_7554 (I131043,I131026,I130817);
nor I_7555 (I131060,I130749,I131043);
DFFARX1 I_7556 (I131060,I2595,I130684,I130667,);
nor I_7557 (I131091,I131026,I130908);
nor I_7558 (I131108,I235135,I235123);
nor I_7559 (I130658,I131108,I131091);
not I_7560 (I131139,I131108);
nand I_7561 (I130661,I130868,I131139);
DFFARX1 I_7562 (I131108,I2595,I130684,I130673,);
DFFARX1 I_7563 (I131108,I2595,I130684,I130670,);
not I_7564 (I131228,I2602);
DFFARX1 I_7565 (I57422,I2595,I131228,I131254,);
DFFARX1 I_7566 (I131254,I2595,I131228,I131271,);
not I_7567 (I131220,I131271);
not I_7568 (I131293,I131254);
nand I_7569 (I131310,I57434,I57413);
and I_7570 (I131327,I131310,I57416);
DFFARX1 I_7571 (I131327,I2595,I131228,I131353,);
not I_7572 (I131361,I131353);
DFFARX1 I_7573 (I57425,I2595,I131228,I131387,);
and I_7574 (I131395,I131387,I57437);
nand I_7575 (I131412,I131387,I57437);
nand I_7576 (I131199,I131361,I131412);
DFFARX1 I_7577 (I57431,I2595,I131228,I131452,);
nor I_7578 (I131460,I131452,I131395);
DFFARX1 I_7579 (I131460,I2595,I131228,I131193,);
nor I_7580 (I131208,I131452,I131353);
nand I_7581 (I131505,I57419,I57416);
and I_7582 (I131522,I131505,I57428);
DFFARX1 I_7583 (I131522,I2595,I131228,I131548,);
nor I_7584 (I131196,I131548,I131452);
not I_7585 (I131570,I131548);
nor I_7586 (I131587,I131570,I131361);
nor I_7587 (I131604,I131293,I131587);
DFFARX1 I_7588 (I131604,I2595,I131228,I131211,);
nor I_7589 (I131635,I131570,I131452);
nor I_7590 (I131652,I57413,I57416);
nor I_7591 (I131202,I131652,I131635);
not I_7592 (I131683,I131652);
nand I_7593 (I131205,I131412,I131683);
DFFARX1 I_7594 (I131652,I2595,I131228,I131217,);
DFFARX1 I_7595 (I131652,I2595,I131228,I131214,);
not I_7596 (I131772,I2602);
DFFARX1 I_7597 (I237234,I2595,I131772,I131798,);
DFFARX1 I_7598 (I131798,I2595,I131772,I131815,);
not I_7599 (I131764,I131815);
not I_7600 (I131837,I131798);
nand I_7601 (I131854,I237228,I237225);
and I_7602 (I131871,I131854,I237240);
DFFARX1 I_7603 (I131871,I2595,I131772,I131897,);
not I_7604 (I131905,I131897);
DFFARX1 I_7605 (I237228,I2595,I131772,I131931,);
and I_7606 (I131939,I131931,I237222);
nand I_7607 (I131956,I131931,I237222);
nand I_7608 (I131743,I131905,I131956);
DFFARX1 I_7609 (I237222,I2595,I131772,I131996,);
nor I_7610 (I132004,I131996,I131939);
DFFARX1 I_7611 (I132004,I2595,I131772,I131737,);
nor I_7612 (I131752,I131996,I131897);
nand I_7613 (I132049,I237237,I237231);
and I_7614 (I132066,I132049,I237225);
DFFARX1 I_7615 (I132066,I2595,I131772,I132092,);
nor I_7616 (I131740,I132092,I131996);
not I_7617 (I132114,I132092);
nor I_7618 (I132131,I132114,I131905);
nor I_7619 (I132148,I131837,I132131);
DFFARX1 I_7620 (I132148,I2595,I131772,I131755,);
nor I_7621 (I132179,I132114,I131996);
nor I_7622 (I132196,I237243,I237231);
nor I_7623 (I131746,I132196,I132179);
not I_7624 (I132227,I132196);
nand I_7625 (I131749,I131956,I132227);
DFFARX1 I_7626 (I132196,I2595,I131772,I131761,);
DFFARX1 I_7627 (I132196,I2595,I131772,I131758,);
not I_7628 (I132316,I2602);
DFFARX1 I_7629 (I83274,I2595,I132316,I132342,);
DFFARX1 I_7630 (I132342,I2595,I132316,I132359,);
not I_7631 (I132308,I132359);
not I_7632 (I132381,I132342);
nand I_7633 (I132398,I83253,I83277);
and I_7634 (I132415,I132398,I83280);
DFFARX1 I_7635 (I132415,I2595,I132316,I132441,);
not I_7636 (I132449,I132441);
DFFARX1 I_7637 (I83262,I2595,I132316,I132475,);
and I_7638 (I132483,I132475,I83268);
nand I_7639 (I132500,I132475,I83268);
nand I_7640 (I132287,I132449,I132500);
DFFARX1 I_7641 (I83256,I2595,I132316,I132540,);
nor I_7642 (I132548,I132540,I132483);
DFFARX1 I_7643 (I132548,I2595,I132316,I132281,);
nor I_7644 (I132296,I132540,I132441);
nand I_7645 (I132593,I83265,I83253);
and I_7646 (I132610,I132593,I83259);
DFFARX1 I_7647 (I132610,I2595,I132316,I132636,);
nor I_7648 (I132284,I132636,I132540);
not I_7649 (I132658,I132636);
nor I_7650 (I132675,I132658,I132449);
nor I_7651 (I132692,I132381,I132675);
DFFARX1 I_7652 (I132692,I2595,I132316,I132299,);
nor I_7653 (I132723,I132658,I132540);
nor I_7654 (I132740,I83271,I83253);
nor I_7655 (I132290,I132740,I132723);
not I_7656 (I132771,I132740);
nand I_7657 (I132293,I132500,I132771);
DFFARX1 I_7658 (I132740,I2595,I132316,I132305,);
DFFARX1 I_7659 (I132740,I2595,I132316,I132302,);
not I_7660 (I132860,I2602);
DFFARX1 I_7661 (I368344,I2595,I132860,I132886,);
DFFARX1 I_7662 (I132886,I2595,I132860,I132903,);
not I_7663 (I132852,I132903);
not I_7664 (I132925,I132886);
nand I_7665 (I132942,I368341,I368338);
and I_7666 (I132959,I132942,I368326);
DFFARX1 I_7667 (I132959,I2595,I132860,I132985,);
not I_7668 (I132993,I132985);
DFFARX1 I_7669 (I368350,I2595,I132860,I133019,);
and I_7670 (I133027,I133019,I368335);
nand I_7671 (I133044,I133019,I368335);
nand I_7672 (I132831,I132993,I133044);
DFFARX1 I_7673 (I368329,I2595,I132860,I133084,);
nor I_7674 (I133092,I133084,I133027);
DFFARX1 I_7675 (I133092,I2595,I132860,I132825,);
nor I_7676 (I132840,I133084,I132985);
nand I_7677 (I133137,I368326,I368332);
and I_7678 (I133154,I133137,I368347);
DFFARX1 I_7679 (I133154,I2595,I132860,I133180,);
nor I_7680 (I132828,I133180,I133084);
not I_7681 (I133202,I133180);
nor I_7682 (I133219,I133202,I132993);
nor I_7683 (I133236,I132925,I133219);
DFFARX1 I_7684 (I133236,I2595,I132860,I132843,);
nor I_7685 (I133267,I133202,I133084);
nor I_7686 (I133284,I368329,I368332);
nor I_7687 (I132834,I133284,I133267);
not I_7688 (I133315,I133284);
nand I_7689 (I132837,I133044,I133315);
DFFARX1 I_7690 (I133284,I2595,I132860,I132849,);
DFFARX1 I_7691 (I133284,I2595,I132860,I132846,);
not I_7692 (I133404,I2602);
DFFARX1 I_7693 (I367188,I2595,I133404,I133430,);
DFFARX1 I_7694 (I133430,I2595,I133404,I133447,);
not I_7695 (I133396,I133447);
not I_7696 (I133469,I133430);
nand I_7697 (I133486,I367185,I367182);
and I_7698 (I133503,I133486,I367170);
DFFARX1 I_7699 (I133503,I2595,I133404,I133529,);
not I_7700 (I133537,I133529);
DFFARX1 I_7701 (I367194,I2595,I133404,I133563,);
and I_7702 (I133571,I133563,I367179);
nand I_7703 (I133588,I133563,I367179);
nand I_7704 (I133375,I133537,I133588);
DFFARX1 I_7705 (I367173,I2595,I133404,I133628,);
nor I_7706 (I133636,I133628,I133571);
DFFARX1 I_7707 (I133636,I2595,I133404,I133369,);
nor I_7708 (I133384,I133628,I133529);
nand I_7709 (I133681,I367170,I367176);
and I_7710 (I133698,I133681,I367191);
DFFARX1 I_7711 (I133698,I2595,I133404,I133724,);
nor I_7712 (I133372,I133724,I133628);
not I_7713 (I133746,I133724);
nor I_7714 (I133763,I133746,I133537);
nor I_7715 (I133780,I133469,I133763);
DFFARX1 I_7716 (I133780,I2595,I133404,I133387,);
nor I_7717 (I133811,I133746,I133628);
nor I_7718 (I133828,I367173,I367176);
nor I_7719 (I133378,I133828,I133811);
not I_7720 (I133859,I133828);
nand I_7721 (I133381,I133588,I133859);
DFFARX1 I_7722 (I133828,I2595,I133404,I133393,);
DFFARX1 I_7723 (I133828,I2595,I133404,I133390,);
not I_7724 (I133948,I2602);
DFFARX1 I_7725 (I216553,I2595,I133948,I133974,);
DFFARX1 I_7726 (I133974,I2595,I133948,I133991,);
not I_7727 (I133940,I133991);
not I_7728 (I134013,I133974);
nand I_7729 (I134030,I216574,I216565);
and I_7730 (I134047,I134030,I216553);
DFFARX1 I_7731 (I134047,I2595,I133948,I134073,);
not I_7732 (I134081,I134073);
DFFARX1 I_7733 (I216559,I2595,I133948,I134107,);
and I_7734 (I134115,I134107,I216556);
nand I_7735 (I134132,I134107,I216556);
nand I_7736 (I133919,I134081,I134132);
DFFARX1 I_7737 (I216550,I2595,I133948,I134172,);
nor I_7738 (I134180,I134172,I134115);
DFFARX1 I_7739 (I134180,I2595,I133948,I133913,);
nor I_7740 (I133928,I134172,I134073);
nand I_7741 (I134225,I216550,I216562);
and I_7742 (I134242,I134225,I216571);
DFFARX1 I_7743 (I134242,I2595,I133948,I134268,);
nor I_7744 (I133916,I134268,I134172);
not I_7745 (I134290,I134268);
nor I_7746 (I134307,I134290,I134081);
nor I_7747 (I134324,I134013,I134307);
DFFARX1 I_7748 (I134324,I2595,I133948,I133931,);
nor I_7749 (I134355,I134290,I134172);
nor I_7750 (I134372,I216568,I216562);
nor I_7751 (I133922,I134372,I134355);
not I_7752 (I134403,I134372);
nand I_7753 (I133925,I134132,I134403);
DFFARX1 I_7754 (I134372,I2595,I133948,I133937,);
DFFARX1 I_7755 (I134372,I2595,I133948,I133934,);
not I_7756 (I134492,I2602);
DFFARX1 I_7757 (I209039,I2595,I134492,I134518,);
DFFARX1 I_7758 (I134518,I2595,I134492,I134535,);
not I_7759 (I134484,I134535);
not I_7760 (I134557,I134518);
nand I_7761 (I134574,I209060,I209051);
and I_7762 (I134591,I134574,I209039);
DFFARX1 I_7763 (I134591,I2595,I134492,I134617,);
not I_7764 (I134625,I134617);
DFFARX1 I_7765 (I209045,I2595,I134492,I134651,);
and I_7766 (I134659,I134651,I209042);
nand I_7767 (I134676,I134651,I209042);
nand I_7768 (I134463,I134625,I134676);
DFFARX1 I_7769 (I209036,I2595,I134492,I134716,);
nor I_7770 (I134724,I134716,I134659);
DFFARX1 I_7771 (I134724,I2595,I134492,I134457,);
nor I_7772 (I134472,I134716,I134617);
nand I_7773 (I134769,I209036,I209048);
and I_7774 (I134786,I134769,I209057);
DFFARX1 I_7775 (I134786,I2595,I134492,I134812,);
nor I_7776 (I134460,I134812,I134716);
not I_7777 (I134834,I134812);
nor I_7778 (I134851,I134834,I134625);
nor I_7779 (I134868,I134557,I134851);
DFFARX1 I_7780 (I134868,I2595,I134492,I134475,);
nor I_7781 (I134899,I134834,I134716);
nor I_7782 (I134916,I209054,I209048);
nor I_7783 (I134466,I134916,I134899);
not I_7784 (I134947,I134916);
nand I_7785 (I134469,I134676,I134947);
DFFARX1 I_7786 (I134916,I2595,I134492,I134481,);
DFFARX1 I_7787 (I134916,I2595,I134492,I134478,);
not I_7788 (I135036,I2602);
DFFARX1 I_7789 (I174937,I2595,I135036,I135062,);
DFFARX1 I_7790 (I135062,I2595,I135036,I135079,);
not I_7791 (I135028,I135079);
not I_7792 (I135101,I135062);
nand I_7793 (I135118,I174934,I174955);
and I_7794 (I135135,I135118,I174958);
DFFARX1 I_7795 (I135135,I2595,I135036,I135161,);
not I_7796 (I135169,I135161);
DFFARX1 I_7797 (I174943,I2595,I135036,I135195,);
and I_7798 (I135203,I135195,I174946);
nand I_7799 (I135220,I135195,I174946);
nand I_7800 (I135007,I135169,I135220);
DFFARX1 I_7801 (I174949,I2595,I135036,I135260,);
nor I_7802 (I135268,I135260,I135203);
DFFARX1 I_7803 (I135268,I2595,I135036,I135001,);
nor I_7804 (I135016,I135260,I135161);
nand I_7805 (I135313,I174934,I174940);
and I_7806 (I135330,I135313,I174952);
DFFARX1 I_7807 (I135330,I2595,I135036,I135356,);
nor I_7808 (I135004,I135356,I135260);
not I_7809 (I135378,I135356);
nor I_7810 (I135395,I135378,I135169);
nor I_7811 (I135412,I135101,I135395);
DFFARX1 I_7812 (I135412,I2595,I135036,I135019,);
nor I_7813 (I135443,I135378,I135260);
nor I_7814 (I135460,I174937,I174940);
nor I_7815 (I135010,I135460,I135443);
not I_7816 (I135491,I135460);
nand I_7817 (I135013,I135220,I135491);
DFFARX1 I_7818 (I135460,I2595,I135036,I135025,);
DFFARX1 I_7819 (I135460,I2595,I135036,I135022,);
not I_7820 (I135580,I2602);
DFFARX1 I_7821 (I105935,I2595,I135580,I135606,);
DFFARX1 I_7822 (I135606,I2595,I135580,I135623,);
not I_7823 (I135572,I135623);
not I_7824 (I135645,I135606);
nand I_7825 (I135662,I105914,I105938);
and I_7826 (I135679,I135662,I105941);
DFFARX1 I_7827 (I135679,I2595,I135580,I135705,);
not I_7828 (I135713,I135705);
DFFARX1 I_7829 (I105923,I2595,I135580,I135739,);
and I_7830 (I135747,I135739,I105929);
nand I_7831 (I135764,I135739,I105929);
nand I_7832 (I135551,I135713,I135764);
DFFARX1 I_7833 (I105917,I2595,I135580,I135804,);
nor I_7834 (I135812,I135804,I135747);
DFFARX1 I_7835 (I135812,I2595,I135580,I135545,);
nor I_7836 (I135560,I135804,I135705);
nand I_7837 (I135857,I105926,I105914);
and I_7838 (I135874,I135857,I105920);
DFFARX1 I_7839 (I135874,I2595,I135580,I135900,);
nor I_7840 (I135548,I135900,I135804);
not I_7841 (I135922,I135900);
nor I_7842 (I135939,I135922,I135713);
nor I_7843 (I135956,I135645,I135939);
DFFARX1 I_7844 (I135956,I2595,I135580,I135563,);
nor I_7845 (I135987,I135922,I135804);
nor I_7846 (I136004,I105932,I105914);
nor I_7847 (I135554,I136004,I135987);
not I_7848 (I136035,I136004);
nand I_7849 (I135557,I135764,I136035);
DFFARX1 I_7850 (I136004,I2595,I135580,I135569,);
DFFARX1 I_7851 (I136004,I2595,I135580,I135566,);
not I_7852 (I136124,I2602);
DFFARX1 I_7853 (I173781,I2595,I136124,I136150,);
DFFARX1 I_7854 (I136150,I2595,I136124,I136167,);
not I_7855 (I136116,I136167);
not I_7856 (I136189,I136150);
nand I_7857 (I136206,I173778,I173799);
and I_7858 (I136223,I136206,I173802);
DFFARX1 I_7859 (I136223,I2595,I136124,I136249,);
not I_7860 (I136257,I136249);
DFFARX1 I_7861 (I173787,I2595,I136124,I136283,);
and I_7862 (I136291,I136283,I173790);
nand I_7863 (I136308,I136283,I173790);
nand I_7864 (I136095,I136257,I136308);
DFFARX1 I_7865 (I173793,I2595,I136124,I136348,);
nor I_7866 (I136356,I136348,I136291);
DFFARX1 I_7867 (I136356,I2595,I136124,I136089,);
nor I_7868 (I136104,I136348,I136249);
nand I_7869 (I136401,I173778,I173784);
and I_7870 (I136418,I136401,I173796);
DFFARX1 I_7871 (I136418,I2595,I136124,I136444,);
nor I_7872 (I136092,I136444,I136348);
not I_7873 (I136466,I136444);
nor I_7874 (I136483,I136466,I136257);
nor I_7875 (I136500,I136189,I136483);
DFFARX1 I_7876 (I136500,I2595,I136124,I136107,);
nor I_7877 (I136531,I136466,I136348);
nor I_7878 (I136548,I173781,I173784);
nor I_7879 (I136098,I136548,I136531);
not I_7880 (I136579,I136548);
nand I_7881 (I136101,I136308,I136579);
DFFARX1 I_7882 (I136548,I2595,I136124,I136113,);
DFFARX1 I_7883 (I136548,I2595,I136124,I136110,);
not I_7884 (I136668,I2602);
DFFARX1 I_7885 (I233018,I2595,I136668,I136694,);
DFFARX1 I_7886 (I136694,I2595,I136668,I136711,);
not I_7887 (I136660,I136711);
not I_7888 (I136733,I136694);
nand I_7889 (I136750,I233012,I233009);
and I_7890 (I136767,I136750,I233024);
DFFARX1 I_7891 (I136767,I2595,I136668,I136793,);
not I_7892 (I136801,I136793);
DFFARX1 I_7893 (I233012,I2595,I136668,I136827,);
and I_7894 (I136835,I136827,I233006);
nand I_7895 (I136852,I136827,I233006);
nand I_7896 (I136639,I136801,I136852);
DFFARX1 I_7897 (I233006,I2595,I136668,I136892,);
nor I_7898 (I136900,I136892,I136835);
DFFARX1 I_7899 (I136900,I2595,I136668,I136633,);
nor I_7900 (I136648,I136892,I136793);
nand I_7901 (I136945,I233021,I233015);
and I_7902 (I136962,I136945,I233009);
DFFARX1 I_7903 (I136962,I2595,I136668,I136988,);
nor I_7904 (I136636,I136988,I136892);
not I_7905 (I137010,I136988);
nor I_7906 (I137027,I137010,I136801);
nor I_7907 (I137044,I136733,I137027);
DFFARX1 I_7908 (I137044,I2595,I136668,I136651,);
nor I_7909 (I137075,I137010,I136892);
nor I_7910 (I137092,I233027,I233015);
nor I_7911 (I136642,I137092,I137075);
not I_7912 (I137123,I137092);
nand I_7913 (I136645,I136852,I137123);
DFFARX1 I_7914 (I137092,I2595,I136668,I136657,);
DFFARX1 I_7915 (I137092,I2595,I136668,I136654,);
not I_7916 (I137212,I2602);
DFFARX1 I_7917 (I37682,I2595,I137212,I137238,);
DFFARX1 I_7918 (I137238,I2595,I137212,I137255,);
not I_7919 (I137204,I137255);
not I_7920 (I137277,I137238);
nand I_7921 (I137294,I37697,I37676);
and I_7922 (I137311,I137294,I37679);
DFFARX1 I_7923 (I137311,I2595,I137212,I137337,);
not I_7924 (I137345,I137337);
DFFARX1 I_7925 (I37685,I2595,I137212,I137371,);
and I_7926 (I137379,I137371,I37679);
nand I_7927 (I137396,I137371,I37679);
nand I_7928 (I137183,I137345,I137396);
DFFARX1 I_7929 (I37694,I2595,I137212,I137436,);
nor I_7930 (I137444,I137436,I137379);
DFFARX1 I_7931 (I137444,I2595,I137212,I137177,);
nor I_7932 (I137192,I137436,I137337);
nand I_7933 (I137489,I37676,I37691);
and I_7934 (I137506,I137489,I37688);
DFFARX1 I_7935 (I137506,I2595,I137212,I137532,);
nor I_7936 (I137180,I137532,I137436);
not I_7937 (I137554,I137532);
nor I_7938 (I137571,I137554,I137345);
nor I_7939 (I137588,I137277,I137571);
DFFARX1 I_7940 (I137588,I2595,I137212,I137195,);
nor I_7941 (I137619,I137554,I137436);
nor I_7942 (I137636,I37700,I37691);
nor I_7943 (I137186,I137636,I137619);
not I_7944 (I137667,I137636);
nand I_7945 (I137189,I137396,I137667);
DFFARX1 I_7946 (I137636,I2595,I137212,I137201,);
DFFARX1 I_7947 (I137636,I2595,I137212,I137198,);
not I_7948 (I137756,I2602);
DFFARX1 I_7949 (I307911,I2595,I137756,I137782,);
DFFARX1 I_7950 (I137782,I2595,I137756,I137799,);
not I_7951 (I137748,I137799);
not I_7952 (I137821,I137782);
nand I_7953 (I137838,I307923,I307911);
and I_7954 (I137855,I137838,I307914);
DFFARX1 I_7955 (I137855,I2595,I137756,I137881,);
not I_7956 (I137889,I137881);
DFFARX1 I_7957 (I307932,I2595,I137756,I137915,);
and I_7958 (I137923,I137915,I307908);
nand I_7959 (I137940,I137915,I307908);
nand I_7960 (I137727,I137889,I137940);
DFFARX1 I_7961 (I307926,I2595,I137756,I137980,);
nor I_7962 (I137988,I137980,I137923);
DFFARX1 I_7963 (I137988,I2595,I137756,I137721,);
nor I_7964 (I137736,I137980,I137881);
nand I_7965 (I138033,I307920,I307917);
and I_7966 (I138050,I138033,I307929);
DFFARX1 I_7967 (I138050,I2595,I137756,I138076,);
nor I_7968 (I137724,I138076,I137980);
not I_7969 (I138098,I138076);
nor I_7970 (I138115,I138098,I137889);
nor I_7971 (I138132,I137821,I138115);
DFFARX1 I_7972 (I138132,I2595,I137756,I137739,);
nor I_7973 (I138163,I138098,I137980);
nor I_7974 (I138180,I307908,I307917);
nor I_7975 (I137730,I138180,I138163);
not I_7976 (I138211,I138180);
nand I_7977 (I137733,I137940,I138211);
DFFARX1 I_7978 (I138180,I2595,I137756,I137745,);
DFFARX1 I_7979 (I138180,I2595,I137756,I137742,);
not I_7980 (I138300,I2602);
DFFARX1 I_7981 (I38736,I2595,I138300,I138326,);
DFFARX1 I_7982 (I138326,I2595,I138300,I138343,);
not I_7983 (I138292,I138343);
not I_7984 (I138365,I138326);
nand I_7985 (I138382,I38751,I38730);
and I_7986 (I138399,I138382,I38733);
DFFARX1 I_7987 (I138399,I2595,I138300,I138425,);
not I_7988 (I138433,I138425);
DFFARX1 I_7989 (I38739,I2595,I138300,I138459,);
and I_7990 (I138467,I138459,I38733);
nand I_7991 (I138484,I138459,I38733);
nand I_7992 (I138271,I138433,I138484);
DFFARX1 I_7993 (I38748,I2595,I138300,I138524,);
nor I_7994 (I138532,I138524,I138467);
DFFARX1 I_7995 (I138532,I2595,I138300,I138265,);
nor I_7996 (I138280,I138524,I138425);
nand I_7997 (I138577,I38730,I38745);
and I_7998 (I138594,I138577,I38742);
DFFARX1 I_7999 (I138594,I2595,I138300,I138620,);
nor I_8000 (I138268,I138620,I138524);
not I_8001 (I138642,I138620);
nor I_8002 (I138659,I138642,I138433);
nor I_8003 (I138676,I138365,I138659);
DFFARX1 I_8004 (I138676,I2595,I138300,I138283,);
nor I_8005 (I138707,I138642,I138524);
nor I_8006 (I138724,I38754,I38745);
nor I_8007 (I138274,I138724,I138707);
not I_8008 (I138755,I138724);
nand I_8009 (I138277,I138484,I138755);
DFFARX1 I_8010 (I138724,I2595,I138300,I138289,);
DFFARX1 I_8011 (I138724,I2595,I138300,I138286,);
not I_8012 (I138844,I2602);
DFFARX1 I_8013 (I247774,I2595,I138844,I138870,);
DFFARX1 I_8014 (I138870,I2595,I138844,I138887,);
not I_8015 (I138836,I138887);
not I_8016 (I138909,I138870);
nand I_8017 (I138926,I247768,I247765);
and I_8018 (I138943,I138926,I247780);
DFFARX1 I_8019 (I138943,I2595,I138844,I138969,);
not I_8020 (I138977,I138969);
DFFARX1 I_8021 (I247768,I2595,I138844,I139003,);
and I_8022 (I139011,I139003,I247762);
nand I_8023 (I139028,I139003,I247762);
nand I_8024 (I138815,I138977,I139028);
DFFARX1 I_8025 (I247762,I2595,I138844,I139068,);
nor I_8026 (I139076,I139068,I139011);
DFFARX1 I_8027 (I139076,I2595,I138844,I138809,);
nor I_8028 (I138824,I139068,I138969);
nand I_8029 (I139121,I247777,I247771);
and I_8030 (I139138,I139121,I247765);
DFFARX1 I_8031 (I139138,I2595,I138844,I139164,);
nor I_8032 (I138812,I139164,I139068);
not I_8033 (I139186,I139164);
nor I_8034 (I139203,I139186,I138977);
nor I_8035 (I139220,I138909,I139203);
DFFARX1 I_8036 (I139220,I2595,I138844,I138827,);
nor I_8037 (I139251,I139186,I139068);
nor I_8038 (I139268,I247783,I247771);
nor I_8039 (I138818,I139268,I139251);
not I_8040 (I139299,I139268);
nand I_8041 (I138821,I139028,I139299);
DFFARX1 I_8042 (I139268,I2595,I138844,I138833,);
DFFARX1 I_8043 (I139268,I2595,I138844,I138830,);
not I_8044 (I139388,I2602);
DFFARX1 I_8045 (I1628,I2595,I139388,I139414,);
DFFARX1 I_8046 (I139414,I2595,I139388,I139431,);
not I_8047 (I139380,I139431);
not I_8048 (I139453,I139414);
nand I_8049 (I139470,I2116,I1700);
and I_8050 (I139487,I139470,I1364);
DFFARX1 I_8051 (I139487,I2595,I139388,I139513,);
not I_8052 (I139521,I139513);
DFFARX1 I_8053 (I1644,I2595,I139388,I139547,);
and I_8054 (I139555,I139547,I1756);
nand I_8055 (I139572,I139547,I1756);
nand I_8056 (I139359,I139521,I139572);
DFFARX1 I_8057 (I2260,I2595,I139388,I139612,);
nor I_8058 (I139620,I139612,I139555);
DFFARX1 I_8059 (I139620,I2595,I139388,I139353,);
nor I_8060 (I139368,I139612,I139513);
nand I_8061 (I139665,I2508,I2268);
and I_8062 (I139682,I139665,I2444);
DFFARX1 I_8063 (I139682,I2595,I139388,I139708,);
nor I_8064 (I139356,I139708,I139612);
not I_8065 (I139730,I139708);
nor I_8066 (I139747,I139730,I139521);
nor I_8067 (I139764,I139453,I139747);
DFFARX1 I_8068 (I139764,I2595,I139388,I139371,);
nor I_8069 (I139795,I139730,I139612);
nor I_8070 (I139812,I1636,I2268);
nor I_8071 (I139362,I139812,I139795);
not I_8072 (I139843,I139812);
nand I_8073 (I139365,I139572,I139843);
DFFARX1 I_8074 (I139812,I2595,I139388,I139377,);
DFFARX1 I_8075 (I139812,I2595,I139388,I139374,);
not I_8076 (I139932,I2602);
DFFARX1 I_8077 (I211351,I2595,I139932,I139958,);
DFFARX1 I_8078 (I139958,I2595,I139932,I139975,);
not I_8079 (I139924,I139975);
not I_8080 (I139997,I139958);
nand I_8081 (I140014,I211372,I211363);
and I_8082 (I140031,I140014,I211351);
DFFARX1 I_8083 (I140031,I2595,I139932,I140057,);
not I_8084 (I140065,I140057);
DFFARX1 I_8085 (I211357,I2595,I139932,I140091,);
and I_8086 (I140099,I140091,I211354);
nand I_8087 (I140116,I140091,I211354);
nand I_8088 (I139903,I140065,I140116);
DFFARX1 I_8089 (I211348,I2595,I139932,I140156,);
nor I_8090 (I140164,I140156,I140099);
DFFARX1 I_8091 (I140164,I2595,I139932,I139897,);
nor I_8092 (I139912,I140156,I140057);
nand I_8093 (I140209,I211348,I211360);
and I_8094 (I140226,I140209,I211369);
DFFARX1 I_8095 (I140226,I2595,I139932,I140252,);
nor I_8096 (I139900,I140252,I140156);
not I_8097 (I140274,I140252);
nor I_8098 (I140291,I140274,I140065);
nor I_8099 (I140308,I139997,I140291);
DFFARX1 I_8100 (I140308,I2595,I139932,I139915,);
nor I_8101 (I140339,I140274,I140156);
nor I_8102 (I140356,I211366,I211360);
nor I_8103 (I139906,I140356,I140339);
not I_8104 (I140387,I140356);
nand I_8105 (I139909,I140116,I140387);
DFFARX1 I_8106 (I140356,I2595,I139932,I139921,);
DFFARX1 I_8107 (I140356,I2595,I139932,I139918,);
not I_8108 (I140476,I2602);
DFFARX1 I_8109 (I178983,I2595,I140476,I140502,);
DFFARX1 I_8110 (I140502,I2595,I140476,I140519,);
not I_8111 (I140468,I140519);
not I_8112 (I140541,I140502);
nand I_8113 (I140558,I178980,I179001);
and I_8114 (I140575,I140558,I179004);
DFFARX1 I_8115 (I140575,I2595,I140476,I140601,);
not I_8116 (I140609,I140601);
DFFARX1 I_8117 (I178989,I2595,I140476,I140635,);
and I_8118 (I140643,I140635,I178992);
nand I_8119 (I140660,I140635,I178992);
nand I_8120 (I140447,I140609,I140660);
DFFARX1 I_8121 (I178995,I2595,I140476,I140700,);
nor I_8122 (I140708,I140700,I140643);
DFFARX1 I_8123 (I140708,I2595,I140476,I140441,);
nor I_8124 (I140456,I140700,I140601);
nand I_8125 (I140753,I178980,I178986);
and I_8126 (I140770,I140753,I178998);
DFFARX1 I_8127 (I140770,I2595,I140476,I140796,);
nor I_8128 (I140444,I140796,I140700);
not I_8129 (I140818,I140796);
nor I_8130 (I140835,I140818,I140609);
nor I_8131 (I140852,I140541,I140835);
DFFARX1 I_8132 (I140852,I2595,I140476,I140459,);
nor I_8133 (I140883,I140818,I140700);
nor I_8134 (I140900,I178983,I178986);
nor I_8135 (I140450,I140900,I140883);
not I_8136 (I140931,I140900);
nand I_8137 (I140453,I140660,I140931);
DFFARX1 I_8138 (I140900,I2595,I140476,I140465,);
DFFARX1 I_8139 (I140900,I2595,I140476,I140462,);
not I_8140 (I141017,I2602);
DFFARX1 I_8141 (I7374,I2595,I141017,I141043,);
DFFARX1 I_8142 (I141043,I2595,I141017,I141060,);
not I_8143 (I141009,I141060);
DFFARX1 I_8144 (I7365,I2595,I141017,I141091,);
not I_8145 (I141099,I7368);
nor I_8146 (I141116,I141043,I141099);
not I_8147 (I141133,I7380);
not I_8148 (I141150,I7365);
nand I_8149 (I141167,I141150,I7380);
nor I_8150 (I141184,I141099,I141167);
nor I_8151 (I141201,I141091,I141184);
DFFARX1 I_8152 (I141150,I2595,I141017,I141006,);
nor I_8153 (I141232,I7365,I7371);
nand I_8154 (I141249,I141232,I7383);
nor I_8155 (I141266,I141249,I141133);
nand I_8156 (I140991,I141266,I7368);
DFFARX1 I_8157 (I141249,I2595,I141017,I141003,);
nand I_8158 (I141311,I141133,I7365);
nor I_8159 (I141328,I141133,I7365);
nand I_8160 (I140997,I141116,I141328);
not I_8161 (I141359,I7386);
nor I_8162 (I141376,I141359,I141311);
DFFARX1 I_8163 (I141376,I2595,I141017,I140985,);
nor I_8164 (I141407,I141359,I7368);
and I_8165 (I141424,I141407,I7377);
or I_8166 (I141441,I141424,I7371);
DFFARX1 I_8167 (I141441,I2595,I141017,I141467,);
nor I_8168 (I141475,I141467,I141091);
nor I_8169 (I140994,I141043,I141475);
not I_8170 (I141506,I141467);
nor I_8171 (I141523,I141506,I141201);
DFFARX1 I_8172 (I141523,I2595,I141017,I141000,);
nand I_8173 (I141554,I141506,I141133);
nor I_8174 (I140988,I141359,I141554);
not I_8175 (I141612,I2602);
DFFARX1 I_8176 (I18704,I2595,I141612,I141638,);
DFFARX1 I_8177 (I141638,I2595,I141612,I141655,);
not I_8178 (I141604,I141655);
DFFARX1 I_8179 (I18704,I2595,I141612,I141686,);
not I_8180 (I141694,I18719);
nor I_8181 (I141711,I141638,I141694);
not I_8182 (I141728,I18722);
not I_8183 (I141745,I18713);
nand I_8184 (I141762,I141745,I18722);
nor I_8185 (I141779,I141694,I141762);
nor I_8186 (I141796,I141686,I141779);
DFFARX1 I_8187 (I141745,I2595,I141612,I141601,);
nor I_8188 (I141827,I18713,I18725);
nand I_8189 (I141844,I141827,I18707);
nor I_8190 (I141861,I141844,I141728);
nand I_8191 (I141586,I141861,I18719);
DFFARX1 I_8192 (I141844,I2595,I141612,I141598,);
nand I_8193 (I141906,I141728,I18713);
nor I_8194 (I141923,I141728,I18713);
nand I_8195 (I141592,I141711,I141923);
not I_8196 (I141954,I18707);
nor I_8197 (I141971,I141954,I141906);
DFFARX1 I_8198 (I141971,I2595,I141612,I141580,);
nor I_8199 (I142002,I141954,I18716);
and I_8200 (I142019,I142002,I18710);
or I_8201 (I142036,I142019,I18728);
DFFARX1 I_8202 (I142036,I2595,I141612,I142062,);
nor I_8203 (I142070,I142062,I141686);
nor I_8204 (I141589,I141638,I142070);
not I_8205 (I142101,I142062);
nor I_8206 (I142118,I142101,I141796);
DFFARX1 I_8207 (I142118,I2595,I141612,I141595,);
nand I_8208 (I142149,I142101,I141728);
nor I_8209 (I141583,I141954,I142149);
not I_8210 (I142207,I2602);
DFFARX1 I_8211 (I124121,I2595,I142207,I142233,);
DFFARX1 I_8212 (I142233,I2595,I142207,I142250,);
not I_8213 (I142199,I142250);
DFFARX1 I_8214 (I124145,I2595,I142207,I142281,);
not I_8215 (I142289,I124124);
nor I_8216 (I142306,I142233,I142289);
not I_8217 (I142323,I124130);
not I_8218 (I142340,I124136);
nand I_8219 (I142357,I142340,I124130);
nor I_8220 (I142374,I142289,I142357);
nor I_8221 (I142391,I142281,I142374);
DFFARX1 I_8222 (I142340,I2595,I142207,I142196,);
nor I_8223 (I142422,I124136,I124148);
nand I_8224 (I142439,I142422,I124142);
nor I_8225 (I142456,I142439,I142323);
nand I_8226 (I142181,I142456,I124124);
DFFARX1 I_8227 (I142439,I2595,I142207,I142193,);
nand I_8228 (I142501,I142323,I124136);
nor I_8229 (I142518,I142323,I124136);
nand I_8230 (I142187,I142306,I142518);
not I_8231 (I142549,I124127);
nor I_8232 (I142566,I142549,I142501);
DFFARX1 I_8233 (I142566,I2595,I142207,I142175,);
nor I_8234 (I142597,I142549,I124121);
and I_8235 (I142614,I142597,I124139);
or I_8236 (I142631,I142614,I124133);
DFFARX1 I_8237 (I142631,I2595,I142207,I142657,);
nor I_8238 (I142665,I142657,I142281);
nor I_8239 (I142184,I142233,I142665);
not I_8240 (I142696,I142657);
nor I_8241 (I142713,I142696,I142391);
DFFARX1 I_8242 (I142713,I2595,I142207,I142190,);
nand I_8243 (I142744,I142696,I142323);
nor I_8244 (I142178,I142549,I142744);
not I_8245 (I142802,I2602);
DFFARX1 I_8246 (I204999,I2595,I142802,I142828,);
DFFARX1 I_8247 (I142828,I2595,I142802,I142845,);
not I_8248 (I142794,I142845);
DFFARX1 I_8249 (I204993,I2595,I142802,I142876,);
not I_8250 (I142884,I204990);
nor I_8251 (I142901,I142828,I142884);
not I_8252 (I142918,I205002);
not I_8253 (I142935,I205005);
nand I_8254 (I142952,I142935,I205002);
nor I_8255 (I142969,I142884,I142952);
nor I_8256 (I142986,I142876,I142969);
DFFARX1 I_8257 (I142935,I2595,I142802,I142791,);
nor I_8258 (I143017,I205005,I205014);
nand I_8259 (I143034,I143017,I205008);
nor I_8260 (I143051,I143034,I142918);
nand I_8261 (I142776,I143051,I204990);
DFFARX1 I_8262 (I143034,I2595,I142802,I142788,);
nand I_8263 (I143096,I142918,I205005);
nor I_8264 (I143113,I142918,I205005);
nand I_8265 (I142782,I142901,I143113);
not I_8266 (I143144,I204996);
nor I_8267 (I143161,I143144,I143096);
DFFARX1 I_8268 (I143161,I2595,I142802,I142770,);
nor I_8269 (I143192,I143144,I205011);
and I_8270 (I143209,I143192,I204990);
or I_8271 (I143226,I143209,I204993);
DFFARX1 I_8272 (I143226,I2595,I142802,I143252,);
nor I_8273 (I143260,I143252,I142876);
nor I_8274 (I142779,I142828,I143260);
not I_8275 (I143291,I143252);
nor I_8276 (I143308,I143291,I142986);
DFFARX1 I_8277 (I143308,I2595,I142802,I142785,);
nand I_8278 (I143339,I143291,I142918);
nor I_8279 (I142773,I143144,I143339);
not I_8280 (I143397,I2602);
DFFARX1 I_8281 (I271254,I2595,I143397,I143423,);
DFFARX1 I_8282 (I143423,I2595,I143397,I143440,);
not I_8283 (I143389,I143440);
DFFARX1 I_8284 (I271242,I2595,I143397,I143471,);
not I_8285 (I143479,I271239);
nor I_8286 (I143496,I143423,I143479);
not I_8287 (I143513,I271251);
not I_8288 (I143530,I271248);
nand I_8289 (I143547,I143530,I271251);
nor I_8290 (I143564,I143479,I143547);
nor I_8291 (I143581,I143471,I143564);
DFFARX1 I_8292 (I143530,I2595,I143397,I143386,);
nor I_8293 (I143612,I271248,I271257);
nand I_8294 (I143629,I143612,I271260);
nor I_8295 (I143646,I143629,I143513);
nand I_8296 (I143371,I143646,I271239);
DFFARX1 I_8297 (I143629,I2595,I143397,I143383,);
nand I_8298 (I143691,I143513,I271248);
nor I_8299 (I143708,I143513,I271248);
nand I_8300 (I143377,I143496,I143708);
not I_8301 (I143739,I271263);
nor I_8302 (I143756,I143739,I143691);
DFFARX1 I_8303 (I143756,I2595,I143397,I143365,);
nor I_8304 (I143787,I143739,I271266);
and I_8305 (I143804,I143787,I271245);
or I_8306 (I143821,I143804,I271239);
DFFARX1 I_8307 (I143821,I2595,I143397,I143847,);
nor I_8308 (I143855,I143847,I143471);
nor I_8309 (I143374,I143423,I143855);
not I_8310 (I143886,I143847);
nor I_8311 (I143903,I143886,I143581);
DFFARX1 I_8312 (I143903,I2595,I143397,I143380,);
nand I_8313 (I143934,I143886,I143513);
nor I_8314 (I143368,I143739,I143934);
not I_8315 (I143992,I2602);
DFFARX1 I_8316 (I125753,I2595,I143992,I144018,);
DFFARX1 I_8317 (I144018,I2595,I143992,I144035,);
not I_8318 (I143984,I144035);
DFFARX1 I_8319 (I125777,I2595,I143992,I144066,);
not I_8320 (I144074,I125756);
nor I_8321 (I144091,I144018,I144074);
not I_8322 (I144108,I125762);
not I_8323 (I144125,I125768);
nand I_8324 (I144142,I144125,I125762);
nor I_8325 (I144159,I144074,I144142);
nor I_8326 (I144176,I144066,I144159);
DFFARX1 I_8327 (I144125,I2595,I143992,I143981,);
nor I_8328 (I144207,I125768,I125780);
nand I_8329 (I144224,I144207,I125774);
nor I_8330 (I144241,I144224,I144108);
nand I_8331 (I143966,I144241,I125756);
DFFARX1 I_8332 (I144224,I2595,I143992,I143978,);
nand I_8333 (I144286,I144108,I125768);
nor I_8334 (I144303,I144108,I125768);
nand I_8335 (I143972,I144091,I144303);
not I_8336 (I144334,I125759);
nor I_8337 (I144351,I144334,I144286);
DFFARX1 I_8338 (I144351,I2595,I143992,I143960,);
nor I_8339 (I144382,I144334,I125753);
and I_8340 (I144399,I144382,I125771);
or I_8341 (I144416,I144399,I125765);
DFFARX1 I_8342 (I144416,I2595,I143992,I144442,);
nor I_8343 (I144450,I144442,I144066);
nor I_8344 (I143969,I144018,I144450);
not I_8345 (I144481,I144442);
nor I_8346 (I144498,I144481,I144176);
DFFARX1 I_8347 (I144498,I2595,I143992,I143975,);
nand I_8348 (I144529,I144481,I144108);
nor I_8349 (I143963,I144334,I144529);
not I_8350 (I144587,I2602);
DFFARX1 I_8351 (I267378,I2595,I144587,I144613,);
DFFARX1 I_8352 (I144613,I2595,I144587,I144630,);
not I_8353 (I144579,I144630);
DFFARX1 I_8354 (I267366,I2595,I144587,I144661,);
not I_8355 (I144669,I267363);
nor I_8356 (I144686,I144613,I144669);
not I_8357 (I144703,I267375);
not I_8358 (I144720,I267372);
nand I_8359 (I144737,I144720,I267375);
nor I_8360 (I144754,I144669,I144737);
nor I_8361 (I144771,I144661,I144754);
DFFARX1 I_8362 (I144720,I2595,I144587,I144576,);
nor I_8363 (I144802,I267372,I267381);
nand I_8364 (I144819,I144802,I267384);
nor I_8365 (I144836,I144819,I144703);
nand I_8366 (I144561,I144836,I267363);
DFFARX1 I_8367 (I144819,I2595,I144587,I144573,);
nand I_8368 (I144881,I144703,I267372);
nor I_8369 (I144898,I144703,I267372);
nand I_8370 (I144567,I144686,I144898);
not I_8371 (I144929,I267387);
nor I_8372 (I144946,I144929,I144881);
DFFARX1 I_8373 (I144946,I2595,I144587,I144555,);
nor I_8374 (I144977,I144929,I267390);
and I_8375 (I144994,I144977,I267369);
or I_8376 (I145011,I144994,I267363);
DFFARX1 I_8377 (I145011,I2595,I144587,I145037,);
nor I_8378 (I145045,I145037,I144661);
nor I_8379 (I144564,I144613,I145045);
not I_8380 (I145076,I145037);
nor I_8381 (I145093,I145076,I144771);
DFFARX1 I_8382 (I145093,I2595,I144587,I144570,);
nand I_8383 (I145124,I145076,I144703);
nor I_8384 (I144558,I144929,I145124);
not I_8385 (I145182,I2602);
DFFARX1 I_8386 (I33469,I2595,I145182,I145208,);
DFFARX1 I_8387 (I145208,I2595,I145182,I145225,);
not I_8388 (I145174,I145225);
DFFARX1 I_8389 (I33481,I2595,I145182,I145256,);
not I_8390 (I145264,I33472);
nor I_8391 (I145281,I145208,I145264);
not I_8392 (I145298,I33463);
not I_8393 (I145315,I33460);
nand I_8394 (I145332,I145315,I33463);
nor I_8395 (I145349,I145264,I145332);
nor I_8396 (I145366,I145256,I145349);
DFFARX1 I_8397 (I145315,I2595,I145182,I145171,);
nor I_8398 (I145397,I33460,I33460);
nand I_8399 (I145414,I145397,I33478);
nor I_8400 (I145431,I145414,I145298);
nand I_8401 (I145156,I145431,I33472);
DFFARX1 I_8402 (I145414,I2595,I145182,I145168,);
nand I_8403 (I145476,I145298,I33460);
nor I_8404 (I145493,I145298,I33460);
nand I_8405 (I145162,I145281,I145493);
not I_8406 (I145524,I33484);
nor I_8407 (I145541,I145524,I145476);
DFFARX1 I_8408 (I145541,I2595,I145182,I145150,);
nor I_8409 (I145572,I145524,I33463);
and I_8410 (I145589,I145572,I33466);
or I_8411 (I145606,I145589,I33475);
DFFARX1 I_8412 (I145606,I2595,I145182,I145632,);
nor I_8413 (I145640,I145632,I145256);
nor I_8414 (I145159,I145208,I145640);
not I_8415 (I145671,I145632);
nor I_8416 (I145688,I145671,I145366);
DFFARX1 I_8417 (I145688,I2595,I145182,I145165,);
nand I_8418 (I145719,I145671,I145298);
nor I_8419 (I145153,I145524,I145719);
not I_8420 (I145777,I2602);
DFFARX1 I_8421 (I293815,I2595,I145777,I145803,);
DFFARX1 I_8422 (I145803,I2595,I145777,I145820,);
not I_8423 (I145769,I145820);
DFFARX1 I_8424 (I293818,I2595,I145777,I145851,);
not I_8425 (I145859,I293821);
nor I_8426 (I145876,I145803,I145859);
not I_8427 (I145893,I293833);
not I_8428 (I145910,I293824);
nand I_8429 (I145927,I145910,I293833);
nor I_8430 (I145944,I145859,I145927);
nor I_8431 (I145961,I145851,I145944);
DFFARX1 I_8432 (I145910,I2595,I145777,I145766,);
nor I_8433 (I145992,I293824,I293830);
nand I_8434 (I146009,I145992,I293818);
nor I_8435 (I146026,I146009,I145893);
nand I_8436 (I145751,I146026,I293821);
DFFARX1 I_8437 (I146009,I2595,I145777,I145763,);
nand I_8438 (I146071,I145893,I293824);
nor I_8439 (I146088,I145893,I293824);
nand I_8440 (I145757,I145876,I146088);
not I_8441 (I146119,I293821);
nor I_8442 (I146136,I146119,I146071);
DFFARX1 I_8443 (I146136,I2595,I145777,I145745,);
nor I_8444 (I146167,I146119,I293827);
and I_8445 (I146184,I146167,I293815);
or I_8446 (I146201,I146184,I293836);
DFFARX1 I_8447 (I146201,I2595,I145777,I146227,);
nor I_8448 (I146235,I146227,I145851);
nor I_8449 (I145754,I145803,I146235);
not I_8450 (I146266,I146227);
nor I_8451 (I146283,I146266,I145961);
DFFARX1 I_8452 (I146283,I2595,I145777,I145760,);
nand I_8453 (I146314,I146266,I145893);
nor I_8454 (I145748,I146119,I146314);
not I_8455 (I146372,I2602);
DFFARX1 I_8456 (I383643,I2595,I146372,I146398,);
DFFARX1 I_8457 (I146398,I2595,I146372,I146415,);
not I_8458 (I146364,I146415);
DFFARX1 I_8459 (I383649,I2595,I146372,I146446,);
not I_8460 (I146454,I383664);
nor I_8461 (I146471,I146398,I146454);
not I_8462 (I146488,I383655);
not I_8463 (I146505,I383652);
nand I_8464 (I146522,I146505,I383655);
nor I_8465 (I146539,I146454,I146522);
nor I_8466 (I146556,I146446,I146539);
DFFARX1 I_8467 (I146505,I2595,I146372,I146361,);
nor I_8468 (I146587,I383652,I383643);
nand I_8469 (I146604,I146587,I383667);
nor I_8470 (I146621,I146604,I146488);
nand I_8471 (I146346,I146621,I383664);
DFFARX1 I_8472 (I146604,I2595,I146372,I146358,);
nand I_8473 (I146666,I146488,I383652);
nor I_8474 (I146683,I146488,I383652);
nand I_8475 (I146352,I146471,I146683);
not I_8476 (I146714,I383661);
nor I_8477 (I146731,I146714,I146666);
DFFARX1 I_8478 (I146731,I2595,I146372,I146340,);
nor I_8479 (I146762,I146714,I383646);
and I_8480 (I146779,I146762,I383658);
or I_8481 (I146796,I146779,I383670);
DFFARX1 I_8482 (I146796,I2595,I146372,I146822,);
nor I_8483 (I146830,I146822,I146446);
nor I_8484 (I146349,I146398,I146830);
not I_8485 (I146861,I146822);
nor I_8486 (I146878,I146861,I146556);
DFFARX1 I_8487 (I146878,I2595,I146372,I146355,);
nand I_8488 (I146909,I146861,I146488);
nor I_8489 (I146343,I146714,I146909);
not I_8490 (I146967,I2602);
DFFARX1 I_8491 (I239339,I2595,I146967,I146993,);
DFFARX1 I_8492 (I146993,I2595,I146967,I147010,);
not I_8493 (I146959,I147010);
DFFARX1 I_8494 (I239336,I2595,I146967,I147041,);
not I_8495 (I147049,I239336);
nor I_8496 (I147066,I146993,I147049);
not I_8497 (I147083,I239333);
not I_8498 (I147100,I239348);
nand I_8499 (I147117,I147100,I239333);
nor I_8500 (I147134,I147049,I147117);
nor I_8501 (I147151,I147041,I147134);
DFFARX1 I_8502 (I147100,I2595,I146967,I146956,);
nor I_8503 (I147182,I239348,I239342);
nand I_8504 (I147199,I147182,I239330);
nor I_8505 (I147216,I147199,I147083);
nand I_8506 (I146941,I147216,I239336);
DFFARX1 I_8507 (I147199,I2595,I146967,I146953,);
nand I_8508 (I147261,I147083,I239348);
nor I_8509 (I147278,I147083,I239348);
nand I_8510 (I146947,I147066,I147278);
not I_8511 (I147309,I239351);
nor I_8512 (I147326,I147309,I147261);
DFFARX1 I_8513 (I147326,I2595,I146967,I146935,);
nor I_8514 (I147357,I147309,I239330);
and I_8515 (I147374,I147357,I239345);
or I_8516 (I147391,I147374,I239333);
DFFARX1 I_8517 (I147391,I2595,I146967,I147417,);
nor I_8518 (I147425,I147417,I147041);
nor I_8519 (I146944,I146993,I147425);
not I_8520 (I147456,I147417);
nor I_8521 (I147473,I147456,I147151);
DFFARX1 I_8522 (I147473,I2595,I146967,I146950,);
nand I_8523 (I147504,I147456,I147083);
nor I_8524 (I146938,I147309,I147504);
not I_8525 (I147562,I2602);
DFFARX1 I_8526 (I248298,I2595,I147562,I147588,);
DFFARX1 I_8527 (I147588,I2595,I147562,I147605,);
not I_8528 (I147554,I147605);
DFFARX1 I_8529 (I248295,I2595,I147562,I147636,);
not I_8530 (I147644,I248295);
nor I_8531 (I147661,I147588,I147644);
not I_8532 (I147678,I248292);
not I_8533 (I147695,I248307);
nand I_8534 (I147712,I147695,I248292);
nor I_8535 (I147729,I147644,I147712);
nor I_8536 (I147746,I147636,I147729);
DFFARX1 I_8537 (I147695,I2595,I147562,I147551,);
nor I_8538 (I147777,I248307,I248301);
nand I_8539 (I147794,I147777,I248289);
nor I_8540 (I147811,I147794,I147678);
nand I_8541 (I147536,I147811,I248295);
DFFARX1 I_8542 (I147794,I2595,I147562,I147548,);
nand I_8543 (I147856,I147678,I248307);
nor I_8544 (I147873,I147678,I248307);
nand I_8545 (I147542,I147661,I147873);
not I_8546 (I147904,I248310);
nor I_8547 (I147921,I147904,I147856);
DFFARX1 I_8548 (I147921,I2595,I147562,I147530,);
nor I_8549 (I147952,I147904,I248289);
and I_8550 (I147969,I147952,I248304);
or I_8551 (I147986,I147969,I248292);
DFFARX1 I_8552 (I147986,I2595,I147562,I148012,);
nor I_8553 (I148020,I148012,I147636);
nor I_8554 (I147539,I147588,I148020);
not I_8555 (I148051,I148012);
nor I_8556 (I148068,I148051,I147746);
DFFARX1 I_8557 (I148068,I2595,I147562,I147545,);
nand I_8558 (I148099,I148051,I147678);
nor I_8559 (I147533,I147904,I148099);
not I_8560 (I148157,I2602);
DFFARX1 I_8561 (I354590,I2595,I148157,I148183,);
DFFARX1 I_8562 (I148183,I2595,I148157,I148200,);
not I_8563 (I148149,I148200);
DFFARX1 I_8564 (I354605,I2595,I148157,I148231,);
not I_8565 (I148239,I354614);
nor I_8566 (I148256,I148183,I148239);
not I_8567 (I148273,I354593);
not I_8568 (I148290,I354599);
nand I_8569 (I148307,I148290,I354593);
nor I_8570 (I148324,I148239,I148307);
nor I_8571 (I148341,I148231,I148324);
DFFARX1 I_8572 (I148290,I2595,I148157,I148146,);
nor I_8573 (I148372,I354599,I354611);
nand I_8574 (I148389,I148372,I354608);
nor I_8575 (I148406,I148389,I148273);
nand I_8576 (I148131,I148406,I354614);
DFFARX1 I_8577 (I148389,I2595,I148157,I148143,);
nand I_8578 (I148451,I148273,I354599);
nor I_8579 (I148468,I148273,I354599);
nand I_8580 (I148137,I148256,I148468);
not I_8581 (I148499,I354590);
nor I_8582 (I148516,I148499,I148451);
DFFARX1 I_8583 (I148516,I2595,I148157,I148125,);
nor I_8584 (I148547,I148499,I354602);
and I_8585 (I148564,I148547,I354596);
or I_8586 (I148581,I148564,I354593);
DFFARX1 I_8587 (I148581,I2595,I148157,I148607,);
nor I_8588 (I148615,I148607,I148231);
nor I_8589 (I148134,I148183,I148615);
not I_8590 (I148646,I148607);
nor I_8591 (I148663,I148646,I148341);
DFFARX1 I_8592 (I148663,I2595,I148157,I148140,);
nand I_8593 (I148694,I148646,I148273);
nor I_8594 (I148128,I148499,I148694);
not I_8595 (I148752,I2602);
DFFARX1 I_8596 (I265440,I2595,I148752,I148778,);
DFFARX1 I_8597 (I148778,I2595,I148752,I148795,);
not I_8598 (I148744,I148795);
DFFARX1 I_8599 (I265428,I2595,I148752,I148826,);
not I_8600 (I148834,I265425);
nor I_8601 (I148851,I148778,I148834);
not I_8602 (I148868,I265437);
not I_8603 (I148885,I265434);
nand I_8604 (I148902,I148885,I265437);
nor I_8605 (I148919,I148834,I148902);
nor I_8606 (I148936,I148826,I148919);
DFFARX1 I_8607 (I148885,I2595,I148752,I148741,);
nor I_8608 (I148967,I265434,I265443);
nand I_8609 (I148984,I148967,I265446);
nor I_8610 (I149001,I148984,I148868);
nand I_8611 (I148726,I149001,I265425);
DFFARX1 I_8612 (I148984,I2595,I148752,I148738,);
nand I_8613 (I149046,I148868,I265434);
nor I_8614 (I149063,I148868,I265434);
nand I_8615 (I148732,I148851,I149063);
not I_8616 (I149094,I265449);
nor I_8617 (I149111,I149094,I149046);
DFFARX1 I_8618 (I149111,I2595,I148752,I148720,);
nor I_8619 (I149142,I149094,I265452);
and I_8620 (I149159,I149142,I265431);
or I_8621 (I149176,I149159,I265425);
DFFARX1 I_8622 (I149176,I2595,I148752,I149202,);
nor I_8623 (I149210,I149202,I148826);
nor I_8624 (I148729,I148778,I149210);
not I_8625 (I149241,I149202);
nor I_8626 (I149258,I149241,I148936);
DFFARX1 I_8627 (I149258,I2595,I148752,I148735,);
nand I_8628 (I149289,I149241,I148868);
nor I_8629 (I148723,I149094,I149289);
not I_8630 (I149347,I2602);
DFFARX1 I_8631 (I236177,I2595,I149347,I149373,);
DFFARX1 I_8632 (I149373,I2595,I149347,I149390,);
not I_8633 (I149339,I149390);
DFFARX1 I_8634 (I236174,I2595,I149347,I149421,);
not I_8635 (I149429,I236174);
nor I_8636 (I149446,I149373,I149429);
not I_8637 (I149463,I236171);
not I_8638 (I149480,I236186);
nand I_8639 (I149497,I149480,I236171);
nor I_8640 (I149514,I149429,I149497);
nor I_8641 (I149531,I149421,I149514);
DFFARX1 I_8642 (I149480,I2595,I149347,I149336,);
nor I_8643 (I149562,I236186,I236180);
nand I_8644 (I149579,I149562,I236168);
nor I_8645 (I149596,I149579,I149463);
nand I_8646 (I149321,I149596,I236174);
DFFARX1 I_8647 (I149579,I2595,I149347,I149333,);
nand I_8648 (I149641,I149463,I236186);
nor I_8649 (I149658,I149463,I236186);
nand I_8650 (I149327,I149446,I149658);
not I_8651 (I149689,I236189);
nor I_8652 (I149706,I149689,I149641);
DFFARX1 I_8653 (I149706,I2595,I149347,I149315,);
nor I_8654 (I149737,I149689,I236168);
and I_8655 (I149754,I149737,I236183);
or I_8656 (I149771,I149754,I236171);
DFFARX1 I_8657 (I149771,I2595,I149347,I149797,);
nor I_8658 (I149805,I149797,I149421);
nor I_8659 (I149324,I149373,I149805);
not I_8660 (I149836,I149797);
nor I_8661 (I149853,I149836,I149531);
DFFARX1 I_8662 (I149853,I2595,I149347,I149330,);
nand I_8663 (I149884,I149836,I149463);
nor I_8664 (I149318,I149689,I149884);
not I_8665 (I149942,I2602);
DFFARX1 I_8666 (I340872,I2595,I149942,I149968,);
DFFARX1 I_8667 (I149968,I2595,I149942,I149985,);
not I_8668 (I149934,I149985);
DFFARX1 I_8669 (I340854,I2595,I149942,I150016,);
not I_8670 (I150024,I340860);
nor I_8671 (I150041,I149968,I150024);
not I_8672 (I150058,I340875);
not I_8673 (I150075,I340866);
nand I_8674 (I150092,I150075,I340875);
nor I_8675 (I150109,I150024,I150092);
nor I_8676 (I150126,I150016,I150109);
DFFARX1 I_8677 (I150075,I2595,I149942,I149931,);
nor I_8678 (I150157,I340866,I340878);
nand I_8679 (I150174,I150157,I340857);
nor I_8680 (I150191,I150174,I150058);
nand I_8681 (I149916,I150191,I340860);
DFFARX1 I_8682 (I150174,I2595,I149942,I149928,);
nand I_8683 (I150236,I150058,I340866);
nor I_8684 (I150253,I150058,I340866);
nand I_8685 (I149922,I150041,I150253);
not I_8686 (I150284,I340863);
nor I_8687 (I150301,I150284,I150236);
DFFARX1 I_8688 (I150301,I2595,I149942,I149910,);
nor I_8689 (I150332,I150284,I340869);
and I_8690 (I150349,I150332,I340854);
or I_8691 (I150366,I150349,I340857);
DFFARX1 I_8692 (I150366,I2595,I149942,I150392,);
nor I_8693 (I150400,I150392,I150016);
nor I_8694 (I149919,I149968,I150400);
not I_8695 (I150431,I150392);
nor I_8696 (I150448,I150431,I150126);
DFFARX1 I_8697 (I150448,I2595,I149942,I149925,);
nand I_8698 (I150479,I150431,I150058);
nor I_8699 (I149913,I150284,I150479);
not I_8700 (I150537,I2602);
DFFARX1 I_8701 (I343166,I2595,I150537,I150563,);
DFFARX1 I_8702 (I150563,I2595,I150537,I150580,);
not I_8703 (I150529,I150580);
DFFARX1 I_8704 (I343181,I2595,I150537,I150611,);
not I_8705 (I150619,I343190);
nor I_8706 (I150636,I150563,I150619);
not I_8707 (I150653,I343169);
not I_8708 (I150670,I343175);
nand I_8709 (I150687,I150670,I343169);
nor I_8710 (I150704,I150619,I150687);
nor I_8711 (I150721,I150611,I150704);
DFFARX1 I_8712 (I150670,I2595,I150537,I150526,);
nor I_8713 (I150752,I343175,I343187);
nand I_8714 (I150769,I150752,I343184);
nor I_8715 (I150786,I150769,I150653);
nand I_8716 (I150511,I150786,I343190);
DFFARX1 I_8717 (I150769,I2595,I150537,I150523,);
nand I_8718 (I150831,I150653,I343175);
nor I_8719 (I150848,I150653,I343175);
nand I_8720 (I150517,I150636,I150848);
not I_8721 (I150879,I343166);
nor I_8722 (I150896,I150879,I150831);
DFFARX1 I_8723 (I150896,I2595,I150537,I150505,);
nor I_8724 (I150927,I150879,I343178);
and I_8725 (I150944,I150927,I343172);
or I_8726 (I150961,I150944,I343169);
DFFARX1 I_8727 (I150961,I2595,I150537,I150987,);
nor I_8728 (I150995,I150987,I150611);
nor I_8729 (I150514,I150563,I150995);
not I_8730 (I151026,I150987);
nor I_8731 (I151043,I151026,I150721);
DFFARX1 I_8732 (I151043,I2595,I150537,I150520,);
nand I_8733 (I151074,I151026,I150653);
nor I_8734 (I150508,I150879,I151074);
not I_8735 (I151132,I2602);
DFFARX1 I_8736 (I196329,I2595,I151132,I151158,);
DFFARX1 I_8737 (I151158,I2595,I151132,I151175,);
not I_8738 (I151124,I151175);
DFFARX1 I_8739 (I196323,I2595,I151132,I151206,);
not I_8740 (I151214,I196320);
nor I_8741 (I151231,I151158,I151214);
not I_8742 (I151248,I196332);
not I_8743 (I151265,I196335);
nand I_8744 (I151282,I151265,I196332);
nor I_8745 (I151299,I151214,I151282);
nor I_8746 (I151316,I151206,I151299);
DFFARX1 I_8747 (I151265,I2595,I151132,I151121,);
nor I_8748 (I151347,I196335,I196344);
nand I_8749 (I151364,I151347,I196338);
nor I_8750 (I151381,I151364,I151248);
nand I_8751 (I151106,I151381,I196320);
DFFARX1 I_8752 (I151364,I2595,I151132,I151118,);
nand I_8753 (I151426,I151248,I196335);
nor I_8754 (I151443,I151248,I196335);
nand I_8755 (I151112,I151231,I151443);
not I_8756 (I151474,I196326);
nor I_8757 (I151491,I151474,I151426);
DFFARX1 I_8758 (I151491,I2595,I151132,I151100,);
nor I_8759 (I151522,I151474,I196341);
and I_8760 (I151539,I151522,I196320);
or I_8761 (I151556,I151539,I196323);
DFFARX1 I_8762 (I151556,I2595,I151132,I151582,);
nor I_8763 (I151590,I151582,I151206);
nor I_8764 (I151109,I151158,I151590);
not I_8765 (I151621,I151582);
nor I_8766 (I151638,I151621,I151316);
DFFARX1 I_8767 (I151638,I2595,I151132,I151115,);
nand I_8768 (I151669,I151621,I151248);
nor I_8769 (I151103,I151474,I151669);
not I_8770 (I151727,I2602);
DFFARX1 I_8771 (I230907,I2595,I151727,I151753,);
DFFARX1 I_8772 (I151753,I2595,I151727,I151770,);
not I_8773 (I151719,I151770);
DFFARX1 I_8774 (I230904,I2595,I151727,I151801,);
not I_8775 (I151809,I230904);
nor I_8776 (I151826,I151753,I151809);
not I_8777 (I151843,I230901);
not I_8778 (I151860,I230916);
nand I_8779 (I151877,I151860,I230901);
nor I_8780 (I151894,I151809,I151877);
nor I_8781 (I151911,I151801,I151894);
DFFARX1 I_8782 (I151860,I2595,I151727,I151716,);
nor I_8783 (I151942,I230916,I230910);
nand I_8784 (I151959,I151942,I230898);
nor I_8785 (I151976,I151959,I151843);
nand I_8786 (I151701,I151976,I230904);
DFFARX1 I_8787 (I151959,I2595,I151727,I151713,);
nand I_8788 (I152021,I151843,I230916);
nor I_8789 (I152038,I151843,I230916);
nand I_8790 (I151707,I151826,I152038);
not I_8791 (I152069,I230919);
nor I_8792 (I152086,I152069,I152021);
DFFARX1 I_8793 (I152086,I2595,I151727,I151695,);
nor I_8794 (I152117,I152069,I230898);
and I_8795 (I152134,I152117,I230913);
or I_8796 (I152151,I152134,I230901);
DFFARX1 I_8797 (I152151,I2595,I151727,I152177,);
nor I_8798 (I152185,I152177,I151801);
nor I_8799 (I151704,I151753,I152185);
not I_8800 (I152216,I152177);
nor I_8801 (I152233,I152216,I151911);
DFFARX1 I_8802 (I152233,I2595,I151727,I151710,);
nand I_8803 (I152264,I152216,I151843);
nor I_8804 (I151698,I152069,I152264);
not I_8805 (I152322,I2602);
DFFARX1 I_8806 (I175515,I2595,I152322,I152348,);
DFFARX1 I_8807 (I152348,I2595,I152322,I152365,);
not I_8808 (I152314,I152365);
DFFARX1 I_8809 (I175527,I2595,I152322,I152396,);
not I_8810 (I152404,I175512);
nor I_8811 (I152421,I152348,I152404);
not I_8812 (I152438,I175530);
not I_8813 (I152455,I175521);
nand I_8814 (I152472,I152455,I175530);
nor I_8815 (I152489,I152404,I152472);
nor I_8816 (I152506,I152396,I152489);
DFFARX1 I_8817 (I152455,I2595,I152322,I152311,);
nor I_8818 (I152537,I175521,I175533);
nand I_8819 (I152554,I152537,I175536);
nor I_8820 (I152571,I152554,I152438);
nand I_8821 (I152296,I152571,I175512);
DFFARX1 I_8822 (I152554,I2595,I152322,I152308,);
nand I_8823 (I152616,I152438,I175521);
nor I_8824 (I152633,I152438,I175521);
nand I_8825 (I152302,I152421,I152633);
not I_8826 (I152664,I175512);
nor I_8827 (I152681,I152664,I152616);
DFFARX1 I_8828 (I152681,I2595,I152322,I152290,);
nor I_8829 (I152712,I152664,I175524);
and I_8830 (I152729,I152712,I175518);
or I_8831 (I152746,I152729,I175515);
DFFARX1 I_8832 (I152746,I2595,I152322,I152772,);
nor I_8833 (I152780,I152772,I152396);
nor I_8834 (I152299,I152348,I152780);
not I_8835 (I152811,I152772);
nor I_8836 (I152828,I152811,I152506);
DFFARX1 I_8837 (I152828,I2595,I152322,I152305,);
nand I_8838 (I152859,I152811,I152438);
nor I_8839 (I152293,I152664,I152859);
not I_8840 (I152917,I2602);
DFFARX1 I_8841 (I39266,I2595,I152917,I152943,);
DFFARX1 I_8842 (I152943,I2595,I152917,I152960,);
not I_8843 (I152909,I152960);
DFFARX1 I_8844 (I39278,I2595,I152917,I152991,);
not I_8845 (I152999,I39269);
nor I_8846 (I153016,I152943,I152999);
not I_8847 (I153033,I39260);
not I_8848 (I153050,I39257);
nand I_8849 (I153067,I153050,I39260);
nor I_8850 (I153084,I152999,I153067);
nor I_8851 (I153101,I152991,I153084);
DFFARX1 I_8852 (I153050,I2595,I152917,I152906,);
nor I_8853 (I153132,I39257,I39257);
nand I_8854 (I153149,I153132,I39275);
nor I_8855 (I153166,I153149,I153033);
nand I_8856 (I152891,I153166,I39269);
DFFARX1 I_8857 (I153149,I2595,I152917,I152903,);
nand I_8858 (I153211,I153033,I39257);
nor I_8859 (I153228,I153033,I39257);
nand I_8860 (I152897,I153016,I153228);
not I_8861 (I153259,I39281);
nor I_8862 (I153276,I153259,I153211);
DFFARX1 I_8863 (I153276,I2595,I152917,I152885,);
nor I_8864 (I153307,I153259,I39260);
and I_8865 (I153324,I153307,I39263);
or I_8866 (I153341,I153324,I39272);
DFFARX1 I_8867 (I153341,I2595,I152917,I153367,);
nor I_8868 (I153375,I153367,I152991);
nor I_8869 (I152894,I152943,I153375);
not I_8870 (I153406,I153367);
nor I_8871 (I153423,I153406,I153101);
DFFARX1 I_8872 (I153423,I2595,I152917,I152900,);
nand I_8873 (I153454,I153406,I153033);
nor I_8874 (I152888,I153259,I153454);
not I_8875 (I153512,I2602);
DFFARX1 I_8876 (I389593,I2595,I153512,I153538,);
DFFARX1 I_8877 (I153538,I2595,I153512,I153555,);
not I_8878 (I153504,I153555);
DFFARX1 I_8879 (I389599,I2595,I153512,I153586,);
not I_8880 (I153594,I389614);
nor I_8881 (I153611,I153538,I153594);
not I_8882 (I153628,I389605);
not I_8883 (I153645,I389602);
nand I_8884 (I153662,I153645,I389605);
nor I_8885 (I153679,I153594,I153662);
nor I_8886 (I153696,I153586,I153679);
DFFARX1 I_8887 (I153645,I2595,I153512,I153501,);
nor I_8888 (I153727,I389602,I389593);
nand I_8889 (I153744,I153727,I389617);
nor I_8890 (I153761,I153744,I153628);
nand I_8891 (I153486,I153761,I389614);
DFFARX1 I_8892 (I153744,I2595,I153512,I153498,);
nand I_8893 (I153806,I153628,I389602);
nor I_8894 (I153823,I153628,I389602);
nand I_8895 (I153492,I153611,I153823);
not I_8896 (I153854,I389611);
nor I_8897 (I153871,I153854,I153806);
DFFARX1 I_8898 (I153871,I2595,I153512,I153480,);
nor I_8899 (I153902,I153854,I389596);
and I_8900 (I153919,I153902,I389608);
or I_8901 (I153936,I153919,I389620);
DFFARX1 I_8902 (I153936,I2595,I153512,I153962,);
nor I_8903 (I153970,I153962,I153586);
nor I_8904 (I153489,I153538,I153970);
not I_8905 (I154001,I153962);
nor I_8906 (I154018,I154001,I153696);
DFFARX1 I_8907 (I154018,I2595,I153512,I153495,);
nand I_8908 (I154049,I154001,I153628);
nor I_8909 (I153483,I153854,I154049);
not I_8910 (I154107,I2602);
DFFARX1 I_8911 (I52058,I2595,I154107,I154133,);
DFFARX1 I_8912 (I154133,I2595,I154107,I154150,);
not I_8913 (I154099,I154150);
DFFARX1 I_8914 (I52082,I2595,I154107,I154181,);
not I_8915 (I154189,I52076);
nor I_8916 (I154206,I154133,I154189);
not I_8917 (I154223,I52070);
not I_8918 (I154240,I52067);
nand I_8919 (I154257,I154240,I52070);
nor I_8920 (I154274,I154189,I154257);
nor I_8921 (I154291,I154181,I154274);
DFFARX1 I_8922 (I154240,I2595,I154107,I154096,);
nor I_8923 (I154322,I52067,I52061);
nand I_8924 (I154339,I154322,I52079);
nor I_8925 (I154356,I154339,I154223);
nand I_8926 (I154081,I154356,I52076);
DFFARX1 I_8927 (I154339,I2595,I154107,I154093,);
nand I_8928 (I154401,I154223,I52067);
nor I_8929 (I154418,I154223,I52067);
nand I_8930 (I154087,I154206,I154418);
not I_8931 (I154449,I52073);
nor I_8932 (I154466,I154449,I154401);
DFFARX1 I_8933 (I154466,I2595,I154107,I154075,);
nor I_8934 (I154497,I154449,I52058);
and I_8935 (I154514,I154497,I52064);
or I_8936 (I154531,I154514,I52061);
DFFARX1 I_8937 (I154531,I2595,I154107,I154557,);
nor I_8938 (I154565,I154557,I154181);
nor I_8939 (I154084,I154133,I154565);
not I_8940 (I154596,I154557);
nor I_8941 (I154613,I154596,I154291);
DFFARX1 I_8942 (I154613,I2595,I154107,I154090,);
nand I_8943 (I154644,I154596,I154223);
nor I_8944 (I154078,I154449,I154644);
not I_8945 (I154702,I2602);
DFFARX1 I_8946 (I92227,I2595,I154702,I154728,);
DFFARX1 I_8947 (I154728,I2595,I154702,I154745,);
not I_8948 (I154694,I154745);
DFFARX1 I_8949 (I92215,I2595,I154702,I154776,);
not I_8950 (I154784,I92218);
nor I_8951 (I154801,I154728,I154784);
not I_8952 (I154818,I92221);
not I_8953 (I154835,I92233);
nand I_8954 (I154852,I154835,I92221);
nor I_8955 (I154869,I154784,I154852);
nor I_8956 (I154886,I154776,I154869);
DFFARX1 I_8957 (I154835,I2595,I154702,I154691,);
nor I_8958 (I154917,I92233,I92224);
nand I_8959 (I154934,I154917,I92212);
nor I_8960 (I154951,I154934,I154818);
nand I_8961 (I154676,I154951,I92218);
DFFARX1 I_8962 (I154934,I2595,I154702,I154688,);
nand I_8963 (I154996,I154818,I92233);
nor I_8964 (I155013,I154818,I92233);
nand I_8965 (I154682,I154801,I155013);
not I_8966 (I155044,I92230);
nor I_8967 (I155061,I155044,I154996);
DFFARX1 I_8968 (I155061,I2595,I154702,I154670,);
nor I_8969 (I155092,I155044,I92236);
and I_8970 (I155109,I155092,I92239);
or I_8971 (I155126,I155109,I92212);
DFFARX1 I_8972 (I155126,I2595,I154702,I155152,);
nor I_8973 (I155160,I155152,I154776);
nor I_8974 (I154679,I154728,I155160);
not I_8975 (I155191,I155152);
nor I_8976 (I155208,I155191,I154886);
DFFARX1 I_8977 (I155208,I2595,I154702,I154685,);
nand I_8978 (I155239,I155191,I154818);
nor I_8979 (I154673,I155044,I155239);
not I_8980 (I155297,I2602);
DFFARX1 I_8981 (I217137,I2595,I155297,I155323,);
DFFARX1 I_8982 (I155323,I2595,I155297,I155340,);
not I_8983 (I155289,I155340);
DFFARX1 I_8984 (I217131,I2595,I155297,I155371,);
not I_8985 (I155379,I217128);
nor I_8986 (I155396,I155323,I155379);
not I_8987 (I155413,I217140);
not I_8988 (I155430,I217143);
nand I_8989 (I155447,I155430,I217140);
nor I_8990 (I155464,I155379,I155447);
nor I_8991 (I155481,I155371,I155464);
DFFARX1 I_8992 (I155430,I2595,I155297,I155286,);
nor I_8993 (I155512,I217143,I217152);
nand I_8994 (I155529,I155512,I217146);
nor I_8995 (I155546,I155529,I155413);
nand I_8996 (I155271,I155546,I217128);
DFFARX1 I_8997 (I155529,I2595,I155297,I155283,);
nand I_8998 (I155591,I155413,I217143);
nor I_8999 (I155608,I155413,I217143);
nand I_9000 (I155277,I155396,I155608);
not I_9001 (I155639,I217134);
nor I_9002 (I155656,I155639,I155591);
DFFARX1 I_9003 (I155656,I2595,I155297,I155265,);
nor I_9004 (I155687,I155639,I217149);
and I_9005 (I155704,I155687,I217128);
or I_9006 (I155721,I155704,I217131);
DFFARX1 I_9007 (I155721,I2595,I155297,I155747,);
nor I_9008 (I155755,I155747,I155371);
nor I_9009 (I155274,I155323,I155755);
not I_9010 (I155786,I155747);
nor I_9011 (I155803,I155786,I155481);
DFFARX1 I_9012 (I155803,I2595,I155297,I155280,);
nand I_9013 (I155834,I155786,I155413);
nor I_9014 (I155268,I155639,I155834);
not I_9015 (I155892,I2602);
DFFARX1 I_9016 (I336230,I2595,I155892,I155918,);
not I_9017 (I155926,I155918);
DFFARX1 I_9018 (I336236,I2595,I155892,I155952,);
not I_9019 (I155960,I336230);
nand I_9020 (I155977,I155960,I336233);
not I_9021 (I155994,I155977);
nor I_9022 (I156011,I155994,I336251);
nor I_9023 (I156028,I155926,I156011);
DFFARX1 I_9024 (I156028,I2595,I155892,I155878,);
not I_9025 (I156059,I336251);
nand I_9026 (I156076,I156059,I155994);
and I_9027 (I156093,I156059,I336254);
nand I_9028 (I156110,I156093,I336233);
nor I_9029 (I155875,I156110,I156059);
and I_9030 (I155866,I155952,I156110);
not I_9031 (I156155,I156110);
nand I_9032 (I155869,I155952,I156155);
nor I_9033 (I155863,I155918,I156110);
not I_9034 (I156200,I336239);
nor I_9035 (I156217,I156200,I336254);
nand I_9036 (I156234,I156217,I156059);
nor I_9037 (I155872,I155977,I156234);
nor I_9038 (I156265,I156200,I336245);
and I_9039 (I156282,I156265,I336242);
or I_9040 (I156299,I156282,I336248);
DFFARX1 I_9041 (I156299,I2595,I155892,I156325,);
nor I_9042 (I156333,I156325,I156076);
DFFARX1 I_9043 (I156333,I2595,I155892,I155860,);
DFFARX1 I_9044 (I156325,I2595,I155892,I155884,);
not I_9045 (I156378,I156325);
nor I_9046 (I156395,I156378,I155952);
nor I_9047 (I156412,I156217,I156395);
DFFARX1 I_9048 (I156412,I2595,I155892,I155881,);
not I_9049 (I156470,I2602);
DFFARX1 I_9050 (I351888,I2595,I156470,I156496,);
not I_9051 (I156504,I156496);
DFFARX1 I_9052 (I351882,I2595,I156470,I156530,);
not I_9053 (I156538,I351891);
nand I_9054 (I156555,I156538,I351870);
not I_9055 (I156572,I156555);
nor I_9056 (I156589,I156572,I351879);
nor I_9057 (I156606,I156504,I156589);
DFFARX1 I_9058 (I156606,I2595,I156470,I156456,);
not I_9059 (I156637,I351879);
nand I_9060 (I156654,I156637,I156572);
and I_9061 (I156671,I156637,I351894);
nand I_9062 (I156688,I156671,I351873);
nor I_9063 (I156453,I156688,I156637);
and I_9064 (I156444,I156530,I156688);
not I_9065 (I156733,I156688);
nand I_9066 (I156447,I156530,I156733);
nor I_9067 (I156441,I156496,I156688);
not I_9068 (I156778,I351876);
nor I_9069 (I156795,I156778,I351894);
nand I_9070 (I156812,I156795,I156637);
nor I_9071 (I156450,I156555,I156812);
nor I_9072 (I156843,I156778,I351885);
and I_9073 (I156860,I156843,I351873);
or I_9074 (I156877,I156860,I351870);
DFFARX1 I_9075 (I156877,I2595,I156470,I156903,);
nor I_9076 (I156911,I156903,I156654);
DFFARX1 I_9077 (I156911,I2595,I156470,I156438,);
DFFARX1 I_9078 (I156903,I2595,I156470,I156462,);
not I_9079 (I156956,I156903);
nor I_9080 (I156973,I156956,I156530);
nor I_9081 (I156990,I156795,I156973);
DFFARX1 I_9082 (I156990,I2595,I156470,I156459,);
not I_9083 (I157048,I2602);
DFFARX1 I_9084 (I143963,I2595,I157048,I157074,);
not I_9085 (I157082,I157074);
DFFARX1 I_9086 (I143975,I2595,I157048,I157108,);
not I_9087 (I157116,I143981);
nand I_9088 (I157133,I157116,I143972);
not I_9089 (I157150,I157133);
nor I_9090 (I157167,I157150,I143978);
nor I_9091 (I157184,I157082,I157167);
DFFARX1 I_9092 (I157184,I2595,I157048,I157034,);
not I_9093 (I157215,I143978);
nand I_9094 (I157232,I157215,I157150);
and I_9095 (I157249,I157215,I143969);
nand I_9096 (I157266,I157249,I143960);
nor I_9097 (I157031,I157266,I157215);
and I_9098 (I157022,I157108,I157266);
not I_9099 (I157311,I157266);
nand I_9100 (I157025,I157108,I157311);
nor I_9101 (I157019,I157074,I157266);
not I_9102 (I157356,I143966);
nor I_9103 (I157373,I157356,I143969);
nand I_9104 (I157390,I157373,I157215);
nor I_9105 (I157028,I157133,I157390);
nor I_9106 (I157421,I157356,I143963);
and I_9107 (I157438,I157421,I143960);
or I_9108 (I157455,I157438,I143984);
DFFARX1 I_9109 (I157455,I2595,I157048,I157481,);
nor I_9110 (I157489,I157481,I157232);
DFFARX1 I_9111 (I157489,I2595,I157048,I157016,);
DFFARX1 I_9112 (I157481,I2595,I157048,I157040,);
not I_9113 (I157534,I157481);
nor I_9114 (I157551,I157534,I157108);
nor I_9115 (I157568,I157373,I157551);
DFFARX1 I_9116 (I157568,I2595,I157048,I157037,);
not I_9117 (I157626,I2602);
DFFARX1 I_9118 (I391973,I2595,I157626,I157652,);
not I_9119 (I157660,I157652);
DFFARX1 I_9120 (I391973,I2595,I157626,I157686,);
not I_9121 (I157694,I391997);
nand I_9122 (I157711,I157694,I391979);
not I_9123 (I157728,I157711);
nor I_9124 (I157745,I157728,I391994);
nor I_9125 (I157762,I157660,I157745);
DFFARX1 I_9126 (I157762,I2595,I157626,I157612,);
not I_9127 (I157793,I391994);
nand I_9128 (I157810,I157793,I157728);
and I_9129 (I157827,I157793,I391976);
nand I_9130 (I157844,I157827,I391985);
nor I_9131 (I157609,I157844,I157793);
and I_9132 (I157600,I157686,I157844);
not I_9133 (I157889,I157844);
nand I_9134 (I157603,I157686,I157889);
nor I_9135 (I157597,I157652,I157844);
not I_9136 (I157934,I391982);
nor I_9137 (I157951,I157934,I391976);
nand I_9138 (I157968,I157951,I157793);
nor I_9139 (I157606,I157711,I157968);
nor I_9140 (I157999,I157934,I391991);
and I_9141 (I158016,I157999,I392000);
or I_9142 (I158033,I158016,I391988);
DFFARX1 I_9143 (I158033,I2595,I157626,I158059,);
nor I_9144 (I158067,I158059,I157810);
DFFARX1 I_9145 (I158067,I2595,I157626,I157594,);
DFFARX1 I_9146 (I158059,I2595,I157626,I157618,);
not I_9147 (I158112,I158059);
nor I_9148 (I158129,I158112,I157686);
nor I_9149 (I158146,I157951,I158129);
DFFARX1 I_9150 (I158146,I2595,I157626,I157615,);
not I_9151 (I158204,I2602);
DFFARX1 I_9152 (I17126,I2595,I158204,I158230,);
not I_9153 (I158238,I158230);
DFFARX1 I_9154 (I17129,I2595,I158204,I158264,);
not I_9155 (I158272,I17123);
nand I_9156 (I158289,I158272,I17147);
not I_9157 (I158306,I158289);
nor I_9158 (I158323,I158306,I17126);
nor I_9159 (I158340,I158238,I158323);
DFFARX1 I_9160 (I158340,I2595,I158204,I158190,);
not I_9161 (I158371,I17126);
nand I_9162 (I158388,I158371,I158306);
and I_9163 (I158405,I158371,I17141);
nand I_9164 (I158422,I158405,I17135);
nor I_9165 (I158187,I158422,I158371);
and I_9166 (I158178,I158264,I158422);
not I_9167 (I158467,I158422);
nand I_9168 (I158181,I158264,I158467);
nor I_9169 (I158175,I158230,I158422);
not I_9170 (I158512,I17144);
nor I_9171 (I158529,I158512,I17141);
nand I_9172 (I158546,I158529,I158371);
nor I_9173 (I158184,I158289,I158546);
nor I_9174 (I158577,I158512,I17123);
and I_9175 (I158594,I158577,I17132);
or I_9176 (I158611,I158594,I17138);
DFFARX1 I_9177 (I158611,I2595,I158204,I158637,);
nor I_9178 (I158645,I158637,I158388);
DFFARX1 I_9179 (I158645,I2595,I158204,I158172,);
DFFARX1 I_9180 (I158637,I2595,I158204,I158196,);
not I_9181 (I158690,I158637);
nor I_9182 (I158707,I158690,I158264);
nor I_9183 (I158724,I158529,I158707);
DFFARX1 I_9184 (I158724,I2595,I158204,I158193,);
not I_9185 (I158782,I2602);
DFFARX1 I_9186 (I246714,I2595,I158782,I158808,);
not I_9187 (I158816,I158808);
DFFARX1 I_9188 (I246714,I2595,I158782,I158842,);
not I_9189 (I158850,I246711);
nand I_9190 (I158867,I158850,I246726);
not I_9191 (I158884,I158867);
nor I_9192 (I158901,I158884,I246720);
nor I_9193 (I158918,I158816,I158901);
DFFARX1 I_9194 (I158918,I2595,I158782,I158768,);
not I_9195 (I158949,I246720);
nand I_9196 (I158966,I158949,I158884);
and I_9197 (I158983,I158949,I246717);
nand I_9198 (I159000,I158983,I246708);
nor I_9199 (I158765,I159000,I158949);
and I_9200 (I158756,I158842,I159000);
not I_9201 (I159045,I159000);
nand I_9202 (I158759,I158842,I159045);
nor I_9203 (I158753,I158808,I159000);
not I_9204 (I159090,I246729);
nor I_9205 (I159107,I159090,I246717);
nand I_9206 (I159124,I159107,I158949);
nor I_9207 (I158762,I158867,I159124);
nor I_9208 (I159155,I159090,I246708);
and I_9209 (I159172,I159155,I246711);
or I_9210 (I159189,I159172,I246723);
DFFARX1 I_9211 (I159189,I2595,I158782,I159215,);
nor I_9212 (I159223,I159215,I158966);
DFFARX1 I_9213 (I159223,I2595,I158782,I158750,);
DFFARX1 I_9214 (I159215,I2595,I158782,I158774,);
not I_9215 (I159268,I159215);
nor I_9216 (I159285,I159268,I158842);
nor I_9217 (I159302,I159107,I159285);
DFFARX1 I_9218 (I159302,I2595,I158782,I158771,);
not I_9219 (I159360,I2602);
DFFARX1 I_9220 (I318890,I2595,I159360,I159386,);
not I_9221 (I159394,I159386);
DFFARX1 I_9222 (I318896,I2595,I159360,I159420,);
not I_9223 (I159428,I318890);
nand I_9224 (I159445,I159428,I318893);
not I_9225 (I159462,I159445);
nor I_9226 (I159479,I159462,I318911);
nor I_9227 (I159496,I159394,I159479);
DFFARX1 I_9228 (I159496,I2595,I159360,I159346,);
not I_9229 (I159527,I318911);
nand I_9230 (I159544,I159527,I159462);
and I_9231 (I159561,I159527,I318914);
nand I_9232 (I159578,I159561,I318893);
nor I_9233 (I159343,I159578,I159527);
and I_9234 (I159334,I159420,I159578);
not I_9235 (I159623,I159578);
nand I_9236 (I159337,I159420,I159623);
nor I_9237 (I159331,I159386,I159578);
not I_9238 (I159668,I318899);
nor I_9239 (I159685,I159668,I318914);
nand I_9240 (I159702,I159685,I159527);
nor I_9241 (I159340,I159445,I159702);
nor I_9242 (I159733,I159668,I318905);
and I_9243 (I159750,I159733,I318902);
or I_9244 (I159767,I159750,I318908);
DFFARX1 I_9245 (I159767,I2595,I159360,I159793,);
nor I_9246 (I159801,I159793,I159544);
DFFARX1 I_9247 (I159801,I2595,I159360,I159328,);
DFFARX1 I_9248 (I159793,I2595,I159360,I159352,);
not I_9249 (I159846,I159793);
nor I_9250 (I159863,I159846,I159420);
nor I_9251 (I159880,I159685,I159863);
DFFARX1 I_9252 (I159880,I2595,I159360,I159349,);
not I_9253 (I159938,I2602);
DFFARX1 I_9254 (I372338,I2595,I159938,I159964,);
not I_9255 (I159972,I159964);
DFFARX1 I_9256 (I372338,I2595,I159938,I159998,);
not I_9257 (I160006,I372362);
nand I_9258 (I160023,I160006,I372344);
not I_9259 (I160040,I160023);
nor I_9260 (I160057,I160040,I372359);
nor I_9261 (I160074,I159972,I160057);
DFFARX1 I_9262 (I160074,I2595,I159938,I159924,);
not I_9263 (I160105,I372359);
nand I_9264 (I160122,I160105,I160040);
and I_9265 (I160139,I160105,I372341);
nand I_9266 (I160156,I160139,I372350);
nor I_9267 (I159921,I160156,I160105);
and I_9268 (I159912,I159998,I160156);
not I_9269 (I160201,I160156);
nand I_9270 (I159915,I159998,I160201);
nor I_9271 (I159909,I159964,I160156);
not I_9272 (I160246,I372347);
nor I_9273 (I160263,I160246,I372341);
nand I_9274 (I160280,I160263,I160105);
nor I_9275 (I159918,I160023,I160280);
nor I_9276 (I160311,I160246,I372356);
and I_9277 (I160328,I160311,I372365);
or I_9278 (I160345,I160328,I372353);
DFFARX1 I_9279 (I160345,I2595,I159938,I160371,);
nor I_9280 (I160379,I160371,I160122);
DFFARX1 I_9281 (I160379,I2595,I159938,I159906,);
DFFARX1 I_9282 (I160371,I2595,I159938,I159930,);
not I_9283 (I160424,I160371);
nor I_9284 (I160441,I160424,I159998);
nor I_9285 (I160458,I160263,I160441);
DFFARX1 I_9286 (I160458,I2595,I159938,I159927,);
not I_9287 (I160516,I2602);
DFFARX1 I_9288 (I104339,I2595,I160516,I160542,);
not I_9289 (I160550,I160542);
DFFARX1 I_9290 (I104354,I2595,I160516,I160576,);
not I_9291 (I160584,I104357);
nand I_9292 (I160601,I160584,I104336);
not I_9293 (I160618,I160601);
nor I_9294 (I160635,I160618,I104360);
nor I_9295 (I160652,I160550,I160635);
DFFARX1 I_9296 (I160652,I2595,I160516,I160502,);
not I_9297 (I160683,I104360);
nand I_9298 (I160700,I160683,I160618);
and I_9299 (I160717,I160683,I104342);
nand I_9300 (I160734,I160717,I104333);
nor I_9301 (I160499,I160734,I160683);
and I_9302 (I160490,I160576,I160734);
not I_9303 (I160779,I160734);
nand I_9304 (I160493,I160576,I160779);
nor I_9305 (I160487,I160542,I160734);
not I_9306 (I160824,I104333);
nor I_9307 (I160841,I160824,I104342);
nand I_9308 (I160858,I160841,I160683);
nor I_9309 (I160496,I160601,I160858);
nor I_9310 (I160889,I160824,I104348);
and I_9311 (I160906,I160889,I104351);
or I_9312 (I160923,I160906,I104345);
DFFARX1 I_9313 (I160923,I2595,I160516,I160949,);
nor I_9314 (I160957,I160949,I160700);
DFFARX1 I_9315 (I160957,I2595,I160516,I160484,);
DFFARX1 I_9316 (I160949,I2595,I160516,I160508,);
not I_9317 (I161002,I160949);
nor I_9318 (I161019,I161002,I160576);
nor I_9319 (I161036,I160841,I161019);
DFFARX1 I_9320 (I161036,I2595,I160516,I160505,);
not I_9321 (I161094,I2602);
DFFARX1 I_9322 (I187650,I2595,I161094,I161120,);
not I_9323 (I161128,I161120);
DFFARX1 I_9324 (I187662,I2595,I161094,I161154,);
not I_9325 (I161162,I187653);
nand I_9326 (I161179,I161162,I187656);
not I_9327 (I161196,I161179);
nor I_9328 (I161213,I161196,I187659);
nor I_9329 (I161230,I161128,I161213);
DFFARX1 I_9330 (I161230,I2595,I161094,I161080,);
not I_9331 (I161261,I187659);
nand I_9332 (I161278,I161261,I161196);
and I_9333 (I161295,I161261,I187653);
nand I_9334 (I161312,I161295,I187665);
nor I_9335 (I161077,I161312,I161261);
and I_9336 (I161068,I161154,I161312);
not I_9337 (I161357,I161312);
nand I_9338 (I161071,I161154,I161357);
nor I_9339 (I161065,I161120,I161312);
not I_9340 (I161402,I187671);
nor I_9341 (I161419,I161402,I187653);
nand I_9342 (I161436,I161419,I161261);
nor I_9343 (I161074,I161179,I161436);
nor I_9344 (I161467,I161402,I187650);
and I_9345 (I161484,I161467,I187668);
or I_9346 (I161501,I161484,I187674);
DFFARX1 I_9347 (I161501,I2595,I161094,I161527,);
nor I_9348 (I161535,I161527,I161278);
DFFARX1 I_9349 (I161535,I2595,I161094,I161062,);
DFFARX1 I_9350 (I161527,I2595,I161094,I161086,);
not I_9351 (I161580,I161527);
nor I_9352 (I161597,I161580,I161154);
nor I_9353 (I161614,I161419,I161597);
DFFARX1 I_9354 (I161614,I2595,I161094,I161083,);
not I_9355 (I161672,I2602);
DFFARX1 I_9356 (I384238,I2595,I161672,I161698,);
not I_9357 (I161706,I161698);
DFFARX1 I_9358 (I384238,I2595,I161672,I161732,);
not I_9359 (I161740,I384262);
nand I_9360 (I161757,I161740,I384244);
not I_9361 (I161774,I161757);
nor I_9362 (I161791,I161774,I384259);
nor I_9363 (I161808,I161706,I161791);
DFFARX1 I_9364 (I161808,I2595,I161672,I161658,);
not I_9365 (I161839,I384259);
nand I_9366 (I161856,I161839,I161774);
and I_9367 (I161873,I161839,I384241);
nand I_9368 (I161890,I161873,I384250);
nor I_9369 (I161655,I161890,I161839);
and I_9370 (I161646,I161732,I161890);
not I_9371 (I161935,I161890);
nand I_9372 (I161649,I161732,I161935);
nor I_9373 (I161643,I161698,I161890);
not I_9374 (I161980,I384247);
nor I_9375 (I161997,I161980,I384241);
nand I_9376 (I162014,I161997,I161839);
nor I_9377 (I161652,I161757,I162014);
nor I_9378 (I162045,I161980,I384256);
and I_9379 (I162062,I162045,I384265);
or I_9380 (I162079,I162062,I384253);
DFFARX1 I_9381 (I162079,I2595,I161672,I162105,);
nor I_9382 (I162113,I162105,I161856);
DFFARX1 I_9383 (I162113,I2595,I161672,I161640,);
DFFARX1 I_9384 (I162105,I2595,I161672,I161664,);
not I_9385 (I162158,I162105);
nor I_9386 (I162175,I162158,I161732);
nor I_9387 (I162192,I161997,I162175);
DFFARX1 I_9388 (I162192,I2595,I161672,I161661,);
not I_9389 (I162250,I2602);
DFFARX1 I_9390 (I68138,I2595,I162250,I162276,);
not I_9391 (I162284,I162276);
DFFARX1 I_9392 (I68123,I2595,I162250,I162310,);
not I_9393 (I162318,I68141);
nand I_9394 (I162335,I162318,I68126);
not I_9395 (I162352,I162335);
nor I_9396 (I162369,I162352,I68123);
nor I_9397 (I162386,I162284,I162369);
DFFARX1 I_9398 (I162386,I2595,I162250,I162236,);
not I_9399 (I162417,I68123);
nand I_9400 (I162434,I162417,I162352);
and I_9401 (I162451,I162417,I68126);
nand I_9402 (I162468,I162451,I68147);
nor I_9403 (I162233,I162468,I162417);
and I_9404 (I162224,I162310,I162468);
not I_9405 (I162513,I162468);
nand I_9406 (I162227,I162310,I162513);
nor I_9407 (I162221,I162276,I162468);
not I_9408 (I162558,I68135);
nor I_9409 (I162575,I162558,I68126);
nand I_9410 (I162592,I162575,I162417);
nor I_9411 (I162230,I162335,I162592);
nor I_9412 (I162623,I162558,I68129);
and I_9413 (I162640,I162623,I68144);
or I_9414 (I162657,I162640,I68132);
DFFARX1 I_9415 (I162657,I2595,I162250,I162683,);
nor I_9416 (I162691,I162683,I162434);
DFFARX1 I_9417 (I162691,I2595,I162250,I162218,);
DFFARX1 I_9418 (I162683,I2595,I162250,I162242,);
not I_9419 (I162736,I162683);
nor I_9420 (I162753,I162736,I162310);
nor I_9421 (I162770,I162575,I162753);
DFFARX1 I_9422 (I162770,I2595,I162250,I162239,);
not I_9423 (I162828,I2602);
DFFARX1 I_9424 (I379478,I2595,I162828,I162854,);
not I_9425 (I162862,I162854);
DFFARX1 I_9426 (I379478,I2595,I162828,I162888,);
not I_9427 (I162896,I379502);
nand I_9428 (I162913,I162896,I379484);
not I_9429 (I162930,I162913);
nor I_9430 (I162947,I162930,I379499);
nor I_9431 (I162964,I162862,I162947);
DFFARX1 I_9432 (I162964,I2595,I162828,I162814,);
not I_9433 (I162995,I379499);
nand I_9434 (I163012,I162995,I162930);
and I_9435 (I163029,I162995,I379481);
nand I_9436 (I163046,I163029,I379490);
nor I_9437 (I162811,I163046,I162995);
and I_9438 (I162802,I162888,I163046);
not I_9439 (I163091,I163046);
nand I_9440 (I162805,I162888,I163091);
nor I_9441 (I162799,I162854,I163046);
not I_9442 (I163136,I379487);
nor I_9443 (I163153,I163136,I379481);
nand I_9444 (I163170,I163153,I162995);
nor I_9445 (I162808,I162913,I163170);
nor I_9446 (I163201,I163136,I379496);
and I_9447 (I163218,I163201,I379505);
or I_9448 (I163235,I163218,I379493);
DFFARX1 I_9449 (I163235,I2595,I162828,I163261,);
nor I_9450 (I163269,I163261,I163012);
DFFARX1 I_9451 (I163269,I2595,I162828,I162796,);
DFFARX1 I_9452 (I163261,I2595,I162828,I162820,);
not I_9453 (I163314,I163261);
nor I_9454 (I163331,I163314,I162888);
nor I_9455 (I163348,I163153,I163331);
DFFARX1 I_9456 (I163348,I2595,I162828,I162817,);
not I_9457 (I163406,I2602);
DFFARX1 I_9458 (I118693,I2595,I163406,I163432,);
not I_9459 (I163440,I163432);
DFFARX1 I_9460 (I118705,I2595,I163406,I163466,);
not I_9461 (I163474,I118681);
nand I_9462 (I163491,I163474,I118708);
not I_9463 (I163508,I163491);
nor I_9464 (I163525,I163508,I118696);
nor I_9465 (I163542,I163440,I163525);
DFFARX1 I_9466 (I163542,I2595,I163406,I163392,);
not I_9467 (I163573,I118696);
nand I_9468 (I163590,I163573,I163508);
and I_9469 (I163607,I163573,I118681);
nand I_9470 (I163624,I163607,I118684);
nor I_9471 (I163389,I163624,I163573);
and I_9472 (I163380,I163466,I163624);
not I_9473 (I163669,I163624);
nand I_9474 (I163383,I163466,I163669);
nor I_9475 (I163377,I163432,I163624);
not I_9476 (I163714,I118690);
nor I_9477 (I163731,I163714,I118681);
nand I_9478 (I163748,I163731,I163573);
nor I_9479 (I163386,I163491,I163748);
nor I_9480 (I163779,I163714,I118699);
and I_9481 (I163796,I163779,I118687);
or I_9482 (I163813,I163796,I118702);
DFFARX1 I_9483 (I163813,I2595,I163406,I163839,);
nor I_9484 (I163847,I163839,I163590);
DFFARX1 I_9485 (I163847,I2595,I163406,I163374,);
DFFARX1 I_9486 (I163839,I2595,I163406,I163398,);
not I_9487 (I163892,I163839);
nor I_9488 (I163909,I163892,I163466);
nor I_9489 (I163926,I163731,I163909);
DFFARX1 I_9490 (I163926,I2595,I163406,I163395,);
not I_9491 (I163984,I2602);
DFFARX1 I_9492 (I91164,I2595,I163984,I164010,);
not I_9493 (I164018,I164010);
DFFARX1 I_9494 (I91179,I2595,I163984,I164044,);
not I_9495 (I164052,I91182);
nand I_9496 (I164069,I164052,I91161);
not I_9497 (I164086,I164069);
nor I_9498 (I164103,I164086,I91185);
nor I_9499 (I164120,I164018,I164103);
DFFARX1 I_9500 (I164120,I2595,I163984,I163970,);
not I_9501 (I164151,I91185);
nand I_9502 (I164168,I164151,I164086);
and I_9503 (I164185,I164151,I91167);
nand I_9504 (I164202,I164185,I91158);
nor I_9505 (I163967,I164202,I164151);
and I_9506 (I163958,I164044,I164202);
not I_9507 (I164247,I164202);
nand I_9508 (I163961,I164044,I164247);
nor I_9509 (I163955,I164010,I164202);
not I_9510 (I164292,I91158);
nor I_9511 (I164309,I164292,I91167);
nand I_9512 (I164326,I164309,I164151);
nor I_9513 (I163964,I164069,I164326);
nor I_9514 (I164357,I164292,I91173);
and I_9515 (I164374,I164357,I91176);
or I_9516 (I164391,I164374,I91170);
DFFARX1 I_9517 (I164391,I2595,I163984,I164417,);
nor I_9518 (I164425,I164417,I164168);
DFFARX1 I_9519 (I164425,I2595,I163984,I163952,);
DFFARX1 I_9520 (I164417,I2595,I163984,I163976,);
not I_9521 (I164470,I164417);
nor I_9522 (I164487,I164470,I164044);
nor I_9523 (I164504,I164309,I164487);
DFFARX1 I_9524 (I164504,I2595,I163984,I163973,);
not I_9525 (I164562,I2602);
DFFARX1 I_9526 (I80624,I2595,I164562,I164588,);
not I_9527 (I164596,I164588);
DFFARX1 I_9528 (I80639,I2595,I164562,I164622,);
not I_9529 (I164630,I80642);
nand I_9530 (I164647,I164630,I80621);
not I_9531 (I164664,I164647);
nor I_9532 (I164681,I164664,I80645);
nor I_9533 (I164698,I164596,I164681);
DFFARX1 I_9534 (I164698,I2595,I164562,I164548,);
not I_9535 (I164729,I80645);
nand I_9536 (I164746,I164729,I164664);
and I_9537 (I164763,I164729,I80627);
nand I_9538 (I164780,I164763,I80618);
nor I_9539 (I164545,I164780,I164729);
and I_9540 (I164536,I164622,I164780);
not I_9541 (I164825,I164780);
nand I_9542 (I164539,I164622,I164825);
nor I_9543 (I164533,I164588,I164780);
not I_9544 (I164870,I80618);
nor I_9545 (I164887,I164870,I80627);
nand I_9546 (I164904,I164887,I164729);
nor I_9547 (I164542,I164647,I164904);
nor I_9548 (I164935,I164870,I80633);
and I_9549 (I164952,I164935,I80636);
or I_9550 (I164969,I164952,I80630);
DFFARX1 I_9551 (I164969,I2595,I164562,I164995,);
nor I_9552 (I165003,I164995,I164746);
DFFARX1 I_9553 (I165003,I2595,I164562,I164530,);
DFFARX1 I_9554 (I164995,I2595,I164562,I164554,);
not I_9555 (I165048,I164995);
nor I_9556 (I165065,I165048,I164622);
nor I_9557 (I165082,I164887,I165065);
DFFARX1 I_9558 (I165082,I2595,I164562,I164551,);
not I_9559 (I165140,I2602);
DFFARX1 I_9560 (I109082,I2595,I165140,I165166,);
not I_9561 (I165174,I165166);
DFFARX1 I_9562 (I109097,I2595,I165140,I165200,);
not I_9563 (I165208,I109100);
nand I_9564 (I165225,I165208,I109079);
not I_9565 (I165242,I165225);
nor I_9566 (I165259,I165242,I109103);
nor I_9567 (I165276,I165174,I165259);
DFFARX1 I_9568 (I165276,I2595,I165140,I165126,);
not I_9569 (I165307,I109103);
nand I_9570 (I165324,I165307,I165242);
and I_9571 (I165341,I165307,I109085);
nand I_9572 (I165358,I165341,I109076);
nor I_9573 (I165123,I165358,I165307);
and I_9574 (I165114,I165200,I165358);
not I_9575 (I165403,I165358);
nand I_9576 (I165117,I165200,I165403);
nor I_9577 (I165111,I165166,I165358);
not I_9578 (I165448,I109076);
nor I_9579 (I165465,I165448,I109085);
nand I_9580 (I165482,I165465,I165307);
nor I_9581 (I165120,I165225,I165482);
nor I_9582 (I165513,I165448,I109091);
and I_9583 (I165530,I165513,I109094);
or I_9584 (I165547,I165530,I109088);
DFFARX1 I_9585 (I165547,I2595,I165140,I165573,);
nor I_9586 (I165581,I165573,I165324);
DFFARX1 I_9587 (I165581,I2595,I165140,I165108,);
DFFARX1 I_9588 (I165573,I2595,I165140,I165132,);
not I_9589 (I165626,I165573);
nor I_9590 (I165643,I165626,I165200);
nor I_9591 (I165660,I165465,I165643);
DFFARX1 I_9592 (I165660,I2595,I165140,I165129,);
not I_9593 (I165718,I2602);
DFFARX1 I_9594 (I38227,I2595,I165718,I165744,);
not I_9595 (I165752,I165744);
DFFARX1 I_9596 (I38206,I2595,I165718,I165778,);
not I_9597 (I165786,I38203);
nand I_9598 (I165803,I165786,I38218);
not I_9599 (I165820,I165803);
nor I_9600 (I165837,I165820,I38206);
nor I_9601 (I165854,I165752,I165837);
DFFARX1 I_9602 (I165854,I2595,I165718,I165704,);
not I_9603 (I165885,I38206);
nand I_9604 (I165902,I165885,I165820);
and I_9605 (I165919,I165885,I38209);
nand I_9606 (I165936,I165919,I38224);
nor I_9607 (I165701,I165936,I165885);
and I_9608 (I165692,I165778,I165936);
not I_9609 (I165981,I165936);
nand I_9610 (I165695,I165778,I165981);
nor I_9611 (I165689,I165744,I165936);
not I_9612 (I166026,I38215);
nor I_9613 (I166043,I166026,I38209);
nand I_9614 (I166060,I166043,I165885);
nor I_9615 (I165698,I165803,I166060);
nor I_9616 (I166091,I166026,I38203);
and I_9617 (I166108,I166091,I38212);
or I_9618 (I166125,I166108,I38221);
DFFARX1 I_9619 (I166125,I2595,I165718,I166151,);
nor I_9620 (I166159,I166151,I165902);
DFFARX1 I_9621 (I166159,I2595,I165718,I165686,);
DFFARX1 I_9622 (I166151,I2595,I165718,I165710,);
not I_9623 (I166204,I166151);
nor I_9624 (I166221,I166204,I165778);
nor I_9625 (I166238,I166043,I166221);
DFFARX1 I_9626 (I166238,I2595,I165718,I165707,);
not I_9627 (I166296,I2602);
DFFARX1 I_9628 (I364870,I2595,I166296,I166322,);
not I_9629 (I166330,I166322);
DFFARX1 I_9630 (I364882,I2595,I166296,I166356,);
not I_9631 (I166364,I364873);
nand I_9632 (I166381,I166364,I364861);
not I_9633 (I166398,I166381);
nor I_9634 (I166415,I166398,I364858);
nor I_9635 (I166432,I166330,I166415);
DFFARX1 I_9636 (I166432,I2595,I166296,I166282,);
not I_9637 (I166463,I364858);
nand I_9638 (I166480,I166463,I166398);
and I_9639 (I166497,I166463,I364864);
nand I_9640 (I166514,I166497,I364861);
nor I_9641 (I166279,I166514,I166463);
and I_9642 (I166270,I166356,I166514);
not I_9643 (I166559,I166514);
nand I_9644 (I166273,I166356,I166559);
nor I_9645 (I166267,I166322,I166514);
not I_9646 (I166604,I364879);
nor I_9647 (I166621,I166604,I364864);
nand I_9648 (I166638,I166621,I166463);
nor I_9649 (I166276,I166381,I166638);
nor I_9650 (I166669,I166604,I364867);
and I_9651 (I166686,I166669,I364858);
or I_9652 (I166703,I166686,I364876);
DFFARX1 I_9653 (I166703,I2595,I166296,I166729,);
nor I_9654 (I166737,I166729,I166480);
DFFARX1 I_9655 (I166737,I2595,I166296,I166264,);
DFFARX1 I_9656 (I166729,I2595,I166296,I166288,);
not I_9657 (I166782,I166729);
nor I_9658 (I166799,I166782,I166356);
nor I_9659 (I166816,I166621,I166799);
DFFARX1 I_9660 (I166816,I2595,I166296,I166285,);
not I_9661 (I166874,I2602);
DFFARX1 I_9662 (I15018,I2595,I166874,I166900,);
not I_9663 (I166908,I166900);
DFFARX1 I_9664 (I15021,I2595,I166874,I166934,);
not I_9665 (I166942,I15015);
nand I_9666 (I166959,I166942,I15039);
not I_9667 (I166976,I166959);
nor I_9668 (I166993,I166976,I15018);
nor I_9669 (I167010,I166908,I166993);
DFFARX1 I_9670 (I167010,I2595,I166874,I166860,);
not I_9671 (I167041,I15018);
nand I_9672 (I167058,I167041,I166976);
and I_9673 (I167075,I167041,I15033);
nand I_9674 (I167092,I167075,I15027);
nor I_9675 (I166857,I167092,I167041);
and I_9676 (I166848,I166934,I167092);
not I_9677 (I167137,I167092);
nand I_9678 (I166851,I166934,I167137);
nor I_9679 (I166845,I166900,I167092);
not I_9680 (I167182,I15036);
nor I_9681 (I167199,I167182,I15033);
nand I_9682 (I167216,I167199,I167041);
nor I_9683 (I166854,I166959,I167216);
nor I_9684 (I167247,I167182,I15015);
and I_9685 (I167264,I167247,I15024);
or I_9686 (I167281,I167264,I15030);
DFFARX1 I_9687 (I167281,I2595,I166874,I167307,);
nor I_9688 (I167315,I167307,I167058);
DFFARX1 I_9689 (I167315,I2595,I166874,I166842,);
DFFARX1 I_9690 (I167307,I2595,I166874,I166866,);
not I_9691 (I167360,I167307);
nor I_9692 (I167377,I167360,I166934);
nor I_9693 (I167394,I167199,I167377);
DFFARX1 I_9694 (I167394,I2595,I166874,I166863,);
not I_9695 (I167452,I2602);
DFFARX1 I_9696 (I268015,I2595,I167452,I167478,);
not I_9697 (I167486,I167478);
DFFARX1 I_9698 (I268012,I2595,I167452,I167512,);
not I_9699 (I167520,I268009);
nand I_9700 (I167537,I167520,I268036);
not I_9701 (I167554,I167537);
nor I_9702 (I167571,I167554,I268024);
nor I_9703 (I167588,I167486,I167571);
DFFARX1 I_9704 (I167588,I2595,I167452,I167438,);
not I_9705 (I167619,I268024);
nand I_9706 (I167636,I167619,I167554);
and I_9707 (I167653,I167619,I268030);
nand I_9708 (I167670,I167653,I268021);
nor I_9709 (I167435,I167670,I167619);
and I_9710 (I167426,I167512,I167670);
not I_9711 (I167715,I167670);
nand I_9712 (I167429,I167512,I167715);
nor I_9713 (I167423,I167478,I167670);
not I_9714 (I167760,I268018);
nor I_9715 (I167777,I167760,I268030);
nand I_9716 (I167794,I167777,I167619);
nor I_9717 (I167432,I167537,I167794);
nor I_9718 (I167825,I167760,I268033);
and I_9719 (I167842,I167825,I268027);
or I_9720 (I167859,I167842,I268009);
DFFARX1 I_9721 (I167859,I2595,I167452,I167885,);
nor I_9722 (I167893,I167885,I167636);
DFFARX1 I_9723 (I167893,I2595,I167452,I167420,);
DFFARX1 I_9724 (I167885,I2595,I167452,I167444,);
not I_9725 (I167938,I167885);
nor I_9726 (I167955,I167938,I167512);
nor I_9727 (I167972,I167777,I167955);
DFFARX1 I_9728 (I167972,I2595,I167452,I167441,);
not I_9729 (I168030,I2602);
DFFARX1 I_9730 (I287395,I2595,I168030,I168056,);
not I_9731 (I168064,I168056);
DFFARX1 I_9732 (I287392,I2595,I168030,I168090,);
not I_9733 (I168098,I287389);
nand I_9734 (I168115,I168098,I287416);
not I_9735 (I168132,I168115);
nor I_9736 (I168149,I168132,I287404);
nor I_9737 (I168166,I168064,I168149);
DFFARX1 I_9738 (I168166,I2595,I168030,I168016,);
not I_9739 (I168197,I287404);
nand I_9740 (I168214,I168197,I168132);
and I_9741 (I168231,I168197,I287410);
nand I_9742 (I168248,I168231,I287401);
nor I_9743 (I168013,I168248,I168197);
and I_9744 (I168004,I168090,I168248);
not I_9745 (I168293,I168248);
nand I_9746 (I168007,I168090,I168293);
nor I_9747 (I168001,I168056,I168248);
not I_9748 (I168338,I287398);
nor I_9749 (I168355,I168338,I287410);
nand I_9750 (I168372,I168355,I168197);
nor I_9751 (I168010,I168115,I168372);
nor I_9752 (I168403,I168338,I287413);
and I_9753 (I168420,I168403,I287407);
or I_9754 (I168437,I168420,I287389);
DFFARX1 I_9755 (I168437,I2595,I168030,I168463,);
nor I_9756 (I168471,I168463,I168214);
DFFARX1 I_9757 (I168471,I2595,I168030,I167998,);
DFFARX1 I_9758 (I168463,I2595,I168030,I168022,);
not I_9759 (I168516,I168463);
nor I_9760 (I168533,I168516,I168090);
nor I_9761 (I168550,I168355,I168533);
DFFARX1 I_9762 (I168550,I2595,I168030,I168019,);
not I_9763 (I168608,I2602);
DFFARX1 I_9764 (I205568,I2595,I168608,I168634,);
not I_9765 (I168642,I168634);
DFFARX1 I_9766 (I205580,I2595,I168608,I168668,);
not I_9767 (I168676,I205571);
nand I_9768 (I168693,I168676,I205574);
not I_9769 (I168710,I168693);
nor I_9770 (I168727,I168710,I205577);
nor I_9771 (I168744,I168642,I168727);
DFFARX1 I_9772 (I168744,I2595,I168608,I168594,);
not I_9773 (I168775,I205577);
nand I_9774 (I168792,I168775,I168710);
and I_9775 (I168809,I168775,I205571);
nand I_9776 (I168826,I168809,I205583);
nor I_9777 (I168591,I168826,I168775);
and I_9778 (I168582,I168668,I168826);
not I_9779 (I168871,I168826);
nand I_9780 (I168585,I168668,I168871);
nor I_9781 (I168579,I168634,I168826);
not I_9782 (I168916,I205589);
nor I_9783 (I168933,I168916,I205571);
nand I_9784 (I168950,I168933,I168775);
nor I_9785 (I168588,I168693,I168950);
nor I_9786 (I168981,I168916,I205568);
and I_9787 (I168998,I168981,I205586);
or I_9788 (I169015,I168998,I205592);
DFFARX1 I_9789 (I169015,I2595,I168608,I169041,);
nor I_9790 (I169049,I169041,I168792);
DFFARX1 I_9791 (I169049,I2595,I168608,I168576,);
DFFARX1 I_9792 (I169041,I2595,I168608,I168600,);
not I_9793 (I169094,I169041);
nor I_9794 (I169111,I169094,I168668);
nor I_9795 (I169128,I168933,I169111);
DFFARX1 I_9796 (I169128,I2595,I168608,I168597,);
not I_9797 (I169186,I2602);
DFFARX1 I_9798 (I366604,I2595,I169186,I169212,);
not I_9799 (I169220,I169212);
DFFARX1 I_9800 (I366616,I2595,I169186,I169246,);
not I_9801 (I169254,I366607);
nand I_9802 (I169271,I169254,I366595);
not I_9803 (I169288,I169271);
nor I_9804 (I169305,I169288,I366592);
nor I_9805 (I169322,I169220,I169305);
DFFARX1 I_9806 (I169322,I2595,I169186,I169172,);
not I_9807 (I169353,I366592);
nand I_9808 (I169370,I169353,I169288);
and I_9809 (I169387,I169353,I366598);
nand I_9810 (I169404,I169387,I366595);
nor I_9811 (I169169,I169404,I169353);
and I_9812 (I169160,I169246,I169404);
not I_9813 (I169449,I169404);
nand I_9814 (I169163,I169246,I169449);
nor I_9815 (I169157,I169212,I169404);
not I_9816 (I169494,I366613);
nor I_9817 (I169511,I169494,I366598);
nand I_9818 (I169528,I169511,I169353);
nor I_9819 (I169166,I169271,I169528);
nor I_9820 (I169559,I169494,I366601);
and I_9821 (I169576,I169559,I366592);
or I_9822 (I169593,I169576,I366610);
DFFARX1 I_9823 (I169593,I2595,I169186,I169619,);
nor I_9824 (I169627,I169619,I169370);
DFFARX1 I_9825 (I169627,I2595,I169186,I169154,);
DFFARX1 I_9826 (I169619,I2595,I169186,I169178,);
not I_9827 (I169672,I169619);
nor I_9828 (I169689,I169672,I169246);
nor I_9829 (I169706,I169511,I169689);
DFFARX1 I_9830 (I169706,I2595,I169186,I169175,);
not I_9831 (I169764,I2602);
DFFARX1 I_9832 (I77658,I2595,I169764,I169790,);
not I_9833 (I169798,I169790);
DFFARX1 I_9834 (I77643,I2595,I169764,I169824,);
not I_9835 (I169832,I77661);
nand I_9836 (I169849,I169832,I77646);
not I_9837 (I169866,I169849);
nor I_9838 (I169883,I169866,I77643);
nor I_9839 (I169900,I169798,I169883);
DFFARX1 I_9840 (I169900,I2595,I169764,I169750,);
not I_9841 (I169931,I77643);
nand I_9842 (I169948,I169931,I169866);
and I_9843 (I169965,I169931,I77646);
nand I_9844 (I169982,I169965,I77667);
nor I_9845 (I169747,I169982,I169931);
and I_9846 (I169738,I169824,I169982);
not I_9847 (I170027,I169982);
nand I_9848 (I169741,I169824,I170027);
nor I_9849 (I169735,I169790,I169982);
not I_9850 (I170072,I77655);
nor I_9851 (I170089,I170072,I77646);
nand I_9852 (I170106,I170089,I169931);
nor I_9853 (I169744,I169849,I170106);
nor I_9854 (I170137,I170072,I77649);
and I_9855 (I170154,I170137,I77664);
or I_9856 (I170171,I170154,I77652);
DFFARX1 I_9857 (I170171,I2595,I169764,I170197,);
nor I_9858 (I170205,I170197,I169948);
DFFARX1 I_9859 (I170205,I2595,I169764,I169732,);
DFFARX1 I_9860 (I170197,I2595,I169764,I169756,);
not I_9861 (I170250,I170197);
nor I_9862 (I170267,I170250,I169824);
nor I_9863 (I170284,I170089,I170267);
DFFARX1 I_9864 (I170284,I2595,I169764,I169753,);
not I_9865 (I170342,I2602);
DFFARX1 I_9866 (I20288,I2595,I170342,I170368,);
not I_9867 (I170376,I170368);
DFFARX1 I_9868 (I20291,I2595,I170342,I170402,);
not I_9869 (I170410,I20285);
nand I_9870 (I170427,I170410,I20309);
not I_9871 (I170444,I170427);
nor I_9872 (I170461,I170444,I20288);
nor I_9873 (I170478,I170376,I170461);
DFFARX1 I_9874 (I170478,I2595,I170342,I170328,);
not I_9875 (I170509,I20288);
nand I_9876 (I170526,I170509,I170444);
and I_9877 (I170543,I170509,I20303);
nand I_9878 (I170560,I170543,I20297);
nor I_9879 (I170325,I170560,I170509);
and I_9880 (I170316,I170402,I170560);
not I_9881 (I170605,I170560);
nand I_9882 (I170319,I170402,I170605);
nor I_9883 (I170313,I170368,I170560);
not I_9884 (I170650,I20306);
nor I_9885 (I170667,I170650,I20303);
nand I_9886 (I170684,I170667,I170509);
nor I_9887 (I170322,I170427,I170684);
nor I_9888 (I170715,I170650,I20285);
and I_9889 (I170732,I170715,I20294);
or I_9890 (I170749,I170732,I20300);
DFFARX1 I_9891 (I170749,I2595,I170342,I170775,);
nor I_9892 (I170783,I170775,I170526);
DFFARX1 I_9893 (I170783,I2595,I170342,I170310,);
DFFARX1 I_9894 (I170775,I2595,I170342,I170334,);
not I_9895 (I170828,I170775);
nor I_9896 (I170845,I170828,I170402);
nor I_9897 (I170862,I170667,I170845);
DFFARX1 I_9898 (I170862,I2595,I170342,I170331,);
not I_9899 (I170920,I2602);
DFFARX1 I_9900 (I44024,I2595,I170920,I170946,);
not I_9901 (I170954,I170946);
DFFARX1 I_9902 (I44003,I2595,I170920,I170980,);
not I_9903 (I170988,I44000);
nand I_9904 (I171005,I170988,I44015);
not I_9905 (I171022,I171005);
nor I_9906 (I171039,I171022,I44003);
nor I_9907 (I171056,I170954,I171039);
DFFARX1 I_9908 (I171056,I2595,I170920,I170906,);
not I_9909 (I171087,I44003);
nand I_9910 (I171104,I171087,I171022);
and I_9911 (I171121,I171087,I44006);
nand I_9912 (I171138,I171121,I44021);
nor I_9913 (I170903,I171138,I171087);
and I_9914 (I170894,I170980,I171138);
not I_9915 (I171183,I171138);
nand I_9916 (I170897,I170980,I171183);
nor I_9917 (I170891,I170946,I171138);
not I_9918 (I171228,I44012);
nor I_9919 (I171245,I171228,I44006);
nand I_9920 (I171262,I171245,I171087);
nor I_9921 (I170900,I171005,I171262);
nor I_9922 (I171293,I171228,I44000);
and I_9923 (I171310,I171293,I44009);
or I_9924 (I171327,I171310,I44018);
DFFARX1 I_9925 (I171327,I2595,I170920,I171353,);
nor I_9926 (I171361,I171353,I171104);
DFFARX1 I_9927 (I171361,I2595,I170920,I170888,);
DFFARX1 I_9928 (I171353,I2595,I170920,I170912,);
not I_9929 (I171406,I171353);
nor I_9930 (I171423,I171406,I170980);
nor I_9931 (I171440,I171245,I171423);
DFFARX1 I_9932 (I171440,I2595,I170920,I170909,);
not I_9933 (I171498,I2602);
DFFARX1 I_9934 (I100123,I2595,I171498,I171524,);
not I_9935 (I171532,I171524);
DFFARX1 I_9936 (I100138,I2595,I171498,I171558,);
not I_9937 (I171566,I100141);
nand I_9938 (I171583,I171566,I100120);
not I_9939 (I171600,I171583);
nor I_9940 (I171617,I171600,I100144);
nor I_9941 (I171634,I171532,I171617);
DFFARX1 I_9942 (I171634,I2595,I171498,I171484,);
not I_9943 (I171665,I100144);
nand I_9944 (I171682,I171665,I171600);
and I_9945 (I171699,I171665,I100126);
nand I_9946 (I171716,I171699,I100117);
nor I_9947 (I171481,I171716,I171665);
and I_9948 (I171472,I171558,I171716);
not I_9949 (I171761,I171716);
nand I_9950 (I171475,I171558,I171761);
nor I_9951 (I171469,I171524,I171716);
not I_9952 (I171806,I100117);
nor I_9953 (I171823,I171806,I100126);
nand I_9954 (I171840,I171823,I171665);
nor I_9955 (I171478,I171583,I171840);
nor I_9956 (I171871,I171806,I100132);
and I_9957 (I171888,I171871,I100135);
or I_9958 (I171905,I171888,I100129);
DFFARX1 I_9959 (I171905,I2595,I171498,I171931,);
nor I_9960 (I171939,I171931,I171682);
DFFARX1 I_9961 (I171939,I2595,I171498,I171466,);
DFFARX1 I_9962 (I171931,I2595,I171498,I171490,);
not I_9963 (I171984,I171931);
nor I_9964 (I172001,I171984,I171558);
nor I_9965 (I172018,I171823,I172001);
DFFARX1 I_9966 (I172018,I2595,I171498,I171487,);
not I_9967 (I172076,I2602);
DFFARX1 I_9968 (I329872,I2595,I172076,I172102,);
not I_9969 (I172110,I172102);
DFFARX1 I_9970 (I329878,I2595,I172076,I172136,);
not I_9971 (I172144,I329872);
nand I_9972 (I172161,I172144,I329875);
not I_9973 (I172178,I172161);
nor I_9974 (I172195,I172178,I329893);
nor I_9975 (I172212,I172110,I172195);
DFFARX1 I_9976 (I172212,I2595,I172076,I172062,);
not I_9977 (I172243,I329893);
nand I_9978 (I172260,I172243,I172178);
and I_9979 (I172277,I172243,I329896);
nand I_9980 (I172294,I172277,I329875);
nor I_9981 (I172059,I172294,I172243);
and I_9982 (I172050,I172136,I172294);
not I_9983 (I172339,I172294);
nand I_9984 (I172053,I172136,I172339);
nor I_9985 (I172047,I172102,I172294);
not I_9986 (I172384,I329881);
nor I_9987 (I172401,I172384,I329896);
nand I_9988 (I172418,I172401,I172243);
nor I_9989 (I172056,I172161,I172418);
nor I_9990 (I172449,I172384,I329887);
and I_9991 (I172466,I172449,I329884);
or I_9992 (I172483,I172466,I329890);
DFFARX1 I_9993 (I172483,I2595,I172076,I172509,);
nor I_9994 (I172517,I172509,I172260);
DFFARX1 I_9995 (I172517,I2595,I172076,I172044,);
DFFARX1 I_9996 (I172509,I2595,I172076,I172068,);
not I_9997 (I172562,I172509);
nor I_9998 (I172579,I172562,I172136);
nor I_9999 (I172596,I172401,I172579);
DFFARX1 I_10000 (I172596,I2595,I172076,I172065,);
not I_10001 (I172654,I2602);
DFFARX1 I_10002 (I250930,I2595,I172654,I172680,);
not I_10003 (I172688,I172680);
DFFARX1 I_10004 (I250930,I2595,I172654,I172714,);
not I_10005 (I172722,I250927);
nand I_10006 (I172739,I172722,I250942);
not I_10007 (I172756,I172739);
nor I_10008 (I172773,I172756,I250936);
nor I_10009 (I172790,I172688,I172773);
DFFARX1 I_10010 (I172790,I2595,I172654,I172640,);
not I_10011 (I172821,I250936);
nand I_10012 (I172838,I172821,I172756);
and I_10013 (I172855,I172821,I250933);
nand I_10014 (I172872,I172855,I250924);
nor I_10015 (I172637,I172872,I172821);
and I_10016 (I172628,I172714,I172872);
not I_10017 (I172917,I172872);
nand I_10018 (I172631,I172714,I172917);
nor I_10019 (I172625,I172680,I172872);
not I_10020 (I172962,I250945);
nor I_10021 (I172979,I172962,I250933);
nand I_10022 (I172996,I172979,I172821);
nor I_10023 (I172634,I172739,I172996);
nor I_10024 (I173027,I172962,I250924);
and I_10025 (I173044,I173027,I250927);
or I_10026 (I173061,I173044,I250939);
DFFARX1 I_10027 (I173061,I2595,I172654,I173087,);
nor I_10028 (I173095,I173087,I172838);
DFFARX1 I_10029 (I173095,I2595,I172654,I172622,);
DFFARX1 I_10030 (I173087,I2595,I172654,I172646,);
not I_10031 (I173140,I173087);
nor I_10032 (I173157,I173140,I172714);
nor I_10033 (I173174,I172979,I173157);
DFFARX1 I_10034 (I173174,I2595,I172654,I172643,);
not I_10035 (I173232,I2602);
DFFARX1 I_10036 (I339120,I2595,I173232,I173258,);
not I_10037 (I173266,I173258);
DFFARX1 I_10038 (I339126,I2595,I173232,I173292,);
not I_10039 (I173300,I339120);
nand I_10040 (I173317,I173300,I339123);
not I_10041 (I173334,I173317);
nor I_10042 (I173351,I173334,I339141);
nor I_10043 (I173368,I173266,I173351);
DFFARX1 I_10044 (I173368,I2595,I173232,I173218,);
not I_10045 (I173399,I339141);
nand I_10046 (I173416,I173399,I173334);
and I_10047 (I173433,I173399,I339144);
nand I_10048 (I173450,I173433,I339123);
nor I_10049 (I173215,I173450,I173399);
and I_10050 (I173206,I173292,I173450);
not I_10051 (I173495,I173450);
nand I_10052 (I173209,I173292,I173495);
nor I_10053 (I173203,I173258,I173450);
not I_10054 (I173540,I339129);
nor I_10055 (I173557,I173540,I339144);
nand I_10056 (I173574,I173557,I173399);
nor I_10057 (I173212,I173317,I173574);
nor I_10058 (I173605,I173540,I339135);
and I_10059 (I173622,I173605,I339132);
or I_10060 (I173639,I173622,I339138);
DFFARX1 I_10061 (I173639,I2595,I173232,I173665,);
nor I_10062 (I173673,I173665,I173416);
DFFARX1 I_10063 (I173673,I2595,I173232,I173200,);
DFFARX1 I_10064 (I173665,I2595,I173232,I173224,);
not I_10065 (I173718,I173665);
nor I_10066 (I173735,I173718,I173292);
nor I_10067 (I173752,I173557,I173735);
DFFARX1 I_10068 (I173752,I2595,I173232,I173221,);
not I_10069 (I173810,I2602);
DFFARX1 I_10070 (I353520,I2595,I173810,I173836,);
not I_10071 (I173844,I173836);
DFFARX1 I_10072 (I353514,I2595,I173810,I173870,);
not I_10073 (I173878,I353523);
nand I_10074 (I173895,I173878,I353502);
not I_10075 (I173912,I173895);
nor I_10076 (I173929,I173912,I353511);
nor I_10077 (I173946,I173844,I173929);
DFFARX1 I_10078 (I173946,I2595,I173810,I173796,);
not I_10079 (I173977,I353511);
nand I_10080 (I173994,I173977,I173912);
and I_10081 (I174011,I173977,I353526);
nand I_10082 (I174028,I174011,I353505);
nor I_10083 (I173793,I174028,I173977);
and I_10084 (I173784,I173870,I174028);
not I_10085 (I174073,I174028);
nand I_10086 (I173787,I173870,I174073);
nor I_10087 (I173781,I173836,I174028);
not I_10088 (I174118,I353508);
nor I_10089 (I174135,I174118,I353526);
nand I_10090 (I174152,I174135,I173977);
nor I_10091 (I173790,I173895,I174152);
nor I_10092 (I174183,I174118,I353517);
and I_10093 (I174200,I174183,I353505);
or I_10094 (I174217,I174200,I353502);
DFFARX1 I_10095 (I174217,I2595,I173810,I174243,);
nor I_10096 (I174251,I174243,I173994);
DFFARX1 I_10097 (I174251,I2595,I173810,I173778,);
DFFARX1 I_10098 (I174243,I2595,I173810,I173802,);
not I_10099 (I174296,I174243);
nor I_10100 (I174313,I174296,I173870);
nor I_10101 (I174330,I174135,I174313);
DFFARX1 I_10102 (I174330,I2595,I173810,I173799,);
not I_10103 (I174388,I2602);
DFFARX1 I_10104 (I214238,I2595,I174388,I174414,);
not I_10105 (I174422,I174414);
DFFARX1 I_10106 (I214250,I2595,I174388,I174448,);
not I_10107 (I174456,I214241);
nand I_10108 (I174473,I174456,I214244);
not I_10109 (I174490,I174473);
nor I_10110 (I174507,I174490,I214247);
nor I_10111 (I174524,I174422,I174507);
DFFARX1 I_10112 (I174524,I2595,I174388,I174374,);
not I_10113 (I174555,I214247);
nand I_10114 (I174572,I174555,I174490);
and I_10115 (I174589,I174555,I214241);
nand I_10116 (I174606,I174589,I214253);
nor I_10117 (I174371,I174606,I174555);
and I_10118 (I174362,I174448,I174606);
not I_10119 (I174651,I174606);
nand I_10120 (I174365,I174448,I174651);
nor I_10121 (I174359,I174414,I174606);
not I_10122 (I174696,I214259);
nor I_10123 (I174713,I174696,I214241);
nand I_10124 (I174730,I174713,I174555);
nor I_10125 (I174368,I174473,I174730);
nor I_10126 (I174761,I174696,I214238);
and I_10127 (I174778,I174761,I214256);
or I_10128 (I174795,I174778,I214262);
DFFARX1 I_10129 (I174795,I2595,I174388,I174821,);
nor I_10130 (I174829,I174821,I174572);
DFFARX1 I_10131 (I174829,I2595,I174388,I174356,);
DFFARX1 I_10132 (I174821,I2595,I174388,I174380,);
not I_10133 (I174874,I174821);
nor I_10134 (I174891,I174874,I174448);
nor I_10135 (I174908,I174713,I174891);
DFFARX1 I_10136 (I174908,I2595,I174388,I174377,);
not I_10137 (I174966,I2602);
DFFARX1 I_10138 (I103812,I2595,I174966,I174992,);
not I_10139 (I175000,I174992);
DFFARX1 I_10140 (I103827,I2595,I174966,I175026,);
not I_10141 (I175034,I103830);
nand I_10142 (I175051,I175034,I103809);
not I_10143 (I175068,I175051);
nor I_10144 (I175085,I175068,I103833);
nor I_10145 (I175102,I175000,I175085);
DFFARX1 I_10146 (I175102,I2595,I174966,I174952,);
not I_10147 (I175133,I103833);
nand I_10148 (I175150,I175133,I175068);
and I_10149 (I175167,I175133,I103815);
nand I_10150 (I175184,I175167,I103806);
nor I_10151 (I174949,I175184,I175133);
and I_10152 (I174940,I175026,I175184);
not I_10153 (I175229,I175184);
nand I_10154 (I174943,I175026,I175229);
nor I_10155 (I174937,I174992,I175184);
not I_10156 (I175274,I103806);
nor I_10157 (I175291,I175274,I103815);
nand I_10158 (I175308,I175291,I175133);
nor I_10159 (I174946,I175051,I175308);
nor I_10160 (I175339,I175274,I103821);
and I_10161 (I175356,I175339,I103824);
or I_10162 (I175373,I175356,I103818);
DFFARX1 I_10163 (I175373,I2595,I174966,I175399,);
nor I_10164 (I175407,I175399,I175150);
DFFARX1 I_10165 (I175407,I2595,I174966,I174934,);
DFFARX1 I_10166 (I175399,I2595,I174966,I174958,);
not I_10167 (I175452,I175399);
nor I_10168 (I175469,I175452,I175026);
nor I_10169 (I175486,I175291,I175469);
DFFARX1 I_10170 (I175486,I2595,I174966,I174955,);
not I_10171 (I175544,I2602);
DFFARX1 I_10172 (I6782,I2595,I175544,I175570,);
not I_10173 (I175578,I175570);
DFFARX1 I_10174 (I6770,I2595,I175544,I175604,);
not I_10175 (I175612,I6779);
nand I_10176 (I175629,I175612,I6776);
not I_10177 (I175646,I175629);
nor I_10178 (I175663,I175646,I6785);
nor I_10179 (I175680,I175578,I175663);
DFFARX1 I_10180 (I175680,I2595,I175544,I175530,);
not I_10181 (I175711,I6785);
nand I_10182 (I175728,I175711,I175646);
and I_10183 (I175745,I175711,I6773);
nand I_10184 (I175762,I175745,I6776);
nor I_10185 (I175527,I175762,I175711);
and I_10186 (I175518,I175604,I175762);
not I_10187 (I175807,I175762);
nand I_10188 (I175521,I175604,I175807);
nor I_10189 (I175515,I175570,I175762);
not I_10190 (I175852,I6791);
nor I_10191 (I175869,I175852,I6773);
nand I_10192 (I175886,I175869,I175711);
nor I_10193 (I175524,I175629,I175886);
nor I_10194 (I175917,I175852,I6773);
and I_10195 (I175934,I175917,I6788);
or I_10196 (I175951,I175934,I6770);
DFFARX1 I_10197 (I175951,I2595,I175544,I175977,);
nor I_10198 (I175985,I175977,I175728);
DFFARX1 I_10199 (I175985,I2595,I175544,I175512,);
DFFARX1 I_10200 (I175977,I2595,I175544,I175536,);
not I_10201 (I176030,I175977);
nor I_10202 (I176047,I176030,I175604);
nor I_10203 (I176064,I175869,I176047);
DFFARX1 I_10204 (I176064,I2595,I175544,I175533,);
not I_10205 (I176122,I2602);
DFFARX1 I_10206 (I220596,I2595,I176122,I176148,);
not I_10207 (I176156,I176148);
DFFARX1 I_10208 (I220608,I2595,I176122,I176182,);
not I_10209 (I176190,I220599);
nand I_10210 (I176207,I176190,I220602);
not I_10211 (I176224,I176207);
nor I_10212 (I176241,I176224,I220605);
nor I_10213 (I176258,I176156,I176241);
DFFARX1 I_10214 (I176258,I2595,I176122,I176108,);
not I_10215 (I176289,I220605);
nand I_10216 (I176306,I176289,I176224);
and I_10217 (I176323,I176289,I220599);
nand I_10218 (I176340,I176323,I220611);
nor I_10219 (I176105,I176340,I176289);
and I_10220 (I176096,I176182,I176340);
not I_10221 (I176385,I176340);
nand I_10222 (I176099,I176182,I176385);
nor I_10223 (I176093,I176148,I176340);
not I_10224 (I176430,I220617);
nor I_10225 (I176447,I176430,I220599);
nand I_10226 (I176464,I176447,I176289);
nor I_10227 (I176102,I176207,I176464);
nor I_10228 (I176495,I176430,I220596);
and I_10229 (I176512,I176495,I220614);
or I_10230 (I176529,I176512,I220620);
DFFARX1 I_10231 (I176529,I2595,I176122,I176555,);
nor I_10232 (I176563,I176555,I176306);
DFFARX1 I_10233 (I176563,I2595,I176122,I176090,);
DFFARX1 I_10234 (I176555,I2595,I176122,I176114,);
not I_10235 (I176608,I176555);
nor I_10236 (I176625,I176608,I176182);
nor I_10237 (I176642,I176447,I176625);
DFFARX1 I_10238 (I176642,I2595,I176122,I176111,);
not I_10239 (I176700,I2602);
DFFARX1 I_10240 (I277059,I2595,I176700,I176726,);
not I_10241 (I176734,I176726);
DFFARX1 I_10242 (I277056,I2595,I176700,I176760,);
not I_10243 (I176768,I277053);
nand I_10244 (I176785,I176768,I277080);
not I_10245 (I176802,I176785);
nor I_10246 (I176819,I176802,I277068);
nor I_10247 (I176836,I176734,I176819);
DFFARX1 I_10248 (I176836,I2595,I176700,I176686,);
not I_10249 (I176867,I277068);
nand I_10250 (I176884,I176867,I176802);
and I_10251 (I176901,I176867,I277074);
nand I_10252 (I176918,I176901,I277065);
nor I_10253 (I176683,I176918,I176867);
and I_10254 (I176674,I176760,I176918);
not I_10255 (I176963,I176918);
nand I_10256 (I176677,I176760,I176963);
nor I_10257 (I176671,I176726,I176918);
not I_10258 (I177008,I277062);
nor I_10259 (I177025,I177008,I277074);
nand I_10260 (I177042,I177025,I176867);
nor I_10261 (I176680,I176785,I177042);
nor I_10262 (I177073,I177008,I277077);
and I_10263 (I177090,I177073,I277071);
or I_10264 (I177107,I177090,I277053);
DFFARX1 I_10265 (I177107,I2595,I176700,I177133,);
nor I_10266 (I177141,I177133,I176884);
DFFARX1 I_10267 (I177141,I2595,I176700,I176668,);
DFFARX1 I_10268 (I177133,I2595,I176700,I176692,);
not I_10269 (I177186,I177133);
nor I_10270 (I177203,I177186,I176760);
nor I_10271 (I177220,I177025,I177203);
DFFARX1 I_10272 (I177220,I2595,I176700,I176689,);
not I_10273 (I177278,I2602);
DFFARX1 I_10274 (I90637,I2595,I177278,I177304,);
not I_10275 (I177312,I177304);
DFFARX1 I_10276 (I90652,I2595,I177278,I177338,);
not I_10277 (I177346,I90655);
nand I_10278 (I177363,I177346,I90634);
not I_10279 (I177380,I177363);
nor I_10280 (I177397,I177380,I90658);
nor I_10281 (I177414,I177312,I177397);
DFFARX1 I_10282 (I177414,I2595,I177278,I177264,);
not I_10283 (I177445,I90658);
nand I_10284 (I177462,I177445,I177380);
and I_10285 (I177479,I177445,I90640);
nand I_10286 (I177496,I177479,I90631);
nor I_10287 (I177261,I177496,I177445);
and I_10288 (I177252,I177338,I177496);
not I_10289 (I177541,I177496);
nand I_10290 (I177255,I177338,I177541);
nor I_10291 (I177249,I177304,I177496);
not I_10292 (I177586,I90631);
nor I_10293 (I177603,I177586,I90640);
nand I_10294 (I177620,I177603,I177445);
nor I_10295 (I177258,I177363,I177620);
nor I_10296 (I177651,I177586,I90646);
and I_10297 (I177668,I177651,I90649);
or I_10298 (I177685,I177668,I90643);
DFFARX1 I_10299 (I177685,I2595,I177278,I177711,);
nor I_10300 (I177719,I177711,I177462);
DFFARX1 I_10301 (I177719,I2595,I177278,I177246,);
DFFARX1 I_10302 (I177711,I2595,I177278,I177270,);
not I_10303 (I177764,I177711);
nor I_10304 (I177781,I177764,I177338);
nor I_10305 (I177798,I177603,I177781);
DFFARX1 I_10306 (I177798,I2595,I177278,I177267,);
not I_10307 (I177856,I2602);
DFFARX1 I_10308 (I113825,I2595,I177856,I177882,);
not I_10309 (I177890,I177882);
DFFARX1 I_10310 (I113840,I2595,I177856,I177916,);
not I_10311 (I177924,I113843);
nand I_10312 (I177941,I177924,I113822);
not I_10313 (I177958,I177941);
nor I_10314 (I177975,I177958,I113846);
nor I_10315 (I177992,I177890,I177975);
DFFARX1 I_10316 (I177992,I2595,I177856,I177842,);
not I_10317 (I178023,I113846);
nand I_10318 (I178040,I178023,I177958);
and I_10319 (I178057,I178023,I113828);
nand I_10320 (I178074,I178057,I113819);
nor I_10321 (I177839,I178074,I178023);
and I_10322 (I177830,I177916,I178074);
not I_10323 (I178119,I178074);
nand I_10324 (I177833,I177916,I178119);
nor I_10325 (I177827,I177882,I178074);
not I_10326 (I178164,I113819);
nor I_10327 (I178181,I178164,I113828);
nand I_10328 (I178198,I178181,I178023);
nor I_10329 (I177836,I177941,I178198);
nor I_10330 (I178229,I178164,I113834);
and I_10331 (I178246,I178229,I113837);
or I_10332 (I178263,I178246,I113831);
DFFARX1 I_10333 (I178263,I2595,I177856,I178289,);
nor I_10334 (I178297,I178289,I178040);
DFFARX1 I_10335 (I178297,I2595,I177856,I177824,);
DFFARX1 I_10336 (I178289,I2595,I177856,I177848,);
not I_10337 (I178342,I178289);
nor I_10338 (I178359,I178342,I177916);
nor I_10339 (I178376,I178181,I178359);
DFFARX1 I_10340 (I178376,I2595,I177856,I177845,);
not I_10341 (I178434,I2602);
DFFARX1 I_10342 (I71113,I2595,I178434,I178460,);
not I_10343 (I178468,I178460);
DFFARX1 I_10344 (I71098,I2595,I178434,I178494,);
not I_10345 (I178502,I71116);
nand I_10346 (I178519,I178502,I71101);
not I_10347 (I178536,I178519);
nor I_10348 (I178553,I178536,I71098);
nor I_10349 (I178570,I178468,I178553);
DFFARX1 I_10350 (I178570,I2595,I178434,I178420,);
not I_10351 (I178601,I71098);
nand I_10352 (I178618,I178601,I178536);
and I_10353 (I178635,I178601,I71101);
nand I_10354 (I178652,I178635,I71122);
nor I_10355 (I178417,I178652,I178601);
and I_10356 (I178408,I178494,I178652);
not I_10357 (I178697,I178652);
nand I_10358 (I178411,I178494,I178697);
nor I_10359 (I178405,I178460,I178652);
not I_10360 (I178742,I71110);
nor I_10361 (I178759,I178742,I71101);
nand I_10362 (I178776,I178759,I178601);
nor I_10363 (I178414,I178519,I178776);
nor I_10364 (I178807,I178742,I71104);
and I_10365 (I178824,I178807,I71119);
or I_10366 (I178841,I178824,I71107);
DFFARX1 I_10367 (I178841,I2595,I178434,I178867,);
nor I_10368 (I178875,I178867,I178618);
DFFARX1 I_10369 (I178875,I2595,I178434,I178402,);
DFFARX1 I_10370 (I178867,I2595,I178434,I178426,);
not I_10371 (I178920,I178867);
nor I_10372 (I178937,I178920,I178494);
nor I_10373 (I178954,I178759,I178937);
DFFARX1 I_10374 (I178954,I2595,I178434,I178423,);
not I_10375 (I179012,I2602);
DFFARX1 I_10376 (I354064,I2595,I179012,I179038,);
not I_10377 (I179046,I179038);
DFFARX1 I_10378 (I354058,I2595,I179012,I179072,);
not I_10379 (I179080,I354067);
nand I_10380 (I179097,I179080,I354046);
not I_10381 (I179114,I179097);
nor I_10382 (I179131,I179114,I354055);
nor I_10383 (I179148,I179046,I179131);
DFFARX1 I_10384 (I179148,I2595,I179012,I178998,);
not I_10385 (I179179,I354055);
nand I_10386 (I179196,I179179,I179114);
and I_10387 (I179213,I179179,I354070);
nand I_10388 (I179230,I179213,I354049);
nor I_10389 (I178995,I179230,I179179);
and I_10390 (I178986,I179072,I179230);
not I_10391 (I179275,I179230);
nand I_10392 (I178989,I179072,I179275);
nor I_10393 (I178983,I179038,I179230);
not I_10394 (I179320,I354052);
nor I_10395 (I179337,I179320,I354070);
nand I_10396 (I179354,I179337,I179179);
nor I_10397 (I178992,I179097,I179354);
nor I_10398 (I179385,I179320,I354061);
and I_10399 (I179402,I179385,I354049);
or I_10400 (I179419,I179402,I354046);
DFFARX1 I_10401 (I179419,I2595,I179012,I179445,);
nor I_10402 (I179453,I179445,I179196);
DFFARX1 I_10403 (I179453,I2595,I179012,I178980,);
DFFARX1 I_10404 (I179445,I2595,I179012,I179004,);
not I_10405 (I179498,I179445);
nor I_10406 (I179515,I179498,I179072);
nor I_10407 (I179532,I179337,I179515);
DFFARX1 I_10408 (I179532,I2595,I179012,I179001,);
not I_10409 (I179590,I2602);
DFFARX1 I_10410 (I54453,I2595,I179590,I179616,);
not I_10411 (I179624,I179616);
DFFARX1 I_10412 (I54438,I2595,I179590,I179650,);
not I_10413 (I179658,I54456);
nand I_10414 (I179675,I179658,I54441);
not I_10415 (I179692,I179675);
nor I_10416 (I179709,I179692,I54438);
nor I_10417 (I179726,I179624,I179709);
DFFARX1 I_10418 (I179726,I2595,I179590,I179576,);
not I_10419 (I179757,I54438);
nand I_10420 (I179774,I179757,I179692);
and I_10421 (I179791,I179757,I54441);
nand I_10422 (I179808,I179791,I54462);
nor I_10423 (I179573,I179808,I179757);
and I_10424 (I179564,I179650,I179808);
not I_10425 (I179853,I179808);
nand I_10426 (I179567,I179650,I179853);
nor I_10427 (I179561,I179616,I179808);
not I_10428 (I179898,I54450);
nor I_10429 (I179915,I179898,I54441);
nand I_10430 (I179932,I179915,I179757);
nor I_10431 (I179570,I179675,I179932);
nor I_10432 (I179963,I179898,I54444);
and I_10433 (I179980,I179963,I54459);
or I_10434 (I179997,I179980,I54447);
DFFARX1 I_10435 (I179997,I2595,I179590,I180023,);
nor I_10436 (I180031,I180023,I179774);
DFFARX1 I_10437 (I180031,I2595,I179590,I179558,);
DFFARX1 I_10438 (I180023,I2595,I179590,I179582,);
not I_10439 (I180076,I180023);
nor I_10440 (I180093,I180076,I179650);
nor I_10441 (I180110,I179915,I180093);
DFFARX1 I_10442 (I180110,I2595,I179590,I179579,);
not I_10443 (I180168,I2602);
DFFARX1 I_10444 (I241444,I2595,I180168,I180194,);
not I_10445 (I180202,I180194);
DFFARX1 I_10446 (I241444,I2595,I180168,I180228,);
not I_10447 (I180236,I241441);
nand I_10448 (I180253,I180236,I241456);
not I_10449 (I180270,I180253);
nor I_10450 (I180287,I180270,I241450);
nor I_10451 (I180304,I180202,I180287);
DFFARX1 I_10452 (I180304,I2595,I180168,I180154,);
not I_10453 (I180335,I241450);
nand I_10454 (I180352,I180335,I180270);
and I_10455 (I180369,I180335,I241447);
nand I_10456 (I180386,I180369,I241438);
nor I_10457 (I180151,I180386,I180335);
and I_10458 (I180142,I180228,I180386);
not I_10459 (I180431,I180386);
nand I_10460 (I180145,I180228,I180431);
nor I_10461 (I180139,I180194,I180386);
not I_10462 (I180476,I241459);
nor I_10463 (I180493,I180476,I241447);
nand I_10464 (I180510,I180493,I180335);
nor I_10465 (I180148,I180253,I180510);
nor I_10466 (I180541,I180476,I241438);
and I_10467 (I180558,I180541,I241441);
or I_10468 (I180575,I180558,I241453);
DFFARX1 I_10469 (I180575,I2595,I180168,I180601,);
nor I_10470 (I180609,I180601,I180352);
DFFARX1 I_10471 (I180609,I2595,I180168,I180136,);
DFFARX1 I_10472 (I180601,I2595,I180168,I180160,);
not I_10473 (I180654,I180601);
nor I_10474 (I180671,I180654,I180228);
nor I_10475 (I180688,I180493,I180671);
DFFARX1 I_10476 (I180688,I2595,I180168,I180157,);
not I_10477 (I180746,I2602);
DFFARX1 I_10478 (I55643,I2595,I180746,I180772,);
not I_10479 (I180780,I180772);
DFFARX1 I_10480 (I55628,I2595,I180746,I180806,);
not I_10481 (I180814,I55646);
nand I_10482 (I180831,I180814,I55631);
not I_10483 (I180848,I180831);
nor I_10484 (I180865,I180848,I55628);
nor I_10485 (I180882,I180780,I180865);
DFFARX1 I_10486 (I180882,I2595,I180746,I180732,);
not I_10487 (I180913,I55628);
nand I_10488 (I180930,I180913,I180848);
and I_10489 (I180947,I180913,I55631);
nand I_10490 (I180964,I180947,I55652);
nor I_10491 (I180729,I180964,I180913);
and I_10492 (I180720,I180806,I180964);
not I_10493 (I181009,I180964);
nand I_10494 (I180723,I180806,I181009);
nor I_10495 (I180717,I180772,I180964);
not I_10496 (I181054,I55640);
nor I_10497 (I181071,I181054,I55631);
nand I_10498 (I181088,I181071,I180913);
nor I_10499 (I180726,I180831,I181088);
nor I_10500 (I181119,I181054,I55634);
and I_10501 (I181136,I181119,I55649);
or I_10502 (I181153,I181136,I55637);
DFFARX1 I_10503 (I181153,I2595,I180746,I181179,);
nor I_10504 (I181187,I181179,I180930);
DFFARX1 I_10505 (I181187,I2595,I180746,I180714,);
DFFARX1 I_10506 (I181179,I2595,I180746,I180738,);
not I_10507 (I181232,I181179);
nor I_10508 (I181249,I181232,I180806);
nor I_10509 (I181266,I181071,I181249);
DFFARX1 I_10510 (I181266,I2595,I180746,I180735,);
not I_10511 (I181324,I2602);
DFFARX1 I_10512 (I14500,I2595,I181324,I181350,);
not I_10513 (I181358,I181350);
nand I_10514 (I181375,I14497,I14488);
and I_10515 (I181392,I181375,I14488);
DFFARX1 I_10516 (I181392,I2595,I181324,I181418,);
not I_10517 (I181426,I14491);
DFFARX1 I_10518 (I14506,I2595,I181324,I181452,);
not I_10519 (I181460,I181452);
nor I_10520 (I181477,I181460,I181358);
and I_10521 (I181494,I181477,I14491);
nor I_10522 (I181511,I181460,I181426);
nor I_10523 (I181307,I181418,I181511);
DFFARX1 I_10524 (I14491,I2595,I181324,I181551,);
nor I_10525 (I181559,I181551,I181418);
not I_10526 (I181576,I181559);
not I_10527 (I181593,I181551);
nor I_10528 (I181610,I181593,I181494);
DFFARX1 I_10529 (I181610,I2595,I181324,I181310,);
nand I_10530 (I181641,I14509,I14494);
and I_10531 (I181658,I181641,I14512);
DFFARX1 I_10532 (I181658,I2595,I181324,I181684,);
nor I_10533 (I181692,I181684,I181551);
DFFARX1 I_10534 (I181692,I2595,I181324,I181292,);
nand I_10535 (I181723,I181684,I181593);
nand I_10536 (I181301,I181576,I181723);
not I_10537 (I181754,I181684);
nor I_10538 (I181771,I181754,I181494);
DFFARX1 I_10539 (I181771,I2595,I181324,I181313,);
nor I_10540 (I181802,I14503,I14494);
or I_10541 (I181304,I181551,I181802);
nor I_10542 (I181295,I181684,I181802);
or I_10543 (I181298,I181418,I181802);
DFFARX1 I_10544 (I181802,I2595,I181324,I181316,);
not I_10545 (I181902,I2602);
DFFARX1 I_10546 (I98033,I2595,I181902,I181928,);
not I_10547 (I181936,I181928);
nand I_10548 (I181953,I98036,I98012);
and I_10549 (I181970,I181953,I98009);
DFFARX1 I_10550 (I181970,I2595,I181902,I181996,);
not I_10551 (I182004,I98015);
DFFARX1 I_10552 (I98009,I2595,I181902,I182030,);
not I_10553 (I182038,I182030);
nor I_10554 (I182055,I182038,I181936);
and I_10555 (I182072,I182055,I98015);
nor I_10556 (I182089,I182038,I182004);
nor I_10557 (I181885,I181996,I182089);
DFFARX1 I_10558 (I98018,I2595,I181902,I182129,);
nor I_10559 (I182137,I182129,I181996);
not I_10560 (I182154,I182137);
not I_10561 (I182171,I182129);
nor I_10562 (I182188,I182171,I182072);
DFFARX1 I_10563 (I182188,I2595,I181902,I181888,);
nand I_10564 (I182219,I98021,I98030);
and I_10565 (I182236,I182219,I98027);
DFFARX1 I_10566 (I182236,I2595,I181902,I182262,);
nor I_10567 (I182270,I182262,I182129);
DFFARX1 I_10568 (I182270,I2595,I181902,I181870,);
nand I_10569 (I182301,I182262,I182171);
nand I_10570 (I181879,I182154,I182301);
not I_10571 (I182332,I182262);
nor I_10572 (I182349,I182332,I182072);
DFFARX1 I_10573 (I182349,I2595,I181902,I181891,);
nor I_10574 (I182380,I98024,I98030);
or I_10575 (I181882,I182129,I182380);
nor I_10576 (I181873,I182262,I182380);
or I_10577 (I181876,I181996,I182380);
DFFARX1 I_10578 (I182380,I2595,I181902,I181894,);
not I_10579 (I182480,I2602);
DFFARX1 I_10580 (I97506,I2595,I182480,I182506,);
not I_10581 (I182514,I182506);
nand I_10582 (I182531,I97509,I97485);
and I_10583 (I182548,I182531,I97482);
DFFARX1 I_10584 (I182548,I2595,I182480,I182574,);
not I_10585 (I182582,I97488);
DFFARX1 I_10586 (I97482,I2595,I182480,I182608,);
not I_10587 (I182616,I182608);
nor I_10588 (I182633,I182616,I182514);
and I_10589 (I182650,I182633,I97488);
nor I_10590 (I182667,I182616,I182582);
nor I_10591 (I182463,I182574,I182667);
DFFARX1 I_10592 (I97491,I2595,I182480,I182707,);
nor I_10593 (I182715,I182707,I182574);
not I_10594 (I182732,I182715);
not I_10595 (I182749,I182707);
nor I_10596 (I182766,I182749,I182650);
DFFARX1 I_10597 (I182766,I2595,I182480,I182466,);
nand I_10598 (I182797,I97494,I97503);
and I_10599 (I182814,I182797,I97500);
DFFARX1 I_10600 (I182814,I2595,I182480,I182840,);
nor I_10601 (I182848,I182840,I182707);
DFFARX1 I_10602 (I182848,I2595,I182480,I182448,);
nand I_10603 (I182879,I182840,I182749);
nand I_10604 (I182457,I182732,I182879);
not I_10605 (I182910,I182840);
nor I_10606 (I182927,I182910,I182650);
DFFARX1 I_10607 (I182927,I2595,I182480,I182469,);
nor I_10608 (I182958,I97497,I97503);
or I_10609 (I182460,I182707,I182958);
nor I_10610 (I182451,I182840,I182958);
or I_10611 (I182454,I182574,I182958);
DFFARX1 I_10612 (I182958,I2595,I182480,I182472,);
not I_10613 (I183058,I2602);
DFFARX1 I_10614 (I146340,I2595,I183058,I183084,);
not I_10615 (I183092,I183084);
nand I_10616 (I183109,I146355,I146340);
and I_10617 (I183126,I183109,I146343);
DFFARX1 I_10618 (I183126,I2595,I183058,I183152,);
not I_10619 (I183160,I146343);
DFFARX1 I_10620 (I146352,I2595,I183058,I183186,);
not I_10621 (I183194,I183186);
nor I_10622 (I183211,I183194,I183092);
and I_10623 (I183228,I183211,I146343);
nor I_10624 (I183245,I183194,I183160);
nor I_10625 (I183041,I183152,I183245);
DFFARX1 I_10626 (I146346,I2595,I183058,I183285,);
nor I_10627 (I183293,I183285,I183152);
not I_10628 (I183310,I183293);
not I_10629 (I183327,I183285);
nor I_10630 (I183344,I183327,I183228);
DFFARX1 I_10631 (I183344,I2595,I183058,I183044,);
nand I_10632 (I183375,I146349,I146358);
and I_10633 (I183392,I183375,I146364);
DFFARX1 I_10634 (I183392,I2595,I183058,I183418,);
nor I_10635 (I183426,I183418,I183285);
DFFARX1 I_10636 (I183426,I2595,I183058,I183026,);
nand I_10637 (I183457,I183418,I183327);
nand I_10638 (I183035,I183310,I183457);
not I_10639 (I183488,I183418);
nor I_10640 (I183505,I183488,I183228);
DFFARX1 I_10641 (I183505,I2595,I183058,I183047,);
nor I_10642 (I183536,I146361,I146358);
or I_10643 (I183038,I183285,I183536);
nor I_10644 (I183029,I183418,I183536);
or I_10645 (I183032,I183152,I183536);
DFFARX1 I_10646 (I183536,I2595,I183058,I183050,);
not I_10647 (I183636,I2602);
DFFARX1 I_10648 (I47310,I2595,I183636,I183662,);
not I_10649 (I183670,I183662);
nand I_10650 (I183687,I47325,I47298);
and I_10651 (I183704,I183687,I47313);
DFFARX1 I_10652 (I183704,I2595,I183636,I183730,);
not I_10653 (I183738,I47316);
DFFARX1 I_10654 (I47301,I2595,I183636,I183764,);
not I_10655 (I183772,I183764);
nor I_10656 (I183789,I183772,I183670);
and I_10657 (I183806,I183789,I47316);
nor I_10658 (I183823,I183772,I183738);
nor I_10659 (I183619,I183730,I183823);
DFFARX1 I_10660 (I47307,I2595,I183636,I183863,);
nor I_10661 (I183871,I183863,I183730);
not I_10662 (I183888,I183871);
not I_10663 (I183905,I183863);
nor I_10664 (I183922,I183905,I183806);
DFFARX1 I_10665 (I183922,I2595,I183636,I183622,);
nand I_10666 (I183953,I47322,I47304);
and I_10667 (I183970,I183953,I47319);
DFFARX1 I_10668 (I183970,I2595,I183636,I183996,);
nor I_10669 (I184004,I183996,I183863);
DFFARX1 I_10670 (I184004,I2595,I183636,I183604,);
nand I_10671 (I184035,I183996,I183905);
nand I_10672 (I183613,I183888,I184035);
not I_10673 (I184066,I183996);
nor I_10674 (I184083,I184066,I183806);
DFFARX1 I_10675 (I184083,I2595,I183636,I183625,);
nor I_10676 (I184114,I47298,I47304);
or I_10677 (I183616,I183863,I184114);
nor I_10678 (I183607,I183996,I184114);
or I_10679 (I183610,I183730,I184114);
DFFARX1 I_10680 (I184114,I2595,I183636,I183628,);
not I_10681 (I184214,I2602);
DFFARX1 I_10682 (I35571,I2595,I184214,I184240,);
not I_10683 (I184248,I184240);
nand I_10684 (I184265,I35580,I35589);
and I_10685 (I184282,I184265,I35568);
DFFARX1 I_10686 (I184282,I2595,I184214,I184308,);
not I_10687 (I184316,I35571);
DFFARX1 I_10688 (I35586,I2595,I184214,I184342,);
not I_10689 (I184350,I184342);
nor I_10690 (I184367,I184350,I184248);
and I_10691 (I184384,I184367,I35571);
nor I_10692 (I184401,I184350,I184316);
nor I_10693 (I184197,I184308,I184401);
DFFARX1 I_10694 (I35577,I2595,I184214,I184441,);
nor I_10695 (I184449,I184441,I184308);
not I_10696 (I184466,I184449);
not I_10697 (I184483,I184441);
nor I_10698 (I184500,I184483,I184384);
DFFARX1 I_10699 (I184500,I2595,I184214,I184200,);
nand I_10700 (I184531,I35592,I35568);
and I_10701 (I184548,I184531,I35574);
DFFARX1 I_10702 (I184548,I2595,I184214,I184574,);
nor I_10703 (I184582,I184574,I184441);
DFFARX1 I_10704 (I184582,I2595,I184214,I184182,);
nand I_10705 (I184613,I184574,I184483);
nand I_10706 (I184191,I184466,I184613);
not I_10707 (I184644,I184574);
nor I_10708 (I184661,I184644,I184384);
DFFARX1 I_10709 (I184661,I2595,I184214,I184203,);
nor I_10710 (I184692,I35583,I35568);
or I_10711 (I184194,I184441,I184692);
nor I_10712 (I184185,I184574,I184692);
or I_10713 (I184188,I184308,I184692);
DFFARX1 I_10714 (I184692,I2595,I184214,I184206,);
not I_10715 (I184792,I2602);
DFFARX1 I_10716 (I174356,I2595,I184792,I184818,);
not I_10717 (I184826,I184818);
nand I_10718 (I184843,I174365,I174374);
and I_10719 (I184860,I184843,I174380);
DFFARX1 I_10720 (I184860,I2595,I184792,I184886,);
not I_10721 (I184894,I174377);
DFFARX1 I_10722 (I174362,I2595,I184792,I184920,);
not I_10723 (I184928,I184920);
nor I_10724 (I184945,I184928,I184826);
and I_10725 (I184962,I184945,I174377);
nor I_10726 (I184979,I184928,I184894);
nor I_10727 (I184775,I184886,I184979);
DFFARX1 I_10728 (I174371,I2595,I184792,I185019,);
nor I_10729 (I185027,I185019,I184886);
not I_10730 (I185044,I185027);
not I_10731 (I185061,I185019);
nor I_10732 (I185078,I185061,I184962);
DFFARX1 I_10733 (I185078,I2595,I184792,I184778,);
nand I_10734 (I185109,I174368,I174359);
and I_10735 (I185126,I185109,I174356);
DFFARX1 I_10736 (I185126,I2595,I184792,I185152,);
nor I_10737 (I185160,I185152,I185019);
DFFARX1 I_10738 (I185160,I2595,I184792,I184760,);
nand I_10739 (I185191,I185152,I185061);
nand I_10740 (I184769,I185044,I185191);
not I_10741 (I185222,I185152);
nor I_10742 (I185239,I185222,I184962);
DFFARX1 I_10743 (I185239,I2595,I184792,I184781,);
nor I_10744 (I185270,I174359,I174359);
or I_10745 (I184772,I185019,I185270);
nor I_10746 (I184763,I185152,I185270);
or I_10747 (I184766,I184886,I185270);
DFFARX1 I_10748 (I185270,I2595,I184792,I184784,);
not I_10749 (I185370,I2602);
DFFARX1 I_10750 (I86966,I2595,I185370,I185396,);
not I_10751 (I185404,I185396);
nand I_10752 (I185421,I86969,I86945);
and I_10753 (I185438,I185421,I86942);
DFFARX1 I_10754 (I185438,I2595,I185370,I185464,);
not I_10755 (I185472,I86948);
DFFARX1 I_10756 (I86942,I2595,I185370,I185498,);
not I_10757 (I185506,I185498);
nor I_10758 (I185523,I185506,I185404);
and I_10759 (I185540,I185523,I86948);
nor I_10760 (I185557,I185506,I185472);
nor I_10761 (I185353,I185464,I185557);
DFFARX1 I_10762 (I86951,I2595,I185370,I185597,);
nor I_10763 (I185605,I185597,I185464);
not I_10764 (I185622,I185605);
not I_10765 (I185639,I185597);
nor I_10766 (I185656,I185639,I185540);
DFFARX1 I_10767 (I185656,I2595,I185370,I185356,);
nand I_10768 (I185687,I86954,I86963);
and I_10769 (I185704,I185687,I86960);
DFFARX1 I_10770 (I185704,I2595,I185370,I185730,);
nor I_10771 (I185738,I185730,I185597);
DFFARX1 I_10772 (I185738,I2595,I185370,I185338,);
nand I_10773 (I185769,I185730,I185639);
nand I_10774 (I185347,I185622,I185769);
not I_10775 (I185800,I185730);
nor I_10776 (I185817,I185800,I185540);
DFFARX1 I_10777 (I185817,I2595,I185370,I185359,);
nor I_10778 (I185848,I86957,I86963);
or I_10779 (I185350,I185597,I185848);
nor I_10780 (I185341,I185730,I185848);
or I_10781 (I185344,I185464,I185848);
DFFARX1 I_10782 (I185848,I2595,I185370,I185362,);
not I_10783 (I185948,I2602);
DFFARX1 I_10784 (I298309,I2595,I185948,I185974,);
not I_10785 (I185982,I185974);
nand I_10786 (I185999,I298306,I298324);
and I_10787 (I186016,I185999,I298321);
DFFARX1 I_10788 (I186016,I2595,I185948,I186042,);
not I_10789 (I186050,I298303);
DFFARX1 I_10790 (I298306,I2595,I185948,I186076,);
not I_10791 (I186084,I186076);
nor I_10792 (I186101,I186084,I185982);
and I_10793 (I186118,I186101,I298303);
nor I_10794 (I186135,I186084,I186050);
nor I_10795 (I185931,I186042,I186135);
DFFARX1 I_10796 (I298315,I2595,I185948,I186175,);
nor I_10797 (I186183,I186175,I186042);
not I_10798 (I186200,I186183);
not I_10799 (I186217,I186175);
nor I_10800 (I186234,I186217,I186118);
DFFARX1 I_10801 (I186234,I2595,I185948,I185934,);
nand I_10802 (I186265,I298318,I298303);
and I_10803 (I186282,I186265,I298309);
DFFARX1 I_10804 (I186282,I2595,I185948,I186308,);
nor I_10805 (I186316,I186308,I186175);
DFFARX1 I_10806 (I186316,I2595,I185948,I185916,);
nand I_10807 (I186347,I186308,I186217);
nand I_10808 (I185925,I186200,I186347);
not I_10809 (I186378,I186308);
nor I_10810 (I186395,I186378,I186118);
DFFARX1 I_10811 (I186395,I2595,I185948,I185937,);
nor I_10812 (I186426,I298312,I298303);
or I_10813 (I185928,I186175,I186426);
nor I_10814 (I185919,I186308,I186426);
or I_10815 (I185922,I186042,I186426);
DFFARX1 I_10816 (I186426,I2595,I185948,I185940,);
not I_10817 (I186526,I2602);
DFFARX1 I_10818 (I374150,I2595,I186526,I186552,);
not I_10819 (I186560,I186552);
nand I_10820 (I186577,I374135,I374123);
and I_10821 (I186594,I186577,I374138);
DFFARX1 I_10822 (I186594,I2595,I186526,I186620,);
not I_10823 (I186628,I374123);
DFFARX1 I_10824 (I374141,I2595,I186526,I186654,);
not I_10825 (I186662,I186654);
nor I_10826 (I186679,I186662,I186560);
and I_10827 (I186696,I186679,I374123);
nor I_10828 (I186713,I186662,I186628);
nor I_10829 (I186509,I186620,I186713);
DFFARX1 I_10830 (I374129,I2595,I186526,I186753,);
nor I_10831 (I186761,I186753,I186620);
not I_10832 (I186778,I186761);
not I_10833 (I186795,I186753);
nor I_10834 (I186812,I186795,I186696);
DFFARX1 I_10835 (I186812,I2595,I186526,I186512,);
nand I_10836 (I186843,I374126,I374132);
and I_10837 (I186860,I186843,I374147);
DFFARX1 I_10838 (I186860,I2595,I186526,I186886,);
nor I_10839 (I186894,I186886,I186753);
DFFARX1 I_10840 (I186894,I2595,I186526,I186494,);
nand I_10841 (I186925,I186886,I186795);
nand I_10842 (I186503,I186778,I186925);
not I_10843 (I186956,I186886);
nor I_10844 (I186973,I186956,I186696);
DFFARX1 I_10845 (I186973,I2595,I186526,I186515,);
nor I_10846 (I187004,I374144,I374132);
or I_10847 (I186506,I186753,I187004);
nor I_10848 (I186497,I186886,I187004);
or I_10849 (I186500,I186620,I187004);
DFFARX1 I_10850 (I187004,I2595,I186526,I186518,);
not I_10851 (I187104,I2602);
DFFARX1 I_10852 (I381885,I2595,I187104,I187130,);
not I_10853 (I187138,I187130);
nand I_10854 (I187155,I381870,I381858);
and I_10855 (I187172,I187155,I381873);
DFFARX1 I_10856 (I187172,I2595,I187104,I187198,);
not I_10857 (I187206,I381858);
DFFARX1 I_10858 (I381876,I2595,I187104,I187232,);
not I_10859 (I187240,I187232);
nor I_10860 (I187257,I187240,I187138);
and I_10861 (I187274,I187257,I381858);
nor I_10862 (I187291,I187240,I187206);
nor I_10863 (I187087,I187198,I187291);
DFFARX1 I_10864 (I381864,I2595,I187104,I187331,);
nor I_10865 (I187339,I187331,I187198);
not I_10866 (I187356,I187339);
not I_10867 (I187373,I187331);
nor I_10868 (I187390,I187373,I187274);
DFFARX1 I_10869 (I187390,I2595,I187104,I187090,);
nand I_10870 (I187421,I381861,I381867);
and I_10871 (I187438,I187421,I381882);
DFFARX1 I_10872 (I187438,I2595,I187104,I187464,);
nor I_10873 (I187472,I187464,I187331);
DFFARX1 I_10874 (I187472,I2595,I187104,I187072,);
nand I_10875 (I187503,I187464,I187373);
nand I_10876 (I187081,I187356,I187503);
not I_10877 (I187534,I187464);
nor I_10878 (I187551,I187534,I187274);
DFFARX1 I_10879 (I187551,I2595,I187104,I187093,);
nor I_10880 (I187582,I381879,I381867);
or I_10881 (I187084,I187331,I187582);
nor I_10882 (I187075,I187464,I187582);
or I_10883 (I187078,I187198,I187582);
DFFARX1 I_10884 (I187582,I2595,I187104,I187096,);
not I_10885 (I187682,I2602);
DFFARX1 I_10886 (I144555,I2595,I187682,I187708,);
not I_10887 (I187716,I187708);
nand I_10888 (I187733,I144570,I144555);
and I_10889 (I187750,I187733,I144558);
DFFARX1 I_10890 (I187750,I2595,I187682,I187776,);
not I_10891 (I187784,I144558);
DFFARX1 I_10892 (I144567,I2595,I187682,I187810,);
not I_10893 (I187818,I187810);
nor I_10894 (I187835,I187818,I187716);
and I_10895 (I187852,I187835,I144558);
nor I_10896 (I187869,I187818,I187784);
nor I_10897 (I187665,I187776,I187869);
DFFARX1 I_10898 (I144561,I2595,I187682,I187909,);
nor I_10899 (I187917,I187909,I187776);
not I_10900 (I187934,I187917);
not I_10901 (I187951,I187909);
nor I_10902 (I187968,I187951,I187852);
DFFARX1 I_10903 (I187968,I2595,I187682,I187668,);
nand I_10904 (I187999,I144564,I144573);
and I_10905 (I188016,I187999,I144579);
DFFARX1 I_10906 (I188016,I2595,I187682,I188042,);
nor I_10907 (I188050,I188042,I187909);
DFFARX1 I_10908 (I188050,I2595,I187682,I187650,);
nand I_10909 (I188081,I188042,I187951);
nand I_10910 (I187659,I187934,I188081);
not I_10911 (I188112,I188042);
nor I_10912 (I188129,I188112,I187852);
DFFARX1 I_10913 (I188129,I2595,I187682,I187671,);
nor I_10914 (I188160,I144576,I144573);
or I_10915 (I187662,I187909,I188160);
nor I_10916 (I187653,I188042,I188160);
or I_10917 (I187656,I187776,I188160);
DFFARX1 I_10918 (I188160,I2595,I187682,I187674,);
not I_10919 (I188260,I2602);
DFFARX1 I_10920 (I255113,I2595,I188260,I188286,);
not I_10921 (I188294,I188286);
nand I_10922 (I188311,I255089,I255104);
and I_10923 (I188328,I188311,I255116);
DFFARX1 I_10924 (I188328,I2595,I188260,I188354,);
not I_10925 (I188362,I255101);
DFFARX1 I_10926 (I255092,I2595,I188260,I188388,);
not I_10927 (I188396,I188388);
nor I_10928 (I188413,I188396,I188294);
and I_10929 (I188430,I188413,I255101);
nor I_10930 (I188447,I188396,I188362);
nor I_10931 (I188243,I188354,I188447);
DFFARX1 I_10932 (I255089,I2595,I188260,I188487,);
nor I_10933 (I188495,I188487,I188354);
not I_10934 (I188512,I188495);
not I_10935 (I188529,I188487);
nor I_10936 (I188546,I188529,I188430);
DFFARX1 I_10937 (I188546,I2595,I188260,I188246,);
nand I_10938 (I188577,I255107,I255098);
and I_10939 (I188594,I188577,I255110);
DFFARX1 I_10940 (I188594,I2595,I188260,I188620,);
nor I_10941 (I188628,I188620,I188487);
DFFARX1 I_10942 (I188628,I2595,I188260,I188228,);
nand I_10943 (I188659,I188620,I188529);
nand I_10944 (I188237,I188512,I188659);
not I_10945 (I188690,I188620);
nor I_10946 (I188707,I188690,I188430);
DFFARX1 I_10947 (I188707,I2595,I188260,I188249,);
nor I_10948 (I188738,I255095,I255098);
or I_10949 (I188240,I188487,I188738);
nor I_10950 (I188231,I188620,I188738);
or I_10951 (I188234,I188354,I188738);
DFFARX1 I_10952 (I188738,I2595,I188260,I188252,);
not I_10953 (I188838,I2602);
DFFARX1 I_10954 (I231967,I2595,I188838,I188864,);
not I_10955 (I188872,I188864);
nand I_10956 (I188889,I231955,I231973);
and I_10957 (I188906,I188889,I231970);
DFFARX1 I_10958 (I188906,I2595,I188838,I188932,);
not I_10959 (I188940,I231961);
DFFARX1 I_10960 (I231958,I2595,I188838,I188966,);
not I_10961 (I188974,I188966);
nor I_10962 (I188991,I188974,I188872);
and I_10963 (I189008,I188991,I231961);
nor I_10964 (I189025,I188974,I188940);
nor I_10965 (I188821,I188932,I189025);
DFFARX1 I_10966 (I231952,I2595,I188838,I189065,);
nor I_10967 (I189073,I189065,I188932);
not I_10968 (I189090,I189073);
not I_10969 (I189107,I189065);
nor I_10970 (I189124,I189107,I189008);
DFFARX1 I_10971 (I189124,I2595,I188838,I188824,);
nand I_10972 (I189155,I231952,I231955);
and I_10973 (I189172,I189155,I231958);
DFFARX1 I_10974 (I189172,I2595,I188838,I189198,);
nor I_10975 (I189206,I189198,I189065);
DFFARX1 I_10976 (I189206,I2595,I188838,I188806,);
nand I_10977 (I189237,I189198,I189107);
nand I_10978 (I188815,I189090,I189237);
not I_10979 (I189268,I189198);
nor I_10980 (I189285,I189268,I189008);
DFFARX1 I_10981 (I189285,I2595,I188838,I188827,);
nor I_10982 (I189316,I231964,I231955);
or I_10983 (I188818,I189065,I189316);
nor I_10984 (I188809,I189198,I189316);
or I_10985 (I188812,I188932,I189316);
DFFARX1 I_10986 (I189316,I2595,I188838,I188830,);
not I_10987 (I189416,I2602);
DFFARX1 I_10988 (I43476,I2595,I189416,I189442,);
not I_10989 (I189450,I189442);
nand I_10990 (I189467,I43485,I43494);
and I_10991 (I189484,I189467,I43473);
DFFARX1 I_10992 (I189484,I2595,I189416,I189510,);
not I_10993 (I189518,I43476);
DFFARX1 I_10994 (I43491,I2595,I189416,I189544,);
not I_10995 (I189552,I189544);
nor I_10996 (I189569,I189552,I189450);
and I_10997 (I189586,I189569,I43476);
nor I_10998 (I189603,I189552,I189518);
nor I_10999 (I189399,I189510,I189603);
DFFARX1 I_11000 (I43482,I2595,I189416,I189643,);
nor I_11001 (I189651,I189643,I189510);
not I_11002 (I189668,I189651);
not I_11003 (I189685,I189643);
nor I_11004 (I189702,I189685,I189586);
DFFARX1 I_11005 (I189702,I2595,I189416,I189402,);
nand I_11006 (I189733,I43497,I43473);
and I_11007 (I189750,I189733,I43479);
DFFARX1 I_11008 (I189750,I2595,I189416,I189776,);
nor I_11009 (I189784,I189776,I189643);
DFFARX1 I_11010 (I189784,I2595,I189416,I189384,);
nand I_11011 (I189815,I189776,I189685);
nand I_11012 (I189393,I189668,I189815);
not I_11013 (I189846,I189776);
nor I_11014 (I189863,I189846,I189586);
DFFARX1 I_11015 (I189863,I2595,I189416,I189405,);
nor I_11016 (I189894,I43488,I43473);
or I_11017 (I189396,I189643,I189894);
nor I_11018 (I189387,I189776,I189894);
or I_11019 (I189390,I189510,I189894);
DFFARX1 I_11020 (I189894,I2595,I189416,I189408,);
not I_11021 (I189994,I2602);
DFFARX1 I_11022 (I81169,I2595,I189994,I190020,);
not I_11023 (I190028,I190020);
nand I_11024 (I190045,I81172,I81148);
and I_11025 (I190062,I190045,I81145);
DFFARX1 I_11026 (I190062,I2595,I189994,I190088,);
not I_11027 (I190096,I81151);
DFFARX1 I_11028 (I81145,I2595,I189994,I190122,);
not I_11029 (I190130,I190122);
nor I_11030 (I190147,I190130,I190028);
and I_11031 (I190164,I190147,I81151);
nor I_11032 (I190181,I190130,I190096);
nor I_11033 (I189977,I190088,I190181);
DFFARX1 I_11034 (I81154,I2595,I189994,I190221,);
nor I_11035 (I190229,I190221,I190088);
not I_11036 (I190246,I190229);
not I_11037 (I190263,I190221);
nor I_11038 (I190280,I190263,I190164);
DFFARX1 I_11039 (I190280,I2595,I189994,I189980,);
nand I_11040 (I190311,I81157,I81166);
and I_11041 (I190328,I190311,I81163);
DFFARX1 I_11042 (I190328,I2595,I189994,I190354,);
nor I_11043 (I190362,I190354,I190221);
DFFARX1 I_11044 (I190362,I2595,I189994,I189962,);
nand I_11045 (I190393,I190354,I190263);
nand I_11046 (I189971,I190246,I190393);
not I_11047 (I190424,I190354);
nor I_11048 (I190441,I190424,I190164);
DFFARX1 I_11049 (I190441,I2595,I189994,I189983,);
nor I_11050 (I190472,I81160,I81166);
or I_11051 (I189974,I190221,I190472);
nor I_11052 (I189965,I190354,I190472);
or I_11053 (I189968,I190088,I190472);
DFFARX1 I_11054 (I190472,I2595,I189994,I189986,);
not I_11055 (I190572,I2602);
DFFARX1 I_11056 (I21351,I2595,I190572,I190598,);
not I_11057 (I190606,I190598);
nand I_11058 (I190623,I21348,I21339);
and I_11059 (I190640,I190623,I21339);
DFFARX1 I_11060 (I190640,I2595,I190572,I190666,);
not I_11061 (I190674,I21342);
DFFARX1 I_11062 (I21357,I2595,I190572,I190700,);
not I_11063 (I190708,I190700);
nor I_11064 (I190725,I190708,I190606);
and I_11065 (I190742,I190725,I21342);
nor I_11066 (I190759,I190708,I190674);
nor I_11067 (I190555,I190666,I190759);
DFFARX1 I_11068 (I21342,I2595,I190572,I190799,);
nor I_11069 (I190807,I190799,I190666);
not I_11070 (I190824,I190807);
not I_11071 (I190841,I190799);
nor I_11072 (I190858,I190841,I190742);
DFFARX1 I_11073 (I190858,I2595,I190572,I190558,);
nand I_11074 (I190889,I21360,I21345);
and I_11075 (I190906,I190889,I21363);
DFFARX1 I_11076 (I190906,I2595,I190572,I190932,);
nor I_11077 (I190940,I190932,I190799);
DFFARX1 I_11078 (I190940,I2595,I190572,I190540,);
nand I_11079 (I190971,I190932,I190841);
nand I_11080 (I190549,I190824,I190971);
not I_11081 (I191002,I190932);
nor I_11082 (I191019,I191002,I190742);
DFFARX1 I_11083 (I191019,I2595,I190572,I190561,);
nor I_11084 (I191050,I21354,I21345);
or I_11085 (I190552,I190799,I191050);
nor I_11086 (I190543,I190932,I191050);
or I_11087 (I190546,I190666,I191050);
DFFARX1 I_11088 (I191050,I2595,I190572,I190564,);
not I_11089 (I191150,I2602);
DFFARX1 I_11090 (I257697,I2595,I191150,I191176,);
not I_11091 (I191184,I191176);
nand I_11092 (I191201,I257673,I257688);
and I_11093 (I191218,I191201,I257700);
DFFARX1 I_11094 (I191218,I2595,I191150,I191244,);
not I_11095 (I191252,I257685);
DFFARX1 I_11096 (I257676,I2595,I191150,I191278,);
not I_11097 (I191286,I191278);
nor I_11098 (I191303,I191286,I191184);
and I_11099 (I191320,I191303,I257685);
nor I_11100 (I191337,I191286,I191252);
nor I_11101 (I191133,I191244,I191337);
DFFARX1 I_11102 (I257673,I2595,I191150,I191377,);
nor I_11103 (I191385,I191377,I191244);
not I_11104 (I191402,I191385);
not I_11105 (I191419,I191377);
nor I_11106 (I191436,I191419,I191320);
DFFARX1 I_11107 (I191436,I2595,I191150,I191136,);
nand I_11108 (I191467,I257691,I257682);
and I_11109 (I191484,I191467,I257694);
DFFARX1 I_11110 (I191484,I2595,I191150,I191510,);
nor I_11111 (I191518,I191510,I191377);
DFFARX1 I_11112 (I191518,I2595,I191150,I191118,);
nand I_11113 (I191549,I191510,I191419);
nand I_11114 (I191127,I191402,I191549);
not I_11115 (I191580,I191510);
nor I_11116 (I191597,I191580,I191320);
DFFARX1 I_11117 (I191597,I2595,I191150,I191139,);
nor I_11118 (I191628,I257679,I257682);
or I_11119 (I191130,I191377,I191628);
nor I_11120 (I191121,I191510,I191628);
or I_11121 (I191124,I191244,I191628);
DFFARX1 I_11122 (I191628,I2595,I191150,I191142,);
not I_11123 (I191728,I2602);
DFFARX1 I_11124 (I128482,I2595,I191728,I191754,);
not I_11125 (I191762,I191754);
nand I_11126 (I191779,I128473,I128491);
and I_11127 (I191796,I191779,I128494);
DFFARX1 I_11128 (I191796,I2595,I191728,I191822,);
not I_11129 (I191830,I128488);
DFFARX1 I_11130 (I128476,I2595,I191728,I191856,);
not I_11131 (I191864,I191856);
nor I_11132 (I191881,I191864,I191762);
and I_11133 (I191898,I191881,I128488);
nor I_11134 (I191915,I191864,I191830);
nor I_11135 (I191711,I191822,I191915);
DFFARX1 I_11136 (I128485,I2595,I191728,I191955,);
nor I_11137 (I191963,I191955,I191822);
not I_11138 (I191980,I191963);
not I_11139 (I191997,I191955);
nor I_11140 (I192014,I191997,I191898);
DFFARX1 I_11141 (I192014,I2595,I191728,I191714,);
nand I_11142 (I192045,I128500,I128497);
and I_11143 (I192062,I192045,I128479);
DFFARX1 I_11144 (I192062,I2595,I191728,I192088,);
nor I_11145 (I192096,I192088,I191955);
DFFARX1 I_11146 (I192096,I2595,I191728,I191696,);
nand I_11147 (I192127,I192088,I191997);
nand I_11148 (I191705,I191980,I192127);
not I_11149 (I192158,I192088);
nor I_11150 (I192175,I192158,I191898);
DFFARX1 I_11151 (I192175,I2595,I191728,I191717,);
nor I_11152 (I192206,I128473,I128497);
or I_11153 (I191708,I191955,I192206);
nor I_11154 (I191699,I192088,I192206);
or I_11155 (I191702,I191822,I192206);
DFFARX1 I_11156 (I192206,I2595,I191728,I191720,);
not I_11157 (I192306,I2602);
DFFARX1 I_11158 (I89601,I2595,I192306,I192332,);
not I_11159 (I192340,I192332);
nand I_11160 (I192357,I89604,I89580);
and I_11161 (I192374,I192357,I89577);
DFFARX1 I_11162 (I192374,I2595,I192306,I192400,);
not I_11163 (I192408,I89583);
DFFARX1 I_11164 (I89577,I2595,I192306,I192434,);
not I_11165 (I192442,I192434);
nor I_11166 (I192459,I192442,I192340);
and I_11167 (I192476,I192459,I89583);
nor I_11168 (I192493,I192442,I192408);
nor I_11169 (I192289,I192400,I192493);
DFFARX1 I_11170 (I89586,I2595,I192306,I192533,);
nor I_11171 (I192541,I192533,I192400);
not I_11172 (I192558,I192541);
not I_11173 (I192575,I192533);
nor I_11174 (I192592,I192575,I192476);
DFFARX1 I_11175 (I192592,I2595,I192306,I192292,);
nand I_11176 (I192623,I89589,I89598);
and I_11177 (I192640,I192623,I89595);
DFFARX1 I_11178 (I192640,I2595,I192306,I192666,);
nor I_11179 (I192674,I192666,I192533);
DFFARX1 I_11180 (I192674,I2595,I192306,I192274,);
nand I_11181 (I192705,I192666,I192575);
nand I_11182 (I192283,I192558,I192705);
not I_11183 (I192736,I192666);
nor I_11184 (I192753,I192736,I192476);
DFFARX1 I_11185 (I192753,I2595,I192306,I192295,);
nor I_11186 (I192784,I89592,I89598);
or I_11187 (I192286,I192533,I192784);
nor I_11188 (I192277,I192666,I192784);
or I_11189 (I192280,I192400,I192784);
DFFARX1 I_11190 (I192784,I2595,I192306,I192298,);
not I_11191 (I192884,I2602);
DFFARX1 I_11192 (I69908,I2595,I192884,I192910,);
not I_11193 (I192918,I192910);
nand I_11194 (I192935,I69911,I69932);
and I_11195 (I192952,I192935,I69920);
DFFARX1 I_11196 (I192952,I2595,I192884,I192978,);
not I_11197 (I192986,I69917);
DFFARX1 I_11198 (I69908,I2595,I192884,I193012,);
not I_11199 (I193020,I193012);
nor I_11200 (I193037,I193020,I192918);
and I_11201 (I193054,I193037,I69917);
nor I_11202 (I193071,I193020,I192986);
nor I_11203 (I192867,I192978,I193071);
DFFARX1 I_11204 (I69926,I2595,I192884,I193111,);
nor I_11205 (I193119,I193111,I192978);
not I_11206 (I193136,I193119);
not I_11207 (I193153,I193111);
nor I_11208 (I193170,I193153,I193054);
DFFARX1 I_11209 (I193170,I2595,I192884,I192870,);
nand I_11210 (I193201,I69911,I69914);
and I_11211 (I193218,I193201,I69923);
DFFARX1 I_11212 (I193218,I2595,I192884,I193244,);
nor I_11213 (I193252,I193244,I193111);
DFFARX1 I_11214 (I193252,I2595,I192884,I192852,);
nand I_11215 (I193283,I193244,I193153);
nand I_11216 (I192861,I193136,I193283);
not I_11217 (I193314,I193244);
nor I_11218 (I193331,I193314,I193054);
DFFARX1 I_11219 (I193331,I2595,I192884,I192873,);
nor I_11220 (I193362,I69929,I69914);
or I_11221 (I192864,I193111,I193362);
nor I_11222 (I192855,I193244,I193362);
or I_11223 (I192858,I192978,I193362);
DFFARX1 I_11224 (I193362,I2595,I192884,I192876,);
not I_11225 (I193462,I2602);
DFFARX1 I_11226 (I309082,I2595,I193462,I193488,);
not I_11227 (I193496,I193488);
nand I_11228 (I193513,I309064,I309076);
and I_11229 (I193530,I193513,I309079);
DFFARX1 I_11230 (I193530,I2595,I193462,I193556,);
not I_11231 (I193564,I309073);
DFFARX1 I_11232 (I309070,I2595,I193462,I193590,);
not I_11233 (I193598,I193590);
nor I_11234 (I193615,I193598,I193496);
and I_11235 (I193632,I193615,I309073);
nor I_11236 (I193649,I193598,I193564);
nor I_11237 (I193445,I193556,I193649);
DFFARX1 I_11238 (I309088,I2595,I193462,I193689,);
nor I_11239 (I193697,I193689,I193556);
not I_11240 (I193714,I193697);
not I_11241 (I193731,I193689);
nor I_11242 (I193748,I193731,I193632);
DFFARX1 I_11243 (I193748,I2595,I193462,I193448,);
nand I_11244 (I193779,I309067,I309067);
and I_11245 (I193796,I193779,I309064);
DFFARX1 I_11246 (I193796,I2595,I193462,I193822,);
nor I_11247 (I193830,I193822,I193689);
DFFARX1 I_11248 (I193830,I2595,I193462,I193430,);
nand I_11249 (I193861,I193822,I193731);
nand I_11250 (I193439,I193714,I193861);
not I_11251 (I193892,I193822);
nor I_11252 (I193909,I193892,I193632);
DFFARX1 I_11253 (I193909,I2595,I193462,I193451,);
nor I_11254 (I193940,I309085,I309067);
or I_11255 (I193442,I193689,I193940);
nor I_11256 (I193433,I193822,I193940);
or I_11257 (I193436,I193556,I193940);
DFFARX1 I_11258 (I193940,I2595,I193462,I193454,);
not I_11259 (I194040,I2602);
DFFARX1 I_11260 (I324688,I2595,I194040,I194066,);
not I_11261 (I194074,I194066);
nand I_11262 (I194091,I324670,I324682);
and I_11263 (I194108,I194091,I324685);
DFFARX1 I_11264 (I194108,I2595,I194040,I194134,);
not I_11265 (I194142,I324679);
DFFARX1 I_11266 (I324676,I2595,I194040,I194168,);
not I_11267 (I194176,I194168);
nor I_11268 (I194193,I194176,I194074);
and I_11269 (I194210,I194193,I324679);
nor I_11270 (I194227,I194176,I194142);
nor I_11271 (I194023,I194134,I194227);
DFFARX1 I_11272 (I324694,I2595,I194040,I194267,);
nor I_11273 (I194275,I194267,I194134);
not I_11274 (I194292,I194275);
not I_11275 (I194309,I194267);
nor I_11276 (I194326,I194309,I194210);
DFFARX1 I_11277 (I194326,I2595,I194040,I194026,);
nand I_11278 (I194357,I324673,I324673);
and I_11279 (I194374,I194357,I324670);
DFFARX1 I_11280 (I194374,I2595,I194040,I194400,);
nor I_11281 (I194408,I194400,I194267);
DFFARX1 I_11282 (I194408,I2595,I194040,I194008,);
nand I_11283 (I194439,I194400,I194309);
nand I_11284 (I194017,I194292,I194439);
not I_11285 (I194470,I194400);
nor I_11286 (I194487,I194470,I194210);
DFFARX1 I_11287 (I194487,I2595,I194040,I194029,);
nor I_11288 (I194518,I324691,I324673);
or I_11289 (I194020,I194267,I194518);
nor I_11290 (I194011,I194400,I194518);
or I_11291 (I194014,I194134,I194518);
DFFARX1 I_11292 (I194518,I2595,I194040,I194032,);
not I_11293 (I194618,I2602);
DFFARX1 I_11294 (I373555,I2595,I194618,I194644,);
not I_11295 (I194652,I194644);
nand I_11296 (I194669,I373540,I373528);
and I_11297 (I194686,I194669,I373543);
DFFARX1 I_11298 (I194686,I2595,I194618,I194712,);
not I_11299 (I194720,I373528);
DFFARX1 I_11300 (I373546,I2595,I194618,I194746,);
not I_11301 (I194754,I194746);
nor I_11302 (I194771,I194754,I194652);
and I_11303 (I194788,I194771,I373528);
nor I_11304 (I194805,I194754,I194720);
nor I_11305 (I194601,I194712,I194805);
DFFARX1 I_11306 (I373534,I2595,I194618,I194845,);
nor I_11307 (I194853,I194845,I194712);
not I_11308 (I194870,I194853);
not I_11309 (I194887,I194845);
nor I_11310 (I194904,I194887,I194788);
DFFARX1 I_11311 (I194904,I2595,I194618,I194604,);
nand I_11312 (I194935,I373531,I373537);
and I_11313 (I194952,I194935,I373552);
DFFARX1 I_11314 (I194952,I2595,I194618,I194978,);
nor I_11315 (I194986,I194978,I194845);
DFFARX1 I_11316 (I194986,I2595,I194618,I194586,);
nand I_11317 (I195017,I194978,I194887);
nand I_11318 (I194595,I194870,I195017);
not I_11319 (I195048,I194978);
nor I_11320 (I195065,I195048,I194788);
DFFARX1 I_11321 (I195065,I2595,I194618,I194607,);
nor I_11322 (I195096,I373549,I373537);
or I_11323 (I194598,I194845,I195096);
nor I_11324 (I194589,I194978,I195096);
or I_11325 (I194592,I194712,I195096);
DFFARX1 I_11326 (I195096,I2595,I194618,I194610,);
not I_11327 (I195196,I2602);
DFFARX1 I_11328 (I350238,I2595,I195196,I195222,);
not I_11329 (I195230,I195222);
nand I_11330 (I195247,I350241,I350250);
and I_11331 (I195264,I195247,I350253);
DFFARX1 I_11332 (I195264,I2595,I195196,I195290,);
not I_11333 (I195298,I350262);
DFFARX1 I_11334 (I350244,I2595,I195196,I195324,);
not I_11335 (I195332,I195324);
nor I_11336 (I195349,I195332,I195230);
and I_11337 (I195366,I195349,I350262);
nor I_11338 (I195383,I195332,I195298);
nor I_11339 (I195179,I195290,I195383);
DFFARX1 I_11340 (I350241,I2595,I195196,I195423,);
nor I_11341 (I195431,I195423,I195290);
not I_11342 (I195448,I195431);
not I_11343 (I195465,I195423);
nor I_11344 (I195482,I195465,I195366);
DFFARX1 I_11345 (I195482,I2595,I195196,I195182,);
nand I_11346 (I195513,I350259,I350238);
and I_11347 (I195530,I195513,I350256);
DFFARX1 I_11348 (I195530,I2595,I195196,I195556,);
nor I_11349 (I195564,I195556,I195423);
DFFARX1 I_11350 (I195564,I2595,I195196,I195164,);
nand I_11351 (I195595,I195556,I195465);
nand I_11352 (I195173,I195448,I195595);
not I_11353 (I195626,I195556);
nor I_11354 (I195643,I195626,I195366);
DFFARX1 I_11355 (I195643,I2595,I195196,I195185,);
nor I_11356 (I195674,I350247,I350238);
or I_11357 (I195176,I195423,I195674);
nor I_11358 (I195167,I195556,I195674);
or I_11359 (I195170,I195290,I195674);
DFFARX1 I_11360 (I195674,I2595,I195196,I195188,);
not I_11361 (I195774,I2602);
DFFARX1 I_11362 (I67528,I2595,I195774,I195800,);
not I_11363 (I195808,I195800);
nand I_11364 (I195825,I67531,I67552);
and I_11365 (I195842,I195825,I67540);
DFFARX1 I_11366 (I195842,I2595,I195774,I195868,);
not I_11367 (I195876,I67537);
DFFARX1 I_11368 (I67528,I2595,I195774,I195902,);
not I_11369 (I195910,I195902);
nor I_11370 (I195927,I195910,I195808);
and I_11371 (I195944,I195927,I67537);
nor I_11372 (I195961,I195910,I195876);
nor I_11373 (I195757,I195868,I195961);
DFFARX1 I_11374 (I67546,I2595,I195774,I196001,);
nor I_11375 (I196009,I196001,I195868);
not I_11376 (I196026,I196009);
not I_11377 (I196043,I196001);
nor I_11378 (I196060,I196043,I195944);
DFFARX1 I_11379 (I196060,I2595,I195774,I195760,);
nand I_11380 (I196091,I67531,I67534);
and I_11381 (I196108,I196091,I67543);
DFFARX1 I_11382 (I196108,I2595,I195774,I196134,);
nor I_11383 (I196142,I196134,I196001);
DFFARX1 I_11384 (I196142,I2595,I195774,I195742,);
nand I_11385 (I196173,I196134,I196043);
nand I_11386 (I195751,I196026,I196173);
not I_11387 (I196204,I196134);
nor I_11388 (I196221,I196204,I195944);
DFFARX1 I_11389 (I196221,I2595,I195774,I195763,);
nor I_11390 (I196252,I67549,I67534);
or I_11391 (I195754,I196001,I196252);
nor I_11392 (I195745,I196134,I196252);
or I_11393 (I195748,I195868,I196252);
DFFARX1 I_11394 (I196252,I2595,I195774,I195766,);
not I_11395 (I196352,I2602);
DFFARX1 I_11396 (I313706,I2595,I196352,I196378,);
not I_11397 (I196386,I196378);
nand I_11398 (I196403,I313688,I313700);
and I_11399 (I196420,I196403,I313703);
DFFARX1 I_11400 (I196420,I2595,I196352,I196446,);
not I_11401 (I196454,I313697);
DFFARX1 I_11402 (I313694,I2595,I196352,I196480,);
not I_11403 (I196488,I196480);
nor I_11404 (I196505,I196488,I196386);
and I_11405 (I196522,I196505,I313697);
nor I_11406 (I196539,I196488,I196454);
nor I_11407 (I196335,I196446,I196539);
DFFARX1 I_11408 (I313712,I2595,I196352,I196579,);
nor I_11409 (I196587,I196579,I196446);
not I_11410 (I196604,I196587);
not I_11411 (I196621,I196579);
nor I_11412 (I196638,I196621,I196522);
DFFARX1 I_11413 (I196638,I2595,I196352,I196338,);
nand I_11414 (I196669,I313691,I313691);
and I_11415 (I196686,I196669,I313688);
DFFARX1 I_11416 (I196686,I2595,I196352,I196712,);
nor I_11417 (I196720,I196712,I196579);
DFFARX1 I_11418 (I196720,I2595,I196352,I196320,);
nand I_11419 (I196751,I196712,I196621);
nand I_11420 (I196329,I196604,I196751);
not I_11421 (I196782,I196712);
nor I_11422 (I196799,I196782,I196522);
DFFARX1 I_11423 (I196799,I2595,I196352,I196341,);
nor I_11424 (I196830,I313709,I313691);
or I_11425 (I196332,I196579,I196830);
nor I_11426 (I196323,I196712,I196830);
or I_11427 (I196326,I196446,I196830);
DFFARX1 I_11428 (I196830,I2595,I196352,I196344,);
not I_11429 (I196930,I2602);
DFFARX1 I_11430 (I323532,I2595,I196930,I196956,);
not I_11431 (I196964,I196956);
nand I_11432 (I196981,I323514,I323526);
and I_11433 (I196998,I196981,I323529);
DFFARX1 I_11434 (I196998,I2595,I196930,I197024,);
not I_11435 (I197032,I323523);
DFFARX1 I_11436 (I323520,I2595,I196930,I197058,);
not I_11437 (I197066,I197058);
nor I_11438 (I197083,I197066,I196964);
and I_11439 (I197100,I197083,I323523);
nor I_11440 (I197117,I197066,I197032);
nor I_11441 (I196913,I197024,I197117);
DFFARX1 I_11442 (I323538,I2595,I196930,I197157,);
nor I_11443 (I197165,I197157,I197024);
not I_11444 (I197182,I197165);
not I_11445 (I197199,I197157);
nor I_11446 (I197216,I197199,I197100);
DFFARX1 I_11447 (I197216,I2595,I196930,I196916,);
nand I_11448 (I197247,I323517,I323517);
and I_11449 (I197264,I197247,I323514);
DFFARX1 I_11450 (I197264,I2595,I196930,I197290,);
nor I_11451 (I197298,I197290,I197157);
DFFARX1 I_11452 (I197298,I2595,I196930,I196898,);
nand I_11453 (I197329,I197290,I197199);
nand I_11454 (I196907,I197182,I197329);
not I_11455 (I197360,I197290);
nor I_11456 (I197377,I197360,I197100);
DFFARX1 I_11457 (I197377,I2595,I196930,I196919,);
nor I_11458 (I197408,I323535,I323517);
or I_11459 (I196910,I197157,I197408);
nor I_11460 (I196901,I197290,I197408);
or I_11461 (I196904,I197024,I197408);
DFFARX1 I_11462 (I197408,I2595,I196930,I196922,);
not I_11463 (I197508,I2602);
DFFARX1 I_11464 (I9757,I2595,I197508,I197534,);
not I_11465 (I197542,I197534);
nand I_11466 (I197559,I9754,I9745);
and I_11467 (I197576,I197559,I9745);
DFFARX1 I_11468 (I197576,I2595,I197508,I197602,);
not I_11469 (I197610,I9748);
DFFARX1 I_11470 (I9763,I2595,I197508,I197636,);
not I_11471 (I197644,I197636);
nor I_11472 (I197661,I197644,I197542);
and I_11473 (I197678,I197661,I9748);
nor I_11474 (I197695,I197644,I197610);
nor I_11475 (I197491,I197602,I197695);
DFFARX1 I_11476 (I9748,I2595,I197508,I197735,);
nor I_11477 (I197743,I197735,I197602);
not I_11478 (I197760,I197743);
not I_11479 (I197777,I197735);
nor I_11480 (I197794,I197777,I197678);
DFFARX1 I_11481 (I197794,I2595,I197508,I197494,);
nand I_11482 (I197825,I9766,I9751);
and I_11483 (I197842,I197825,I9769);
DFFARX1 I_11484 (I197842,I2595,I197508,I197868,);
nor I_11485 (I197876,I197868,I197735);
DFFARX1 I_11486 (I197876,I2595,I197508,I197476,);
nand I_11487 (I197907,I197868,I197777);
nand I_11488 (I197485,I197760,I197907);
not I_11489 (I197938,I197868);
nor I_11490 (I197955,I197938,I197678);
DFFARX1 I_11491 (I197955,I2595,I197508,I197497,);
nor I_11492 (I197986,I9760,I9751);
or I_11493 (I197488,I197735,I197986);
nor I_11494 (I197479,I197868,I197986);
or I_11495 (I197482,I197602,I197986);
DFFARX1 I_11496 (I197986,I2595,I197508,I197500,);
not I_11497 (I198086,I2602);
DFFARX1 I_11498 (I364280,I2595,I198086,I198112,);
not I_11499 (I198120,I198112);
nand I_11500 (I198137,I364304,I364286);
and I_11501 (I198154,I198137,I364292);
DFFARX1 I_11502 (I198154,I2595,I198086,I198180,);
not I_11503 (I198188,I364298);
DFFARX1 I_11504 (I364283,I2595,I198086,I198214,);
not I_11505 (I198222,I198214);
nor I_11506 (I198239,I198222,I198120);
and I_11507 (I198256,I198239,I364298);
nor I_11508 (I198273,I198222,I198188);
nor I_11509 (I198069,I198180,I198273);
DFFARX1 I_11510 (I364295,I2595,I198086,I198313,);
nor I_11511 (I198321,I198313,I198180);
not I_11512 (I198338,I198321);
not I_11513 (I198355,I198313);
nor I_11514 (I198372,I198355,I198256);
DFFARX1 I_11515 (I198372,I2595,I198086,I198072,);
nand I_11516 (I198403,I364301,I364289);
and I_11517 (I198420,I198403,I364283);
DFFARX1 I_11518 (I198420,I2595,I198086,I198446,);
nor I_11519 (I198454,I198446,I198313);
DFFARX1 I_11520 (I198454,I2595,I198086,I198054,);
nand I_11521 (I198485,I198446,I198355);
nand I_11522 (I198063,I198338,I198485);
not I_11523 (I198516,I198446);
nor I_11524 (I198533,I198516,I198256);
DFFARX1 I_11525 (I198533,I2595,I198086,I198075,);
nor I_11526 (I198564,I364280,I364289);
or I_11527 (I198066,I198313,I198564);
nor I_11528 (I198057,I198446,I198564);
or I_11529 (I198060,I198180,I198564);
DFFARX1 I_11530 (I198564,I2595,I198086,I198078,);
not I_11531 (I198664,I2602);
DFFARX1 I_11532 (I260281,I2595,I198664,I198690,);
not I_11533 (I198698,I198690);
nand I_11534 (I198715,I260257,I260272);
and I_11535 (I198732,I198715,I260284);
DFFARX1 I_11536 (I198732,I2595,I198664,I198758,);
not I_11537 (I198766,I260269);
DFFARX1 I_11538 (I260260,I2595,I198664,I198792,);
not I_11539 (I198800,I198792);
nor I_11540 (I198817,I198800,I198698);
and I_11541 (I198834,I198817,I260269);
nor I_11542 (I198851,I198800,I198766);
nor I_11543 (I198647,I198758,I198851);
DFFARX1 I_11544 (I260257,I2595,I198664,I198891,);
nor I_11545 (I198899,I198891,I198758);
not I_11546 (I198916,I198899);
not I_11547 (I198933,I198891);
nor I_11548 (I198950,I198933,I198834);
DFFARX1 I_11549 (I198950,I2595,I198664,I198650,);
nand I_11550 (I198981,I260275,I260266);
and I_11551 (I198998,I198981,I260278);
DFFARX1 I_11552 (I198998,I2595,I198664,I199024,);
nor I_11553 (I199032,I199024,I198891);
DFFARX1 I_11554 (I199032,I2595,I198664,I198632,);
nand I_11555 (I199063,I199024,I198933);
nand I_11556 (I198641,I198916,I199063);
not I_11557 (I199094,I199024);
nor I_11558 (I199111,I199094,I198834);
DFFARX1 I_11559 (I199111,I2595,I198664,I198653,);
nor I_11560 (I199142,I260263,I260266);
or I_11561 (I198644,I198891,I199142);
nor I_11562 (I198635,I199024,I199142);
or I_11563 (I198638,I198758,I199142);
DFFARX1 I_11564 (I199142,I2595,I198664,I198656,);
not I_11565 (I199242,I2602);
DFFARX1 I_11566 (I68718,I2595,I199242,I199268,);
not I_11567 (I199276,I199268);
nand I_11568 (I199293,I68721,I68742);
and I_11569 (I199310,I199293,I68730);
DFFARX1 I_11570 (I199310,I2595,I199242,I199336,);
not I_11571 (I199344,I68727);
DFFARX1 I_11572 (I68718,I2595,I199242,I199370,);
not I_11573 (I199378,I199370);
nor I_11574 (I199395,I199378,I199276);
and I_11575 (I199412,I199395,I68727);
nor I_11576 (I199429,I199378,I199344);
nor I_11577 (I199225,I199336,I199429);
DFFARX1 I_11578 (I68736,I2595,I199242,I199469,);
nor I_11579 (I199477,I199469,I199336);
not I_11580 (I199494,I199477);
not I_11581 (I199511,I199469);
nor I_11582 (I199528,I199511,I199412);
DFFARX1 I_11583 (I199528,I2595,I199242,I199228,);
nand I_11584 (I199559,I68721,I68724);
and I_11585 (I199576,I199559,I68733);
DFFARX1 I_11586 (I199576,I2595,I199242,I199602,);
nor I_11587 (I199610,I199602,I199469);
DFFARX1 I_11588 (I199610,I2595,I199242,I199210,);
nand I_11589 (I199641,I199602,I199511);
nand I_11590 (I199219,I199494,I199641);
not I_11591 (I199672,I199602);
nor I_11592 (I199689,I199672,I199412);
DFFARX1 I_11593 (I199689,I2595,I199242,I199231,);
nor I_11594 (I199720,I68739,I68724);
or I_11595 (I199222,I199469,I199720);
nor I_11596 (I199213,I199602,I199720);
or I_11597 (I199216,I199336,I199720);
DFFARX1 I_11598 (I199720,I2595,I199242,I199234,);
not I_11599 (I199820,I2602);
DFFARX1 I_11600 (I93290,I2595,I199820,I199846,);
not I_11601 (I199854,I199846);
nand I_11602 (I199871,I93293,I93269);
and I_11603 (I199888,I199871,I93266);
DFFARX1 I_11604 (I199888,I2595,I199820,I199914,);
not I_11605 (I199922,I93272);
DFFARX1 I_11606 (I93266,I2595,I199820,I199948,);
not I_11607 (I199956,I199948);
nor I_11608 (I199973,I199956,I199854);
and I_11609 (I199990,I199973,I93272);
nor I_11610 (I200007,I199956,I199922);
nor I_11611 (I199803,I199914,I200007);
DFFARX1 I_11612 (I93275,I2595,I199820,I200047,);
nor I_11613 (I200055,I200047,I199914);
not I_11614 (I200072,I200055);
not I_11615 (I200089,I200047);
nor I_11616 (I200106,I200089,I199990);
DFFARX1 I_11617 (I200106,I2595,I199820,I199806,);
nand I_11618 (I200137,I93278,I93287);
and I_11619 (I200154,I200137,I93284);
DFFARX1 I_11620 (I200154,I2595,I199820,I200180,);
nor I_11621 (I200188,I200180,I200047);
DFFARX1 I_11622 (I200188,I2595,I199820,I199788,);
nand I_11623 (I200219,I200180,I200089);
nand I_11624 (I199797,I200072,I200219);
not I_11625 (I200250,I200180);
nor I_11626 (I200267,I200250,I199990);
DFFARX1 I_11627 (I200267,I2595,I199820,I199809,);
nor I_11628 (I200298,I93281,I93287);
or I_11629 (I199800,I200047,I200298);
nor I_11630 (I199791,I200180,I200298);
or I_11631 (I199794,I199914,I200298);
DFFARX1 I_11632 (I200298,I2595,I199820,I199812,);
not I_11633 (I200398,I2602);
DFFARX1 I_11634 (I136642,I2595,I200398,I200424,);
not I_11635 (I200432,I200424);
nand I_11636 (I200449,I136633,I136651);
and I_11637 (I200466,I200449,I136654);
DFFARX1 I_11638 (I200466,I2595,I200398,I200492,);
not I_11639 (I200500,I136648);
DFFARX1 I_11640 (I136636,I2595,I200398,I200526,);
not I_11641 (I200534,I200526);
nor I_11642 (I200551,I200534,I200432);
and I_11643 (I200568,I200551,I136648);
nor I_11644 (I200585,I200534,I200500);
nor I_11645 (I200381,I200492,I200585);
DFFARX1 I_11646 (I136645,I2595,I200398,I200625,);
nor I_11647 (I200633,I200625,I200492);
not I_11648 (I200650,I200633);
not I_11649 (I200667,I200625);
nor I_11650 (I200684,I200667,I200568);
DFFARX1 I_11651 (I200684,I2595,I200398,I200384,);
nand I_11652 (I200715,I136660,I136657);
and I_11653 (I200732,I200715,I136639);
DFFARX1 I_11654 (I200732,I2595,I200398,I200758,);
nor I_11655 (I200766,I200758,I200625);
DFFARX1 I_11656 (I200766,I2595,I200398,I200366,);
nand I_11657 (I200797,I200758,I200667);
nand I_11658 (I200375,I200650,I200797);
not I_11659 (I200828,I200758);
nor I_11660 (I200845,I200828,I200568);
DFFARX1 I_11661 (I200845,I2595,I200398,I200387,);
nor I_11662 (I200876,I136633,I136657);
or I_11663 (I200378,I200625,I200876);
nor I_11664 (I200369,I200758,I200876);
or I_11665 (I200372,I200492,I200876);
DFFARX1 I_11666 (I200876,I2595,I200398,I200390,);
not I_11667 (I200976,I2602);
DFFARX1 I_11668 (I66338,I2595,I200976,I201002,);
not I_11669 (I201010,I201002);
nand I_11670 (I201027,I66341,I66362);
and I_11671 (I201044,I201027,I66350);
DFFARX1 I_11672 (I201044,I2595,I200976,I201070,);
not I_11673 (I201078,I66347);
DFFARX1 I_11674 (I66338,I2595,I200976,I201104,);
not I_11675 (I201112,I201104);
nor I_11676 (I201129,I201112,I201010);
and I_11677 (I201146,I201129,I66347);
nor I_11678 (I201163,I201112,I201078);
nor I_11679 (I200959,I201070,I201163);
DFFARX1 I_11680 (I66356,I2595,I200976,I201203,);
nor I_11681 (I201211,I201203,I201070);
not I_11682 (I201228,I201211);
not I_11683 (I201245,I201203);
nor I_11684 (I201262,I201245,I201146);
DFFARX1 I_11685 (I201262,I2595,I200976,I200962,);
nand I_11686 (I201293,I66341,I66344);
and I_11687 (I201310,I201293,I66353);
DFFARX1 I_11688 (I201310,I2595,I200976,I201336,);
nor I_11689 (I201344,I201336,I201203);
DFFARX1 I_11690 (I201344,I2595,I200976,I200944,);
nand I_11691 (I201375,I201336,I201245);
nand I_11692 (I200953,I201228,I201375);
not I_11693 (I201406,I201336);
nor I_11694 (I201423,I201406,I201146);
DFFARX1 I_11695 (I201423,I2595,I200976,I200965,);
nor I_11696 (I201454,I66359,I66344);
or I_11697 (I200956,I201203,I201454);
nor I_11698 (I200947,I201336,I201454);
or I_11699 (I200950,I201070,I201454);
DFFARX1 I_11700 (I201454,I2595,I200976,I200968,);
not I_11701 (I201554,I2602);
DFFARX1 I_11702 (I1940,I2595,I201554,I201580,);
not I_11703 (I201588,I201580);
nand I_11704 (I201605,I2164,I1524);
and I_11705 (I201622,I201605,I2156);
DFFARX1 I_11706 (I201622,I2595,I201554,I201648,);
not I_11707 (I201656,I2004);
DFFARX1 I_11708 (I2100,I2595,I201554,I201682,);
not I_11709 (I201690,I201682);
nor I_11710 (I201707,I201690,I201588);
and I_11711 (I201724,I201707,I2004);
nor I_11712 (I201741,I201690,I201656);
nor I_11713 (I201537,I201648,I201741);
DFFARX1 I_11714 (I2540,I2595,I201554,I201781,);
nor I_11715 (I201789,I201781,I201648);
not I_11716 (I201806,I201789);
not I_11717 (I201823,I201781);
nor I_11718 (I201840,I201823,I201724);
DFFARX1 I_11719 (I201840,I2595,I201554,I201540,);
nand I_11720 (I201871,I2396,I2308);
and I_11721 (I201888,I201871,I2500);
DFFARX1 I_11722 (I201888,I2595,I201554,I201914,);
nor I_11723 (I201922,I201914,I201781);
DFFARX1 I_11724 (I201922,I2595,I201554,I201522,);
nand I_11725 (I201953,I201914,I201823);
nand I_11726 (I201531,I201806,I201953);
not I_11727 (I201984,I201914);
nor I_11728 (I202001,I201984,I201724);
DFFARX1 I_11729 (I202001,I2595,I201554,I201543,);
nor I_11730 (I202032,I1388,I2308);
or I_11731 (I201534,I201781,I202032);
nor I_11732 (I201525,I201914,I202032);
or I_11733 (I201528,I201648,I202032);
DFFARX1 I_11734 (I202032,I2595,I201554,I201546,);
not I_11735 (I202132,I2602);
DFFARX1 I_11736 (I159906,I2595,I202132,I202158,);
not I_11737 (I202166,I202158);
nand I_11738 (I202183,I159915,I159924);
and I_11739 (I202200,I202183,I159930);
DFFARX1 I_11740 (I202200,I2595,I202132,I202226,);
not I_11741 (I202234,I159927);
DFFARX1 I_11742 (I159912,I2595,I202132,I202260,);
not I_11743 (I202268,I202260);
nor I_11744 (I202285,I202268,I202166);
and I_11745 (I202302,I202285,I159927);
nor I_11746 (I202319,I202268,I202234);
nor I_11747 (I202115,I202226,I202319);
DFFARX1 I_11748 (I159921,I2595,I202132,I202359,);
nor I_11749 (I202367,I202359,I202226);
not I_11750 (I202384,I202367);
not I_11751 (I202401,I202359);
nor I_11752 (I202418,I202401,I202302);
DFFARX1 I_11753 (I202418,I2595,I202132,I202118,);
nand I_11754 (I202449,I159918,I159909);
and I_11755 (I202466,I202449,I159906);
DFFARX1 I_11756 (I202466,I2595,I202132,I202492,);
nor I_11757 (I202500,I202492,I202359);
DFFARX1 I_11758 (I202500,I2595,I202132,I202100,);
nand I_11759 (I202531,I202492,I202401);
nand I_11760 (I202109,I202384,I202531);
not I_11761 (I202562,I202492);
nor I_11762 (I202579,I202562,I202302);
DFFARX1 I_11763 (I202579,I2595,I202132,I202121,);
nor I_11764 (I202610,I159909,I159909);
or I_11765 (I202112,I202359,I202610);
nor I_11766 (I202103,I202492,I202610);
or I_11767 (I202106,I202226,I202610);
DFFARX1 I_11768 (I202610,I2595,I202132,I202124,);
not I_11769 (I202710,I2602);
DFFARX1 I_11770 (I117058,I2595,I202710,I202736,);
not I_11771 (I202744,I202736);
nand I_11772 (I202761,I117049,I117067);
and I_11773 (I202778,I202761,I117070);
DFFARX1 I_11774 (I202778,I2595,I202710,I202804,);
not I_11775 (I202812,I117064);
DFFARX1 I_11776 (I117052,I2595,I202710,I202838,);
not I_11777 (I202846,I202838);
nor I_11778 (I202863,I202846,I202744);
and I_11779 (I202880,I202863,I117064);
nor I_11780 (I202897,I202846,I202812);
nor I_11781 (I202693,I202804,I202897);
DFFARX1 I_11782 (I117061,I2595,I202710,I202937,);
nor I_11783 (I202945,I202937,I202804);
not I_11784 (I202962,I202945);
not I_11785 (I202979,I202937);
nor I_11786 (I202996,I202979,I202880);
DFFARX1 I_11787 (I202996,I2595,I202710,I202696,);
nand I_11788 (I203027,I117076,I117073);
and I_11789 (I203044,I203027,I117055);
DFFARX1 I_11790 (I203044,I2595,I202710,I203070,);
nor I_11791 (I203078,I203070,I202937);
DFFARX1 I_11792 (I203078,I2595,I202710,I202678,);
nand I_11793 (I203109,I203070,I202979);
nand I_11794 (I202687,I202962,I203109);
not I_11795 (I203140,I203070);
nor I_11796 (I203157,I203140,I202880);
DFFARX1 I_11797 (I203157,I2595,I202710,I202699,);
nor I_11798 (I203188,I117049,I117073);
or I_11799 (I202690,I202937,I203188);
nor I_11800 (I202681,I203070,I203188);
or I_11801 (I202684,I202804,I203188);
DFFARX1 I_11802 (I203188,I2595,I202710,I202702,);
not I_11803 (I203288,I2602);
DFFARX1 I_11804 (I26085,I2595,I203288,I203314,);
not I_11805 (I203322,I203314);
nand I_11806 (I203339,I26094,I26103);
and I_11807 (I203356,I203339,I26082);
DFFARX1 I_11808 (I203356,I2595,I203288,I203382,);
not I_11809 (I203390,I26085);
DFFARX1 I_11810 (I26100,I2595,I203288,I203416,);
not I_11811 (I203424,I203416);
nor I_11812 (I203441,I203424,I203322);
and I_11813 (I203458,I203441,I26085);
nor I_11814 (I203475,I203424,I203390);
nor I_11815 (I203271,I203382,I203475);
DFFARX1 I_11816 (I26091,I2595,I203288,I203515,);
nor I_11817 (I203523,I203515,I203382);
not I_11818 (I203540,I203523);
not I_11819 (I203557,I203515);
nor I_11820 (I203574,I203557,I203458);
DFFARX1 I_11821 (I203574,I2595,I203288,I203274,);
nand I_11822 (I203605,I26106,I26082);
and I_11823 (I203622,I203605,I26088);
DFFARX1 I_11824 (I203622,I2595,I203288,I203648,);
nor I_11825 (I203656,I203648,I203515);
DFFARX1 I_11826 (I203656,I2595,I203288,I203256,);
nand I_11827 (I203687,I203648,I203557);
nand I_11828 (I203265,I203540,I203687);
not I_11829 (I203718,I203648);
nor I_11830 (I203735,I203718,I203458);
DFFARX1 I_11831 (I203735,I2595,I203288,I203277,);
nor I_11832 (I203766,I26097,I26082);
or I_11833 (I203268,I203515,I203766);
nor I_11834 (I203259,I203648,I203766);
or I_11835 (I203262,I203382,I203766);
DFFARX1 I_11836 (I203766,I2595,I203288,I203280,);
not I_11837 (I203866,I2602);
DFFARX1 I_11838 (I2588,I2595,I203866,I203892,);
not I_11839 (I203900,I203892);
nand I_11840 (I203917,I2172,I1468);
and I_11841 (I203934,I203917,I1540);
DFFARX1 I_11842 (I203934,I2595,I203866,I203960,);
not I_11843 (I203968,I1532);
DFFARX1 I_11844 (I2180,I2595,I203866,I203994,);
not I_11845 (I204002,I203994);
nor I_11846 (I204019,I204002,I203900);
and I_11847 (I204036,I204019,I1532);
nor I_11848 (I204053,I204002,I203968);
nor I_11849 (I203849,I203960,I204053);
DFFARX1 I_11850 (I2340,I2595,I203866,I204093,);
nor I_11851 (I204101,I204093,I203960);
not I_11852 (I204118,I204101);
not I_11853 (I204135,I204093);
nor I_11854 (I204152,I204135,I204036);
DFFARX1 I_11855 (I204152,I2595,I203866,I203852,);
nand I_11856 (I204183,I1564,I1380);
and I_11857 (I204200,I204183,I2076);
DFFARX1 I_11858 (I204200,I2595,I203866,I204226,);
nor I_11859 (I204234,I204226,I204093);
DFFARX1 I_11860 (I204234,I2595,I203866,I203834,);
nand I_11861 (I204265,I204226,I204135);
nand I_11862 (I203843,I204118,I204265);
not I_11863 (I204296,I204226);
nor I_11864 (I204313,I204296,I204036);
DFFARX1 I_11865 (I204313,I2595,I203866,I203855,);
nor I_11866 (I204344,I1676,I1380);
or I_11867 (I203846,I204093,I204344);
nor I_11868 (I203837,I204226,I204344);
or I_11869 (I203840,I203960,I204344);
DFFARX1 I_11870 (I204344,I2595,I203866,I203858,);
not I_11871 (I204444,I2602);
DFFARX1 I_11872 (I125218,I2595,I204444,I204470,);
not I_11873 (I204478,I204470);
nand I_11874 (I204495,I125209,I125227);
and I_11875 (I204512,I204495,I125230);
DFFARX1 I_11876 (I204512,I2595,I204444,I204538,);
not I_11877 (I204546,I125224);
DFFARX1 I_11878 (I125212,I2595,I204444,I204572,);
not I_11879 (I204580,I204572);
nor I_11880 (I204597,I204580,I204478);
and I_11881 (I204614,I204597,I125224);
nor I_11882 (I204631,I204580,I204546);
nor I_11883 (I204427,I204538,I204631);
DFFARX1 I_11884 (I125221,I2595,I204444,I204671,);
nor I_11885 (I204679,I204671,I204538);
not I_11886 (I204696,I204679);
not I_11887 (I204713,I204671);
nor I_11888 (I204730,I204713,I204614);
DFFARX1 I_11889 (I204730,I2595,I204444,I204430,);
nand I_11890 (I204761,I125236,I125233);
and I_11891 (I204778,I204761,I125215);
DFFARX1 I_11892 (I204778,I2595,I204444,I204804,);
nor I_11893 (I204812,I204804,I204671);
DFFARX1 I_11894 (I204812,I2595,I204444,I204412,);
nand I_11895 (I204843,I204804,I204713);
nand I_11896 (I204421,I204696,I204843);
not I_11897 (I204874,I204804);
nor I_11898 (I204891,I204874,I204614);
DFFARX1 I_11899 (I204891,I2595,I204444,I204433,);
nor I_11900 (I204922,I125209,I125233);
or I_11901 (I204424,I204671,I204922);
nor I_11902 (I204415,I204804,I204922);
or I_11903 (I204418,I204538,I204922);
DFFARX1 I_11904 (I204922,I2595,I204444,I204436,);
not I_11905 (I205022,I2602);
DFFARX1 I_11906 (I286767,I2595,I205022,I205048,);
not I_11907 (I205056,I205048);
nand I_11908 (I205073,I286743,I286758);
and I_11909 (I205090,I205073,I286770);
DFFARX1 I_11910 (I205090,I2595,I205022,I205116,);
not I_11911 (I205124,I286755);
DFFARX1 I_11912 (I286746,I2595,I205022,I205150,);
not I_11913 (I205158,I205150);
nor I_11914 (I205175,I205158,I205056);
and I_11915 (I205192,I205175,I286755);
nor I_11916 (I205209,I205158,I205124);
nor I_11917 (I205005,I205116,I205209);
DFFARX1 I_11918 (I286743,I2595,I205022,I205249,);
nor I_11919 (I205257,I205249,I205116);
not I_11920 (I205274,I205257);
not I_11921 (I205291,I205249);
nor I_11922 (I205308,I205291,I205192);
DFFARX1 I_11923 (I205308,I2595,I205022,I205008,);
nand I_11924 (I205339,I286761,I286752);
and I_11925 (I205356,I205339,I286764);
DFFARX1 I_11926 (I205356,I2595,I205022,I205382,);
nor I_11927 (I205390,I205382,I205249);
DFFARX1 I_11928 (I205390,I2595,I205022,I204990,);
nand I_11929 (I205421,I205382,I205291);
nand I_11930 (I204999,I205274,I205421);
not I_11931 (I205452,I205382);
nor I_11932 (I205469,I205452,I205192);
DFFARX1 I_11933 (I205469,I2595,I205022,I205011,);
nor I_11934 (I205500,I286749,I286752);
or I_11935 (I205002,I205249,I205500);
nor I_11936 (I204993,I205382,I205500);
or I_11937 (I204996,I205116,I205500);
DFFARX1 I_11938 (I205500,I2595,I205022,I205014,);
not I_11939 (I205600,I2602);
DFFARX1 I_11940 (I264803,I2595,I205600,I205626,);
not I_11941 (I205634,I205626);
nand I_11942 (I205651,I264779,I264794);
and I_11943 (I205668,I205651,I264806);
DFFARX1 I_11944 (I205668,I2595,I205600,I205694,);
not I_11945 (I205702,I264791);
DFFARX1 I_11946 (I264782,I2595,I205600,I205728,);
not I_11947 (I205736,I205728);
nor I_11948 (I205753,I205736,I205634);
and I_11949 (I205770,I205753,I264791);
nor I_11950 (I205787,I205736,I205702);
nor I_11951 (I205583,I205694,I205787);
DFFARX1 I_11952 (I264779,I2595,I205600,I205827,);
nor I_11953 (I205835,I205827,I205694);
not I_11954 (I205852,I205835);
not I_11955 (I205869,I205827);
nor I_11956 (I205886,I205869,I205770);
DFFARX1 I_11957 (I205886,I2595,I205600,I205586,);
nand I_11958 (I205917,I264797,I264788);
and I_11959 (I205934,I205917,I264800);
DFFARX1 I_11960 (I205934,I2595,I205600,I205960,);
nor I_11961 (I205968,I205960,I205827);
DFFARX1 I_11962 (I205968,I2595,I205600,I205568,);
nand I_11963 (I205999,I205960,I205869);
nand I_11964 (I205577,I205852,I205999);
not I_11965 (I206030,I205960);
nor I_11966 (I206047,I206030,I205770);
DFFARX1 I_11967 (I206047,I2595,I205600,I205589,);
nor I_11968 (I206078,I264785,I264788);
or I_11969 (I205580,I205827,I206078);
nor I_11970 (I205571,I205960,I206078);
or I_11971 (I205574,I205694,I206078);
DFFARX1 I_11972 (I206078,I2595,I205600,I205592,);
not I_11973 (I206178,I2602);
DFFARX1 I_11974 (I20824,I2595,I206178,I206204,);
not I_11975 (I206212,I206204);
nand I_11976 (I206229,I20821,I20812);
and I_11977 (I206246,I206229,I20812);
DFFARX1 I_11978 (I206246,I2595,I206178,I206272,);
not I_11979 (I206280,I20815);
DFFARX1 I_11980 (I20830,I2595,I206178,I206306,);
not I_11981 (I206314,I206306);
nor I_11982 (I206331,I206314,I206212);
and I_11983 (I206348,I206331,I20815);
nor I_11984 (I206365,I206314,I206280);
nor I_11985 (I206161,I206272,I206365);
DFFARX1 I_11986 (I20815,I2595,I206178,I206405,);
nor I_11987 (I206413,I206405,I206272);
not I_11988 (I206430,I206413);
not I_11989 (I206447,I206405);
nor I_11990 (I206464,I206447,I206348);
DFFARX1 I_11991 (I206464,I2595,I206178,I206164,);
nand I_11992 (I206495,I20833,I20818);
and I_11993 (I206512,I206495,I20836);
DFFARX1 I_11994 (I206512,I2595,I206178,I206538,);
nor I_11995 (I206546,I206538,I206405);
DFFARX1 I_11996 (I206546,I2595,I206178,I206146,);
nand I_11997 (I206577,I206538,I206447);
nand I_11998 (I206155,I206430,I206577);
not I_11999 (I206608,I206538);
nor I_12000 (I206625,I206608,I206348);
DFFARX1 I_12001 (I206625,I2595,I206178,I206167,);
nor I_12002 (I206656,I20827,I20818);
or I_12003 (I206158,I206405,I206656);
nor I_12004 (I206149,I206538,I206656);
or I_12005 (I206152,I206272,I206656);
DFFARX1 I_12006 (I206656,I2595,I206178,I206170,);
not I_12007 (I206756,I2602);
DFFARX1 I_12008 (I258989,I2595,I206756,I206782,);
not I_12009 (I206790,I206782);
nand I_12010 (I206807,I258965,I258980);
and I_12011 (I206824,I206807,I258992);
DFFARX1 I_12012 (I206824,I2595,I206756,I206850,);
not I_12013 (I206858,I258977);
DFFARX1 I_12014 (I258968,I2595,I206756,I206884,);
not I_12015 (I206892,I206884);
nor I_12016 (I206909,I206892,I206790);
and I_12017 (I206926,I206909,I258977);
nor I_12018 (I206943,I206892,I206858);
nor I_12019 (I206739,I206850,I206943);
DFFARX1 I_12020 (I258965,I2595,I206756,I206983,);
nor I_12021 (I206991,I206983,I206850);
not I_12022 (I207008,I206991);
not I_12023 (I207025,I206983);
nor I_12024 (I207042,I207025,I206926);
DFFARX1 I_12025 (I207042,I2595,I206756,I206742,);
nand I_12026 (I207073,I258983,I258974);
and I_12027 (I207090,I207073,I258986);
DFFARX1 I_12028 (I207090,I2595,I206756,I207116,);
nor I_12029 (I207124,I207116,I206983);
DFFARX1 I_12030 (I207124,I2595,I206756,I206724,);
nand I_12031 (I207155,I207116,I207025);
nand I_12032 (I206733,I207008,I207155);
not I_12033 (I207186,I207116);
nor I_12034 (I207203,I207186,I206926);
DFFARX1 I_12035 (I207203,I2595,I206756,I206745,);
nor I_12036 (I207234,I258971,I258974);
or I_12037 (I206736,I206983,I207234);
nor I_12038 (I206727,I207116,I207234);
or I_12039 (I206730,I206850,I207234);
DFFARX1 I_12040 (I207234,I2595,I206756,I206748,);
not I_12041 (I207334,I2602);
DFFARX1 I_12042 (I333936,I2595,I207334,I207360,);
not I_12043 (I207368,I207360);
nand I_12044 (I207385,I333918,I333930);
and I_12045 (I207402,I207385,I333933);
DFFARX1 I_12046 (I207402,I2595,I207334,I207428,);
not I_12047 (I207436,I333927);
DFFARX1 I_12048 (I333924,I2595,I207334,I207462,);
not I_12049 (I207470,I207462);
nor I_12050 (I207487,I207470,I207368);
and I_12051 (I207504,I207487,I333927);
nor I_12052 (I207521,I207470,I207436);
nor I_12053 (I207317,I207428,I207521);
DFFARX1 I_12054 (I333942,I2595,I207334,I207561,);
nor I_12055 (I207569,I207561,I207428);
not I_12056 (I207586,I207569);
not I_12057 (I207603,I207561);
nor I_12058 (I207620,I207603,I207504);
DFFARX1 I_12059 (I207620,I2595,I207334,I207320,);
nand I_12060 (I207651,I333921,I333921);
and I_12061 (I207668,I207651,I333918);
DFFARX1 I_12062 (I207668,I2595,I207334,I207694,);
nor I_12063 (I207702,I207694,I207561);
DFFARX1 I_12064 (I207702,I2595,I207334,I207302,);
nand I_12065 (I207733,I207694,I207603);
nand I_12066 (I207311,I207586,I207733);
not I_12067 (I207764,I207694);
nor I_12068 (I207781,I207764,I207504);
DFFARX1 I_12069 (I207781,I2595,I207334,I207323,);
nor I_12070 (I207812,I333939,I333921);
or I_12071 (I207314,I207561,I207812);
nor I_12072 (I207305,I207694,I207812);
or I_12073 (I207308,I207428,I207812);
DFFARX1 I_12074 (I207812,I2595,I207334,I207326,);
not I_12075 (I207912,I2602);
DFFARX1 I_12076 (I279661,I2595,I207912,I207938,);
not I_12077 (I207946,I207938);
nand I_12078 (I207963,I279637,I279652);
and I_12079 (I207980,I207963,I279664);
DFFARX1 I_12080 (I207980,I2595,I207912,I208006,);
not I_12081 (I208014,I279649);
DFFARX1 I_12082 (I279640,I2595,I207912,I208040,);
not I_12083 (I208048,I208040);
nor I_12084 (I208065,I208048,I207946);
and I_12085 (I208082,I208065,I279649);
nor I_12086 (I208099,I208048,I208014);
nor I_12087 (I207895,I208006,I208099);
DFFARX1 I_12088 (I279637,I2595,I207912,I208139,);
nor I_12089 (I208147,I208139,I208006);
not I_12090 (I208164,I208147);
not I_12091 (I208181,I208139);
nor I_12092 (I208198,I208181,I208082);
DFFARX1 I_12093 (I208198,I2595,I207912,I207898,);
nand I_12094 (I208229,I279655,I279646);
and I_12095 (I208246,I208229,I279658);
DFFARX1 I_12096 (I208246,I2595,I207912,I208272,);
nor I_12097 (I208280,I208272,I208139);
DFFARX1 I_12098 (I208280,I2595,I207912,I207880,);
nand I_12099 (I208311,I208272,I208181);
nand I_12100 (I207889,I208164,I208311);
not I_12101 (I208342,I208272);
nor I_12102 (I208359,I208342,I208082);
DFFARX1 I_12103 (I208359,I2595,I207912,I207901,);
nor I_12104 (I208390,I279643,I279646);
or I_12105 (I207892,I208139,I208390);
nor I_12106 (I207883,I208272,I208390);
or I_12107 (I207886,I208006,I208390);
DFFARX1 I_12108 (I208390,I2595,I207912,I207904,);
not I_12109 (I208490,I2602);
DFFARX1 I_12110 (I342028,I2595,I208490,I208516,);
not I_12111 (I208524,I208516);
nand I_12112 (I208541,I342010,I342022);
and I_12113 (I208558,I208541,I342025);
DFFARX1 I_12114 (I208558,I2595,I208490,I208584,);
not I_12115 (I208592,I342019);
DFFARX1 I_12116 (I342016,I2595,I208490,I208618,);
not I_12117 (I208626,I208618);
nor I_12118 (I208643,I208626,I208524);
and I_12119 (I208660,I208643,I342019);
nor I_12120 (I208677,I208626,I208592);
nor I_12121 (I208473,I208584,I208677);
DFFARX1 I_12122 (I342034,I2595,I208490,I208717,);
nor I_12123 (I208725,I208717,I208584);
not I_12124 (I208742,I208725);
not I_12125 (I208759,I208717);
nor I_12126 (I208776,I208759,I208660);
DFFARX1 I_12127 (I208776,I2595,I208490,I208476,);
nand I_12128 (I208807,I342013,I342013);
and I_12129 (I208824,I208807,I342010);
DFFARX1 I_12130 (I208824,I2595,I208490,I208850,);
nor I_12131 (I208858,I208850,I208717);
DFFARX1 I_12132 (I208858,I2595,I208490,I208458,);
nand I_12133 (I208889,I208850,I208759);
nand I_12134 (I208467,I208742,I208889);
not I_12135 (I208920,I208850);
nor I_12136 (I208937,I208920,I208660);
DFFARX1 I_12137 (I208937,I2595,I208490,I208479,);
nor I_12138 (I208968,I342031,I342013);
or I_12139 (I208470,I208717,I208968);
nor I_12140 (I208461,I208850,I208968);
or I_12141 (I208464,I208584,I208968);
DFFARX1 I_12142 (I208968,I2595,I208490,I208482,);
not I_12143 (I209068,I2602);
DFFARX1 I_12144 (I150505,I2595,I209068,I209094,);
not I_12145 (I209102,I209094);
nand I_12146 (I209119,I150520,I150505);
and I_12147 (I209136,I209119,I150508);
DFFARX1 I_12148 (I209136,I2595,I209068,I209162,);
not I_12149 (I209170,I150508);
DFFARX1 I_12150 (I150517,I2595,I209068,I209196,);
not I_12151 (I209204,I209196);
nor I_12152 (I209221,I209204,I209102);
and I_12153 (I209238,I209221,I150508);
nor I_12154 (I209255,I209204,I209170);
nor I_12155 (I209051,I209162,I209255);
DFFARX1 I_12156 (I150511,I2595,I209068,I209295,);
nor I_12157 (I209303,I209295,I209162);
not I_12158 (I209320,I209303);
not I_12159 (I209337,I209295);
nor I_12160 (I209354,I209337,I209238);
DFFARX1 I_12161 (I209354,I2595,I209068,I209054,);
nand I_12162 (I209385,I150514,I150523);
and I_12163 (I209402,I209385,I150529);
DFFARX1 I_12164 (I209402,I2595,I209068,I209428,);
nor I_12165 (I209436,I209428,I209295);
DFFARX1 I_12166 (I209436,I2595,I209068,I209036,);
nand I_12167 (I209467,I209428,I209337);
nand I_12168 (I209045,I209320,I209467);
not I_12169 (I209498,I209428);
nor I_12170 (I209515,I209498,I209238);
DFFARX1 I_12171 (I209515,I2595,I209068,I209057,);
nor I_12172 (I209546,I150526,I150523);
or I_12173 (I209048,I209295,I209546);
nor I_12174 (I209039,I209428,I209546);
or I_12175 (I209042,I209162,I209546);
DFFARX1 I_12176 (I209546,I2595,I209068,I209060,);
not I_12177 (I209646,I2602);
DFFARX1 I_12178 (I317174,I2595,I209646,I209672,);
not I_12179 (I209680,I209672);
nand I_12180 (I209697,I317156,I317168);
and I_12181 (I209714,I209697,I317171);
DFFARX1 I_12182 (I209714,I2595,I209646,I209740,);
not I_12183 (I209748,I317165);
DFFARX1 I_12184 (I317162,I2595,I209646,I209774,);
not I_12185 (I209782,I209774);
nor I_12186 (I209799,I209782,I209680);
and I_12187 (I209816,I209799,I317165);
nor I_12188 (I209833,I209782,I209748);
nor I_12189 (I209629,I209740,I209833);
DFFARX1 I_12190 (I317180,I2595,I209646,I209873,);
nor I_12191 (I209881,I209873,I209740);
not I_12192 (I209898,I209881);
not I_12193 (I209915,I209873);
nor I_12194 (I209932,I209915,I209816);
DFFARX1 I_12195 (I209932,I2595,I209646,I209632,);
nand I_12196 (I209963,I317159,I317159);
and I_12197 (I209980,I209963,I317156);
DFFARX1 I_12198 (I209980,I2595,I209646,I210006,);
nor I_12199 (I210014,I210006,I209873);
DFFARX1 I_12200 (I210014,I2595,I209646,I209614,);
nand I_12201 (I210045,I210006,I209915);
nand I_12202 (I209623,I209898,I210045);
not I_12203 (I210076,I210006);
nor I_12204 (I210093,I210076,I209816);
DFFARX1 I_12205 (I210093,I2595,I209646,I209635,);
nor I_12206 (I210124,I317177,I317159);
or I_12207 (I209626,I209873,I210124);
nor I_12208 (I209617,I210006,I210124);
or I_12209 (I209620,I209740,I210124);
DFFARX1 I_12210 (I210124,I2595,I209646,I209638,);
not I_12211 (I210224,I2602);
DFFARX1 I_12212 (I170888,I2595,I210224,I210250,);
not I_12213 (I210258,I210250);
nand I_12214 (I210275,I170897,I170906);
and I_12215 (I210292,I210275,I170912);
DFFARX1 I_12216 (I210292,I2595,I210224,I210318,);
not I_12217 (I210326,I170909);
DFFARX1 I_12218 (I170894,I2595,I210224,I210352,);
not I_12219 (I210360,I210352);
nor I_12220 (I210377,I210360,I210258);
and I_12221 (I210394,I210377,I170909);
nor I_12222 (I210411,I210360,I210326);
nor I_12223 (I210207,I210318,I210411);
DFFARX1 I_12224 (I170903,I2595,I210224,I210451,);
nor I_12225 (I210459,I210451,I210318);
not I_12226 (I210476,I210459);
not I_12227 (I210493,I210451);
nor I_12228 (I210510,I210493,I210394);
DFFARX1 I_12229 (I210510,I2595,I210224,I210210,);
nand I_12230 (I210541,I170900,I170891);
and I_12231 (I210558,I210541,I170888);
DFFARX1 I_12232 (I210558,I2595,I210224,I210584,);
nor I_12233 (I210592,I210584,I210451);
DFFARX1 I_12234 (I210592,I2595,I210224,I210192,);
nand I_12235 (I210623,I210584,I210493);
nand I_12236 (I210201,I210476,I210623);
not I_12237 (I210654,I210584);
nor I_12238 (I210671,I210654,I210394);
DFFARX1 I_12239 (I210671,I2595,I210224,I210213,);
nor I_12240 (I210702,I170891,I170891);
or I_12241 (I210204,I210451,I210702);
nor I_12242 (I210195,I210584,I210702);
or I_12243 (I210198,I210318,I210702);
DFFARX1 I_12244 (I210702,I2595,I210224,I210216,);
not I_12245 (I210802,I2602);
DFFARX1 I_12246 (I275139,I2595,I210802,I210828,);
not I_12247 (I210836,I210828);
nand I_12248 (I210853,I275115,I275130);
and I_12249 (I210870,I210853,I275142);
DFFARX1 I_12250 (I210870,I2595,I210802,I210896,);
not I_12251 (I210904,I275127);
DFFARX1 I_12252 (I275118,I2595,I210802,I210930,);
not I_12253 (I210938,I210930);
nor I_12254 (I210955,I210938,I210836);
and I_12255 (I210972,I210955,I275127);
nor I_12256 (I210989,I210938,I210904);
nor I_12257 (I210785,I210896,I210989);
DFFARX1 I_12258 (I275115,I2595,I210802,I211029,);
nor I_12259 (I211037,I211029,I210896);
not I_12260 (I211054,I211037);
not I_12261 (I211071,I211029);
nor I_12262 (I211088,I211071,I210972);
DFFARX1 I_12263 (I211088,I2595,I210802,I210788,);
nand I_12264 (I211119,I275133,I275124);
and I_12265 (I211136,I211119,I275136);
DFFARX1 I_12266 (I211136,I2595,I210802,I211162,);
nor I_12267 (I211170,I211162,I211029);
DFFARX1 I_12268 (I211170,I2595,I210802,I210770,);
nand I_12269 (I211201,I211162,I211071);
nand I_12270 (I210779,I211054,I211201);
not I_12271 (I211232,I211162);
nor I_12272 (I211249,I211232,I210972);
DFFARX1 I_12273 (I211249,I2595,I210802,I210791,);
nor I_12274 (I211280,I275121,I275124);
or I_12275 (I210782,I211029,I211280);
nor I_12276 (I210773,I211162,I211280);
or I_12277 (I210776,I210896,I211280);
DFFARX1 I_12278 (I211280,I2595,I210802,I210794,);
not I_12279 (I211380,I2602);
DFFARX1 I_12280 (I104884,I2595,I211380,I211406,);
not I_12281 (I211414,I211406);
nand I_12282 (I211431,I104887,I104863);
and I_12283 (I211448,I211431,I104860);
DFFARX1 I_12284 (I211448,I2595,I211380,I211474,);
not I_12285 (I211482,I104866);
DFFARX1 I_12286 (I104860,I2595,I211380,I211508,);
not I_12287 (I211516,I211508);
nor I_12288 (I211533,I211516,I211414);
and I_12289 (I211550,I211533,I104866);
nor I_12290 (I211567,I211516,I211482);
nor I_12291 (I211363,I211474,I211567);
DFFARX1 I_12292 (I104869,I2595,I211380,I211607,);
nor I_12293 (I211615,I211607,I211474);
not I_12294 (I211632,I211615);
not I_12295 (I211649,I211607);
nor I_12296 (I211666,I211649,I211550);
DFFARX1 I_12297 (I211666,I2595,I211380,I211366,);
nand I_12298 (I211697,I104872,I104881);
and I_12299 (I211714,I211697,I104878);
DFFARX1 I_12300 (I211714,I2595,I211380,I211740,);
nor I_12301 (I211748,I211740,I211607);
DFFARX1 I_12302 (I211748,I2595,I211380,I211348,);
nand I_12303 (I211779,I211740,I211649);
nand I_12304 (I211357,I211632,I211779);
not I_12305 (I211810,I211740);
nor I_12306 (I211827,I211810,I211550);
DFFARX1 I_12307 (I211827,I2595,I211380,I211369,);
nor I_12308 (I211858,I104875,I104881);
or I_12309 (I211360,I211607,I211858);
nor I_12310 (I211351,I211740,I211858);
or I_12311 (I211354,I211474,I211858);
DFFARX1 I_12312 (I211858,I2595,I211380,I211372,);
not I_12313 (I211958,I2602);
DFFARX1 I_12314 (I40841,I2595,I211958,I211984,);
not I_12315 (I211992,I211984);
nand I_12316 (I212009,I40850,I40859);
and I_12317 (I212026,I212009,I40838);
DFFARX1 I_12318 (I212026,I2595,I211958,I212052,);
not I_12319 (I212060,I40841);
DFFARX1 I_12320 (I40856,I2595,I211958,I212086,);
not I_12321 (I212094,I212086);
nor I_12322 (I212111,I212094,I211992);
and I_12323 (I212128,I212111,I40841);
nor I_12324 (I212145,I212094,I212060);
nor I_12325 (I211941,I212052,I212145);
DFFARX1 I_12326 (I40847,I2595,I211958,I212185,);
nor I_12327 (I212193,I212185,I212052);
not I_12328 (I212210,I212193);
not I_12329 (I212227,I212185);
nor I_12330 (I212244,I212227,I212128);
DFFARX1 I_12331 (I212244,I2595,I211958,I211944,);
nand I_12332 (I212275,I40862,I40838);
and I_12333 (I212292,I212275,I40844);
DFFARX1 I_12334 (I212292,I2595,I211958,I212318,);
nor I_12335 (I212326,I212318,I212185);
DFFARX1 I_12336 (I212326,I2595,I211958,I211926,);
nand I_12337 (I212357,I212318,I212227);
nand I_12338 (I211935,I212210,I212357);
not I_12339 (I212388,I212318);
nor I_12340 (I212405,I212388,I212128);
DFFARX1 I_12341 (I212405,I2595,I211958,I211947,);
nor I_12342 (I212436,I40853,I40838);
or I_12343 (I211938,I212185,I212436);
nor I_12344 (I211929,I212318,I212436);
or I_12345 (I211932,I212052,I212436);
DFFARX1 I_12346 (I212436,I2595,I211958,I211950,);
not I_12347 (I212536,I2602);
DFFARX1 I_12348 (I247250,I2595,I212536,I212562,);
not I_12349 (I212570,I212562);
nand I_12350 (I212587,I247238,I247256);
and I_12351 (I212604,I212587,I247253);
DFFARX1 I_12352 (I212604,I2595,I212536,I212630,);
not I_12353 (I212638,I247244);
DFFARX1 I_12354 (I247241,I2595,I212536,I212664,);
not I_12355 (I212672,I212664);
nor I_12356 (I212689,I212672,I212570);
and I_12357 (I212706,I212689,I247244);
nor I_12358 (I212723,I212672,I212638);
nor I_12359 (I212519,I212630,I212723);
DFFARX1 I_12360 (I247235,I2595,I212536,I212763,);
nor I_12361 (I212771,I212763,I212630);
not I_12362 (I212788,I212771);
not I_12363 (I212805,I212763);
nor I_12364 (I212822,I212805,I212706);
DFFARX1 I_12365 (I212822,I2595,I212536,I212522,);
nand I_12366 (I212853,I247235,I247238);
and I_12367 (I212870,I212853,I247241);
DFFARX1 I_12368 (I212870,I2595,I212536,I212896,);
nor I_12369 (I212904,I212896,I212763);
DFFARX1 I_12370 (I212904,I2595,I212536,I212504,);
nand I_12371 (I212935,I212896,I212805);
nand I_12372 (I212513,I212788,I212935);
not I_12373 (I212966,I212896);
nor I_12374 (I212983,I212966,I212706);
DFFARX1 I_12375 (I212983,I2595,I212536,I212525,);
nor I_12376 (I213014,I247247,I247238);
or I_12377 (I212516,I212763,I213014);
nor I_12378 (I212507,I212896,I213014);
or I_12379 (I212510,I212630,I213014);
DFFARX1 I_12380 (I213014,I2595,I212536,I212528,);
not I_12381 (I213114,I2602);
DFFARX1 I_12382 (I259635,I2595,I213114,I213140,);
not I_12383 (I213148,I213140);
nand I_12384 (I213165,I259611,I259626);
and I_12385 (I213182,I213165,I259638);
DFFARX1 I_12386 (I213182,I2595,I213114,I213208,);
not I_12387 (I213216,I259623);
DFFARX1 I_12388 (I259614,I2595,I213114,I213242,);
not I_12389 (I213250,I213242);
nor I_12390 (I213267,I213250,I213148);
and I_12391 (I213284,I213267,I259623);
nor I_12392 (I213301,I213250,I213216);
nor I_12393 (I213097,I213208,I213301);
DFFARX1 I_12394 (I259611,I2595,I213114,I213341,);
nor I_12395 (I213349,I213341,I213208);
not I_12396 (I213366,I213349);
not I_12397 (I213383,I213341);
nor I_12398 (I213400,I213383,I213284);
DFFARX1 I_12399 (I213400,I2595,I213114,I213100,);
nand I_12400 (I213431,I259629,I259620);
and I_12401 (I213448,I213431,I259632);
DFFARX1 I_12402 (I213448,I2595,I213114,I213474,);
nor I_12403 (I213482,I213474,I213341);
DFFARX1 I_12404 (I213482,I2595,I213114,I213082,);
nand I_12405 (I213513,I213474,I213383);
nand I_12406 (I213091,I213366,I213513);
not I_12407 (I213544,I213474);
nor I_12408 (I213561,I213544,I213284);
DFFARX1 I_12409 (I213561,I2595,I213114,I213103,);
nor I_12410 (I213592,I259617,I259620);
or I_12411 (I213094,I213341,I213592);
nor I_12412 (I213085,I213474,I213592);
or I_12413 (I213088,I213208,I213592);
DFFARX1 I_12414 (I213592,I2595,I213114,I213106,);
not I_12415 (I213692,I2602);
DFFARX1 I_12416 (I101195,I2595,I213692,I213718,);
not I_12417 (I213726,I213718);
nand I_12418 (I213743,I101198,I101174);
and I_12419 (I213760,I213743,I101171);
DFFARX1 I_12420 (I213760,I2595,I213692,I213786,);
not I_12421 (I213794,I101177);
DFFARX1 I_12422 (I101171,I2595,I213692,I213820,);
not I_12423 (I213828,I213820);
nor I_12424 (I213845,I213828,I213726);
and I_12425 (I213862,I213845,I101177);
nor I_12426 (I213879,I213828,I213794);
nor I_12427 (I213675,I213786,I213879);
DFFARX1 I_12428 (I101180,I2595,I213692,I213919,);
nor I_12429 (I213927,I213919,I213786);
not I_12430 (I213944,I213927);
not I_12431 (I213961,I213919);
nor I_12432 (I213978,I213961,I213862);
DFFARX1 I_12433 (I213978,I2595,I213692,I213678,);
nand I_12434 (I214009,I101183,I101192);
and I_12435 (I214026,I214009,I101189);
DFFARX1 I_12436 (I214026,I2595,I213692,I214052,);
nor I_12437 (I214060,I214052,I213919);
DFFARX1 I_12438 (I214060,I2595,I213692,I213660,);
nand I_12439 (I214091,I214052,I213961);
nand I_12440 (I213669,I213944,I214091);
not I_12441 (I214122,I214052);
nor I_12442 (I214139,I214122,I213862);
DFFARX1 I_12443 (I214139,I2595,I213692,I213681,);
nor I_12444 (I214170,I101186,I101192);
or I_12445 (I213672,I213919,I214170);
nor I_12446 (I213663,I214052,I214170);
or I_12447 (I213666,I213786,I214170);
DFFARX1 I_12448 (I214170,I2595,I213692,I213684,);
not I_12449 (I214270,I2602);
DFFARX1 I_12450 (I79428,I2595,I214270,I214296,);
not I_12451 (I214304,I214296);
nand I_12452 (I214321,I79431,I79452);
and I_12453 (I214338,I214321,I79440);
DFFARX1 I_12454 (I214338,I2595,I214270,I214364,);
not I_12455 (I214372,I79437);
DFFARX1 I_12456 (I79428,I2595,I214270,I214398,);
not I_12457 (I214406,I214398);
nor I_12458 (I214423,I214406,I214304);
and I_12459 (I214440,I214423,I79437);
nor I_12460 (I214457,I214406,I214372);
nor I_12461 (I214253,I214364,I214457);
DFFARX1 I_12462 (I79446,I2595,I214270,I214497,);
nor I_12463 (I214505,I214497,I214364);
not I_12464 (I214522,I214505);
not I_12465 (I214539,I214497);
nor I_12466 (I214556,I214539,I214440);
DFFARX1 I_12467 (I214556,I2595,I214270,I214256,);
nand I_12468 (I214587,I79431,I79434);
and I_12469 (I214604,I214587,I79443);
DFFARX1 I_12470 (I214604,I2595,I214270,I214630,);
nor I_12471 (I214638,I214630,I214497);
DFFARX1 I_12472 (I214638,I2595,I214270,I214238,);
nand I_12473 (I214669,I214630,I214539);
nand I_12474 (I214247,I214522,I214669);
not I_12475 (I214700,I214630);
nor I_12476 (I214717,I214700,I214440);
DFFARX1 I_12477 (I214717,I2595,I214270,I214259,);
nor I_12478 (I214748,I79449,I79434);
or I_12479 (I214250,I214497,I214748);
nor I_12480 (I214241,I214630,I214748);
or I_12481 (I214244,I214364,I214748);
DFFARX1 I_12482 (I214748,I2595,I214270,I214262,);
not I_12483 (I214848,I2602);
DFFARX1 I_12484 (I380100,I2595,I214848,I214874,);
not I_12485 (I214882,I214874);
nand I_12486 (I214899,I380085,I380073);
and I_12487 (I214916,I214899,I380088);
DFFARX1 I_12488 (I214916,I2595,I214848,I214942,);
not I_12489 (I214950,I380073);
DFFARX1 I_12490 (I380091,I2595,I214848,I214976,);
not I_12491 (I214984,I214976);
nor I_12492 (I215001,I214984,I214882);
and I_12493 (I215018,I215001,I380073);
nor I_12494 (I215035,I214984,I214950);
nor I_12495 (I214831,I214942,I215035);
DFFARX1 I_12496 (I380079,I2595,I214848,I215075,);
nor I_12497 (I215083,I215075,I214942);
not I_12498 (I215100,I215083);
not I_12499 (I215117,I215075);
nor I_12500 (I215134,I215117,I215018);
DFFARX1 I_12501 (I215134,I2595,I214848,I214834,);
nand I_12502 (I215165,I380076,I380082);
and I_12503 (I215182,I215165,I380097);
DFFARX1 I_12504 (I215182,I2595,I214848,I215208,);
nor I_12505 (I215216,I215208,I215075);
DFFARX1 I_12506 (I215216,I2595,I214848,I214816,);
nand I_12507 (I215247,I215208,I215117);
nand I_12508 (I214825,I215100,I215247);
not I_12509 (I215278,I215208);
nor I_12510 (I215295,I215278,I215018);
DFFARX1 I_12511 (I215295,I2595,I214848,I214837,);
nor I_12512 (I215326,I380094,I380082);
or I_12513 (I214828,I215075,I215326);
nor I_12514 (I214819,I215208,I215326);
or I_12515 (I214822,I214942,I215326);
DFFARX1 I_12516 (I215326,I2595,I214848,I214840,);
not I_12517 (I215426,I2602);
DFFARX1 I_12518 (I119234,I2595,I215426,I215452,);
not I_12519 (I215460,I215452);
nand I_12520 (I215477,I119225,I119243);
and I_12521 (I215494,I215477,I119246);
DFFARX1 I_12522 (I215494,I2595,I215426,I215520,);
not I_12523 (I215528,I119240);
DFFARX1 I_12524 (I119228,I2595,I215426,I215554,);
not I_12525 (I215562,I215554);
nor I_12526 (I215579,I215562,I215460);
and I_12527 (I215596,I215579,I119240);
nor I_12528 (I215613,I215562,I215528);
nor I_12529 (I215409,I215520,I215613);
DFFARX1 I_12530 (I119237,I2595,I215426,I215653,);
nor I_12531 (I215661,I215653,I215520);
not I_12532 (I215678,I215661);
not I_12533 (I215695,I215653);
nor I_12534 (I215712,I215695,I215596);
DFFARX1 I_12535 (I215712,I2595,I215426,I215412,);
nand I_12536 (I215743,I119252,I119249);
and I_12537 (I215760,I215743,I119231);
DFFARX1 I_12538 (I215760,I2595,I215426,I215786,);
nor I_12539 (I215794,I215786,I215653);
DFFARX1 I_12540 (I215794,I2595,I215426,I215394,);
nand I_12541 (I215825,I215786,I215695);
nand I_12542 (I215403,I215678,I215825);
not I_12543 (I215856,I215786);
nor I_12544 (I215873,I215856,I215596);
DFFARX1 I_12545 (I215873,I2595,I215426,I215415,);
nor I_12546 (I215904,I119225,I119249);
or I_12547 (I215406,I215653,I215904);
nor I_12548 (I215397,I215786,I215904);
or I_12549 (I215400,I215520,I215904);
DFFARX1 I_12550 (I215904,I2595,I215426,I215418,);
not I_12551 (I216004,I2602);
DFFARX1 I_12552 (I29774,I2595,I216004,I216030,);
not I_12553 (I216038,I216030);
nand I_12554 (I216055,I29783,I29792);
and I_12555 (I216072,I216055,I29771);
DFFARX1 I_12556 (I216072,I2595,I216004,I216098,);
not I_12557 (I216106,I29774);
DFFARX1 I_12558 (I29789,I2595,I216004,I216132,);
not I_12559 (I216140,I216132);
nor I_12560 (I216157,I216140,I216038);
and I_12561 (I216174,I216157,I29774);
nor I_12562 (I216191,I216140,I216106);
nor I_12563 (I215987,I216098,I216191);
DFFARX1 I_12564 (I29780,I2595,I216004,I216231,);
nor I_12565 (I216239,I216231,I216098);
not I_12566 (I216256,I216239);
not I_12567 (I216273,I216231);
nor I_12568 (I216290,I216273,I216174);
DFFARX1 I_12569 (I216290,I2595,I216004,I215990,);
nand I_12570 (I216321,I29795,I29771);
and I_12571 (I216338,I216321,I29777);
DFFARX1 I_12572 (I216338,I2595,I216004,I216364,);
nor I_12573 (I216372,I216364,I216231);
DFFARX1 I_12574 (I216372,I2595,I216004,I215972,);
nand I_12575 (I216403,I216364,I216273);
nand I_12576 (I215981,I216256,I216403);
not I_12577 (I216434,I216364);
nor I_12578 (I216451,I216434,I216174);
DFFARX1 I_12579 (I216451,I2595,I216004,I215993,);
nor I_12580 (I216482,I29786,I29771);
or I_12581 (I215984,I216231,I216482);
nor I_12582 (I215975,I216364,I216482);
or I_12583 (I215978,I216098,I216482);
DFFARX1 I_12584 (I216482,I2595,I216004,I215996,);
not I_12585 (I216582,I2602);
DFFARX1 I_12586 (I28193,I2595,I216582,I216608,);
not I_12587 (I216616,I216608);
nand I_12588 (I216633,I28202,I28211);
and I_12589 (I216650,I216633,I28190);
DFFARX1 I_12590 (I216650,I2595,I216582,I216676,);
not I_12591 (I216684,I28193);
DFFARX1 I_12592 (I28208,I2595,I216582,I216710,);
not I_12593 (I216718,I216710);
nor I_12594 (I216735,I216718,I216616);
and I_12595 (I216752,I216735,I28193);
nor I_12596 (I216769,I216718,I216684);
nor I_12597 (I216565,I216676,I216769);
DFFARX1 I_12598 (I28199,I2595,I216582,I216809,);
nor I_12599 (I216817,I216809,I216676);
not I_12600 (I216834,I216817);
not I_12601 (I216851,I216809);
nor I_12602 (I216868,I216851,I216752);
DFFARX1 I_12603 (I216868,I2595,I216582,I216568,);
nand I_12604 (I216899,I28214,I28190);
and I_12605 (I216916,I216899,I28196);
DFFARX1 I_12606 (I216916,I2595,I216582,I216942,);
nor I_12607 (I216950,I216942,I216809);
DFFARX1 I_12608 (I216950,I2595,I216582,I216550,);
nand I_12609 (I216981,I216942,I216851);
nand I_12610 (I216559,I216834,I216981);
not I_12611 (I217012,I216942);
nor I_12612 (I217029,I217012,I216752);
DFFARX1 I_12613 (I217029,I2595,I216582,I216571,);
nor I_12614 (I217060,I28205,I28190);
or I_12615 (I216562,I216809,I217060);
nor I_12616 (I216553,I216942,I217060);
or I_12617 (I216556,I216676,I217060);
DFFARX1 I_12618 (I217060,I2595,I216582,I216574,);
not I_12619 (I217160,I2602);
DFFARX1 I_12620 (I253175,I2595,I217160,I217186,);
not I_12621 (I217194,I217186);
nand I_12622 (I217211,I253151,I253166);
and I_12623 (I217228,I217211,I253178);
DFFARX1 I_12624 (I217228,I2595,I217160,I217254,);
not I_12625 (I217262,I253163);
DFFARX1 I_12626 (I253154,I2595,I217160,I217288,);
not I_12627 (I217296,I217288);
nor I_12628 (I217313,I217296,I217194);
and I_12629 (I217330,I217313,I253163);
nor I_12630 (I217347,I217296,I217262);
nor I_12631 (I217143,I217254,I217347);
DFFARX1 I_12632 (I253151,I2595,I217160,I217387,);
nor I_12633 (I217395,I217387,I217254);
not I_12634 (I217412,I217395);
not I_12635 (I217429,I217387);
nor I_12636 (I217446,I217429,I217330);
DFFARX1 I_12637 (I217446,I2595,I217160,I217146,);
nand I_12638 (I217477,I253169,I253160);
and I_12639 (I217494,I217477,I253172);
DFFARX1 I_12640 (I217494,I2595,I217160,I217520,);
nor I_12641 (I217528,I217520,I217387);
DFFARX1 I_12642 (I217528,I2595,I217160,I217128,);
nand I_12643 (I217559,I217520,I217429);
nand I_12644 (I217137,I217412,I217559);
not I_12645 (I217590,I217520);
nor I_12646 (I217607,I217590,I217330);
DFFARX1 I_12647 (I217607,I2595,I217160,I217149,);
nor I_12648 (I217638,I253157,I253160);
or I_12649 (I217140,I217387,I217638);
nor I_12650 (I217131,I217520,I217638);
or I_12651 (I217134,I217254,I217638);
DFFARX1 I_12652 (I217638,I2595,I217160,I217152,);
not I_12653 (I217738,I2602);
DFFARX1 I_12654 (I377720,I2595,I217738,I217764,);
not I_12655 (I217772,I217764);
nand I_12656 (I217789,I377705,I377693);
and I_12657 (I217806,I217789,I377708);
DFFARX1 I_12658 (I217806,I2595,I217738,I217832,);
not I_12659 (I217840,I377693);
DFFARX1 I_12660 (I377711,I2595,I217738,I217866,);
not I_12661 (I217874,I217866);
nor I_12662 (I217891,I217874,I217772);
and I_12663 (I217908,I217891,I377693);
nor I_12664 (I217925,I217874,I217840);
nor I_12665 (I217721,I217832,I217925);
DFFARX1 I_12666 (I377699,I2595,I217738,I217965,);
nor I_12667 (I217973,I217965,I217832);
not I_12668 (I217990,I217973);
not I_12669 (I218007,I217965);
nor I_12670 (I218024,I218007,I217908);
DFFARX1 I_12671 (I218024,I2595,I217738,I217724,);
nand I_12672 (I218055,I377696,I377702);
and I_12673 (I218072,I218055,I377717);
DFFARX1 I_12674 (I218072,I2595,I217738,I218098,);
nor I_12675 (I218106,I218098,I217965);
DFFARX1 I_12676 (I218106,I2595,I217738,I217706,);
nand I_12677 (I218137,I218098,I218007);
nand I_12678 (I217715,I217990,I218137);
not I_12679 (I218168,I218098);
nor I_12680 (I218185,I218168,I217908);
DFFARX1 I_12681 (I218185,I2595,I217738,I217727,);
nor I_12682 (I218216,I377714,I377702);
or I_12683 (I217718,I217965,I218216);
nor I_12684 (I217709,I218098,I218216);
or I_12685 (I217712,I217832,I218216);
DFFARX1 I_12686 (I218216,I2595,I217738,I217730,);
not I_12687 (I218316,I2602);
DFFARX1 I_12688 (I370602,I2595,I218316,I218342,);
not I_12689 (I218350,I218342);
nand I_12690 (I218367,I370590,I370608);
and I_12691 (I218384,I218367,I370599);
DFFARX1 I_12692 (I218384,I2595,I218316,I218410,);
not I_12693 (I218418,I370614);
DFFARX1 I_12694 (I370611,I2595,I218316,I218444,);
not I_12695 (I218452,I218444);
nor I_12696 (I218469,I218452,I218350);
and I_12697 (I218486,I218469,I370614);
nor I_12698 (I218503,I218452,I218418);
nor I_12699 (I218299,I218410,I218503);
DFFARX1 I_12700 (I370593,I2595,I218316,I218543,);
nor I_12701 (I218551,I218543,I218410);
not I_12702 (I218568,I218551);
not I_12703 (I218585,I218543);
nor I_12704 (I218602,I218585,I218486);
DFFARX1 I_12705 (I218602,I2595,I218316,I218302,);
nand I_12706 (I218633,I370587,I370587);
and I_12707 (I218650,I218633,I370596);
DFFARX1 I_12708 (I218650,I2595,I218316,I218676,);
nor I_12709 (I218684,I218676,I218543);
DFFARX1 I_12710 (I218684,I2595,I218316,I218284,);
nand I_12711 (I218715,I218676,I218585);
nand I_12712 (I218293,I218568,I218715);
not I_12713 (I218746,I218676);
nor I_12714 (I218763,I218746,I218486);
DFFARX1 I_12715 (I218763,I2595,I218316,I218305,);
nor I_12716 (I218794,I370605,I370587);
or I_12717 (I218296,I218543,I218794);
nor I_12718 (I218287,I218676,I218794);
or I_12719 (I218290,I218410,I218794);
DFFARX1 I_12720 (I218794,I2595,I218316,I218308,);
not I_12721 (I218894,I2602);
DFFARX1 I_12722 (I335092,I2595,I218894,I218920,);
not I_12723 (I218928,I218920);
nand I_12724 (I218945,I335074,I335086);
and I_12725 (I218962,I218945,I335089);
DFFARX1 I_12726 (I218962,I2595,I218894,I218988,);
not I_12727 (I218996,I335083);
DFFARX1 I_12728 (I335080,I2595,I218894,I219022,);
not I_12729 (I219030,I219022);
nor I_12730 (I219047,I219030,I218928);
and I_12731 (I219064,I219047,I335083);
nor I_12732 (I219081,I219030,I218996);
nor I_12733 (I218877,I218988,I219081);
DFFARX1 I_12734 (I335098,I2595,I218894,I219121,);
nor I_12735 (I219129,I219121,I218988);
not I_12736 (I219146,I219129);
not I_12737 (I219163,I219121);
nor I_12738 (I219180,I219163,I219064);
DFFARX1 I_12739 (I219180,I2595,I218894,I218880,);
nand I_12740 (I219211,I335077,I335077);
and I_12741 (I219228,I219211,I335074);
DFFARX1 I_12742 (I219228,I2595,I218894,I219254,);
nor I_12743 (I219262,I219254,I219121);
DFFARX1 I_12744 (I219262,I2595,I218894,I218862,);
nand I_12745 (I219293,I219254,I219163);
nand I_12746 (I218871,I219146,I219293);
not I_12747 (I219324,I219254);
nor I_12748 (I219341,I219324,I219064);
DFFARX1 I_12749 (I219341,I2595,I218894,I218883,);
nor I_12750 (I219372,I335095,I335077);
or I_12751 (I218874,I219121,I219372);
nor I_12752 (I218865,I219254,I219372);
or I_12753 (I218868,I218988,I219372);
DFFARX1 I_12754 (I219372,I2595,I218894,I218886,);
not I_12755 (I219472,I2602);
DFFARX1 I_12756 (I137730,I2595,I219472,I219498,);
not I_12757 (I219506,I219498);
nand I_12758 (I219523,I137721,I137739);
and I_12759 (I219540,I219523,I137742);
DFFARX1 I_12760 (I219540,I2595,I219472,I219566,);
not I_12761 (I219574,I137736);
DFFARX1 I_12762 (I137724,I2595,I219472,I219600,);
not I_12763 (I219608,I219600);
nor I_12764 (I219625,I219608,I219506);
and I_12765 (I219642,I219625,I137736);
nor I_12766 (I219659,I219608,I219574);
nor I_12767 (I219455,I219566,I219659);
DFFARX1 I_12768 (I137733,I2595,I219472,I219699,);
nor I_12769 (I219707,I219699,I219566);
not I_12770 (I219724,I219707);
not I_12771 (I219741,I219699);
nor I_12772 (I219758,I219741,I219642);
DFFARX1 I_12773 (I219758,I2595,I219472,I219458,);
nand I_12774 (I219789,I137748,I137745);
and I_12775 (I219806,I219789,I137727);
DFFARX1 I_12776 (I219806,I2595,I219472,I219832,);
nor I_12777 (I219840,I219832,I219699);
DFFARX1 I_12778 (I219840,I2595,I219472,I219440,);
nand I_12779 (I219871,I219832,I219741);
nand I_12780 (I219449,I219724,I219871);
not I_12781 (I219902,I219832);
nor I_12782 (I219919,I219902,I219642);
DFFARX1 I_12783 (I219919,I2595,I219472,I219461,);
nor I_12784 (I219950,I137721,I137745);
or I_12785 (I219452,I219699,I219950);
nor I_12786 (I219443,I219832,I219950);
or I_12787 (I219446,I219566,I219950);
DFFARX1 I_12788 (I219950,I2595,I219472,I219464,);
not I_12789 (I220050,I2602);
DFFARX1 I_12790 (I114882,I2595,I220050,I220076,);
not I_12791 (I220084,I220076);
nand I_12792 (I220101,I114873,I114891);
and I_12793 (I220118,I220101,I114894);
DFFARX1 I_12794 (I220118,I2595,I220050,I220144,);
not I_12795 (I220152,I114888);
DFFARX1 I_12796 (I114876,I2595,I220050,I220178,);
not I_12797 (I220186,I220178);
nor I_12798 (I220203,I220186,I220084);
and I_12799 (I220220,I220203,I114888);
nor I_12800 (I220237,I220186,I220152);
nor I_12801 (I220033,I220144,I220237);
DFFARX1 I_12802 (I114885,I2595,I220050,I220277,);
nor I_12803 (I220285,I220277,I220144);
not I_12804 (I220302,I220285);
not I_12805 (I220319,I220277);
nor I_12806 (I220336,I220319,I220220);
DFFARX1 I_12807 (I220336,I2595,I220050,I220036,);
nand I_12808 (I220367,I114900,I114897);
and I_12809 (I220384,I220367,I114879);
DFFARX1 I_12810 (I220384,I2595,I220050,I220410,);
nor I_12811 (I220418,I220410,I220277);
DFFARX1 I_12812 (I220418,I2595,I220050,I220018,);
nand I_12813 (I220449,I220410,I220319);
nand I_12814 (I220027,I220302,I220449);
not I_12815 (I220480,I220410);
nor I_12816 (I220497,I220480,I220220);
DFFARX1 I_12817 (I220497,I2595,I220050,I220039,);
nor I_12818 (I220528,I114873,I114897);
or I_12819 (I220030,I220277,I220528);
nor I_12820 (I220021,I220410,I220528);
or I_12821 (I220024,I220144,I220528);
DFFARX1 I_12822 (I220528,I2595,I220050,I220042,);
not I_12823 (I220628,I2602);
DFFARX1 I_12824 (I146935,I2595,I220628,I220654,);
not I_12825 (I220662,I220654);
nand I_12826 (I220679,I146950,I146935);
and I_12827 (I220696,I220679,I146938);
DFFARX1 I_12828 (I220696,I2595,I220628,I220722,);
not I_12829 (I220730,I146938);
DFFARX1 I_12830 (I146947,I2595,I220628,I220756,);
not I_12831 (I220764,I220756);
nor I_12832 (I220781,I220764,I220662);
and I_12833 (I220798,I220781,I146938);
nor I_12834 (I220815,I220764,I220730);
nor I_12835 (I220611,I220722,I220815);
DFFARX1 I_12836 (I146941,I2595,I220628,I220855,);
nor I_12837 (I220863,I220855,I220722);
not I_12838 (I220880,I220863);
not I_12839 (I220897,I220855);
nor I_12840 (I220914,I220897,I220798);
DFFARX1 I_12841 (I220914,I2595,I220628,I220614,);
nand I_12842 (I220945,I146944,I146953);
and I_12843 (I220962,I220945,I146959);
DFFARX1 I_12844 (I220962,I2595,I220628,I220988,);
nor I_12845 (I220996,I220988,I220855);
DFFARX1 I_12846 (I220996,I2595,I220628,I220596,);
nand I_12847 (I221027,I220988,I220897);
nand I_12848 (I220605,I220880,I221027);
not I_12849 (I221058,I220988);
nor I_12850 (I221075,I221058,I220798);
DFFARX1 I_12851 (I221075,I2595,I220628,I220617,);
nor I_12852 (I221106,I146956,I146953);
or I_12853 (I220608,I220855,I221106);
nor I_12854 (I220599,I220988,I221106);
or I_12855 (I220602,I220722,I221106);
DFFARX1 I_12856 (I221106,I2595,I220628,I220620,);
not I_12857 (I221206,I2602);
DFFARX1 I_12858 (I384860,I2595,I221206,I221232,);
not I_12859 (I221240,I221232);
nand I_12860 (I221257,I384845,I384833);
and I_12861 (I221274,I221257,I384848);
DFFARX1 I_12862 (I221274,I2595,I221206,I221300,);
not I_12863 (I221308,I384833);
DFFARX1 I_12864 (I384851,I2595,I221206,I221334,);
not I_12865 (I221342,I221334);
nor I_12866 (I221359,I221342,I221240);
and I_12867 (I221376,I221359,I384833);
nor I_12868 (I221393,I221342,I221308);
nor I_12869 (I221189,I221300,I221393);
DFFARX1 I_12870 (I384839,I2595,I221206,I221433,);
nor I_12871 (I221441,I221433,I221300);
not I_12872 (I221458,I221441);
not I_12873 (I221475,I221433);
nor I_12874 (I221492,I221475,I221376);
DFFARX1 I_12875 (I221492,I2595,I221206,I221192,);
nand I_12876 (I221523,I384836,I384842);
and I_12877 (I221540,I221523,I384857);
DFFARX1 I_12878 (I221540,I2595,I221206,I221566,);
nor I_12879 (I221574,I221566,I221433);
DFFARX1 I_12880 (I221574,I2595,I221206,I221174,);
nand I_12881 (I221605,I221566,I221475);
nand I_12882 (I221183,I221458,I221605);
not I_12883 (I221636,I221566);
nor I_12884 (I221653,I221636,I221376);
DFFARX1 I_12885 (I221653,I2595,I221206,I221195,);
nor I_12886 (I221684,I384854,I384842);
or I_12887 (I221186,I221433,I221684);
nor I_12888 (I221177,I221566,I221684);
or I_12889 (I221180,I221300,I221684);
DFFARX1 I_12890 (I221684,I2595,I221206,I221198,);
not I_12891 (I221784,I2602);
DFFARX1 I_12892 (I94871,I2595,I221784,I221810,);
not I_12893 (I221818,I221810);
nand I_12894 (I221835,I94874,I94850);
and I_12895 (I221852,I221835,I94847);
DFFARX1 I_12896 (I221852,I2595,I221784,I221878,);
not I_12897 (I221886,I94853);
DFFARX1 I_12898 (I94847,I2595,I221784,I221912,);
not I_12899 (I221920,I221912);
nor I_12900 (I221937,I221920,I221818);
and I_12901 (I221954,I221937,I94853);
nor I_12902 (I221971,I221920,I221886);
nor I_12903 (I221767,I221878,I221971);
DFFARX1 I_12904 (I94856,I2595,I221784,I222011,);
nor I_12905 (I222019,I222011,I221878);
not I_12906 (I222036,I222019);
not I_12907 (I222053,I222011);
nor I_12908 (I222070,I222053,I221954);
DFFARX1 I_12909 (I222070,I2595,I221784,I221770,);
nand I_12910 (I222101,I94859,I94868);
and I_12911 (I222118,I222101,I94865);
DFFARX1 I_12912 (I222118,I2595,I221784,I222144,);
nor I_12913 (I222152,I222144,I222011);
DFFARX1 I_12914 (I222152,I2595,I221784,I221752,);
nand I_12915 (I222183,I222144,I222053);
nand I_12916 (I221761,I222036,I222183);
not I_12917 (I222214,I222144);
nor I_12918 (I222231,I222214,I221954);
DFFARX1 I_12919 (I222231,I2595,I221784,I221773,);
nor I_12920 (I222262,I94862,I94868);
or I_12921 (I221764,I222011,I222262);
nor I_12922 (I221755,I222144,I222262);
or I_12923 (I221758,I221878,I222262);
DFFARX1 I_12924 (I222262,I2595,I221784,I221776,);
not I_12925 (I222362,I2602);
DFFARX1 I_12926 (I120866,I2595,I222362,I222388,);
not I_12927 (I222396,I222388);
nand I_12928 (I222413,I120857,I120875);
and I_12929 (I222430,I222413,I120878);
DFFARX1 I_12930 (I222430,I2595,I222362,I222456,);
not I_12931 (I222464,I120872);
DFFARX1 I_12932 (I120860,I2595,I222362,I222490,);
not I_12933 (I222498,I222490);
nor I_12934 (I222515,I222498,I222396);
and I_12935 (I222532,I222515,I120872);
nor I_12936 (I222549,I222498,I222464);
nor I_12937 (I222345,I222456,I222549);
DFFARX1 I_12938 (I120869,I2595,I222362,I222589,);
nor I_12939 (I222597,I222589,I222456);
not I_12940 (I222614,I222597);
not I_12941 (I222631,I222589);
nor I_12942 (I222648,I222631,I222532);
DFFARX1 I_12943 (I222648,I2595,I222362,I222348,);
nand I_12944 (I222679,I120884,I120881);
and I_12945 (I222696,I222679,I120863);
DFFARX1 I_12946 (I222696,I2595,I222362,I222722,);
nor I_12947 (I222730,I222722,I222589);
DFFARX1 I_12948 (I222730,I2595,I222362,I222330,);
nand I_12949 (I222761,I222722,I222631);
nand I_12950 (I222339,I222614,I222761);
not I_12951 (I222792,I222722);
nor I_12952 (I222809,I222792,I222532);
DFFARX1 I_12953 (I222809,I2595,I222362,I222351,);
nor I_12954 (I222840,I120857,I120881);
or I_12955 (I222342,I222589,I222840);
nor I_12956 (I222333,I222722,I222840);
or I_12957 (I222336,I222456,I222840);
DFFARX1 I_12958 (I222840,I2595,I222362,I222354,);
not I_12959 (I222940,I2602);
DFFARX1 I_12960 (I66933,I2595,I222940,I222966,);
not I_12961 (I222974,I222966);
nand I_12962 (I222991,I66936,I66957);
and I_12963 (I223008,I222991,I66945);
DFFARX1 I_12964 (I223008,I2595,I222940,I223034,);
not I_12965 (I223042,I66942);
DFFARX1 I_12966 (I66933,I2595,I222940,I223068,);
not I_12967 (I223076,I223068);
nor I_12968 (I223093,I223076,I222974);
and I_12969 (I223110,I223093,I66942);
nor I_12970 (I223127,I223076,I223042);
nor I_12971 (I222923,I223034,I223127);
DFFARX1 I_12972 (I66951,I2595,I222940,I223167,);
nor I_12973 (I223175,I223167,I223034);
not I_12974 (I223192,I223175);
not I_12975 (I223209,I223167);
nor I_12976 (I223226,I223209,I223110);
DFFARX1 I_12977 (I223226,I2595,I222940,I222926,);
nand I_12978 (I223257,I66936,I66939);
and I_12979 (I223274,I223257,I66948);
DFFARX1 I_12980 (I223274,I2595,I222940,I223300,);
nor I_12981 (I223308,I223300,I223167);
DFFARX1 I_12982 (I223308,I2595,I222940,I222908,);
nand I_12983 (I223339,I223300,I223209);
nand I_12984 (I222917,I223192,I223339);
not I_12985 (I223370,I223300);
nor I_12986 (I223387,I223370,I223110);
DFFARX1 I_12987 (I223387,I2595,I222940,I222929,);
nor I_12988 (I223418,I66954,I66939);
or I_12989 (I222920,I223167,I223418);
nor I_12990 (I222911,I223300,I223418);
or I_12991 (I222914,I223034,I223418);
DFFARX1 I_12992 (I223418,I2595,I222940,I222932,);
not I_12993 (I223518,I2602);
DFFARX1 I_12994 (I24504,I2595,I223518,I223544,);
not I_12995 (I223552,I223544);
nand I_12996 (I223569,I24513,I24522);
and I_12997 (I223586,I223569,I24501);
DFFARX1 I_12998 (I223586,I2595,I223518,I223612,);
not I_12999 (I223620,I24504);
DFFARX1 I_13000 (I24519,I2595,I223518,I223646,);
not I_13001 (I223654,I223646);
nor I_13002 (I223671,I223654,I223552);
and I_13003 (I223688,I223671,I24504);
nor I_13004 (I223705,I223654,I223620);
nor I_13005 (I223501,I223612,I223705);
DFFARX1 I_13006 (I24510,I2595,I223518,I223745,);
nor I_13007 (I223753,I223745,I223612);
not I_13008 (I223770,I223753);
not I_13009 (I223787,I223745);
nor I_13010 (I223804,I223787,I223688);
DFFARX1 I_13011 (I223804,I2595,I223518,I223504,);
nand I_13012 (I223835,I24525,I24501);
and I_13013 (I223852,I223835,I24507);
DFFARX1 I_13014 (I223852,I2595,I223518,I223878,);
nor I_13015 (I223886,I223878,I223745);
DFFARX1 I_13016 (I223886,I2595,I223518,I223486,);
nand I_13017 (I223917,I223878,I223787);
nand I_13018 (I223495,I223770,I223917);
not I_13019 (I223948,I223878);
nor I_13020 (I223965,I223948,I223688);
DFFARX1 I_13021 (I223965,I2595,I223518,I223507,);
nor I_13022 (I223996,I24516,I24501);
or I_13023 (I223498,I223745,I223996);
nor I_13024 (I223489,I223878,I223996);
or I_13025 (I223492,I223612,I223996);
DFFARX1 I_13026 (I223996,I2595,I223518,I223510,);
not I_13027 (I224096,I2602);
DFFARX1 I_13028 (I135010,I2595,I224096,I224122,);
not I_13029 (I224130,I224122);
nand I_13030 (I224147,I135001,I135019);
and I_13031 (I224164,I224147,I135022);
DFFARX1 I_13032 (I224164,I2595,I224096,I224190,);
not I_13033 (I224198,I135016);
DFFARX1 I_13034 (I135004,I2595,I224096,I224224,);
not I_13035 (I224232,I224224);
nor I_13036 (I224249,I224232,I224130);
and I_13037 (I224266,I224249,I135016);
nor I_13038 (I224283,I224232,I224198);
nor I_13039 (I224079,I224190,I224283);
DFFARX1 I_13040 (I135013,I2595,I224096,I224323,);
nor I_13041 (I224331,I224323,I224190);
not I_13042 (I224348,I224331);
not I_13043 (I224365,I224323);
nor I_13044 (I224382,I224365,I224266);
DFFARX1 I_13045 (I224382,I2595,I224096,I224082,);
nand I_13046 (I224413,I135028,I135025);
and I_13047 (I224430,I224413,I135007);
DFFARX1 I_13048 (I224430,I2595,I224096,I224456,);
nor I_13049 (I224464,I224456,I224323);
DFFARX1 I_13050 (I224464,I2595,I224096,I224064,);
nand I_13051 (I224495,I224456,I224365);
nand I_13052 (I224073,I224348,I224495);
not I_13053 (I224526,I224456);
nor I_13054 (I224543,I224526,I224266);
DFFARX1 I_13055 (I224543,I2595,I224096,I224085,);
nor I_13056 (I224574,I135001,I135025);
or I_13057 (I224076,I224323,I224574);
nor I_13058 (I224067,I224456,I224574);
or I_13059 (I224070,I224190,I224574);
DFFARX1 I_13060 (I224574,I2595,I224096,I224088,);
not I_13061 (I224674,I2602);
DFFARX1 I_13062 (I352414,I2595,I224674,I224700,);
not I_13063 (I224708,I224700);
nand I_13064 (I224725,I352417,I352426);
and I_13065 (I224742,I224725,I352429);
DFFARX1 I_13066 (I224742,I2595,I224674,I224768,);
not I_13067 (I224776,I352438);
DFFARX1 I_13068 (I352420,I2595,I224674,I224802,);
not I_13069 (I224810,I224802);
nor I_13070 (I224827,I224810,I224708);
and I_13071 (I224844,I224827,I352438);
nor I_13072 (I224861,I224810,I224776);
nor I_13073 (I224657,I224768,I224861);
DFFARX1 I_13074 (I352417,I2595,I224674,I224901,);
nor I_13075 (I224909,I224901,I224768);
not I_13076 (I224926,I224909);
not I_13077 (I224943,I224901);
nor I_13078 (I224960,I224943,I224844);
DFFARX1 I_13079 (I224960,I2595,I224674,I224660,);
nand I_13080 (I224991,I352435,I352414);
and I_13081 (I225008,I224991,I352432);
DFFARX1 I_13082 (I225008,I2595,I224674,I225034,);
nor I_13083 (I225042,I225034,I224901);
DFFARX1 I_13084 (I225042,I2595,I224674,I224642,);
nand I_13085 (I225073,I225034,I224943);
nand I_13086 (I224651,I224926,I225073);
not I_13087 (I225104,I225034);
nor I_13088 (I225121,I225104,I224844);
DFFARX1 I_13089 (I225121,I2595,I224674,I224663,);
nor I_13090 (I225152,I352423,I352414);
or I_13091 (I224654,I224901,I225152);
nor I_13092 (I224645,I225034,I225152);
or I_13093 (I224648,I224768,I225152);
DFFARX1 I_13094 (I225152,I2595,I224674,I224666,);
not I_13095 (I225252,I2602);
DFFARX1 I_13096 (I371770,I2595,I225252,I225278,);
not I_13097 (I225286,I225278);
nand I_13098 (I225303,I371755,I371743);
and I_13099 (I225320,I225303,I371758);
DFFARX1 I_13100 (I225320,I2595,I225252,I225346,);
not I_13101 (I225354,I371743);
DFFARX1 I_13102 (I371761,I2595,I225252,I225380,);
not I_13103 (I225388,I225380);
nor I_13104 (I225405,I225388,I225286);
and I_13105 (I225422,I225405,I371743);
nor I_13106 (I225439,I225388,I225354);
nor I_13107 (I225235,I225346,I225439);
DFFARX1 I_13108 (I371749,I2595,I225252,I225479,);
nor I_13109 (I225487,I225479,I225346);
not I_13110 (I225504,I225487);
not I_13111 (I225521,I225479);
nor I_13112 (I225538,I225521,I225422);
DFFARX1 I_13113 (I225538,I2595,I225252,I225238,);
nand I_13114 (I225569,I371746,I371752);
and I_13115 (I225586,I225569,I371767);
DFFARX1 I_13116 (I225586,I2595,I225252,I225612,);
nor I_13117 (I225620,I225612,I225479);
DFFARX1 I_13118 (I225620,I2595,I225252,I225220,);
nand I_13119 (I225651,I225612,I225521);
nand I_13120 (I225229,I225504,I225651);
not I_13121 (I225682,I225612);
nor I_13122 (I225699,I225682,I225422);
DFFARX1 I_13123 (I225699,I2595,I225252,I225241,);
nor I_13124 (I225730,I371764,I371752);
or I_13125 (I225232,I225479,I225730);
nor I_13126 (I225223,I225612,I225730);
or I_13127 (I225226,I225346,I225730);
DFFARX1 I_13128 (I225730,I2595,I225252,I225244,);
not I_13129 (I225830,I2602);
DFFARX1 I_13130 (I50868,I2595,I225830,I225856,);
not I_13131 (I225864,I225856);
nand I_13132 (I225881,I50871,I50892);
and I_13133 (I225898,I225881,I50880);
DFFARX1 I_13134 (I225898,I2595,I225830,I225924,);
not I_13135 (I225932,I50877);
DFFARX1 I_13136 (I50868,I2595,I225830,I225958,);
not I_13137 (I225966,I225958);
nor I_13138 (I225983,I225966,I225864);
and I_13139 (I226000,I225983,I50877);
nor I_13140 (I226017,I225966,I225932);
nor I_13141 (I225813,I225924,I226017);
DFFARX1 I_13142 (I50886,I2595,I225830,I226057,);
nor I_13143 (I226065,I226057,I225924);
not I_13144 (I226082,I226065);
not I_13145 (I226099,I226057);
nor I_13146 (I226116,I226099,I226000);
DFFARX1 I_13147 (I226116,I2595,I225830,I225816,);
nand I_13148 (I226147,I50871,I50874);
and I_13149 (I226164,I226147,I50883);
DFFARX1 I_13150 (I226164,I2595,I225830,I226190,);
nor I_13151 (I226198,I226190,I226057);
DFFARX1 I_13152 (I226198,I2595,I225830,I225798,);
nand I_13153 (I226229,I226190,I226099);
nand I_13154 (I225807,I226082,I226229);
not I_13155 (I226260,I226190);
nor I_13156 (I226277,I226260,I226000);
DFFARX1 I_13157 (I226277,I2595,I225830,I225819,);
nor I_13158 (I226308,I50889,I50874);
or I_13159 (I225810,I226057,I226308);
nor I_13160 (I225801,I226190,I226308);
or I_13161 (I225804,I225924,I226308);
DFFARX1 I_13162 (I226308,I2595,I225830,I225822,);
not I_13163 (I226408,I2602);
DFFARX1 I_13164 (I152290,I2595,I226408,I226434,);
not I_13165 (I226442,I226434);
nand I_13166 (I226459,I152305,I152290);
and I_13167 (I226476,I226459,I152293);
DFFARX1 I_13168 (I226476,I2595,I226408,I226502,);
not I_13169 (I226510,I152293);
DFFARX1 I_13170 (I152302,I2595,I226408,I226536,);
not I_13171 (I226544,I226536);
nor I_13172 (I226561,I226544,I226442);
and I_13173 (I226578,I226561,I152293);
nor I_13174 (I226595,I226544,I226510);
nor I_13175 (I226391,I226502,I226595);
DFFARX1 I_13176 (I152296,I2595,I226408,I226635,);
nor I_13177 (I226643,I226635,I226502);
not I_13178 (I226660,I226643);
not I_13179 (I226677,I226635);
nor I_13180 (I226694,I226677,I226578);
DFFARX1 I_13181 (I226694,I2595,I226408,I226394,);
nand I_13182 (I226725,I152299,I152308);
and I_13183 (I226742,I226725,I152314);
DFFARX1 I_13184 (I226742,I2595,I226408,I226768,);
nor I_13185 (I226776,I226768,I226635);
DFFARX1 I_13186 (I226776,I2595,I226408,I226376,);
nand I_13187 (I226807,I226768,I226677);
nand I_13188 (I226385,I226660,I226807);
not I_13189 (I226838,I226768);
nor I_13190 (I226855,I226838,I226578);
DFFARX1 I_13191 (I226855,I2595,I226408,I226397,);
nor I_13192 (I226886,I152311,I152308);
or I_13193 (I226388,I226635,I226886);
nor I_13194 (I226379,I226768,I226886);
or I_13195 (I226382,I226502,I226886);
DFFARX1 I_13196 (I226886,I2595,I226408,I226400,);
not I_13197 (I226986,I2602);
DFFARX1 I_13198 (I284183,I2595,I226986,I227012,);
not I_13199 (I227020,I227012);
nand I_13200 (I227037,I284159,I284174);
and I_13201 (I227054,I227037,I284186);
DFFARX1 I_13202 (I227054,I2595,I226986,I227080,);
not I_13203 (I227088,I284171);
DFFARX1 I_13204 (I284162,I2595,I226986,I227114,);
not I_13205 (I227122,I227114);
nor I_13206 (I227139,I227122,I227020);
and I_13207 (I227156,I227139,I284171);
nor I_13208 (I227173,I227122,I227088);
nor I_13209 (I226969,I227080,I227173);
DFFARX1 I_13210 (I284159,I2595,I226986,I227213,);
nor I_13211 (I227221,I227213,I227080);
not I_13212 (I227238,I227221);
not I_13213 (I227255,I227213);
nor I_13214 (I227272,I227255,I227156);
DFFARX1 I_13215 (I227272,I2595,I226986,I226972,);
nand I_13216 (I227303,I284177,I284168);
and I_13217 (I227320,I227303,I284180);
DFFARX1 I_13218 (I227320,I2595,I226986,I227346,);
nor I_13219 (I227354,I227346,I227213);
DFFARX1 I_13220 (I227354,I2595,I226986,I226954,);
nand I_13221 (I227385,I227346,I227255);
nand I_13222 (I226963,I227238,I227385);
not I_13223 (I227416,I227346);
nor I_13224 (I227433,I227416,I227156);
DFFARX1 I_13225 (I227433,I2595,I226986,I226975,);
nor I_13226 (I227464,I284165,I284168);
or I_13227 (I226966,I227213,I227464);
nor I_13228 (I226957,I227346,I227464);
or I_13229 (I226960,I227080,I227464);
DFFARX1 I_13230 (I227464,I2595,I226986,I226978,);
not I_13231 (I227564,I2602);
DFFARX1 I_13232 (I340294,I2595,I227564,I227590,);
not I_13233 (I227598,I227590);
nand I_13234 (I227615,I340276,I340288);
and I_13235 (I227632,I227615,I340291);
DFFARX1 I_13236 (I227632,I2595,I227564,I227658,);
not I_13237 (I227666,I340285);
DFFARX1 I_13238 (I340282,I2595,I227564,I227692,);
not I_13239 (I227700,I227692);
nor I_13240 (I227717,I227700,I227598);
and I_13241 (I227734,I227717,I340285);
nor I_13242 (I227751,I227700,I227666);
nor I_13243 (I227547,I227658,I227751);
DFFARX1 I_13244 (I340300,I2595,I227564,I227791,);
nor I_13245 (I227799,I227791,I227658);
not I_13246 (I227816,I227799);
not I_13247 (I227833,I227791);
nor I_13248 (I227850,I227833,I227734);
DFFARX1 I_13249 (I227850,I2595,I227564,I227550,);
nand I_13250 (I227881,I340279,I340279);
and I_13251 (I227898,I227881,I340276);
DFFARX1 I_13252 (I227898,I2595,I227564,I227924,);
nor I_13253 (I227932,I227924,I227791);
DFFARX1 I_13254 (I227932,I2595,I227564,I227532,);
nand I_13255 (I227963,I227924,I227833);
nand I_13256 (I227541,I227816,I227963);
not I_13257 (I227994,I227924);
nor I_13258 (I228011,I227994,I227734);
DFFARX1 I_13259 (I228011,I2595,I227564,I227553,);
nor I_13260 (I228042,I340297,I340279);
or I_13261 (I227544,I227791,I228042);
nor I_13262 (I227535,I227924,I228042);
or I_13263 (I227538,I227658,I228042);
DFFARX1 I_13264 (I228042,I2595,I227564,I227556,);
not I_13265 (I228142,I2602);
DFFARX1 I_13266 (I279015,I2595,I228142,I228168,);
not I_13267 (I228176,I228168);
nand I_13268 (I228193,I278991,I279006);
and I_13269 (I228210,I228193,I279018);
DFFARX1 I_13270 (I228210,I2595,I228142,I228236,);
not I_13271 (I228244,I279003);
DFFARX1 I_13272 (I278994,I2595,I228142,I228270,);
not I_13273 (I228278,I228270);
nor I_13274 (I228295,I228278,I228176);
and I_13275 (I228312,I228295,I279003);
nor I_13276 (I228329,I228278,I228244);
nor I_13277 (I228125,I228236,I228329);
DFFARX1 I_13278 (I278991,I2595,I228142,I228369,);
nor I_13279 (I228377,I228369,I228236);
not I_13280 (I228394,I228377);
not I_13281 (I228411,I228369);
nor I_13282 (I228428,I228411,I228312);
DFFARX1 I_13283 (I228428,I2595,I228142,I228128,);
nand I_13284 (I228459,I279009,I279000);
and I_13285 (I228476,I228459,I279012);
DFFARX1 I_13286 (I228476,I2595,I228142,I228502,);
nor I_13287 (I228510,I228502,I228369);
DFFARX1 I_13288 (I228510,I2595,I228142,I228110,);
nand I_13289 (I228541,I228502,I228411);
nand I_13290 (I228119,I228394,I228541);
not I_13291 (I228572,I228502);
nor I_13292 (I228589,I228572,I228312);
DFFARX1 I_13293 (I228589,I2595,I228142,I228131,);
nor I_13294 (I228620,I278997,I279000);
or I_13295 (I228122,I228369,I228620);
nor I_13296 (I228113,I228502,I228620);
or I_13297 (I228116,I228236,I228620);
DFFARX1 I_13298 (I228620,I2595,I228142,I228134,);
not I_13299 (I228720,I2602);
DFFARX1 I_13300 (I89074,I2595,I228720,I228746,);
not I_13301 (I228754,I228746);
nand I_13302 (I228771,I89077,I89053);
and I_13303 (I228788,I228771,I89050);
DFFARX1 I_13304 (I228788,I2595,I228720,I228814,);
not I_13305 (I228822,I89056);
DFFARX1 I_13306 (I89050,I2595,I228720,I228848,);
not I_13307 (I228856,I228848);
nor I_13308 (I228873,I228856,I228754);
and I_13309 (I228890,I228873,I89056);
nor I_13310 (I228907,I228856,I228822);
nor I_13311 (I228703,I228814,I228907);
DFFARX1 I_13312 (I89059,I2595,I228720,I228947,);
nor I_13313 (I228955,I228947,I228814);
not I_13314 (I228972,I228955);
not I_13315 (I228989,I228947);
nor I_13316 (I229006,I228989,I228890);
DFFARX1 I_13317 (I229006,I2595,I228720,I228706,);
nand I_13318 (I229037,I89062,I89071);
and I_13319 (I229054,I229037,I89068);
DFFARX1 I_13320 (I229054,I2595,I228720,I229080,);
nor I_13321 (I229088,I229080,I228947);
DFFARX1 I_13322 (I229088,I2595,I228720,I228688,);
nand I_13323 (I229119,I229080,I228989);
nand I_13324 (I228697,I228972,I229119);
not I_13325 (I229150,I229080);
nor I_13326 (I229167,I229150,I228890);
DFFARX1 I_13327 (I229167,I2595,I228720,I228709,);
nor I_13328 (I229198,I89065,I89071);
or I_13329 (I228700,I228947,I229198);
nor I_13330 (I228691,I229080,I229198);
or I_13331 (I228694,I228814,I229198);
DFFARX1 I_13332 (I229198,I2595,I228720,I228712,);
not I_13333 (I229298,I2602);
DFFARX1 I_13334 (I317752,I2595,I229298,I229324,);
not I_13335 (I229332,I229324);
nand I_13336 (I229349,I317734,I317746);
and I_13337 (I229366,I229349,I317749);
DFFARX1 I_13338 (I229366,I2595,I229298,I229392,);
not I_13339 (I229400,I317743);
DFFARX1 I_13340 (I317740,I2595,I229298,I229426,);
not I_13341 (I229434,I229426);
nor I_13342 (I229451,I229434,I229332);
and I_13343 (I229468,I229451,I317743);
nor I_13344 (I229485,I229434,I229400);
nor I_13345 (I229281,I229392,I229485);
DFFARX1 I_13346 (I317758,I2595,I229298,I229525,);
nor I_13347 (I229533,I229525,I229392);
not I_13348 (I229550,I229533);
not I_13349 (I229567,I229525);
nor I_13350 (I229584,I229567,I229468);
DFFARX1 I_13351 (I229584,I2595,I229298,I229284,);
nand I_13352 (I229615,I317737,I317737);
and I_13353 (I229632,I229615,I317734);
DFFARX1 I_13354 (I229632,I2595,I229298,I229658,);
nor I_13355 (I229666,I229658,I229525);
DFFARX1 I_13356 (I229666,I2595,I229298,I229266,);
nand I_13357 (I229697,I229658,I229567);
nand I_13358 (I229275,I229550,I229697);
not I_13359 (I229728,I229658);
nor I_13360 (I229745,I229728,I229468);
DFFARX1 I_13361 (I229745,I2595,I229298,I229287,);
nor I_13362 (I229776,I317755,I317737);
or I_13363 (I229278,I229525,I229776);
nor I_13364 (I229269,I229658,I229776);
or I_13365 (I229272,I229392,I229776);
DFFARX1 I_13366 (I229776,I2595,I229298,I229290,);
not I_13367 (I229873,I2602);
DFFARX1 I_13368 (I257030,I2595,I229873,I229899,);
not I_13369 (I229907,I229899);
nand I_13370 (I229924,I257045,I257027);
and I_13371 (I229941,I229924,I257027);
DFFARX1 I_13372 (I229941,I2595,I229873,I229967,);
DFFARX1 I_13373 (I229967,I2595,I229873,I229862,);
DFFARX1 I_13374 (I257036,I2595,I229873,I229998,);
nand I_13375 (I230006,I229998,I257054);
not I_13376 (I230023,I230006);
DFFARX1 I_13377 (I230023,I2595,I229873,I230049,);
not I_13378 (I230057,I230049);
nor I_13379 (I229865,I229907,I230057);
DFFARX1 I_13380 (I257051,I2595,I229873,I230097,);
nor I_13381 (I229856,I230097,I229967);
nor I_13382 (I229847,I230097,I230023);
nand I_13383 (I230133,I257048,I257039);
and I_13384 (I230150,I230133,I257033);
DFFARX1 I_13385 (I230150,I2595,I229873,I230176,);
not I_13386 (I230184,I230176);
nand I_13387 (I230201,I230184,I230097);
nand I_13388 (I229850,I230184,I230006);
nor I_13389 (I230232,I257042,I257039);
and I_13390 (I230249,I230097,I230232);
nor I_13391 (I230266,I230184,I230249);
DFFARX1 I_13392 (I230266,I2595,I229873,I229859,);
nor I_13393 (I230297,I229899,I230232);
DFFARX1 I_13394 (I230297,I2595,I229873,I229844,);
nor I_13395 (I230328,I230176,I230232);
not I_13396 (I230345,I230328);
nand I_13397 (I229853,I230345,I230201);
not I_13398 (I230400,I2602);
DFFARX1 I_13399 (I203834,I2595,I230400,I230426,);
not I_13400 (I230434,I230426);
nand I_13401 (I230451,I203837,I203834);
and I_13402 (I230468,I230451,I203846);
DFFARX1 I_13403 (I230468,I2595,I230400,I230494,);
DFFARX1 I_13404 (I230494,I2595,I230400,I230389,);
DFFARX1 I_13405 (I203843,I2595,I230400,I230525,);
nand I_13406 (I230533,I230525,I203849);
not I_13407 (I230550,I230533);
DFFARX1 I_13408 (I230550,I2595,I230400,I230576,);
not I_13409 (I230584,I230576);
nor I_13410 (I230392,I230434,I230584);
DFFARX1 I_13411 (I203858,I2595,I230400,I230624,);
nor I_13412 (I230383,I230624,I230494);
nor I_13413 (I230374,I230624,I230550);
nand I_13414 (I230660,I203852,I203840);
and I_13415 (I230677,I230660,I203837);
DFFARX1 I_13416 (I230677,I2595,I230400,I230703,);
not I_13417 (I230711,I230703);
nand I_13418 (I230728,I230711,I230624);
nand I_13419 (I230377,I230711,I230533);
nor I_13420 (I230759,I203855,I203840);
and I_13421 (I230776,I230624,I230759);
nor I_13422 (I230793,I230711,I230776);
DFFARX1 I_13423 (I230793,I2595,I230400,I230386,);
nor I_13424 (I230824,I230426,I230759);
DFFARX1 I_13425 (I230824,I2595,I230400,I230371,);
nor I_13426 (I230855,I230703,I230759);
not I_13427 (I230872,I230855);
nand I_13428 (I230380,I230872,I230728);
not I_13429 (I230927,I2602);
DFFARX1 I_13430 (I172059,I2595,I230927,I230953,);
not I_13431 (I230961,I230953);
nand I_13432 (I230978,I172044,I172065);
and I_13433 (I230995,I230978,I172053);
DFFARX1 I_13434 (I230995,I2595,I230927,I231021,);
DFFARX1 I_13435 (I231021,I2595,I230927,I230916,);
DFFARX1 I_13436 (I172047,I2595,I230927,I231052,);
nand I_13437 (I231060,I231052,I172056);
not I_13438 (I231077,I231060);
DFFARX1 I_13439 (I231077,I2595,I230927,I231103,);
not I_13440 (I231111,I231103);
nor I_13441 (I230919,I230961,I231111);
DFFARX1 I_13442 (I172062,I2595,I230927,I231151,);
nor I_13443 (I230910,I231151,I231021);
nor I_13444 (I230901,I231151,I231077);
nand I_13445 (I231187,I172044,I172047);
and I_13446 (I231204,I231187,I172068);
DFFARX1 I_13447 (I231204,I2595,I230927,I231230,);
not I_13448 (I231238,I231230);
nand I_13449 (I231255,I231238,I231151);
nand I_13450 (I230904,I231238,I231060);
nor I_13451 (I231286,I172050,I172047);
and I_13452 (I231303,I231151,I231286);
nor I_13453 (I231320,I231238,I231303);
DFFARX1 I_13454 (I231320,I2595,I230927,I230913,);
nor I_13455 (I231351,I230953,I231286);
DFFARX1 I_13456 (I231351,I2595,I230927,I230898,);
nor I_13457 (I231382,I231230,I231286);
not I_13458 (I231399,I231382);
nand I_13459 (I230907,I231399,I231255);
not I_13460 (I231454,I2602);
DFFARX1 I_13461 (I302239,I2595,I231454,I231480,);
not I_13462 (I231488,I231480);
nand I_13463 (I231505,I302248,I302236);
and I_13464 (I231522,I231505,I302233);
DFFARX1 I_13465 (I231522,I2595,I231454,I231548,);
DFFARX1 I_13466 (I231548,I2595,I231454,I231443,);
DFFARX1 I_13467 (I302233,I2595,I231454,I231579,);
nand I_13468 (I231587,I231579,I302230);
not I_13469 (I231604,I231587);
DFFARX1 I_13470 (I231604,I2595,I231454,I231630,);
not I_13471 (I231638,I231630);
nor I_13472 (I231446,I231488,I231638);
DFFARX1 I_13473 (I302236,I2595,I231454,I231678,);
nor I_13474 (I231437,I231678,I231548);
nor I_13475 (I231428,I231678,I231604);
nand I_13476 (I231714,I302251,I302242);
and I_13477 (I231731,I231714,I302245);
DFFARX1 I_13478 (I231731,I2595,I231454,I231757,);
not I_13479 (I231765,I231757);
nand I_13480 (I231782,I231765,I231678);
nand I_13481 (I231431,I231765,I231587);
nor I_13482 (I231813,I302230,I302242);
and I_13483 (I231830,I231678,I231813);
nor I_13484 (I231847,I231765,I231830);
DFFARX1 I_13485 (I231847,I2595,I231454,I231440,);
nor I_13486 (I231878,I231480,I231813);
DFFARX1 I_13487 (I231878,I2595,I231454,I231425,);
nor I_13488 (I231909,I231757,I231813);
not I_13489 (I231926,I231909);
nand I_13490 (I231434,I231926,I231782);
not I_13491 (I231981,I2602);
DFFARX1 I_13492 (I53254,I2595,I231981,I232007,);
not I_13493 (I232015,I232007);
nand I_13494 (I232032,I53251,I53269);
and I_13495 (I232049,I232032,I53260);
DFFARX1 I_13496 (I232049,I2595,I231981,I232075,);
DFFARX1 I_13497 (I232075,I2595,I231981,I231970,);
DFFARX1 I_13498 (I53266,I2595,I231981,I232106,);
nand I_13499 (I232114,I232106,I53263);
not I_13500 (I232131,I232114);
DFFARX1 I_13501 (I232131,I2595,I231981,I232157,);
not I_13502 (I232165,I232157);
nor I_13503 (I231973,I232015,I232165);
DFFARX1 I_13504 (I53257,I2595,I231981,I232205,);
nor I_13505 (I231964,I232205,I232075);
nor I_13506 (I231955,I232205,I232131);
nand I_13507 (I232241,I53248,I53272);
and I_13508 (I232258,I232241,I53251);
DFFARX1 I_13509 (I232258,I2595,I231981,I232284,);
not I_13510 (I232292,I232284);
nand I_13511 (I232309,I232292,I232205);
nand I_13512 (I231958,I232292,I232114);
nor I_13513 (I232340,I53248,I53272);
and I_13514 (I232357,I232205,I232340);
nor I_13515 (I232374,I232292,I232357);
DFFARX1 I_13516 (I232374,I2595,I231981,I231967,);
nor I_13517 (I232405,I232007,I232340);
DFFARX1 I_13518 (I232405,I2595,I231981,I231952,);
nor I_13519 (I232436,I232284,I232340);
not I_13520 (I232453,I232436);
nand I_13521 (I231961,I232453,I232309);
not I_13522 (I232508,I2602);
DFFARX1 I_13523 (I191696,I2595,I232508,I232534,);
not I_13524 (I232542,I232534);
nand I_13525 (I232559,I191699,I191696);
and I_13526 (I232576,I232559,I191708);
DFFARX1 I_13527 (I232576,I2595,I232508,I232602,);
DFFARX1 I_13528 (I232602,I2595,I232508,I232497,);
DFFARX1 I_13529 (I191705,I2595,I232508,I232633,);
nand I_13530 (I232641,I232633,I191711);
not I_13531 (I232658,I232641);
DFFARX1 I_13532 (I232658,I2595,I232508,I232684,);
not I_13533 (I232692,I232684);
nor I_13534 (I232500,I232542,I232692);
DFFARX1 I_13535 (I191720,I2595,I232508,I232732,);
nor I_13536 (I232491,I232732,I232602);
nor I_13537 (I232482,I232732,I232658);
nand I_13538 (I232768,I191714,I191702);
and I_13539 (I232785,I232768,I191699);
DFFARX1 I_13540 (I232785,I2595,I232508,I232811,);
not I_13541 (I232819,I232811);
nand I_13542 (I232836,I232819,I232732);
nand I_13543 (I232485,I232819,I232641);
nor I_13544 (I232867,I191717,I191702);
and I_13545 (I232884,I232732,I232867);
nor I_13546 (I232901,I232819,I232884);
DFFARX1 I_13547 (I232901,I2595,I232508,I232494,);
nor I_13548 (I232932,I232534,I232867);
DFFARX1 I_13549 (I232932,I2595,I232508,I232479,);
nor I_13550 (I232963,I232811,I232867);
not I_13551 (I232980,I232963);
nand I_13552 (I232488,I232980,I232836);
not I_13553 (I233035,I2602);
DFFARX1 I_13554 (I338560,I2595,I233035,I233061,);
not I_13555 (I233069,I233061);
nand I_13556 (I233086,I338542,I338542);
and I_13557 (I233103,I233086,I338548);
DFFARX1 I_13558 (I233103,I2595,I233035,I233129,);
DFFARX1 I_13559 (I233129,I2595,I233035,I233024,);
DFFARX1 I_13560 (I338545,I2595,I233035,I233160,);
nand I_13561 (I233168,I233160,I338554);
not I_13562 (I233185,I233168);
DFFARX1 I_13563 (I233185,I2595,I233035,I233211,);
not I_13564 (I233219,I233211);
nor I_13565 (I233027,I233069,I233219);
DFFARX1 I_13566 (I338566,I2595,I233035,I233259,);
nor I_13567 (I233018,I233259,I233129);
nor I_13568 (I233009,I233259,I233185);
nand I_13569 (I233295,I338557,I338551);
and I_13570 (I233312,I233295,I338545);
DFFARX1 I_13571 (I233312,I2595,I233035,I233338,);
not I_13572 (I233346,I233338);
nand I_13573 (I233363,I233346,I233259);
nand I_13574 (I233012,I233346,I233168);
nor I_13575 (I233394,I338563,I338551);
and I_13576 (I233411,I233259,I233394);
nor I_13577 (I233428,I233346,I233411);
DFFARX1 I_13578 (I233428,I2595,I233035,I233021,);
nor I_13579 (I233459,I233061,I233394);
DFFARX1 I_13580 (I233459,I2595,I233035,I233006,);
nor I_13581 (I233490,I233338,I233394);
not I_13582 (I233507,I233490);
nand I_13583 (I233015,I233507,I233363);
not I_13584 (I233562,I2602);
DFFARX1 I_13585 (I260906,I2595,I233562,I233588,);
not I_13586 (I233596,I233588);
nand I_13587 (I233613,I260921,I260903);
and I_13588 (I233630,I233613,I260903);
DFFARX1 I_13589 (I233630,I2595,I233562,I233656,);
DFFARX1 I_13590 (I233656,I2595,I233562,I233551,);
DFFARX1 I_13591 (I260912,I2595,I233562,I233687,);
nand I_13592 (I233695,I233687,I260930);
not I_13593 (I233712,I233695);
DFFARX1 I_13594 (I233712,I2595,I233562,I233738,);
not I_13595 (I233746,I233738);
nor I_13596 (I233554,I233596,I233746);
DFFARX1 I_13597 (I260927,I2595,I233562,I233786,);
nor I_13598 (I233545,I233786,I233656);
nor I_13599 (I233536,I233786,I233712);
nand I_13600 (I233822,I260924,I260915);
and I_13601 (I233839,I233822,I260909);
DFFARX1 I_13602 (I233839,I2595,I233562,I233865,);
not I_13603 (I233873,I233865);
nand I_13604 (I233890,I233873,I233786);
nand I_13605 (I233539,I233873,I233695);
nor I_13606 (I233921,I260918,I260915);
and I_13607 (I233938,I233786,I233921);
nor I_13608 (I233955,I233873,I233938);
DFFARX1 I_13609 (I233955,I2595,I233562,I233548,);
nor I_13610 (I233986,I233588,I233921);
DFFARX1 I_13611 (I233986,I2595,I233562,I233533,);
nor I_13612 (I234017,I233865,I233921);
not I_13613 (I234034,I234017);
nand I_13614 (I233542,I234034,I233890);
not I_13615 (I234089,I2602);
DFFARX1 I_13616 (I93802,I2595,I234089,I234115,);
not I_13617 (I234123,I234115);
nand I_13618 (I234140,I93793,I93793);
and I_13619 (I234157,I234140,I93811);
DFFARX1 I_13620 (I234157,I2595,I234089,I234183,);
DFFARX1 I_13621 (I234183,I2595,I234089,I234078,);
DFFARX1 I_13622 (I93814,I2595,I234089,I234214,);
nand I_13623 (I234222,I234214,I93796);
not I_13624 (I234239,I234222);
DFFARX1 I_13625 (I234239,I2595,I234089,I234265,);
not I_13626 (I234273,I234265);
nor I_13627 (I234081,I234123,I234273);
DFFARX1 I_13628 (I93808,I2595,I234089,I234313,);
nor I_13629 (I234072,I234313,I234183);
nor I_13630 (I234063,I234313,I234239);
nand I_13631 (I234349,I93820,I93799);
and I_13632 (I234366,I234349,I93805);
DFFARX1 I_13633 (I234366,I2595,I234089,I234392,);
not I_13634 (I234400,I234392);
nand I_13635 (I234417,I234400,I234313);
nand I_13636 (I234066,I234400,I234222);
nor I_13637 (I234448,I93817,I93799);
and I_13638 (I234465,I234313,I234448);
nor I_13639 (I234482,I234400,I234465);
DFFARX1 I_13640 (I234482,I2595,I234089,I234075,);
nor I_13641 (I234513,I234115,I234448);
DFFARX1 I_13642 (I234513,I2595,I234089,I234060,);
nor I_13643 (I234544,I234392,I234448);
not I_13644 (I234561,I234544);
nand I_13645 (I234069,I234561,I234417);
not I_13646 (I234616,I2602);
DFFARX1 I_13647 (I391393,I2595,I234616,I234642,);
not I_13648 (I234650,I234642);
nand I_13649 (I234667,I391390,I391399);
and I_13650 (I234684,I234667,I391378);
DFFARX1 I_13651 (I234684,I2595,I234616,I234710,);
DFFARX1 I_13652 (I234710,I2595,I234616,I234605,);
DFFARX1 I_13653 (I391381,I2595,I234616,I234741,);
nand I_13654 (I234749,I234741,I391396);
not I_13655 (I234766,I234749);
DFFARX1 I_13656 (I234766,I2595,I234616,I234792,);
not I_13657 (I234800,I234792);
nor I_13658 (I234608,I234650,I234800);
DFFARX1 I_13659 (I391402,I2595,I234616,I234840,);
nor I_13660 (I234599,I234840,I234710);
nor I_13661 (I234590,I234840,I234766);
nand I_13662 (I234876,I391384,I391405);
and I_13663 (I234893,I234876,I391387);
DFFARX1 I_13664 (I234893,I2595,I234616,I234919,);
not I_13665 (I234927,I234919);
nand I_13666 (I234944,I234927,I234840);
nand I_13667 (I234593,I234927,I234749);
nor I_13668 (I234975,I391378,I391405);
and I_13669 (I234992,I234840,I234975);
nor I_13670 (I235009,I234927,I234992);
DFFARX1 I_13671 (I235009,I2595,I234616,I234602,);
nor I_13672 (I235040,I234642,I234975);
DFFARX1 I_13673 (I235040,I2595,I234616,I234587,);
nor I_13674 (I235071,I234919,I234975);
not I_13675 (I235088,I235071);
nand I_13676 (I234596,I235088,I234944);
not I_13677 (I235143,I2602);
DFFARX1 I_13678 (I151701,I2595,I235143,I235169,);
not I_13679 (I235177,I235169);
nand I_13680 (I235194,I151719,I151710);
and I_13681 (I235211,I235194,I151713);
DFFARX1 I_13682 (I235211,I2595,I235143,I235237,);
DFFARX1 I_13683 (I235237,I2595,I235143,I235132,);
DFFARX1 I_13684 (I151707,I2595,I235143,I235268,);
nand I_13685 (I235276,I235268,I151698);
not I_13686 (I235293,I235276);
DFFARX1 I_13687 (I235293,I2595,I235143,I235319,);
not I_13688 (I235327,I235319);
nor I_13689 (I235135,I235177,I235327);
DFFARX1 I_13690 (I151704,I2595,I235143,I235367,);
nor I_13691 (I235126,I235367,I235237);
nor I_13692 (I235117,I235367,I235293);
nand I_13693 (I235403,I151698,I151695);
and I_13694 (I235420,I235403,I151716);
DFFARX1 I_13695 (I235420,I2595,I235143,I235446,);
not I_13696 (I235454,I235446);
nand I_13697 (I235471,I235454,I235367);
nand I_13698 (I235120,I235454,I235276);
nor I_13699 (I235502,I151695,I151695);
and I_13700 (I235519,I235367,I235502);
nor I_13701 (I235536,I235454,I235519);
DFFARX1 I_13702 (I235536,I2595,I235143,I235129,);
nor I_13703 (I235567,I235169,I235502);
DFFARX1 I_13704 (I235567,I2595,I235143,I235114,);
nor I_13705 (I235598,I235446,I235502);
not I_13706 (I235615,I235598);
nand I_13707 (I235123,I235615,I235471);
not I_13708 (I235670,I2602);
DFFARX1 I_13709 (I194586,I2595,I235670,I235696,);
not I_13710 (I235704,I235696);
nand I_13711 (I235721,I194589,I194586);
and I_13712 (I235738,I235721,I194598);
DFFARX1 I_13713 (I235738,I2595,I235670,I235764,);
DFFARX1 I_13714 (I235764,I2595,I235670,I235659,);
DFFARX1 I_13715 (I194595,I2595,I235670,I235795,);
nand I_13716 (I235803,I235795,I194601);
not I_13717 (I235820,I235803);
DFFARX1 I_13718 (I235820,I2595,I235670,I235846,);
not I_13719 (I235854,I235846);
nor I_13720 (I235662,I235704,I235854);
DFFARX1 I_13721 (I194610,I2595,I235670,I235894,);
nor I_13722 (I235653,I235894,I235764);
nor I_13723 (I235644,I235894,I235820);
nand I_13724 (I235930,I194604,I194592);
and I_13725 (I235947,I235930,I194589);
DFFARX1 I_13726 (I235947,I2595,I235670,I235973,);
not I_13727 (I235981,I235973);
nand I_13728 (I235998,I235981,I235894);
nand I_13729 (I235647,I235981,I235803);
nor I_13730 (I236029,I194607,I194592);
and I_13731 (I236046,I235894,I236029);
nor I_13732 (I236063,I235981,I236046);
DFFARX1 I_13733 (I236063,I2595,I235670,I235656,);
nor I_13734 (I236094,I235696,I236029);
DFFARX1 I_13735 (I236094,I2595,I235670,I235641,);
nor I_13736 (I236125,I235973,I236029);
not I_13737 (I236142,I236125);
nand I_13738 (I235650,I236142,I235998);
not I_13739 (I236197,I2602);
DFFARX1 I_13740 (I224642,I2595,I236197,I236223,);
not I_13741 (I236231,I236223);
nand I_13742 (I236248,I224645,I224642);
and I_13743 (I236265,I236248,I224654);
DFFARX1 I_13744 (I236265,I2595,I236197,I236291,);
DFFARX1 I_13745 (I236291,I2595,I236197,I236186,);
DFFARX1 I_13746 (I224651,I2595,I236197,I236322,);
nand I_13747 (I236330,I236322,I224657);
not I_13748 (I236347,I236330);
DFFARX1 I_13749 (I236347,I2595,I236197,I236373,);
not I_13750 (I236381,I236373);
nor I_13751 (I236189,I236231,I236381);
DFFARX1 I_13752 (I224666,I2595,I236197,I236421,);
nor I_13753 (I236180,I236421,I236291);
nor I_13754 (I236171,I236421,I236347);
nand I_13755 (I236457,I224660,I224648);
and I_13756 (I236474,I236457,I224645);
DFFARX1 I_13757 (I236474,I2595,I236197,I236500,);
not I_13758 (I236508,I236500);
nand I_13759 (I236525,I236508,I236421);
nand I_13760 (I236174,I236508,I236330);
nor I_13761 (I236556,I224663,I224648);
and I_13762 (I236573,I236421,I236556);
nor I_13763 (I236590,I236508,I236573);
DFFARX1 I_13764 (I236590,I2595,I236197,I236183,);
nor I_13765 (I236621,I236223,I236556);
DFFARX1 I_13766 (I236621,I2595,I236197,I236168,);
nor I_13767 (I236652,I236500,I236556);
not I_13768 (I236669,I236652);
nand I_13769 (I236177,I236669,I236525);
not I_13770 (I236724,I2602);
DFFARX1 I_13771 (I158187,I2595,I236724,I236750,);
not I_13772 (I236758,I236750);
nand I_13773 (I236775,I158172,I158193);
and I_13774 (I236792,I236775,I158181);
DFFARX1 I_13775 (I236792,I2595,I236724,I236818,);
DFFARX1 I_13776 (I236818,I2595,I236724,I236713,);
DFFARX1 I_13777 (I158175,I2595,I236724,I236849,);
nand I_13778 (I236857,I236849,I158184);
not I_13779 (I236874,I236857);
DFFARX1 I_13780 (I236874,I2595,I236724,I236900,);
not I_13781 (I236908,I236900);
nor I_13782 (I236716,I236758,I236908);
DFFARX1 I_13783 (I158190,I2595,I236724,I236948,);
nor I_13784 (I236707,I236948,I236818);
nor I_13785 (I236698,I236948,I236874);
nand I_13786 (I236984,I158172,I158175);
and I_13787 (I237001,I236984,I158196);
DFFARX1 I_13788 (I237001,I2595,I236724,I237027,);
not I_13789 (I237035,I237027);
nand I_13790 (I237052,I237035,I236948);
nand I_13791 (I236701,I237035,I236857);
nor I_13792 (I237083,I158178,I158175);
and I_13793 (I237100,I236948,I237083);
nor I_13794 (I237117,I237035,I237100);
DFFARX1 I_13795 (I237117,I2595,I236724,I236710,);
nor I_13796 (I237148,I236750,I237083);
DFFARX1 I_13797 (I237148,I2595,I236724,I236695,);
nor I_13798 (I237179,I237027,I237083);
not I_13799 (I237196,I237179);
nand I_13800 (I236704,I237196,I237052);
not I_13801 (I237251,I2602);
DFFARX1 I_13802 (I60989,I2595,I237251,I237277,);
not I_13803 (I237285,I237277);
nand I_13804 (I237302,I60986,I61004);
and I_13805 (I237319,I237302,I60995);
DFFARX1 I_13806 (I237319,I2595,I237251,I237345,);
DFFARX1 I_13807 (I237345,I2595,I237251,I237240,);
DFFARX1 I_13808 (I61001,I2595,I237251,I237376,);
nand I_13809 (I237384,I237376,I60998);
not I_13810 (I237401,I237384);
DFFARX1 I_13811 (I237401,I2595,I237251,I237427,);
not I_13812 (I237435,I237427);
nor I_13813 (I237243,I237285,I237435);
DFFARX1 I_13814 (I60992,I2595,I237251,I237475,);
nor I_13815 (I237234,I237475,I237345);
nor I_13816 (I237225,I237475,I237401);
nand I_13817 (I237511,I60983,I61007);
and I_13818 (I237528,I237511,I60986);
DFFARX1 I_13819 (I237528,I2595,I237251,I237554,);
not I_13820 (I237562,I237554);
nand I_13821 (I237579,I237562,I237475);
nand I_13822 (I237228,I237562,I237384);
nor I_13823 (I237610,I60983,I61007);
and I_13824 (I237627,I237475,I237610);
nor I_13825 (I237644,I237562,I237627);
DFFARX1 I_13826 (I237644,I2595,I237251,I237237,);
nor I_13827 (I237675,I237277,I237610);
DFFARX1 I_13828 (I237675,I2595,I237251,I237222,);
nor I_13829 (I237706,I237554,I237610);
not I_13830 (I237723,I237706);
nand I_13831 (I237231,I237723,I237579);
not I_13832 (I237778,I2602);
DFFARX1 I_13833 (I261552,I2595,I237778,I237804,);
not I_13834 (I237812,I237804);
nand I_13835 (I237829,I261567,I261549);
and I_13836 (I237846,I237829,I261549);
DFFARX1 I_13837 (I237846,I2595,I237778,I237872,);
DFFARX1 I_13838 (I237872,I2595,I237778,I237767,);
DFFARX1 I_13839 (I261558,I2595,I237778,I237903,);
nand I_13840 (I237911,I237903,I261576);
not I_13841 (I237928,I237911);
DFFARX1 I_13842 (I237928,I2595,I237778,I237954,);
not I_13843 (I237962,I237954);
nor I_13844 (I237770,I237812,I237962);
DFFARX1 I_13845 (I261573,I2595,I237778,I238002,);
nor I_13846 (I237761,I238002,I237872);
nor I_13847 (I237752,I238002,I237928);
nand I_13848 (I238038,I261570,I261561);
and I_13849 (I238055,I238038,I261555);
DFFARX1 I_13850 (I238055,I2595,I237778,I238081,);
not I_13851 (I238089,I238081);
nand I_13852 (I238106,I238089,I238002);
nand I_13853 (I237755,I238089,I237911);
nor I_13854 (I238137,I261564,I261561);
and I_13855 (I238154,I238002,I238137);
nor I_13856 (I238171,I238089,I238154);
DFFARX1 I_13857 (I238171,I2595,I237778,I237764,);
nor I_13858 (I238202,I237804,I238137);
DFFARX1 I_13859 (I238202,I2595,I237778,I237749,);
nor I_13860 (I238233,I238081,I238137);
not I_13861 (I238250,I238233);
nand I_13862 (I237758,I238250,I238106);
not I_13863 (I238305,I2602);
DFFARX1 I_13864 (I76459,I2595,I238305,I238331,);
not I_13865 (I238339,I238331);
nand I_13866 (I238356,I76456,I76474);
and I_13867 (I238373,I238356,I76465);
DFFARX1 I_13868 (I238373,I2595,I238305,I238399,);
DFFARX1 I_13869 (I238399,I2595,I238305,I238294,);
DFFARX1 I_13870 (I76471,I2595,I238305,I238430,);
nand I_13871 (I238438,I238430,I76468);
not I_13872 (I238455,I238438);
DFFARX1 I_13873 (I238455,I2595,I238305,I238481,);
not I_13874 (I238489,I238481);
nor I_13875 (I238297,I238339,I238489);
DFFARX1 I_13876 (I76462,I2595,I238305,I238529,);
nor I_13877 (I238288,I238529,I238399);
nor I_13878 (I238279,I238529,I238455);
nand I_13879 (I238565,I76453,I76477);
and I_13880 (I238582,I238565,I76456);
DFFARX1 I_13881 (I238582,I2595,I238305,I238608,);
not I_13882 (I238616,I238608);
nand I_13883 (I238633,I238616,I238529);
nand I_13884 (I238282,I238616,I238438);
nor I_13885 (I238664,I76453,I76477);
and I_13886 (I238681,I238529,I238664);
nor I_13887 (I238698,I238616,I238681);
DFFARX1 I_13888 (I238698,I2595,I238305,I238291,);
nor I_13889 (I238729,I238331,I238664);
DFFARX1 I_13890 (I238729,I2595,I238305,I238276,);
nor I_13891 (I238760,I238608,I238664);
not I_13892 (I238777,I238760);
nand I_13893 (I238285,I238777,I238633);
not I_13894 (I238832,I2602);
DFFARX1 I_13895 (I296629,I2595,I238832,I238858,);
not I_13896 (I238866,I238858);
nand I_13897 (I238883,I296638,I296626);
and I_13898 (I238900,I238883,I296623);
DFFARX1 I_13899 (I238900,I2595,I238832,I238926,);
DFFARX1 I_13900 (I238926,I2595,I238832,I238821,);
DFFARX1 I_13901 (I296623,I2595,I238832,I238957,);
nand I_13902 (I238965,I238957,I296620);
not I_13903 (I238982,I238965);
DFFARX1 I_13904 (I238982,I2595,I238832,I239008,);
not I_13905 (I239016,I239008);
nor I_13906 (I238824,I238866,I239016);
DFFARX1 I_13907 (I296626,I2595,I238832,I239056,);
nor I_13908 (I238815,I239056,I238926);
nor I_13909 (I238806,I239056,I238982);
nand I_13910 (I239092,I296641,I296632);
and I_13911 (I239109,I239092,I296635);
DFFARX1 I_13912 (I239109,I2595,I238832,I239135,);
not I_13913 (I239143,I239135);
nand I_13914 (I239160,I239143,I239056);
nand I_13915 (I238809,I239143,I238965);
nor I_13916 (I239191,I296620,I296632);
and I_13917 (I239208,I239056,I239191);
nor I_13918 (I239225,I239143,I239208);
DFFARX1 I_13919 (I239225,I2595,I238832,I238818,);
nor I_13920 (I239256,I238858,I239191);
DFFARX1 I_13921 (I239256,I2595,I238832,I238803,);
nor I_13922 (I239287,I239135,I239191);
not I_13923 (I239304,I239287);
nand I_13924 (I238812,I239304,I239160);
not I_13925 (I239359,I2602);
DFFARX1 I_13926 (I213082,I2595,I239359,I239385,);
not I_13927 (I239393,I239385);
nand I_13928 (I239410,I213085,I213082);
and I_13929 (I239427,I239410,I213094);
DFFARX1 I_13930 (I239427,I2595,I239359,I239453,);
DFFARX1 I_13931 (I239453,I2595,I239359,I239348,);
DFFARX1 I_13932 (I213091,I2595,I239359,I239484,);
nand I_13933 (I239492,I239484,I213097);
not I_13934 (I239509,I239492);
DFFARX1 I_13935 (I239509,I2595,I239359,I239535,);
not I_13936 (I239543,I239535);
nor I_13937 (I239351,I239393,I239543);
DFFARX1 I_13938 (I213106,I2595,I239359,I239583,);
nor I_13939 (I239342,I239583,I239453);
nor I_13940 (I239333,I239583,I239509);
nand I_13941 (I239619,I213100,I213088);
and I_13942 (I239636,I239619,I213085);
DFFARX1 I_13943 (I239636,I2595,I239359,I239662,);
not I_13944 (I239670,I239662);
nand I_13945 (I239687,I239670,I239583);
nand I_13946 (I239336,I239670,I239492);
nor I_13947 (I239718,I213103,I213088);
and I_13948 (I239735,I239583,I239718);
nor I_13949 (I239752,I239670,I239735);
DFFARX1 I_13950 (I239752,I2595,I239359,I239345,);
nor I_13951 (I239783,I239385,I239718);
DFFARX1 I_13952 (I239783,I2595,I239359,I239330,);
nor I_13953 (I239814,I239662,I239718);
not I_13954 (I239831,I239814);
nand I_13955 (I239339,I239831,I239687);
not I_13956 (I239886,I2602);
DFFARX1 I_13957 (I221174,I2595,I239886,I239912,);
not I_13958 (I239920,I239912);
nand I_13959 (I239937,I221177,I221174);
and I_13960 (I239954,I239937,I221186);
DFFARX1 I_13961 (I239954,I2595,I239886,I239980,);
DFFARX1 I_13962 (I239980,I2595,I239886,I239875,);
DFFARX1 I_13963 (I221183,I2595,I239886,I240011,);
nand I_13964 (I240019,I240011,I221189);
not I_13965 (I240036,I240019);
DFFARX1 I_13966 (I240036,I2595,I239886,I240062,);
not I_13967 (I240070,I240062);
nor I_13968 (I239878,I239920,I240070);
DFFARX1 I_13969 (I221198,I2595,I239886,I240110,);
nor I_13970 (I239869,I240110,I239980);
nor I_13971 (I239860,I240110,I240036);
nand I_13972 (I240146,I221192,I221180);
and I_13973 (I240163,I240146,I221177);
DFFARX1 I_13974 (I240163,I2595,I239886,I240189,);
not I_13975 (I240197,I240189);
nand I_13976 (I240214,I240197,I240110);
nand I_13977 (I239863,I240197,I240019);
nor I_13978 (I240245,I221195,I221180);
and I_13979 (I240262,I240110,I240245);
nor I_13980 (I240279,I240197,I240262);
DFFARX1 I_13981 (I240279,I2595,I239886,I239872,);
nor I_13982 (I240310,I239912,I240245);
DFFARX1 I_13983 (I240310,I2595,I239886,I239857,);
nor I_13984 (I240341,I240189,I240245);
not I_13985 (I240358,I240341);
nand I_13986 (I239866,I240358,I240214);
not I_13987 (I240413,I2602);
DFFARX1 I_13988 (I322376,I2595,I240413,I240439,);
not I_13989 (I240447,I240439);
nand I_13990 (I240464,I322358,I322358);
and I_13991 (I240481,I240464,I322364);
DFFARX1 I_13992 (I240481,I2595,I240413,I240507,);
DFFARX1 I_13993 (I240507,I2595,I240413,I240402,);
DFFARX1 I_13994 (I322361,I2595,I240413,I240538,);
nand I_13995 (I240546,I240538,I322370);
not I_13996 (I240563,I240546);
DFFARX1 I_13997 (I240563,I2595,I240413,I240589,);
not I_13998 (I240597,I240589);
nor I_13999 (I240405,I240447,I240597);
DFFARX1 I_14000 (I322382,I2595,I240413,I240637,);
nor I_14001 (I240396,I240637,I240507);
nor I_14002 (I240387,I240637,I240563);
nand I_14003 (I240673,I322373,I322367);
and I_14004 (I240690,I240673,I322361);
DFFARX1 I_14005 (I240690,I2595,I240413,I240716,);
not I_14006 (I240724,I240716);
nand I_14007 (I240741,I240724,I240637);
nand I_14008 (I240390,I240724,I240546);
nor I_14009 (I240772,I322379,I322367);
and I_14010 (I240789,I240637,I240772);
nor I_14011 (I240806,I240724,I240789);
DFFARX1 I_14012 (I240806,I2595,I240413,I240399,);
nor I_14013 (I240837,I240439,I240772);
DFFARX1 I_14014 (I240837,I2595,I240413,I240384,);
nor I_14015 (I240868,I240716,I240772);
not I_14016 (I240885,I240868);
nand I_14017 (I240393,I240885,I240741);
not I_14018 (I240940,I2602);
DFFARX1 I_14019 (I32430,I2595,I240940,I240966,);
not I_14020 (I240974,I240966);
nand I_14021 (I240991,I32406,I32415);
and I_14022 (I241008,I240991,I32409);
DFFARX1 I_14023 (I241008,I2595,I240940,I241034,);
DFFARX1 I_14024 (I241034,I2595,I240940,I240929,);
DFFARX1 I_14025 (I32427,I2595,I240940,I241065,);
nand I_14026 (I241073,I241065,I32418);
not I_14027 (I241090,I241073);
DFFARX1 I_14028 (I241090,I2595,I240940,I241116,);
not I_14029 (I241124,I241116);
nor I_14030 (I240932,I240974,I241124);
DFFARX1 I_14031 (I32412,I2595,I240940,I241164,);
nor I_14032 (I240923,I241164,I241034);
nor I_14033 (I240914,I241164,I241090);
nand I_14034 (I241200,I32424,I32421);
and I_14035 (I241217,I241200,I32409);
DFFARX1 I_14036 (I241217,I2595,I240940,I241243,);
not I_14037 (I241251,I241243);
nand I_14038 (I241268,I241251,I241164);
nand I_14039 (I240917,I241251,I241073);
nor I_14040 (I241299,I32406,I32421);
and I_14041 (I241316,I241164,I241299);
nor I_14042 (I241333,I241251,I241316);
DFFARX1 I_14043 (I241333,I2595,I240940,I240926,);
nor I_14044 (I241364,I240966,I241299);
DFFARX1 I_14045 (I241364,I2595,I240940,I240911,);
nor I_14046 (I241395,I241243,I241299);
not I_14047 (I241412,I241395);
nand I_14048 (I240920,I241412,I241268);
not I_14049 (I241467,I2602);
DFFARX1 I_14050 (I313128,I2595,I241467,I241493,);
not I_14051 (I241501,I241493);
nand I_14052 (I241518,I313110,I313110);
and I_14053 (I241535,I241518,I313116);
DFFARX1 I_14054 (I241535,I2595,I241467,I241561,);
DFFARX1 I_14055 (I241561,I2595,I241467,I241456,);
DFFARX1 I_14056 (I313113,I2595,I241467,I241592,);
nand I_14057 (I241600,I241592,I313122);
not I_14058 (I241617,I241600);
DFFARX1 I_14059 (I241617,I2595,I241467,I241643,);
not I_14060 (I241651,I241643);
nor I_14061 (I241459,I241501,I241651);
DFFARX1 I_14062 (I313134,I2595,I241467,I241691,);
nor I_14063 (I241450,I241691,I241561);
nor I_14064 (I241441,I241691,I241617);
nand I_14065 (I241727,I313125,I313119);
and I_14066 (I241744,I241727,I313113);
DFFARX1 I_14067 (I241744,I2595,I241467,I241770,);
not I_14068 (I241778,I241770);
nand I_14069 (I241795,I241778,I241691);
nand I_14070 (I241444,I241778,I241600);
nor I_14071 (I241826,I313131,I313119);
and I_14072 (I241843,I241691,I241826);
nor I_14073 (I241860,I241778,I241843);
DFFARX1 I_14074 (I241860,I2595,I241467,I241453,);
nor I_14075 (I241891,I241493,I241826);
DFFARX1 I_14076 (I241891,I2595,I241467,I241438,);
nor I_14077 (I241922,I241770,I241826);
not I_14078 (I241939,I241922);
nand I_14079 (I241447,I241939,I241795);
not I_14080 (I241994,I2602);
DFFARX1 I_14081 (I374733,I2595,I241994,I242020,);
not I_14082 (I242028,I242020);
nand I_14083 (I242045,I374730,I374739);
and I_14084 (I242062,I242045,I374718);
DFFARX1 I_14085 (I242062,I2595,I241994,I242088,);
DFFARX1 I_14086 (I242088,I2595,I241994,I241983,);
DFFARX1 I_14087 (I374721,I2595,I241994,I242119,);
nand I_14088 (I242127,I242119,I374736);
not I_14089 (I242144,I242127);
DFFARX1 I_14090 (I242144,I2595,I241994,I242170,);
not I_14091 (I242178,I242170);
nor I_14092 (I241986,I242028,I242178);
DFFARX1 I_14093 (I374742,I2595,I241994,I242218,);
nor I_14094 (I241977,I242218,I242088);
nor I_14095 (I241968,I242218,I242144);
nand I_14096 (I242254,I374724,I374745);
and I_14097 (I242271,I242254,I374727);
DFFARX1 I_14098 (I242271,I2595,I241994,I242297,);
not I_14099 (I242305,I242297);
nand I_14100 (I242322,I242305,I242218);
nand I_14101 (I241971,I242305,I242127);
nor I_14102 (I242353,I374718,I374745);
and I_14103 (I242370,I242218,I242353);
nor I_14104 (I242387,I242305,I242370);
DFFARX1 I_14105 (I242387,I2595,I241994,I241980,);
nor I_14106 (I242418,I242020,I242353);
DFFARX1 I_14107 (I242418,I2595,I241994,I241965,);
nor I_14108 (I242449,I242297,I242353);
not I_14109 (I242466,I242449);
nand I_14110 (I241974,I242466,I242322);
not I_14111 (I242521,I2602);
DFFARX1 I_14112 (I192274,I2595,I242521,I242547,);
not I_14113 (I242555,I242547);
nand I_14114 (I242572,I192277,I192274);
and I_14115 (I242589,I242572,I192286);
DFFARX1 I_14116 (I242589,I2595,I242521,I242615,);
DFFARX1 I_14117 (I242615,I2595,I242521,I242510,);
DFFARX1 I_14118 (I192283,I2595,I242521,I242646,);
nand I_14119 (I242654,I242646,I192289);
not I_14120 (I242671,I242654);
DFFARX1 I_14121 (I242671,I2595,I242521,I242697,);
not I_14122 (I242705,I242697);
nor I_14123 (I242513,I242555,I242705);
DFFARX1 I_14124 (I192298,I2595,I242521,I242745,);
nor I_14125 (I242504,I242745,I242615);
nor I_14126 (I242495,I242745,I242671);
nand I_14127 (I242781,I192292,I192280);
and I_14128 (I242798,I242781,I192277);
DFFARX1 I_14129 (I242798,I2595,I242521,I242824,);
not I_14130 (I242832,I242824);
nand I_14131 (I242849,I242832,I242745);
nand I_14132 (I242498,I242832,I242654);
nor I_14133 (I242880,I192295,I192280);
and I_14134 (I242897,I242745,I242880);
nor I_14135 (I242914,I242832,I242897);
DFFARX1 I_14136 (I242914,I2595,I242521,I242507,);
nor I_14137 (I242945,I242547,I242880);
DFFARX1 I_14138 (I242945,I2595,I242521,I242492,);
nor I_14139 (I242976,I242824,I242880);
not I_14140 (I242993,I242976);
nand I_14141 (I242501,I242993,I242849);
not I_14142 (I243048,I2602);
DFFARX1 I_14143 (I376518,I2595,I243048,I243074,);
not I_14144 (I243082,I243074);
nand I_14145 (I243099,I376515,I376524);
and I_14146 (I243116,I243099,I376503);
DFFARX1 I_14147 (I243116,I2595,I243048,I243142,);
DFFARX1 I_14148 (I243142,I2595,I243048,I243037,);
DFFARX1 I_14149 (I376506,I2595,I243048,I243173,);
nand I_14150 (I243181,I243173,I376521);
not I_14151 (I243198,I243181);
DFFARX1 I_14152 (I243198,I2595,I243048,I243224,);
not I_14153 (I243232,I243224);
nor I_14154 (I243040,I243082,I243232);
DFFARX1 I_14155 (I376527,I2595,I243048,I243272,);
nor I_14156 (I243031,I243272,I243142);
nor I_14157 (I243022,I243272,I243198);
nand I_14158 (I243308,I376509,I376530);
and I_14159 (I243325,I243308,I376512);
DFFARX1 I_14160 (I243325,I2595,I243048,I243351,);
not I_14161 (I243359,I243351);
nand I_14162 (I243376,I243359,I243272);
nand I_14163 (I243025,I243359,I243181);
nor I_14164 (I243407,I376503,I376530);
and I_14165 (I243424,I243272,I243407);
nor I_14166 (I243441,I243359,I243424);
DFFARX1 I_14167 (I243441,I2595,I243048,I243034,);
nor I_14168 (I243472,I243074,I243407);
DFFARX1 I_14169 (I243472,I2595,I243048,I243019,);
nor I_14170 (I243503,I243351,I243407);
not I_14171 (I243520,I243503);
nand I_14172 (I243028,I243520,I243376);
not I_14173 (I243575,I2602);
DFFARX1 I_14174 (I214816,I2595,I243575,I243601,);
not I_14175 (I243609,I243601);
nand I_14176 (I243626,I214819,I214816);
and I_14177 (I243643,I243626,I214828);
DFFARX1 I_14178 (I243643,I2595,I243575,I243669,);
DFFARX1 I_14179 (I243669,I2595,I243575,I243564,);
DFFARX1 I_14180 (I214825,I2595,I243575,I243700,);
nand I_14181 (I243708,I243700,I214831);
not I_14182 (I243725,I243708);
DFFARX1 I_14183 (I243725,I2595,I243575,I243751,);
not I_14184 (I243759,I243751);
nor I_14185 (I243567,I243609,I243759);
DFFARX1 I_14186 (I214840,I2595,I243575,I243799,);
nor I_14187 (I243558,I243799,I243669);
nor I_14188 (I243549,I243799,I243725);
nand I_14189 (I243835,I214834,I214822);
and I_14190 (I243852,I243835,I214819);
DFFARX1 I_14191 (I243852,I2595,I243575,I243878,);
not I_14192 (I243886,I243878);
nand I_14193 (I243903,I243886,I243799);
nand I_14194 (I243552,I243886,I243708);
nor I_14195 (I243934,I214837,I214822);
and I_14196 (I243951,I243799,I243934);
nor I_14197 (I243968,I243886,I243951);
DFFARX1 I_14198 (I243968,I2595,I243575,I243561,);
nor I_14199 (I243999,I243601,I243934);
DFFARX1 I_14200 (I243999,I2595,I243575,I243546,);
nor I_14201 (I244030,I243878,I243934);
not I_14202 (I244047,I244030);
nand I_14203 (I243555,I244047,I243903);
not I_14204 (I244102,I2602);
DFFARX1 I_14205 (I301117,I2595,I244102,I244128,);
not I_14206 (I244136,I244128);
nand I_14207 (I244153,I301126,I301114);
and I_14208 (I244170,I244153,I301111);
DFFARX1 I_14209 (I244170,I2595,I244102,I244196,);
DFFARX1 I_14210 (I244196,I2595,I244102,I244091,);
DFFARX1 I_14211 (I301111,I2595,I244102,I244227,);
nand I_14212 (I244235,I244227,I301108);
not I_14213 (I244252,I244235);
DFFARX1 I_14214 (I244252,I2595,I244102,I244278,);
not I_14215 (I244286,I244278);
nor I_14216 (I244094,I244136,I244286);
DFFARX1 I_14217 (I301114,I2595,I244102,I244326,);
nor I_14218 (I244085,I244326,I244196);
nor I_14219 (I244076,I244326,I244252);
nand I_14220 (I244362,I301129,I301120);
and I_14221 (I244379,I244362,I301123);
DFFARX1 I_14222 (I244379,I2595,I244102,I244405,);
not I_14223 (I244413,I244405);
nand I_14224 (I244430,I244413,I244326);
nand I_14225 (I244079,I244413,I244235);
nor I_14226 (I244461,I301108,I301120);
and I_14227 (I244478,I244326,I244461);
nor I_14228 (I244495,I244413,I244478);
DFFARX1 I_14229 (I244495,I2595,I244102,I244088,);
nor I_14230 (I244526,I244128,I244461);
DFFARX1 I_14231 (I244526,I2595,I244102,I244073,);
nor I_14232 (I244557,I244405,I244461);
not I_14233 (I244574,I244557);
nand I_14234 (I244082,I244574,I244430);
not I_14235 (I244629,I2602);
DFFARX1 I_14236 (I157609,I2595,I244629,I244655,);
not I_14237 (I244663,I244655);
nand I_14238 (I244680,I157594,I157615);
and I_14239 (I244697,I244680,I157603);
DFFARX1 I_14240 (I244697,I2595,I244629,I244723,);
DFFARX1 I_14241 (I244723,I2595,I244629,I244618,);
DFFARX1 I_14242 (I157597,I2595,I244629,I244754,);
nand I_14243 (I244762,I244754,I157606);
not I_14244 (I244779,I244762);
DFFARX1 I_14245 (I244779,I2595,I244629,I244805,);
not I_14246 (I244813,I244805);
nor I_14247 (I244621,I244663,I244813);
DFFARX1 I_14248 (I157612,I2595,I244629,I244853,);
nor I_14249 (I244612,I244853,I244723);
nor I_14250 (I244603,I244853,I244779);
nand I_14251 (I244889,I157594,I157597);
and I_14252 (I244906,I244889,I157618);
DFFARX1 I_14253 (I244906,I2595,I244629,I244932,);
not I_14254 (I244940,I244932);
nand I_14255 (I244957,I244940,I244853);
nand I_14256 (I244606,I244940,I244762);
nor I_14257 (I244988,I157600,I157597);
and I_14258 (I245005,I244853,I244988);
nor I_14259 (I245022,I244940,I245005);
DFFARX1 I_14260 (I245022,I2595,I244629,I244615,);
nor I_14261 (I245053,I244655,I244988);
DFFARX1 I_14262 (I245053,I2595,I244629,I244600,);
nor I_14263 (I245084,I244932,I244988);
not I_14264 (I245101,I245084);
nand I_14265 (I244609,I245101,I244957);
not I_14266 (I245156,I2602);
DFFARX1 I_14267 (I172637,I2595,I245156,I245182,);
not I_14268 (I245190,I245182);
nand I_14269 (I245207,I172622,I172643);
and I_14270 (I245224,I245207,I172631);
DFFARX1 I_14271 (I245224,I2595,I245156,I245250,);
DFFARX1 I_14272 (I245250,I2595,I245156,I245145,);
DFFARX1 I_14273 (I172625,I2595,I245156,I245281,);
nand I_14274 (I245289,I245281,I172634);
not I_14275 (I245306,I245289);
DFFARX1 I_14276 (I245306,I2595,I245156,I245332,);
not I_14277 (I245340,I245332);
nor I_14278 (I245148,I245190,I245340);
DFFARX1 I_14279 (I172640,I2595,I245156,I245380,);
nor I_14280 (I245139,I245380,I245250);
nor I_14281 (I245130,I245380,I245306);
nand I_14282 (I245416,I172622,I172625);
and I_14283 (I245433,I245416,I172646);
DFFARX1 I_14284 (I245433,I2595,I245156,I245459,);
not I_14285 (I245467,I245459);
nand I_14286 (I245484,I245467,I245380);
nand I_14287 (I245133,I245467,I245289);
nor I_14288 (I245515,I172628,I172625);
and I_14289 (I245532,I245380,I245515);
nor I_14290 (I245549,I245467,I245532);
DFFARX1 I_14291 (I245549,I2595,I245156,I245142,);
nor I_14292 (I245580,I245182,I245515);
DFFARX1 I_14293 (I245580,I2595,I245156,I245127,);
nor I_14294 (I245611,I245459,I245515);
not I_14295 (I245628,I245611);
nand I_14296 (I245136,I245628,I245484);
not I_14297 (I245683,I2602);
DFFARX1 I_14298 (I314284,I2595,I245683,I245709,);
not I_14299 (I245717,I245709);
nand I_14300 (I245734,I314266,I314266);
and I_14301 (I245751,I245734,I314272);
DFFARX1 I_14302 (I245751,I2595,I245683,I245777,);
DFFARX1 I_14303 (I245777,I2595,I245683,I245672,);
DFFARX1 I_14304 (I314269,I2595,I245683,I245808,);
nand I_14305 (I245816,I245808,I314278);
not I_14306 (I245833,I245816);
DFFARX1 I_14307 (I245833,I2595,I245683,I245859,);
not I_14308 (I245867,I245859);
nor I_14309 (I245675,I245717,I245867);
DFFARX1 I_14310 (I314290,I2595,I245683,I245907,);
nor I_14311 (I245666,I245907,I245777);
nor I_14312 (I245657,I245907,I245833);
nand I_14313 (I245943,I314281,I314275);
and I_14314 (I245960,I245943,I314269);
DFFARX1 I_14315 (I245960,I2595,I245683,I245986,);
not I_14316 (I245994,I245986);
nand I_14317 (I246011,I245994,I245907);
nand I_14318 (I245660,I245994,I245816);
nor I_14319 (I246042,I314287,I314275);
and I_14320 (I246059,I245907,I246042);
nor I_14321 (I246076,I245994,I246059);
DFFARX1 I_14322 (I246076,I2595,I245683,I245669,);
nor I_14323 (I246107,I245709,I246042);
DFFARX1 I_14324 (I246107,I2595,I245683,I245654,);
nor I_14325 (I246138,I245986,I246042);
not I_14326 (I246155,I246138);
nand I_14327 (I245663,I246155,I246011);
not I_14328 (I246210,I2602);
DFFARX1 I_14329 (I330468,I2595,I246210,I246236,);
not I_14330 (I246244,I246236);
nand I_14331 (I246261,I330450,I330450);
and I_14332 (I246278,I246261,I330456);
DFFARX1 I_14333 (I246278,I2595,I246210,I246304,);
DFFARX1 I_14334 (I246304,I2595,I246210,I246199,);
DFFARX1 I_14335 (I330453,I2595,I246210,I246335,);
nand I_14336 (I246343,I246335,I330462);
not I_14337 (I246360,I246343);
DFFARX1 I_14338 (I246360,I2595,I246210,I246386,);
not I_14339 (I246394,I246386);
nor I_14340 (I246202,I246244,I246394);
DFFARX1 I_14341 (I330474,I2595,I246210,I246434,);
nor I_14342 (I246193,I246434,I246304);
nor I_14343 (I246184,I246434,I246360);
nand I_14344 (I246470,I330465,I330459);
and I_14345 (I246487,I246470,I330453);
DFFARX1 I_14346 (I246487,I2595,I246210,I246513,);
not I_14347 (I246521,I246513);
nand I_14348 (I246538,I246521,I246434);
nand I_14349 (I246187,I246521,I246343);
nor I_14350 (I246569,I330471,I330459);
and I_14351 (I246586,I246434,I246569);
nor I_14352 (I246603,I246521,I246586);
DFFARX1 I_14353 (I246603,I2595,I246210,I246196,);
nor I_14354 (I246634,I246236,I246569);
DFFARX1 I_14355 (I246634,I2595,I246210,I246181,);
nor I_14356 (I246665,I246513,I246569);
not I_14357 (I246682,I246665);
nand I_14358 (I246190,I246682,I246538);
not I_14359 (I246737,I2602);
DFFARX1 I_14360 (I264136,I2595,I246737,I246763,);
not I_14361 (I246771,I246763);
nand I_14362 (I246788,I264151,I264133);
and I_14363 (I246805,I246788,I264133);
DFFARX1 I_14364 (I246805,I2595,I246737,I246831,);
DFFARX1 I_14365 (I246831,I2595,I246737,I246726,);
DFFARX1 I_14366 (I264142,I2595,I246737,I246862,);
nand I_14367 (I246870,I246862,I264160);
not I_14368 (I246887,I246870);
DFFARX1 I_14369 (I246887,I2595,I246737,I246913,);
not I_14370 (I246921,I246913);
nor I_14371 (I246729,I246771,I246921);
DFFARX1 I_14372 (I264157,I2595,I246737,I246961,);
nor I_14373 (I246720,I246961,I246831);
nor I_14374 (I246711,I246961,I246887);
nand I_14375 (I246997,I264154,I264145);
and I_14376 (I247014,I246997,I264139);
DFFARX1 I_14377 (I247014,I2595,I246737,I247040,);
not I_14378 (I247048,I247040);
nand I_14379 (I247065,I247048,I246961);
nand I_14380 (I246714,I247048,I246870);
nor I_14381 (I247096,I264148,I264145);
and I_14382 (I247113,I246961,I247096);
nor I_14383 (I247130,I247048,I247113);
DFFARX1 I_14384 (I247130,I2595,I246737,I246723,);
nor I_14385 (I247161,I246763,I247096);
DFFARX1 I_14386 (I247161,I2595,I246737,I246708,);
nor I_14387 (I247192,I247040,I247096);
not I_14388 (I247209,I247192);
nand I_14389 (I246717,I247209,I247065);
not I_14390 (I247264,I2602);
DFFARX1 I_14391 (I121407,I2595,I247264,I247290,);
not I_14392 (I247298,I247290);
nand I_14393 (I247315,I121404,I121413);
and I_14394 (I247332,I247315,I121422);
DFFARX1 I_14395 (I247332,I2595,I247264,I247358,);
DFFARX1 I_14396 (I247358,I2595,I247264,I247253,);
DFFARX1 I_14397 (I121425,I2595,I247264,I247389,);
nand I_14398 (I247397,I247389,I121428);
not I_14399 (I247414,I247397);
DFFARX1 I_14400 (I247414,I2595,I247264,I247440,);
not I_14401 (I247448,I247440);
nor I_14402 (I247256,I247298,I247448);
DFFARX1 I_14403 (I121401,I2595,I247264,I247488,);
nor I_14404 (I247247,I247488,I247358);
nor I_14405 (I247238,I247488,I247414);
nand I_14406 (I247524,I121416,I121419);
and I_14407 (I247541,I247524,I121410);
DFFARX1 I_14408 (I247541,I2595,I247264,I247567,);
not I_14409 (I247575,I247567);
nand I_14410 (I247592,I247575,I247488);
nand I_14411 (I247241,I247575,I247397);
nor I_14412 (I247623,I121401,I121419);
and I_14413 (I247640,I247488,I247623);
nor I_14414 (I247657,I247575,I247640);
DFFARX1 I_14415 (I247657,I2595,I247264,I247250,);
nor I_14416 (I247688,I247290,I247623);
DFFARX1 I_14417 (I247688,I2595,I247264,I247235,);
nor I_14418 (I247719,I247567,I247623);
not I_14419 (I247736,I247719);
nand I_14420 (I247244,I247736,I247592);
not I_14421 (I247791,I2602);
DFFARX1 I_14422 (I375923,I2595,I247791,I247817,);
not I_14423 (I247825,I247817);
nand I_14424 (I247842,I375920,I375929);
and I_14425 (I247859,I247842,I375908);
DFFARX1 I_14426 (I247859,I2595,I247791,I247885,);
DFFARX1 I_14427 (I247885,I2595,I247791,I247780,);
DFFARX1 I_14428 (I375911,I2595,I247791,I247916,);
nand I_14429 (I247924,I247916,I375926);
not I_14430 (I247941,I247924);
DFFARX1 I_14431 (I247941,I2595,I247791,I247967,);
not I_14432 (I247975,I247967);
nor I_14433 (I247783,I247825,I247975);
DFFARX1 I_14434 (I375932,I2595,I247791,I248015,);
nor I_14435 (I247774,I248015,I247885);
nor I_14436 (I247765,I248015,I247941);
nand I_14437 (I248051,I375914,I375935);
and I_14438 (I248068,I248051,I375917);
DFFARX1 I_14439 (I248068,I2595,I247791,I248094,);
not I_14440 (I248102,I248094);
nand I_14441 (I248119,I248102,I248015);
nand I_14442 (I247768,I248102,I247924);
nor I_14443 (I248150,I375908,I375935);
and I_14444 (I248167,I248015,I248150);
nor I_14445 (I248184,I248102,I248167);
DFFARX1 I_14446 (I248184,I2595,I247791,I247777,);
nor I_14447 (I248215,I247817,I248150);
DFFARX1 I_14448 (I248215,I2595,I247791,I247762,);
nor I_14449 (I248246,I248094,I248150);
not I_14450 (I248263,I248246);
nand I_14451 (I247771,I248263,I248119);
not I_14452 (I248318,I2602);
DFFARX1 I_14453 (I348074,I2595,I248318,I248344,);
not I_14454 (I248352,I248344);
nand I_14455 (I248369,I348080,I348062);
and I_14456 (I248386,I248369,I348071);
DFFARX1 I_14457 (I248386,I2595,I248318,I248412,);
DFFARX1 I_14458 (I248412,I2595,I248318,I248307,);
DFFARX1 I_14459 (I348077,I2595,I248318,I248443,);
nand I_14460 (I248451,I248443,I348065);
not I_14461 (I248468,I248451);
DFFARX1 I_14462 (I248468,I2595,I248318,I248494,);
not I_14463 (I248502,I248494);
nor I_14464 (I248310,I248352,I248502);
DFFARX1 I_14465 (I348083,I2595,I248318,I248542,);
nor I_14466 (I248301,I248542,I248412);
nor I_14467 (I248292,I248542,I248468);
nand I_14468 (I248578,I348062,I348068);
and I_14469 (I248595,I248578,I348086);
DFFARX1 I_14470 (I248595,I2595,I248318,I248621,);
not I_14471 (I248629,I248621);
nand I_14472 (I248646,I248629,I248542);
nand I_14473 (I248295,I248629,I248451);
nor I_14474 (I248677,I348065,I348068);
and I_14475 (I248694,I248542,I248677);
nor I_14476 (I248711,I248629,I248694);
DFFARX1 I_14477 (I248711,I2595,I248318,I248304,);
nor I_14478 (I248742,I248344,I248677);
DFFARX1 I_14479 (I248742,I2595,I248318,I248289,);
nor I_14480 (I248773,I248621,I248677);
not I_14481 (I248790,I248773);
nand I_14482 (I248298,I248790,I248646);
not I_14483 (I248845,I2602);
DFFARX1 I_14484 (I300556,I2595,I248845,I248871,);
not I_14485 (I248879,I248871);
nand I_14486 (I248896,I300565,I300553);
and I_14487 (I248913,I248896,I300550);
DFFARX1 I_14488 (I248913,I2595,I248845,I248939,);
DFFARX1 I_14489 (I248939,I2595,I248845,I248834,);
DFFARX1 I_14490 (I300550,I2595,I248845,I248970,);
nand I_14491 (I248978,I248970,I300547);
not I_14492 (I248995,I248978);
DFFARX1 I_14493 (I248995,I2595,I248845,I249021,);
not I_14494 (I249029,I249021);
nor I_14495 (I248837,I248879,I249029);
DFFARX1 I_14496 (I300553,I2595,I248845,I249069,);
nor I_14497 (I248828,I249069,I248939);
nor I_14498 (I248819,I249069,I248995);
nand I_14499 (I249105,I300568,I300559);
and I_14500 (I249122,I249105,I300562);
DFFARX1 I_14501 (I249122,I2595,I248845,I249148,);
not I_14502 (I249156,I249148);
nand I_14503 (I249173,I249156,I249069);
nand I_14504 (I248822,I249156,I248978);
nor I_14505 (I249204,I300547,I300559);
and I_14506 (I249221,I249069,I249204);
nor I_14507 (I249238,I249156,I249221);
DFFARX1 I_14508 (I249238,I2595,I248845,I248831,);
nor I_14509 (I249269,I248871,I249204);
DFFARX1 I_14510 (I249269,I2595,I248845,I248816,);
nor I_14511 (I249300,I249148,I249204);
not I_14512 (I249317,I249300);
nand I_14513 (I248825,I249317,I249173);
not I_14514 (I249372,I2602);
DFFARX1 I_14515 (I34011,I2595,I249372,I249398,);
not I_14516 (I249406,I249398);
nand I_14517 (I249423,I33987,I33996);
and I_14518 (I249440,I249423,I33990);
DFFARX1 I_14519 (I249440,I2595,I249372,I249466,);
DFFARX1 I_14520 (I249466,I2595,I249372,I249361,);
DFFARX1 I_14521 (I34008,I2595,I249372,I249497,);
nand I_14522 (I249505,I249497,I33999);
not I_14523 (I249522,I249505);
DFFARX1 I_14524 (I249522,I2595,I249372,I249548,);
not I_14525 (I249556,I249548);
nor I_14526 (I249364,I249406,I249556);
DFFARX1 I_14527 (I33993,I2595,I249372,I249596,);
nor I_14528 (I249355,I249596,I249466);
nor I_14529 (I249346,I249596,I249522);
nand I_14530 (I249632,I34005,I34002);
and I_14531 (I249649,I249632,I33990);
DFFARX1 I_14532 (I249649,I2595,I249372,I249675,);
not I_14533 (I249683,I249675);
nand I_14534 (I249700,I249683,I249596);
nand I_14535 (I249349,I249683,I249505);
nor I_14536 (I249731,I33987,I34002);
and I_14537 (I249748,I249596,I249731);
nor I_14538 (I249765,I249683,I249748);
DFFARX1 I_14539 (I249765,I2595,I249372,I249358,);
nor I_14540 (I249796,I249398,I249731);
DFFARX1 I_14541 (I249796,I2595,I249372,I249343,);
nor I_14542 (I249827,I249675,I249731);
not I_14543 (I249844,I249827);
nand I_14544 (I249352,I249844,I249700);
not I_14545 (I249899,I2602);
DFFARX1 I_14546 (I27160,I2595,I249899,I249925,);
not I_14547 (I249933,I249925);
nand I_14548 (I249950,I27136,I27145);
and I_14549 (I249967,I249950,I27139);
DFFARX1 I_14550 (I249967,I2595,I249899,I249993,);
DFFARX1 I_14551 (I249993,I2595,I249899,I249888,);
DFFARX1 I_14552 (I27157,I2595,I249899,I250024,);
nand I_14553 (I250032,I250024,I27148);
not I_14554 (I250049,I250032);
DFFARX1 I_14555 (I250049,I2595,I249899,I250075,);
not I_14556 (I250083,I250075);
nor I_14557 (I249891,I249933,I250083);
DFFARX1 I_14558 (I27142,I2595,I249899,I250123,);
nor I_14559 (I249882,I250123,I249993);
nor I_14560 (I249873,I250123,I250049);
nand I_14561 (I250159,I27154,I27151);
and I_14562 (I250176,I250159,I27139);
DFFARX1 I_14563 (I250176,I2595,I249899,I250202,);
not I_14564 (I250210,I250202);
nand I_14565 (I250227,I250210,I250123);
nand I_14566 (I249876,I250210,I250032);
nor I_14567 (I250258,I27136,I27151);
and I_14568 (I250275,I250123,I250258);
nor I_14569 (I250292,I250210,I250275);
DFFARX1 I_14570 (I250292,I2595,I249899,I249885,);
nor I_14571 (I250323,I249925,I250258);
DFFARX1 I_14572 (I250323,I2595,I249899,I249870,);
nor I_14573 (I250354,I250202,I250258);
not I_14574 (I250371,I250354);
nand I_14575 (I249879,I250371,I250227);
not I_14576 (I250426,I2602);
DFFARX1 I_14577 (I352970,I2595,I250426,I250452,);
not I_14578 (I250460,I250452);
nand I_14579 (I250477,I352976,I352958);
and I_14580 (I250494,I250477,I352967);
DFFARX1 I_14581 (I250494,I2595,I250426,I250520,);
DFFARX1 I_14582 (I250520,I2595,I250426,I250415,);
DFFARX1 I_14583 (I352973,I2595,I250426,I250551,);
nand I_14584 (I250559,I250551,I352961);
not I_14585 (I250576,I250559);
DFFARX1 I_14586 (I250576,I2595,I250426,I250602,);
not I_14587 (I250610,I250602);
nor I_14588 (I250418,I250460,I250610);
DFFARX1 I_14589 (I352979,I2595,I250426,I250650,);
nor I_14590 (I250409,I250650,I250520);
nor I_14591 (I250400,I250650,I250576);
nand I_14592 (I250686,I352958,I352964);
and I_14593 (I250703,I250686,I352982);
DFFARX1 I_14594 (I250703,I2595,I250426,I250729,);
not I_14595 (I250737,I250729);
nand I_14596 (I250754,I250737,I250650);
nand I_14597 (I250403,I250737,I250559);
nor I_14598 (I250785,I352961,I352964);
and I_14599 (I250802,I250650,I250785);
nor I_14600 (I250819,I250737,I250802);
DFFARX1 I_14601 (I250819,I2595,I250426,I250412,);
nor I_14602 (I250850,I250452,I250785);
DFFARX1 I_14603 (I250850,I2595,I250426,I250397,);
nor I_14604 (I250881,I250729,I250785);
not I_14605 (I250898,I250881);
nand I_14606 (I250406,I250898,I250754);
not I_14607 (I250953,I2602);
DFFARX1 I_14608 (I142776,I2595,I250953,I250979,);
not I_14609 (I250987,I250979);
nand I_14610 (I251004,I142794,I142785);
and I_14611 (I251021,I251004,I142788);
DFFARX1 I_14612 (I251021,I2595,I250953,I251047,);
DFFARX1 I_14613 (I251047,I2595,I250953,I250942,);
DFFARX1 I_14614 (I142782,I2595,I250953,I251078,);
nand I_14615 (I251086,I251078,I142773);
not I_14616 (I251103,I251086);
DFFARX1 I_14617 (I251103,I2595,I250953,I251129,);
not I_14618 (I251137,I251129);
nor I_14619 (I250945,I250987,I251137);
DFFARX1 I_14620 (I142779,I2595,I250953,I251177,);
nor I_14621 (I250936,I251177,I251047);
nor I_14622 (I250927,I251177,I251103);
nand I_14623 (I251213,I142773,I142770);
and I_14624 (I251230,I251213,I142791);
DFFARX1 I_14625 (I251230,I2595,I250953,I251256,);
not I_14626 (I251264,I251256);
nand I_14627 (I251281,I251264,I251177);
nand I_14628 (I250930,I251264,I251086);
nor I_14629 (I251312,I142770,I142770);
and I_14630 (I251329,I251177,I251312);
nor I_14631 (I251346,I251264,I251329);
DFFARX1 I_14632 (I251346,I2595,I250953,I250939,);
nor I_14633 (I251377,I250979,I251312);
DFFARX1 I_14634 (I251377,I2595,I250953,I250924,);
nor I_14635 (I251408,I251256,I251312);
not I_14636 (I251425,I251408);
nand I_14637 (I250933,I251425,I251281);
not I_14638 (I251480,I2602);
DFFARX1 I_14639 (I269304,I2595,I251480,I251506,);
not I_14640 (I251514,I251506);
nand I_14641 (I251531,I269319,I269301);
and I_14642 (I251548,I251531,I269301);
DFFARX1 I_14643 (I251548,I2595,I251480,I251574,);
DFFARX1 I_14644 (I251574,I2595,I251480,I251469,);
DFFARX1 I_14645 (I269310,I2595,I251480,I251605,);
nand I_14646 (I251613,I251605,I269328);
not I_14647 (I251630,I251613);
DFFARX1 I_14648 (I251630,I2595,I251480,I251656,);
not I_14649 (I251664,I251656);
nor I_14650 (I251472,I251514,I251664);
DFFARX1 I_14651 (I269325,I2595,I251480,I251704,);
nor I_14652 (I251463,I251704,I251574);
nor I_14653 (I251454,I251704,I251630);
nand I_14654 (I251740,I269322,I269313);
and I_14655 (I251757,I251740,I269307);
DFFARX1 I_14656 (I251757,I2595,I251480,I251783,);
not I_14657 (I251791,I251783);
nand I_14658 (I251808,I251791,I251704);
nand I_14659 (I251457,I251791,I251613);
nor I_14660 (I251839,I269316,I269313);
and I_14661 (I251856,I251704,I251839);
nor I_14662 (I251873,I251791,I251856);
DFFARX1 I_14663 (I251873,I2595,I251480,I251466,);
nor I_14664 (I251904,I251506,I251839);
DFFARX1 I_14665 (I251904,I2595,I251480,I251451,);
nor I_14666 (I251935,I251783,I251839);
not I_14667 (I251952,I251935);
nand I_14668 (I251460,I251952,I251808);
not I_14669 (I252007,I2602);
DFFARX1 I_14670 (I95910,I2595,I252007,I252033,);
not I_14671 (I252041,I252033);
nand I_14672 (I252058,I95901,I95901);
and I_14673 (I252075,I252058,I95919);
DFFARX1 I_14674 (I252075,I2595,I252007,I252101,);
DFFARX1 I_14675 (I252101,I2595,I252007,I251996,);
DFFARX1 I_14676 (I95922,I2595,I252007,I252132,);
nand I_14677 (I252140,I252132,I95904);
not I_14678 (I252157,I252140);
DFFARX1 I_14679 (I252157,I2595,I252007,I252183,);
not I_14680 (I252191,I252183);
nor I_14681 (I251999,I252041,I252191);
DFFARX1 I_14682 (I95916,I2595,I252007,I252231,);
nor I_14683 (I251990,I252231,I252101);
nor I_14684 (I251981,I252231,I252157);
nand I_14685 (I252267,I95928,I95907);
and I_14686 (I252284,I252267,I95913);
DFFARX1 I_14687 (I252284,I2595,I252007,I252310,);
not I_14688 (I252318,I252310);
nand I_14689 (I252335,I252318,I252231);
nand I_14690 (I251984,I252318,I252140);
nor I_14691 (I252366,I95925,I95907);
and I_14692 (I252383,I252231,I252366);
nor I_14693 (I252400,I252318,I252383);
DFFARX1 I_14694 (I252400,I2595,I252007,I251993,);
nor I_14695 (I252431,I252033,I252366);
DFFARX1 I_14696 (I252431,I2595,I252007,I251978,);
nor I_14697 (I252462,I252310,I252366);
not I_14698 (I252479,I252462);
nand I_14699 (I251987,I252479,I252335);
not I_14700 (I252540,I2602);
DFFARX1 I_14701 (I58014,I2595,I252540,I252566,);
DFFARX1 I_14702 (I58026,I2595,I252540,I252583,);
not I_14703 (I252591,I252583);
not I_14704 (I252608,I58032);
nor I_14705 (I252625,I252608,I58017);
not I_14706 (I252642,I58008);
nor I_14707 (I252659,I252625,I58029);
nor I_14708 (I252676,I252583,I252659);
DFFARX1 I_14709 (I252676,I2595,I252540,I252526,);
nor I_14710 (I252707,I58029,I58017);
nand I_14711 (I252724,I252707,I58032);
DFFARX1 I_14712 (I252724,I2595,I252540,I252529,);
nor I_14713 (I252755,I252642,I58029);
nand I_14714 (I252772,I252755,I58011);
nor I_14715 (I252789,I252566,I252772);
DFFARX1 I_14716 (I252789,I2595,I252540,I252505,);
not I_14717 (I252820,I252772);
nand I_14718 (I252517,I252583,I252820);
DFFARX1 I_14719 (I252772,I2595,I252540,I252860,);
not I_14720 (I252868,I252860);
not I_14721 (I252885,I58029);
not I_14722 (I252902,I58020);
nor I_14723 (I252919,I252902,I58008);
nor I_14724 (I252532,I252868,I252919);
nor I_14725 (I252950,I252902,I58023);
and I_14726 (I252967,I252950,I58011);
or I_14727 (I252984,I252967,I58008);
DFFARX1 I_14728 (I252984,I2595,I252540,I253010,);
nor I_14729 (I252520,I253010,I252566);
not I_14730 (I253032,I253010);
and I_14731 (I253049,I253032,I252566);
nor I_14732 (I252514,I252591,I253049);
nand I_14733 (I253080,I253032,I252642);
nor I_14734 (I252508,I252902,I253080);
nand I_14735 (I252511,I253032,I252820);
nand I_14736 (I253125,I252642,I58020);
nor I_14737 (I252523,I252885,I253125);
not I_14738 (I253186,I2602);
DFFARX1 I_14739 (I251457,I2595,I253186,I253212,);
DFFARX1 I_14740 (I251454,I2595,I253186,I253229,);
not I_14741 (I253237,I253229);
not I_14742 (I253254,I251454);
nor I_14743 (I253271,I253254,I251457);
not I_14744 (I253288,I251469);
nor I_14745 (I253305,I253271,I251463);
nor I_14746 (I253322,I253229,I253305);
DFFARX1 I_14747 (I253322,I2595,I253186,I253172,);
nor I_14748 (I253353,I251463,I251457);
nand I_14749 (I253370,I253353,I251454);
DFFARX1 I_14750 (I253370,I2595,I253186,I253175,);
nor I_14751 (I253401,I253288,I251463);
nand I_14752 (I253418,I253401,I251451);
nor I_14753 (I253435,I253212,I253418);
DFFARX1 I_14754 (I253435,I2595,I253186,I253151,);
not I_14755 (I253466,I253418);
nand I_14756 (I253163,I253229,I253466);
DFFARX1 I_14757 (I253418,I2595,I253186,I253506,);
not I_14758 (I253514,I253506);
not I_14759 (I253531,I251463);
not I_14760 (I253548,I251460);
nor I_14761 (I253565,I253548,I251469);
nor I_14762 (I253178,I253514,I253565);
nor I_14763 (I253596,I253548,I251466);
and I_14764 (I253613,I253596,I251472);
or I_14765 (I253630,I253613,I251451);
DFFARX1 I_14766 (I253630,I2595,I253186,I253656,);
nor I_14767 (I253166,I253656,I253212);
not I_14768 (I253678,I253656);
and I_14769 (I253695,I253678,I253212);
nor I_14770 (I253160,I253237,I253695);
nand I_14771 (I253726,I253678,I253288);
nor I_14772 (I253154,I253548,I253726);
nand I_14773 (I253157,I253678,I253466);
nand I_14774 (I253771,I253288,I251460);
nor I_14775 (I253169,I253531,I253771);
not I_14776 (I253832,I2602);
DFFARX1 I_14777 (I303352,I2595,I253832,I253858,);
DFFARX1 I_14778 (I303355,I2595,I253832,I253875,);
not I_14779 (I253883,I253875);
not I_14780 (I253900,I303352);
nor I_14781 (I253917,I253900,I303364);
not I_14782 (I253934,I303373);
nor I_14783 (I253951,I253917,I303361);
nor I_14784 (I253968,I253875,I253951);
DFFARX1 I_14785 (I253968,I2595,I253832,I253818,);
nor I_14786 (I253999,I303361,I303364);
nand I_14787 (I254016,I253999,I303352);
DFFARX1 I_14788 (I254016,I2595,I253832,I253821,);
nor I_14789 (I254047,I253934,I303361);
nand I_14790 (I254064,I254047,I303367);
nor I_14791 (I254081,I253858,I254064);
DFFARX1 I_14792 (I254081,I2595,I253832,I253797,);
not I_14793 (I254112,I254064);
nand I_14794 (I253809,I253875,I254112);
DFFARX1 I_14795 (I254064,I2595,I253832,I254152,);
not I_14796 (I254160,I254152);
not I_14797 (I254177,I303361);
not I_14798 (I254194,I303358);
nor I_14799 (I254211,I254194,I303373);
nor I_14800 (I253824,I254160,I254211);
nor I_14801 (I254242,I254194,I303370);
and I_14802 (I254259,I254242,I303358);
or I_14803 (I254276,I254259,I303355);
DFFARX1 I_14804 (I254276,I2595,I253832,I254302,);
nor I_14805 (I253812,I254302,I253858);
not I_14806 (I254324,I254302);
and I_14807 (I254341,I254324,I253858);
nor I_14808 (I253806,I253883,I254341);
nand I_14809 (I254372,I254324,I253934);
nor I_14810 (I253800,I254194,I254372);
nand I_14811 (I253803,I254324,I254112);
nand I_14812 (I254417,I253934,I303358);
nor I_14813 (I253815,I254177,I254417);
not I_14814 (I254478,I2602);
DFFARX1 I_14815 (I2228,I2595,I254478,I254504,);
DFFARX1 I_14816 (I2220,I2595,I254478,I254521,);
not I_14817 (I254529,I254521);
not I_14818 (I254546,I2428);
nor I_14819 (I254563,I254546,I1484);
not I_14820 (I254580,I1372);
nor I_14821 (I254597,I254563,I2300);
nor I_14822 (I254614,I254521,I254597);
DFFARX1 I_14823 (I254614,I2595,I254478,I254464,);
nor I_14824 (I254645,I2300,I1484);
nand I_14825 (I254662,I254645,I2428);
DFFARX1 I_14826 (I254662,I2595,I254478,I254467,);
nor I_14827 (I254693,I254580,I2300);
nand I_14828 (I254710,I254693,I1684);
nor I_14829 (I254727,I254504,I254710);
DFFARX1 I_14830 (I254727,I2595,I254478,I254443,);
not I_14831 (I254758,I254710);
nand I_14832 (I254455,I254521,I254758);
DFFARX1 I_14833 (I254710,I2595,I254478,I254798,);
not I_14834 (I254806,I254798);
not I_14835 (I254823,I2300);
not I_14836 (I254840,I1412);
nor I_14837 (I254857,I254840,I1372);
nor I_14838 (I254470,I254806,I254857);
nor I_14839 (I254888,I254840,I2316);
and I_14840 (I254905,I254888,I1420);
or I_14841 (I254922,I254905,I2284);
DFFARX1 I_14842 (I254922,I2595,I254478,I254948,);
nor I_14843 (I254458,I254948,I254504);
not I_14844 (I254970,I254948);
and I_14845 (I254987,I254970,I254504);
nor I_14846 (I254452,I254529,I254987);
nand I_14847 (I255018,I254970,I254580);
nor I_14848 (I254446,I254840,I255018);
nand I_14849 (I254449,I254970,I254758);
nand I_14850 (I255063,I254580,I1412);
nor I_14851 (I254461,I254823,I255063);
not I_14852 (I255124,I2602);
DFFARX1 I_14853 (I218290,I2595,I255124,I255150,);
DFFARX1 I_14854 (I218284,I2595,I255124,I255167,);
not I_14855 (I255175,I255167);
not I_14856 (I255192,I218299);
nor I_14857 (I255209,I255192,I218284);
not I_14858 (I255226,I218293);
nor I_14859 (I255243,I255209,I218302);
nor I_14860 (I255260,I255167,I255243);
DFFARX1 I_14861 (I255260,I2595,I255124,I255110,);
nor I_14862 (I255291,I218302,I218284);
nand I_14863 (I255308,I255291,I218299);
DFFARX1 I_14864 (I255308,I2595,I255124,I255113,);
nor I_14865 (I255339,I255226,I218302);
nand I_14866 (I255356,I255339,I218287);
nor I_14867 (I255373,I255150,I255356);
DFFARX1 I_14868 (I255373,I2595,I255124,I255089,);
not I_14869 (I255404,I255356);
nand I_14870 (I255101,I255167,I255404);
DFFARX1 I_14871 (I255356,I2595,I255124,I255444,);
not I_14872 (I255452,I255444);
not I_14873 (I255469,I218302);
not I_14874 (I255486,I218296);
nor I_14875 (I255503,I255486,I218293);
nor I_14876 (I255116,I255452,I255503);
nor I_14877 (I255534,I255486,I218305);
and I_14878 (I255551,I255534,I218308);
or I_14879 (I255568,I255551,I218287);
DFFARX1 I_14880 (I255568,I2595,I255124,I255594,);
nor I_14881 (I255104,I255594,I255150);
not I_14882 (I255616,I255594);
and I_14883 (I255633,I255616,I255150);
nor I_14884 (I255098,I255175,I255633);
nand I_14885 (I255664,I255616,I255226);
nor I_14886 (I255092,I255486,I255664);
nand I_14887 (I255095,I255616,I255404);
nand I_14888 (I255709,I255226,I218296);
nor I_14889 (I255107,I255469,I255709);
not I_14890 (I255770,I2602);
DFFARX1 I_14891 (I162799,I2595,I255770,I255796,);
DFFARX1 I_14892 (I162811,I2595,I255770,I255813,);
not I_14893 (I255821,I255813);
not I_14894 (I255838,I162820);
nor I_14895 (I255855,I255838,I162796);
not I_14896 (I255872,I162814);
nor I_14897 (I255889,I255855,I162808);
nor I_14898 (I255906,I255813,I255889);
DFFARX1 I_14899 (I255906,I2595,I255770,I255756,);
nor I_14900 (I255937,I162808,I162796);
nand I_14901 (I255954,I255937,I162820);
DFFARX1 I_14902 (I255954,I2595,I255770,I255759,);
nor I_14903 (I255985,I255872,I162808);
nand I_14904 (I256002,I255985,I162802);
nor I_14905 (I256019,I255796,I256002);
DFFARX1 I_14906 (I256019,I2595,I255770,I255735,);
not I_14907 (I256050,I256002);
nand I_14908 (I255747,I255813,I256050);
DFFARX1 I_14909 (I256002,I2595,I255770,I256090,);
not I_14910 (I256098,I256090);
not I_14911 (I256115,I162808);
not I_14912 (I256132,I162817);
nor I_14913 (I256149,I256132,I162814);
nor I_14914 (I255762,I256098,I256149);
nor I_14915 (I256180,I256132,I162799);
and I_14916 (I256197,I256180,I162796);
or I_14917 (I256214,I256197,I162805);
DFFARX1 I_14918 (I256214,I2595,I255770,I256240,);
nor I_14919 (I255750,I256240,I255796);
not I_14920 (I256262,I256240);
and I_14921 (I256279,I256262,I255796);
nor I_14922 (I255744,I255821,I256279);
nand I_14923 (I256310,I256262,I255872);
nor I_14924 (I255738,I256132,I256310);
nand I_14925 (I255741,I256262,I256050);
nand I_14926 (I256355,I255872,I162817);
nor I_14927 (I255753,I256115,I256355);
not I_14928 (I256416,I2602);
DFFARX1 I_14929 (I2380,I2595,I256416,I256442,);
DFFARX1 I_14930 (I1796,I2595,I256416,I256459,);
not I_14931 (I256467,I256459);
not I_14932 (I256484,I1996);
nor I_14933 (I256501,I256484,I1900);
not I_14934 (I256518,I2468);
nor I_14935 (I256535,I256501,I2324);
nor I_14936 (I256552,I256459,I256535);
DFFARX1 I_14937 (I256552,I2595,I256416,I256402,);
nor I_14938 (I256583,I2324,I1900);
nand I_14939 (I256600,I256583,I1996);
DFFARX1 I_14940 (I256600,I2595,I256416,I256405,);
nor I_14941 (I256631,I256518,I2324);
nand I_14942 (I256648,I256631,I2036);
nor I_14943 (I256665,I256442,I256648);
DFFARX1 I_14944 (I256665,I2595,I256416,I256381,);
not I_14945 (I256696,I256648);
nand I_14946 (I256393,I256459,I256696);
DFFARX1 I_14947 (I256648,I2595,I256416,I256736,);
not I_14948 (I256744,I256736);
not I_14949 (I256761,I2324);
not I_14950 (I256778,I2348);
nor I_14951 (I256795,I256778,I2468);
nor I_14952 (I256408,I256744,I256795);
nor I_14953 (I256826,I256778,I2276);
and I_14954 (I256843,I256826,I2332);
or I_14955 (I256860,I256843,I2460);
DFFARX1 I_14956 (I256860,I2595,I256416,I256886,);
nor I_14957 (I256396,I256886,I256442);
not I_14958 (I256908,I256886);
and I_14959 (I256925,I256908,I256442);
nor I_14960 (I256390,I256467,I256925);
nand I_14961 (I256956,I256908,I256518);
nor I_14962 (I256384,I256778,I256956);
nand I_14963 (I256387,I256908,I256696);
nand I_14964 (I257001,I256518,I2348);
nor I_14965 (I256399,I256761,I257001);
not I_14966 (I257062,I2602);
DFFARX1 I_14967 (I123583,I2595,I257062,I257088,);
DFFARX1 I_14968 (I123580,I2595,I257062,I257105,);
not I_14969 (I257113,I257105);
not I_14970 (I257130,I123595);
nor I_14971 (I257147,I257130,I123598);
not I_14972 (I257164,I123586);
nor I_14973 (I257181,I257147,I123592);
nor I_14974 (I257198,I257105,I257181);
DFFARX1 I_14975 (I257198,I2595,I257062,I257048,);
nor I_14976 (I257229,I123592,I123598);
nand I_14977 (I257246,I257229,I123595);
DFFARX1 I_14978 (I257246,I2595,I257062,I257051,);
nor I_14979 (I257277,I257164,I123592);
nand I_14980 (I257294,I257277,I123604);
nor I_14981 (I257311,I257088,I257294);
DFFARX1 I_14982 (I257311,I2595,I257062,I257027,);
not I_14983 (I257342,I257294);
nand I_14984 (I257039,I257105,I257342);
DFFARX1 I_14985 (I257294,I2595,I257062,I257382,);
not I_14986 (I257390,I257382);
not I_14987 (I257407,I123592);
not I_14988 (I257424,I123577);
nor I_14989 (I257441,I257424,I123586);
nor I_14990 (I257054,I257390,I257441);
nor I_14991 (I257472,I257424,I123589);
and I_14992 (I257489,I257472,I123577);
or I_14993 (I257506,I257489,I123601);
DFFARX1 I_14994 (I257506,I2595,I257062,I257532,);
nor I_14995 (I257042,I257532,I257088);
not I_14996 (I257554,I257532);
and I_14997 (I257571,I257554,I257088);
nor I_14998 (I257036,I257113,I257571);
nand I_14999 (I257602,I257554,I257164);
nor I_15000 (I257030,I257424,I257602);
nand I_15001 (I257033,I257554,I257342);
nand I_15002 (I257647,I257164,I123577);
nor I_15003 (I257045,I257407,I257647);
not I_15004 (I257708,I2602);
DFFARX1 I_15005 (I130111,I2595,I257708,I257734,);
DFFARX1 I_15006 (I130108,I2595,I257708,I257751,);
not I_15007 (I257759,I257751);
not I_15008 (I257776,I130123);
nor I_15009 (I257793,I257776,I130126);
not I_15010 (I257810,I130114);
nor I_15011 (I257827,I257793,I130120);
nor I_15012 (I257844,I257751,I257827);
DFFARX1 I_15013 (I257844,I2595,I257708,I257694,);
nor I_15014 (I257875,I130120,I130126);
nand I_15015 (I257892,I257875,I130123);
DFFARX1 I_15016 (I257892,I2595,I257708,I257697,);
nor I_15017 (I257923,I257810,I130120);
nand I_15018 (I257940,I257923,I130132);
nor I_15019 (I257957,I257734,I257940);
DFFARX1 I_15020 (I257957,I2595,I257708,I257673,);
not I_15021 (I257988,I257940);
nand I_15022 (I257685,I257751,I257988);
DFFARX1 I_15023 (I257940,I2595,I257708,I258028,);
not I_15024 (I258036,I258028);
not I_15025 (I258053,I130120);
not I_15026 (I258070,I130105);
nor I_15027 (I258087,I258070,I130114);
nor I_15028 (I257700,I258036,I258087);
nor I_15029 (I258118,I258070,I130117);
and I_15030 (I258135,I258118,I130105);
or I_15031 (I258152,I258135,I130129);
DFFARX1 I_15032 (I258152,I2595,I257708,I258178,);
nor I_15033 (I257688,I258178,I257734);
not I_15034 (I258200,I258178);
and I_15035 (I258217,I258200,I257734);
nor I_15036 (I257682,I257759,I258217);
nand I_15037 (I258248,I258200,I257810);
nor I_15038 (I257676,I258070,I258248);
nand I_15039 (I257679,I258200,I257988);
nand I_15040 (I258293,I257810,I130105);
nor I_15041 (I257691,I258053,I258293);
not I_15042 (I258354,I2602);
DFFARX1 I_15043 (I238809,I2595,I258354,I258380,);
DFFARX1 I_15044 (I238806,I2595,I258354,I258397,);
not I_15045 (I258405,I258397);
not I_15046 (I258422,I238806);
nor I_15047 (I258439,I258422,I238809);
not I_15048 (I258456,I238821);
nor I_15049 (I258473,I258439,I238815);
nor I_15050 (I258490,I258397,I258473);
DFFARX1 I_15051 (I258490,I2595,I258354,I258340,);
nor I_15052 (I258521,I238815,I238809);
nand I_15053 (I258538,I258521,I238806);
DFFARX1 I_15054 (I258538,I2595,I258354,I258343,);
nor I_15055 (I258569,I258456,I238815);
nand I_15056 (I258586,I258569,I238803);
nor I_15057 (I258603,I258380,I258586);
DFFARX1 I_15058 (I258603,I2595,I258354,I258319,);
not I_15059 (I258634,I258586);
nand I_15060 (I258331,I258397,I258634);
DFFARX1 I_15061 (I258586,I2595,I258354,I258674,);
not I_15062 (I258682,I258674);
not I_15063 (I258699,I238815);
not I_15064 (I258716,I238812);
nor I_15065 (I258733,I258716,I238821);
nor I_15066 (I258346,I258682,I258733);
nor I_15067 (I258764,I258716,I238818);
and I_15068 (I258781,I258764,I238824);
or I_15069 (I258798,I258781,I238803);
DFFARX1 I_15070 (I258798,I2595,I258354,I258824,);
nor I_15071 (I258334,I258824,I258380);
not I_15072 (I258846,I258824);
and I_15073 (I258863,I258846,I258380);
nor I_15074 (I258328,I258405,I258863);
nand I_15075 (I258894,I258846,I258456);
nor I_15076 (I258322,I258716,I258894);
nand I_15077 (I258325,I258846,I258634);
nand I_15078 (I258939,I258456,I238812);
nor I_15079 (I258337,I258699,I258939);
not I_15080 (I259000,I2602);
DFFARX1 I_15081 (I110130,I2595,I259000,I259026,);
DFFARX1 I_15082 (I110136,I2595,I259000,I259043,);
not I_15083 (I259051,I259043);
not I_15084 (I259068,I110157);
nor I_15085 (I259085,I259068,I110145);
not I_15086 (I259102,I110154);
nor I_15087 (I259119,I259085,I110139);
nor I_15088 (I259136,I259043,I259119);
DFFARX1 I_15089 (I259136,I2595,I259000,I258986,);
nor I_15090 (I259167,I110139,I110145);
nand I_15091 (I259184,I259167,I110157);
DFFARX1 I_15092 (I259184,I2595,I259000,I258989,);
nor I_15093 (I259215,I259102,I110139);
nand I_15094 (I259232,I259215,I110130);
nor I_15095 (I259249,I259026,I259232);
DFFARX1 I_15096 (I259249,I2595,I259000,I258965,);
not I_15097 (I259280,I259232);
nand I_15098 (I258977,I259043,I259280);
DFFARX1 I_15099 (I259232,I2595,I259000,I259320,);
not I_15100 (I259328,I259320);
not I_15101 (I259345,I110139);
not I_15102 (I259362,I110142);
nor I_15103 (I259379,I259362,I110154);
nor I_15104 (I258992,I259328,I259379);
nor I_15105 (I259410,I259362,I110151);
and I_15106 (I259427,I259410,I110133);
or I_15107 (I259444,I259427,I110148);
DFFARX1 I_15108 (I259444,I2595,I259000,I259470,);
nor I_15109 (I258980,I259470,I259026);
not I_15110 (I259492,I259470);
and I_15111 (I259509,I259492,I259026);
nor I_15112 (I258974,I259051,I259509);
nand I_15113 (I259540,I259492,I259102);
nor I_15114 (I258968,I259362,I259540);
nand I_15115 (I258971,I259492,I259280);
nand I_15116 (I259585,I259102,I110142);
nor I_15117 (I258983,I259345,I259585);
not I_15118 (I259646,I2602);
DFFARX1 I_15119 (I390188,I2595,I259646,I259672,);
DFFARX1 I_15120 (I390212,I2595,I259646,I259689,);
not I_15121 (I259697,I259689);
not I_15122 (I259714,I390194);
nor I_15123 (I259731,I259714,I390203);
not I_15124 (I259748,I390188);
nor I_15125 (I259765,I259731,I390209);
nor I_15126 (I259782,I259689,I259765);
DFFARX1 I_15127 (I259782,I2595,I259646,I259632,);
nor I_15128 (I259813,I390209,I390203);
nand I_15129 (I259830,I259813,I390194);
DFFARX1 I_15130 (I259830,I2595,I259646,I259635,);
nor I_15131 (I259861,I259748,I390209);
nand I_15132 (I259878,I259861,I390206);
nor I_15133 (I259895,I259672,I259878);
DFFARX1 I_15134 (I259895,I2595,I259646,I259611,);
not I_15135 (I259926,I259878);
nand I_15136 (I259623,I259689,I259926);
DFFARX1 I_15137 (I259878,I2595,I259646,I259966,);
not I_15138 (I259974,I259966);
not I_15139 (I259991,I390209);
not I_15140 (I260008,I390200);
nor I_15141 (I260025,I260008,I390188);
nor I_15142 (I259638,I259974,I260025);
nor I_15143 (I260056,I260008,I390191);
and I_15144 (I260073,I260056,I390215);
or I_15145 (I260090,I260073,I390197);
DFFARX1 I_15146 (I260090,I2595,I259646,I260116,);
nor I_15147 (I259626,I260116,I259672);
not I_15148 (I260138,I260116);
and I_15149 (I260155,I260138,I259672);
nor I_15150 (I259620,I259697,I260155);
nand I_15151 (I260186,I260138,I259748);
nor I_15152 (I259614,I260008,I260186);
nand I_15153 (I259617,I260138,I259926);
nand I_15154 (I260231,I259748,I390200);
nor I_15155 (I259629,I259991,I260231);
not I_15156 (I260292,I2602);
DFFARX1 I_15157 (I95374,I2595,I260292,I260318,);
DFFARX1 I_15158 (I95380,I2595,I260292,I260335,);
not I_15159 (I260343,I260335);
not I_15160 (I260360,I95401);
nor I_15161 (I260377,I260360,I95389);
not I_15162 (I260394,I95398);
nor I_15163 (I260411,I260377,I95383);
nor I_15164 (I260428,I260335,I260411);
DFFARX1 I_15165 (I260428,I2595,I260292,I260278,);
nor I_15166 (I260459,I95383,I95389);
nand I_15167 (I260476,I260459,I95401);
DFFARX1 I_15168 (I260476,I2595,I260292,I260281,);
nor I_15169 (I260507,I260394,I95383);
nand I_15170 (I260524,I260507,I95374);
nor I_15171 (I260541,I260318,I260524);
DFFARX1 I_15172 (I260541,I2595,I260292,I260257,);
not I_15173 (I260572,I260524);
nand I_15174 (I260269,I260335,I260572);
DFFARX1 I_15175 (I260524,I2595,I260292,I260612,);
not I_15176 (I260620,I260612);
not I_15177 (I260637,I95383);
not I_15178 (I260654,I95386);
nor I_15179 (I260671,I260654,I95398);
nor I_15180 (I260284,I260620,I260671);
nor I_15181 (I260702,I260654,I95395);
and I_15182 (I260719,I260702,I95377);
or I_15183 (I260736,I260719,I95392);
DFFARX1 I_15184 (I260736,I2595,I260292,I260762,);
nor I_15185 (I260272,I260762,I260318);
not I_15186 (I260784,I260762);
and I_15187 (I260801,I260784,I260318);
nor I_15188 (I260266,I260343,I260801);
nand I_15189 (I260832,I260784,I260394);
nor I_15190 (I260260,I260654,I260832);
nand I_15191 (I260263,I260784,I260572);
nand I_15192 (I260877,I260394,I95386);
nor I_15193 (I260275,I260637,I260877);
not I_15194 (I260938,I2602);
DFFARX1 I_15195 (I228694,I2595,I260938,I260964,);
DFFARX1 I_15196 (I228688,I2595,I260938,I260981,);
not I_15197 (I260989,I260981);
not I_15198 (I261006,I228703);
nor I_15199 (I261023,I261006,I228688);
not I_15200 (I261040,I228697);
nor I_15201 (I261057,I261023,I228706);
nor I_15202 (I261074,I260981,I261057);
DFFARX1 I_15203 (I261074,I2595,I260938,I260924,);
nor I_15204 (I261105,I228706,I228688);
nand I_15205 (I261122,I261105,I228703);
DFFARX1 I_15206 (I261122,I2595,I260938,I260927,);
nor I_15207 (I261153,I261040,I228706);
nand I_15208 (I261170,I261153,I228691);
nor I_15209 (I261187,I260964,I261170);
DFFARX1 I_15210 (I261187,I2595,I260938,I260903,);
not I_15211 (I261218,I261170);
nand I_15212 (I260915,I260981,I261218);
DFFARX1 I_15213 (I261170,I2595,I260938,I261258,);
not I_15214 (I261266,I261258);
not I_15215 (I261283,I228706);
not I_15216 (I261300,I228700);
nor I_15217 (I261317,I261300,I228697);
nor I_15218 (I260930,I261266,I261317);
nor I_15219 (I261348,I261300,I228709);
and I_15220 (I261365,I261348,I228712);
or I_15221 (I261382,I261365,I228691);
DFFARX1 I_15222 (I261382,I2595,I260938,I261408,);
nor I_15223 (I260918,I261408,I260964);
not I_15224 (I261430,I261408);
and I_15225 (I261447,I261430,I260964);
nor I_15226 (I260912,I260989,I261447);
nand I_15227 (I261478,I261430,I261040);
nor I_15228 (I260906,I261300,I261478);
nand I_15229 (I260909,I261430,I261218);
nand I_15230 (I261523,I261040,I228700);
nor I_15231 (I260921,I261283,I261523);
not I_15232 (I261584,I2602);
DFFARX1 I_15233 (I2532,I2595,I261584,I261610,);
DFFARX1 I_15234 (I2140,I2595,I261584,I261627,);
not I_15235 (I261635,I261627);
not I_15236 (I261652,I2132);
nor I_15237 (I261669,I261652,I2548);
not I_15238 (I261686,I1556);
nor I_15239 (I261703,I261669,I2580);
nor I_15240 (I261720,I261627,I261703);
DFFARX1 I_15241 (I261720,I2595,I261584,I261570,);
nor I_15242 (I261751,I2580,I2548);
nand I_15243 (I261768,I261751,I2132);
DFFARX1 I_15244 (I261768,I2595,I261584,I261573,);
nor I_15245 (I261799,I261686,I2580);
nand I_15246 (I261816,I261799,I2012);
nor I_15247 (I261833,I261610,I261816);
DFFARX1 I_15248 (I261833,I2595,I261584,I261549,);
not I_15249 (I261864,I261816);
nand I_15250 (I261561,I261627,I261864);
DFFARX1 I_15251 (I261816,I2595,I261584,I261904,);
not I_15252 (I261912,I261904);
not I_15253 (I261929,I2580);
not I_15254 (I261946,I1804);
nor I_15255 (I261963,I261946,I1556);
nor I_15256 (I261576,I261912,I261963);
nor I_15257 (I261994,I261946,I1788);
and I_15258 (I262011,I261994,I1772);
or I_15259 (I262028,I262011,I2388);
DFFARX1 I_15260 (I262028,I2595,I261584,I262054,);
nor I_15261 (I261564,I262054,I261610);
not I_15262 (I262076,I262054);
and I_15263 (I262093,I262076,I261610);
nor I_15264 (I261558,I261635,I262093);
nand I_15265 (I262124,I262076,I261686);
nor I_15266 (I261552,I261946,I262124);
nand I_15267 (I261555,I262076,I261864);
nand I_15268 (I262169,I261686,I1804);
nor I_15269 (I261567,I261929,I262169);
not I_15270 (I262230,I2602);
DFFARX1 I_15271 (I294376,I2595,I262230,I262256,);
DFFARX1 I_15272 (I294379,I2595,I262230,I262273,);
not I_15273 (I262281,I262273);
not I_15274 (I262298,I294376);
nor I_15275 (I262315,I262298,I294388);
not I_15276 (I262332,I294397);
nor I_15277 (I262349,I262315,I294385);
nor I_15278 (I262366,I262273,I262349);
DFFARX1 I_15279 (I262366,I2595,I262230,I262216,);
nor I_15280 (I262397,I294385,I294388);
nand I_15281 (I262414,I262397,I294376);
DFFARX1 I_15282 (I262414,I2595,I262230,I262219,);
nor I_15283 (I262445,I262332,I294385);
nand I_15284 (I262462,I262445,I294391);
nor I_15285 (I262479,I262256,I262462);
DFFARX1 I_15286 (I262479,I2595,I262230,I262195,);
not I_15287 (I262510,I262462);
nand I_15288 (I262207,I262273,I262510);
DFFARX1 I_15289 (I262462,I2595,I262230,I262550,);
not I_15290 (I262558,I262550);
not I_15291 (I262575,I294385);
not I_15292 (I262592,I294382);
nor I_15293 (I262609,I262592,I294397);
nor I_15294 (I262222,I262558,I262609);
nor I_15295 (I262640,I262592,I294394);
and I_15296 (I262657,I262640,I294382);
or I_15297 (I262674,I262657,I294379);
DFFARX1 I_15298 (I262674,I2595,I262230,I262700,);
nor I_15299 (I262210,I262700,I262256);
not I_15300 (I262722,I262700);
and I_15301 (I262739,I262722,I262256);
nor I_15302 (I262204,I262281,I262739);
nand I_15303 (I262770,I262722,I262332);
nor I_15304 (I262198,I262592,I262770);
nand I_15305 (I262201,I262722,I262510);
nand I_15306 (I262815,I262332,I294382);
nor I_15307 (I262213,I262575,I262815);
not I_15308 (I262876,I2602);
DFFARX1 I_15309 (I332780,I2595,I262876,I262902,);
DFFARX1 I_15310 (I332762,I2595,I262876,I262919,);
not I_15311 (I262927,I262919);
not I_15312 (I262944,I332771);
nor I_15313 (I262961,I262944,I332783);
not I_15314 (I262978,I332765);
nor I_15315 (I262995,I262961,I332774);
nor I_15316 (I263012,I262919,I262995);
DFFARX1 I_15317 (I263012,I2595,I262876,I262862,);
nor I_15318 (I263043,I332774,I332783);
nand I_15319 (I263060,I263043,I332771);
DFFARX1 I_15320 (I263060,I2595,I262876,I262865,);
nor I_15321 (I263091,I262978,I332774);
nand I_15322 (I263108,I263091,I332786);
nor I_15323 (I263125,I262902,I263108);
DFFARX1 I_15324 (I263125,I2595,I262876,I262841,);
not I_15325 (I263156,I263108);
nand I_15326 (I262853,I262919,I263156);
DFFARX1 I_15327 (I263108,I2595,I262876,I263196,);
not I_15328 (I263204,I263196);
not I_15329 (I263221,I332774);
not I_15330 (I263238,I332762);
nor I_15331 (I263255,I263238,I332765);
nor I_15332 (I262868,I263204,I263255);
nor I_15333 (I263286,I263238,I332768);
and I_15334 (I263303,I263286,I332777);
or I_15335 (I263320,I263303,I332765);
DFFARX1 I_15336 (I263320,I2595,I262876,I263346,);
nor I_15337 (I262856,I263346,I262902);
not I_15338 (I263368,I263346);
and I_15339 (I263385,I263368,I262902);
nor I_15340 (I262850,I262927,I263385);
nand I_15341 (I263416,I263368,I262978);
nor I_15342 (I262844,I263238,I263416);
nand I_15343 (I262847,I263368,I263156);
nand I_15344 (I263461,I262978,I332762);
nor I_15345 (I262859,I263221,I263461);
not I_15346 (I263522,I2602);
DFFARX1 I_15347 (I23974,I2595,I263522,I263548,);
DFFARX1 I_15348 (I23980,I2595,I263522,I263565,);
not I_15349 (I263573,I263565);
not I_15350 (I263590,I23998);
nor I_15351 (I263607,I263590,I23977);
not I_15352 (I263624,I23983);
nor I_15353 (I263641,I263607,I23989);
nor I_15354 (I263658,I263565,I263641);
DFFARX1 I_15355 (I263658,I2595,I263522,I263508,);
nor I_15356 (I263689,I23989,I23977);
nand I_15357 (I263706,I263689,I23998);
DFFARX1 I_15358 (I263706,I2595,I263522,I263511,);
nor I_15359 (I263737,I263624,I23989);
nand I_15360 (I263754,I263737,I23995);
nor I_15361 (I263771,I263548,I263754);
DFFARX1 I_15362 (I263771,I2595,I263522,I263487,);
not I_15363 (I263802,I263754);
nand I_15364 (I263499,I263565,I263802);
DFFARX1 I_15365 (I263754,I2595,I263522,I263842,);
not I_15366 (I263850,I263842);
not I_15367 (I263867,I23989);
not I_15368 (I263884,I23977);
nor I_15369 (I263901,I263884,I23983);
nor I_15370 (I263514,I263850,I263901);
nor I_15371 (I263932,I263884,I23986);
and I_15372 (I263949,I263932,I23974);
or I_15373 (I263966,I263949,I23992);
DFFARX1 I_15374 (I263966,I2595,I263522,I263992,);
nor I_15375 (I263502,I263992,I263548);
not I_15376 (I264014,I263992);
and I_15377 (I264031,I264014,I263548);
nor I_15378 (I263496,I263573,I264031);
nand I_15379 (I264062,I264014,I263624);
nor I_15380 (I263490,I263884,I264062);
nand I_15381 (I263493,I264014,I263802);
nand I_15382 (I264107,I263624,I23977);
nor I_15383 (I263505,I263867,I264107);
not I_15384 (I264168,I2602);
DFFARX1 I_15385 (I167423,I2595,I264168,I264194,);
DFFARX1 I_15386 (I167435,I2595,I264168,I264211,);
not I_15387 (I264219,I264211);
not I_15388 (I264236,I167444);
nor I_15389 (I264253,I264236,I167420);
not I_15390 (I264270,I167438);
nor I_15391 (I264287,I264253,I167432);
nor I_15392 (I264304,I264211,I264287);
DFFARX1 I_15393 (I264304,I2595,I264168,I264154,);
nor I_15394 (I264335,I167432,I167420);
nand I_15395 (I264352,I264335,I167444);
DFFARX1 I_15396 (I264352,I2595,I264168,I264157,);
nor I_15397 (I264383,I264270,I167432);
nand I_15398 (I264400,I264383,I167426);
nor I_15399 (I264417,I264194,I264400);
DFFARX1 I_15400 (I264417,I2595,I264168,I264133,);
not I_15401 (I264448,I264400);
nand I_15402 (I264145,I264211,I264448);
DFFARX1 I_15403 (I264400,I2595,I264168,I264488,);
not I_15404 (I264496,I264488);
not I_15405 (I264513,I167432);
not I_15406 (I264530,I167441);
nor I_15407 (I264547,I264530,I167438);
nor I_15408 (I264160,I264496,I264547);
nor I_15409 (I264578,I264530,I167423);
and I_15410 (I264595,I264578,I167420);
or I_15411 (I264612,I264595,I167429);
DFFARX1 I_15412 (I264612,I2595,I264168,I264638,);
nor I_15413 (I264148,I264638,I264194);
not I_15414 (I264660,I264638);
and I_15415 (I264677,I264660,I264194);
nor I_15416 (I264142,I264219,I264677);
nand I_15417 (I264708,I264660,I264270);
nor I_15418 (I264136,I264530,I264708);
nand I_15419 (I264139,I264660,I264448);
nand I_15420 (I264753,I264270,I167441);
nor I_15421 (I264151,I264513,I264753);
not I_15422 (I264814,I2602);
DFFARX1 I_15423 (I80029,I2595,I264814,I264840,);
DFFARX1 I_15424 (I80041,I2595,I264814,I264857,);
not I_15425 (I264865,I264857);
not I_15426 (I264882,I80047);
nor I_15427 (I264899,I264882,I80032);
not I_15428 (I264916,I80023);
nor I_15429 (I264933,I264899,I80044);
nor I_15430 (I264950,I264857,I264933);
DFFARX1 I_15431 (I264950,I2595,I264814,I264800,);
nor I_15432 (I264981,I80044,I80032);
nand I_15433 (I264998,I264981,I80047);
DFFARX1 I_15434 (I264998,I2595,I264814,I264803,);
nor I_15435 (I265029,I264916,I80044);
nand I_15436 (I265046,I265029,I80026);
nor I_15437 (I265063,I264840,I265046);
DFFARX1 I_15438 (I265063,I2595,I264814,I264779,);
not I_15439 (I265094,I265046);
nand I_15440 (I264791,I264857,I265094);
DFFARX1 I_15441 (I265046,I2595,I264814,I265134,);
not I_15442 (I265142,I265134);
not I_15443 (I265159,I80044);
not I_15444 (I265176,I80035);
nor I_15445 (I265193,I265176,I80023);
nor I_15446 (I264806,I265142,I265193);
nor I_15447 (I265224,I265176,I80038);
and I_15448 (I265241,I265224,I80026);
or I_15449 (I265258,I265241,I80023);
DFFARX1 I_15450 (I265258,I2595,I264814,I265284,);
nor I_15451 (I264794,I265284,I264840);
not I_15452 (I265306,I265284);
and I_15453 (I265323,I265306,I264840);
nor I_15454 (I264788,I264865,I265323);
nand I_15455 (I265354,I265306,I264916);
nor I_15456 (I264782,I265176,I265354);
nand I_15457 (I264785,I265306,I265094);
nand I_15458 (I265399,I264916,I80035);
nor I_15459 (I264797,I265159,I265399);
not I_15460 (I265460,I2602);
DFFARX1 I_15461 (I59204,I2595,I265460,I265486,);
DFFARX1 I_15462 (I59216,I2595,I265460,I265503,);
not I_15463 (I265511,I265503);
not I_15464 (I265528,I59222);
nor I_15465 (I265545,I265528,I59207);
not I_15466 (I265562,I59198);
nor I_15467 (I265579,I265545,I59219);
nor I_15468 (I265596,I265503,I265579);
DFFARX1 I_15469 (I265596,I2595,I265460,I265446,);
nor I_15470 (I265627,I59219,I59207);
nand I_15471 (I265644,I265627,I59222);
DFFARX1 I_15472 (I265644,I2595,I265460,I265449,);
nor I_15473 (I265675,I265562,I59219);
nand I_15474 (I265692,I265675,I59201);
nor I_15475 (I265709,I265486,I265692);
DFFARX1 I_15476 (I265709,I2595,I265460,I265425,);
not I_15477 (I265740,I265692);
nand I_15478 (I265437,I265503,I265740);
DFFARX1 I_15479 (I265692,I2595,I265460,I265780,);
not I_15480 (I265788,I265780);
not I_15481 (I265805,I59219);
not I_15482 (I265822,I59210);
nor I_15483 (I265839,I265822,I59198);
nor I_15484 (I265452,I265788,I265839);
nor I_15485 (I265870,I265822,I59213);
and I_15486 (I265887,I265870,I59201);
or I_15487 (I265904,I265887,I59198);
DFFARX1 I_15488 (I265904,I2595,I265460,I265930,);
nor I_15489 (I265440,I265930,I265486);
not I_15490 (I265952,I265930);
and I_15491 (I265969,I265952,I265486);
nor I_15492 (I265434,I265511,I265969);
nand I_15493 (I266000,I265952,I265562);
nor I_15494 (I265428,I265822,I266000);
nand I_15495 (I265431,I265952,I265740);
nand I_15496 (I266045,I265562,I59210);
nor I_15497 (I265443,I265805,I266045);
not I_15498 (I266106,I2602);
DFFARX1 I_15499 (I118143,I2595,I266106,I266132,);
DFFARX1 I_15500 (I118140,I2595,I266106,I266149,);
not I_15501 (I266157,I266149);
not I_15502 (I266174,I118155);
nor I_15503 (I266191,I266174,I118158);
not I_15504 (I266208,I118146);
nor I_15505 (I266225,I266191,I118152);
nor I_15506 (I266242,I266149,I266225);
DFFARX1 I_15507 (I266242,I2595,I266106,I266092,);
nor I_15508 (I266273,I118152,I118158);
nand I_15509 (I266290,I266273,I118155);
DFFARX1 I_15510 (I266290,I2595,I266106,I266095,);
nor I_15511 (I266321,I266208,I118152);
nand I_15512 (I266338,I266321,I118164);
nor I_15513 (I266355,I266132,I266338);
DFFARX1 I_15514 (I266355,I2595,I266106,I266071,);
not I_15515 (I266386,I266338);
nand I_15516 (I266083,I266149,I266386);
DFFARX1 I_15517 (I266338,I2595,I266106,I266426,);
not I_15518 (I266434,I266426);
not I_15519 (I266451,I118152);
not I_15520 (I266468,I118137);
nor I_15521 (I266485,I266468,I118146);
nor I_15522 (I266098,I266434,I266485);
nor I_15523 (I266516,I266468,I118149);
and I_15524 (I266533,I266516,I118137);
or I_15525 (I266550,I266533,I118161);
DFFARX1 I_15526 (I266550,I2595,I266106,I266576,);
nor I_15527 (I266086,I266576,I266132);
not I_15528 (I266598,I266576);
and I_15529 (I266615,I266598,I266132);
nor I_15530 (I266080,I266157,I266615);
nand I_15531 (I266646,I266598,I266208);
nor I_15532 (I266074,I266468,I266646);
nand I_15533 (I266077,I266598,I266386);
nand I_15534 (I266691,I266208,I118137);
nor I_15535 (I266089,I266451,I266691);
not I_15536 (I266752,I2602);
DFFARX1 I_15537 (I304474,I2595,I266752,I266778,);
DFFARX1 I_15538 (I304477,I2595,I266752,I266795,);
not I_15539 (I266803,I266795);
not I_15540 (I266820,I304474);
nor I_15541 (I266837,I266820,I304486);
not I_15542 (I266854,I304495);
nor I_15543 (I266871,I266837,I304483);
nor I_15544 (I266888,I266795,I266871);
DFFARX1 I_15545 (I266888,I2595,I266752,I266738,);
nor I_15546 (I266919,I304483,I304486);
nand I_15547 (I266936,I266919,I304474);
DFFARX1 I_15548 (I266936,I2595,I266752,I266741,);
nor I_15549 (I266967,I266854,I304483);
nand I_15550 (I266984,I266967,I304489);
nor I_15551 (I267001,I266778,I266984);
DFFARX1 I_15552 (I267001,I2595,I266752,I266717,);
not I_15553 (I267032,I266984);
nand I_15554 (I266729,I266795,I267032);
DFFARX1 I_15555 (I266984,I2595,I266752,I267072,);
not I_15556 (I267080,I267072);
not I_15557 (I267097,I304483);
not I_15558 (I267114,I304480);
nor I_15559 (I267131,I267114,I304495);
nor I_15560 (I266744,I267080,I267131);
nor I_15561 (I267162,I267114,I304492);
and I_15562 (I267179,I267162,I304480);
or I_15563 (I267196,I267179,I304477);
DFFARX1 I_15564 (I267196,I2595,I266752,I267222,);
nor I_15565 (I266732,I267222,I266778);
not I_15566 (I267244,I267222);
and I_15567 (I267261,I267244,I266778);
nor I_15568 (I266726,I266803,I267261);
nand I_15569 (I267292,I267244,I266854);
nor I_15570 (I266720,I267114,I267292);
nand I_15571 (I266723,I267244,I267032);
nand I_15572 (I267337,I266854,I304480);
nor I_15573 (I266735,I267097,I267337);
not I_15574 (I267398,I2602);
DFFARX1 I_15575 (I65154,I2595,I267398,I267424,);
DFFARX1 I_15576 (I65166,I2595,I267398,I267441,);
not I_15577 (I267449,I267441);
not I_15578 (I267466,I65172);
nor I_15579 (I267483,I267466,I65157);
not I_15580 (I267500,I65148);
nor I_15581 (I267517,I267483,I65169);
nor I_15582 (I267534,I267441,I267517);
DFFARX1 I_15583 (I267534,I2595,I267398,I267384,);
nor I_15584 (I267565,I65169,I65157);
nand I_15585 (I267582,I267565,I65172);
DFFARX1 I_15586 (I267582,I2595,I267398,I267387,);
nor I_15587 (I267613,I267500,I65169);
nand I_15588 (I267630,I267613,I65151);
nor I_15589 (I267647,I267424,I267630);
DFFARX1 I_15590 (I267647,I2595,I267398,I267363,);
not I_15591 (I267678,I267630);
nand I_15592 (I267375,I267441,I267678);
DFFARX1 I_15593 (I267630,I2595,I267398,I267718,);
not I_15594 (I267726,I267718);
not I_15595 (I267743,I65169);
not I_15596 (I267760,I65160);
nor I_15597 (I267777,I267760,I65148);
nor I_15598 (I267390,I267726,I267777);
nor I_15599 (I267808,I267760,I65163);
and I_15600 (I267825,I267808,I65151);
or I_15601 (I267842,I267825,I65148);
DFFARX1 I_15602 (I267842,I2595,I267398,I267868,);
nor I_15603 (I267378,I267868,I267424);
not I_15604 (I267890,I267868);
and I_15605 (I267907,I267890,I267424);
nor I_15606 (I267372,I267449,I267907);
nand I_15607 (I267938,I267890,I267500);
nor I_15608 (I267366,I267760,I267938);
nand I_15609 (I267369,I267890,I267678);
nand I_15610 (I267983,I267500,I65160);
nor I_15611 (I267381,I267743,I267983);
not I_15612 (I268044,I2602);
DFFARX1 I_15613 (I157019,I2595,I268044,I268070,);
DFFARX1 I_15614 (I157031,I2595,I268044,I268087,);
not I_15615 (I268095,I268087);
not I_15616 (I268112,I157040);
nor I_15617 (I268129,I268112,I157016);
not I_15618 (I268146,I157034);
nor I_15619 (I268163,I268129,I157028);
nor I_15620 (I268180,I268087,I268163);
DFFARX1 I_15621 (I268180,I2595,I268044,I268030,);
nor I_15622 (I268211,I157028,I157016);
nand I_15623 (I268228,I268211,I157040);
DFFARX1 I_15624 (I268228,I2595,I268044,I268033,);
nor I_15625 (I268259,I268146,I157028);
nand I_15626 (I268276,I268259,I157022);
nor I_15627 (I268293,I268070,I268276);
DFFARX1 I_15628 (I268293,I2595,I268044,I268009,);
not I_15629 (I268324,I268276);
nand I_15630 (I268021,I268087,I268324);
DFFARX1 I_15631 (I268276,I2595,I268044,I268364,);
not I_15632 (I268372,I268364);
not I_15633 (I268389,I157028);
not I_15634 (I268406,I157037);
nor I_15635 (I268423,I268406,I157034);
nor I_15636 (I268036,I268372,I268423);
nor I_15637 (I268454,I268406,I157019);
and I_15638 (I268471,I268454,I157016);
or I_15639 (I268488,I268471,I157025);
DFFARX1 I_15640 (I268488,I2595,I268044,I268514,);
nor I_15641 (I268024,I268514,I268070);
not I_15642 (I268536,I268514);
and I_15643 (I268553,I268536,I268070);
nor I_15644 (I268018,I268095,I268553);
nand I_15645 (I268584,I268536,I268146);
nor I_15646 (I268012,I268406,I268584);
nand I_15647 (I268015,I268536,I268324);
nand I_15648 (I268629,I268146,I157037);
nor I_15649 (I268027,I268389,I268629);
not I_15650 (I268690,I2602);
DFFARX1 I_15651 (I45581,I2595,I268690,I268716,);
DFFARX1 I_15652 (I45587,I2595,I268690,I268733,);
not I_15653 (I268741,I268733);
not I_15654 (I268758,I45605);
nor I_15655 (I268775,I268758,I45584);
not I_15656 (I268792,I45590);
nor I_15657 (I268809,I268775,I45596);
nor I_15658 (I268826,I268733,I268809);
DFFARX1 I_15659 (I268826,I2595,I268690,I268676,);
nor I_15660 (I268857,I45596,I45584);
nand I_15661 (I268874,I268857,I45605);
DFFARX1 I_15662 (I268874,I2595,I268690,I268679,);
nor I_15663 (I268905,I268792,I45596);
nand I_15664 (I268922,I268905,I45602);
nor I_15665 (I268939,I268716,I268922);
DFFARX1 I_15666 (I268939,I2595,I268690,I268655,);
not I_15667 (I268970,I268922);
nand I_15668 (I268667,I268733,I268970);
DFFARX1 I_15669 (I268922,I2595,I268690,I269010,);
not I_15670 (I269018,I269010);
not I_15671 (I269035,I45596);
not I_15672 (I269052,I45584);
nor I_15673 (I269069,I269052,I45590);
nor I_15674 (I268682,I269018,I269069);
nor I_15675 (I269100,I269052,I45593);
and I_15676 (I269117,I269100,I45581);
or I_15677 (I269134,I269117,I45599);
DFFARX1 I_15678 (I269134,I2595,I268690,I269160,);
nor I_15679 (I268670,I269160,I268716);
not I_15680 (I269182,I269160);
and I_15681 (I269199,I269182,I268716);
nor I_15682 (I268664,I268741,I269199);
nand I_15683 (I269230,I269182,I268792);
nor I_15684 (I268658,I269052,I269230);
nand I_15685 (I268661,I269182,I268970);
nand I_15686 (I269275,I268792,I45584);
nor I_15687 (I268673,I269035,I269275);
not I_15688 (I269336,I2602);
DFFARX1 I_15689 (I130655,I2595,I269336,I269362,);
DFFARX1 I_15690 (I130652,I2595,I269336,I269379,);
not I_15691 (I269387,I269379);
not I_15692 (I269404,I130667);
nor I_15693 (I269421,I269404,I130670);
not I_15694 (I269438,I130658);
nor I_15695 (I269455,I269421,I130664);
nor I_15696 (I269472,I269379,I269455);
DFFARX1 I_15697 (I269472,I2595,I269336,I269322,);
nor I_15698 (I269503,I130664,I130670);
nand I_15699 (I269520,I269503,I130667);
DFFARX1 I_15700 (I269520,I2595,I269336,I269325,);
nor I_15701 (I269551,I269438,I130664);
nand I_15702 (I269568,I269551,I130676);
nor I_15703 (I269585,I269362,I269568);
DFFARX1 I_15704 (I269585,I2595,I269336,I269301,);
not I_15705 (I269616,I269568);
nand I_15706 (I269313,I269379,I269616);
DFFARX1 I_15707 (I269568,I2595,I269336,I269656,);
not I_15708 (I269664,I269656);
not I_15709 (I269681,I130664);
not I_15710 (I269698,I130649);
nor I_15711 (I269715,I269698,I130658);
nor I_15712 (I269328,I269664,I269715);
nor I_15713 (I269746,I269698,I130661);
and I_15714 (I269763,I269746,I130649);
or I_15715 (I269780,I269763,I130673);
DFFARX1 I_15716 (I269780,I2595,I269336,I269806,);
nor I_15717 (I269316,I269806,I269362);
not I_15718 (I269828,I269806);
and I_15719 (I269845,I269828,I269362);
nor I_15720 (I269310,I269387,I269845);
nand I_15721 (I269876,I269828,I269438);
nor I_15722 (I269304,I269698,I269876);
nand I_15723 (I269307,I269828,I269616);
nand I_15724 (I269921,I269438,I130649);
nor I_15725 (I269319,I269681,I269921);
not I_15726 (I269982,I2602);
DFFARX1 I_15727 (I148128,I2595,I269982,I270008,);
DFFARX1 I_15728 (I148140,I2595,I269982,I270025,);
not I_15729 (I270033,I270025);
not I_15730 (I270050,I148125);
nor I_15731 (I270067,I270050,I148143);
not I_15732 (I270084,I148149);
nor I_15733 (I270101,I270067,I148131);
nor I_15734 (I270118,I270025,I270101);
DFFARX1 I_15735 (I270118,I2595,I269982,I269968,);
nor I_15736 (I270149,I148131,I148143);
nand I_15737 (I270166,I270149,I148125);
DFFARX1 I_15738 (I270166,I2595,I269982,I269971,);
nor I_15739 (I270197,I270084,I148131);
nand I_15740 (I270214,I270197,I148134);
nor I_15741 (I270231,I270008,I270214);
DFFARX1 I_15742 (I270231,I2595,I269982,I269947,);
not I_15743 (I270262,I270214);
nand I_15744 (I269959,I270025,I270262);
DFFARX1 I_15745 (I270214,I2595,I269982,I270302,);
not I_15746 (I270310,I270302);
not I_15747 (I270327,I148131);
not I_15748 (I270344,I148137);
nor I_15749 (I270361,I270344,I148149);
nor I_15750 (I269974,I270310,I270361);
nor I_15751 (I270392,I270344,I148146);
and I_15752 (I270409,I270392,I148125);
or I_15753 (I270426,I270409,I148128);
DFFARX1 I_15754 (I270426,I2595,I269982,I270452,);
nor I_15755 (I269962,I270452,I270008);
not I_15756 (I270474,I270452);
and I_15757 (I270491,I270474,I270008);
nor I_15758 (I269956,I270033,I270491);
nand I_15759 (I270522,I270474,I270084);
nor I_15760 (I269950,I270344,I270522);
nand I_15761 (I269953,I270474,I270262);
nand I_15762 (I270567,I270084,I148137);
nor I_15763 (I269965,I270327,I270567);
not I_15764 (I270628,I2602);
DFFARX1 I_15765 (I311972,I2595,I270628,I270654,);
DFFARX1 I_15766 (I311954,I2595,I270628,I270671,);
not I_15767 (I270679,I270671);
not I_15768 (I270696,I311963);
nor I_15769 (I270713,I270696,I311975);
not I_15770 (I270730,I311957);
nor I_15771 (I270747,I270713,I311966);
nor I_15772 (I270764,I270671,I270747);
DFFARX1 I_15773 (I270764,I2595,I270628,I270614,);
nor I_15774 (I270795,I311966,I311975);
nand I_15775 (I270812,I270795,I311963);
DFFARX1 I_15776 (I270812,I2595,I270628,I270617,);
nor I_15777 (I270843,I270730,I311966);
nand I_15778 (I270860,I270843,I311978);
nor I_15779 (I270877,I270654,I270860);
DFFARX1 I_15780 (I270877,I2595,I270628,I270593,);
not I_15781 (I270908,I270860);
nand I_15782 (I270605,I270671,I270908);
DFFARX1 I_15783 (I270860,I2595,I270628,I270948,);
not I_15784 (I270956,I270948);
not I_15785 (I270973,I311966);
not I_15786 (I270990,I311954);
nor I_15787 (I271007,I270990,I311957);
nor I_15788 (I270620,I270956,I271007);
nor I_15789 (I271038,I270990,I311960);
and I_15790 (I271055,I271038,I311969);
or I_15791 (I271072,I271055,I311957);
DFFARX1 I_15792 (I271072,I2595,I270628,I271098,);
nor I_15793 (I270608,I271098,I270654);
not I_15794 (I271120,I271098);
and I_15795 (I271137,I271120,I270654);
nor I_15796 (I270602,I270679,I271137);
nand I_15797 (I271168,I271120,I270730);
nor I_15798 (I270596,I270990,I271168);
nand I_15799 (I270599,I271120,I270908);
nand I_15800 (I271213,I270730,I311954);
nor I_15801 (I270611,I270973,I271213);
not I_15802 (I271274,I2602);
DFFARX1 I_15803 (I392568,I2595,I271274,I271300,);
DFFARX1 I_15804 (I392592,I2595,I271274,I271317,);
not I_15805 (I271325,I271317);
not I_15806 (I271342,I392574);
nor I_15807 (I271359,I271342,I392583);
not I_15808 (I271376,I392568);
nor I_15809 (I271393,I271359,I392589);
nor I_15810 (I271410,I271317,I271393);
DFFARX1 I_15811 (I271410,I2595,I271274,I271260,);
nor I_15812 (I271441,I392589,I392583);
nand I_15813 (I271458,I271441,I392574);
DFFARX1 I_15814 (I271458,I2595,I271274,I271263,);
nor I_15815 (I271489,I271376,I392589);
nand I_15816 (I271506,I271489,I392586);
nor I_15817 (I271523,I271300,I271506);
DFFARX1 I_15818 (I271523,I2595,I271274,I271239,);
not I_15819 (I271554,I271506);
nand I_15820 (I271251,I271317,I271554);
DFFARX1 I_15821 (I271506,I2595,I271274,I271594,);
not I_15822 (I271602,I271594);
not I_15823 (I271619,I392589);
not I_15824 (I271636,I392580);
nor I_15825 (I271653,I271636,I392568);
nor I_15826 (I271266,I271602,I271653);
nor I_15827 (I271684,I271636,I392571);
and I_15828 (I271701,I271684,I392595);
or I_15829 (I271718,I271701,I392577);
DFFARX1 I_15830 (I271718,I2595,I271274,I271744,);
nor I_15831 (I271254,I271744,I271300);
not I_15832 (I271766,I271744);
and I_15833 (I271783,I271766,I271300);
nor I_15834 (I271248,I271325,I271783);
nand I_15835 (I271814,I271766,I271376);
nor I_15836 (I271242,I271636,I271814);
nand I_15837 (I271245,I271766,I271554);
nand I_15838 (I271859,I271376,I392580);
nor I_15839 (I271257,I271619,I271859);
not I_15840 (I271920,I2602);
DFFARX1 I_15841 (I26609,I2595,I271920,I271946,);
DFFARX1 I_15842 (I26615,I2595,I271920,I271963,);
not I_15843 (I271971,I271963);
not I_15844 (I271988,I26633);
nor I_15845 (I272005,I271988,I26612);
not I_15846 (I272022,I26618);
nor I_15847 (I272039,I272005,I26624);
nor I_15848 (I272056,I271963,I272039);
DFFARX1 I_15849 (I272056,I2595,I271920,I271906,);
nor I_15850 (I272087,I26624,I26612);
nand I_15851 (I272104,I272087,I26633);
DFFARX1 I_15852 (I272104,I2595,I271920,I271909,);
nor I_15853 (I272135,I272022,I26624);
nand I_15854 (I272152,I272135,I26630);
nor I_15855 (I272169,I271946,I272152);
DFFARX1 I_15856 (I272169,I2595,I271920,I271885,);
not I_15857 (I272200,I272152);
nand I_15858 (I271897,I271963,I272200);
DFFARX1 I_15859 (I272152,I2595,I271920,I272240,);
not I_15860 (I272248,I272240);
not I_15861 (I272265,I26624);
not I_15862 (I272282,I26612);
nor I_15863 (I272299,I272282,I26618);
nor I_15864 (I271912,I272248,I272299);
nor I_15865 (I272330,I272282,I26621);
and I_15866 (I272347,I272330,I26609);
or I_15867 (I272364,I272347,I26627);
DFFARX1 I_15868 (I272364,I2595,I271920,I272390,);
nor I_15869 (I271900,I272390,I271946);
not I_15870 (I272412,I272390);
and I_15871 (I272429,I272412,I271946);
nor I_15872 (I271894,I271971,I272429);
nand I_15873 (I272460,I272412,I272022);
nor I_15874 (I271888,I272282,I272460);
nand I_15875 (I271891,I272412,I272200);
nand I_15876 (I272505,I272022,I26612);
nor I_15877 (I271903,I272265,I272505);
not I_15878 (I272566,I2602);
DFFARX1 I_15879 (I109603,I2595,I272566,I272592,);
DFFARX1 I_15880 (I109609,I2595,I272566,I272609,);
not I_15881 (I272617,I272609);
not I_15882 (I272634,I109630);
nor I_15883 (I272651,I272634,I109618);
not I_15884 (I272668,I109627);
nor I_15885 (I272685,I272651,I109612);
nor I_15886 (I272702,I272609,I272685);
DFFARX1 I_15887 (I272702,I2595,I272566,I272552,);
nor I_15888 (I272733,I109612,I109618);
nand I_15889 (I272750,I272733,I109630);
DFFARX1 I_15890 (I272750,I2595,I272566,I272555,);
nor I_15891 (I272781,I272668,I109612);
nand I_15892 (I272798,I272781,I109603);
nor I_15893 (I272815,I272592,I272798);
DFFARX1 I_15894 (I272815,I2595,I272566,I272531,);
not I_15895 (I272846,I272798);
nand I_15896 (I272543,I272609,I272846);
DFFARX1 I_15897 (I272798,I2595,I272566,I272886,);
not I_15898 (I272894,I272886);
not I_15899 (I272911,I109612);
not I_15900 (I272928,I109615);
nor I_15901 (I272945,I272928,I109627);
nor I_15902 (I272558,I272894,I272945);
nor I_15903 (I272976,I272928,I109624);
and I_15904 (I272993,I272976,I109606);
or I_15905 (I273010,I272993,I109621);
DFFARX1 I_15906 (I273010,I2595,I272566,I273036,);
nor I_15907 (I272546,I273036,I272592);
not I_15908 (I273058,I273036);
and I_15909 (I273075,I273058,I272592);
nor I_15910 (I272540,I272617,I273075);
nand I_15911 (I273106,I273058,I272668);
nor I_15912 (I272534,I272928,I273106);
nand I_15913 (I272537,I273058,I272846);
nand I_15914 (I273151,I272668,I109615);
nor I_15915 (I272549,I272911,I273151);
not I_15916 (I273212,I2602);
DFFARX1 I_15917 (I387808,I2595,I273212,I273238,);
DFFARX1 I_15918 (I387832,I2595,I273212,I273255,);
not I_15919 (I273263,I273255);
not I_15920 (I273280,I387814);
nor I_15921 (I273297,I273280,I387823);
not I_15922 (I273314,I387808);
nor I_15923 (I273331,I273297,I387829);
nor I_15924 (I273348,I273255,I273331);
DFFARX1 I_15925 (I273348,I2595,I273212,I273198,);
nor I_15926 (I273379,I387829,I387823);
nand I_15927 (I273396,I273379,I387814);
DFFARX1 I_15928 (I273396,I2595,I273212,I273201,);
nor I_15929 (I273427,I273314,I387829);
nand I_15930 (I273444,I273427,I387826);
nor I_15931 (I273461,I273238,I273444);
DFFARX1 I_15932 (I273461,I2595,I273212,I273177,);
not I_15933 (I273492,I273444);
nand I_15934 (I273189,I273255,I273492);
DFFARX1 I_15935 (I273444,I2595,I273212,I273532,);
not I_15936 (I273540,I273532);
not I_15937 (I273557,I387829);
not I_15938 (I273574,I387820);
nor I_15939 (I273591,I273574,I387808);
nor I_15940 (I273204,I273540,I273591);
nor I_15941 (I273622,I273574,I387811);
and I_15942 (I273639,I273622,I387835);
or I_15943 (I273656,I273639,I387817);
DFFARX1 I_15944 (I273656,I2595,I273212,I273682,);
nor I_15945 (I273192,I273682,I273238);
not I_15946 (I273704,I273682);
and I_15947 (I273721,I273704,I273238);
nor I_15948 (I273186,I273263,I273721);
nand I_15949 (I273752,I273704,I273314);
nor I_15950 (I273180,I273574,I273752);
nand I_15951 (I273183,I273704,I273492);
nand I_15952 (I273797,I273314,I387820);
nor I_15953 (I273195,I273557,I273797);
not I_15954 (I273858,I2602);
DFFARX1 I_15955 (I363711,I2595,I273858,I273884,);
DFFARX1 I_15956 (I363705,I2595,I273858,I273901,);
not I_15957 (I273909,I273901);
not I_15958 (I273926,I363714);
nor I_15959 (I273943,I273926,I363726);
not I_15960 (I273960,I363708);
nor I_15961 (I273977,I273943,I363705);
nor I_15962 (I273994,I273901,I273977);
DFFARX1 I_15963 (I273994,I2595,I273858,I273844,);
nor I_15964 (I274025,I363705,I363726);
nand I_15965 (I274042,I274025,I363714);
DFFARX1 I_15966 (I274042,I2595,I273858,I273847,);
nor I_15967 (I274073,I273960,I363705);
nand I_15968 (I274090,I274073,I363702);
nor I_15969 (I274107,I273884,I274090);
DFFARX1 I_15970 (I274107,I2595,I273858,I273823,);
not I_15971 (I274138,I274090);
nand I_15972 (I273835,I273901,I274138);
DFFARX1 I_15973 (I274090,I2595,I273858,I274178,);
not I_15974 (I274186,I274178);
not I_15975 (I274203,I363705);
not I_15976 (I274220,I363723);
nor I_15977 (I274237,I274220,I363708);
nor I_15978 (I273850,I274186,I274237);
nor I_15979 (I274268,I274220,I363717);
and I_15980 (I274285,I274268,I363702);
or I_15981 (I274302,I274285,I363720);
DFFARX1 I_15982 (I274302,I2595,I273858,I274328,);
nor I_15983 (I273838,I274328,I273884);
not I_15984 (I274350,I274328);
and I_15985 (I274367,I274350,I273884);
nor I_15986 (I273832,I273909,I274367);
nand I_15987 (I274398,I274350,I273960);
nor I_15988 (I273826,I274220,I274398);
nand I_15989 (I273829,I274350,I274138);
nand I_15990 (I274443,I273960,I363723);
nor I_15991 (I273841,I274203,I274443);
not I_15992 (I274504,I2602);
DFFARX1 I_15993 (I169157,I2595,I274504,I274530,);
DFFARX1 I_15994 (I169169,I2595,I274504,I274547,);
not I_15995 (I274555,I274547);
not I_15996 (I274572,I169178);
nor I_15997 (I274589,I274572,I169154);
not I_15998 (I274606,I169172);
nor I_15999 (I274623,I274589,I169166);
nor I_16000 (I274640,I274547,I274623);
DFFARX1 I_16001 (I274640,I2595,I274504,I274490,);
nor I_16002 (I274671,I169166,I169154);
nand I_16003 (I274688,I274671,I169178);
DFFARX1 I_16004 (I274688,I2595,I274504,I274493,);
nor I_16005 (I274719,I274606,I169166);
nand I_16006 (I274736,I274719,I169160);
nor I_16007 (I274753,I274530,I274736);
DFFARX1 I_16008 (I274753,I2595,I274504,I274469,);
not I_16009 (I274784,I274736);
nand I_16010 (I274481,I274547,I274784);
DFFARX1 I_16011 (I274736,I2595,I274504,I274824,);
not I_16012 (I274832,I274824);
not I_16013 (I274849,I169166);
not I_16014 (I274866,I169175);
nor I_16015 (I274883,I274866,I169172);
nor I_16016 (I274496,I274832,I274883);
nor I_16017 (I274914,I274866,I169157);
and I_16018 (I274931,I274914,I169154);
or I_16019 (I274948,I274931,I169163);
DFFARX1 I_16020 (I274948,I2595,I274504,I274974,);
nor I_16021 (I274484,I274974,I274530);
not I_16022 (I274996,I274974);
and I_16023 (I275013,I274996,I274530);
nor I_16024 (I274478,I274555,I275013);
nand I_16025 (I275044,I274996,I274606);
nor I_16026 (I274472,I274866,I275044);
nand I_16027 (I274475,I274996,I274784);
nand I_16028 (I275089,I274606,I169175);
nor I_16029 (I274487,I274849,I275089);
not I_16030 (I275150,I2602);
DFFARX1 I_16031 (I13434,I2595,I275150,I275176,);
DFFARX1 I_16032 (I13440,I2595,I275150,I275193,);
not I_16033 (I275201,I275193);
not I_16034 (I275218,I13434);
nor I_16035 (I275235,I275218,I13446);
not I_16036 (I275252,I13458);
nor I_16037 (I275269,I275235,I13452);
nor I_16038 (I275286,I275193,I275269);
DFFARX1 I_16039 (I275286,I2595,I275150,I275136,);
nor I_16040 (I275317,I13452,I13446);
nand I_16041 (I275334,I275317,I13434);
DFFARX1 I_16042 (I275334,I2595,I275150,I275139,);
nor I_16043 (I275365,I275252,I13452);
nand I_16044 (I275382,I275365,I13437);
nor I_16045 (I275399,I275176,I275382);
DFFARX1 I_16046 (I275399,I2595,I275150,I275115,);
not I_16047 (I275430,I275382);
nand I_16048 (I275127,I275193,I275430);
DFFARX1 I_16049 (I275382,I2595,I275150,I275470,);
not I_16050 (I275478,I275470);
not I_16051 (I275495,I13452);
not I_16052 (I275512,I13437);
nor I_16053 (I275529,I275512,I13458);
nor I_16054 (I275142,I275478,I275529);
nor I_16055 (I275560,I275512,I13455);
and I_16056 (I275577,I275560,I13449);
or I_16057 (I275594,I275577,I13443);
DFFARX1 I_16058 (I275594,I2595,I275150,I275620,);
nor I_16059 (I275130,I275620,I275176);
not I_16060 (I275642,I275620);
and I_16061 (I275659,I275642,I275176);
nor I_16062 (I275124,I275201,I275659);
nand I_16063 (I275690,I275642,I275252);
nor I_16064 (I275118,I275512,I275690);
nand I_16065 (I275121,I275642,I275430);
nand I_16066 (I275735,I275252,I13437);
nor I_16067 (I275133,I275495,I275735);
not I_16068 (I275796,I2602);
DFFARX1 I_16069 (I336826,I2595,I275796,I275822,);
DFFARX1 I_16070 (I336808,I2595,I275796,I275839,);
not I_16071 (I275847,I275839);
not I_16072 (I275864,I336817);
nor I_16073 (I275881,I275864,I336829);
not I_16074 (I275898,I336811);
nor I_16075 (I275915,I275881,I336820);
nor I_16076 (I275932,I275839,I275915);
DFFARX1 I_16077 (I275932,I2595,I275796,I275782,);
nor I_16078 (I275963,I336820,I336829);
nand I_16079 (I275980,I275963,I336817);
DFFARX1 I_16080 (I275980,I2595,I275796,I275785,);
nor I_16081 (I276011,I275898,I336820);
nand I_16082 (I276028,I276011,I336832);
nor I_16083 (I276045,I275822,I276028);
DFFARX1 I_16084 (I276045,I2595,I275796,I275761,);
not I_16085 (I276076,I276028);
nand I_16086 (I275773,I275839,I276076);
DFFARX1 I_16087 (I276028,I2595,I275796,I276116,);
not I_16088 (I276124,I276116);
not I_16089 (I276141,I336820);
not I_16090 (I276158,I336808);
nor I_16091 (I276175,I276158,I336811);
nor I_16092 (I275788,I276124,I276175);
nor I_16093 (I276206,I276158,I336814);
and I_16094 (I276223,I276206,I336823);
or I_16095 (I276240,I276223,I336811);
DFFARX1 I_16096 (I276240,I2595,I275796,I276266,);
nor I_16097 (I275776,I276266,I275822);
not I_16098 (I276288,I276266);
and I_16099 (I276305,I276288,I275822);
nor I_16100 (I275770,I275847,I276305);
nand I_16101 (I276336,I276288,I275898);
nor I_16102 (I275764,I276158,I276336);
nand I_16103 (I275767,I276288,I276076);
nand I_16104 (I276381,I275898,I336808);
nor I_16105 (I275779,I276141,I276381);
not I_16106 (I276442,I2602);
DFFARX1 I_16107 (I84307,I2595,I276442,I276468,);
DFFARX1 I_16108 (I84313,I2595,I276442,I276485,);
not I_16109 (I276493,I276485);
not I_16110 (I276510,I84334);
nor I_16111 (I276527,I276510,I84322);
not I_16112 (I276544,I84331);
nor I_16113 (I276561,I276527,I84316);
nor I_16114 (I276578,I276485,I276561);
DFFARX1 I_16115 (I276578,I2595,I276442,I276428,);
nor I_16116 (I276609,I84316,I84322);
nand I_16117 (I276626,I276609,I84334);
DFFARX1 I_16118 (I276626,I2595,I276442,I276431,);
nor I_16119 (I276657,I276544,I84316);
nand I_16120 (I276674,I276657,I84307);
nor I_16121 (I276691,I276468,I276674);
DFFARX1 I_16122 (I276691,I2595,I276442,I276407,);
not I_16123 (I276722,I276674);
nand I_16124 (I276419,I276485,I276722);
DFFARX1 I_16125 (I276674,I2595,I276442,I276762,);
not I_16126 (I276770,I276762);
not I_16127 (I276787,I84316);
not I_16128 (I276804,I84319);
nor I_16129 (I276821,I276804,I84331);
nor I_16130 (I276434,I276770,I276821);
nor I_16131 (I276852,I276804,I84328);
and I_16132 (I276869,I276852,I84310);
or I_16133 (I276886,I276869,I84325);
DFFARX1 I_16134 (I276886,I2595,I276442,I276912,);
nor I_16135 (I276422,I276912,I276468);
not I_16136 (I276934,I276912);
and I_16137 (I276951,I276934,I276468);
nor I_16138 (I276416,I276493,I276951);
nand I_16139 (I276982,I276934,I276544);
nor I_16140 (I276410,I276804,I276982);
nand I_16141 (I276413,I276934,I276722);
nand I_16142 (I277027,I276544,I84319);
nor I_16143 (I276425,I276787,I277027);
not I_16144 (I277088,I2602);
DFFARX1 I_16145 (I112765,I2595,I277088,I277114,);
DFFARX1 I_16146 (I112771,I2595,I277088,I277131,);
not I_16147 (I277139,I277131);
not I_16148 (I277156,I112792);
nor I_16149 (I277173,I277156,I112780);
not I_16150 (I277190,I112789);
nor I_16151 (I277207,I277173,I112774);
nor I_16152 (I277224,I277131,I277207);
DFFARX1 I_16153 (I277224,I2595,I277088,I277074,);
nor I_16154 (I277255,I112774,I112780);
nand I_16155 (I277272,I277255,I112792);
DFFARX1 I_16156 (I277272,I2595,I277088,I277077,);
nor I_16157 (I277303,I277190,I112774);
nand I_16158 (I277320,I277303,I112765);
nor I_16159 (I277337,I277114,I277320);
DFFARX1 I_16160 (I277337,I2595,I277088,I277053,);
not I_16161 (I277368,I277320);
nand I_16162 (I277065,I277131,I277368);
DFFARX1 I_16163 (I277320,I2595,I277088,I277408,);
not I_16164 (I277416,I277408);
not I_16165 (I277433,I112774);
not I_16166 (I277450,I112777);
nor I_16167 (I277467,I277450,I112789);
nor I_16168 (I277080,I277416,I277467);
nor I_16169 (I277498,I277450,I112786);
and I_16170 (I277515,I277498,I112768);
or I_16171 (I277532,I277515,I112783);
DFFARX1 I_16172 (I277532,I2595,I277088,I277558,);
nor I_16173 (I277068,I277558,I277114);
not I_16174 (I277580,I277558);
and I_16175 (I277597,I277580,I277114);
nor I_16176 (I277062,I277139,I277597);
nand I_16177 (I277628,I277580,I277190);
nor I_16178 (I277056,I277450,I277628);
nand I_16179 (I277059,I277580,I277368);
nand I_16180 (I277673,I277190,I112777);
nor I_16181 (I277071,I277433,I277673);
not I_16182 (I277734,I2602);
DFFARX1 I_16183 (I191124,I2595,I277734,I277760,);
DFFARX1 I_16184 (I191118,I2595,I277734,I277777,);
not I_16185 (I277785,I277777);
not I_16186 (I277802,I191133);
nor I_16187 (I277819,I277802,I191118);
not I_16188 (I277836,I191127);
nor I_16189 (I277853,I277819,I191136);
nor I_16190 (I277870,I277777,I277853);
DFFARX1 I_16191 (I277870,I2595,I277734,I277720,);
nor I_16192 (I277901,I191136,I191118);
nand I_16193 (I277918,I277901,I191133);
DFFARX1 I_16194 (I277918,I2595,I277734,I277723,);
nor I_16195 (I277949,I277836,I191136);
nand I_16196 (I277966,I277949,I191121);
nor I_16197 (I277983,I277760,I277966);
DFFARX1 I_16198 (I277983,I2595,I277734,I277699,);
not I_16199 (I278014,I277966);
nand I_16200 (I277711,I277777,I278014);
DFFARX1 I_16201 (I277966,I2595,I277734,I278054,);
not I_16202 (I278062,I278054);
not I_16203 (I278079,I191136);
not I_16204 (I278096,I191130);
nor I_16205 (I278113,I278096,I191127);
nor I_16206 (I277726,I278062,I278113);
nor I_16207 (I278144,I278096,I191139);
and I_16208 (I278161,I278144,I191142);
or I_16209 (I278178,I278161,I191121);
DFFARX1 I_16210 (I278178,I2595,I277734,I278204,);
nor I_16211 (I277714,I278204,I277760);
not I_16212 (I278226,I278204);
and I_16213 (I278243,I278226,I277760);
nor I_16214 (I277708,I277785,I278243);
nand I_16215 (I278274,I278226,I277836);
nor I_16216 (I277702,I278096,I278274);
nand I_16217 (I277705,I278226,I278014);
nand I_16218 (I278319,I277836,I191130);
nor I_16219 (I277717,I278079,I278319);
not I_16220 (I278380,I2602);
DFFARX1 I_16221 (I290449,I2595,I278380,I278406,);
DFFARX1 I_16222 (I290452,I2595,I278380,I278423,);
not I_16223 (I278431,I278423);
not I_16224 (I278448,I290449);
nor I_16225 (I278465,I278448,I290461);
not I_16226 (I278482,I290470);
nor I_16227 (I278499,I278465,I290458);
nor I_16228 (I278516,I278423,I278499);
DFFARX1 I_16229 (I278516,I2595,I278380,I278366,);
nor I_16230 (I278547,I290458,I290461);
nand I_16231 (I278564,I278547,I290449);
DFFARX1 I_16232 (I278564,I2595,I278380,I278369,);
nor I_16233 (I278595,I278482,I290458);
nand I_16234 (I278612,I278595,I290464);
nor I_16235 (I278629,I278406,I278612);
DFFARX1 I_16236 (I278629,I2595,I278380,I278345,);
not I_16237 (I278660,I278612);
nand I_16238 (I278357,I278423,I278660);
DFFARX1 I_16239 (I278612,I2595,I278380,I278700,);
not I_16240 (I278708,I278700);
not I_16241 (I278725,I290458);
not I_16242 (I278742,I290455);
nor I_16243 (I278759,I278742,I290470);
nor I_16244 (I278372,I278708,I278759);
nor I_16245 (I278790,I278742,I290467);
and I_16246 (I278807,I278790,I290455);
or I_16247 (I278824,I278807,I290452);
DFFARX1 I_16248 (I278824,I2595,I278380,I278850,);
nor I_16249 (I278360,I278850,I278406);
not I_16250 (I278872,I278850);
and I_16251 (I278889,I278872,I278406);
nor I_16252 (I278354,I278431,I278889);
nand I_16253 (I278920,I278872,I278482);
nor I_16254 (I278348,I278742,I278920);
nand I_16255 (I278351,I278872,I278660);
nand I_16256 (I278965,I278482,I290455);
nor I_16257 (I278363,I278725,I278965);
not I_16258 (I279026,I2602);
DFFARX1 I_16259 (I106441,I2595,I279026,I279052,);
DFFARX1 I_16260 (I106447,I2595,I279026,I279069,);
not I_16261 (I279077,I279069);
not I_16262 (I279094,I106468);
nor I_16263 (I279111,I279094,I106456);
not I_16264 (I279128,I106465);
nor I_16265 (I279145,I279111,I106450);
nor I_16266 (I279162,I279069,I279145);
DFFARX1 I_16267 (I279162,I2595,I279026,I279012,);
nor I_16268 (I279193,I106450,I106456);
nand I_16269 (I279210,I279193,I106468);
DFFARX1 I_16270 (I279210,I2595,I279026,I279015,);
nor I_16271 (I279241,I279128,I106450);
nand I_16272 (I279258,I279241,I106441);
nor I_16273 (I279275,I279052,I279258);
DFFARX1 I_16274 (I279275,I2595,I279026,I278991,);
not I_16275 (I279306,I279258);
nand I_16276 (I279003,I279069,I279306);
DFFARX1 I_16277 (I279258,I2595,I279026,I279346,);
not I_16278 (I279354,I279346);
not I_16279 (I279371,I106450);
not I_16280 (I279388,I106453);
nor I_16281 (I279405,I279388,I106465);
nor I_16282 (I279018,I279354,I279405);
nor I_16283 (I279436,I279388,I106462);
and I_16284 (I279453,I279436,I106444);
or I_16285 (I279470,I279453,I106459);
DFFARX1 I_16286 (I279470,I2595,I279026,I279496,);
nor I_16287 (I279006,I279496,I279052);
not I_16288 (I279518,I279496);
and I_16289 (I279535,I279518,I279052);
nor I_16290 (I279000,I279077,I279535);
nand I_16291 (I279566,I279518,I279128);
nor I_16292 (I278994,I279388,I279566);
nand I_16293 (I278997,I279518,I279306);
nand I_16294 (I279611,I279128,I106453);
nor I_16295 (I279009,I279371,I279611);
not I_16296 (I279672,I2602);
DFFARX1 I_16297 (I345904,I2595,I279672,I279698,);
DFFARX1 I_16298 (I345910,I2595,I279672,I279715,);
not I_16299 (I279723,I279715);
not I_16300 (I279740,I345907);
nor I_16301 (I279757,I279740,I345886);
not I_16302 (I279774,I345889);
nor I_16303 (I279791,I279757,I345895);
nor I_16304 (I279808,I279715,I279791);
DFFARX1 I_16305 (I279808,I2595,I279672,I279658,);
nor I_16306 (I279839,I345895,I345886);
nand I_16307 (I279856,I279839,I345907);
DFFARX1 I_16308 (I279856,I2595,I279672,I279661,);
nor I_16309 (I279887,I279774,I345895);
nand I_16310 (I279904,I279887,I345889);
nor I_16311 (I279921,I279698,I279904);
DFFARX1 I_16312 (I279921,I2595,I279672,I279637,);
not I_16313 (I279952,I279904);
nand I_16314 (I279649,I279715,I279952);
DFFARX1 I_16315 (I279904,I2595,I279672,I279992,);
not I_16316 (I280000,I279992);
not I_16317 (I280017,I345895);
not I_16318 (I280034,I345898);
nor I_16319 (I280051,I280034,I345889);
nor I_16320 (I279664,I280000,I280051);
nor I_16321 (I280082,I280034,I345886);
and I_16322 (I280099,I280082,I345892);
or I_16323 (I280116,I280099,I345901);
DFFARX1 I_16324 (I280116,I2595,I279672,I280142,);
nor I_16325 (I279652,I280142,I279698);
not I_16326 (I280164,I280142);
and I_16327 (I280181,I280164,I279698);
nor I_16328 (I279646,I279723,I280181);
nand I_16329 (I280212,I280164,I279774);
nor I_16330 (I279640,I280034,I280212);
nand I_16331 (I279643,I280164,I279952);
nand I_16332 (I280257,I279774,I345898);
nor I_16333 (I279655,I280017,I280257);
not I_16334 (I280318,I2602);
DFFARX1 I_16335 (I1508,I2595,I280318,I280344,);
DFFARX1 I_16336 (I1892,I2595,I280318,I280361,);
not I_16337 (I280369,I280361);
not I_16338 (I280386,I2412);
nor I_16339 (I280403,I280386,I1596);
not I_16340 (I280420,I1548);
nor I_16341 (I280437,I280403,I1732);
nor I_16342 (I280454,I280361,I280437);
DFFARX1 I_16343 (I280454,I2595,I280318,I280304,);
nor I_16344 (I280485,I1732,I1596);
nand I_16345 (I280502,I280485,I2412);
DFFARX1 I_16346 (I280502,I2595,I280318,I280307,);
nor I_16347 (I280533,I280420,I1732);
nand I_16348 (I280550,I280533,I1692);
nor I_16349 (I280567,I280344,I280550);
DFFARX1 I_16350 (I280567,I2595,I280318,I280283,);
not I_16351 (I280598,I280550);
nand I_16352 (I280295,I280361,I280598);
DFFARX1 I_16353 (I280550,I2595,I280318,I280638,);
not I_16354 (I280646,I280638);
not I_16355 (I280663,I1732);
not I_16356 (I280680,I1924);
nor I_16357 (I280697,I280680,I1548);
nor I_16358 (I280310,I280646,I280697);
nor I_16359 (I280728,I280680,I2044);
and I_16360 (I280745,I280728,I1852);
or I_16361 (I280762,I280745,I1580);
DFFARX1 I_16362 (I280762,I2595,I280318,I280788,);
nor I_16363 (I280298,I280788,I280344);
not I_16364 (I280810,I280788);
and I_16365 (I280827,I280810,I280344);
nor I_16366 (I280292,I280369,I280827);
nand I_16367 (I280858,I280810,I280420);
nor I_16368 (I280286,I280680,I280858);
nand I_16369 (I280289,I280810,I280598);
nand I_16370 (I280903,I280420,I1924);
nor I_16371 (I280301,I280663,I280903);
not I_16372 (I280964,I2602);
DFFARX1 I_16373 (I75864,I2595,I280964,I280990,);
DFFARX1 I_16374 (I75876,I2595,I280964,I281007,);
not I_16375 (I281015,I281007);
not I_16376 (I281032,I75882);
nor I_16377 (I281049,I281032,I75867);
not I_16378 (I281066,I75858);
nor I_16379 (I281083,I281049,I75879);
nor I_16380 (I281100,I281007,I281083);
DFFARX1 I_16381 (I281100,I2595,I280964,I280950,);
nor I_16382 (I281131,I75879,I75867);
nand I_16383 (I281148,I281131,I75882);
DFFARX1 I_16384 (I281148,I2595,I280964,I280953,);
nor I_16385 (I281179,I281066,I75879);
nand I_16386 (I281196,I281179,I75861);
nor I_16387 (I281213,I280990,I281196);
DFFARX1 I_16388 (I281213,I2595,I280964,I280929,);
not I_16389 (I281244,I281196);
nand I_16390 (I280941,I281007,I281244);
DFFARX1 I_16391 (I281196,I2595,I280964,I281284,);
not I_16392 (I281292,I281284);
not I_16393 (I281309,I75879);
not I_16394 (I281326,I75870);
nor I_16395 (I281343,I281326,I75858);
nor I_16396 (I280956,I281292,I281343);
nor I_16397 (I281374,I281326,I75873);
and I_16398 (I281391,I281374,I75861);
or I_16399 (I281408,I281391,I75858);
DFFARX1 I_16400 (I281408,I2595,I280964,I281434,);
nor I_16401 (I280944,I281434,I280990);
not I_16402 (I281456,I281434);
and I_16403 (I281473,I281456,I280990);
nor I_16404 (I280938,I281015,I281473);
nand I_16405 (I281504,I281456,I281066);
nor I_16406 (I280932,I281326,I281504);
nand I_16407 (I280935,I281456,I281244);
nand I_16408 (I281549,I281066,I75870);
nor I_16409 (I280947,I281309,I281549);
not I_16410 (I281610,I2602);
DFFARX1 I_16411 (I6178,I2595,I281610,I281636,);
DFFARX1 I_16412 (I6175,I2595,I281610,I281653,);
not I_16413 (I281661,I281653);
not I_16414 (I281678,I6187);
nor I_16415 (I281695,I281678,I6184);
not I_16416 (I281712,I6193);
nor I_16417 (I281729,I281695,I6190);
nor I_16418 (I281746,I281653,I281729);
DFFARX1 I_16419 (I281746,I2595,I281610,I281596,);
nor I_16420 (I281777,I6190,I6184);
nand I_16421 (I281794,I281777,I6187);
DFFARX1 I_16422 (I281794,I2595,I281610,I281599,);
nor I_16423 (I281825,I281712,I6190);
nand I_16424 (I281842,I281825,I6181);
nor I_16425 (I281859,I281636,I281842);
DFFARX1 I_16426 (I281859,I2595,I281610,I281575,);
not I_16427 (I281890,I281842);
nand I_16428 (I281587,I281653,I281890);
DFFARX1 I_16429 (I281842,I2595,I281610,I281930,);
not I_16430 (I281938,I281930);
not I_16431 (I281955,I6190);
not I_16432 (I281972,I6181);
nor I_16433 (I281989,I281972,I6193);
nor I_16434 (I281602,I281938,I281989);
nor I_16435 (I282020,I281972,I6175);
and I_16436 (I282037,I282020,I6196);
or I_16437 (I282054,I282037,I6178);
DFFARX1 I_16438 (I282054,I2595,I281610,I282080,);
nor I_16439 (I281590,I282080,I281636);
not I_16440 (I282102,I282080);
and I_16441 (I282119,I282102,I281636);
nor I_16442 (I281584,I281661,I282119);
nand I_16443 (I282150,I282102,I281712);
nor I_16444 (I281578,I281972,I282150);
nand I_16445 (I281581,I282102,I281890);
nand I_16446 (I282195,I281712,I6181);
nor I_16447 (I281593,I281955,I282195);
not I_16448 (I282256,I2602);
DFFARX1 I_16449 (I349168,I2595,I282256,I282282,);
DFFARX1 I_16450 (I349174,I2595,I282256,I282299,);
not I_16451 (I282307,I282299);
not I_16452 (I282324,I349171);
nor I_16453 (I282341,I282324,I349150);
not I_16454 (I282358,I349153);
nor I_16455 (I282375,I282341,I349159);
nor I_16456 (I282392,I282299,I282375);
DFFARX1 I_16457 (I282392,I2595,I282256,I282242,);
nor I_16458 (I282423,I349159,I349150);
nand I_16459 (I282440,I282423,I349171);
DFFARX1 I_16460 (I282440,I2595,I282256,I282245,);
nor I_16461 (I282471,I282358,I349159);
nand I_16462 (I282488,I282471,I349153);
nor I_16463 (I282505,I282282,I282488);
DFFARX1 I_16464 (I282505,I2595,I282256,I282221,);
not I_16465 (I282536,I282488);
nand I_16466 (I282233,I282299,I282536);
DFFARX1 I_16467 (I282488,I2595,I282256,I282576,);
not I_16468 (I282584,I282576);
not I_16469 (I282601,I349159);
not I_16470 (I282618,I349162);
nor I_16471 (I282635,I282618,I349153);
nor I_16472 (I282248,I282584,I282635);
nor I_16473 (I282666,I282618,I349150);
and I_16474 (I282683,I282666,I349156);
or I_16475 (I282700,I282683,I349165);
DFFARX1 I_16476 (I282700,I2595,I282256,I282726,);
nor I_16477 (I282236,I282726,I282282);
not I_16478 (I282748,I282726);
and I_16479 (I282765,I282748,I282282);
nor I_16480 (I282230,I282307,I282765);
nand I_16481 (I282796,I282748,I282358);
nor I_16482 (I282224,I282618,I282796);
nand I_16483 (I282227,I282748,I282536);
nand I_16484 (I282841,I282358,I349162);
nor I_16485 (I282239,I282601,I282841);
not I_16486 (I282902,I2602);
DFFARX1 I_16487 (I314862,I2595,I282902,I282928,);
DFFARX1 I_16488 (I314844,I2595,I282902,I282945,);
not I_16489 (I282953,I282945);
not I_16490 (I282970,I314853);
nor I_16491 (I282987,I282970,I314865);
not I_16492 (I283004,I314847);
nor I_16493 (I283021,I282987,I314856);
nor I_16494 (I283038,I282945,I283021);
DFFARX1 I_16495 (I283038,I2595,I282902,I282888,);
nor I_16496 (I283069,I314856,I314865);
nand I_16497 (I283086,I283069,I314853);
DFFARX1 I_16498 (I283086,I2595,I282902,I282891,);
nor I_16499 (I283117,I283004,I314856);
nand I_16500 (I283134,I283117,I314868);
nor I_16501 (I283151,I282928,I283134);
DFFARX1 I_16502 (I283151,I2595,I282902,I282867,);
not I_16503 (I283182,I283134);
nand I_16504 (I282879,I282945,I283182);
DFFARX1 I_16505 (I283134,I2595,I282902,I283222,);
not I_16506 (I283230,I283222);
not I_16507 (I283247,I314856);
not I_16508 (I283264,I314844);
nor I_16509 (I283281,I283264,I314847);
nor I_16510 (I282894,I283230,I283281);
nor I_16511 (I283312,I283264,I314850);
and I_16512 (I283329,I283312,I314859);
or I_16513 (I283346,I283329,I314847);
DFFARX1 I_16514 (I283346,I2595,I282902,I283372,);
nor I_16515 (I282882,I283372,I282928);
not I_16516 (I283394,I283372);
and I_16517 (I283411,I283394,I282928);
nor I_16518 (I282876,I282953,I283411);
nand I_16519 (I283442,I283394,I283004);
nor I_16520 (I282870,I283264,I283442);
nand I_16521 (I282873,I283394,I283182);
nand I_16522 (I283487,I283004,I314844);
nor I_16523 (I282885,I283247,I283487);
not I_16524 (I283548,I2602);
DFFARX1 I_16525 (I220024,I2595,I283548,I283574,);
DFFARX1 I_16526 (I220018,I2595,I283548,I283591,);
not I_16527 (I283599,I283591);
not I_16528 (I283616,I220033);
nor I_16529 (I283633,I283616,I220018);
not I_16530 (I283650,I220027);
nor I_16531 (I283667,I283633,I220036);
nor I_16532 (I283684,I283591,I283667);
DFFARX1 I_16533 (I283684,I2595,I283548,I283534,);
nor I_16534 (I283715,I220036,I220018);
nand I_16535 (I283732,I283715,I220033);
DFFARX1 I_16536 (I283732,I2595,I283548,I283537,);
nor I_16537 (I283763,I283650,I220036);
nand I_16538 (I283780,I283763,I220021);
nor I_16539 (I283797,I283574,I283780);
DFFARX1 I_16540 (I283797,I2595,I283548,I283513,);
not I_16541 (I283828,I283780);
nand I_16542 (I283525,I283591,I283828);
DFFARX1 I_16543 (I283780,I2595,I283548,I283868,);
not I_16544 (I283876,I283868);
not I_16545 (I283893,I220036);
not I_16546 (I283910,I220030);
nor I_16547 (I283927,I283910,I220027);
nor I_16548 (I283540,I283876,I283927);
nor I_16549 (I283958,I283910,I220039);
and I_16550 (I283975,I283958,I220042);
or I_16551 (I283992,I283975,I220021);
DFFARX1 I_16552 (I283992,I2595,I283548,I284018,);
nor I_16553 (I283528,I284018,I283574);
not I_16554 (I284040,I284018);
and I_16555 (I284057,I284040,I283574);
nor I_16556 (I283522,I283599,I284057);
nand I_16557 (I284088,I284040,I283650);
nor I_16558 (I283516,I283910,I284088);
nand I_16559 (I283519,I284040,I283828);
nand I_16560 (I284133,I283650,I220030);
nor I_16561 (I283531,I283893,I284133);
not I_16562 (I284194,I2602);
DFFARX1 I_16563 (I81672,I2595,I284194,I284220,);
DFFARX1 I_16564 (I81678,I2595,I284194,I284237,);
not I_16565 (I284245,I284237);
not I_16566 (I284262,I81699);
nor I_16567 (I284279,I284262,I81687);
not I_16568 (I284296,I81696);
nor I_16569 (I284313,I284279,I81681);
nor I_16570 (I284330,I284237,I284313);
DFFARX1 I_16571 (I284330,I2595,I284194,I284180,);
nor I_16572 (I284361,I81681,I81687);
nand I_16573 (I284378,I284361,I81699);
DFFARX1 I_16574 (I284378,I2595,I284194,I284183,);
nor I_16575 (I284409,I284296,I81681);
nand I_16576 (I284426,I284409,I81672);
nor I_16577 (I284443,I284220,I284426);
DFFARX1 I_16578 (I284443,I2595,I284194,I284159,);
not I_16579 (I284474,I284426);
nand I_16580 (I284171,I284237,I284474);
DFFARX1 I_16581 (I284426,I2595,I284194,I284514,);
not I_16582 (I284522,I284514);
not I_16583 (I284539,I81681);
not I_16584 (I284556,I81684);
nor I_16585 (I284573,I284556,I81696);
nor I_16586 (I284186,I284522,I284573);
nor I_16587 (I284604,I284556,I81693);
and I_16588 (I284621,I284604,I81675);
or I_16589 (I284638,I284621,I81690);
DFFARX1 I_16590 (I284638,I2595,I284194,I284664,);
nor I_16591 (I284174,I284664,I284220);
not I_16592 (I284686,I284664);
and I_16593 (I284703,I284686,I284220);
nor I_16594 (I284168,I284245,I284703);
nand I_16595 (I284734,I284686,I284296);
nor I_16596 (I284162,I284556,I284734);
nand I_16597 (I284165,I284686,I284474);
nand I_16598 (I284779,I284296,I81684);
nor I_16599 (I284177,I284539,I284779);
not I_16600 (I284840,I2602);
DFFARX1 I_16601 (I223492,I2595,I284840,I284866,);
DFFARX1 I_16602 (I223486,I2595,I284840,I284883,);
not I_16603 (I284891,I284883);
not I_16604 (I284908,I223501);
nor I_16605 (I284925,I284908,I223486);
not I_16606 (I284942,I223495);
nor I_16607 (I284959,I284925,I223504);
nor I_16608 (I284976,I284883,I284959);
DFFARX1 I_16609 (I284976,I2595,I284840,I284826,);
nor I_16610 (I285007,I223504,I223486);
nand I_16611 (I285024,I285007,I223501);
DFFARX1 I_16612 (I285024,I2595,I284840,I284829,);
nor I_16613 (I285055,I284942,I223504);
nand I_16614 (I285072,I285055,I223489);
nor I_16615 (I285089,I284866,I285072);
DFFARX1 I_16616 (I285089,I2595,I284840,I284805,);
not I_16617 (I285120,I285072);
nand I_16618 (I284817,I284883,I285120);
DFFARX1 I_16619 (I285072,I2595,I284840,I285160,);
not I_16620 (I285168,I285160);
not I_16621 (I285185,I223504);
not I_16622 (I285202,I223498);
nor I_16623 (I285219,I285202,I223495);
nor I_16624 (I284832,I285168,I285219);
nor I_16625 (I285250,I285202,I223507);
and I_16626 (I285267,I285250,I223510);
or I_16627 (I285284,I285267,I223489);
DFFARX1 I_16628 (I285284,I2595,I284840,I285310,);
nor I_16629 (I284820,I285310,I284866);
not I_16630 (I285332,I285310);
and I_16631 (I285349,I285332,I284866);
nor I_16632 (I284814,I284891,I285349);
nand I_16633 (I285380,I285332,I284942);
nor I_16634 (I284808,I285202,I285380);
nand I_16635 (I284811,I285332,I285120);
nand I_16636 (I285425,I284942,I223498);
nor I_16637 (I284823,I285185,I285425);
not I_16638 (I285486,I2602);
DFFARX1 I_16639 (I4393,I2595,I285486,I285512,);
DFFARX1 I_16640 (I4390,I2595,I285486,I285529,);
not I_16641 (I285537,I285529);
not I_16642 (I285554,I4402);
nor I_16643 (I285571,I285554,I4399);
not I_16644 (I285588,I4408);
nor I_16645 (I285605,I285571,I4405);
nor I_16646 (I285622,I285529,I285605);
DFFARX1 I_16647 (I285622,I2595,I285486,I285472,);
nor I_16648 (I285653,I4405,I4399);
nand I_16649 (I285670,I285653,I4402);
DFFARX1 I_16650 (I285670,I2595,I285486,I285475,);
nor I_16651 (I285701,I285588,I4405);
nand I_16652 (I285718,I285701,I4396);
nor I_16653 (I285735,I285512,I285718);
DFFARX1 I_16654 (I285735,I2595,I285486,I285451,);
not I_16655 (I285766,I285718);
nand I_16656 (I285463,I285529,I285766);
DFFARX1 I_16657 (I285718,I2595,I285486,I285806,);
not I_16658 (I285814,I285806);
not I_16659 (I285831,I4405);
not I_16660 (I285848,I4396);
nor I_16661 (I285865,I285848,I4408);
nor I_16662 (I285478,I285814,I285865);
nor I_16663 (I285896,I285848,I4390);
and I_16664 (I285913,I285896,I4411);
or I_16665 (I285930,I285913,I4393);
DFFARX1 I_16666 (I285930,I2595,I285486,I285956,);
nor I_16667 (I285466,I285956,I285512);
not I_16668 (I285978,I285956);
and I_16669 (I285995,I285978,I285512);
nor I_16670 (I285460,I285537,I285995);
nand I_16671 (I286026,I285978,I285588);
nor I_16672 (I285454,I285848,I286026);
nand I_16673 (I285457,I285978,I285766);
nand I_16674 (I286071,I285588,I4396);
nor I_16675 (I285469,I285831,I286071);
not I_16676 (I286132,I2602);
DFFARX1 I_16677 (I292693,I2595,I286132,I286158,);
DFFARX1 I_16678 (I292696,I2595,I286132,I286175,);
not I_16679 (I286183,I286175);
not I_16680 (I286200,I292693);
nor I_16681 (I286217,I286200,I292705);
not I_16682 (I286234,I292714);
nor I_16683 (I286251,I286217,I292702);
nor I_16684 (I286268,I286175,I286251);
DFFARX1 I_16685 (I286268,I2595,I286132,I286118,);
nor I_16686 (I286299,I292702,I292705);
nand I_16687 (I286316,I286299,I292693);
DFFARX1 I_16688 (I286316,I2595,I286132,I286121,);
nor I_16689 (I286347,I286234,I292702);
nand I_16690 (I286364,I286347,I292708);
nor I_16691 (I286381,I286158,I286364);
DFFARX1 I_16692 (I286381,I2595,I286132,I286097,);
not I_16693 (I286412,I286364);
nand I_16694 (I286109,I286175,I286412);
DFFARX1 I_16695 (I286364,I2595,I286132,I286452,);
not I_16696 (I286460,I286452);
not I_16697 (I286477,I292702);
not I_16698 (I286494,I292699);
nor I_16699 (I286511,I286494,I292714);
nor I_16700 (I286124,I286460,I286511);
nor I_16701 (I286542,I286494,I292711);
and I_16702 (I286559,I286542,I292699);
or I_16703 (I286576,I286559,I292696);
DFFARX1 I_16704 (I286576,I2595,I286132,I286602,);
nor I_16705 (I286112,I286602,I286158);
not I_16706 (I286624,I286602);
and I_16707 (I286641,I286624,I286158);
nor I_16708 (I286106,I286183,I286641);
nand I_16709 (I286672,I286624,I286234);
nor I_16710 (I286100,I286494,I286672);
nand I_16711 (I286103,I286624,I286412);
nand I_16712 (I286717,I286234,I292699);
nor I_16713 (I286115,I286477,I286717);
not I_16714 (I286778,I2602);
DFFARX1 I_16715 (I388403,I2595,I286778,I286804,);
DFFARX1 I_16716 (I388427,I2595,I286778,I286821,);
not I_16717 (I286829,I286821);
not I_16718 (I286846,I388409);
nor I_16719 (I286863,I286846,I388418);
not I_16720 (I286880,I388403);
nor I_16721 (I286897,I286863,I388424);
nor I_16722 (I286914,I286821,I286897);
DFFARX1 I_16723 (I286914,I2595,I286778,I286764,);
nor I_16724 (I286945,I388424,I388418);
nand I_16725 (I286962,I286945,I388409);
DFFARX1 I_16726 (I286962,I2595,I286778,I286767,);
nor I_16727 (I286993,I286880,I388424);
nand I_16728 (I287010,I286993,I388421);
nor I_16729 (I287027,I286804,I287010);
DFFARX1 I_16730 (I287027,I2595,I286778,I286743,);
not I_16731 (I287058,I287010);
nand I_16732 (I286755,I286821,I287058);
DFFARX1 I_16733 (I287010,I2595,I286778,I287098,);
not I_16734 (I287106,I287098);
not I_16735 (I287123,I388424);
not I_16736 (I287140,I388415);
nor I_16737 (I287157,I287140,I388403);
nor I_16738 (I286770,I287106,I287157);
nor I_16739 (I287188,I287140,I388406);
and I_16740 (I287205,I287188,I388430);
or I_16741 (I287222,I287205,I388412);
DFFARX1 I_16742 (I287222,I2595,I286778,I287248,);
nor I_16743 (I286758,I287248,I286804);
not I_16744 (I287270,I287248);
and I_16745 (I287287,I287270,I286804);
nor I_16746 (I286752,I286829,I287287);
nand I_16747 (I287318,I287270,I286880);
nor I_16748 (I286746,I287140,I287318);
nand I_16749 (I286749,I287270,I287058);
nand I_16750 (I287363,I286880,I388415);
nor I_16751 (I286761,I287123,I287363);
not I_16752 (I287424,I2602);
DFFARX1 I_16753 (I358509,I2595,I287424,I287450,);
DFFARX1 I_16754 (I358503,I2595,I287424,I287467,);
not I_16755 (I287475,I287467);
not I_16756 (I287492,I358512);
nor I_16757 (I287509,I287492,I358524);
not I_16758 (I287526,I358506);
nor I_16759 (I287543,I287509,I358503);
nor I_16760 (I287560,I287467,I287543);
DFFARX1 I_16761 (I287560,I2595,I287424,I287410,);
nor I_16762 (I287591,I358503,I358524);
nand I_16763 (I287608,I287591,I358512);
DFFARX1 I_16764 (I287608,I2595,I287424,I287413,);
nor I_16765 (I287639,I287526,I358503);
nand I_16766 (I287656,I287639,I358500);
nor I_16767 (I287673,I287450,I287656);
DFFARX1 I_16768 (I287673,I2595,I287424,I287389,);
not I_16769 (I287704,I287656);
nand I_16770 (I287401,I287467,I287704);
DFFARX1 I_16771 (I287656,I2595,I287424,I287744,);
not I_16772 (I287752,I287744);
not I_16773 (I287769,I358503);
not I_16774 (I287786,I358521);
nor I_16775 (I287803,I287786,I358506);
nor I_16776 (I287416,I287752,I287803);
nor I_16777 (I287834,I287786,I358515);
and I_16778 (I287851,I287834,I358500);
or I_16779 (I287868,I287851,I358518);
DFFARX1 I_16780 (I287868,I2595,I287424,I287894,);
nor I_16781 (I287404,I287894,I287450);
not I_16782 (I287916,I287894);
and I_16783 (I287933,I287916,I287450);
nor I_16784 (I287398,I287475,I287933);
nand I_16785 (I287964,I287916,I287526);
nor I_16786 (I287392,I287786,I287964);
nand I_16787 (I287395,I287916,I287704);
nand I_16788 (I288009,I287526,I358521);
nor I_16789 (I287407,I287769,I288009);
not I_16790 (I288070,I2602);
DFFARX1 I_16791 (I46126,I2595,I288070,I288096,);
DFFARX1 I_16792 (I46129,I2595,I288070,I288113,);
not I_16793 (I288121,I288113);
not I_16794 (I288138,I46114);
nor I_16795 (I288155,I288138,I46108);
not I_16796 (I288172,I46117);
nor I_16797 (I288189,I288155,I46132);
nor I_16798 (I288206,I288113,I288189);
DFFARX1 I_16799 (I288206,I2595,I288070,I288056,);
nor I_16800 (I288237,I46132,I46108);
nand I_16801 (I288254,I288237,I46114);
DFFARX1 I_16802 (I288254,I2595,I288070,I288059,);
nor I_16803 (I288285,I288172,I46132);
nand I_16804 (I288302,I288285,I46135);
nor I_16805 (I288319,I288096,I288302);
DFFARX1 I_16806 (I288319,I2595,I288070,I288035,);
not I_16807 (I288350,I288302);
nand I_16808 (I288047,I288113,I288350);
DFFARX1 I_16809 (I288302,I2595,I288070,I288390,);
not I_16810 (I288398,I288390);
not I_16811 (I288415,I46132);
not I_16812 (I288432,I46111);
nor I_16813 (I288449,I288432,I46117);
nor I_16814 (I288062,I288398,I288449);
nor I_16815 (I288480,I288432,I46120);
and I_16816 (I288497,I288480,I46108);
or I_16817 (I288514,I288497,I46123);
DFFARX1 I_16818 (I288514,I2595,I288070,I288540,);
nor I_16819 (I288050,I288540,I288096);
not I_16820 (I288562,I288540);
and I_16821 (I288579,I288562,I288096);
nor I_16822 (I288044,I288121,I288579);
nand I_16823 (I288610,I288562,I288172);
nor I_16824 (I288038,I288432,I288610);
nand I_16825 (I288041,I288562,I288350);
nand I_16826 (I288655,I288172,I46111);
nor I_16827 (I288053,I288415,I288655);
not I_16828 (I288716,I2602);
DFFARX1 I_16829 (I219446,I2595,I288716,I288742,);
DFFARX1 I_16830 (I219440,I2595,I288716,I288759,);
not I_16831 (I288767,I288759);
not I_16832 (I288784,I219455);
nor I_16833 (I288801,I288784,I219440);
not I_16834 (I288818,I219449);
nor I_16835 (I288835,I288801,I219458);
nor I_16836 (I288852,I288759,I288835);
DFFARX1 I_16837 (I288852,I2595,I288716,I288702,);
nor I_16838 (I288883,I219458,I219440);
nand I_16839 (I288900,I288883,I219455);
DFFARX1 I_16840 (I288900,I2595,I288716,I288705,);
nor I_16841 (I288931,I288818,I219458);
nand I_16842 (I288948,I288931,I219443);
nor I_16843 (I288965,I288742,I288948);
DFFARX1 I_16844 (I288965,I2595,I288716,I288681,);
not I_16845 (I288996,I288948);
nand I_16846 (I288693,I288759,I288996);
DFFARX1 I_16847 (I288948,I2595,I288716,I289036,);
not I_16848 (I289044,I289036);
not I_16849 (I289061,I219458);
not I_16850 (I289078,I219452);
nor I_16851 (I289095,I289078,I219449);
nor I_16852 (I288708,I289044,I289095);
nor I_16853 (I289126,I289078,I219461);
and I_16854 (I289143,I289126,I219464);
or I_16855 (I289160,I289143,I219443);
DFFARX1 I_16856 (I289160,I2595,I288716,I289186,);
nor I_16857 (I288696,I289186,I288742);
not I_16858 (I289208,I289186);
and I_16859 (I289225,I289208,I288742);
nor I_16860 (I288690,I288767,I289225);
nand I_16861 (I289256,I289208,I288818);
nor I_16862 (I288684,I289078,I289256);
nand I_16863 (I288687,I289208,I288996);
nand I_16864 (I289301,I288818,I219452);
nor I_16865 (I288699,I289061,I289301);
not I_16866 (I289356,I2602);
DFFARX1 I_16867 (I19776,I2595,I289356,I289382,);
DFFARX1 I_16868 (I289382,I2595,I289356,I289399,);
not I_16869 (I289348,I289399);
not I_16870 (I289421,I289382);
DFFARX1 I_16871 (I19761,I2595,I289356,I289447,);
nand I_16872 (I289455,I289447,I19773);
not I_16873 (I289472,I19773);
not I_16874 (I289489,I19779);
nand I_16875 (I289506,I19767,I19758);
and I_16876 (I289523,I19767,I19758);
not I_16877 (I289540,I19764);
nand I_16878 (I289557,I289540,I289489);
nor I_16879 (I289330,I289557,I289455);
nor I_16880 (I289588,I289472,I289557);
nand I_16881 (I289333,I289523,I289588);
not I_16882 (I289619,I19770);
nor I_16883 (I289636,I289619,I19767);
nor I_16884 (I289653,I289636,I19764);
nor I_16885 (I289670,I289421,I289653);
DFFARX1 I_16886 (I289670,I2595,I289356,I289342,);
not I_16887 (I289701,I289636);
DFFARX1 I_16888 (I289701,I2595,I289356,I289345,);
and I_16889 (I289339,I289447,I289636);
nor I_16890 (I289746,I289619,I19758);
and I_16891 (I289763,I289746,I19782);
or I_16892 (I289780,I289763,I19761);
DFFARX1 I_16893 (I289780,I2595,I289356,I289806,);
nor I_16894 (I289814,I289806,I289540);
DFFARX1 I_16895 (I289814,I2595,I289356,I289327,);
nand I_16896 (I289845,I289806,I289447);
nand I_16897 (I289862,I289540,I289845);
nor I_16898 (I289336,I289862,I289506);
not I_16899 (I289917,I2602);
DFFARX1 I_16900 (I254443,I2595,I289917,I289943,);
DFFARX1 I_16901 (I289943,I2595,I289917,I289960,);
not I_16902 (I289909,I289960);
not I_16903 (I289982,I289943);
DFFARX1 I_16904 (I254470,I2595,I289917,I290008,);
nand I_16905 (I290016,I290008,I254461);
not I_16906 (I290033,I254461);
not I_16907 (I290050,I254443);
nand I_16908 (I290067,I254455,I254458);
and I_16909 (I290084,I254455,I254458);
not I_16910 (I290101,I254467);
nand I_16911 (I290118,I290101,I290050);
nor I_16912 (I289891,I290118,I290016);
nor I_16913 (I290149,I290033,I290118);
nand I_16914 (I289894,I290084,I290149);
not I_16915 (I290180,I254452);
nor I_16916 (I290197,I290180,I254455);
nor I_16917 (I290214,I290197,I254467);
nor I_16918 (I290231,I289982,I290214);
DFFARX1 I_16919 (I290231,I2595,I289917,I289903,);
not I_16920 (I290262,I290197);
DFFARX1 I_16921 (I290262,I2595,I289917,I289906,);
and I_16922 (I289900,I290008,I290197);
nor I_16923 (I290307,I290180,I254446);
and I_16924 (I290324,I290307,I254449);
or I_16925 (I290341,I290324,I254464);
DFFARX1 I_16926 (I290341,I2595,I289917,I290367,);
nor I_16927 (I290375,I290367,I290101);
DFFARX1 I_16928 (I290375,I2595,I289917,I289888,);
nand I_16929 (I290406,I290367,I290008);
nand I_16930 (I290423,I290101,I290406);
nor I_16931 (I289897,I290423,I290067);
not I_16932 (I290478,I2602);
DFFARX1 I_16933 (I228113,I2595,I290478,I290504,);
DFFARX1 I_16934 (I290504,I2595,I290478,I290521,);
not I_16935 (I290470,I290521);
not I_16936 (I290543,I290504);
DFFARX1 I_16937 (I228125,I2595,I290478,I290569,);
nand I_16938 (I290577,I290569,I228134);
not I_16939 (I290594,I228134);
not I_16940 (I290611,I228116);
nand I_16941 (I290628,I228119,I228110);
and I_16942 (I290645,I228119,I228110);
not I_16943 (I290662,I228128);
nand I_16944 (I290679,I290662,I290611);
nor I_16945 (I290452,I290679,I290577);
nor I_16946 (I290710,I290594,I290679);
nand I_16947 (I290455,I290645,I290710);
not I_16948 (I290741,I228131);
nor I_16949 (I290758,I290741,I228119);
nor I_16950 (I290775,I290758,I228128);
nor I_16951 (I290792,I290543,I290775);
DFFARX1 I_16952 (I290792,I2595,I290478,I290464,);
not I_16953 (I290823,I290758);
DFFARX1 I_16954 (I290823,I2595,I290478,I290467,);
and I_16955 (I290461,I290569,I290758);
nor I_16956 (I290868,I290741,I228110);
and I_16957 (I290885,I290868,I228122);
or I_16958 (I290902,I290885,I228113);
DFFARX1 I_16959 (I290902,I2595,I290478,I290928,);
nor I_16960 (I290936,I290928,I290662);
DFFARX1 I_16961 (I290936,I2595,I290478,I290449,);
nand I_16962 (I290967,I290928,I290569);
nand I_16963 (I290984,I290662,I290967);
nor I_16964 (I290458,I290984,I290628);
not I_16965 (I291039,I2602);
DFFARX1 I_16966 (I230380,I2595,I291039,I291065,);
DFFARX1 I_16967 (I291065,I2595,I291039,I291082,);
not I_16968 (I291031,I291082);
not I_16969 (I291104,I291065);
DFFARX1 I_16970 (I230377,I2595,I291039,I291130,);
nand I_16971 (I291138,I291130,I230392);
not I_16972 (I291155,I230392);
not I_16973 (I291172,I230389);
nand I_16974 (I291189,I230386,I230374);
and I_16975 (I291206,I230386,I230374);
not I_16976 (I291223,I230371);
nand I_16977 (I291240,I291223,I291172);
nor I_16978 (I291013,I291240,I291138);
nor I_16979 (I291271,I291155,I291240);
nand I_16980 (I291016,I291206,I291271);
not I_16981 (I291302,I230377);
nor I_16982 (I291319,I291302,I230386);
nor I_16983 (I291336,I291319,I230371);
nor I_16984 (I291353,I291104,I291336);
DFFARX1 I_16985 (I291353,I2595,I291039,I291025,);
not I_16986 (I291384,I291319);
DFFARX1 I_16987 (I291384,I2595,I291039,I291028,);
and I_16988 (I291022,I291130,I291319);
nor I_16989 (I291429,I291302,I230383);
and I_16990 (I291446,I291429,I230371);
or I_16991 (I291463,I291446,I230374);
DFFARX1 I_16992 (I291463,I2595,I291039,I291489,);
nor I_16993 (I291497,I291489,I291223);
DFFARX1 I_16994 (I291497,I2595,I291039,I291010,);
nand I_16995 (I291528,I291489,I291130);
nand I_16996 (I291545,I291223,I291528);
nor I_16997 (I291019,I291545,I291189);
not I_16998 (I291600,I2602);
DFFARX1 I_16999 (I351332,I2595,I291600,I291626,);
DFFARX1 I_17000 (I291626,I2595,I291600,I291643,);
not I_17001 (I291592,I291643);
not I_17002 (I291665,I291626);
DFFARX1 I_17003 (I351338,I2595,I291600,I291691,);
nand I_17004 (I291699,I291691,I351347);
not I_17005 (I291716,I351347);
not I_17006 (I291733,I351326);
nand I_17007 (I291750,I351329,I351329);
and I_17008 (I291767,I351329,I351329);
not I_17009 (I291784,I351341);
nand I_17010 (I291801,I291784,I291733);
nor I_17011 (I291574,I291801,I291699);
nor I_17012 (I291832,I291716,I291801);
nand I_17013 (I291577,I291767,I291832);
not I_17014 (I291863,I351335);
nor I_17015 (I291880,I291863,I351329);
nor I_17016 (I291897,I291880,I351341);
nor I_17017 (I291914,I291665,I291897);
DFFARX1 I_17018 (I291914,I2595,I291600,I291586,);
not I_17019 (I291945,I291880);
DFFARX1 I_17020 (I291945,I2595,I291600,I291589,);
and I_17021 (I291583,I291691,I291880);
nor I_17022 (I291990,I291863,I351350);
and I_17023 (I292007,I291990,I351326);
or I_17024 (I292024,I292007,I351344);
DFFARX1 I_17025 (I292024,I2595,I291600,I292050,);
nor I_17026 (I292058,I292050,I291784);
DFFARX1 I_17027 (I292058,I2595,I291600,I291571,);
nand I_17028 (I292089,I292050,I291691);
nand I_17029 (I292106,I291784,I292089);
nor I_17030 (I291580,I292106,I291750);
not I_17031 (I292161,I2602);
DFFARX1 I_17032 (I4991,I2595,I292161,I292187,);
DFFARX1 I_17033 (I292187,I2595,I292161,I292204,);
not I_17034 (I292153,I292204);
not I_17035 (I292226,I292187);
DFFARX1 I_17036 (I5003,I2595,I292161,I292252,);
nand I_17037 (I292260,I292252,I5000);
not I_17038 (I292277,I5000);
not I_17039 (I292294,I4991);
nand I_17040 (I292311,I4985,I4985);
and I_17041 (I292328,I4985,I4985);
not I_17042 (I292345,I5006);
nand I_17043 (I292362,I292345,I292294);
nor I_17044 (I292135,I292362,I292260);
nor I_17045 (I292393,I292277,I292362);
nand I_17046 (I292138,I292328,I292393);
not I_17047 (I292424,I4997);
nor I_17048 (I292441,I292424,I4985);
nor I_17049 (I292458,I292441,I5006);
nor I_17050 (I292475,I292226,I292458);
DFFARX1 I_17051 (I292475,I2595,I292161,I292147,);
not I_17052 (I292506,I292441);
DFFARX1 I_17053 (I292506,I2595,I292161,I292150,);
and I_17054 (I292144,I292252,I292441);
nor I_17055 (I292551,I292424,I4988);
and I_17056 (I292568,I292551,I4988);
or I_17057 (I292585,I292568,I4994);
DFFARX1 I_17058 (I292585,I2595,I292161,I292611,);
nor I_17059 (I292619,I292611,I292345);
DFFARX1 I_17060 (I292619,I2595,I292161,I292132,);
nand I_17061 (I292650,I292611,I292252);
nand I_17062 (I292667,I292345,I292650);
nor I_17063 (I292141,I292667,I292311);
not I_17064 (I292722,I2602);
DFFARX1 I_17065 (I366017,I2595,I292722,I292748,);
DFFARX1 I_17066 (I292748,I2595,I292722,I292765,);
not I_17067 (I292714,I292765);
not I_17068 (I292787,I292748);
DFFARX1 I_17069 (I366014,I2595,I292722,I292813,);
nand I_17070 (I292821,I292813,I366020);
not I_17071 (I292838,I366020);
not I_17072 (I292855,I366029);
nand I_17073 (I292872,I366023,I366017);
and I_17074 (I292889,I366023,I366017);
not I_17075 (I292906,I366035);
nand I_17076 (I292923,I292906,I292855);
nor I_17077 (I292696,I292923,I292821);
nor I_17078 (I292954,I292838,I292923);
nand I_17079 (I292699,I292889,I292954);
not I_17080 (I292985,I366032);
nor I_17081 (I293002,I292985,I366023);
nor I_17082 (I293019,I293002,I366035);
nor I_17083 (I293036,I292787,I293019);
DFFARX1 I_17084 (I293036,I2595,I292722,I292708,);
not I_17085 (I293067,I293002);
DFFARX1 I_17086 (I293067,I2595,I292722,I292711,);
and I_17087 (I292705,I292813,I293002);
nor I_17088 (I293112,I292985,I366026);
and I_17089 (I293129,I293112,I366038);
or I_17090 (I293146,I293129,I366014);
DFFARX1 I_17091 (I293146,I2595,I292722,I293172,);
nor I_17092 (I293180,I293172,I292906);
DFFARX1 I_17093 (I293180,I2595,I292722,I292693,);
nand I_17094 (I293211,I293172,I292813);
nand I_17095 (I293228,I292906,I293211);
nor I_17096 (I292702,I293228,I292872);
not I_17097 (I293283,I2602);
DFFARX1 I_17098 (I177246,I2595,I293283,I293309,);
DFFARX1 I_17099 (I293309,I2595,I293283,I293326,);
not I_17100 (I293275,I293326);
not I_17101 (I293348,I293309);
DFFARX1 I_17102 (I177261,I2595,I293283,I293374,);
nand I_17103 (I293382,I293374,I177252);
not I_17104 (I293399,I177252);
not I_17105 (I293416,I177258);
nand I_17106 (I293433,I177255,I177264);
and I_17107 (I293450,I177255,I177264);
not I_17108 (I293467,I177249);
nand I_17109 (I293484,I293467,I293416);
nor I_17110 (I293257,I293484,I293382);
nor I_17111 (I293515,I293399,I293484);
nand I_17112 (I293260,I293450,I293515);
not I_17113 (I293546,I177246);
nor I_17114 (I293563,I293546,I177255);
nor I_17115 (I293580,I293563,I177249);
nor I_17116 (I293597,I293348,I293580);
DFFARX1 I_17117 (I293597,I2595,I293283,I293269,);
not I_17118 (I293628,I293563);
DFFARX1 I_17119 (I293628,I2595,I293283,I293272,);
and I_17120 (I293266,I293374,I293563);
nor I_17121 (I293673,I293546,I177270);
and I_17122 (I293690,I293673,I177249);
or I_17123 (I293707,I293690,I177267);
DFFARX1 I_17124 (I293707,I2595,I293283,I293733,);
nor I_17125 (I293741,I293733,I293467);
DFFARX1 I_17126 (I293741,I2595,I293283,I293254,);
nand I_17127 (I293772,I293733,I293374);
nand I_17128 (I293789,I293467,I293772);
nor I_17129 (I293263,I293789,I293433);
not I_17130 (I293844,I2602);
DFFARX1 I_17131 (I148738,I2595,I293844,I293870,);
DFFARX1 I_17132 (I293870,I2595,I293844,I293887,);
not I_17133 (I293836,I293887);
not I_17134 (I293909,I293870);
DFFARX1 I_17135 (I148735,I2595,I293844,I293935,);
nand I_17136 (I293943,I293935,I148729);
not I_17137 (I293960,I148729);
not I_17138 (I293977,I148741);
nand I_17139 (I293994,I148744,I148723);
and I_17140 (I294011,I148744,I148723);
not I_17141 (I294028,I148720);
nand I_17142 (I294045,I294028,I293977);
nor I_17143 (I293818,I294045,I293943);
nor I_17144 (I294076,I293960,I294045);
nand I_17145 (I293821,I294011,I294076);
not I_17146 (I294107,I148726);
nor I_17147 (I294124,I294107,I148744);
nor I_17148 (I294141,I294124,I148720);
nor I_17149 (I294158,I293909,I294141);
DFFARX1 I_17150 (I294158,I2595,I293844,I293830,);
not I_17151 (I294189,I294124);
DFFARX1 I_17152 (I294189,I2595,I293844,I293833,);
and I_17153 (I293827,I293935,I294124);
nor I_17154 (I294234,I294107,I148720);
and I_17155 (I294251,I294234,I148732);
or I_17156 (I294268,I294251,I148723);
DFFARX1 I_17157 (I294268,I2595,I293844,I294294,);
nor I_17158 (I294302,I294294,I294028);
DFFARX1 I_17159 (I294302,I2595,I293844,I293815,);
nand I_17160 (I294333,I294294,I293935);
nand I_17161 (I294350,I294028,I294333);
nor I_17162 (I293824,I294350,I293994);
not I_17163 (I294405,I2602);
DFFARX1 I_17164 (I166842,I2595,I294405,I294431,);
DFFARX1 I_17165 (I294431,I2595,I294405,I294448,);
not I_17166 (I294397,I294448);
not I_17167 (I294470,I294431);
DFFARX1 I_17168 (I166857,I2595,I294405,I294496,);
nand I_17169 (I294504,I294496,I166848);
not I_17170 (I294521,I166848);
not I_17171 (I294538,I166854);
nand I_17172 (I294555,I166851,I166860);
and I_17173 (I294572,I166851,I166860);
not I_17174 (I294589,I166845);
nand I_17175 (I294606,I294589,I294538);
nor I_17176 (I294379,I294606,I294504);
nor I_17177 (I294637,I294521,I294606);
nand I_17178 (I294382,I294572,I294637);
not I_17179 (I294668,I166842);
nor I_17180 (I294685,I294668,I166851);
nor I_17181 (I294702,I294685,I166845);
nor I_17182 (I294719,I294470,I294702);
DFFARX1 I_17183 (I294719,I2595,I294405,I294391,);
not I_17184 (I294750,I294685);
DFFARX1 I_17185 (I294750,I2595,I294405,I294394,);
and I_17186 (I294388,I294496,I294685);
nor I_17187 (I294795,I294668,I166866);
and I_17188 (I294812,I294795,I166845);
or I_17189 (I294829,I294812,I166863);
DFFARX1 I_17190 (I294829,I2595,I294405,I294855,);
nor I_17191 (I294863,I294855,I294589);
DFFARX1 I_17192 (I294863,I2595,I294405,I294376,);
nand I_17193 (I294894,I294855,I294496);
nand I_17194 (I294911,I294589,I294894);
nor I_17195 (I294385,I294911,I294555);
not I_17196 (I294966,I2602);
DFFARX1 I_17197 (I329309,I2595,I294966,I294992,);
DFFARX1 I_17198 (I294992,I2595,I294966,I295009,);
not I_17199 (I294958,I295009);
not I_17200 (I295031,I294992);
DFFARX1 I_17201 (I329300,I2595,I294966,I295057,);
nand I_17202 (I295065,I295057,I329297);
not I_17203 (I295082,I329297);
not I_17204 (I295099,I329306);
nand I_17205 (I295116,I329315,I329297);
and I_17206 (I295133,I329315,I329297);
not I_17207 (I295150,I329294);
nand I_17208 (I295167,I295150,I295099);
nor I_17209 (I294940,I295167,I295065);
nor I_17210 (I295198,I295082,I295167);
nand I_17211 (I294943,I295133,I295198);
not I_17212 (I295229,I329303);
nor I_17213 (I295246,I295229,I329315);
nor I_17214 (I295263,I295246,I329294);
nor I_17215 (I295280,I295031,I295263);
DFFARX1 I_17216 (I295280,I2595,I294966,I294952,);
not I_17217 (I295311,I295246);
DFFARX1 I_17218 (I295311,I2595,I294966,I294955,);
and I_17219 (I294949,I295057,I295246);
nor I_17220 (I295356,I295229,I329318);
and I_17221 (I295373,I295356,I329294);
or I_17222 (I295390,I295373,I329312);
DFFARX1 I_17223 (I295390,I2595,I294966,I295416,);
nor I_17224 (I295424,I295416,I295150);
DFFARX1 I_17225 (I295424,I2595,I294966,I294937,);
nand I_17226 (I295455,I295416,I295057);
nand I_17227 (I295472,I295150,I295455);
nor I_17228 (I294946,I295472,I295116);
not I_17229 (I295527,I2602);
DFFARX1 I_17230 (I383063,I2595,I295527,I295553,);
DFFARX1 I_17231 (I295553,I2595,I295527,I295570,);
not I_17232 (I295519,I295570);
not I_17233 (I295592,I295553);
DFFARX1 I_17234 (I383057,I2595,I295527,I295618,);
nand I_17235 (I295626,I295618,I383048);
not I_17236 (I295643,I383048);
not I_17237 (I295660,I383075);
nand I_17238 (I295677,I383060,I383069);
and I_17239 (I295694,I383060,I383069);
not I_17240 (I295711,I383054);
nand I_17241 (I295728,I295711,I295660);
nor I_17242 (I295501,I295728,I295626);
nor I_17243 (I295759,I295643,I295728);
nand I_17244 (I295504,I295694,I295759);
not I_17245 (I295790,I383072);
nor I_17246 (I295807,I295790,I383060);
nor I_17247 (I295824,I295807,I383054);
nor I_17248 (I295841,I295592,I295824);
DFFARX1 I_17249 (I295841,I2595,I295527,I295513,);
not I_17250 (I295872,I295807);
DFFARX1 I_17251 (I295872,I2595,I295527,I295516,);
and I_17252 (I295510,I295618,I295807);
nor I_17253 (I295917,I295790,I383066);
and I_17254 (I295934,I295917,I383048);
or I_17255 (I295951,I295934,I383051);
DFFARX1 I_17256 (I295951,I2595,I295527,I295977,);
nor I_17257 (I295985,I295977,I295711);
DFFARX1 I_17258 (I295985,I2595,I295527,I295498,);
nand I_17259 (I296016,I295977,I295618);
nand I_17260 (I296033,I295711,I296016);
nor I_17261 (I295507,I296033,I295677);
not I_17262 (I296088,I2602);
DFFARX1 I_17263 (I47917,I2595,I296088,I296114,);
DFFARX1 I_17264 (I296114,I2595,I296088,I296131,);
not I_17265 (I296080,I296131);
not I_17266 (I296153,I296114);
DFFARX1 I_17267 (I47899,I2595,I296088,I296179,);
nand I_17268 (I296187,I296179,I47893);
not I_17269 (I296204,I47893);
not I_17270 (I296221,I47896);
nand I_17271 (I296238,I47911,I47902);
and I_17272 (I296255,I47911,I47902);
not I_17273 (I296272,I47914);
nand I_17274 (I296289,I296272,I296221);
nor I_17275 (I296062,I296289,I296187);
nor I_17276 (I296320,I296204,I296289);
nand I_17277 (I296065,I296255,I296320);
not I_17278 (I296351,I47908);
nor I_17279 (I296368,I296351,I47911);
nor I_17280 (I296385,I296368,I47914);
nor I_17281 (I296402,I296153,I296385);
DFFARX1 I_17282 (I296402,I2595,I296088,I296074,);
not I_17283 (I296433,I296368);
DFFARX1 I_17284 (I296433,I2595,I296088,I296077,);
and I_17285 (I296071,I296179,I296368);
nor I_17286 (I296478,I296351,I47920);
and I_17287 (I296495,I296478,I47893);
or I_17288 (I296512,I296495,I47905);
DFFARX1 I_17289 (I296512,I2595,I296088,I296538,);
nor I_17290 (I296546,I296538,I296272);
DFFARX1 I_17291 (I296546,I2595,I296088,I296059,);
nand I_17292 (I296577,I296538,I296179);
nand I_17293 (I296594,I296272,I296577);
nor I_17294 (I296068,I296594,I296238);
not I_17295 (I296649,I2602);
DFFARX1 I_17296 (I141003,I2595,I296649,I296675,);
DFFARX1 I_17297 (I296675,I2595,I296649,I296692,);
not I_17298 (I296641,I296692);
not I_17299 (I296714,I296675);
DFFARX1 I_17300 (I141000,I2595,I296649,I296740,);
nand I_17301 (I296748,I296740,I140994);
not I_17302 (I296765,I140994);
not I_17303 (I296782,I141006);
nand I_17304 (I296799,I141009,I140988);
and I_17305 (I296816,I141009,I140988);
not I_17306 (I296833,I140985);
nand I_17307 (I296850,I296833,I296782);
nor I_17308 (I296623,I296850,I296748);
nor I_17309 (I296881,I296765,I296850);
nand I_17310 (I296626,I296816,I296881);
not I_17311 (I296912,I140991);
nor I_17312 (I296929,I296912,I141009);
nor I_17313 (I296946,I296929,I140985);
nor I_17314 (I296963,I296714,I296946);
DFFARX1 I_17315 (I296963,I2595,I296649,I296635,);
not I_17316 (I296994,I296929);
DFFARX1 I_17317 (I296994,I2595,I296649,I296638,);
and I_17318 (I296632,I296740,I296929);
nor I_17319 (I297039,I296912,I140985);
and I_17320 (I297056,I297039,I140997);
or I_17321 (I297073,I297056,I140988);
DFFARX1 I_17322 (I297073,I2595,I296649,I297099,);
nor I_17323 (I297107,I297099,I296833);
DFFARX1 I_17324 (I297107,I2595,I296649,I296620,);
nand I_17325 (I297138,I297099,I296740);
nand I_17326 (I297155,I296833,I297138);
nor I_17327 (I296629,I297155,I296799);
not I_17328 (I297210,I2602);
DFFARX1 I_17329 (I357925,I2595,I297210,I297236,);
DFFARX1 I_17330 (I297236,I2595,I297210,I297253,);
not I_17331 (I297202,I297253);
not I_17332 (I297275,I297236);
DFFARX1 I_17333 (I357922,I2595,I297210,I297301,);
nand I_17334 (I297309,I297301,I357928);
not I_17335 (I297326,I357928);
not I_17336 (I297343,I357937);
nand I_17337 (I297360,I357931,I357925);
and I_17338 (I297377,I357931,I357925);
not I_17339 (I297394,I357943);
nand I_17340 (I297411,I297394,I297343);
nor I_17341 (I297184,I297411,I297309);
nor I_17342 (I297442,I297326,I297411);
nand I_17343 (I297187,I297377,I297442);
not I_17344 (I297473,I357940);
nor I_17345 (I297490,I297473,I357931);
nor I_17346 (I297507,I297490,I357943);
nor I_17347 (I297524,I297275,I297507);
DFFARX1 I_17348 (I297524,I2595,I297210,I297196,);
not I_17349 (I297555,I297490);
DFFARX1 I_17350 (I297555,I2595,I297210,I297199,);
and I_17351 (I297193,I297301,I297490);
nor I_17352 (I297600,I297473,I357934);
and I_17353 (I297617,I297600,I357946);
or I_17354 (I297634,I297617,I357922);
DFFARX1 I_17355 (I297634,I2595,I297210,I297660,);
nor I_17356 (I297668,I297660,I297394);
DFFARX1 I_17357 (I297668,I2595,I297210,I297181,);
nand I_17358 (I297699,I297660,I297301);
nand I_17359 (I297716,I297394,I297699);
nor I_17360 (I297190,I297716,I297360);
not I_17361 (I297771,I2602);
DFFARX1 I_17362 (I185341,I2595,I297771,I297797,);
DFFARX1 I_17363 (I297797,I2595,I297771,I297814,);
not I_17364 (I297763,I297814);
not I_17365 (I297836,I297797);
DFFARX1 I_17366 (I185353,I2595,I297771,I297862,);
nand I_17367 (I297870,I297862,I185362);
not I_17368 (I297887,I185362);
not I_17369 (I297904,I185344);
nand I_17370 (I297921,I185347,I185338);
and I_17371 (I297938,I185347,I185338);
not I_17372 (I297955,I185356);
nand I_17373 (I297972,I297955,I297904);
nor I_17374 (I297745,I297972,I297870);
nor I_17375 (I298003,I297887,I297972);
nand I_17376 (I297748,I297938,I298003);
not I_17377 (I298034,I185359);
nor I_17378 (I298051,I298034,I185347);
nor I_17379 (I298068,I298051,I185356);
nor I_17380 (I298085,I297836,I298068);
DFFARX1 I_17381 (I298085,I2595,I297771,I297757,);
not I_17382 (I298116,I298051);
DFFARX1 I_17383 (I298116,I2595,I297771,I297760,);
and I_17384 (I297754,I297862,I298051);
nor I_17385 (I298161,I298034,I185338);
and I_17386 (I298178,I298161,I185350);
or I_17387 (I298195,I298178,I185341);
DFFARX1 I_17388 (I298195,I2595,I297771,I298221,);
nor I_17389 (I298229,I298221,I297955);
DFFARX1 I_17390 (I298229,I2595,I297771,I297742,);
nand I_17391 (I298260,I298221,I297862);
nand I_17392 (I298277,I297955,I298260);
nor I_17393 (I297751,I298277,I297921);
not I_17394 (I298332,I2602);
DFFARX1 I_17395 (I11344,I2595,I298332,I298358,);
DFFARX1 I_17396 (I298358,I2595,I298332,I298375,);
not I_17397 (I298324,I298375);
not I_17398 (I298397,I298358);
DFFARX1 I_17399 (I11329,I2595,I298332,I298423,);
nand I_17400 (I298431,I298423,I11341);
not I_17401 (I298448,I11341);
not I_17402 (I298465,I11347);
nand I_17403 (I298482,I11335,I11326);
and I_17404 (I298499,I11335,I11326);
not I_17405 (I298516,I11332);
nand I_17406 (I298533,I298516,I298465);
nor I_17407 (I298306,I298533,I298431);
nor I_17408 (I298564,I298448,I298533);
nand I_17409 (I298309,I298499,I298564);
not I_17410 (I298595,I11338);
nor I_17411 (I298612,I298595,I11335);
nor I_17412 (I298629,I298612,I11332);
nor I_17413 (I298646,I298397,I298629);
DFFARX1 I_17414 (I298646,I2595,I298332,I298318,);
not I_17415 (I298677,I298612);
DFFARX1 I_17416 (I298677,I2595,I298332,I298321,);
and I_17417 (I298315,I298423,I298612);
nor I_17418 (I298722,I298595,I11326);
and I_17419 (I298739,I298722,I11350);
or I_17420 (I298756,I298739,I11329);
DFFARX1 I_17421 (I298756,I2595,I298332,I298782,);
nor I_17422 (I298790,I298782,I298516);
DFFARX1 I_17423 (I298790,I2595,I298332,I298303,);
nand I_17424 (I298821,I298782,I298423);
nand I_17425 (I298838,I298516,I298821);
nor I_17426 (I298312,I298838,I298482);
not I_17427 (I298893,I2602);
DFFARX1 I_17428 (I182451,I2595,I298893,I298919,);
DFFARX1 I_17429 (I298919,I2595,I298893,I298936,);
not I_17430 (I298885,I298936);
not I_17431 (I298958,I298919);
DFFARX1 I_17432 (I182463,I2595,I298893,I298984,);
nand I_17433 (I298992,I298984,I182472);
not I_17434 (I299009,I182472);
not I_17435 (I299026,I182454);
nand I_17436 (I299043,I182457,I182448);
and I_17437 (I299060,I182457,I182448);
not I_17438 (I299077,I182466);
nand I_17439 (I299094,I299077,I299026);
nor I_17440 (I298867,I299094,I298992);
nor I_17441 (I299125,I299009,I299094);
nand I_17442 (I298870,I299060,I299125);
not I_17443 (I299156,I182469);
nor I_17444 (I299173,I299156,I182457);
nor I_17445 (I299190,I299173,I182466);
nor I_17446 (I299207,I298958,I299190);
DFFARX1 I_17447 (I299207,I2595,I298893,I298879,);
not I_17448 (I299238,I299173);
DFFARX1 I_17449 (I299238,I2595,I298893,I298882,);
and I_17450 (I298876,I298984,I299173);
nor I_17451 (I299283,I299156,I182448);
and I_17452 (I299300,I299283,I182460);
or I_17453 (I299317,I299300,I182451);
DFFARX1 I_17454 (I299317,I2595,I298893,I299343,);
nor I_17455 (I299351,I299343,I299077);
DFFARX1 I_17456 (I299351,I2595,I298893,I298864,);
nand I_17457 (I299382,I299343,I298984);
nand I_17458 (I299399,I299077,I299382);
nor I_17459 (I298873,I299399,I299043);
not I_17460 (I299454,I2602);
DFFARX1 I_17461 (I207305,I2595,I299454,I299480,);
DFFARX1 I_17462 (I299480,I2595,I299454,I299497,);
not I_17463 (I299446,I299497);
not I_17464 (I299519,I299480);
DFFARX1 I_17465 (I207317,I2595,I299454,I299545,);
nand I_17466 (I299553,I299545,I207326);
not I_17467 (I299570,I207326);
not I_17468 (I299587,I207308);
nand I_17469 (I299604,I207311,I207302);
and I_17470 (I299621,I207311,I207302);
not I_17471 (I299638,I207320);
nand I_17472 (I299655,I299638,I299587);
nor I_17473 (I299428,I299655,I299553);
nor I_17474 (I299686,I299570,I299655);
nand I_17475 (I299431,I299621,I299686);
not I_17476 (I299717,I207323);
nor I_17477 (I299734,I299717,I207311);
nor I_17478 (I299751,I299734,I207320);
nor I_17479 (I299768,I299519,I299751);
DFFARX1 I_17480 (I299768,I2595,I299454,I299440,);
not I_17481 (I299799,I299734);
DFFARX1 I_17482 (I299799,I2595,I299454,I299443,);
and I_17483 (I299437,I299545,I299734);
nor I_17484 (I299844,I299717,I207302);
and I_17485 (I299861,I299844,I207314);
or I_17486 (I299878,I299861,I207305);
DFFARX1 I_17487 (I299878,I2595,I299454,I299904,);
nor I_17488 (I299912,I299904,I299638);
DFFARX1 I_17489 (I299912,I2595,I299454,I299425,);
nand I_17490 (I299943,I299904,I299545);
nand I_17491 (I299960,I299638,I299943);
nor I_17492 (I299434,I299960,I299604);
not I_17493 (I300015,I2602);
DFFARX1 I_17494 (I2292,I2595,I300015,I300041,);
DFFARX1 I_17495 (I300041,I2595,I300015,I300058,);
not I_17496 (I300007,I300058);
not I_17497 (I300080,I300041);
DFFARX1 I_17498 (I1972,I2595,I300015,I300106,);
nand I_17499 (I300114,I300106,I2084);
not I_17500 (I300131,I2084);
not I_17501 (I300148,I1572);
nand I_17502 (I300165,I2108,I2244);
and I_17503 (I300182,I2108,I2244);
not I_17504 (I300199,I1780);
nand I_17505 (I300216,I300199,I300148);
nor I_17506 (I299989,I300216,I300114);
nor I_17507 (I300247,I300131,I300216);
nand I_17508 (I299992,I300182,I300247);
not I_17509 (I300278,I1516);
nor I_17510 (I300295,I300278,I2108);
nor I_17511 (I300312,I300295,I1780);
nor I_17512 (I300329,I300080,I300312);
DFFARX1 I_17513 (I300329,I2595,I300015,I300001,);
not I_17514 (I300360,I300295);
DFFARX1 I_17515 (I300360,I2595,I300015,I300004,);
and I_17516 (I299998,I300106,I300295);
nor I_17517 (I300405,I300278,I2092);
and I_17518 (I300422,I300405,I2356);
or I_17519 (I300439,I300422,I2364);
DFFARX1 I_17520 (I300439,I2595,I300015,I300465,);
nor I_17521 (I300473,I300465,I300199);
DFFARX1 I_17522 (I300473,I2595,I300015,I299986,);
nand I_17523 (I300504,I300465,I300106);
nand I_17524 (I300521,I300199,I300504);
nor I_17525 (I299995,I300521,I300165);
not I_17526 (I300576,I2602);
DFFARX1 I_17527 (I229269,I2595,I300576,I300602,);
DFFARX1 I_17528 (I300602,I2595,I300576,I300619,);
not I_17529 (I300568,I300619);
not I_17530 (I300641,I300602);
DFFARX1 I_17531 (I229281,I2595,I300576,I300667,);
nand I_17532 (I300675,I300667,I229290);
not I_17533 (I300692,I229290);
not I_17534 (I300709,I229272);
nand I_17535 (I300726,I229275,I229266);
and I_17536 (I300743,I229275,I229266);
not I_17537 (I300760,I229284);
nand I_17538 (I300777,I300760,I300709);
nor I_17539 (I300550,I300777,I300675);
nor I_17540 (I300808,I300692,I300777);
nand I_17541 (I300553,I300743,I300808);
not I_17542 (I300839,I229287);
nor I_17543 (I300856,I300839,I229275);
nor I_17544 (I300873,I300856,I229284);
nor I_17545 (I300890,I300641,I300873);
DFFARX1 I_17546 (I300890,I2595,I300576,I300562,);
not I_17547 (I300921,I300856);
DFFARX1 I_17548 (I300921,I2595,I300576,I300565,);
and I_17549 (I300559,I300667,I300856);
nor I_17550 (I300966,I300839,I229266);
and I_17551 (I300983,I300966,I229278);
or I_17552 (I301000,I300983,I229269);
DFFARX1 I_17553 (I301000,I2595,I300576,I301026,);
nor I_17554 (I301034,I301026,I300760);
DFFARX1 I_17555 (I301034,I2595,I300576,I300547,);
nand I_17556 (I301065,I301026,I300667);
nand I_17557 (I301082,I300760,I301065);
nor I_17558 (I300556,I301082,I300726);
not I_17559 (I301137,I2602);
DFFARX1 I_17560 (I281575,I2595,I301137,I301163,);
DFFARX1 I_17561 (I301163,I2595,I301137,I301180,);
not I_17562 (I301129,I301180);
not I_17563 (I301202,I301163);
DFFARX1 I_17564 (I281602,I2595,I301137,I301228,);
nand I_17565 (I301236,I301228,I281593);
not I_17566 (I301253,I281593);
not I_17567 (I301270,I281575);
nand I_17568 (I301287,I281587,I281590);
and I_17569 (I301304,I281587,I281590);
not I_17570 (I301321,I281599);
nand I_17571 (I301338,I301321,I301270);
nor I_17572 (I301111,I301338,I301236);
nor I_17573 (I301369,I301253,I301338);
nand I_17574 (I301114,I301304,I301369);
not I_17575 (I301400,I281584);
nor I_17576 (I301417,I301400,I281587);
nor I_17577 (I301434,I301417,I281599);
nor I_17578 (I301451,I301202,I301434);
DFFARX1 I_17579 (I301451,I2595,I301137,I301123,);
not I_17580 (I301482,I301417);
DFFARX1 I_17581 (I301482,I2595,I301137,I301126,);
and I_17582 (I301120,I301228,I301417);
nor I_17583 (I301527,I301400,I281578);
and I_17584 (I301544,I301527,I281581);
or I_17585 (I301561,I301544,I281596);
DFFARX1 I_17586 (I301561,I2595,I301137,I301587,);
nor I_17587 (I301595,I301587,I301321);
DFFARX1 I_17588 (I301595,I2595,I301137,I301108,);
nand I_17589 (I301626,I301587,I301228);
nand I_17590 (I301643,I301321,I301626);
nor I_17591 (I301117,I301643,I301287);
not I_17592 (I301698,I2602);
DFFARX1 I_17593 (I243028,I2595,I301698,I301724,);
DFFARX1 I_17594 (I301724,I2595,I301698,I301741,);
not I_17595 (I301690,I301741);
not I_17596 (I301763,I301724);
DFFARX1 I_17597 (I243025,I2595,I301698,I301789,);
nand I_17598 (I301797,I301789,I243040);
not I_17599 (I301814,I243040);
not I_17600 (I301831,I243037);
nand I_17601 (I301848,I243034,I243022);
and I_17602 (I301865,I243034,I243022);
not I_17603 (I301882,I243019);
nand I_17604 (I301899,I301882,I301831);
nor I_17605 (I301672,I301899,I301797);
nor I_17606 (I301930,I301814,I301899);
nand I_17607 (I301675,I301865,I301930);
not I_17608 (I301961,I243025);
nor I_17609 (I301978,I301961,I243034);
nor I_17610 (I301995,I301978,I243019);
nor I_17611 (I302012,I301763,I301995);
DFFARX1 I_17612 (I302012,I2595,I301698,I301684,);
not I_17613 (I302043,I301978);
DFFARX1 I_17614 (I302043,I2595,I301698,I301687,);
and I_17615 (I301681,I301789,I301978);
nor I_17616 (I302088,I301961,I243031);
and I_17617 (I302105,I302088,I243019);
or I_17618 (I302122,I302105,I243022);
DFFARX1 I_17619 (I302122,I2595,I301698,I302148,);
nor I_17620 (I302156,I302148,I301882);
DFFARX1 I_17621 (I302156,I2595,I301698,I301669,);
nand I_17622 (I302187,I302148,I301789);
nand I_17623 (I302204,I301882,I302187);
nor I_17624 (I301678,I302204,I301848);
not I_17625 (I302259,I2602);
DFFARX1 I_17626 (I266071,I2595,I302259,I302285,);
DFFARX1 I_17627 (I302285,I2595,I302259,I302302,);
not I_17628 (I302251,I302302);
not I_17629 (I302324,I302285);
DFFARX1 I_17630 (I266098,I2595,I302259,I302350,);
nand I_17631 (I302358,I302350,I266089);
not I_17632 (I302375,I266089);
not I_17633 (I302392,I266071);
nand I_17634 (I302409,I266083,I266086);
and I_17635 (I302426,I266083,I266086);
not I_17636 (I302443,I266095);
nand I_17637 (I302460,I302443,I302392);
nor I_17638 (I302233,I302460,I302358);
nor I_17639 (I302491,I302375,I302460);
nand I_17640 (I302236,I302426,I302491);
not I_17641 (I302522,I266080);
nor I_17642 (I302539,I302522,I266083);
nor I_17643 (I302556,I302539,I266095);
nor I_17644 (I302573,I302324,I302556);
DFFARX1 I_17645 (I302573,I2595,I302259,I302245,);
not I_17646 (I302604,I302539);
DFFARX1 I_17647 (I302604,I2595,I302259,I302248,);
and I_17648 (I302242,I302350,I302539);
nor I_17649 (I302649,I302522,I266074);
and I_17650 (I302666,I302649,I266077);
or I_17651 (I302683,I302666,I266092);
DFFARX1 I_17652 (I302683,I2595,I302259,I302709,);
nor I_17653 (I302717,I302709,I302443);
DFFARX1 I_17654 (I302717,I2595,I302259,I302230,);
nand I_17655 (I302748,I302709,I302350);
nand I_17656 (I302765,I302443,I302748);
nor I_17657 (I302239,I302765,I302409);
not I_17658 (I302820,I2602);
DFFARX1 I_17659 (I310235,I2595,I302820,I302846,);
DFFARX1 I_17660 (I302846,I2595,I302820,I302863,);
not I_17661 (I302812,I302863);
not I_17662 (I302885,I302846);
DFFARX1 I_17663 (I310226,I2595,I302820,I302911,);
nand I_17664 (I302919,I302911,I310223);
not I_17665 (I302936,I310223);
not I_17666 (I302953,I310232);
nand I_17667 (I302970,I310241,I310223);
and I_17668 (I302987,I310241,I310223);
not I_17669 (I303004,I310220);
nand I_17670 (I303021,I303004,I302953);
nor I_17671 (I302794,I303021,I302919);
nor I_17672 (I303052,I302936,I303021);
nand I_17673 (I302797,I302987,I303052);
not I_17674 (I303083,I310229);
nor I_17675 (I303100,I303083,I310241);
nor I_17676 (I303117,I303100,I310220);
nor I_17677 (I303134,I302885,I303117);
DFFARX1 I_17678 (I303134,I2595,I302820,I302806,);
not I_17679 (I303165,I303100);
DFFARX1 I_17680 (I303165,I2595,I302820,I302809,);
and I_17681 (I302803,I302911,I303100);
nor I_17682 (I303210,I303083,I310244);
and I_17683 (I303227,I303210,I310220);
or I_17684 (I303244,I303227,I310238);
DFFARX1 I_17685 (I303244,I2595,I302820,I303270,);
nor I_17686 (I303278,I303270,I303004);
DFFARX1 I_17687 (I303278,I2595,I302820,I302791,);
nand I_17688 (I303309,I303270,I302911);
nand I_17689 (I303326,I303004,I303309);
nor I_17690 (I302800,I303326,I302970);
not I_17691 (I303381,I2602);
DFFARX1 I_17692 (I166264,I2595,I303381,I303407,);
DFFARX1 I_17693 (I303407,I2595,I303381,I303424,);
not I_17694 (I303373,I303424);
not I_17695 (I303446,I303407);
DFFARX1 I_17696 (I166279,I2595,I303381,I303472,);
nand I_17697 (I303480,I303472,I166270);
not I_17698 (I303497,I166270);
not I_17699 (I303514,I166276);
nand I_17700 (I303531,I166273,I166282);
and I_17701 (I303548,I166273,I166282);
not I_17702 (I303565,I166267);
nand I_17703 (I303582,I303565,I303514);
nor I_17704 (I303355,I303582,I303480);
nor I_17705 (I303613,I303497,I303582);
nand I_17706 (I303358,I303548,I303613);
not I_17707 (I303644,I166264);
nor I_17708 (I303661,I303644,I166273);
nor I_17709 (I303678,I303661,I166267);
nor I_17710 (I303695,I303446,I303678);
DFFARX1 I_17711 (I303695,I2595,I303381,I303367,);
not I_17712 (I303726,I303661);
DFFARX1 I_17713 (I303726,I2595,I303381,I303370,);
and I_17714 (I303364,I303472,I303661);
nor I_17715 (I303771,I303644,I166288);
and I_17716 (I303788,I303771,I166267);
or I_17717 (I303805,I303788,I166285);
DFFARX1 I_17718 (I303805,I2595,I303381,I303831,);
nor I_17719 (I303839,I303831,I303565);
DFFARX1 I_17720 (I303839,I2595,I303381,I303352,);
nand I_17721 (I303870,I303831,I303472);
nand I_17722 (I303887,I303565,I303870);
nor I_17723 (I303361,I303887,I303531);
not I_17724 (I303942,I2602);
DFFARX1 I_17725 (I386038,I2595,I303942,I303968,);
DFFARX1 I_17726 (I303968,I2595,I303942,I303985,);
not I_17727 (I303934,I303985);
not I_17728 (I304007,I303968);
DFFARX1 I_17729 (I386032,I2595,I303942,I304033,);
nand I_17730 (I304041,I304033,I386023);
not I_17731 (I304058,I386023);
not I_17732 (I304075,I386050);
nand I_17733 (I304092,I386035,I386044);
and I_17734 (I304109,I386035,I386044);
not I_17735 (I304126,I386029);
nand I_17736 (I304143,I304126,I304075);
nor I_17737 (I303916,I304143,I304041);
nor I_17738 (I304174,I304058,I304143);
nand I_17739 (I303919,I304109,I304174);
not I_17740 (I304205,I386047);
nor I_17741 (I304222,I304205,I386035);
nor I_17742 (I304239,I304222,I386029);
nor I_17743 (I304256,I304007,I304239);
DFFARX1 I_17744 (I304256,I2595,I303942,I303928,);
not I_17745 (I304287,I304222);
DFFARX1 I_17746 (I304287,I2595,I303942,I303931,);
and I_17747 (I303925,I304033,I304222);
nor I_17748 (I304332,I304205,I386041);
and I_17749 (I304349,I304332,I386023);
or I_17750 (I304366,I304349,I386026);
DFFARX1 I_17751 (I304366,I2595,I303942,I304392,);
nor I_17752 (I304400,I304392,I304126);
DFFARX1 I_17753 (I304400,I2595,I303942,I303913,);
nand I_17754 (I304431,I304392,I304033);
nand I_17755 (I304448,I304126,I304431);
nor I_17756 (I303922,I304448,I304092);
not I_17757 (I304503,I2602);
DFFARX1 I_17758 (I389013,I2595,I304503,I304529,);
DFFARX1 I_17759 (I304529,I2595,I304503,I304546,);
not I_17760 (I304495,I304546);
not I_17761 (I304568,I304529);
DFFARX1 I_17762 (I389007,I2595,I304503,I304594,);
nand I_17763 (I304602,I304594,I388998);
not I_17764 (I304619,I388998);
not I_17765 (I304636,I389025);
nand I_17766 (I304653,I389010,I389019);
and I_17767 (I304670,I389010,I389019);
not I_17768 (I304687,I389004);
nand I_17769 (I304704,I304687,I304636);
nor I_17770 (I304477,I304704,I304602);
nor I_17771 (I304735,I304619,I304704);
nand I_17772 (I304480,I304670,I304735);
not I_17773 (I304766,I389022);
nor I_17774 (I304783,I304766,I389010);
nor I_17775 (I304800,I304783,I389004);
nor I_17776 (I304817,I304568,I304800);
DFFARX1 I_17777 (I304817,I2595,I304503,I304489,);
not I_17778 (I304848,I304783);
DFFARX1 I_17779 (I304848,I2595,I304503,I304492,);
and I_17780 (I304486,I304594,I304783);
nor I_17781 (I304893,I304766,I389016);
and I_17782 (I304910,I304893,I388998);
or I_17783 (I304927,I304910,I389001);
DFFARX1 I_17784 (I304927,I2595,I304503,I304953,);
nor I_17785 (I304961,I304953,I304687);
DFFARX1 I_17786 (I304961,I2595,I304503,I304474,);
nand I_17787 (I304992,I304953,I304594);
nand I_17788 (I305009,I304687,I304992);
nor I_17789 (I304483,I305009,I304653);
not I_17790 (I305064,I2602);
DFFARX1 I_17791 (I271885,I2595,I305064,I305090,);
DFFARX1 I_17792 (I305090,I2595,I305064,I305107,);
not I_17793 (I305056,I305107);
not I_17794 (I305129,I305090);
DFFARX1 I_17795 (I271912,I2595,I305064,I305155,);
nand I_17796 (I305163,I305155,I271903);
not I_17797 (I305180,I271903);
not I_17798 (I305197,I271885);
nand I_17799 (I305214,I271897,I271900);
and I_17800 (I305231,I271897,I271900);
not I_17801 (I305248,I271909);
nand I_17802 (I305265,I305248,I305197);
nor I_17803 (I305038,I305265,I305163);
nor I_17804 (I305296,I305180,I305265);
nand I_17805 (I305041,I305231,I305296);
not I_17806 (I305327,I271894);
nor I_17807 (I305344,I305327,I271897);
nor I_17808 (I305361,I305344,I271909);
nor I_17809 (I305378,I305129,I305361);
DFFARX1 I_17810 (I305378,I2595,I305064,I305050,);
not I_17811 (I305409,I305344);
DFFARX1 I_17812 (I305409,I2595,I305064,I305053,);
and I_17813 (I305047,I305155,I305344);
nor I_17814 (I305454,I305327,I271888);
and I_17815 (I305471,I305454,I271891);
or I_17816 (I305488,I305471,I271906);
DFFARX1 I_17817 (I305488,I2595,I305064,I305514,);
nor I_17818 (I305522,I305514,I305248);
DFFARX1 I_17819 (I305522,I2595,I305064,I305035,);
nand I_17820 (I305553,I305514,I305155);
nand I_17821 (I305570,I305248,I305553);
nor I_17822 (I305044,I305570,I305214);
not I_17823 (I305628,I2602);
DFFARX1 I_17824 (I269953,I2595,I305628,I305654,);
and I_17825 (I305662,I305654,I269947);
DFFARX1 I_17826 (I305662,I2595,I305628,I305611,);
DFFARX1 I_17827 (I269965,I2595,I305628,I305702,);
not I_17828 (I305710,I269956);
not I_17829 (I305727,I269968);
nand I_17830 (I305744,I305727,I305710);
nor I_17831 (I305599,I305702,I305744);
DFFARX1 I_17832 (I305744,I2595,I305628,I305784,);
not I_17833 (I305620,I305784);
not I_17834 (I305806,I269974);
nand I_17835 (I305823,I305727,I305806);
DFFARX1 I_17836 (I305823,I2595,I305628,I305849,);
not I_17837 (I305857,I305849);
not I_17838 (I305874,I269950);
nand I_17839 (I305891,I305874,I269971);
and I_17840 (I305908,I305710,I305891);
nor I_17841 (I305925,I305823,I305908);
DFFARX1 I_17842 (I305925,I2595,I305628,I305596,);
DFFARX1 I_17843 (I305908,I2595,I305628,I305617,);
nor I_17844 (I305970,I269950,I269962);
nor I_17845 (I305608,I305823,I305970);
or I_17846 (I306001,I269950,I269962);
nor I_17847 (I306018,I269947,I269959);
DFFARX1 I_17848 (I306018,I2595,I305628,I306044,);
not I_17849 (I306052,I306044);
nor I_17850 (I305614,I306052,I305857);
nand I_17851 (I306083,I306052,I305702);
not I_17852 (I306100,I269947);
nand I_17853 (I306117,I306100,I305806);
nand I_17854 (I306134,I306052,I306117);
nand I_17855 (I305605,I306134,I306083);
nand I_17856 (I305602,I306117,I306001);
not I_17857 (I306206,I2602);
DFFARX1 I_17858 (I189977,I2595,I306206,I306232,);
and I_17859 (I306240,I306232,I189965);
DFFARX1 I_17860 (I306240,I2595,I306206,I306189,);
DFFARX1 I_17861 (I189968,I2595,I306206,I306280,);
not I_17862 (I306288,I189962);
not I_17863 (I306305,I189986);
nand I_17864 (I306322,I306305,I306288);
nor I_17865 (I306177,I306280,I306322);
DFFARX1 I_17866 (I306322,I2595,I306206,I306362,);
not I_17867 (I306198,I306362);
not I_17868 (I306384,I189974);
nand I_17869 (I306401,I306305,I306384);
DFFARX1 I_17870 (I306401,I2595,I306206,I306427,);
not I_17871 (I306435,I306427);
not I_17872 (I306452,I189983);
nand I_17873 (I306469,I306452,I189980);
and I_17874 (I306486,I306288,I306469);
nor I_17875 (I306503,I306401,I306486);
DFFARX1 I_17876 (I306503,I2595,I306206,I306174,);
DFFARX1 I_17877 (I306486,I2595,I306206,I306195,);
nor I_17878 (I306548,I189983,I189971);
nor I_17879 (I306186,I306401,I306548);
or I_17880 (I306579,I189983,I189971);
nor I_17881 (I306596,I189962,I189965);
DFFARX1 I_17882 (I306596,I2595,I306206,I306622,);
not I_17883 (I306630,I306622);
nor I_17884 (I306192,I306630,I306435);
nand I_17885 (I306661,I306630,I306280);
not I_17886 (I306678,I189962);
nand I_17887 (I306695,I306678,I306384);
nand I_17888 (I306712,I306630,I306695);
nand I_17889 (I306183,I306712,I306661);
nand I_17890 (I306180,I306695,I306579);
not I_17891 (I306784,I2602);
DFFARX1 I_17892 (I262201,I2595,I306784,I306810,);
and I_17893 (I306818,I306810,I262195);
DFFARX1 I_17894 (I306818,I2595,I306784,I306767,);
DFFARX1 I_17895 (I262213,I2595,I306784,I306858,);
not I_17896 (I306866,I262204);
not I_17897 (I306883,I262216);
nand I_17898 (I306900,I306883,I306866);
nor I_17899 (I306755,I306858,I306900);
DFFARX1 I_17900 (I306900,I2595,I306784,I306940,);
not I_17901 (I306776,I306940);
not I_17902 (I306962,I262222);
nand I_17903 (I306979,I306883,I306962);
DFFARX1 I_17904 (I306979,I2595,I306784,I307005,);
not I_17905 (I307013,I307005);
not I_17906 (I307030,I262198);
nand I_17907 (I307047,I307030,I262219);
and I_17908 (I307064,I306866,I307047);
nor I_17909 (I307081,I306979,I307064);
DFFARX1 I_17910 (I307081,I2595,I306784,I306752,);
DFFARX1 I_17911 (I307064,I2595,I306784,I306773,);
nor I_17912 (I307126,I262198,I262210);
nor I_17913 (I306764,I306979,I307126);
or I_17914 (I307157,I262198,I262210);
nor I_17915 (I307174,I262195,I262207);
DFFARX1 I_17916 (I307174,I2595,I306784,I307200,);
not I_17917 (I307208,I307200);
nor I_17918 (I306770,I307208,I307013);
nand I_17919 (I307239,I307208,I306858);
not I_17920 (I307256,I262195);
nand I_17921 (I307273,I307256,I306962);
nand I_17922 (I307290,I307208,I307273);
nand I_17923 (I306761,I307290,I307239);
nand I_17924 (I306758,I307273,I307157);
not I_17925 (I307362,I2602);
DFFARX1 I_17926 (I136089,I2595,I307362,I307388,);
and I_17927 (I307396,I307388,I136104);
DFFARX1 I_17928 (I307396,I2595,I307362,I307345,);
DFFARX1 I_17929 (I136107,I2595,I307362,I307436,);
not I_17930 (I307444,I136101);
not I_17931 (I307461,I136116);
nand I_17932 (I307478,I307461,I307444);
nor I_17933 (I307333,I307436,I307478);
DFFARX1 I_17934 (I307478,I2595,I307362,I307518,);
not I_17935 (I307354,I307518);
not I_17936 (I307540,I136092);
nand I_17937 (I307557,I307461,I307540);
DFFARX1 I_17938 (I307557,I2595,I307362,I307583,);
not I_17939 (I307591,I307583);
not I_17940 (I307608,I136095);
nand I_17941 (I307625,I307608,I136089);
and I_17942 (I307642,I307444,I307625);
nor I_17943 (I307659,I307557,I307642);
DFFARX1 I_17944 (I307659,I2595,I307362,I307330,);
DFFARX1 I_17945 (I307642,I2595,I307362,I307351,);
nor I_17946 (I307704,I136095,I136098);
nor I_17947 (I307342,I307557,I307704);
or I_17948 (I307735,I136095,I136098);
nor I_17949 (I307752,I136113,I136110);
DFFARX1 I_17950 (I307752,I2595,I307362,I307778,);
not I_17951 (I307786,I307778);
nor I_17952 (I307348,I307786,I307591);
nand I_17953 (I307817,I307786,I307436);
not I_17954 (I307834,I136113);
nand I_17955 (I307851,I307834,I307540);
nand I_17956 (I307868,I307786,I307851);
nand I_17957 (I307339,I307868,I307817);
nand I_17958 (I307336,I307851,I307735);
not I_17959 (I307940,I2602);
DFFARX1 I_17960 (I286103,I2595,I307940,I307966,);
and I_17961 (I307974,I307966,I286097);
DFFARX1 I_17962 (I307974,I2595,I307940,I307923,);
DFFARX1 I_17963 (I286115,I2595,I307940,I308014,);
not I_17964 (I308022,I286106);
not I_17965 (I308039,I286118);
nand I_17966 (I308056,I308039,I308022);
nor I_17967 (I307911,I308014,I308056);
DFFARX1 I_17968 (I308056,I2595,I307940,I308096,);
not I_17969 (I307932,I308096);
not I_17970 (I308118,I286124);
nand I_17971 (I308135,I308039,I308118);
DFFARX1 I_17972 (I308135,I2595,I307940,I308161,);
not I_17973 (I308169,I308161);
not I_17974 (I308186,I286100);
nand I_17975 (I308203,I308186,I286121);
and I_17976 (I308220,I308022,I308203);
nor I_17977 (I308237,I308135,I308220);
DFFARX1 I_17978 (I308237,I2595,I307940,I307908,);
DFFARX1 I_17979 (I308220,I2595,I307940,I307929,);
nor I_17980 (I308282,I286100,I286112);
nor I_17981 (I307920,I308135,I308282);
or I_17982 (I308313,I286100,I286112);
nor I_17983 (I308330,I286097,I286109);
DFFARX1 I_17984 (I308330,I2595,I307940,I308356,);
not I_17985 (I308364,I308356);
nor I_17986 (I307926,I308364,I308169);
nand I_17987 (I308395,I308364,I308014);
not I_17988 (I308412,I286097);
nand I_17989 (I308429,I308412,I308118);
nand I_17990 (I308446,I308364,I308429);
nand I_17991 (I307917,I308446,I308395);
nand I_17992 (I307914,I308429,I308313);
not I_17993 (I308518,I2602);
DFFARX1 I_17994 (I380695,I2595,I308518,I308544,);
and I_17995 (I308552,I308544,I380677);
DFFARX1 I_17996 (I308552,I2595,I308518,I308501,);
DFFARX1 I_17997 (I380668,I2595,I308518,I308592,);
not I_17998 (I308600,I380683);
not I_17999 (I308617,I380671);
nand I_18000 (I308634,I308617,I308600);
nor I_18001 (I308489,I308592,I308634);
DFFARX1 I_18002 (I308634,I2595,I308518,I308674,);
not I_18003 (I308510,I308674);
not I_18004 (I308696,I380680);
nand I_18005 (I308713,I308617,I308696);
DFFARX1 I_18006 (I308713,I2595,I308518,I308739,);
not I_18007 (I308747,I308739);
not I_18008 (I308764,I380689);
nand I_18009 (I308781,I308764,I380668);
and I_18010 (I308798,I308600,I308781);
nor I_18011 (I308815,I308713,I308798);
DFFARX1 I_18012 (I308815,I2595,I308518,I308486,);
DFFARX1 I_18013 (I308798,I2595,I308518,I308507,);
nor I_18014 (I308860,I380689,I380692);
nor I_18015 (I308498,I308713,I308860);
or I_18016 (I308891,I380689,I380692);
nor I_18017 (I308908,I380686,I380674);
DFFARX1 I_18018 (I308908,I2595,I308518,I308934,);
not I_18019 (I308942,I308934);
nor I_18020 (I308504,I308942,I308747);
nand I_18021 (I308973,I308942,I308592);
not I_18022 (I308990,I380686);
nand I_18023 (I309007,I308990,I308696);
nand I_18024 (I309024,I308942,I309007);
nand I_18025 (I308495,I309024,I308973);
nand I_18026 (I308492,I309007,I308891);
not I_18027 (I309096,I2602);
DFFARX1 I_18028 (I3215,I2595,I309096,I309122,);
and I_18029 (I309130,I309122,I3221);
DFFARX1 I_18030 (I309130,I2595,I309096,I309079,);
DFFARX1 I_18031 (I3200,I2595,I309096,I309170,);
not I_18032 (I309178,I3206);
not I_18033 (I309195,I3212);
nand I_18034 (I309212,I309195,I309178);
nor I_18035 (I309067,I309170,I309212);
DFFARX1 I_18036 (I309212,I2595,I309096,I309252,);
not I_18037 (I309088,I309252);
not I_18038 (I309274,I3203);
nand I_18039 (I309291,I309195,I309274);
DFFARX1 I_18040 (I309291,I2595,I309096,I309317,);
not I_18041 (I309325,I309317);
not I_18042 (I309342,I3218);
nand I_18043 (I309359,I309342,I3203);
and I_18044 (I309376,I309178,I309359);
nor I_18045 (I309393,I309291,I309376);
DFFARX1 I_18046 (I309393,I2595,I309096,I309064,);
DFFARX1 I_18047 (I309376,I2595,I309096,I309085,);
nor I_18048 (I309438,I3218,I3206);
nor I_18049 (I309076,I309291,I309438);
or I_18050 (I309469,I3218,I3206);
nor I_18051 (I309486,I3209,I3200);
DFFARX1 I_18052 (I309486,I2595,I309096,I309512,);
not I_18053 (I309520,I309512);
nor I_18054 (I309082,I309520,I309325);
nand I_18055 (I309551,I309520,I309170);
not I_18056 (I309568,I3209);
nand I_18057 (I309585,I309568,I309274);
nand I_18058 (I309602,I309520,I309585);
nand I_18059 (I309073,I309602,I309551);
nand I_18060 (I309070,I309585,I309469);
not I_18061 (I309674,I2602);
DFFARX1 I_18062 (I156453,I2595,I309674,I309700,);
and I_18063 (I309708,I309700,I156441);
DFFARX1 I_18064 (I309708,I2595,I309674,I309657,);
DFFARX1 I_18065 (I156456,I2595,I309674,I309748,);
not I_18066 (I309756,I156447);
not I_18067 (I309773,I156438);
nand I_18068 (I309790,I309773,I309756);
nor I_18069 (I309645,I309748,I309790);
DFFARX1 I_18070 (I309790,I2595,I309674,I309830,);
not I_18071 (I309666,I309830);
not I_18072 (I309852,I156444);
nand I_18073 (I309869,I309773,I309852);
DFFARX1 I_18074 (I309869,I2595,I309674,I309895,);
not I_18075 (I309903,I309895);
not I_18076 (I309920,I156459);
nand I_18077 (I309937,I309920,I156462);
and I_18078 (I309954,I309756,I309937);
nor I_18079 (I309971,I309869,I309954);
DFFARX1 I_18080 (I309971,I2595,I309674,I309642,);
DFFARX1 I_18081 (I309954,I2595,I309674,I309663,);
nor I_18082 (I310016,I156459,I156438);
nor I_18083 (I309654,I309869,I310016);
or I_18084 (I310047,I156459,I156438);
nor I_18085 (I310064,I156450,I156441);
DFFARX1 I_18086 (I310064,I2595,I309674,I310090,);
not I_18087 (I310098,I310090);
nor I_18088 (I309660,I310098,I309903);
nand I_18089 (I310129,I310098,I309748);
not I_18090 (I310146,I156450);
nand I_18091 (I310163,I310146,I309852);
nand I_18092 (I310180,I310098,I310163);
nand I_18093 (I309651,I310180,I310129);
nand I_18094 (I309648,I310163,I310047);
not I_18095 (I310252,I2602);
DFFARX1 I_18096 (I292135,I2595,I310252,I310278,);
and I_18097 (I310286,I310278,I292132);
DFFARX1 I_18098 (I310286,I2595,I310252,I310235,);
DFFARX1 I_18099 (I292138,I2595,I310252,I310326,);
not I_18100 (I310334,I292141);
not I_18101 (I310351,I292135);
nand I_18102 (I310368,I310351,I310334);
nor I_18103 (I310223,I310326,I310368);
DFFARX1 I_18104 (I310368,I2595,I310252,I310408,);
not I_18105 (I310244,I310408);
not I_18106 (I310430,I292150);
nand I_18107 (I310447,I310351,I310430);
DFFARX1 I_18108 (I310447,I2595,I310252,I310473,);
not I_18109 (I310481,I310473);
not I_18110 (I310498,I292147);
nand I_18111 (I310515,I310498,I292153);
and I_18112 (I310532,I310334,I310515);
nor I_18113 (I310549,I310447,I310532);
DFFARX1 I_18114 (I310549,I2595,I310252,I310220,);
DFFARX1 I_18115 (I310532,I2595,I310252,I310241,);
nor I_18116 (I310594,I292147,I292132);
nor I_18117 (I310232,I310447,I310594);
or I_18118 (I310625,I292147,I292132);
nor I_18119 (I310642,I292144,I292138);
DFFARX1 I_18120 (I310642,I2595,I310252,I310668,);
not I_18121 (I310676,I310668);
nor I_18122 (I310238,I310676,I310481);
nand I_18123 (I310707,I310676,I310326);
not I_18124 (I310724,I292144);
nand I_18125 (I310741,I310724,I310430);
nand I_18126 (I310758,I310676,I310741);
nand I_18127 (I310229,I310758,I310707);
nand I_18128 (I310226,I310741,I310625);
not I_18129 (I310830,I2602);
DFFARX1 I_18130 (I153483,I2595,I310830,I310856,);
and I_18131 (I310864,I310856,I153498);
DFFARX1 I_18132 (I310864,I2595,I310830,I310813,);
DFFARX1 I_18133 (I153489,I2595,I310830,I310904,);
not I_18134 (I310912,I153483);
not I_18135 (I310929,I153501);
nand I_18136 (I310946,I310929,I310912);
nor I_18137 (I310801,I310904,I310946);
DFFARX1 I_18138 (I310946,I2595,I310830,I310986,);
not I_18139 (I310822,I310986);
not I_18140 (I311008,I153492);
nand I_18141 (I311025,I310929,I311008);
DFFARX1 I_18142 (I311025,I2595,I310830,I311051,);
not I_18143 (I311059,I311051);
not I_18144 (I311076,I153504);
nand I_18145 (I311093,I311076,I153480);
and I_18146 (I311110,I310912,I311093);
nor I_18147 (I311127,I311025,I311110);
DFFARX1 I_18148 (I311127,I2595,I310830,I310798,);
DFFARX1 I_18149 (I311110,I2595,I310830,I310819,);
nor I_18150 (I311172,I153504,I153480);
nor I_18151 (I310810,I311025,I311172);
or I_18152 (I311203,I153504,I153480);
nor I_18153 (I311220,I153486,I153495);
DFFARX1 I_18154 (I311220,I2595,I310830,I311246,);
not I_18155 (I311254,I311246);
nor I_18156 (I310816,I311254,I311059);
nand I_18157 (I311285,I311254,I310904);
not I_18158 (I311302,I153486);
nand I_18159 (I311319,I311302,I311008);
nand I_18160 (I311336,I311254,I311319);
nand I_18161 (I310807,I311336,I311285);
nand I_18162 (I310804,I311319,I311203);
not I_18163 (I311408,I2602);
DFFARX1 I_18164 (I96982,I2595,I311408,I311434,);
and I_18165 (I311442,I311434,I96967);
DFFARX1 I_18166 (I311442,I2595,I311408,I311391,);
DFFARX1 I_18167 (I96973,I2595,I311408,I311482,);
not I_18168 (I311490,I96955);
not I_18169 (I311507,I96976);
nand I_18170 (I311524,I311507,I311490);
nor I_18171 (I311379,I311482,I311524);
DFFARX1 I_18172 (I311524,I2595,I311408,I311564,);
not I_18173 (I311400,I311564);
not I_18174 (I311586,I96979);
nand I_18175 (I311603,I311507,I311586);
DFFARX1 I_18176 (I311603,I2595,I311408,I311629,);
not I_18177 (I311637,I311629);
not I_18178 (I311654,I96970);
nand I_18179 (I311671,I311654,I96958);
and I_18180 (I311688,I311490,I311671);
nor I_18181 (I311705,I311603,I311688);
DFFARX1 I_18182 (I311705,I2595,I311408,I311376,);
DFFARX1 I_18183 (I311688,I2595,I311408,I311397,);
nor I_18184 (I311750,I96970,I96964);
nor I_18185 (I311388,I311603,I311750);
or I_18186 (I311781,I96970,I96964);
nor I_18187 (I311798,I96961,I96955);
DFFARX1 I_18188 (I311798,I2595,I311408,I311824,);
not I_18189 (I311832,I311824);
nor I_18190 (I311394,I311832,I311637);
nand I_18191 (I311863,I311832,I311482);
not I_18192 (I311880,I96961);
nand I_18193 (I311897,I311880,I311586);
nand I_18194 (I311914,I311832,I311897);
nand I_18195 (I311385,I311914,I311863);
nand I_18196 (I311382,I311897,I311781);
not I_18197 (I311986,I2602);
DFFARX1 I_18198 (I243549,I2595,I311986,I312012,);
and I_18199 (I312020,I312012,I243555);
DFFARX1 I_18200 (I312020,I2595,I311986,I311969,);
DFFARX1 I_18201 (I243561,I2595,I311986,I312060,);
not I_18202 (I312068,I243546);
not I_18203 (I312085,I243546);
nand I_18204 (I312102,I312085,I312068);
nor I_18205 (I311957,I312060,I312102);
DFFARX1 I_18206 (I312102,I2595,I311986,I312142,);
not I_18207 (I311978,I312142);
not I_18208 (I312164,I243564);
nand I_18209 (I312181,I312085,I312164);
DFFARX1 I_18210 (I312181,I2595,I311986,I312207,);
not I_18211 (I312215,I312207);
not I_18212 (I312232,I243558);
nand I_18213 (I312249,I312232,I243549);
and I_18214 (I312266,I312068,I312249);
nor I_18215 (I312283,I312181,I312266);
DFFARX1 I_18216 (I312283,I2595,I311986,I311954,);
DFFARX1 I_18217 (I312266,I2595,I311986,I311975,);
nor I_18218 (I312328,I243558,I243567);
nor I_18219 (I311966,I312181,I312328);
or I_18220 (I312359,I243558,I243567);
nor I_18221 (I312376,I243552,I243552);
DFFARX1 I_18222 (I312376,I2595,I311986,I312402,);
not I_18223 (I312410,I312402);
nor I_18224 (I311972,I312410,I312215);
nand I_18225 (I312441,I312410,I312060);
not I_18226 (I312458,I243552);
nand I_18227 (I312475,I312458,I312164);
nand I_18228 (I312492,I312410,I312475);
nand I_18229 (I311963,I312492,I312441);
nand I_18230 (I311960,I312475,I312359);
not I_18231 (I312564,I2602);
DFFARX1 I_18232 (I16069,I2595,I312564,I312590,);
and I_18233 (I312598,I312590,I16072);
DFFARX1 I_18234 (I312598,I2595,I312564,I312547,);
DFFARX1 I_18235 (I16072,I2595,I312564,I312638,);
not I_18236 (I312646,I16075);
not I_18237 (I312663,I16090);
nand I_18238 (I312680,I312663,I312646);
nor I_18239 (I312535,I312638,I312680);
DFFARX1 I_18240 (I312680,I2595,I312564,I312720,);
not I_18241 (I312556,I312720);
not I_18242 (I312742,I16084);
nand I_18243 (I312759,I312663,I312742);
DFFARX1 I_18244 (I312759,I2595,I312564,I312785,);
not I_18245 (I312793,I312785);
not I_18246 (I312810,I16087);
nand I_18247 (I312827,I312810,I16069);
and I_18248 (I312844,I312646,I312827);
nor I_18249 (I312861,I312759,I312844);
DFFARX1 I_18250 (I312861,I2595,I312564,I312532,);
DFFARX1 I_18251 (I312844,I2595,I312564,I312553,);
nor I_18252 (I312906,I16087,I16081);
nor I_18253 (I312544,I312759,I312906);
or I_18254 (I312937,I16087,I16081);
nor I_18255 (I312954,I16078,I16093);
DFFARX1 I_18256 (I312954,I2595,I312564,I312980,);
not I_18257 (I312988,I312980);
nor I_18258 (I312550,I312988,I312793);
nand I_18259 (I313019,I312988,I312638);
not I_18260 (I313036,I16078);
nand I_18261 (I313053,I313036,I312742);
nand I_18262 (I313070,I312988,I313053);
nand I_18263 (I312541,I313070,I313019);
nand I_18264 (I312538,I313053,I312937);
not I_18265 (I313142,I2602);
DFFARX1 I_18266 (I190555,I2595,I313142,I313168,);
and I_18267 (I313176,I313168,I190543);
DFFARX1 I_18268 (I313176,I2595,I313142,I313125,);
DFFARX1 I_18269 (I190546,I2595,I313142,I313216,);
not I_18270 (I313224,I190540);
not I_18271 (I313241,I190564);
nand I_18272 (I313258,I313241,I313224);
nor I_18273 (I313113,I313216,I313258);
DFFARX1 I_18274 (I313258,I2595,I313142,I313298,);
not I_18275 (I313134,I313298);
not I_18276 (I313320,I190552);
nand I_18277 (I313337,I313241,I313320);
DFFARX1 I_18278 (I313337,I2595,I313142,I313363,);
not I_18279 (I313371,I313363);
not I_18280 (I313388,I190561);
nand I_18281 (I313405,I313388,I190558);
and I_18282 (I313422,I313224,I313405);
nor I_18283 (I313439,I313337,I313422);
DFFARX1 I_18284 (I313439,I2595,I313142,I313110,);
DFFARX1 I_18285 (I313422,I2595,I313142,I313131,);
nor I_18286 (I313484,I190561,I190549);
nor I_18287 (I313122,I313337,I313484);
or I_18288 (I313515,I190561,I190549);
nor I_18289 (I313532,I190540,I190543);
DFFARX1 I_18290 (I313532,I2595,I313142,I313558,);
not I_18291 (I313566,I313558);
nor I_18292 (I313128,I313566,I313371);
nand I_18293 (I313597,I313566,I313216);
not I_18294 (I313614,I190540);
nand I_18295 (I313631,I313614,I313320);
nand I_18296 (I313648,I313566,I313631);
nand I_18297 (I313119,I313648,I313597);
nand I_18298 (I313116,I313631,I313515);
not I_18299 (I313720,I2602);
DFFARX1 I_18300 (I231428,I2595,I313720,I313746,);
and I_18301 (I313754,I313746,I231434);
DFFARX1 I_18302 (I313754,I2595,I313720,I313703,);
DFFARX1 I_18303 (I231440,I2595,I313720,I313794,);
not I_18304 (I313802,I231425);
not I_18305 (I313819,I231425);
nand I_18306 (I313836,I313819,I313802);
nor I_18307 (I313691,I313794,I313836);
DFFARX1 I_18308 (I313836,I2595,I313720,I313876,);
not I_18309 (I313712,I313876);
not I_18310 (I313898,I231443);
nand I_18311 (I313915,I313819,I313898);
DFFARX1 I_18312 (I313915,I2595,I313720,I313941,);
not I_18313 (I313949,I313941);
not I_18314 (I313966,I231437);
nand I_18315 (I313983,I313966,I231428);
and I_18316 (I314000,I313802,I313983);
nor I_18317 (I314017,I313915,I314000);
DFFARX1 I_18318 (I314017,I2595,I313720,I313688,);
DFFARX1 I_18319 (I314000,I2595,I313720,I313709,);
nor I_18320 (I314062,I231437,I231446);
nor I_18321 (I313700,I313915,I314062);
or I_18322 (I314093,I231437,I231446);
nor I_18323 (I314110,I231431,I231431);
DFFARX1 I_18324 (I314110,I2595,I313720,I314136,);
not I_18325 (I314144,I314136);
nor I_18326 (I313706,I314144,I313949);
nand I_18327 (I314175,I314144,I313794);
not I_18328 (I314192,I231431);
nand I_18329 (I314209,I314192,I313898);
nand I_18330 (I314226,I314144,I314209);
nand I_18331 (I313697,I314226,I314175);
nand I_18332 (I313694,I314209,I314093);
not I_18333 (I314298,I2602);
DFFARX1 I_18334 (I92766,I2595,I314298,I314324,);
and I_18335 (I314332,I314324,I92751);
DFFARX1 I_18336 (I314332,I2595,I314298,I314281,);
DFFARX1 I_18337 (I92757,I2595,I314298,I314372,);
not I_18338 (I314380,I92739);
not I_18339 (I314397,I92760);
nand I_18340 (I314414,I314397,I314380);
nor I_18341 (I314269,I314372,I314414);
DFFARX1 I_18342 (I314414,I2595,I314298,I314454,);
not I_18343 (I314290,I314454);
not I_18344 (I314476,I92763);
nand I_18345 (I314493,I314397,I314476);
DFFARX1 I_18346 (I314493,I2595,I314298,I314519,);
not I_18347 (I314527,I314519);
not I_18348 (I314544,I92754);
nand I_18349 (I314561,I314544,I92742);
and I_18350 (I314578,I314380,I314561);
nor I_18351 (I314595,I314493,I314578);
DFFARX1 I_18352 (I314595,I2595,I314298,I314266,);
DFFARX1 I_18353 (I314578,I2595,I314298,I314287,);
nor I_18354 (I314640,I92754,I92748);
nor I_18355 (I314278,I314493,I314640);
or I_18356 (I314671,I92754,I92748);
nor I_18357 (I314688,I92745,I92739);
DFFARX1 I_18358 (I314688,I2595,I314298,I314714,);
not I_18359 (I314722,I314714);
nor I_18360 (I314284,I314722,I314527);
nand I_18361 (I314753,I314722,I314372);
not I_18362 (I314770,I92745);
nand I_18363 (I314787,I314770,I314476);
nand I_18364 (I314804,I314722,I314787);
nand I_18365 (I314275,I314804,I314753);
nand I_18366 (I314272,I314787,I314671);
not I_18367 (I314876,I2602);
DFFARX1 I_18368 (I301672,I2595,I314876,I314902,);
and I_18369 (I314910,I314902,I301669);
DFFARX1 I_18370 (I314910,I2595,I314876,I314859,);
DFFARX1 I_18371 (I301675,I2595,I314876,I314950,);
not I_18372 (I314958,I301678);
not I_18373 (I314975,I301672);
nand I_18374 (I314992,I314975,I314958);
nor I_18375 (I314847,I314950,I314992);
DFFARX1 I_18376 (I314992,I2595,I314876,I315032,);
not I_18377 (I314868,I315032);
not I_18378 (I315054,I301687);
nand I_18379 (I315071,I314975,I315054);
DFFARX1 I_18380 (I315071,I2595,I314876,I315097,);
not I_18381 (I315105,I315097);
not I_18382 (I315122,I301684);
nand I_18383 (I315139,I315122,I301690);
and I_18384 (I315156,I314958,I315139);
nor I_18385 (I315173,I315071,I315156);
DFFARX1 I_18386 (I315173,I2595,I314876,I314844,);
DFFARX1 I_18387 (I315156,I2595,I314876,I314865,);
nor I_18388 (I315218,I301684,I301669);
nor I_18389 (I314856,I315071,I315218);
or I_18390 (I315249,I301684,I301669);
nor I_18391 (I315266,I301681,I301675);
DFFARX1 I_18392 (I315266,I2595,I314876,I315292,);
not I_18393 (I315300,I315292);
nor I_18394 (I314862,I315300,I315105);
nand I_18395 (I315331,I315300,I314950);
not I_18396 (I315348,I301681);
nand I_18397 (I315365,I315348,I315054);
nand I_18398 (I315382,I315300,I315365);
nand I_18399 (I314853,I315382,I315331);
nand I_18400 (I314850,I315365,I315249);
not I_18401 (I315454,I2602);
DFFARX1 I_18402 (I213675,I2595,I315454,I315480,);
and I_18403 (I315488,I315480,I213663);
DFFARX1 I_18404 (I315488,I2595,I315454,I315437,);
DFFARX1 I_18405 (I213666,I2595,I315454,I315528,);
not I_18406 (I315536,I213660);
not I_18407 (I315553,I213684);
nand I_18408 (I315570,I315553,I315536);
nor I_18409 (I315425,I315528,I315570);
DFFARX1 I_18410 (I315570,I2595,I315454,I315610,);
not I_18411 (I315446,I315610);
not I_18412 (I315632,I213672);
nand I_18413 (I315649,I315553,I315632);
DFFARX1 I_18414 (I315649,I2595,I315454,I315675,);
not I_18415 (I315683,I315675);
not I_18416 (I315700,I213681);
nand I_18417 (I315717,I315700,I213678);
and I_18418 (I315734,I315536,I315717);
nor I_18419 (I315751,I315649,I315734);
DFFARX1 I_18420 (I315751,I2595,I315454,I315422,);
DFFARX1 I_18421 (I315734,I2595,I315454,I315443,);
nor I_18422 (I315796,I213681,I213669);
nor I_18423 (I315434,I315649,I315796);
or I_18424 (I315827,I213681,I213669);
nor I_18425 (I315844,I213660,I213663);
DFFARX1 I_18426 (I315844,I2595,I315454,I315870,);
not I_18427 (I315878,I315870);
nor I_18428 (I315440,I315878,I315683);
nand I_18429 (I315909,I315878,I315528);
not I_18430 (I315926,I213660);
nand I_18431 (I315943,I315926,I315632);
nand I_18432 (I315960,I315878,I315943);
nand I_18433 (I315431,I315960,I315909);
nand I_18434 (I315428,I315943,I315827);
not I_18435 (I316032,I2602);
DFFARX1 I_18436 (I72883,I2595,I316032,I316058,);
and I_18437 (I316066,I316058,I72886);
DFFARX1 I_18438 (I316066,I2595,I316032,I316015,);
DFFARX1 I_18439 (I72886,I2595,I316032,I316106,);
not I_18440 (I316114,I72901);
not I_18441 (I316131,I72907);
nand I_18442 (I316148,I316131,I316114);
nor I_18443 (I316003,I316106,I316148);
DFFARX1 I_18444 (I316148,I2595,I316032,I316188,);
not I_18445 (I316024,I316188);
not I_18446 (I316210,I72895);
nand I_18447 (I316227,I316131,I316210);
DFFARX1 I_18448 (I316227,I2595,I316032,I316253,);
not I_18449 (I316261,I316253);
not I_18450 (I316278,I72892);
nand I_18451 (I316295,I316278,I72889);
and I_18452 (I316312,I316114,I316295);
nor I_18453 (I316329,I316227,I316312);
DFFARX1 I_18454 (I316329,I2595,I316032,I316000,);
DFFARX1 I_18455 (I316312,I2595,I316032,I316021,);
nor I_18456 (I316374,I72892,I72883);
nor I_18457 (I316012,I316227,I316374);
or I_18458 (I316405,I72892,I72883);
nor I_18459 (I316422,I72898,I72904);
DFFARX1 I_18460 (I316422,I2595,I316032,I316448,);
not I_18461 (I316456,I316448);
nor I_18462 (I316018,I316456,I316261);
nand I_18463 (I316487,I316456,I316106);
not I_18464 (I316504,I72898);
nand I_18465 (I316521,I316504,I316210);
nand I_18466 (I316538,I316456,I316521);
nand I_18467 (I316009,I316538,I316487);
nand I_18468 (I316006,I316521,I316405);
not I_18469 (I316610,I2602);
DFFARX1 I_18470 (I375340,I2595,I316610,I316636,);
and I_18471 (I316644,I316636,I375322);
DFFARX1 I_18472 (I316644,I2595,I316610,I316593,);
DFFARX1 I_18473 (I375313,I2595,I316610,I316684,);
not I_18474 (I316692,I375328);
not I_18475 (I316709,I375316);
nand I_18476 (I316726,I316709,I316692);
nor I_18477 (I316581,I316684,I316726);
DFFARX1 I_18478 (I316726,I2595,I316610,I316766,);
not I_18479 (I316602,I316766);
not I_18480 (I316788,I375325);
nand I_18481 (I316805,I316709,I316788);
DFFARX1 I_18482 (I316805,I2595,I316610,I316831,);
not I_18483 (I316839,I316831);
not I_18484 (I316856,I375334);
nand I_18485 (I316873,I316856,I375313);
and I_18486 (I316890,I316692,I316873);
nor I_18487 (I316907,I316805,I316890);
DFFARX1 I_18488 (I316907,I2595,I316610,I316578,);
DFFARX1 I_18489 (I316890,I2595,I316610,I316599,);
nor I_18490 (I316952,I375334,I375337);
nor I_18491 (I316590,I316805,I316952);
or I_18492 (I316983,I375334,I375337);
nor I_18493 (I317000,I375331,I375319);
DFFARX1 I_18494 (I317000,I2595,I316610,I317026,);
not I_18495 (I317034,I317026);
nor I_18496 (I316596,I317034,I316839);
nand I_18497 (I317065,I317034,I316684);
not I_18498 (I317082,I375331);
nand I_18499 (I317099,I317082,I316788);
nand I_18500 (I317116,I317034,I317099);
nand I_18501 (I316587,I317116,I317065);
nand I_18502 (I316584,I317099,I316983);
not I_18503 (I317188,I2602);
DFFARX1 I_18504 (I147533,I2595,I317188,I317214,);
and I_18505 (I317222,I317214,I147548);
DFFARX1 I_18506 (I317222,I2595,I317188,I317171,);
DFFARX1 I_18507 (I147539,I2595,I317188,I317262,);
not I_18508 (I317270,I147533);
not I_18509 (I317287,I147551);
nand I_18510 (I317304,I317287,I317270);
nor I_18511 (I317159,I317262,I317304);
DFFARX1 I_18512 (I317304,I2595,I317188,I317344,);
not I_18513 (I317180,I317344);
not I_18514 (I317366,I147542);
nand I_18515 (I317383,I317287,I317366);
DFFARX1 I_18516 (I317383,I2595,I317188,I317409,);
not I_18517 (I317417,I317409);
not I_18518 (I317434,I147554);
nand I_18519 (I317451,I317434,I147530);
and I_18520 (I317468,I317270,I317451);
nor I_18521 (I317485,I317383,I317468);
DFFARX1 I_18522 (I317485,I2595,I317188,I317156,);
DFFARX1 I_18523 (I317468,I2595,I317188,I317177,);
nor I_18524 (I317530,I147554,I147530);
nor I_18525 (I317168,I317383,I317530);
or I_18526 (I317561,I147554,I147530);
nor I_18527 (I317578,I147536,I147545);
DFFARX1 I_18528 (I317578,I2595,I317188,I317604,);
not I_18529 (I317612,I317604);
nor I_18530 (I317174,I317612,I317417);
nand I_18531 (I317643,I317612,I317262);
not I_18532 (I317660,I147536);
nand I_18533 (I317677,I317660,I317366);
nand I_18534 (I317694,I317612,I317677);
nand I_18535 (I317165,I317694,I317643);
nand I_18536 (I317162,I317677,I317561);
not I_18537 (I317766,I2602);
DFFARX1 I_18538 (I143368,I2595,I317766,I317792,);
and I_18539 (I317800,I317792,I143383);
DFFARX1 I_18540 (I317800,I2595,I317766,I317749,);
DFFARX1 I_18541 (I143374,I2595,I317766,I317840,);
not I_18542 (I317848,I143368);
not I_18543 (I317865,I143386);
nand I_18544 (I317882,I317865,I317848);
nor I_18545 (I317737,I317840,I317882);
DFFARX1 I_18546 (I317882,I2595,I317766,I317922,);
not I_18547 (I317758,I317922);
not I_18548 (I317944,I143377);
nand I_18549 (I317961,I317865,I317944);
DFFARX1 I_18550 (I317961,I2595,I317766,I317987,);
not I_18551 (I317995,I317987);
not I_18552 (I318012,I143389);
nand I_18553 (I318029,I318012,I143365);
and I_18554 (I318046,I317848,I318029);
nor I_18555 (I318063,I317961,I318046);
DFFARX1 I_18556 (I318063,I2595,I317766,I317734,);
DFFARX1 I_18557 (I318046,I2595,I317766,I317755,);
nor I_18558 (I318108,I143389,I143365);
nor I_18559 (I317746,I317961,I318108);
or I_18560 (I318139,I143389,I143365);
nor I_18561 (I318156,I143371,I143380);
DFFARX1 I_18562 (I318156,I2595,I317766,I318182,);
not I_18563 (I318190,I318182);
nor I_18564 (I317752,I318190,I317995);
nand I_18565 (I318221,I318190,I317840);
not I_18566 (I318238,I143371);
nand I_18567 (I318255,I318238,I317944);
nand I_18568 (I318272,I318190,I318255);
nand I_18569 (I317743,I318272,I318221);
nand I_18570 (I317740,I318255,I318139);
not I_18571 (I318344,I2602);
DFFARX1 I_18572 (I145153,I2595,I318344,I318370,);
and I_18573 (I318378,I318370,I145168);
DFFARX1 I_18574 (I318378,I2595,I318344,I318327,);
DFFARX1 I_18575 (I145159,I2595,I318344,I318418,);
not I_18576 (I318426,I145153);
not I_18577 (I318443,I145171);
nand I_18578 (I318460,I318443,I318426);
nor I_18579 (I318315,I318418,I318460);
DFFARX1 I_18580 (I318460,I2595,I318344,I318500,);
not I_18581 (I318336,I318500);
not I_18582 (I318522,I145162);
nand I_18583 (I318539,I318443,I318522);
DFFARX1 I_18584 (I318539,I2595,I318344,I318565,);
not I_18585 (I318573,I318565);
not I_18586 (I318590,I145174);
nand I_18587 (I318607,I318590,I145150);
and I_18588 (I318624,I318426,I318607);
nor I_18589 (I318641,I318539,I318624);
DFFARX1 I_18590 (I318641,I2595,I318344,I318312,);
DFFARX1 I_18591 (I318624,I2595,I318344,I318333,);
nor I_18592 (I318686,I145174,I145150);
nor I_18593 (I318324,I318539,I318686);
or I_18594 (I318717,I145174,I145150);
nor I_18595 (I318734,I145156,I145165);
DFFARX1 I_18596 (I318734,I2595,I318344,I318760,);
not I_18597 (I318768,I318760);
nor I_18598 (I318330,I318768,I318573);
nand I_18599 (I318799,I318768,I318418);
not I_18600 (I318816,I145156);
nand I_18601 (I318833,I318816,I318522);
nand I_18602 (I318850,I318768,I318833);
nand I_18603 (I318321,I318850,I318799);
nand I_18604 (I318318,I318833,I318717);
not I_18605 (I318922,I2602);
DFFARX1 I_18606 (I184197,I2595,I318922,I318948,);
and I_18607 (I318956,I318948,I184185);
DFFARX1 I_18608 (I318956,I2595,I318922,I318905,);
DFFARX1 I_18609 (I184188,I2595,I318922,I318996,);
not I_18610 (I319004,I184182);
not I_18611 (I319021,I184206);
nand I_18612 (I319038,I319021,I319004);
nor I_18613 (I318893,I318996,I319038);
DFFARX1 I_18614 (I319038,I2595,I318922,I319078,);
not I_18615 (I318914,I319078);
not I_18616 (I319100,I184194);
nand I_18617 (I319117,I319021,I319100);
DFFARX1 I_18618 (I319117,I2595,I318922,I319143,);
not I_18619 (I319151,I319143);
not I_18620 (I319168,I184203);
nand I_18621 (I319185,I319168,I184200);
and I_18622 (I319202,I319004,I319185);
nor I_18623 (I319219,I319117,I319202);
DFFARX1 I_18624 (I319219,I2595,I318922,I318890,);
DFFARX1 I_18625 (I319202,I2595,I318922,I318911,);
nor I_18626 (I319264,I184203,I184191);
nor I_18627 (I318902,I319117,I319264);
or I_18628 (I319295,I184203,I184191);
nor I_18629 (I319312,I184182,I184185);
DFFARX1 I_18630 (I319312,I2595,I318922,I319338,);
not I_18631 (I319346,I319338);
nor I_18632 (I318908,I319346,I319151);
nand I_18633 (I319377,I319346,I318996);
not I_18634 (I319394,I184182);
nand I_18635 (I319411,I319394,I319100);
nand I_18636 (I319428,I319346,I319411);
nand I_18637 (I318899,I319428,I319377);
nand I_18638 (I318896,I319411,I319295);
not I_18639 (I319500,I2602);
DFFARX1 I_18640 (I258325,I2595,I319500,I319526,);
and I_18641 (I319534,I319526,I258319);
DFFARX1 I_18642 (I319534,I2595,I319500,I319483,);
DFFARX1 I_18643 (I258337,I2595,I319500,I319574,);
not I_18644 (I319582,I258328);
not I_18645 (I319599,I258340);
nand I_18646 (I319616,I319599,I319582);
nor I_18647 (I319471,I319574,I319616);
DFFARX1 I_18648 (I319616,I2595,I319500,I319656,);
not I_18649 (I319492,I319656);
not I_18650 (I319678,I258346);
nand I_18651 (I319695,I319599,I319678);
DFFARX1 I_18652 (I319695,I2595,I319500,I319721,);
not I_18653 (I319729,I319721);
not I_18654 (I319746,I258322);
nand I_18655 (I319763,I319746,I258343);
and I_18656 (I319780,I319582,I319763);
nor I_18657 (I319797,I319695,I319780);
DFFARX1 I_18658 (I319797,I2595,I319500,I319468,);
DFFARX1 I_18659 (I319780,I2595,I319500,I319489,);
nor I_18660 (I319842,I258322,I258334);
nor I_18661 (I319480,I319695,I319842);
or I_18662 (I319873,I258322,I258334);
nor I_18663 (I319890,I258319,I258331);
DFFARX1 I_18664 (I319890,I2595,I319500,I319916,);
not I_18665 (I319924,I319916);
nor I_18666 (I319486,I319924,I319729);
nand I_18667 (I319955,I319924,I319574);
not I_18668 (I319972,I258319);
nand I_18669 (I319989,I319972,I319678);
nand I_18670 (I320006,I319924,I319989);
nand I_18671 (I319477,I320006,I319955);
nand I_18672 (I319474,I319989,I319873);
not I_18673 (I320078,I2602);
DFFARX1 I_18674 (I141583,I2595,I320078,I320104,);
and I_18675 (I320112,I320104,I141598);
DFFARX1 I_18676 (I320112,I2595,I320078,I320061,);
DFFARX1 I_18677 (I141589,I2595,I320078,I320152,);
not I_18678 (I320160,I141583);
not I_18679 (I320177,I141601);
nand I_18680 (I320194,I320177,I320160);
nor I_18681 (I320049,I320152,I320194);
DFFARX1 I_18682 (I320194,I2595,I320078,I320234,);
not I_18683 (I320070,I320234);
not I_18684 (I320256,I141592);
nand I_18685 (I320273,I320177,I320256);
DFFARX1 I_18686 (I320273,I2595,I320078,I320299,);
not I_18687 (I320307,I320299);
not I_18688 (I320324,I141604);
nand I_18689 (I320341,I320324,I141580);
and I_18690 (I320358,I320160,I320341);
nor I_18691 (I320375,I320273,I320358);
DFFARX1 I_18692 (I320375,I2595,I320078,I320046,);
DFFARX1 I_18693 (I320358,I2595,I320078,I320067,);
nor I_18694 (I320420,I141604,I141580);
nor I_18695 (I320058,I320273,I320420);
or I_18696 (I320451,I141604,I141580);
nor I_18697 (I320468,I141586,I141595);
DFFARX1 I_18698 (I320468,I2595,I320078,I320494,);
not I_18699 (I320502,I320494);
nor I_18700 (I320064,I320502,I320307);
nand I_18701 (I320533,I320502,I320152);
not I_18702 (I320550,I141586);
nand I_18703 (I320567,I320550,I320256);
nand I_18704 (I320584,I320502,I320567);
nand I_18705 (I320055,I320584,I320533);
nand I_18706 (I320052,I320567,I320451);
not I_18707 (I320656,I2602);
DFFARX1 I_18708 (I110684,I2595,I320656,I320682,);
and I_18709 (I320690,I320682,I110669);
DFFARX1 I_18710 (I320690,I2595,I320656,I320639,);
DFFARX1 I_18711 (I110675,I2595,I320656,I320730,);
not I_18712 (I320738,I110657);
not I_18713 (I320755,I110678);
nand I_18714 (I320772,I320755,I320738);
nor I_18715 (I320627,I320730,I320772);
DFFARX1 I_18716 (I320772,I2595,I320656,I320812,);
not I_18717 (I320648,I320812);
not I_18718 (I320834,I110681);
nand I_18719 (I320851,I320755,I320834);
DFFARX1 I_18720 (I320851,I2595,I320656,I320877,);
not I_18721 (I320885,I320877);
not I_18722 (I320902,I110672);
nand I_18723 (I320919,I320902,I110660);
and I_18724 (I320936,I320738,I320919);
nor I_18725 (I320953,I320851,I320936);
DFFARX1 I_18726 (I320953,I2595,I320656,I320624,);
DFFARX1 I_18727 (I320936,I2595,I320656,I320645,);
nor I_18728 (I320998,I110672,I110666);
nor I_18729 (I320636,I320851,I320998);
or I_18730 (I321029,I110672,I110666);
nor I_18731 (I321046,I110663,I110657);
DFFARX1 I_18732 (I321046,I2595,I320656,I321072,);
not I_18733 (I321080,I321072);
nor I_18734 (I320642,I321080,I320885);
nand I_18735 (I321111,I321080,I320730);
not I_18736 (I321128,I110663);
nand I_18737 (I321145,I321128,I320834);
nand I_18738 (I321162,I321080,I321145);
nand I_18739 (I320633,I321162,I321111);
nand I_18740 (I320630,I321145,I321029);
not I_18741 (I321234,I2602);
DFFARX1 I_18742 (I63958,I2595,I321234,I321260,);
and I_18743 (I321268,I321260,I63961);
DFFARX1 I_18744 (I321268,I2595,I321234,I321217,);
DFFARX1 I_18745 (I63961,I2595,I321234,I321308,);
not I_18746 (I321316,I63976);
not I_18747 (I321333,I63982);
nand I_18748 (I321350,I321333,I321316);
nor I_18749 (I321205,I321308,I321350);
DFFARX1 I_18750 (I321350,I2595,I321234,I321390,);
not I_18751 (I321226,I321390);
not I_18752 (I321412,I63970);
nand I_18753 (I321429,I321333,I321412);
DFFARX1 I_18754 (I321429,I2595,I321234,I321455,);
not I_18755 (I321463,I321455);
not I_18756 (I321480,I63967);
nand I_18757 (I321497,I321480,I63964);
and I_18758 (I321514,I321316,I321497);
nor I_18759 (I321531,I321429,I321514);
DFFARX1 I_18760 (I321531,I2595,I321234,I321202,);
DFFARX1 I_18761 (I321514,I2595,I321234,I321223,);
nor I_18762 (I321576,I63967,I63958);
nor I_18763 (I321214,I321429,I321576);
or I_18764 (I321607,I63967,I63958);
nor I_18765 (I321624,I63973,I63979);
DFFARX1 I_18766 (I321624,I2595,I321234,I321650,);
not I_18767 (I321658,I321650);
nor I_18768 (I321220,I321658,I321463);
nand I_18769 (I321689,I321658,I321308);
not I_18770 (I321706,I63973);
nand I_18771 (I321723,I321706,I321412);
nand I_18772 (I321740,I321658,I321723);
nand I_18773 (I321211,I321740,I321689);
nand I_18774 (I321208,I321723,I321607);
not I_18775 (I321812,I2602);
DFFARX1 I_18776 (I23471,I2595,I321812,I321838,);
and I_18777 (I321846,I321838,I23447);
DFFARX1 I_18778 (I321846,I2595,I321812,I321795,);
DFFARX1 I_18779 (I23465,I2595,I321812,I321886,);
not I_18780 (I321894,I23453);
not I_18781 (I321911,I23450);
nand I_18782 (I321928,I321911,I321894);
nor I_18783 (I321783,I321886,I321928);
DFFARX1 I_18784 (I321928,I2595,I321812,I321968,);
not I_18785 (I321804,I321968);
not I_18786 (I321990,I23459);
nand I_18787 (I322007,I321911,I321990);
DFFARX1 I_18788 (I322007,I2595,I321812,I322033,);
not I_18789 (I322041,I322033);
not I_18790 (I322058,I23450);
nand I_18791 (I322075,I322058,I23468);
and I_18792 (I322092,I321894,I322075);
nor I_18793 (I322109,I322007,I322092);
DFFARX1 I_18794 (I322109,I2595,I321812,I321780,);
DFFARX1 I_18795 (I322092,I2595,I321812,I321801,);
nor I_18796 (I322154,I23450,I23462);
nor I_18797 (I321792,I322007,I322154);
or I_18798 (I322185,I23450,I23462);
nor I_18799 (I322202,I23456,I23447);
DFFARX1 I_18800 (I322202,I2595,I321812,I322228,);
not I_18801 (I322236,I322228);
nor I_18802 (I321798,I322236,I322041);
nand I_18803 (I322267,I322236,I321886);
not I_18804 (I322284,I23456);
nand I_18805 (I322301,I322284,I321990);
nand I_18806 (I322318,I322236,I322301);
nand I_18807 (I321789,I322318,I322267);
nand I_18808 (I321786,I322301,I322185);
not I_18809 (I322390,I2602);
DFFARX1 I_18810 (I296062,I2595,I322390,I322416,);
and I_18811 (I322424,I322416,I296059);
DFFARX1 I_18812 (I322424,I2595,I322390,I322373,);
DFFARX1 I_18813 (I296065,I2595,I322390,I322464,);
not I_18814 (I322472,I296068);
not I_18815 (I322489,I296062);
nand I_18816 (I322506,I322489,I322472);
nor I_18817 (I322361,I322464,I322506);
DFFARX1 I_18818 (I322506,I2595,I322390,I322546,);
not I_18819 (I322382,I322546);
not I_18820 (I322568,I296077);
nand I_18821 (I322585,I322489,I322568);
DFFARX1 I_18822 (I322585,I2595,I322390,I322611,);
not I_18823 (I322619,I322611);
not I_18824 (I322636,I296074);
nand I_18825 (I322653,I322636,I296080);
and I_18826 (I322670,I322472,I322653);
nor I_18827 (I322687,I322585,I322670);
DFFARX1 I_18828 (I322687,I2595,I322390,I322358,);
DFFARX1 I_18829 (I322670,I2595,I322390,I322379,);
nor I_18830 (I322732,I296074,I296059);
nor I_18831 (I322370,I322585,I322732);
or I_18832 (I322763,I296074,I296059);
nor I_18833 (I322780,I296071,I296065);
DFFARX1 I_18834 (I322780,I2595,I322390,I322806,);
not I_18835 (I322814,I322806);
nor I_18836 (I322376,I322814,I322619);
nand I_18837 (I322845,I322814,I322464);
not I_18838 (I322862,I296071);
nand I_18839 (I322879,I322862,I322568);
nand I_18840 (I322896,I322814,I322879);
nand I_18841 (I322367,I322896,I322845);
nand I_18842 (I322364,I322879,I322763);
not I_18843 (I322968,I2602);
DFFARX1 I_18844 (I124665,I2595,I322968,I322994,);
and I_18845 (I323002,I322994,I124680);
DFFARX1 I_18846 (I323002,I2595,I322968,I322951,);
DFFARX1 I_18847 (I124683,I2595,I322968,I323042,);
not I_18848 (I323050,I124677);
not I_18849 (I323067,I124692);
nand I_18850 (I323084,I323067,I323050);
nor I_18851 (I322939,I323042,I323084);
DFFARX1 I_18852 (I323084,I2595,I322968,I323124,);
not I_18853 (I322960,I323124);
not I_18854 (I323146,I124668);
nand I_18855 (I323163,I323067,I323146);
DFFARX1 I_18856 (I323163,I2595,I322968,I323189,);
not I_18857 (I323197,I323189);
not I_18858 (I323214,I124671);
nand I_18859 (I323231,I323214,I124665);
and I_18860 (I323248,I323050,I323231);
nor I_18861 (I323265,I323163,I323248);
DFFARX1 I_18862 (I323265,I2595,I322968,I322936,);
DFFARX1 I_18863 (I323248,I2595,I322968,I322957,);
nor I_18864 (I323310,I124671,I124674);
nor I_18865 (I322948,I323163,I323310);
or I_18866 (I323341,I124671,I124674);
nor I_18867 (I323358,I124689,I124686);
DFFARX1 I_18868 (I323358,I2595,I322968,I323384,);
not I_18869 (I323392,I323384);
nor I_18870 (I322954,I323392,I323197);
nand I_18871 (I323423,I323392,I323042);
not I_18872 (I323440,I124689);
nand I_18873 (I323457,I323440,I323146);
nand I_18874 (I323474,I323392,I323457);
nand I_18875 (I322945,I323474,I323423);
nand I_18876 (I322942,I323457,I323341);
not I_18877 (I323546,I2602);
DFFARX1 I_18878 (I46703,I2595,I323546,I323572,);
and I_18879 (I323580,I323572,I46727);
DFFARX1 I_18880 (I323580,I2595,I323546,I323529,);
DFFARX1 I_18881 (I46703,I2595,I323546,I323620,);
not I_18882 (I323628,I46721);
not I_18883 (I323645,I46706);
nand I_18884 (I323662,I323645,I323628);
nor I_18885 (I323517,I323620,I323662);
DFFARX1 I_18886 (I323662,I2595,I323546,I323702,);
not I_18887 (I323538,I323702);
not I_18888 (I323724,I46715);
nand I_18889 (I323741,I323645,I323724);
DFFARX1 I_18890 (I323741,I2595,I323546,I323767,);
not I_18891 (I323775,I323767);
not I_18892 (I323792,I46712);
nand I_18893 (I323809,I323792,I46709);
and I_18894 (I323826,I323628,I323809);
nor I_18895 (I323843,I323741,I323826);
DFFARX1 I_18896 (I323843,I2595,I323546,I323514,);
DFFARX1 I_18897 (I323826,I2595,I323546,I323535,);
nor I_18898 (I323888,I46712,I46718);
nor I_18899 (I323526,I323741,I323888);
or I_18900 (I323919,I46712,I46718);
nor I_18901 (I323936,I46724,I46730);
DFFARX1 I_18902 (I323936,I2595,I323546,I323962,);
not I_18903 (I323970,I323962);
nor I_18904 (I323532,I323970,I323775);
nand I_18905 (I324001,I323970,I323620);
not I_18906 (I324018,I46724);
nand I_18907 (I324035,I324018,I323724);
nand I_18908 (I324052,I323970,I324035);
nand I_18909 (I323523,I324052,I324001);
nand I_18910 (I323520,I324035,I323919);
not I_18911 (I324124,I2602);
DFFARX1 I_18912 (I278351,I2595,I324124,I324150,);
and I_18913 (I324158,I324150,I278345);
DFFARX1 I_18914 (I324158,I2595,I324124,I324107,);
DFFARX1 I_18915 (I278363,I2595,I324124,I324198,);
not I_18916 (I324206,I278354);
not I_18917 (I324223,I278366);
nand I_18918 (I324240,I324223,I324206);
nor I_18919 (I324095,I324198,I324240);
DFFARX1 I_18920 (I324240,I2595,I324124,I324280,);
not I_18921 (I324116,I324280);
not I_18922 (I324302,I278372);
nand I_18923 (I324319,I324223,I324302);
DFFARX1 I_18924 (I324319,I2595,I324124,I324345,);
not I_18925 (I324353,I324345);
not I_18926 (I324370,I278348);
nand I_18927 (I324387,I324370,I278369);
and I_18928 (I324404,I324206,I324387);
nor I_18929 (I324421,I324319,I324404);
DFFARX1 I_18930 (I324421,I2595,I324124,I324092,);
DFFARX1 I_18931 (I324404,I2595,I324124,I324113,);
nor I_18932 (I324466,I278348,I278360);
nor I_18933 (I324104,I324319,I324466);
or I_18934 (I324497,I278348,I278360);
nor I_18935 (I324514,I278345,I278357);
DFFARX1 I_18936 (I324514,I2595,I324124,I324540,);
not I_18937 (I324548,I324540);
nor I_18938 (I324110,I324548,I324353);
nand I_18939 (I324579,I324548,I324198);
not I_18940 (I324596,I278345);
nand I_18941 (I324613,I324596,I324302);
nand I_18942 (I324630,I324548,I324613);
nand I_18943 (I324101,I324630,I324579);
nand I_18944 (I324098,I324613,I324497);
not I_18945 (I324702,I2602);
DFFARX1 I_18946 (I238279,I2595,I324702,I324728,);
and I_18947 (I324736,I324728,I238285);
DFFARX1 I_18948 (I324736,I2595,I324702,I324685,);
DFFARX1 I_18949 (I238291,I2595,I324702,I324776,);
not I_18950 (I324784,I238276);
not I_18951 (I324801,I238276);
nand I_18952 (I324818,I324801,I324784);
nor I_18953 (I324673,I324776,I324818);
DFFARX1 I_18954 (I324818,I2595,I324702,I324858,);
not I_18955 (I324694,I324858);
not I_18956 (I324880,I238294);
nand I_18957 (I324897,I324801,I324880);
DFFARX1 I_18958 (I324897,I2595,I324702,I324923,);
not I_18959 (I324931,I324923);
not I_18960 (I324948,I238288);
nand I_18961 (I324965,I324948,I238279);
and I_18962 (I324982,I324784,I324965);
nor I_18963 (I324999,I324897,I324982);
DFFARX1 I_18964 (I324999,I2595,I324702,I324670,);
DFFARX1 I_18965 (I324982,I2595,I324702,I324691,);
nor I_18966 (I325044,I238288,I238297);
nor I_18967 (I324682,I324897,I325044);
or I_18968 (I325075,I238288,I238297);
nor I_18969 (I325092,I238282,I238282);
DFFARX1 I_18970 (I325092,I2595,I324702,I325118,);
not I_18971 (I325126,I325118);
nor I_18972 (I324688,I325126,I324931);
nand I_18973 (I325157,I325126,I324776);
not I_18974 (I325174,I238282);
nand I_18975 (I325191,I325174,I324880);
nand I_18976 (I325208,I325126,I325191);
nand I_18977 (I324679,I325208,I325157);
nand I_18978 (I324676,I325191,I325075);
not I_18979 (I325280,I2602);
DFFARX1 I_18980 (I215987,I2595,I325280,I325306,);
and I_18981 (I325314,I325306,I215975);
DFFARX1 I_18982 (I325314,I2595,I325280,I325263,);
DFFARX1 I_18983 (I215978,I2595,I325280,I325354,);
not I_18984 (I325362,I215972);
not I_18985 (I325379,I215996);
nand I_18986 (I325396,I325379,I325362);
nor I_18987 (I325251,I325354,I325396);
DFFARX1 I_18988 (I325396,I2595,I325280,I325436,);
not I_18989 (I325272,I325436);
not I_18990 (I325458,I215984);
nand I_18991 (I325475,I325379,I325458);
DFFARX1 I_18992 (I325475,I2595,I325280,I325501,);
not I_18993 (I325509,I325501);
not I_18994 (I325526,I215993);
nand I_18995 (I325543,I325526,I215990);
and I_18996 (I325560,I325362,I325543);
nor I_18997 (I325577,I325475,I325560);
DFFARX1 I_18998 (I325577,I2595,I325280,I325248,);
DFFARX1 I_18999 (I325560,I2595,I325280,I325269,);
nor I_19000 (I325622,I215993,I215981);
nor I_19001 (I325260,I325475,I325622);
or I_19002 (I325653,I215993,I215981);
nor I_19003 (I325670,I215972,I215975);
DFFARX1 I_19004 (I325670,I2595,I325280,I325696,);
not I_19005 (I325704,I325696);
nor I_19006 (I325266,I325704,I325509);
nand I_19007 (I325735,I325704,I325354);
not I_19008 (I325752,I215972);
nand I_19009 (I325769,I325752,I325458);
nand I_19010 (I325786,I325704,I325769);
nand I_19011 (I325257,I325786,I325735);
nand I_19012 (I325254,I325769,I325653);
not I_19013 (I325858,I2602);
DFFARX1 I_19014 (I107522,I2595,I325858,I325884,);
and I_19015 (I325892,I325884,I107507);
DFFARX1 I_19016 (I325892,I2595,I325858,I325841,);
DFFARX1 I_19017 (I107513,I2595,I325858,I325932,);
not I_19018 (I325940,I107495);
not I_19019 (I325957,I107516);
nand I_19020 (I325974,I325957,I325940);
nor I_19021 (I325829,I325932,I325974);
DFFARX1 I_19022 (I325974,I2595,I325858,I326014,);
not I_19023 (I325850,I326014);
not I_19024 (I326036,I107519);
nand I_19025 (I326053,I325957,I326036);
DFFARX1 I_19026 (I326053,I2595,I325858,I326079,);
not I_19027 (I326087,I326079);
not I_19028 (I326104,I107510);
nand I_19029 (I326121,I326104,I107498);
and I_19030 (I326138,I325940,I326121);
nor I_19031 (I326155,I326053,I326138);
DFFARX1 I_19032 (I326155,I2595,I325858,I325826,);
DFFARX1 I_19033 (I326138,I2595,I325858,I325847,);
nor I_19034 (I326200,I107510,I107504);
nor I_19035 (I325838,I326053,I326200);
or I_19036 (I326231,I107510,I107504);
nor I_19037 (I326248,I107501,I107495);
DFFARX1 I_19038 (I326248,I2595,I325858,I326274,);
not I_19039 (I326282,I326274);
nor I_19040 (I325844,I326282,I326087);
nand I_19041 (I326313,I326282,I325932);
not I_19042 (I326330,I107501);
nand I_19043 (I326347,I326330,I326036);
nand I_19044 (I326364,I326282,I326347);
nand I_19045 (I325835,I326364,I326313);
nand I_19046 (I325832,I326347,I326231);
not I_19047 (I326436,I2602);
DFFARX1 I_19048 (I359102,I2595,I326436,I326462,);
and I_19049 (I326470,I326462,I359084);
DFFARX1 I_19050 (I326470,I2595,I326436,I326419,);
DFFARX1 I_19051 (I359093,I2595,I326436,I326510,);
not I_19052 (I326518,I359078);
not I_19053 (I326535,I359090);
nand I_19054 (I326552,I326535,I326518);
nor I_19055 (I326407,I326510,I326552);
DFFARX1 I_19056 (I326552,I2595,I326436,I326592,);
not I_19057 (I326428,I326592);
not I_19058 (I326614,I359081);
nand I_19059 (I326631,I326535,I326614);
DFFARX1 I_19060 (I326631,I2595,I326436,I326657,);
not I_19061 (I326665,I326657);
not I_19062 (I326682,I359078);
nand I_19063 (I326699,I326682,I359081);
and I_19064 (I326716,I326518,I326699);
nor I_19065 (I326733,I326631,I326716);
DFFARX1 I_19066 (I326733,I2595,I326436,I326404,);
DFFARX1 I_19067 (I326716,I2595,I326436,I326425,);
nor I_19068 (I326778,I359078,I359099);
nor I_19069 (I326416,I326631,I326778);
or I_19070 (I326809,I359078,I359099);
nor I_19071 (I326826,I359087,I359096);
DFFARX1 I_19072 (I326826,I2595,I326436,I326852,);
not I_19073 (I326860,I326852);
nor I_19074 (I326422,I326860,I326665);
nand I_19075 (I326891,I326860,I326510);
not I_19076 (I326908,I359087);
nand I_19077 (I326925,I326908,I326614);
nand I_19078 (I326942,I326860,I326925);
nand I_19079 (I326413,I326942,I326891);
nand I_19080 (I326410,I326925,I326809);
not I_19081 (I327014,I2602);
DFFARX1 I_19082 (I123033,I2595,I327014,I327040,);
and I_19083 (I327048,I327040,I123048);
DFFARX1 I_19084 (I327048,I2595,I327014,I326997,);
DFFARX1 I_19085 (I123051,I2595,I327014,I327088,);
not I_19086 (I327096,I123045);
not I_19087 (I327113,I123060);
nand I_19088 (I327130,I327113,I327096);
nor I_19089 (I326985,I327088,I327130);
DFFARX1 I_19090 (I327130,I2595,I327014,I327170,);
not I_19091 (I327006,I327170);
not I_19092 (I327192,I123036);
nand I_19093 (I327209,I327113,I327192);
DFFARX1 I_19094 (I327209,I2595,I327014,I327235,);
not I_19095 (I327243,I327235);
not I_19096 (I327260,I123039);
nand I_19097 (I327277,I327260,I123033);
and I_19098 (I327294,I327096,I327277);
nor I_19099 (I327311,I327209,I327294);
DFFARX1 I_19100 (I327311,I2595,I327014,I326982,);
DFFARX1 I_19101 (I327294,I2595,I327014,I327003,);
nor I_19102 (I327356,I123039,I123042);
nor I_19103 (I326994,I327209,I327356);
or I_19104 (I327387,I123039,I123042);
nor I_19105 (I327404,I123057,I123054);
DFFARX1 I_19106 (I327404,I2595,I327014,I327430,);
not I_19107 (I327438,I327430);
nor I_19108 (I327000,I327438,I327243);
nand I_19109 (I327469,I327438,I327088);
not I_19110 (I327486,I123057);
nand I_19111 (I327503,I327486,I327192);
nand I_19112 (I327520,I327438,I327503);
nand I_19113 (I326991,I327520,I327469);
nand I_19114 (I326988,I327503,I327387);
not I_19115 (I327592,I2602);
DFFARX1 I_19116 (I117593,I2595,I327592,I327618,);
and I_19117 (I327626,I327618,I117608);
DFFARX1 I_19118 (I327626,I2595,I327592,I327575,);
DFFARX1 I_19119 (I117611,I2595,I327592,I327666,);
not I_19120 (I327674,I117605);
not I_19121 (I327691,I117620);
nand I_19122 (I327708,I327691,I327674);
nor I_19123 (I327563,I327666,I327708);
DFFARX1 I_19124 (I327708,I2595,I327592,I327748,);
not I_19125 (I327584,I327748);
not I_19126 (I327770,I117596);
nand I_19127 (I327787,I327691,I327770);
DFFARX1 I_19128 (I327787,I2595,I327592,I327813,);
not I_19129 (I327821,I327813);
not I_19130 (I327838,I117599);
nand I_19131 (I327855,I327838,I117593);
and I_19132 (I327872,I327674,I327855);
nor I_19133 (I327889,I327787,I327872);
DFFARX1 I_19134 (I327889,I2595,I327592,I327560,);
DFFARX1 I_19135 (I327872,I2595,I327592,I327581,);
nor I_19136 (I327934,I117599,I117602);
nor I_19137 (I327572,I327787,I327934);
or I_19138 (I327965,I117599,I117602);
nor I_19139 (I327982,I117617,I117614);
DFFARX1 I_19140 (I327982,I2595,I327592,I328008,);
not I_19141 (I328016,I328008);
nor I_19142 (I327578,I328016,I327821);
nand I_19143 (I328047,I328016,I327666);
not I_19144 (I328064,I117617);
nand I_19145 (I328081,I328064,I327770);
nand I_19146 (I328098,I328016,I328081);
nand I_19147 (I327569,I328098,I328047);
nand I_19148 (I327566,I328081,I327965);
not I_19149 (I328170,I2602);
DFFARX1 I_19150 (I56223,I2595,I328170,I328196,);
and I_19151 (I328204,I328196,I56226);
DFFARX1 I_19152 (I328204,I2595,I328170,I328153,);
DFFARX1 I_19153 (I56226,I2595,I328170,I328244,);
not I_19154 (I328252,I56241);
not I_19155 (I328269,I56247);
nand I_19156 (I328286,I328269,I328252);
nor I_19157 (I328141,I328244,I328286);
DFFARX1 I_19158 (I328286,I2595,I328170,I328326,);
not I_19159 (I328162,I328326);
not I_19160 (I328348,I56235);
nand I_19161 (I328365,I328269,I328348);
DFFARX1 I_19162 (I328365,I2595,I328170,I328391,);
not I_19163 (I328399,I328391);
not I_19164 (I328416,I56232);
nand I_19165 (I328433,I328416,I56229);
and I_19166 (I328450,I328252,I328433);
nor I_19167 (I328467,I328365,I328450);
DFFARX1 I_19168 (I328467,I2595,I328170,I328138,);
DFFARX1 I_19169 (I328450,I2595,I328170,I328159,);
nor I_19170 (I328512,I56232,I56223);
nor I_19171 (I328150,I328365,I328512);
or I_19172 (I328543,I56232,I56223);
nor I_19173 (I328560,I56238,I56244);
DFFARX1 I_19174 (I328560,I2595,I328170,I328586,);
not I_19175 (I328594,I328586);
nor I_19176 (I328156,I328594,I328399);
nand I_19177 (I328625,I328594,I328244);
not I_19178 (I328642,I56238);
nand I_19179 (I328659,I328642,I328348);
nand I_19180 (I328676,I328594,I328659);
nand I_19181 (I328147,I328676,I328625);
nand I_19182 (I328144,I328659,I328543);
not I_19183 (I328748,I2602);
DFFARX1 I_19184 (I192867,I2595,I328748,I328774,);
and I_19185 (I328782,I328774,I192855);
DFFARX1 I_19186 (I328782,I2595,I328748,I328731,);
DFFARX1 I_19187 (I192858,I2595,I328748,I328822,);
not I_19188 (I328830,I192852);
not I_19189 (I328847,I192876);
nand I_19190 (I328864,I328847,I328830);
nor I_19191 (I328719,I328822,I328864);
DFFARX1 I_19192 (I328864,I2595,I328748,I328904,);
not I_19193 (I328740,I328904);
not I_19194 (I328926,I192864);
nand I_19195 (I328943,I328847,I328926);
DFFARX1 I_19196 (I328943,I2595,I328748,I328969,);
not I_19197 (I328977,I328969);
not I_19198 (I328994,I192873);
nand I_19199 (I329011,I328994,I192870);
and I_19200 (I329028,I328830,I329011);
nor I_19201 (I329045,I328943,I329028);
DFFARX1 I_19202 (I329045,I2595,I328748,I328716,);
DFFARX1 I_19203 (I329028,I2595,I328748,I328737,);
nor I_19204 (I329090,I192873,I192861);
nor I_19205 (I328728,I328943,I329090);
or I_19206 (I329121,I192873,I192861);
nor I_19207 (I329138,I192852,I192855);
DFFARX1 I_19208 (I329138,I2595,I328748,I329164,);
not I_19209 (I329172,I329164);
nor I_19210 (I328734,I329172,I328977);
nand I_19211 (I329203,I329172,I328822);
not I_19212 (I329220,I192852);
nand I_19213 (I329237,I329220,I328926);
nand I_19214 (I329254,I329172,I329237);
nand I_19215 (I328725,I329254,I329203);
nand I_19216 (I328722,I329237,I329121);
not I_19217 (I329326,I2602);
DFFARX1 I_19218 (I70503,I2595,I329326,I329352,);
and I_19219 (I329360,I329352,I70506);
DFFARX1 I_19220 (I329360,I2595,I329326,I329309,);
DFFARX1 I_19221 (I70506,I2595,I329326,I329400,);
not I_19222 (I329408,I70521);
not I_19223 (I329425,I70527);
nand I_19224 (I329442,I329425,I329408);
nor I_19225 (I329297,I329400,I329442);
DFFARX1 I_19226 (I329442,I2595,I329326,I329482,);
not I_19227 (I329318,I329482);
not I_19228 (I329504,I70515);
nand I_19229 (I329521,I329425,I329504);
DFFARX1 I_19230 (I329521,I2595,I329326,I329547,);
not I_19231 (I329555,I329547);
not I_19232 (I329572,I70512);
nand I_19233 (I329589,I329572,I70509);
and I_19234 (I329606,I329408,I329589);
nor I_19235 (I329623,I329521,I329606);
DFFARX1 I_19236 (I329623,I2595,I329326,I329294,);
DFFARX1 I_19237 (I329606,I2595,I329326,I329315,);
nor I_19238 (I329668,I70512,I70503);
nor I_19239 (I329306,I329521,I329668);
or I_19240 (I329699,I70512,I70503);
nor I_19241 (I329716,I70518,I70524);
DFFARX1 I_19242 (I329716,I2595,I329326,I329742,);
not I_19243 (I329750,I329742);
nor I_19244 (I329312,I329750,I329555);
nand I_19245 (I329781,I329750,I329400);
not I_19246 (I329798,I70518);
nand I_19247 (I329815,I329798,I329504);
nand I_19248 (I329832,I329750,I329815);
nand I_19249 (I329303,I329832,I329781);
nand I_19250 (I329300,I329815,I329699);
not I_19251 (I329904,I2602);
DFFARX1 I_19252 (I188821,I2595,I329904,I329930,);
and I_19253 (I329938,I329930,I188809);
DFFARX1 I_19254 (I329938,I2595,I329904,I329887,);
DFFARX1 I_19255 (I188812,I2595,I329904,I329978,);
not I_19256 (I329986,I188806);
not I_19257 (I330003,I188830);
nand I_19258 (I330020,I330003,I329986);
nor I_19259 (I329875,I329978,I330020);
DFFARX1 I_19260 (I330020,I2595,I329904,I330060,);
not I_19261 (I329896,I330060);
not I_19262 (I330082,I188818);
nand I_19263 (I330099,I330003,I330082);
DFFARX1 I_19264 (I330099,I2595,I329904,I330125,);
not I_19265 (I330133,I330125);
not I_19266 (I330150,I188827);
nand I_19267 (I330167,I330150,I188824);
and I_19268 (I330184,I329986,I330167);
nor I_19269 (I330201,I330099,I330184);
DFFARX1 I_19270 (I330201,I2595,I329904,I329872,);
DFFARX1 I_19271 (I330184,I2595,I329904,I329893,);
nor I_19272 (I330246,I188827,I188815);
nor I_19273 (I329884,I330099,I330246);
or I_19274 (I330277,I188827,I188815);
nor I_19275 (I330294,I188806,I188809);
DFFARX1 I_19276 (I330294,I2595,I329904,I330320,);
not I_19277 (I330328,I330320);
nor I_19278 (I329890,I330328,I330133);
nand I_19279 (I330359,I330328,I329978);
not I_19280 (I330376,I188806);
nand I_19281 (I330393,I330376,I330082);
nand I_19282 (I330410,I330328,I330393);
nand I_19283 (I329881,I330410,I330359);
nand I_19284 (I329878,I330393,I330277);
not I_19285 (I330482,I2602);
DFFARX1 I_19286 (I371175,I2595,I330482,I330508,);
and I_19287 (I330516,I330508,I371157);
DFFARX1 I_19288 (I330516,I2595,I330482,I330465,);
DFFARX1 I_19289 (I371148,I2595,I330482,I330556,);
not I_19290 (I330564,I371163);
not I_19291 (I330581,I371151);
nand I_19292 (I330598,I330581,I330564);
nor I_19293 (I330453,I330556,I330598);
DFFARX1 I_19294 (I330598,I2595,I330482,I330638,);
not I_19295 (I330474,I330638);
not I_19296 (I330660,I371160);
nand I_19297 (I330677,I330581,I330660);
DFFARX1 I_19298 (I330677,I2595,I330482,I330703,);
not I_19299 (I330711,I330703);
not I_19300 (I330728,I371169);
nand I_19301 (I330745,I330728,I371148);
and I_19302 (I330762,I330564,I330745);
nor I_19303 (I330779,I330677,I330762);
DFFARX1 I_19304 (I330779,I2595,I330482,I330450,);
DFFARX1 I_19305 (I330762,I2595,I330482,I330471,);
nor I_19306 (I330824,I371169,I371172);
nor I_19307 (I330462,I330677,I330824);
or I_19308 (I330855,I371169,I371172);
nor I_19309 (I330872,I371166,I371154);
DFFARX1 I_19310 (I330872,I2595,I330482,I330898,);
not I_19311 (I330906,I330898);
nor I_19312 (I330468,I330906,I330711);
nand I_19313 (I330937,I330906,I330556);
not I_19314 (I330954,I371166);
nand I_19315 (I330971,I330954,I330660);
nand I_19316 (I330988,I330906,I330971);
nand I_19317 (I330459,I330988,I330937);
nand I_19318 (I330456,I330971,I330855);
not I_19319 (I331060,I2602);
DFFARX1 I_19320 (I234063,I2595,I331060,I331086,);
and I_19321 (I331094,I331086,I234069);
DFFARX1 I_19322 (I331094,I2595,I331060,I331043,);
DFFARX1 I_19323 (I234075,I2595,I331060,I331134,);
not I_19324 (I331142,I234060);
not I_19325 (I331159,I234060);
nand I_19326 (I331176,I331159,I331142);
nor I_19327 (I331031,I331134,I331176);
DFFARX1 I_19328 (I331176,I2595,I331060,I331216,);
not I_19329 (I331052,I331216);
not I_19330 (I331238,I234078);
nand I_19331 (I331255,I331159,I331238);
DFFARX1 I_19332 (I331255,I2595,I331060,I331281,);
not I_19333 (I331289,I331281);
not I_19334 (I331306,I234072);
nand I_19335 (I331323,I331306,I234063);
and I_19336 (I331340,I331142,I331323);
nor I_19337 (I331357,I331255,I331340);
DFFARX1 I_19338 (I331357,I2595,I331060,I331028,);
DFFARX1 I_19339 (I331340,I2595,I331060,I331049,);
nor I_19340 (I331402,I234072,I234081);
nor I_19341 (I331040,I331255,I331402);
or I_19342 (I331433,I234072,I234081);
nor I_19343 (I331450,I234066,I234066);
DFFARX1 I_19344 (I331450,I2595,I331060,I331476,);
not I_19345 (I331484,I331476);
nor I_19346 (I331046,I331484,I331289);
nand I_19347 (I331515,I331484,I331134);
not I_19348 (I331532,I234066);
nand I_19349 (I331549,I331532,I331238);
nand I_19350 (I331566,I331484,I331549);
nand I_19351 (I331037,I331566,I331515);
nand I_19352 (I331034,I331549,I331433);
not I_19353 (I331638,I2602);
DFFARX1 I_19354 (I85388,I2595,I331638,I331664,);
and I_19355 (I331672,I331664,I85373);
DFFARX1 I_19356 (I331672,I2595,I331638,I331621,);
DFFARX1 I_19357 (I85379,I2595,I331638,I331712,);
not I_19358 (I331720,I85361);
not I_19359 (I331737,I85382);
nand I_19360 (I331754,I331737,I331720);
nor I_19361 (I331609,I331712,I331754);
DFFARX1 I_19362 (I331754,I2595,I331638,I331794,);
not I_19363 (I331630,I331794);
not I_19364 (I331816,I85385);
nand I_19365 (I331833,I331737,I331816);
DFFARX1 I_19366 (I331833,I2595,I331638,I331859,);
not I_19367 (I331867,I331859);
not I_19368 (I331884,I85376);
nand I_19369 (I331901,I331884,I85364);
and I_19370 (I331918,I331720,I331901);
nor I_19371 (I331935,I331833,I331918);
DFFARX1 I_19372 (I331935,I2595,I331638,I331606,);
DFFARX1 I_19373 (I331918,I2595,I331638,I331627,);
nor I_19374 (I331980,I85376,I85370);
nor I_19375 (I331618,I331833,I331980);
or I_19376 (I332011,I85376,I85370);
nor I_19377 (I332028,I85367,I85361);
DFFARX1 I_19378 (I332028,I2595,I331638,I332054,);
not I_19379 (I332062,I332054);
nor I_19380 (I331624,I332062,I331867);
nand I_19381 (I332093,I332062,I331712);
not I_19382 (I332110,I85367);
nand I_19383 (I332127,I332110,I331816);
nand I_19384 (I332144,I332062,I332127);
nand I_19385 (I331615,I332144,I332093);
nand I_19386 (I331612,I332127,I332011);
not I_19387 (I332216,I2602);
DFFARX1 I_19388 (I163389,I2595,I332216,I332242,);
and I_19389 (I332250,I332242,I163377);
DFFARX1 I_19390 (I332250,I2595,I332216,I332199,);
DFFARX1 I_19391 (I163392,I2595,I332216,I332290,);
not I_19392 (I332298,I163383);
not I_19393 (I332315,I163374);
nand I_19394 (I332332,I332315,I332298);
nor I_19395 (I332187,I332290,I332332);
DFFARX1 I_19396 (I332332,I2595,I332216,I332372,);
not I_19397 (I332208,I332372);
not I_19398 (I332394,I163380);
nand I_19399 (I332411,I332315,I332394);
DFFARX1 I_19400 (I332411,I2595,I332216,I332437,);
not I_19401 (I332445,I332437);
not I_19402 (I332462,I163395);
nand I_19403 (I332479,I332462,I163398);
and I_19404 (I332496,I332298,I332479);
nor I_19405 (I332513,I332411,I332496);
DFFARX1 I_19406 (I332513,I2595,I332216,I332184,);
DFFARX1 I_19407 (I332496,I2595,I332216,I332205,);
nor I_19408 (I332558,I163395,I163374);
nor I_19409 (I332196,I332411,I332558);
or I_19410 (I332589,I163395,I163374);
nor I_19411 (I332606,I163386,I163377);
DFFARX1 I_19412 (I332606,I2595,I332216,I332632,);
not I_19413 (I332640,I332632);
nor I_19414 (I332202,I332640,I332445);
nand I_19415 (I332671,I332640,I332290);
not I_19416 (I332688,I163386);
nand I_19417 (I332705,I332688,I332394);
nand I_19418 (I332722,I332640,I332705);
nand I_19419 (I332193,I332722,I332671);
nand I_19420 (I332190,I332705,I332589);
not I_19421 (I332794,I2602);
DFFARX1 I_19422 (I103306,I2595,I332794,I332820,);
and I_19423 (I332828,I332820,I103291);
DFFARX1 I_19424 (I332828,I2595,I332794,I332777,);
DFFARX1 I_19425 (I103297,I2595,I332794,I332868,);
not I_19426 (I332876,I103279);
not I_19427 (I332893,I103300);
nand I_19428 (I332910,I332893,I332876);
nor I_19429 (I332765,I332868,I332910);
DFFARX1 I_19430 (I332910,I2595,I332794,I332950,);
not I_19431 (I332786,I332950);
not I_19432 (I332972,I103303);
nand I_19433 (I332989,I332893,I332972);
DFFARX1 I_19434 (I332989,I2595,I332794,I333015,);
not I_19435 (I333023,I333015);
not I_19436 (I333040,I103294);
nand I_19437 (I333057,I333040,I103282);
and I_19438 (I333074,I332876,I333057);
nor I_19439 (I333091,I332989,I333074);
DFFARX1 I_19440 (I333091,I2595,I332794,I332762,);
DFFARX1 I_19441 (I333074,I2595,I332794,I332783,);
nor I_19442 (I333136,I103294,I103288);
nor I_19443 (I332774,I332989,I333136);
or I_19444 (I333167,I103294,I103288);
nor I_19445 (I333184,I103285,I103279);
DFFARX1 I_19446 (I333184,I2595,I332794,I333210,);
not I_19447 (I333218,I333210);
nor I_19448 (I332780,I333218,I333023);
nand I_19449 (I333249,I333218,I332868);
not I_19450 (I333266,I103285);
nand I_19451 (I333283,I333266,I332972);
nand I_19452 (I333300,I333218,I333283);
nand I_19453 (I332771,I333300,I333249);
nand I_19454 (I332768,I333283,I333167);
not I_19455 (I333372,I2602);
DFFARX1 I_19456 (I72288,I2595,I333372,I333398,);
and I_19457 (I333406,I333398,I72291);
DFFARX1 I_19458 (I333406,I2595,I333372,I333355,);
DFFARX1 I_19459 (I72291,I2595,I333372,I333446,);
not I_19460 (I333454,I72306);
not I_19461 (I333471,I72312);
nand I_19462 (I333488,I333471,I333454);
nor I_19463 (I333343,I333446,I333488);
DFFARX1 I_19464 (I333488,I2595,I333372,I333528,);
not I_19465 (I333364,I333528);
not I_19466 (I333550,I72300);
nand I_19467 (I333567,I333471,I333550);
DFFARX1 I_19468 (I333567,I2595,I333372,I333593,);
not I_19469 (I333601,I333593);
not I_19470 (I333618,I72297);
nand I_19471 (I333635,I333618,I72294);
and I_19472 (I333652,I333454,I333635);
nor I_19473 (I333669,I333567,I333652);
DFFARX1 I_19474 (I333669,I2595,I333372,I333340,);
DFFARX1 I_19475 (I333652,I2595,I333372,I333361,);
nor I_19476 (I333714,I72297,I72288);
nor I_19477 (I333352,I333567,I333714);
or I_19478 (I333745,I72297,I72288);
nor I_19479 (I333762,I72303,I72309);
DFFARX1 I_19480 (I333762,I2595,I333372,I333788,);
not I_19481 (I333796,I333788);
nor I_19482 (I333358,I333796,I333601);
nand I_19483 (I333827,I333796,I333446);
not I_19484 (I333844,I72303);
nand I_19485 (I333861,I333844,I333550);
nand I_19486 (I333878,I333796,I333861);
nand I_19487 (I333349,I333878,I333827);
nand I_19488 (I333346,I333861,I333745);
not I_19489 (I333950,I2602);
DFFARX1 I_19490 (I39808,I2595,I333950,I333976,);
and I_19491 (I333984,I333976,I39784);
DFFARX1 I_19492 (I333984,I2595,I333950,I333933,);
DFFARX1 I_19493 (I39802,I2595,I333950,I334024,);
not I_19494 (I334032,I39790);
not I_19495 (I334049,I39787);
nand I_19496 (I334066,I334049,I334032);
nor I_19497 (I333921,I334024,I334066);
DFFARX1 I_19498 (I334066,I2595,I333950,I334106,);
not I_19499 (I333942,I334106);
not I_19500 (I334128,I39796);
nand I_19501 (I334145,I334049,I334128);
DFFARX1 I_19502 (I334145,I2595,I333950,I334171,);
not I_19503 (I334179,I334171);
not I_19504 (I334196,I39787);
nand I_19505 (I334213,I334196,I39805);
and I_19506 (I334230,I334032,I334213);
nor I_19507 (I334247,I334145,I334230);
DFFARX1 I_19508 (I334247,I2595,I333950,I333918,);
DFFARX1 I_19509 (I334230,I2595,I333950,I333939,);
nor I_19510 (I334292,I39787,I39799);
nor I_19511 (I333930,I334145,I334292);
or I_19512 (I334323,I39787,I39799);
nor I_19513 (I334340,I39793,I39784);
DFFARX1 I_19514 (I334340,I2595,I333950,I334366,);
not I_19515 (I334374,I334366);
nor I_19516 (I333936,I334374,I334179);
nand I_19517 (I334405,I334374,I334024);
not I_19518 (I334422,I39793);
nand I_19519 (I334439,I334422,I334128);
nand I_19520 (I334456,I334374,I334439);
nand I_19521 (I333927,I334456,I334405);
nand I_19522 (I333924,I334439,I334323);
not I_19523 (I334528,I2602);
DFFARX1 I_19524 (I132281,I2595,I334528,I334554,);
and I_19525 (I334562,I334554,I132296);
DFFARX1 I_19526 (I334562,I2595,I334528,I334511,);
DFFARX1 I_19527 (I132299,I2595,I334528,I334602,);
not I_19528 (I334610,I132293);
not I_19529 (I334627,I132308);
nand I_19530 (I334644,I334627,I334610);
nor I_19531 (I334499,I334602,I334644);
DFFARX1 I_19532 (I334644,I2595,I334528,I334684,);
not I_19533 (I334520,I334684);
not I_19534 (I334706,I132284);
nand I_19535 (I334723,I334627,I334706);
DFFARX1 I_19536 (I334723,I2595,I334528,I334749,);
not I_19537 (I334757,I334749);
not I_19538 (I334774,I132287);
nand I_19539 (I334791,I334774,I132281);
and I_19540 (I334808,I334610,I334791);
nor I_19541 (I334825,I334723,I334808);
DFFARX1 I_19542 (I334825,I2595,I334528,I334496,);
DFFARX1 I_19543 (I334808,I2595,I334528,I334517,);
nor I_19544 (I334870,I132287,I132290);
nor I_19545 (I334508,I334723,I334870);
or I_19546 (I334901,I132287,I132290);
nor I_19547 (I334918,I132305,I132302);
DFFARX1 I_19548 (I334918,I2595,I334528,I334944,);
not I_19549 (I334952,I334944);
nor I_19550 (I334514,I334952,I334757);
nand I_19551 (I334983,I334952,I334602);
not I_19552 (I335000,I132305);
nand I_19553 (I335017,I335000,I334706);
nand I_19554 (I335034,I334952,I335017);
nand I_19555 (I334505,I335034,I334983);
nand I_19556 (I334502,I335017,I334901);
not I_19557 (I335106,I2602);
DFFARX1 I_19558 (I199803,I2595,I335106,I335132,);
and I_19559 (I335140,I335132,I199791);
DFFARX1 I_19560 (I335140,I2595,I335106,I335089,);
DFFARX1 I_19561 (I199794,I2595,I335106,I335180,);
not I_19562 (I335188,I199788);
not I_19563 (I335205,I199812);
nand I_19564 (I335222,I335205,I335188);
nor I_19565 (I335077,I335180,I335222);
DFFARX1 I_19566 (I335222,I2595,I335106,I335262,);
not I_19567 (I335098,I335262);
not I_19568 (I335284,I199800);
nand I_19569 (I335301,I335205,I335284);
DFFARX1 I_19570 (I335301,I2595,I335106,I335327,);
not I_19571 (I335335,I335327);
not I_19572 (I335352,I199809);
nand I_19573 (I335369,I335352,I199806);
and I_19574 (I335386,I335188,I335369);
nor I_19575 (I335403,I335301,I335386);
DFFARX1 I_19576 (I335403,I2595,I335106,I335074,);
DFFARX1 I_19577 (I335386,I2595,I335106,I335095,);
nor I_19578 (I335448,I199809,I199797);
nor I_19579 (I335086,I335301,I335448);
or I_19580 (I335479,I199809,I199797);
nor I_19581 (I335496,I199788,I199791);
DFFARX1 I_19582 (I335496,I2595,I335106,I335522,);
not I_19583 (I335530,I335522);
nor I_19584 (I335092,I335530,I335335);
nand I_19585 (I335561,I335530,I335180);
not I_19586 (I335578,I199788);
nand I_19587 (I335595,I335578,I335284);
nand I_19588 (I335612,I335530,I335595);
nand I_19589 (I335083,I335612,I335561);
nand I_19590 (I335080,I335595,I335479);
not I_19591 (I335684,I2602);
DFFARX1 I_19592 (I28741,I2595,I335684,I335710,);
and I_19593 (I335718,I335710,I28717);
DFFARX1 I_19594 (I335718,I2595,I335684,I335667,);
DFFARX1 I_19595 (I28735,I2595,I335684,I335758,);
not I_19596 (I335766,I28723);
not I_19597 (I335783,I28720);
nand I_19598 (I335800,I335783,I335766);
nor I_19599 (I335655,I335758,I335800);
DFFARX1 I_19600 (I335800,I2595,I335684,I335840,);
not I_19601 (I335676,I335840);
not I_19602 (I335862,I28729);
nand I_19603 (I335879,I335783,I335862);
DFFARX1 I_19604 (I335879,I2595,I335684,I335905,);
not I_19605 (I335913,I335905);
not I_19606 (I335930,I28720);
nand I_19607 (I335947,I335930,I28738);
and I_19608 (I335964,I335766,I335947);
nor I_19609 (I335981,I335879,I335964);
DFFARX1 I_19610 (I335981,I2595,I335684,I335652,);
DFFARX1 I_19611 (I335964,I2595,I335684,I335673,);
nor I_19612 (I336026,I28720,I28732);
nor I_19613 (I335664,I335879,I336026);
or I_19614 (I336057,I28720,I28732);
nor I_19615 (I336074,I28726,I28717);
DFFARX1 I_19616 (I336074,I2595,I335684,I336100,);
not I_19617 (I336108,I336100);
nor I_19618 (I335670,I336108,I335913);
nand I_19619 (I336139,I336108,I335758);
not I_19620 (I336156,I28726);
nand I_19621 (I336173,I336156,I335862);
nand I_19622 (I336190,I336108,I336173);
nand I_19623 (I335661,I336190,I336139);
nand I_19624 (I335658,I336173,I336057);
not I_19625 (I336262,I2602);
DFFARX1 I_19626 (I49083,I2595,I336262,I336288,);
and I_19627 (I336296,I336288,I49086);
DFFARX1 I_19628 (I336296,I2595,I336262,I336245,);
DFFARX1 I_19629 (I49086,I2595,I336262,I336336,);
not I_19630 (I336344,I49101);
not I_19631 (I336361,I49107);
nand I_19632 (I336378,I336361,I336344);
nor I_19633 (I336233,I336336,I336378);
DFFARX1 I_19634 (I336378,I2595,I336262,I336418,);
not I_19635 (I336254,I336418);
not I_19636 (I336440,I49095);
nand I_19637 (I336457,I336361,I336440);
DFFARX1 I_19638 (I336457,I2595,I336262,I336483,);
not I_19639 (I336491,I336483);
not I_19640 (I336508,I49092);
nand I_19641 (I336525,I336508,I49089);
and I_19642 (I336542,I336344,I336525);
nor I_19643 (I336559,I336457,I336542);
DFFARX1 I_19644 (I336559,I2595,I336262,I336230,);
DFFARX1 I_19645 (I336542,I2595,I336262,I336251,);
nor I_19646 (I336604,I49092,I49083);
nor I_19647 (I336242,I336457,I336604);
or I_19648 (I336635,I49092,I49083);
nor I_19649 (I336652,I49098,I49104);
DFFARX1 I_19650 (I336652,I2595,I336262,I336678,);
not I_19651 (I336686,I336678);
nor I_19652 (I336248,I336686,I336491);
nand I_19653 (I336717,I336686,I336336);
not I_19654 (I336734,I49098);
nand I_19655 (I336751,I336734,I336440);
nand I_19656 (I336768,I336686,I336751);
nand I_19657 (I336239,I336768,I336717);
nand I_19658 (I336236,I336751,I336635);
not I_19659 (I336840,I2602);
DFFARX1 I_19660 (I256387,I2595,I336840,I336866,);
and I_19661 (I336874,I336866,I256381);
DFFARX1 I_19662 (I336874,I2595,I336840,I336823,);
DFFARX1 I_19663 (I256399,I2595,I336840,I336914,);
not I_19664 (I336922,I256390);
not I_19665 (I336939,I256402);
nand I_19666 (I336956,I336939,I336922);
nor I_19667 (I336811,I336914,I336956);
DFFARX1 I_19668 (I336956,I2595,I336840,I336996,);
not I_19669 (I336832,I336996);
not I_19670 (I337018,I256408);
nand I_19671 (I337035,I336939,I337018);
DFFARX1 I_19672 (I337035,I2595,I336840,I337061,);
not I_19673 (I337069,I337061);
not I_19674 (I337086,I256384);
nand I_19675 (I337103,I337086,I256405);
and I_19676 (I337120,I336922,I337103);
nor I_19677 (I337137,I337035,I337120);
DFFARX1 I_19678 (I337137,I2595,I336840,I336808,);
DFFARX1 I_19679 (I337120,I2595,I336840,I336829,);
nor I_19680 (I337182,I256384,I256396);
nor I_19681 (I336820,I337035,I337182);
or I_19682 (I337213,I256384,I256396);
nor I_19683 (I337230,I256381,I256393);
DFFARX1 I_19684 (I337230,I2595,I336840,I337256,);
not I_19685 (I337264,I337256);
nor I_19686 (I336826,I337264,I337069);
nand I_19687 (I337295,I337264,I336914);
not I_19688 (I337312,I256381);
nand I_19689 (I337329,I337312,I337018);
nand I_19690 (I337346,I337264,I337329);
nand I_19691 (I336817,I337346,I337295);
nand I_19692 (I336814,I337329,I337213);
not I_19693 (I337418,I2602);
DFFARX1 I_19694 (I163967,I2595,I337418,I337444,);
and I_19695 (I337452,I337444,I163955);
DFFARX1 I_19696 (I337452,I2595,I337418,I337401,);
DFFARX1 I_19697 (I163970,I2595,I337418,I337492,);
not I_19698 (I337500,I163961);
not I_19699 (I337517,I163952);
nand I_19700 (I337534,I337517,I337500);
nor I_19701 (I337389,I337492,I337534);
DFFARX1 I_19702 (I337534,I2595,I337418,I337574,);
not I_19703 (I337410,I337574);
not I_19704 (I337596,I163958);
nand I_19705 (I337613,I337517,I337596);
DFFARX1 I_19706 (I337613,I2595,I337418,I337639,);
not I_19707 (I337647,I337639);
not I_19708 (I337664,I163973);
nand I_19709 (I337681,I337664,I163976);
and I_19710 (I337698,I337500,I337681);
nor I_19711 (I337715,I337613,I337698);
DFFARX1 I_19712 (I337715,I2595,I337418,I337386,);
DFFARX1 I_19713 (I337698,I2595,I337418,I337407,);
nor I_19714 (I337760,I163973,I163952);
nor I_19715 (I337398,I337613,I337760);
or I_19716 (I337791,I163973,I163952);
nor I_19717 (I337808,I163964,I163955);
DFFARX1 I_19718 (I337808,I2595,I337418,I337834,);
not I_19719 (I337842,I337834);
nor I_19720 (I337404,I337842,I337647);
nand I_19721 (I337873,I337842,I337492);
not I_19722 (I337890,I163964);
nand I_19723 (I337907,I337890,I337596);
nand I_19724 (I337924,I337842,I337907);
nand I_19725 (I337395,I337924,I337873);
nand I_19726 (I337392,I337907,I337791);
not I_19727 (I337996,I2602);
DFFARX1 I_19728 (I102252,I2595,I337996,I338022,);
and I_19729 (I338030,I338022,I102237);
DFFARX1 I_19730 (I338030,I2595,I337996,I337979,);
DFFARX1 I_19731 (I102243,I2595,I337996,I338070,);
not I_19732 (I338078,I102225);
not I_19733 (I338095,I102246);
nand I_19734 (I338112,I338095,I338078);
nor I_19735 (I337967,I338070,I338112);
DFFARX1 I_19736 (I338112,I2595,I337996,I338152,);
not I_19737 (I337988,I338152);
not I_19738 (I338174,I102249);
nand I_19739 (I338191,I338095,I338174);
DFFARX1 I_19740 (I338191,I2595,I337996,I338217,);
not I_19741 (I338225,I338217);
not I_19742 (I338242,I102240);
nand I_19743 (I338259,I338242,I102228);
and I_19744 (I338276,I338078,I338259);
nor I_19745 (I338293,I338191,I338276);
DFFARX1 I_19746 (I338293,I2595,I337996,I337964,);
DFFARX1 I_19747 (I338276,I2595,I337996,I337985,);
nor I_19748 (I338338,I102240,I102234);
nor I_19749 (I337976,I338191,I338338);
or I_19750 (I338369,I102240,I102234);
nor I_19751 (I338386,I102231,I102225);
DFFARX1 I_19752 (I338386,I2595,I337996,I338412,);
not I_19753 (I338420,I338412);
nor I_19754 (I337982,I338420,I338225);
nand I_19755 (I338451,I338420,I338070);
not I_19756 (I338468,I102231);
nand I_19757 (I338485,I338468,I338174);
nand I_19758 (I338502,I338420,I338485);
nand I_19759 (I337973,I338502,I338451);
nand I_19760 (I337970,I338485,I338369);
not I_19761 (I338574,I2602);
DFFARX1 I_19762 (I120313,I2595,I338574,I338600,);
and I_19763 (I338608,I338600,I120328);
DFFARX1 I_19764 (I338608,I2595,I338574,I338557,);
DFFARX1 I_19765 (I120331,I2595,I338574,I338648,);
not I_19766 (I338656,I120325);
not I_19767 (I338673,I120340);
nand I_19768 (I338690,I338673,I338656);
nor I_19769 (I338545,I338648,I338690);
DFFARX1 I_19770 (I338690,I2595,I338574,I338730,);
not I_19771 (I338566,I338730);
not I_19772 (I338752,I120316);
nand I_19773 (I338769,I338673,I338752);
DFFARX1 I_19774 (I338769,I2595,I338574,I338795,);
not I_19775 (I338803,I338795);
not I_19776 (I338820,I120319);
nand I_19777 (I338837,I338820,I120313);
and I_19778 (I338854,I338656,I338837);
nor I_19779 (I338871,I338769,I338854);
DFFARX1 I_19780 (I338871,I2595,I338574,I338542,);
DFFARX1 I_19781 (I338854,I2595,I338574,I338563,);
nor I_19782 (I338916,I120319,I120322);
nor I_19783 (I338554,I338769,I338916);
or I_19784 (I338947,I120319,I120322);
nor I_19785 (I338964,I120337,I120334);
DFFARX1 I_19786 (I338964,I2595,I338574,I338990,);
not I_19787 (I338998,I338990);
nor I_19788 (I338560,I338998,I338803);
nand I_19789 (I339029,I338998,I338648);
not I_19790 (I339046,I120337);
nand I_19791 (I339063,I339046,I338752);
nand I_19792 (I339080,I338998,I339063);
nand I_19793 (I338551,I339080,I339029);
nand I_19794 (I338548,I339063,I338947);
not I_19795 (I339152,I2602);
DFFARX1 I_19796 (I246184,I2595,I339152,I339178,);
and I_19797 (I339186,I339178,I246190);
DFFARX1 I_19798 (I339186,I2595,I339152,I339135,);
DFFARX1 I_19799 (I246196,I2595,I339152,I339226,);
not I_19800 (I339234,I246181);
not I_19801 (I339251,I246181);
nand I_19802 (I339268,I339251,I339234);
nor I_19803 (I339123,I339226,I339268);
DFFARX1 I_19804 (I339268,I2595,I339152,I339308,);
not I_19805 (I339144,I339308);
not I_19806 (I339330,I246199);
nand I_19807 (I339347,I339251,I339330);
DFFARX1 I_19808 (I339347,I2595,I339152,I339373,);
not I_19809 (I339381,I339373);
not I_19810 (I339398,I246193);
nand I_19811 (I339415,I339398,I246184);
and I_19812 (I339432,I339234,I339415);
nor I_19813 (I339449,I339347,I339432);
DFFARX1 I_19814 (I339449,I2595,I339152,I339120,);
DFFARX1 I_19815 (I339432,I2595,I339152,I339141,);
nor I_19816 (I339494,I246193,I246202);
nor I_19817 (I339132,I339347,I339494);
or I_19818 (I339525,I246193,I246202);
nor I_19819 (I339542,I246187,I246187);
DFFARX1 I_19820 (I339542,I2595,I339152,I339568,);
not I_19821 (I339576,I339568);
nor I_19822 (I339138,I339576,I339381);
nand I_19823 (I339607,I339576,I339226);
not I_19824 (I339624,I246187);
nand I_19825 (I339641,I339624,I339330);
nand I_19826 (I339658,I339576,I339641);
nand I_19827 (I339129,I339658,I339607);
nand I_19828 (I339126,I339641,I339525);
not I_19829 (I339730,I2602);
DFFARX1 I_19830 (I284811,I2595,I339730,I339756,);
and I_19831 (I339764,I339756,I284805);
DFFARX1 I_19832 (I339764,I2595,I339730,I339713,);
DFFARX1 I_19833 (I284823,I2595,I339730,I339804,);
not I_19834 (I339812,I284814);
not I_19835 (I339829,I284826);
nand I_19836 (I339846,I339829,I339812);
nor I_19837 (I339701,I339804,I339846);
DFFARX1 I_19838 (I339846,I2595,I339730,I339886,);
not I_19839 (I339722,I339886);
not I_19840 (I339908,I284832);
nand I_19841 (I339925,I339829,I339908);
DFFARX1 I_19842 (I339925,I2595,I339730,I339951,);
not I_19843 (I339959,I339951);
not I_19844 (I339976,I284808);
nand I_19845 (I339993,I339976,I284829);
and I_19846 (I340010,I339812,I339993);
nor I_19847 (I340027,I339925,I340010);
DFFARX1 I_19848 (I340027,I2595,I339730,I339698,);
DFFARX1 I_19849 (I340010,I2595,I339730,I339719,);
nor I_19850 (I340072,I284808,I284820);
nor I_19851 (I339710,I339925,I340072);
or I_19852 (I340103,I284808,I284820);
nor I_19853 (I340120,I284805,I284817);
DFFARX1 I_19854 (I340120,I2595,I339730,I340146,);
not I_19855 (I340154,I340146);
nor I_19856 (I339716,I340154,I339959);
nand I_19857 (I340185,I340154,I339804);
not I_19858 (I340202,I284805);
nand I_19859 (I340219,I340202,I339908);
nand I_19860 (I340236,I340154,I340219);
nand I_19861 (I339707,I340236,I340185);
nand I_19862 (I339704,I340219,I340103);
not I_19863 (I340308,I2602);
DFFARX1 I_19864 (I378910,I2595,I340308,I340334,);
and I_19865 (I340342,I340334,I378892);
DFFARX1 I_19866 (I340342,I2595,I340308,I340291,);
DFFARX1 I_19867 (I378883,I2595,I340308,I340382,);
not I_19868 (I340390,I378898);
not I_19869 (I340407,I378886);
nand I_19870 (I340424,I340407,I340390);
nor I_19871 (I340279,I340382,I340424);
DFFARX1 I_19872 (I340424,I2595,I340308,I340464,);
not I_19873 (I340300,I340464);
not I_19874 (I340486,I378895);
nand I_19875 (I340503,I340407,I340486);
DFFARX1 I_19876 (I340503,I2595,I340308,I340529,);
not I_19877 (I340537,I340529);
not I_19878 (I340554,I378904);
nand I_19879 (I340571,I340554,I378883);
and I_19880 (I340588,I340390,I340571);
nor I_19881 (I340605,I340503,I340588);
DFFARX1 I_19882 (I340605,I2595,I340308,I340276,);
DFFARX1 I_19883 (I340588,I2595,I340308,I340297,);
nor I_19884 (I340650,I378904,I378907);
nor I_19885 (I340288,I340503,I340650);
or I_19886 (I340681,I378904,I378907);
nor I_19887 (I340698,I378901,I378889);
DFFARX1 I_19888 (I340698,I2595,I340308,I340724,);
not I_19889 (I340732,I340724);
nor I_19890 (I340294,I340732,I340537);
nand I_19891 (I340763,I340732,I340382);
not I_19892 (I340780,I378901);
nand I_19893 (I340797,I340780,I340486);
nand I_19894 (I340814,I340732,I340797);
nand I_19895 (I340285,I340814,I340763);
nand I_19896 (I340282,I340797,I340681);
not I_19897 (I340886,I2602);
DFFARX1 I_19898 (I82226,I2595,I340886,I340912,);
and I_19899 (I340920,I340912,I82211);
DFFARX1 I_19900 (I340920,I2595,I340886,I340869,);
DFFARX1 I_19901 (I82217,I2595,I340886,I340960,);
not I_19902 (I340968,I82199);
not I_19903 (I340985,I82220);
nand I_19904 (I341002,I340985,I340968);
nor I_19905 (I340857,I340960,I341002);
DFFARX1 I_19906 (I341002,I2595,I340886,I341042,);
not I_19907 (I340878,I341042);
not I_19908 (I341064,I82223);
nand I_19909 (I341081,I340985,I341064);
DFFARX1 I_19910 (I341081,I2595,I340886,I341107,);
not I_19911 (I341115,I341107);
not I_19912 (I341132,I82214);
nand I_19913 (I341149,I341132,I82202);
and I_19914 (I341166,I340968,I341149);
nor I_19915 (I341183,I341081,I341166);
DFFARX1 I_19916 (I341183,I2595,I340886,I340854,);
DFFARX1 I_19917 (I341166,I2595,I340886,I340875,);
nor I_19918 (I341228,I82214,I82208);
nor I_19919 (I340866,I341081,I341228);
or I_19920 (I341259,I82214,I82208);
nor I_19921 (I341276,I82205,I82199);
DFFARX1 I_19922 (I341276,I2595,I340886,I341302,);
not I_19923 (I341310,I341302);
nor I_19924 (I340872,I341310,I341115);
nand I_19925 (I341341,I341310,I340960);
not I_19926 (I341358,I82205);
nand I_19927 (I341375,I341358,I341064);
nand I_19928 (I341392,I341310,I341375);
nand I_19929 (I340863,I341392,I341341);
nand I_19930 (I340860,I341375,I341259);
not I_19931 (I341464,I2602);
DFFARX1 I_19932 (I305038,I2595,I341464,I341490,);
and I_19933 (I341498,I341490,I305035);
DFFARX1 I_19934 (I341498,I2595,I341464,I341447,);
DFFARX1 I_19935 (I305041,I2595,I341464,I341538,);
not I_19936 (I341546,I305044);
not I_19937 (I341563,I305038);
nand I_19938 (I341580,I341563,I341546);
nor I_19939 (I341435,I341538,I341580);
DFFARX1 I_19940 (I341580,I2595,I341464,I341620,);
not I_19941 (I341456,I341620);
not I_19942 (I341642,I305053);
nand I_19943 (I341659,I341563,I341642);
DFFARX1 I_19944 (I341659,I2595,I341464,I341685,);
not I_19945 (I341693,I341685);
not I_19946 (I341710,I305050);
nand I_19947 (I341727,I341710,I305056);
and I_19948 (I341744,I341546,I341727);
nor I_19949 (I341761,I341659,I341744);
DFFARX1 I_19950 (I341761,I2595,I341464,I341432,);
DFFARX1 I_19951 (I341744,I2595,I341464,I341453,);
nor I_19952 (I341806,I305050,I305035);
nor I_19953 (I341444,I341659,I341806);
or I_19954 (I341837,I305050,I305035);
nor I_19955 (I341854,I305047,I305041);
DFFARX1 I_19956 (I341854,I2595,I341464,I341880,);
not I_19957 (I341888,I341880);
nor I_19958 (I341450,I341888,I341693);
nand I_19959 (I341919,I341888,I341538);
not I_19960 (I341936,I305047);
nand I_19961 (I341953,I341936,I341642);
nand I_19962 (I341970,I341888,I341953);
nand I_19963 (I341441,I341970,I341919);
nand I_19964 (I341438,I341953,I341837);
not I_19965 (I342042,I2602);
DFFARX1 I_19966 (I112265,I2595,I342042,I342068,);
and I_19967 (I342076,I342068,I112250);
DFFARX1 I_19968 (I342076,I2595,I342042,I342025,);
DFFARX1 I_19969 (I112256,I2595,I342042,I342116,);
not I_19970 (I342124,I112238);
not I_19971 (I342141,I112259);
nand I_19972 (I342158,I342141,I342124);
nor I_19973 (I342013,I342116,I342158);
DFFARX1 I_19974 (I342158,I2595,I342042,I342198,);
not I_19975 (I342034,I342198);
not I_19976 (I342220,I112262);
nand I_19977 (I342237,I342141,I342220);
DFFARX1 I_19978 (I342237,I2595,I342042,I342263,);
not I_19979 (I342271,I342263);
not I_19980 (I342288,I112253);
nand I_19981 (I342305,I342288,I112241);
and I_19982 (I342322,I342124,I342305);
nor I_19983 (I342339,I342237,I342322);
DFFARX1 I_19984 (I342339,I2595,I342042,I342010,);
DFFARX1 I_19985 (I342322,I2595,I342042,I342031,);
nor I_19986 (I342384,I112253,I112247);
nor I_19987 (I342022,I342237,I342384);
or I_19988 (I342415,I112253,I112247);
nor I_19989 (I342432,I112244,I112238);
DFFARX1 I_19990 (I342432,I2595,I342042,I342458,);
not I_19991 (I342466,I342458);
nor I_19992 (I342028,I342466,I342271);
nand I_19993 (I342497,I342466,I342116);
not I_19994 (I342514,I112244);
nand I_19995 (I342531,I342514,I342220);
nand I_19996 (I342548,I342466,I342531);
nand I_19997 (I342019,I342548,I342497);
nand I_19998 (I342016,I342531,I342415);
not I_19999 (I342620,I2602);
DFFARX1 I_20000 (I161077,I2595,I342620,I342646,);
and I_20001 (I342654,I342646,I161065);
DFFARX1 I_20002 (I342654,I2595,I342620,I342603,);
DFFARX1 I_20003 (I161080,I2595,I342620,I342694,);
not I_20004 (I342702,I161071);
not I_20005 (I342719,I161062);
nand I_20006 (I342736,I342719,I342702);
nor I_20007 (I342591,I342694,I342736);
DFFARX1 I_20008 (I342736,I2595,I342620,I342776,);
not I_20009 (I342612,I342776);
not I_20010 (I342798,I161068);
nand I_20011 (I342815,I342719,I342798);
DFFARX1 I_20012 (I342815,I2595,I342620,I342841,);
not I_20013 (I342849,I342841);
not I_20014 (I342866,I161083);
nand I_20015 (I342883,I342866,I161086);
and I_20016 (I342900,I342702,I342883);
nor I_20017 (I342917,I342815,I342900);
DFFARX1 I_20018 (I342917,I2595,I342620,I342588,);
DFFARX1 I_20019 (I342900,I2595,I342620,I342609,);
nor I_20020 (I342962,I161083,I161062);
nor I_20021 (I342600,I342815,I342962);
or I_20022 (I342993,I161083,I161062);
nor I_20023 (I343010,I161074,I161065);
DFFARX1 I_20024 (I343010,I2595,I342620,I343036,);
not I_20025 (I343044,I343036);
nor I_20026 (I342606,I343044,I342849);
nand I_20027 (I343075,I343044,I342694);
not I_20028 (I343092,I161074);
nand I_20029 (I343109,I343092,I342798);
nand I_20030 (I343126,I343044,I343109);
nand I_20031 (I342597,I343126,I343075);
nand I_20032 (I342594,I343109,I342993);
not I_20033 (I343198,I2602);
DFFARX1 I_20034 (I316024,I2595,I343198,I343224,);
nand I_20035 (I343232,I343224,I316003);
DFFARX1 I_20036 (I316000,I2595,I343198,I343258,);
DFFARX1 I_20037 (I343258,I2595,I343198,I343275,);
not I_20038 (I343190,I343275);
not I_20039 (I343297,I316012);
nor I_20040 (I343314,I316012,I316021);
not I_20041 (I343331,I316009);
nand I_20042 (I343348,I343297,I343331);
nor I_20043 (I343365,I316009,I316012);
and I_20044 (I343169,I343365,I343232);
not I_20045 (I343396,I316018);
nand I_20046 (I343413,I343396,I316015);
nor I_20047 (I343430,I316018,I316000);
not I_20048 (I343447,I343430);
nand I_20049 (I343172,I343314,I343447);
DFFARX1 I_20050 (I343430,I2595,I343198,I343187,);
nor I_20051 (I343492,I316003,I316009);
nor I_20052 (I343509,I343492,I316021);
and I_20053 (I343526,I343509,I343413);
DFFARX1 I_20054 (I343526,I2595,I343198,I343184,);
nor I_20055 (I343181,I343492,I343348);
or I_20056 (I343178,I343430,I343492);
nor I_20057 (I343585,I316003,I316006);
DFFARX1 I_20058 (I343585,I2595,I343198,I343611,);
not I_20059 (I343619,I343611);
nand I_20060 (I343636,I343619,I343297);
nor I_20061 (I343653,I343636,I316021);
DFFARX1 I_20062 (I343653,I2595,I343198,I343166,);
nor I_20063 (I343684,I343619,I343348);
nor I_20064 (I343175,I343492,I343684);
not I_20065 (I343742,I2602);
DFFARX1 I_20066 (I311400,I2595,I343742,I343768,);
nand I_20067 (I343776,I343768,I311379);
DFFARX1 I_20068 (I311376,I2595,I343742,I343802,);
DFFARX1 I_20069 (I343802,I2595,I343742,I343819,);
not I_20070 (I343734,I343819);
not I_20071 (I343841,I311388);
nor I_20072 (I343858,I311388,I311397);
not I_20073 (I343875,I311385);
nand I_20074 (I343892,I343841,I343875);
nor I_20075 (I343909,I311385,I311388);
and I_20076 (I343713,I343909,I343776);
not I_20077 (I343940,I311394);
nand I_20078 (I343957,I343940,I311391);
nor I_20079 (I343974,I311394,I311376);
not I_20080 (I343991,I343974);
nand I_20081 (I343716,I343858,I343991);
DFFARX1 I_20082 (I343974,I2595,I343742,I343731,);
nor I_20083 (I344036,I311379,I311385);
nor I_20084 (I344053,I344036,I311397);
and I_20085 (I344070,I344053,I343957);
DFFARX1 I_20086 (I344070,I2595,I343742,I343728,);
nor I_20087 (I343725,I344036,I343892);
or I_20088 (I343722,I343974,I344036);
nor I_20089 (I344129,I311379,I311382);
DFFARX1 I_20090 (I344129,I2595,I343742,I344155,);
not I_20091 (I344163,I344155);
nand I_20092 (I344180,I344163,I343841);
nor I_20093 (I344197,I344180,I311397);
DFFARX1 I_20094 (I344197,I2595,I343742,I343710,);
nor I_20095 (I344228,I344163,I343892);
nor I_20096 (I343719,I344036,I344228);
not I_20097 (I344286,I2602);
DFFARX1 I_20098 (I86427,I2595,I344286,I344312,);
nand I_20099 (I344320,I344312,I86430);
DFFARX1 I_20100 (I86424,I2595,I344286,I344346,);
DFFARX1 I_20101 (I344346,I2595,I344286,I344363,);
not I_20102 (I344278,I344363);
not I_20103 (I344385,I86433);
nor I_20104 (I344402,I86433,I86418);
not I_20105 (I344419,I86442);
nand I_20106 (I344436,I344385,I344419);
nor I_20107 (I344453,I86442,I86433);
and I_20108 (I344257,I344453,I344320);
not I_20109 (I344484,I86421);
nand I_20110 (I344501,I344484,I86439);
nor I_20111 (I344518,I86421,I86415);
not I_20112 (I344535,I344518);
nand I_20113 (I344260,I344402,I344535);
DFFARX1 I_20114 (I344518,I2595,I344286,I344275,);
nor I_20115 (I344580,I86436,I86442);
nor I_20116 (I344597,I344580,I86418);
and I_20117 (I344614,I344597,I344501);
DFFARX1 I_20118 (I344614,I2595,I344286,I344272,);
nor I_20119 (I344269,I344580,I344436);
or I_20120 (I344266,I344518,I344580);
nor I_20121 (I344673,I86436,I86415);
DFFARX1 I_20122 (I344673,I2595,I344286,I344699,);
not I_20123 (I344707,I344699);
nand I_20124 (I344724,I344707,I344385);
nor I_20125 (I344741,I344724,I86418);
DFFARX1 I_20126 (I344741,I2595,I344286,I344254,);
nor I_20127 (I344772,I344707,I344436);
nor I_20128 (I344263,I344580,I344772);
not I_20129 (I344830,I2602);
DFFARX1 I_20130 (I2068,I2595,I344830,I344856,);
nand I_20131 (I344864,I344856,I1980);
DFFARX1 I_20132 (I1908,I2595,I344830,I344890,);
DFFARX1 I_20133 (I344890,I2595,I344830,I344907,);
not I_20134 (I344822,I344907);
not I_20135 (I344929,I2236);
nor I_20136 (I344946,I2236,I1716);
not I_20137 (I344963,I2372);
nand I_20138 (I344980,I344929,I344963);
nor I_20139 (I344997,I2372,I2236);
and I_20140 (I344801,I344997,I344864);
not I_20141 (I345028,I2524);
nand I_20142 (I345045,I345028,I1988);
nor I_20143 (I345062,I2524,I2492);
not I_20144 (I345079,I345062);
nand I_20145 (I344804,I344946,I345079);
DFFARX1 I_20146 (I345062,I2595,I344830,I344819,);
nor I_20147 (I345124,I1724,I2372);
nor I_20148 (I345141,I345124,I1716);
and I_20149 (I345158,I345141,I345045);
DFFARX1 I_20150 (I345158,I2595,I344830,I344816,);
nor I_20151 (I344813,I345124,I344980);
or I_20152 (I344810,I345062,I345124);
nor I_20153 (I345217,I1724,I2572);
DFFARX1 I_20154 (I345217,I2595,I344830,I345243,);
not I_20155 (I345251,I345243);
nand I_20156 (I345268,I345251,I344929);
nor I_20157 (I345285,I345268,I1716);
DFFARX1 I_20158 (I345285,I2595,I344830,I344798,);
nor I_20159 (I345316,I345251,I344980);
nor I_20160 (I344807,I345124,I345316);
not I_20161 (I345374,I2602);
DFFARX1 I_20162 (I12916,I2595,I345374,I345400,);
nand I_20163 (I345408,I345400,I12910);
DFFARX1 I_20164 (I12931,I2595,I345374,I345434,);
DFFARX1 I_20165 (I345434,I2595,I345374,I345451,);
not I_20166 (I345366,I345451);
not I_20167 (I345473,I12919);
nor I_20168 (I345490,I12919,I12928);
not I_20169 (I345507,I12907);
nand I_20170 (I345524,I345473,I345507);
nor I_20171 (I345541,I12907,I12919);
and I_20172 (I345345,I345541,I345408);
not I_20173 (I345572,I12925);
nand I_20174 (I345589,I345572,I12913);
nor I_20175 (I345606,I12925,I12907);
not I_20176 (I345623,I345606);
nand I_20177 (I345348,I345490,I345623);
DFFARX1 I_20178 (I345606,I2595,I345374,I345363,);
nor I_20179 (I345668,I12910,I12907);
nor I_20180 (I345685,I345668,I12928);
and I_20181 (I345702,I345685,I345589);
DFFARX1 I_20182 (I345702,I2595,I345374,I345360,);
nor I_20183 (I345357,I345668,I345524);
or I_20184 (I345354,I345606,I345668);
nor I_20185 (I345761,I12910,I12922);
DFFARX1 I_20186 (I345761,I2595,I345374,I345787,);
not I_20187 (I345795,I345787);
nand I_20188 (I345812,I345795,I345473);
nor I_20189 (I345829,I345812,I12928);
DFFARX1 I_20190 (I345829,I2595,I345374,I345342,);
nor I_20191 (I345860,I345795,I345524);
nor I_20192 (I345351,I345668,I345860);
not I_20193 (I345918,I2602);
DFFARX1 I_20194 (I161661,I2595,I345918,I345944,);
nand I_20195 (I345952,I345944,I161649);
DFFARX1 I_20196 (I161655,I2595,I345918,I345978,);
DFFARX1 I_20197 (I345978,I2595,I345918,I345995,);
not I_20198 (I345910,I345995);
not I_20199 (I346017,I161640);
nor I_20200 (I346034,I161640,I161652);
not I_20201 (I346051,I161643);
nand I_20202 (I346068,I346017,I346051);
nor I_20203 (I346085,I161643,I161640);
and I_20204 (I345889,I346085,I345952);
not I_20205 (I346116,I161658);
nand I_20206 (I346133,I346116,I161640);
nor I_20207 (I346150,I161658,I161664);
not I_20208 (I346167,I346150);
nand I_20209 (I345892,I346034,I346167);
DFFARX1 I_20210 (I346150,I2595,I345918,I345907,);
nor I_20211 (I346212,I161646,I161643);
nor I_20212 (I346229,I346212,I161652);
and I_20213 (I346246,I346229,I346133);
DFFARX1 I_20214 (I346246,I2595,I345918,I345904,);
nor I_20215 (I345901,I346212,I346068);
or I_20216 (I345898,I346150,I346212);
nor I_20217 (I346305,I161646,I161643);
DFFARX1 I_20218 (I346305,I2595,I345918,I346331,);
not I_20219 (I346339,I346331);
nand I_20220 (I346356,I346339,I346017);
nor I_20221 (I346373,I346356,I161652);
DFFARX1 I_20222 (I346373,I2595,I345918,I345886,);
nor I_20223 (I346404,I346339,I346068);
nor I_20224 (I345895,I346212,I346404);
not I_20225 (I346462,I2602);
DFFARX1 I_20226 (I78247,I2595,I346462,I346488,);
nand I_20227 (I346496,I346488,I78262);
DFFARX1 I_20228 (I78259,I2595,I346462,I346522,);
DFFARX1 I_20229 (I346522,I2595,I346462,I346539,);
not I_20230 (I346454,I346539);
not I_20231 (I346561,I78238);
nor I_20232 (I346578,I78238,I78244);
not I_20233 (I346595,I78250);
nand I_20234 (I346612,I346561,I346595);
nor I_20235 (I346629,I78250,I78238);
and I_20236 (I346433,I346629,I346496);
not I_20237 (I346660,I78256);
nand I_20238 (I346677,I346660,I78238);
nor I_20239 (I346694,I78256,I78241);
not I_20240 (I346711,I346694);
nand I_20241 (I346436,I346578,I346711);
DFFARX1 I_20242 (I346694,I2595,I346462,I346451,);
nor I_20243 (I346756,I78241,I78250);
nor I_20244 (I346773,I346756,I78244);
and I_20245 (I346790,I346773,I346677);
DFFARX1 I_20246 (I346790,I2595,I346462,I346448,);
nor I_20247 (I346445,I346756,I346612);
or I_20248 (I346442,I346694,I346756);
nor I_20249 (I346849,I78241,I78253);
DFFARX1 I_20250 (I346849,I2595,I346462,I346875,);
not I_20251 (I346883,I346875);
nand I_20252 (I346900,I346883,I346561);
nor I_20253 (I346917,I346900,I78244);
DFFARX1 I_20254 (I346917,I2595,I346462,I346430,);
nor I_20255 (I346948,I346883,I346612);
nor I_20256 (I346439,I346756,I346948);
not I_20257 (I347006,I2602);
DFFARX1 I_20258 (I196901,I2595,I347006,I347032,);
nand I_20259 (I347040,I347032,I196916);
DFFARX1 I_20260 (I196910,I2595,I347006,I347066,);
DFFARX1 I_20261 (I347066,I2595,I347006,I347083,);
not I_20262 (I346998,I347083);
not I_20263 (I347105,I196913);
nor I_20264 (I347122,I196913,I196919);
not I_20265 (I347139,I196901);
nand I_20266 (I347156,I347105,I347139);
nor I_20267 (I347173,I196901,I196913);
and I_20268 (I346977,I347173,I347040);
not I_20269 (I347204,I196898);
nand I_20270 (I347221,I347204,I196904);
nor I_20271 (I347238,I196898,I196898);
not I_20272 (I347255,I347238);
nand I_20273 (I346980,I347122,I347255);
DFFARX1 I_20274 (I347238,I2595,I347006,I346995,);
nor I_20275 (I347300,I196907,I196901);
nor I_20276 (I347317,I347300,I196919);
and I_20277 (I347334,I347317,I347221);
DFFARX1 I_20278 (I347334,I2595,I347006,I346992,);
nor I_20279 (I346989,I347300,I347156);
or I_20280 (I346986,I347238,I347300);
nor I_20281 (I347393,I196907,I196922);
DFFARX1 I_20282 (I347393,I2595,I347006,I347419,);
not I_20283 (I347427,I347419);
nand I_20284 (I347444,I347427,I347105);
nor I_20285 (I347461,I347444,I196919);
DFFARX1 I_20286 (I347461,I2595,I347006,I346974,);
nor I_20287 (I347492,I347427,I347156);
nor I_20288 (I346983,I347300,I347492);
not I_20289 (I347550,I2602);
DFFARX1 I_20290 (I310822,I2595,I347550,I347576,);
nand I_20291 (I347584,I347576,I310801);
DFFARX1 I_20292 (I310798,I2595,I347550,I347610,);
DFFARX1 I_20293 (I347610,I2595,I347550,I347627,);
not I_20294 (I347542,I347627);
not I_20295 (I347649,I310810);
nor I_20296 (I347666,I310810,I310819);
not I_20297 (I347683,I310807);
nand I_20298 (I347700,I347649,I347683);
nor I_20299 (I347717,I310807,I310810);
and I_20300 (I347521,I347717,I347584);
not I_20301 (I347748,I310816);
nand I_20302 (I347765,I347748,I310813);
nor I_20303 (I347782,I310816,I310798);
not I_20304 (I347799,I347782);
nand I_20305 (I347524,I347666,I347799);
DFFARX1 I_20306 (I347782,I2595,I347550,I347539,);
nor I_20307 (I347844,I310801,I310807);
nor I_20308 (I347861,I347844,I310819);
and I_20309 (I347878,I347861,I347765);
DFFARX1 I_20310 (I347878,I2595,I347550,I347536,);
nor I_20311 (I347533,I347844,I347700);
or I_20312 (I347530,I347782,I347844);
nor I_20313 (I347937,I310801,I310804);
DFFARX1 I_20314 (I347937,I2595,I347550,I347963,);
not I_20315 (I347971,I347963);
nand I_20316 (I347988,I347971,I347649);
nor I_20317 (I348005,I347988,I310819);
DFFARX1 I_20318 (I348005,I2595,I347550,I347518,);
nor I_20319 (I348036,I347971,I347700);
nor I_20320 (I347527,I347844,I348036);
not I_20321 (I348094,I2602);
DFFARX1 I_20322 (I10281,I2595,I348094,I348120,);
nand I_20323 (I348128,I348120,I10275);
DFFARX1 I_20324 (I10296,I2595,I348094,I348154,);
DFFARX1 I_20325 (I348154,I2595,I348094,I348171,);
not I_20326 (I348086,I348171);
not I_20327 (I348193,I10284);
nor I_20328 (I348210,I10284,I10293);
not I_20329 (I348227,I10272);
nand I_20330 (I348244,I348193,I348227);
nor I_20331 (I348261,I10272,I10284);
and I_20332 (I348065,I348261,I348128);
not I_20333 (I348292,I10290);
nand I_20334 (I348309,I348292,I10278);
nor I_20335 (I348326,I10290,I10272);
not I_20336 (I348343,I348326);
nand I_20337 (I348068,I348210,I348343);
DFFARX1 I_20338 (I348326,I2595,I348094,I348083,);
nor I_20339 (I348388,I10275,I10272);
nor I_20340 (I348405,I348388,I10293);
and I_20341 (I348422,I348405,I348309);
DFFARX1 I_20342 (I348422,I2595,I348094,I348080,);
nor I_20343 (I348077,I348388,I348244);
or I_20344 (I348074,I348326,I348388);
nor I_20345 (I348481,I10275,I10287);
DFFARX1 I_20346 (I348481,I2595,I348094,I348507,);
not I_20347 (I348515,I348507);
nand I_20348 (I348532,I348515,I348193);
nor I_20349 (I348549,I348532,I10293);
DFFARX1 I_20350 (I348549,I2595,I348094,I348062,);
nor I_20351 (I348580,I348515,I348244);
nor I_20352 (I348071,I348388,I348580);
not I_20353 (I348638,I2602);
DFFARX1 I_20354 (I337410,I2595,I348638,I348664,);
nand I_20355 (I348672,I348664,I337389);
DFFARX1 I_20356 (I337386,I2595,I348638,I348698,);
DFFARX1 I_20357 (I348698,I2595,I348638,I348715,);
not I_20358 (I348630,I348715);
not I_20359 (I348737,I337398);
nor I_20360 (I348754,I337398,I337407);
not I_20361 (I348771,I337395);
nand I_20362 (I348788,I348737,I348771);
nor I_20363 (I348805,I337395,I337398);
and I_20364 (I348609,I348805,I348672);
not I_20365 (I348836,I337404);
nand I_20366 (I348853,I348836,I337401);
nor I_20367 (I348870,I337404,I337386);
not I_20368 (I348887,I348870);
nand I_20369 (I348612,I348754,I348887);
DFFARX1 I_20370 (I348870,I2595,I348638,I348627,);
nor I_20371 (I348932,I337389,I337395);
nor I_20372 (I348949,I348932,I337407);
and I_20373 (I348966,I348949,I348853);
DFFARX1 I_20374 (I348966,I2595,I348638,I348624,);
nor I_20375 (I348621,I348932,I348788);
or I_20376 (I348618,I348870,I348932);
nor I_20377 (I349025,I337389,I337392);
DFFARX1 I_20378 (I349025,I2595,I348638,I349051,);
not I_20379 (I349059,I349051);
nand I_20380 (I349076,I349059,I348737);
nor I_20381 (I349093,I349076,I337407);
DFFARX1 I_20382 (I349093,I2595,I348638,I348606,);
nor I_20383 (I349124,I349059,I348788);
nor I_20384 (I348615,I348932,I349124);
not I_20385 (I349182,I2602);
DFFARX1 I_20386 (I140465,I2595,I349182,I349208,);
nand I_20387 (I349216,I349208,I140462);
DFFARX1 I_20388 (I140441,I2595,I349182,I349242,);
DFFARX1 I_20389 (I349242,I2595,I349182,I349259,);
not I_20390 (I349174,I349259);
not I_20391 (I349281,I140456);
nor I_20392 (I349298,I140456,I140459);
not I_20393 (I349315,I140450);
nand I_20394 (I349332,I349281,I349315);
nor I_20395 (I349349,I140450,I140456);
and I_20396 (I349153,I349349,I349216);
not I_20397 (I349380,I140447);
nand I_20398 (I349397,I349380,I140468);
nor I_20399 (I349414,I140447,I140444);
not I_20400 (I349431,I349414);
nand I_20401 (I349156,I349298,I349431);
DFFARX1 I_20402 (I349414,I2595,I349182,I349171,);
nor I_20403 (I349476,I140453,I140450);
nor I_20404 (I349493,I349476,I140459);
and I_20405 (I349510,I349493,I349397);
DFFARX1 I_20406 (I349510,I2595,I349182,I349168,);
nor I_20407 (I349165,I349476,I349332);
or I_20408 (I349162,I349414,I349476);
nor I_20409 (I349569,I140453,I140441);
DFFARX1 I_20410 (I349569,I2595,I349182,I349595,);
not I_20411 (I349603,I349595);
nand I_20412 (I349620,I349603,I349281);
nor I_20413 (I349637,I349620,I140459);
DFFARX1 I_20414 (I349637,I2595,I349182,I349150,);
nor I_20415 (I349668,I349603,I349332);
nor I_20416 (I349159,I349476,I349668);
not I_20417 (I349726,I2602);
DFFARX1 I_20418 (I36116,I2595,I349726,I349752,);
nand I_20419 (I349760,I349752,I36098);
DFFARX1 I_20420 (I36095,I2595,I349726,I349786,);
DFFARX1 I_20421 (I349786,I2595,I349726,I349803,);
not I_20422 (I349718,I349803);
not I_20423 (I349825,I36113);
nor I_20424 (I349842,I36113,I36107);
not I_20425 (I349859,I36095);
nand I_20426 (I349876,I349825,I349859);
nor I_20427 (I349893,I36095,I36113);
and I_20428 (I349697,I349893,I349760);
not I_20429 (I349924,I36104);
nand I_20430 (I349941,I349924,I36110);
nor I_20431 (I349958,I36104,I36098);
not I_20432 (I349975,I349958);
nand I_20433 (I349700,I349842,I349975);
DFFARX1 I_20434 (I349958,I2595,I349726,I349715,);
nor I_20435 (I350020,I36101,I36095);
nor I_20436 (I350037,I350020,I36107);
and I_20437 (I350054,I350037,I349941);
DFFARX1 I_20438 (I350054,I2595,I349726,I349712,);
nor I_20439 (I349709,I350020,I349876);
or I_20440 (I349706,I349958,I350020);
nor I_20441 (I350113,I36101,I36119);
DFFARX1 I_20442 (I350113,I2595,I349726,I350139,);
not I_20443 (I350147,I350139);
nand I_20444 (I350164,I350147,I349825);
nor I_20445 (I350181,I350164,I36107);
DFFARX1 I_20446 (I350181,I2595,I349726,I349694,);
nor I_20447 (I350212,I350147,I349876);
nor I_20448 (I349703,I350020,I350212);
not I_20449 (I350270,I2602);
DFFARX1 I_20450 (I356775,I2595,I350270,I350296,);
nand I_20451 (I350304,I350296,I356784);
DFFARX1 I_20452 (I356787,I2595,I350270,I350330,);
DFFARX1 I_20453 (I350330,I2595,I350270,I350347,);
not I_20454 (I350262,I350347);
not I_20455 (I350369,I356781);
nor I_20456 (I350386,I356781,I356778);
not I_20457 (I350403,I356772);
nand I_20458 (I350420,I350369,I350403);
nor I_20459 (I350437,I356772,I356781);
and I_20460 (I350241,I350437,I350304);
not I_20461 (I350468,I356769);
nand I_20462 (I350485,I350468,I356766);
nor I_20463 (I350502,I356769,I356766);
not I_20464 (I350519,I350502);
nand I_20465 (I350244,I350386,I350519);
DFFARX1 I_20466 (I350502,I2595,I350270,I350259,);
nor I_20467 (I350564,I356769,I356772);
nor I_20468 (I350581,I350564,I356778);
and I_20469 (I350598,I350581,I350485);
DFFARX1 I_20470 (I350598,I2595,I350270,I350256,);
nor I_20471 (I350253,I350564,I350420);
or I_20472 (I350250,I350502,I350564);
nor I_20473 (I350657,I356769,I356790);
DFFARX1 I_20474 (I350657,I2595,I350270,I350683,);
not I_20475 (I350691,I350683);
nand I_20476 (I350708,I350691,I350369);
nor I_20477 (I350725,I350708,I356778);
DFFARX1 I_20478 (I350725,I2595,I350270,I350238,);
nor I_20479 (I350756,I350691,I350420);
nor I_20480 (I350247,I350564,I350756);
not I_20481 (I350814,I2602);
DFFARX1 I_20482 (I48497,I2595,I350814,I350840,);
nand I_20483 (I350848,I350840,I48512);
DFFARX1 I_20484 (I48509,I2595,I350814,I350874,);
DFFARX1 I_20485 (I350874,I2595,I350814,I350891,);
not I_20486 (I350806,I350891);
not I_20487 (I350913,I48488);
nor I_20488 (I350930,I48488,I48494);
not I_20489 (I350947,I48500);
nand I_20490 (I350964,I350913,I350947);
nor I_20491 (I350981,I48500,I48488);
and I_20492 (I350785,I350981,I350848);
not I_20493 (I351012,I48506);
nand I_20494 (I351029,I351012,I48488);
nor I_20495 (I351046,I48506,I48491);
not I_20496 (I351063,I351046);
nand I_20497 (I350788,I350930,I351063);
DFFARX1 I_20498 (I351046,I2595,I350814,I350803,);
nor I_20499 (I351108,I48491,I48500);
nor I_20500 (I351125,I351108,I48494);
and I_20501 (I351142,I351125,I351029);
DFFARX1 I_20502 (I351142,I2595,I350814,I350800,);
nor I_20503 (I350797,I351108,I350964);
or I_20504 (I350794,I351046,I351108);
nor I_20505 (I351201,I48491,I48503);
DFFARX1 I_20506 (I351201,I2595,I350814,I351227,);
not I_20507 (I351235,I351227);
nand I_20508 (I351252,I351235,I350913);
nor I_20509 (I351269,I351252,I48494);
DFFARX1 I_20510 (I351269,I2595,I350814,I350782,);
nor I_20511 (I351300,I351235,I350964);
nor I_20512 (I350791,I351108,I351300);
not I_20513 (I351358,I2602);
DFFARX1 I_20514 (I129585,I2595,I351358,I351384,);
nand I_20515 (I351392,I351384,I129582);
DFFARX1 I_20516 (I129561,I2595,I351358,I351418,);
DFFARX1 I_20517 (I351418,I2595,I351358,I351435,);
not I_20518 (I351350,I351435);
not I_20519 (I351457,I129576);
nor I_20520 (I351474,I129576,I129579);
not I_20521 (I351491,I129570);
nand I_20522 (I351508,I351457,I351491);
nor I_20523 (I351525,I129570,I129576);
and I_20524 (I351329,I351525,I351392);
not I_20525 (I351556,I129567);
nand I_20526 (I351573,I351556,I129588);
nor I_20527 (I351590,I129567,I129564);
not I_20528 (I351607,I351590);
nand I_20529 (I351332,I351474,I351607);
DFFARX1 I_20530 (I351590,I2595,I351358,I351347,);
nor I_20531 (I351652,I129573,I129570);
nor I_20532 (I351669,I351652,I129579);
and I_20533 (I351686,I351669,I351573);
DFFARX1 I_20534 (I351686,I2595,I351358,I351344,);
nor I_20535 (I351341,I351652,I351508);
or I_20536 (I351338,I351590,I351652);
nor I_20537 (I351745,I129573,I129561);
DFFARX1 I_20538 (I351745,I2595,I351358,I351771,);
not I_20539 (I351779,I351771);
nand I_20540 (I351796,I351779,I351457);
nor I_20541 (I351813,I351796,I129579);
DFFARX1 I_20542 (I351813,I2595,I351358,I351326,);
nor I_20543 (I351844,I351779,I351508);
nor I_20544 (I351335,I351652,I351844);
not I_20545 (I351902,I2602);
DFFARX1 I_20546 (I77057,I2595,I351902,I351928,);
nand I_20547 (I351936,I351928,I77072);
DFFARX1 I_20548 (I77069,I2595,I351902,I351962,);
DFFARX1 I_20549 (I351962,I2595,I351902,I351979,);
not I_20550 (I351894,I351979);
not I_20551 (I352001,I77048);
nor I_20552 (I352018,I77048,I77054);
not I_20553 (I352035,I77060);
nand I_20554 (I352052,I352001,I352035);
nor I_20555 (I352069,I77060,I77048);
and I_20556 (I351873,I352069,I351936);
not I_20557 (I352100,I77066);
nand I_20558 (I352117,I352100,I77048);
nor I_20559 (I352134,I77066,I77051);
not I_20560 (I352151,I352134);
nand I_20561 (I351876,I352018,I352151);
DFFARX1 I_20562 (I352134,I2595,I351902,I351891,);
nor I_20563 (I352196,I77051,I77060);
nor I_20564 (I352213,I352196,I77054);
and I_20565 (I352230,I352213,I352117);
DFFARX1 I_20566 (I352230,I2595,I351902,I351888,);
nor I_20567 (I351885,I352196,I352052);
or I_20568 (I351882,I352134,I352196);
nor I_20569 (I352289,I77051,I77063);
DFFARX1 I_20570 (I352289,I2595,I351902,I352315,);
not I_20571 (I352323,I352315);
nand I_20572 (I352340,I352323,I352001);
nor I_20573 (I352357,I352340,I77054);
DFFARX1 I_20574 (I352357,I2595,I351902,I351870,);
nor I_20575 (I352388,I352323,I352052);
nor I_20576 (I351879,I352196,I352388);
not I_20577 (I352446,I2602);
DFFARX1 I_20578 (I363133,I2595,I352446,I352472,);
nand I_20579 (I352480,I352472,I363142);
DFFARX1 I_20580 (I363145,I2595,I352446,I352506,);
DFFARX1 I_20581 (I352506,I2595,I352446,I352523,);
not I_20582 (I352438,I352523);
not I_20583 (I352545,I363139);
nor I_20584 (I352562,I363139,I363136);
not I_20585 (I352579,I363130);
nand I_20586 (I352596,I352545,I352579);
nor I_20587 (I352613,I363130,I363139);
and I_20588 (I352417,I352613,I352480);
not I_20589 (I352644,I363127);
nand I_20590 (I352661,I352644,I363124);
nor I_20591 (I352678,I363127,I363124);
not I_20592 (I352695,I352678);
nand I_20593 (I352420,I352562,I352695);
DFFARX1 I_20594 (I352678,I2595,I352446,I352435,);
nor I_20595 (I352740,I363127,I363130);
nor I_20596 (I352757,I352740,I363136);
and I_20597 (I352774,I352757,I352661);
DFFARX1 I_20598 (I352774,I2595,I352446,I352432,);
nor I_20599 (I352429,I352740,I352596);
or I_20600 (I352426,I352678,I352740);
nor I_20601 (I352833,I363127,I363148);
DFFARX1 I_20602 (I352833,I2595,I352446,I352859,);
not I_20603 (I352867,I352859);
nand I_20604 (I352884,I352867,I352545);
nor I_20605 (I352901,I352884,I363136);
DFFARX1 I_20606 (I352901,I2595,I352446,I352414,);
nor I_20607 (I352932,I352867,I352596);
nor I_20608 (I352423,I352740,I352932);
not I_20609 (I352990,I2602);
DFFARX1 I_20610 (I25049,I2595,I352990,I353016,);
nand I_20611 (I353024,I353016,I25031);
DFFARX1 I_20612 (I25028,I2595,I352990,I353050,);
DFFARX1 I_20613 (I353050,I2595,I352990,I353067,);
not I_20614 (I352982,I353067);
not I_20615 (I353089,I25046);
nor I_20616 (I353106,I25046,I25040);
not I_20617 (I353123,I25028);
nand I_20618 (I353140,I353089,I353123);
nor I_20619 (I353157,I25028,I25046);
and I_20620 (I352961,I353157,I353024);
not I_20621 (I353188,I25037);
nand I_20622 (I353205,I353188,I25043);
nor I_20623 (I353222,I25037,I25031);
not I_20624 (I353239,I353222);
nand I_20625 (I352964,I353106,I353239);
DFFARX1 I_20626 (I353222,I2595,I352990,I352979,);
nor I_20627 (I353284,I25034,I25028);
nor I_20628 (I353301,I353284,I25040);
and I_20629 (I353318,I353301,I353205);
DFFARX1 I_20630 (I353318,I2595,I352990,I352976,);
nor I_20631 (I352973,I353284,I353140);
or I_20632 (I352970,I353222,I353284);
nor I_20633 (I353377,I25034,I25052);
DFFARX1 I_20634 (I353377,I2595,I352990,I353403,);
not I_20635 (I353411,I353403);
nand I_20636 (I353428,I353411,I353089);
nor I_20637 (I353445,I353428,I25040);
DFFARX1 I_20638 (I353445,I2595,I352990,I352958,);
nor I_20639 (I353476,I353411,I353140);
nor I_20640 (I352967,I353284,I353476);
not I_20641 (I353534,I2602);
DFFARX1 I_20642 (I274469,I2595,I353534,I353560,);
nand I_20643 (I353568,I353560,I274469);
DFFARX1 I_20644 (I274481,I2595,I353534,I353594,);
DFFARX1 I_20645 (I353594,I2595,I353534,I353611,);
not I_20646 (I353526,I353611);
not I_20647 (I353633,I274475);
nor I_20648 (I353650,I274475,I274496);
not I_20649 (I353667,I274484);
nand I_20650 (I353684,I353633,I353667);
nor I_20651 (I353701,I274484,I274475);
and I_20652 (I353505,I353701,I353568);
not I_20653 (I353732,I274478);
nand I_20654 (I353749,I353732,I274493);
nor I_20655 (I353766,I274478,I274487);
not I_20656 (I353783,I353766);
nand I_20657 (I353508,I353650,I353783);
DFFARX1 I_20658 (I353766,I2595,I353534,I353523,);
nor I_20659 (I353828,I274490,I274484);
nor I_20660 (I353845,I353828,I274496);
and I_20661 (I353862,I353845,I353749);
DFFARX1 I_20662 (I353862,I2595,I353534,I353520,);
nor I_20663 (I353517,I353828,I353684);
or I_20664 (I353514,I353766,I353828);
nor I_20665 (I353921,I274490,I274472);
DFFARX1 I_20666 (I353921,I2595,I353534,I353947,);
not I_20667 (I353955,I353947);
nand I_20668 (I353972,I353955,I353633);
nor I_20669 (I353989,I353972,I274496);
DFFARX1 I_20670 (I353989,I2595,I353534,I353502,);
nor I_20671 (I354020,I353955,I353684);
nor I_20672 (I353511,I353828,I354020);
not I_20673 (I354078,I2602);
DFFARX1 I_20674 (I176689,I2595,I354078,I354104,);
nand I_20675 (I354112,I354104,I176677);
DFFARX1 I_20676 (I176683,I2595,I354078,I354138,);
DFFARX1 I_20677 (I354138,I2595,I354078,I354155,);
not I_20678 (I354070,I354155);
not I_20679 (I354177,I176668);
nor I_20680 (I354194,I176668,I176680);
not I_20681 (I354211,I176671);
nand I_20682 (I354228,I354177,I354211);
nor I_20683 (I354245,I176671,I176668);
and I_20684 (I354049,I354245,I354112);
not I_20685 (I354276,I176686);
nand I_20686 (I354293,I354276,I176668);
nor I_20687 (I354310,I176686,I176692);
not I_20688 (I354327,I354310);
nand I_20689 (I354052,I354194,I354327);
DFFARX1 I_20690 (I354310,I2595,I354078,I354067,);
nor I_20691 (I354372,I176674,I176671);
nor I_20692 (I354389,I354372,I176680);
and I_20693 (I354406,I354389,I354293);
DFFARX1 I_20694 (I354406,I2595,I354078,I354064,);
nor I_20695 (I354061,I354372,I354228);
or I_20696 (I354058,I354310,I354372);
nor I_20697 (I354465,I176674,I176671);
DFFARX1 I_20698 (I354465,I2595,I354078,I354491,);
not I_20699 (I354499,I354491);
nand I_20700 (I354516,I354499,I354177);
nor I_20701 (I354533,I354516,I176680);
DFFARX1 I_20702 (I354533,I2595,I354078,I354046,);
nor I_20703 (I354564,I354499,I354228);
nor I_20704 (I354055,I354372,I354564);
not I_20705 (I354622,I2602);
DFFARX1 I_20706 (I273177,I2595,I354622,I354648,);
nand I_20707 (I354656,I354648,I273177);
DFFARX1 I_20708 (I273189,I2595,I354622,I354682,);
DFFARX1 I_20709 (I354682,I2595,I354622,I354699,);
not I_20710 (I354614,I354699);
not I_20711 (I354721,I273183);
nor I_20712 (I354738,I273183,I273204);
not I_20713 (I354755,I273192);
nand I_20714 (I354772,I354721,I354755);
nor I_20715 (I354789,I273192,I273183);
and I_20716 (I354593,I354789,I354656);
not I_20717 (I354820,I273186);
nand I_20718 (I354837,I354820,I273201);
nor I_20719 (I354854,I273186,I273195);
not I_20720 (I354871,I354854);
nand I_20721 (I354596,I354738,I354871);
DFFARX1 I_20722 (I354854,I2595,I354622,I354611,);
nor I_20723 (I354916,I273198,I273192);
nor I_20724 (I354933,I354916,I273204);
and I_20725 (I354950,I354933,I354837);
DFFARX1 I_20726 (I354950,I2595,I354622,I354608,);
nor I_20727 (I354605,I354916,I354772);
or I_20728 (I354602,I354854,I354916);
nor I_20729 (I355009,I273198,I273180);
DFFARX1 I_20730 (I355009,I2595,I354622,I355035,);
not I_20731 (I355043,I355035);
nand I_20732 (I355060,I355043,I354721);
nor I_20733 (I355077,I355060,I273204);
DFFARX1 I_20734 (I355077,I2595,I354622,I354590,);
nor I_20735 (I355108,I355043,I354772);
nor I_20736 (I354599,I354916,I355108);
not I_20737 (I355166,I2602);
DFFARX1 I_20738 (I263487,I2595,I355166,I355192,);
nand I_20739 (I355200,I355192,I263487);
DFFARX1 I_20740 (I263499,I2595,I355166,I355226,);
DFFARX1 I_20741 (I355226,I2595,I355166,I355243,);
not I_20742 (I355158,I355243);
not I_20743 (I355265,I263493);
nor I_20744 (I355282,I263493,I263514);
not I_20745 (I355299,I263502);
nand I_20746 (I355316,I355265,I355299);
nor I_20747 (I355333,I263502,I263493);
and I_20748 (I355137,I355333,I355200);
not I_20749 (I355364,I263496);
nand I_20750 (I355381,I355364,I263511);
nor I_20751 (I355398,I263496,I263505);
not I_20752 (I355415,I355398);
nand I_20753 (I355140,I355282,I355415);
DFFARX1 I_20754 (I355398,I2595,I355166,I355155,);
nor I_20755 (I355460,I263508,I263502);
nor I_20756 (I355477,I355460,I263514);
and I_20757 (I355494,I355477,I355381);
DFFARX1 I_20758 (I355494,I2595,I355166,I355152,);
nor I_20759 (I355149,I355460,I355316);
or I_20760 (I355146,I355398,I355460);
nor I_20761 (I355553,I263508,I263490);
DFFARX1 I_20762 (I355553,I2595,I355166,I355579,);
not I_20763 (I355587,I355579);
nand I_20764 (I355604,I355587,I355265);
nor I_20765 (I355621,I355604,I263514);
DFFARX1 I_20766 (I355621,I2595,I355166,I355134,);
nor I_20767 (I355652,I355587,I355316);
nor I_20768 (I355143,I355460,I355652);
not I_20769 (I355710,I2602);
DFFARX1 I_20770 (I198635,I2595,I355710,I355736,);
nand I_20771 (I355744,I355736,I198650);
DFFARX1 I_20772 (I198644,I2595,I355710,I355770,);
DFFARX1 I_20773 (I355770,I2595,I355710,I355787,);
not I_20774 (I355702,I355787);
not I_20775 (I355809,I198647);
nor I_20776 (I355826,I198647,I198653);
not I_20777 (I355843,I198635);
nand I_20778 (I355860,I355809,I355843);
nor I_20779 (I355877,I198635,I198647);
and I_20780 (I355681,I355877,I355744);
not I_20781 (I355908,I198632);
nand I_20782 (I355925,I355908,I198638);
nor I_20783 (I355942,I198632,I198632);
not I_20784 (I355959,I355942);
nand I_20785 (I355684,I355826,I355959);
DFFARX1 I_20786 (I355942,I2595,I355710,I355699,);
nor I_20787 (I356004,I198641,I198635);
nor I_20788 (I356021,I356004,I198653);
and I_20789 (I356038,I356021,I355925);
DFFARX1 I_20790 (I356038,I2595,I355710,I355696,);
nor I_20791 (I355693,I356004,I355860);
or I_20792 (I355690,I355942,I356004);
nor I_20793 (I356097,I198641,I198656);
DFFARX1 I_20794 (I356097,I2595,I355710,I356123,);
not I_20795 (I356131,I356123);
nand I_20796 (I356148,I356131,I355809);
nor I_20797 (I356165,I356148,I198653);
DFFARX1 I_20798 (I356165,I2595,I355710,I355678,);
nor I_20799 (I356196,I356131,I355860);
nor I_20800 (I355687,I356004,I356196);
not I_20801 (I356254,I2602);
DFFARX1 I_20802 (I53852,I2595,I356254,I356280,);
nand I_20803 (I356288,I356280,I53867);
DFFARX1 I_20804 (I53864,I2595,I356254,I356314,);
DFFARX1 I_20805 (I356314,I2595,I356254,I356331,);
not I_20806 (I356246,I356331);
not I_20807 (I356353,I53843);
nor I_20808 (I356370,I53843,I53849);
not I_20809 (I356387,I53855);
nand I_20810 (I356404,I356353,I356387);
nor I_20811 (I356421,I53855,I53843);
and I_20812 (I356225,I356421,I356288);
not I_20813 (I356452,I53861);
nand I_20814 (I356469,I356452,I53843);
nor I_20815 (I356486,I53861,I53846);
not I_20816 (I356503,I356486);
nand I_20817 (I356228,I356370,I356503);
DFFARX1 I_20818 (I356486,I2595,I356254,I356243,);
nor I_20819 (I356548,I53846,I53855);
nor I_20820 (I356565,I356548,I53849);
and I_20821 (I356582,I356565,I356469);
DFFARX1 I_20822 (I356582,I2595,I356254,I356240,);
nor I_20823 (I356237,I356548,I356404);
or I_20824 (I356234,I356486,I356548);
nor I_20825 (I356641,I53846,I53858);
DFFARX1 I_20826 (I356641,I2595,I356254,I356667,);
not I_20827 (I356675,I356667);
nand I_20828 (I356692,I356675,I356353);
nor I_20829 (I356709,I356692,I53849);
DFFARX1 I_20830 (I356709,I2595,I356254,I356222,);
nor I_20831 (I356740,I356675,I356404);
nor I_20832 (I356231,I356548,I356740);
not I_20833 (I356798,I2602);
DFFARX1 I_20834 (I135548,I2595,I356798,I356824,);
nand I_20835 (I356832,I356824,I135557);
not I_20836 (I356849,I356832);
DFFARX1 I_20837 (I135545,I2595,I356798,I356875,);
not I_20838 (I356883,I356875);
not I_20839 (I356900,I135551);
or I_20840 (I356917,I135545,I135551);
nor I_20841 (I356934,I135545,I135551);
or I_20842 (I356951,I135560,I135545);
DFFARX1 I_20843 (I356951,I2595,I356798,I356790,);
not I_20844 (I356982,I135554);
nand I_20845 (I356999,I356982,I135569);
nand I_20846 (I357016,I356900,I356999);
and I_20847 (I356769,I356883,I357016);
nor I_20848 (I357047,I135554,I135572);
and I_20849 (I357064,I356883,I357047);
nor I_20850 (I356775,I356849,I357064);
DFFARX1 I_20851 (I357047,I2595,I356798,I357104,);
not I_20852 (I357112,I357104);
nor I_20853 (I356784,I356883,I357112);
or I_20854 (I357143,I356951,I135563);
nor I_20855 (I357160,I135563,I135560);
nand I_20856 (I357177,I357016,I357160);
nand I_20857 (I357194,I357143,I357177);
DFFARX1 I_20858 (I357194,I2595,I356798,I356787,);
nor I_20859 (I357225,I357160,I356917);
DFFARX1 I_20860 (I357225,I2595,I356798,I356766,);
nor I_20861 (I357256,I135563,I135566);
DFFARX1 I_20862 (I357256,I2595,I356798,I357282,);
DFFARX1 I_20863 (I357282,I2595,I356798,I356781,);
not I_20864 (I357304,I357282);
nand I_20865 (I356778,I357304,I356832);
nand I_20866 (I356772,I357304,I356934);
not I_20867 (I357376,I2602);
DFFARX1 I_20868 (I168579,I2595,I357376,I357402,);
nand I_20869 (I357410,I357402,I168594);
not I_20870 (I357427,I357410);
DFFARX1 I_20871 (I168576,I2595,I357376,I357453,);
not I_20872 (I357461,I357453);
not I_20873 (I357478,I168585);
or I_20874 (I357495,I168579,I168585);
nor I_20875 (I357512,I168579,I168585);
or I_20876 (I357529,I168576,I168579);
DFFARX1 I_20877 (I357529,I2595,I357376,I357368,);
not I_20878 (I357560,I168597);
nand I_20879 (I357577,I357560,I168600);
nand I_20880 (I357594,I357478,I357577);
and I_20881 (I357347,I357461,I357594);
nor I_20882 (I357625,I168597,I168582);
and I_20883 (I357642,I357461,I357625);
nor I_20884 (I357353,I357427,I357642);
DFFARX1 I_20885 (I357625,I2595,I357376,I357682,);
not I_20886 (I357690,I357682);
nor I_20887 (I357362,I357461,I357690);
or I_20888 (I357721,I357529,I168588);
nor I_20889 (I357738,I168588,I168576);
nand I_20890 (I357755,I357594,I357738);
nand I_20891 (I357772,I357721,I357755);
DFFARX1 I_20892 (I357772,I2595,I357376,I357365,);
nor I_20893 (I357803,I357738,I357495);
DFFARX1 I_20894 (I357803,I2595,I357376,I357344,);
nor I_20895 (I357834,I168588,I168591);
DFFARX1 I_20896 (I357834,I2595,I357376,I357860,);
DFFARX1 I_20897 (I357860,I2595,I357376,I357359,);
not I_20898 (I357882,I357860);
nand I_20899 (I357356,I357882,I357410);
nand I_20900 (I357350,I357882,I357512);
not I_20901 (I357954,I2602);
DFFARX1 I_20902 (I186494,I2595,I357954,I357980,);
nand I_20903 (I357988,I357980,I186497);
not I_20904 (I358005,I357988);
DFFARX1 I_20905 (I186509,I2595,I357954,I358031,);
not I_20906 (I358039,I358031);
not I_20907 (I358056,I186494);
or I_20908 (I358073,I186503,I186494);
nor I_20909 (I358090,I186503,I186494);
or I_20910 (I358107,I186512,I186503);
DFFARX1 I_20911 (I358107,I2595,I357954,I357946,);
not I_20912 (I358138,I186515);
nand I_20913 (I358155,I358138,I186497);
nand I_20914 (I358172,I358056,I358155);
and I_20915 (I357925,I358039,I358172);
nor I_20916 (I358203,I186515,I186500);
and I_20917 (I358220,I358039,I358203);
nor I_20918 (I357931,I358005,I358220);
DFFARX1 I_20919 (I358203,I2595,I357954,I358260,);
not I_20920 (I358268,I358260);
nor I_20921 (I357940,I358039,I358268);
or I_20922 (I358299,I358107,I186506);
nor I_20923 (I358316,I186506,I186512);
nand I_20924 (I358333,I358172,I358316);
nand I_20925 (I358350,I358299,I358333);
DFFARX1 I_20926 (I358350,I2595,I357954,I357943,);
nor I_20927 (I358381,I358316,I358073);
DFFARX1 I_20928 (I358381,I2595,I357954,I357922,);
nor I_20929 (I358412,I186506,I186518);
DFFARX1 I_20930 (I358412,I2595,I357954,I358438,);
DFFARX1 I_20931 (I358438,I2595,I357954,I357937,);
not I_20932 (I358460,I358438);
nand I_20933 (I357934,I358460,I357988);
nand I_20934 (I357928,I358460,I358090);
not I_20935 (I358532,I2602);
DFFARX1 I_20936 (I41377,I2595,I358532,I358558,);
nand I_20937 (I358566,I358558,I41368);
not I_20938 (I358583,I358566);
DFFARX1 I_20939 (I41365,I2595,I358532,I358609,);
not I_20940 (I358617,I358609);
not I_20941 (I358634,I41374);
or I_20942 (I358651,I41365,I41374);
nor I_20943 (I358668,I41365,I41374);
or I_20944 (I358685,I41371,I41365);
DFFARX1 I_20945 (I358685,I2595,I358532,I358524,);
not I_20946 (I358716,I41380);
nand I_20947 (I358733,I358716,I41389);
nand I_20948 (I358750,I358634,I358733);
and I_20949 (I358503,I358617,I358750);
nor I_20950 (I358781,I41380,I41383);
and I_20951 (I358798,I358617,I358781);
nor I_20952 (I358509,I358583,I358798);
DFFARX1 I_20953 (I358781,I2595,I358532,I358838,);
not I_20954 (I358846,I358838);
nor I_20955 (I358518,I358617,I358846);
or I_20956 (I358877,I358685,I41368);
nor I_20957 (I358894,I41368,I41371);
nand I_20958 (I358911,I358750,I358894);
nand I_20959 (I358928,I358877,I358911);
DFFARX1 I_20960 (I358928,I2595,I358532,I358521,);
nor I_20961 (I358959,I358894,I358651);
DFFARX1 I_20962 (I358959,I2595,I358532,I358500,);
nor I_20963 (I358990,I41368,I41386);
DFFARX1 I_20964 (I358990,I2595,I358532,I359016,);
DFFARX1 I_20965 (I359016,I2595,I358532,I358515,);
not I_20966 (I359038,I359016);
nand I_20967 (I358512,I359038,I358566);
nand I_20968 (I358506,I359038,I358668);
not I_20969 (I359110,I2602);
DFFARX1 I_20970 (I226954,I2595,I359110,I359136,);
nand I_20971 (I359144,I359136,I226957);
not I_20972 (I359161,I359144);
DFFARX1 I_20973 (I226969,I2595,I359110,I359187,);
not I_20974 (I359195,I359187);
not I_20975 (I359212,I226954);
or I_20976 (I359229,I226963,I226954);
nor I_20977 (I359246,I226963,I226954);
or I_20978 (I359263,I226972,I226963);
DFFARX1 I_20979 (I359263,I2595,I359110,I359102,);
not I_20980 (I359294,I226975);
nand I_20981 (I359311,I359294,I226957);
nand I_20982 (I359328,I359212,I359311);
and I_20983 (I359081,I359195,I359328);
nor I_20984 (I359359,I226975,I226960);
and I_20985 (I359376,I359195,I359359);
nor I_20986 (I359087,I359161,I359376);
DFFARX1 I_20987 (I359359,I2595,I359110,I359416,);
not I_20988 (I359424,I359416);
nor I_20989 (I359096,I359195,I359424);
or I_20990 (I359455,I359263,I226966);
nor I_20991 (I359472,I226966,I226972);
nand I_20992 (I359489,I359328,I359472);
nand I_20993 (I359506,I359455,I359489);
DFFARX1 I_20994 (I359506,I2595,I359110,I359099,);
nor I_20995 (I359537,I359472,I359229);
DFFARX1 I_20996 (I359537,I2595,I359110,I359078,);
nor I_20997 (I359568,I226966,I226978);
DFFARX1 I_20998 (I359568,I2595,I359110,I359594,);
DFFARX1 I_20999 (I359594,I2595,I359110,I359093,);
not I_21000 (I359616,I359594);
nand I_21001 (I359090,I359616,I359144);
nand I_21002 (I359084,I359616,I359246);
not I_21003 (I359688,I2602);
DFFARX1 I_21004 (I98542,I2595,I359688,I359714,);
nand I_21005 (I359722,I359714,I98563);
not I_21006 (I359739,I359722);
DFFARX1 I_21007 (I98557,I2595,I359688,I359765,);
not I_21008 (I359773,I359765);
not I_21009 (I359790,I98545);
or I_21010 (I359807,I98560,I98545);
nor I_21011 (I359824,I98560,I98545);
or I_21012 (I359841,I98551,I98560);
DFFARX1 I_21013 (I359841,I2595,I359688,I359680,);
not I_21014 (I359872,I98539);
nand I_21015 (I359889,I359872,I98536);
nand I_21016 (I359906,I359790,I359889);
and I_21017 (I359659,I359773,I359906);
nor I_21018 (I359937,I98539,I98548);
and I_21019 (I359954,I359773,I359937);
nor I_21020 (I359665,I359739,I359954);
DFFARX1 I_21021 (I359937,I2595,I359688,I359994,);
not I_21022 (I360002,I359994);
nor I_21023 (I359674,I359773,I360002);
or I_21024 (I360033,I359841,I98554);
nor I_21025 (I360050,I98554,I98551);
nand I_21026 (I360067,I359906,I360050);
nand I_21027 (I360084,I360033,I360067);
DFFARX1 I_21028 (I360084,I2595,I359688,I359677,);
nor I_21029 (I360115,I360050,I359807);
DFFARX1 I_21030 (I360115,I2595,I359688,I359656,);
nor I_21031 (I360146,I98554,I98536);
DFFARX1 I_21032 (I360146,I2595,I359688,I360172,);
DFFARX1 I_21033 (I360172,I2595,I359688,I359671,);
not I_21034 (I360194,I360172);
nand I_21035 (I359668,I360194,I359722);
nand I_21036 (I359662,I360194,I359824);
not I_21037 (I360266,I2602);
DFFARX1 I_21038 (I198054,I2595,I360266,I360292,);
nand I_21039 (I360300,I360292,I198057);
not I_21040 (I360317,I360300);
DFFARX1 I_21041 (I198069,I2595,I360266,I360343,);
not I_21042 (I360351,I360343);
not I_21043 (I360368,I198054);
or I_21044 (I360385,I198063,I198054);
nor I_21045 (I360402,I198063,I198054);
or I_21046 (I360419,I198072,I198063);
DFFARX1 I_21047 (I360419,I2595,I360266,I360258,);
not I_21048 (I360450,I198075);
nand I_21049 (I360467,I360450,I198057);
nand I_21050 (I360484,I360368,I360467);
and I_21051 (I360237,I360351,I360484);
nor I_21052 (I360515,I198075,I198060);
and I_21053 (I360532,I360351,I360515);
nor I_21054 (I360243,I360317,I360532);
DFFARX1 I_21055 (I360515,I2595,I360266,I360572,);
not I_21056 (I360580,I360572);
nor I_21057 (I360252,I360351,I360580);
or I_21058 (I360611,I360419,I198066);
nor I_21059 (I360628,I198066,I198072);
nand I_21060 (I360645,I360484,I360628);
nand I_21061 (I360662,I360611,I360645);
DFFARX1 I_21062 (I360662,I2595,I360266,I360255,);
nor I_21063 (I360693,I360628,I360385);
DFFARX1 I_21064 (I360693,I2595,I360266,I360234,);
nor I_21065 (I360724,I198066,I198078);
DFFARX1 I_21066 (I360724,I2595,I360266,I360750,);
DFFARX1 I_21067 (I360750,I2595,I360266,I360249,);
not I_21068 (I360772,I360750);
nand I_21069 (I360246,I360772,I360300);
nand I_21070 (I360240,I360772,I360402);
not I_21071 (I360844,I2602);
DFFARX1 I_21072 (I232482,I2595,I360844,I360870,);
nand I_21073 (I360878,I360870,I232482);
not I_21074 (I360895,I360878);
DFFARX1 I_21075 (I232488,I2595,I360844,I360921,);
not I_21076 (I360929,I360921);
not I_21077 (I360946,I232500);
or I_21078 (I360963,I232485,I232500);
nor I_21079 (I360980,I232485,I232500);
or I_21080 (I360997,I232479,I232485);
DFFARX1 I_21081 (I360997,I2595,I360844,I360836,);
not I_21082 (I361028,I232497);
nand I_21083 (I361045,I361028,I232491);
nand I_21084 (I361062,I360946,I361045);
and I_21085 (I360815,I360929,I361062);
nor I_21086 (I361093,I232497,I232479);
and I_21087 (I361110,I360929,I361093);
nor I_21088 (I360821,I360895,I361110);
DFFARX1 I_21089 (I361093,I2595,I360844,I361150,);
not I_21090 (I361158,I361150);
nor I_21091 (I360830,I360929,I361158);
or I_21092 (I361189,I360997,I232494);
nor I_21093 (I361206,I232494,I232479);
nand I_21094 (I361223,I361062,I361206);
nand I_21095 (I361240,I361189,I361223);
DFFARX1 I_21096 (I361240,I2595,I360844,I360833,);
nor I_21097 (I361271,I361206,I360963);
DFFARX1 I_21098 (I361271,I2595,I360844,I360812,);
nor I_21099 (I361302,I232494,I232485);
DFFARX1 I_21100 (I361302,I2595,I360844,I361328,);
DFFARX1 I_21101 (I361328,I2595,I360844,I360827,);
not I_21102 (I361350,I361328);
nand I_21103 (I360824,I361350,I360878);
nand I_21104 (I360818,I361350,I360980);
not I_21105 (I361422,I2602);
DFFARX1 I_21106 (I1748,I2595,I361422,I361448,);
nand I_21107 (I361456,I361448,I1452);
not I_21108 (I361473,I361456);
DFFARX1 I_21109 (I2436,I2595,I361422,I361499,);
not I_21110 (I361507,I361499);
not I_21111 (I361524,I2516);
or I_21112 (I361541,I1820,I2516);
nor I_21113 (I361558,I1820,I2516);
or I_21114 (I361575,I2020,I1820);
DFFARX1 I_21115 (I361575,I2595,I361422,I361414,);
not I_21116 (I361606,I1836);
nand I_21117 (I361623,I361606,I1868);
nand I_21118 (I361640,I361524,I361623);
and I_21119 (I361393,I361507,I361640);
nor I_21120 (I361671,I1836,I1668);
and I_21121 (I361688,I361507,I361671);
nor I_21122 (I361399,I361473,I361688);
DFFARX1 I_21123 (I361671,I2595,I361422,I361728,);
not I_21124 (I361736,I361728);
nor I_21125 (I361408,I361507,I361736);
or I_21126 (I361767,I361575,I1956);
nor I_21127 (I361784,I1956,I2020);
nand I_21128 (I361801,I361640,I361784);
nand I_21129 (I361818,I361767,I361801);
DFFARX1 I_21130 (I361818,I2595,I361422,I361411,);
nor I_21131 (I361849,I361784,I361541);
DFFARX1 I_21132 (I361849,I2595,I361422,I361390,);
nor I_21133 (I361880,I1956,I1740);
DFFARX1 I_21134 (I361880,I2595,I361422,I361906,);
DFFARX1 I_21135 (I361906,I2595,I361422,I361405,);
not I_21136 (I361928,I361906);
nand I_21137 (I361402,I361928,I361456);
nand I_21138 (I361396,I361928,I361558);
not I_21139 (I362000,I2602);
DFFARX1 I_21140 (I30310,I2595,I362000,I362026,);
nand I_21141 (I362034,I362026,I30301);
not I_21142 (I362051,I362034);
DFFARX1 I_21143 (I30298,I2595,I362000,I362077,);
not I_21144 (I362085,I362077);
not I_21145 (I362102,I30307);
or I_21146 (I362119,I30298,I30307);
nor I_21147 (I362136,I30298,I30307);
or I_21148 (I362153,I30304,I30298);
DFFARX1 I_21149 (I362153,I2595,I362000,I361992,);
not I_21150 (I362184,I30313);
nand I_21151 (I362201,I362184,I30322);
nand I_21152 (I362218,I362102,I362201);
and I_21153 (I361971,I362085,I362218);
nor I_21154 (I362249,I30313,I30316);
and I_21155 (I362266,I362085,I362249);
nor I_21156 (I361977,I362051,I362266);
DFFARX1 I_21157 (I362249,I2595,I362000,I362306,);
not I_21158 (I362314,I362306);
nor I_21159 (I361986,I362085,I362314);
or I_21160 (I362345,I362153,I30301);
nor I_21161 (I362362,I30301,I30304);
nand I_21162 (I362379,I362218,I362362);
nand I_21163 (I362396,I362345,I362379);
DFFARX1 I_21164 (I362396,I2595,I362000,I361989,);
nor I_21165 (I362427,I362362,I362119);
DFFARX1 I_21166 (I362427,I2595,I362000,I361968,);
nor I_21167 (I362458,I30301,I30319);
DFFARX1 I_21168 (I362458,I2595,I362000,I362484,);
DFFARX1 I_21169 (I362484,I2595,I362000,I361983,);
not I_21170 (I362506,I362484);
nand I_21171 (I361980,I362506,I362034);
nand I_21172 (I361974,I362506,I362136);
not I_21173 (I362578,I2602);
DFFARX1 I_21174 (I332202,I2595,I362578,I362604,);
nand I_21175 (I362612,I362604,I332187);
not I_21176 (I362629,I362612);
DFFARX1 I_21177 (I332190,I2595,I362578,I362655,);
not I_21178 (I362663,I362655);
not I_21179 (I362680,I332205);
or I_21180 (I362697,I332208,I332205);
nor I_21181 (I362714,I332208,I332205);
or I_21182 (I362731,I332184,I332208);
DFFARX1 I_21183 (I362731,I2595,I362578,I362570,);
not I_21184 (I362762,I332196);
nand I_21185 (I362779,I362762,I332199);
nand I_21186 (I362796,I362680,I362779);
and I_21187 (I362549,I362663,I362796);
nor I_21188 (I362827,I332196,I332193);
and I_21189 (I362844,I362663,I362827);
nor I_21190 (I362555,I362629,I362844);
DFFARX1 I_21191 (I362827,I2595,I362578,I362884,);
not I_21192 (I362892,I362884);
nor I_21193 (I362564,I362663,I362892);
or I_21194 (I362923,I362731,I332184);
nor I_21195 (I362940,I332184,I332184);
nand I_21196 (I362957,I362796,I362940);
nand I_21197 (I362974,I362923,I362957);
DFFARX1 I_21198 (I362974,I2595,I362578,I362567,);
nor I_21199 (I363005,I362940,I362697);
DFFARX1 I_21200 (I363005,I2595,I362578,I362546,);
nor I_21201 (I363036,I332184,I332187);
DFFARX1 I_21202 (I363036,I2595,I362578,I363062,);
DFFARX1 I_21203 (I363062,I2595,I362578,I362561,);
not I_21204 (I363084,I363062);
nand I_21205 (I362558,I363084,I362612);
nand I_21206 (I362552,I363084,I362714);
not I_21207 (I363156,I2602);
DFFARX1 I_21208 (I52653,I2595,I363156,I363182,);
nand I_21209 (I363190,I363182,I52656);
not I_21210 (I363207,I363190);
DFFARX1 I_21211 (I52665,I2595,I363156,I363233,);
not I_21212 (I363241,I363233);
not I_21213 (I363258,I52668);
or I_21214 (I363275,I52659,I52668);
nor I_21215 (I363292,I52659,I52668);
or I_21216 (I363309,I52671,I52659);
DFFARX1 I_21217 (I363309,I2595,I363156,I363148,);
not I_21218 (I363340,I52656);
nand I_21219 (I363357,I363340,I52662);
nand I_21220 (I363374,I363258,I363357);
and I_21221 (I363127,I363241,I363374);
nor I_21222 (I363405,I52656,I52674);
and I_21223 (I363422,I363241,I363405);
nor I_21224 (I363133,I363207,I363422);
DFFARX1 I_21225 (I363405,I2595,I363156,I363462,);
not I_21226 (I363470,I363462);
nor I_21227 (I363142,I363241,I363470);
or I_21228 (I363501,I363309,I52653);
nor I_21229 (I363518,I52653,I52671);
nand I_21230 (I363535,I363374,I363518);
nand I_21231 (I363552,I363501,I363535);
DFFARX1 I_21232 (I363552,I2595,I363156,I363145,);
nor I_21233 (I363583,I363518,I363275);
DFFARX1 I_21234 (I363583,I2595,I363156,I363124,);
nor I_21235 (I363614,I52653,I52677);
DFFARX1 I_21236 (I363614,I2595,I363156,I363640,);
DFFARX1 I_21237 (I363640,I2595,I363156,I363139,);
not I_21238 (I363662,I363640);
nand I_21239 (I363136,I363662,I363190);
nand I_21240 (I363130,I363662,I363292);
not I_21241 (I363734,I2602);
DFFARX1 I_21242 (I334514,I2595,I363734,I363760,);
nand I_21243 (I363768,I363760,I334499);
not I_21244 (I363785,I363768);
DFFARX1 I_21245 (I334502,I2595,I363734,I363811,);
not I_21246 (I363819,I363811);
not I_21247 (I363836,I334517);
or I_21248 (I363853,I334520,I334517);
nor I_21249 (I363870,I334520,I334517);
or I_21250 (I363887,I334496,I334520);
DFFARX1 I_21251 (I363887,I2595,I363734,I363726,);
not I_21252 (I363918,I334508);
nand I_21253 (I363935,I363918,I334511);
nand I_21254 (I363952,I363836,I363935);
and I_21255 (I363705,I363819,I363952);
nor I_21256 (I363983,I334508,I334505);
and I_21257 (I364000,I363819,I363983);
nor I_21258 (I363711,I363785,I364000);
DFFARX1 I_21259 (I363983,I2595,I363734,I364040,);
not I_21260 (I364048,I364040);
nor I_21261 (I363720,I363819,I364048);
or I_21262 (I364079,I363887,I334496);
nor I_21263 (I364096,I334496,I334496);
nand I_21264 (I364113,I363952,I364096);
nand I_21265 (I364130,I364079,I364113);
DFFARX1 I_21266 (I364130,I2595,I363734,I363723,);
nor I_21267 (I364161,I364096,I363853);
DFFARX1 I_21268 (I364161,I2595,I363734,I363702,);
nor I_21269 (I364192,I334496,I334499);
DFFARX1 I_21270 (I364192,I2595,I363734,I364218,);
DFFARX1 I_21271 (I364218,I2595,I363734,I363717,);
not I_21272 (I364240,I364218);
nand I_21273 (I363714,I364240,I363768);
nand I_21274 (I363708,I364240,I363870);
not I_21275 (I364312,I2602);
DFFARX1 I_21276 (I244076,I2595,I364312,I364338,);
nand I_21277 (I364346,I364338,I244076);
not I_21278 (I364363,I364346);
DFFARX1 I_21279 (I244082,I2595,I364312,I364389,);
not I_21280 (I364397,I364389);
not I_21281 (I364414,I244094);
or I_21282 (I364431,I244079,I244094);
nor I_21283 (I364448,I244079,I244094);
or I_21284 (I364465,I244073,I244079);
DFFARX1 I_21285 (I364465,I2595,I364312,I364304,);
not I_21286 (I364496,I244091);
nand I_21287 (I364513,I364496,I244085);
nand I_21288 (I364530,I364414,I364513);
and I_21289 (I364283,I364397,I364530);
nor I_21290 (I364561,I244091,I244073);
and I_21291 (I364578,I364397,I364561);
nor I_21292 (I364289,I364363,I364578);
DFFARX1 I_21293 (I364561,I2595,I364312,I364618,);
not I_21294 (I364626,I364618);
nor I_21295 (I364298,I364397,I364626);
or I_21296 (I364657,I364465,I244088);
nor I_21297 (I364674,I244088,I244073);
nand I_21298 (I364691,I364530,I364674);
nand I_21299 (I364708,I364657,I364691);
DFFARX1 I_21300 (I364708,I2595,I364312,I364301,);
nor I_21301 (I364739,I364674,I364431);
DFFARX1 I_21302 (I364739,I2595,I364312,I364280,);
nor I_21303 (I364770,I244088,I244079);
DFFARX1 I_21304 (I364770,I2595,I364312,I364796,);
DFFARX1 I_21305 (I364796,I2595,I364312,I364295,);
not I_21306 (I364818,I364796);
nand I_21307 (I364292,I364818,I364346);
nand I_21308 (I364286,I364818,I364448);
not I_21309 (I364890,I2602);
DFFARX1 I_21310 (I73478,I2595,I364890,I364916,);
nand I_21311 (I364924,I364916,I73481);
not I_21312 (I364941,I364924);
DFFARX1 I_21313 (I73490,I2595,I364890,I364967,);
not I_21314 (I364975,I364967);
not I_21315 (I364992,I73493);
or I_21316 (I365009,I73484,I73493);
nor I_21317 (I365026,I73484,I73493);
or I_21318 (I365043,I73496,I73484);
DFFARX1 I_21319 (I365043,I2595,I364890,I364882,);
not I_21320 (I365074,I73481);
nand I_21321 (I365091,I365074,I73487);
nand I_21322 (I365108,I364992,I365091);
and I_21323 (I364861,I364975,I365108);
nor I_21324 (I365139,I73481,I73499);
and I_21325 (I365156,I364975,I365139);
nor I_21326 (I364867,I364941,I365156);
DFFARX1 I_21327 (I365139,I2595,I364890,I365196,);
not I_21328 (I365204,I365196);
nor I_21329 (I364876,I364975,I365204);
or I_21330 (I365235,I365043,I73478);
nor I_21331 (I365252,I73478,I73496);
nand I_21332 (I365269,I365108,I365252);
nand I_21333 (I365286,I365235,I365269);
DFFARX1 I_21334 (I365286,I2595,I364890,I364879,);
nor I_21335 (I365317,I365252,I365009);
DFFARX1 I_21336 (I365317,I2595,I364890,I364858,);
nor I_21337 (I365348,I73478,I73502);
DFFARX1 I_21338 (I365348,I2595,I364890,I365374,);
DFFARX1 I_21339 (I365374,I2595,I364890,I364873,);
not I_21340 (I365396,I365374);
nand I_21341 (I364870,I365396,I364924);
nand I_21342 (I364864,I365396,I365026);
not I_21343 (I365468,I2602);
DFFARX1 I_21344 (I13967,I2595,I365468,I365494,);
nand I_21345 (I365502,I365494,I13961);
not I_21346 (I365519,I365502);
DFFARX1 I_21347 (I13979,I2595,I365468,I365545,);
not I_21348 (I365553,I365545);
not I_21349 (I365570,I13982);
or I_21350 (I365587,I13985,I13982);
nor I_21351 (I365604,I13985,I13982);
or I_21352 (I365621,I13970,I13985);
DFFARX1 I_21353 (I365621,I2595,I365468,I365460,);
not I_21354 (I365652,I13973);
nand I_21355 (I365669,I365652,I13976);
nand I_21356 (I365686,I365570,I365669);
and I_21357 (I365439,I365553,I365686);
nor I_21358 (I365717,I13973,I13964);
and I_21359 (I365734,I365553,I365717);
nor I_21360 (I365445,I365519,I365734);
DFFARX1 I_21361 (I365717,I2595,I365468,I365774,);
not I_21362 (I365782,I365774);
nor I_21363 (I365454,I365553,I365782);
or I_21364 (I365813,I365621,I13964);
nor I_21365 (I365830,I13964,I13970);
nand I_21366 (I365847,I365686,I365830);
nand I_21367 (I365864,I365813,I365847);
DFFARX1 I_21368 (I365864,I2595,I365468,I365457,);
nor I_21369 (I365895,I365830,I365587);
DFFARX1 I_21370 (I365895,I2595,I365468,I365436,);
nor I_21371 (I365926,I13964,I13961);
DFFARX1 I_21372 (I365926,I2595,I365468,I365952,);
DFFARX1 I_21373 (I365952,I2595,I365468,I365451,);
not I_21374 (I365974,I365952);
nand I_21375 (I365448,I365974,I365502);
nand I_21376 (I365442,I365974,I365604);
not I_21377 (I366046,I2602);
DFFARX1 I_21378 (I280935,I2595,I366046,I366072,);
nand I_21379 (I366080,I366072,I280956);
not I_21380 (I366097,I366080);
DFFARX1 I_21381 (I280929,I2595,I366046,I366123,);
not I_21382 (I366131,I366123);
not I_21383 (I366148,I280950);
or I_21384 (I366165,I280941,I280950);
nor I_21385 (I366182,I280941,I280950);
or I_21386 (I366199,I280944,I280941);
DFFARX1 I_21387 (I366199,I2595,I366046,I366038,);
not I_21388 (I366230,I280932);
nand I_21389 (I366247,I366230,I280947);
nand I_21390 (I366264,I366148,I366247);
and I_21391 (I366017,I366131,I366264);
nor I_21392 (I366295,I280932,I280929);
and I_21393 (I366312,I366131,I366295);
nor I_21394 (I366023,I366097,I366312);
DFFARX1 I_21395 (I366295,I2595,I366046,I366352,);
not I_21396 (I366360,I366352);
nor I_21397 (I366032,I366131,I366360);
or I_21398 (I366391,I366199,I280953);
nor I_21399 (I366408,I280953,I280944);
nand I_21400 (I366425,I366264,I366408);
nand I_21401 (I366442,I366391,I366425);
DFFARX1 I_21402 (I366442,I2595,I366046,I366035,);
nor I_21403 (I366473,I366408,I366165);
DFFARX1 I_21404 (I366473,I2595,I366046,I366014,);
nor I_21405 (I366504,I280953,I280938);
DFFARX1 I_21406 (I366504,I2595,I366046,I366530,);
DFFARX1 I_21407 (I366530,I2595,I366046,I366029,);
not I_21408 (I366552,I366530);
nand I_21409 (I366026,I366552,I366080);
nand I_21410 (I366020,I366552,I366182);
not I_21411 (I366624,I2602);
DFFARX1 I_21412 (I187072,I2595,I366624,I366650,);
nand I_21413 (I366658,I366650,I187075);
not I_21414 (I366675,I366658);
DFFARX1 I_21415 (I187087,I2595,I366624,I366701,);
not I_21416 (I366709,I366701);
not I_21417 (I366726,I187072);
or I_21418 (I366743,I187081,I187072);
nor I_21419 (I366760,I187081,I187072);
or I_21420 (I366777,I187090,I187081);
DFFARX1 I_21421 (I366777,I2595,I366624,I366616,);
not I_21422 (I366808,I187093);
nand I_21423 (I366825,I366808,I187075);
nand I_21424 (I366842,I366726,I366825);
and I_21425 (I366595,I366709,I366842);
nor I_21426 (I366873,I187093,I187078);
and I_21427 (I366890,I366709,I366873);
nor I_21428 (I366601,I366675,I366890);
DFFARX1 I_21429 (I366873,I2595,I366624,I366930,);
not I_21430 (I366938,I366930);
nor I_21431 (I366610,I366709,I366938);
or I_21432 (I366969,I366777,I187084);
nor I_21433 (I366986,I187084,I187090);
nand I_21434 (I367003,I366842,I366986);
nand I_21435 (I367020,I366969,I367003);
DFFARX1 I_21436 (I367020,I2595,I366624,I366613,);
nor I_21437 (I367051,I366986,I366743);
DFFARX1 I_21438 (I367051,I2595,I366624,I366592,);
nor I_21439 (I367082,I187084,I187096);
DFFARX1 I_21440 (I367082,I2595,I366624,I367108,);
DFFARX1 I_21441 (I367108,I2595,I366624,I366607,);
not I_21442 (I367130,I367108);
nand I_21443 (I366604,I367130,I366658);
nand I_21444 (I366598,I367130,I366760);
not I_21445 (I367202,I2602);
DFFARX1 I_21446 (I88529,I2595,I367202,I367228,);
nand I_21447 (I367236,I367228,I88550);
not I_21448 (I367253,I367236);
DFFARX1 I_21449 (I88544,I2595,I367202,I367279,);
not I_21450 (I367287,I367279);
not I_21451 (I367304,I88532);
or I_21452 (I367321,I88547,I88532);
nor I_21453 (I367338,I88547,I88532);
or I_21454 (I367355,I88538,I88547);
DFFARX1 I_21455 (I367355,I2595,I367202,I367194,);
not I_21456 (I367386,I88526);
nand I_21457 (I367403,I367386,I88523);
nand I_21458 (I367420,I367304,I367403);
and I_21459 (I367173,I367287,I367420);
nor I_21460 (I367451,I88526,I88535);
and I_21461 (I367468,I367287,I367451);
nor I_21462 (I367179,I367253,I367468);
DFFARX1 I_21463 (I367451,I2595,I367202,I367508,);
not I_21464 (I367516,I367508);
nor I_21465 (I367188,I367287,I367516);
or I_21466 (I367547,I367355,I88541);
nor I_21467 (I367564,I88541,I88538);
nand I_21468 (I367581,I367420,I367564);
nand I_21469 (I367598,I367547,I367581);
DFFARX1 I_21470 (I367598,I2595,I367202,I367191,);
nor I_21471 (I367629,I367564,I367321);
DFFARX1 I_21472 (I367629,I2595,I367202,I367170,);
nor I_21473 (I367660,I88541,I88523);
DFFARX1 I_21474 (I367660,I2595,I367202,I367686,);
DFFARX1 I_21475 (I367686,I2595,I367202,I367185,);
not I_21476 (I367708,I367686);
nand I_21477 (I367182,I367708,I367236);
nand I_21478 (I367176,I367708,I367338);
not I_21479 (I367780,I2602);
DFFARX1 I_21480 (I7963,I2595,I367780,I367806,);
nand I_21481 (I367814,I367806,I7960);
not I_21482 (I367831,I367814);
DFFARX1 I_21483 (I7981,I2595,I367780,I367857,);
not I_21484 (I367865,I367857);
not I_21485 (I367882,I7966);
or I_21486 (I367899,I7975,I7966);
nor I_21487 (I367916,I7975,I7966);
or I_21488 (I367933,I7960,I7975);
DFFARX1 I_21489 (I367933,I2595,I367780,I367772,);
not I_21490 (I367964,I7972);
nand I_21491 (I367981,I367964,I7978);
nand I_21492 (I367998,I367882,I367981);
and I_21493 (I367751,I367865,I367998);
nor I_21494 (I368029,I7972,I7966);
and I_21495 (I368046,I367865,I368029);
nor I_21496 (I367757,I367831,I368046);
DFFARX1 I_21497 (I368029,I2595,I367780,I368086,);
not I_21498 (I368094,I368086);
nor I_21499 (I367766,I367865,I368094);
or I_21500 (I368125,I367933,I7963);
nor I_21501 (I368142,I7963,I7960);
nand I_21502 (I368159,I367998,I368142);
nand I_21503 (I368176,I368125,I368159);
DFFARX1 I_21504 (I368176,I2595,I367780,I367769,);
nor I_21505 (I368207,I368142,I367899);
DFFARX1 I_21506 (I368207,I2595,I367780,I367748,);
nor I_21507 (I368238,I7963,I7969);
DFFARX1 I_21508 (I368238,I2595,I367780,I368264,);
DFFARX1 I_21509 (I368264,I2595,I367780,I367763,);
not I_21510 (I368286,I368264);
nand I_21511 (I367760,I368286,I367814);
nand I_21512 (I367754,I368286,I367916);
not I_21513 (I368358,I2602);
DFFARX1 I_21514 (I5583,I2595,I368358,I368384,);
nand I_21515 (I368392,I368384,I5580);
not I_21516 (I368409,I368392);
DFFARX1 I_21517 (I5601,I2595,I368358,I368435,);
not I_21518 (I368443,I368435);
not I_21519 (I368460,I5586);
or I_21520 (I368477,I5595,I5586);
nor I_21521 (I368494,I5595,I5586);
or I_21522 (I368511,I5580,I5595);
DFFARX1 I_21523 (I368511,I2595,I368358,I368350,);
not I_21524 (I368542,I5592);
nand I_21525 (I368559,I368542,I5598);
nand I_21526 (I368576,I368460,I368559);
and I_21527 (I368329,I368443,I368576);
nor I_21528 (I368607,I5592,I5586);
and I_21529 (I368624,I368443,I368607);
nor I_21530 (I368335,I368409,I368624);
DFFARX1 I_21531 (I368607,I2595,I368358,I368664,);
not I_21532 (I368672,I368664);
nor I_21533 (I368344,I368443,I368672);
or I_21534 (I368703,I368511,I5583);
nor I_21535 (I368720,I5583,I5580);
nand I_21536 (I368737,I368576,I368720);
nand I_21537 (I368754,I368703,I368737);
DFFARX1 I_21538 (I368754,I2595,I368358,I368347,);
nor I_21539 (I368785,I368720,I368477);
DFFARX1 I_21540 (I368785,I2595,I368358,I368326,);
nor I_21541 (I368816,I5583,I5589);
DFFARX1 I_21542 (I368816,I2595,I368358,I368842,);
DFFARX1 I_21543 (I368842,I2595,I368358,I368341,);
not I_21544 (I368864,I368842);
nand I_21545 (I368338,I368864,I368392);
nand I_21546 (I368332,I368864,I368494);
not I_21547 (I368939,I2602);
DFFARX1 I_21548 (I55033,I2595,I368939,I368965,);
nand I_21549 (I368973,I368965,I55057);
not I_21550 (I368990,I368973);
DFFARX1 I_21551 (I55045,I2595,I368939,I369016,);
not I_21552 (I369024,I369016);
nor I_21553 (I369041,I55036,I55054);
not I_21554 (I369058,I369041);
DFFARX1 I_21555 (I369058,I2595,I368939,I368925,);
or I_21556 (I369089,I55048,I55036);
DFFARX1 I_21557 (I369089,I2595,I368939,I368928,);
not I_21558 (I369120,I55036);
nor I_21559 (I369137,I369120,I55051);
nor I_21560 (I369154,I369137,I55054);
nor I_21561 (I369171,I55051,I55042);
nor I_21562 (I369188,I369024,I369171);
nor I_21563 (I368913,I368990,I369188);
not I_21564 (I369219,I369171);
nand I_21565 (I368916,I369219,I368973);
nand I_21566 (I368910,I369219,I369041);
nor I_21567 (I368907,I369171,I369154);
nor I_21568 (I369278,I55039,I55048);
not I_21569 (I369295,I369278);
DFFARX1 I_21570 (I369278,I2595,I368939,I369321,);
not I_21571 (I368931,I369321);
nor I_21572 (I369343,I55039,I55033);
DFFARX1 I_21573 (I369343,I2595,I368939,I369369,);
and I_21574 (I369377,I369369,I55036);
nor I_21575 (I369394,I369377,I369295);
DFFARX1 I_21576 (I369394,I2595,I368939,I368922,);
nor I_21577 (I369425,I369369,I369154);
DFFARX1 I_21578 (I369425,I2595,I368939,I368904,);
nor I_21579 (I368919,I369369,I369058);
not I_21580 (I369500,I2602);
DFFARX1 I_21581 (I64553,I2595,I369500,I369526,);
nand I_21582 (I369534,I369526,I64577);
not I_21583 (I369551,I369534);
DFFARX1 I_21584 (I64565,I2595,I369500,I369577,);
not I_21585 (I369585,I369577);
nor I_21586 (I369602,I64556,I64574);
not I_21587 (I369619,I369602);
DFFARX1 I_21588 (I369619,I2595,I369500,I369486,);
or I_21589 (I369650,I64568,I64556);
DFFARX1 I_21590 (I369650,I2595,I369500,I369489,);
not I_21591 (I369681,I64556);
nor I_21592 (I369698,I369681,I64571);
nor I_21593 (I369715,I369698,I64574);
nor I_21594 (I369732,I64571,I64562);
nor I_21595 (I369749,I369585,I369732);
nor I_21596 (I369474,I369551,I369749);
not I_21597 (I369780,I369732);
nand I_21598 (I369477,I369780,I369534);
nand I_21599 (I369471,I369780,I369602);
nor I_21600 (I369468,I369732,I369715);
nor I_21601 (I369839,I64559,I64568);
not I_21602 (I369856,I369839);
DFFARX1 I_21603 (I369839,I2595,I369500,I369882,);
not I_21604 (I369492,I369882);
nor I_21605 (I369904,I64559,I64553);
DFFARX1 I_21606 (I369904,I2595,I369500,I369930,);
and I_21607 (I369938,I369930,I64556);
nor I_21608 (I369955,I369938,I369856);
DFFARX1 I_21609 (I369955,I2595,I369500,I369483,);
nor I_21610 (I369986,I369930,I369715);
DFFARX1 I_21611 (I369986,I2595,I369500,I369465,);
nor I_21612 (I369480,I369930,I369619);
not I_21613 (I370061,I2602);
DFFARX1 I_21614 (I324095,I2595,I370061,I370087,);
nand I_21615 (I370095,I370087,I324092);
not I_21616 (I370112,I370095);
DFFARX1 I_21617 (I324095,I2595,I370061,I370138,);
not I_21618 (I370146,I370138);
nor I_21619 (I370163,I324113,I324107);
not I_21620 (I370180,I370163);
DFFARX1 I_21621 (I370180,I2595,I370061,I370047,);
or I_21622 (I370211,I324116,I324113);
DFFARX1 I_21623 (I370211,I2595,I370061,I370050,);
not I_21624 (I370242,I324104);
nor I_21625 (I370259,I370242,I324101);
nor I_21626 (I370276,I370259,I324107);
nor I_21627 (I370293,I324101,I324092);
nor I_21628 (I370310,I370146,I370293);
nor I_21629 (I370035,I370112,I370310);
not I_21630 (I370341,I370293);
nand I_21631 (I370038,I370341,I370095);
nand I_21632 (I370032,I370341,I370163);
nor I_21633 (I370029,I370293,I370276);
nor I_21634 (I370400,I324098,I324116);
not I_21635 (I370417,I370400);
DFFARX1 I_21636 (I370400,I2595,I370061,I370443,);
not I_21637 (I370053,I370443);
nor I_21638 (I370465,I324098,I324110);
DFFARX1 I_21639 (I370465,I2595,I370061,I370491,);
and I_21640 (I370499,I370491,I324113);
nor I_21641 (I370516,I370499,I370417);
DFFARX1 I_21642 (I370516,I2595,I370061,I370044,);
nor I_21643 (I370547,I370491,I370276);
DFFARX1 I_21644 (I370547,I2595,I370061,I370026,);
nor I_21645 (I370041,I370491,I370180);
not I_21646 (I370622,I2602);
DFFARX1 I_21647 (I105408,I2595,I370622,I370648,);
nand I_21648 (I370656,I370648,I105387);
not I_21649 (I370673,I370656);
DFFARX1 I_21650 (I105396,I2595,I370622,I370699,);
not I_21651 (I370707,I370699);
nor I_21652 (I370724,I105390,I105402);
not I_21653 (I370741,I370724);
DFFARX1 I_21654 (I370741,I2595,I370622,I370608,);
or I_21655 (I370772,I105393,I105390);
DFFARX1 I_21656 (I370772,I2595,I370622,I370611,);
not I_21657 (I370803,I105414);
nor I_21658 (I370820,I370803,I105399);
nor I_21659 (I370837,I370820,I105402);
nor I_21660 (I370854,I105399,I105387);
nor I_21661 (I370871,I370707,I370854);
nor I_21662 (I370596,I370673,I370871);
not I_21663 (I370902,I370854);
nand I_21664 (I370599,I370902,I370656);
nand I_21665 (I370593,I370902,I370724);
nor I_21666 (I370590,I370854,I370837);
nor I_21667 (I370961,I105405,I105393);
not I_21668 (I370978,I370961);
DFFARX1 I_21669 (I370961,I2595,I370622,I371004,);
not I_21670 (I370614,I371004);
nor I_21671 (I371026,I105405,I105411);
DFFARX1 I_21672 (I371026,I2595,I370622,I371052,);
and I_21673 (I371060,I371052,I105390);
nor I_21674 (I371077,I371060,I370978);
DFFARX1 I_21675 (I371077,I2595,I370622,I370605,);
nor I_21676 (I371108,I371052,I370837);
DFFARX1 I_21677 (I371108,I2595,I370622,I370587,);
nor I_21678 (I370602,I371052,I370741);
not I_21679 (I371183,I2602);
DFFARX1 I_21680 (I183625,I2595,I371183,I371209,);
DFFARX1 I_21681 (I183607,I2595,I371183,I371226,);
not I_21682 (I371234,I371226);
nor I_21683 (I371151,I371209,I371234);
DFFARX1 I_21684 (I371234,I2595,I371183,I371166,);
nor I_21685 (I371279,I183613,I183616);
and I_21686 (I371296,I371279,I183604);
nor I_21687 (I371313,I371296,I183613);
not I_21688 (I371330,I183613);
and I_21689 (I371347,I371330,I183622);
nand I_21690 (I371364,I371347,I183610);
nor I_21691 (I371381,I371330,I371364);
DFFARX1 I_21692 (I371381,I2595,I371183,I371148,);
not I_21693 (I371412,I371364);
nand I_21694 (I371429,I371234,I371412);
nand I_21695 (I371160,I371296,I371412);
DFFARX1 I_21696 (I371330,I2595,I371183,I371175,);
not I_21697 (I371474,I183607);
nor I_21698 (I371491,I371474,I183622);
nor I_21699 (I371508,I371491,I371313);
DFFARX1 I_21700 (I371508,I2595,I371183,I371172,);
not I_21701 (I371539,I371491);
DFFARX1 I_21702 (I371539,I2595,I371183,I371565,);
not I_21703 (I371573,I371565);
nor I_21704 (I371169,I371573,I371491);
nor I_21705 (I371604,I371474,I183619);
and I_21706 (I371621,I371604,I183628);
or I_21707 (I371638,I371621,I183604);
DFFARX1 I_21708 (I371638,I2595,I371183,I371664,);
not I_21709 (I371672,I371664);
nand I_21710 (I371689,I371672,I371412);
not I_21711 (I371163,I371689);
nand I_21712 (I371157,I371689,I371429);
nand I_21713 (I371154,I371672,I371296);
not I_21714 (I371778,I2602);
DFFARX1 I_21715 (I184781,I2595,I371778,I371804,);
DFFARX1 I_21716 (I184763,I2595,I371778,I371821,);
not I_21717 (I371829,I371821);
nor I_21718 (I371746,I371804,I371829);
DFFARX1 I_21719 (I371829,I2595,I371778,I371761,);
nor I_21720 (I371874,I184769,I184772);
and I_21721 (I371891,I371874,I184760);
nor I_21722 (I371908,I371891,I184769);
not I_21723 (I371925,I184769);
and I_21724 (I371942,I371925,I184778);
nand I_21725 (I371959,I371942,I184766);
nor I_21726 (I371976,I371925,I371959);
DFFARX1 I_21727 (I371976,I2595,I371778,I371743,);
not I_21728 (I372007,I371959);
nand I_21729 (I372024,I371829,I372007);
nand I_21730 (I371755,I371891,I372007);
DFFARX1 I_21731 (I371925,I2595,I371778,I371770,);
not I_21732 (I372069,I184763);
nor I_21733 (I372086,I372069,I184778);
nor I_21734 (I372103,I372086,I371908);
DFFARX1 I_21735 (I372103,I2595,I371778,I371767,);
not I_21736 (I372134,I372086);
DFFARX1 I_21737 (I372134,I2595,I371778,I372160,);
not I_21738 (I372168,I372160);
nor I_21739 (I371764,I372168,I372086);
nor I_21740 (I372199,I372069,I184775);
and I_21741 (I372216,I372199,I184784);
or I_21742 (I372233,I372216,I184760);
DFFARX1 I_21743 (I372233,I2595,I371778,I372259,);
not I_21744 (I372267,I372259);
nand I_21745 (I372284,I372267,I372007);
not I_21746 (I371758,I372284);
nand I_21747 (I371752,I372284,I372024);
nand I_21748 (I371749,I372267,I371891);
not I_21749 (I372373,I2602);
DFFARX1 I_21750 (I137177,I2595,I372373,I372399,);
DFFARX1 I_21751 (I137183,I2595,I372373,I372416,);
not I_21752 (I372424,I372416);
nor I_21753 (I372341,I372399,I372424);
DFFARX1 I_21754 (I372424,I2595,I372373,I372356,);
nor I_21755 (I372469,I137192,I137177);
and I_21756 (I372486,I372469,I137204);
nor I_21757 (I372503,I372486,I137192);
not I_21758 (I372520,I137192);
and I_21759 (I372537,I372520,I137180);
nand I_21760 (I372554,I372537,I137201);
nor I_21761 (I372571,I372520,I372554);
DFFARX1 I_21762 (I372571,I2595,I372373,I372338,);
not I_21763 (I372602,I372554);
nand I_21764 (I372619,I372424,I372602);
nand I_21765 (I372350,I372486,I372602);
DFFARX1 I_21766 (I372520,I2595,I372373,I372365,);
not I_21767 (I372664,I137189);
nor I_21768 (I372681,I372664,I137180);
nor I_21769 (I372698,I372681,I372503);
DFFARX1 I_21770 (I372698,I2595,I372373,I372362,);
not I_21771 (I372729,I372681);
DFFARX1 I_21772 (I372729,I2595,I372373,I372755,);
not I_21773 (I372763,I372755);
nor I_21774 (I372359,I372763,I372681);
nor I_21775 (I372794,I372664,I137186);
and I_21776 (I372811,I372794,I137198);
or I_21777 (I372828,I372811,I137195);
DFFARX1 I_21778 (I372828,I2595,I372373,I372854,);
not I_21779 (I372862,I372854);
nand I_21780 (I372879,I372862,I372602);
not I_21781 (I372353,I372879);
nand I_21782 (I372347,I372879,I372619);
nand I_21783 (I372344,I372862,I372486);
not I_21784 (I372968,I2602);
DFFARX1 I_21785 (I45075,I2595,I372968,I372994,);
DFFARX1 I_21786 (I45063,I2595,I372968,I373011,);
not I_21787 (I373019,I373011);
nor I_21788 (I372936,I372994,I373019);
DFFARX1 I_21789 (I373019,I2595,I372968,I372951,);
nor I_21790 (I373064,I45054,I45078);
and I_21791 (I373081,I373064,I45057);
nor I_21792 (I373098,I373081,I45054);
not I_21793 (I373115,I45054);
and I_21794 (I373132,I373115,I45060);
nand I_21795 (I373149,I373132,I45072);
nor I_21796 (I373166,I373115,I373149);
DFFARX1 I_21797 (I373166,I2595,I372968,I372933,);
not I_21798 (I373197,I373149);
nand I_21799 (I373214,I373019,I373197);
nand I_21800 (I372945,I373081,I373197);
DFFARX1 I_21801 (I373115,I2595,I372968,I372960,);
not I_21802 (I373259,I45054);
nor I_21803 (I373276,I373259,I45060);
nor I_21804 (I373293,I373276,I373098);
DFFARX1 I_21805 (I373293,I2595,I372968,I372957,);
not I_21806 (I373324,I373276);
DFFARX1 I_21807 (I373324,I2595,I372968,I373350,);
not I_21808 (I373358,I373350);
nor I_21809 (I372954,I373358,I373276);
nor I_21810 (I373389,I373259,I45057);
and I_21811 (I373406,I373389,I45066);
or I_21812 (I373423,I373406,I45069);
DFFARX1 I_21813 (I373423,I2595,I372968,I373449,);
not I_21814 (I373457,I373449);
nand I_21815 (I373474,I373457,I373197);
not I_21816 (I372948,I373474);
nand I_21817 (I372942,I373474,I373214);
nand I_21818 (I372939,I373457,I373081);
not I_21819 (I373563,I2602);
DFFARX1 I_21820 (I15560,I2595,I373563,I373589,);
DFFARX1 I_21821 (I15542,I2595,I373563,I373606,);
not I_21822 (I373614,I373606);
nor I_21823 (I373531,I373589,I373614);
DFFARX1 I_21824 (I373614,I2595,I373563,I373546,);
nor I_21825 (I373659,I15542,I15557);
and I_21826 (I373676,I373659,I15551);
nor I_21827 (I373693,I373676,I15542);
not I_21828 (I373710,I15542);
and I_21829 (I373727,I373710,I15545);
nand I_21830 (I373744,I373727,I15548);
nor I_21831 (I373761,I373710,I373744);
DFFARX1 I_21832 (I373761,I2595,I373563,I373528,);
not I_21833 (I373792,I373744);
nand I_21834 (I373809,I373614,I373792);
nand I_21835 (I373540,I373676,I373792);
DFFARX1 I_21836 (I373710,I2595,I373563,I373555,);
not I_21837 (I373854,I15554);
nor I_21838 (I373871,I373854,I15545);
nor I_21839 (I373888,I373871,I373693);
DFFARX1 I_21840 (I373888,I2595,I373563,I373552,);
not I_21841 (I373919,I373871);
DFFARX1 I_21842 (I373919,I2595,I373563,I373945,);
not I_21843 (I373953,I373945);
nor I_21844 (I373549,I373953,I373871);
nor I_21845 (I373984,I373854,I15566);
and I_21846 (I374001,I373984,I15563);
or I_21847 (I374018,I374001,I15545);
DFFARX1 I_21848 (I374018,I2595,I373563,I374044,);
not I_21849 (I374052,I374044);
nand I_21850 (I374069,I374052,I373792);
not I_21851 (I373543,I374069);
nand I_21852 (I373537,I374069,I373809);
nand I_21853 (I373534,I374052,I373676);
not I_21854 (I374158,I2602);
DFFARX1 I_21855 (I235650,I2595,I374158,I374184,);
DFFARX1 I_21856 (I235647,I2595,I374158,I374201,);
not I_21857 (I374209,I374201);
nor I_21858 (I374126,I374184,I374209);
DFFARX1 I_21859 (I374209,I2595,I374158,I374141,);
nor I_21860 (I374254,I235662,I235644);
and I_21861 (I374271,I374254,I235641);
nor I_21862 (I374288,I374271,I235662);
not I_21863 (I374305,I235662);
and I_21864 (I374322,I374305,I235647);
nand I_21865 (I374339,I374322,I235659);
nor I_21866 (I374356,I374305,I374339);
DFFARX1 I_21867 (I374356,I2595,I374158,I374123,);
not I_21868 (I374387,I374339);
nand I_21869 (I374404,I374209,I374387);
nand I_21870 (I374135,I374271,I374387);
DFFARX1 I_21871 (I374305,I2595,I374158,I374150,);
not I_21872 (I374449,I235653);
nor I_21873 (I374466,I374449,I235647);
nor I_21874 (I374483,I374466,I374288);
DFFARX1 I_21875 (I374483,I2595,I374158,I374147,);
not I_21876 (I374514,I374466);
DFFARX1 I_21877 (I374514,I2595,I374158,I374540,);
not I_21878 (I374548,I374540);
nor I_21879 (I374144,I374548,I374466);
nor I_21880 (I374579,I374449,I235641);
and I_21881 (I374596,I374579,I235656);
or I_21882 (I374613,I374596,I235644);
DFFARX1 I_21883 (I374613,I2595,I374158,I374639,);
not I_21884 (I374647,I374639);
nand I_21885 (I374664,I374647,I374387);
not I_21886 (I374138,I374664);
nand I_21887 (I374132,I374664,I374404);
nand I_21888 (I374129,I374647,I374271);
not I_21889 (I374753,I2602);
DFFARX1 I_21890 (I206167,I2595,I374753,I374779,);
DFFARX1 I_21891 (I206149,I2595,I374753,I374796,);
not I_21892 (I374804,I374796);
nor I_21893 (I374721,I374779,I374804);
DFFARX1 I_21894 (I374804,I2595,I374753,I374736,);
nor I_21895 (I374849,I206155,I206158);
and I_21896 (I374866,I374849,I206146);
nor I_21897 (I374883,I374866,I206155);
not I_21898 (I374900,I206155);
and I_21899 (I374917,I374900,I206164);
nand I_21900 (I374934,I374917,I206152);
nor I_21901 (I374951,I374900,I374934);
DFFARX1 I_21902 (I374951,I2595,I374753,I374718,);
not I_21903 (I374982,I374934);
nand I_21904 (I374999,I374804,I374982);
nand I_21905 (I374730,I374866,I374982);
DFFARX1 I_21906 (I374900,I2595,I374753,I374745,);
not I_21907 (I375044,I206149);
nor I_21908 (I375061,I375044,I206164);
nor I_21909 (I375078,I375061,I374883);
DFFARX1 I_21910 (I375078,I2595,I374753,I374742,);
not I_21911 (I375109,I375061);
DFFARX1 I_21912 (I375109,I2595,I374753,I375135,);
not I_21913 (I375143,I375135);
nor I_21914 (I374739,I375143,I375061);
nor I_21915 (I375174,I375044,I206161);
and I_21916 (I375191,I375174,I206170);
or I_21917 (I375208,I375191,I206146);
DFFARX1 I_21918 (I375208,I2595,I374753,I375234,);
not I_21919 (I375242,I375234);
nand I_21920 (I375259,I375242,I374982);
not I_21921 (I374733,I375259);
nand I_21922 (I374727,I375259,I374999);
nand I_21923 (I374724,I375242,I374866);
not I_21924 (I375348,I2602);
DFFARX1 I_21925 (I61578,I2595,I375348,I375374,);
DFFARX1 I_21926 (I61581,I2595,I375348,I375391,);
not I_21927 (I375399,I375391);
nor I_21928 (I375316,I375374,I375399);
DFFARX1 I_21929 (I375399,I2595,I375348,I375331,);
nor I_21930 (I375444,I61587,I61581);
and I_21931 (I375461,I375444,I61584);
nor I_21932 (I375478,I375461,I61587);
not I_21933 (I375495,I61587);
and I_21934 (I375512,I375495,I61578);
nand I_21935 (I375529,I375512,I61596);
nor I_21936 (I375546,I375495,I375529);
DFFARX1 I_21937 (I375546,I2595,I375348,I375313,);
not I_21938 (I375577,I375529);
nand I_21939 (I375594,I375399,I375577);
nand I_21940 (I375325,I375461,I375577);
DFFARX1 I_21941 (I375495,I2595,I375348,I375340,);
not I_21942 (I375639,I61590);
nor I_21943 (I375656,I375639,I61578);
nor I_21944 (I375673,I375656,I375478);
DFFARX1 I_21945 (I375673,I2595,I375348,I375337,);
not I_21946 (I375704,I375656);
DFFARX1 I_21947 (I375704,I2595,I375348,I375730,);
not I_21948 (I375738,I375730);
nor I_21949 (I375334,I375738,I375656);
nor I_21950 (I375769,I375639,I61593);
and I_21951 (I375786,I375769,I61599);
or I_21952 (I375803,I375786,I61602);
DFFARX1 I_21953 (I375803,I2595,I375348,I375829,);
not I_21954 (I375837,I375829);
nand I_21955 (I375854,I375837,I375577);
not I_21956 (I375328,I375854);
nand I_21957 (I375322,I375854,I375594);
nand I_21958 (I375319,I375837,I375461);
not I_21959 (I375943,I2602);
DFFARX1 I_21960 (I253803,I2595,I375943,I375969,);
DFFARX1 I_21961 (I253821,I2595,I375943,I375986,);
not I_21962 (I375994,I375986);
nor I_21963 (I375911,I375969,I375994);
DFFARX1 I_21964 (I375994,I2595,I375943,I375926,);
nor I_21965 (I376039,I253800,I253812);
and I_21966 (I376056,I376039,I253797);
nor I_21967 (I376073,I376056,I253800);
not I_21968 (I376090,I253800);
and I_21969 (I376107,I376090,I253806);
nand I_21970 (I376124,I376107,I253818);
nor I_21971 (I376141,I376090,I376124);
DFFARX1 I_21972 (I376141,I2595,I375943,I375908,);
not I_21973 (I376172,I376124);
nand I_21974 (I376189,I375994,I376172);
nand I_21975 (I375920,I376056,I376172);
DFFARX1 I_21976 (I376090,I2595,I375943,I375935,);
not I_21977 (I376234,I253809);
nor I_21978 (I376251,I376234,I253806);
nor I_21979 (I376268,I376251,I376073);
DFFARX1 I_21980 (I376268,I2595,I375943,I375932,);
not I_21981 (I376299,I376251);
DFFARX1 I_21982 (I376299,I2595,I375943,I376325,);
not I_21983 (I376333,I376325);
nor I_21984 (I375929,I376333,I376251);
nor I_21985 (I376364,I376234,I253797);
and I_21986 (I376381,I376364,I253824);
or I_21987 (I376398,I376381,I253815);
DFFARX1 I_21988 (I376398,I2595,I375943,I376424,);
not I_21989 (I376432,I376424);
nand I_21990 (I376449,I376432,I376172);
not I_21991 (I375923,I376449);
nand I_21992 (I375917,I376449,I376189);
nand I_21993 (I375914,I376432,I376056);
not I_21994 (I376538,I2602);
DFFARX1 I_21995 (I96449,I2595,I376538,I376564,);
DFFARX1 I_21996 (I96443,I2595,I376538,I376581,);
not I_21997 (I376589,I376581);
nor I_21998 (I376506,I376564,I376589);
DFFARX1 I_21999 (I376589,I2595,I376538,I376521,);
nor I_22000 (I376634,I96431,I96452);
and I_22001 (I376651,I376634,I96446);
nor I_22002 (I376668,I376651,I96431);
not I_22003 (I376685,I96431);
and I_22004 (I376702,I376685,I96428);
nand I_22005 (I376719,I376702,I96440);
nor I_22006 (I376736,I376685,I376719);
DFFARX1 I_22007 (I376736,I2595,I376538,I376503,);
not I_22008 (I376767,I376719);
nand I_22009 (I376784,I376589,I376767);
nand I_22010 (I376515,I376651,I376767);
DFFARX1 I_22011 (I376685,I2595,I376538,I376530,);
not I_22012 (I376829,I96455);
nor I_22013 (I376846,I376829,I96428);
nor I_22014 (I376863,I376846,I376668);
DFFARX1 I_22015 (I376863,I2595,I376538,I376527,);
not I_22016 (I376894,I376846);
DFFARX1 I_22017 (I376894,I2595,I376538,I376920,);
not I_22018 (I376928,I376920);
nor I_22019 (I376524,I376928,I376846);
nor I_22020 (I376959,I376829,I96437);
and I_22021 (I376976,I376959,I96434);
or I_22022 (I376993,I376976,I96428);
DFFARX1 I_22023 (I376993,I2595,I376538,I377019,);
not I_22024 (I377027,I377019);
nand I_22025 (I377044,I377027,I376767);
not I_22026 (I376518,I377044);
nand I_22027 (I376512,I377044,I376784);
nand I_22028 (I376509,I377027,I376651);
not I_22029 (I377133,I2602);
DFFARX1 I_22030 (I327563,I2595,I377133,I377159,);
DFFARX1 I_22031 (I327575,I2595,I377133,I377176,);
not I_22032 (I377184,I377176);
nor I_22033 (I377101,I377159,I377184);
DFFARX1 I_22034 (I377184,I2595,I377133,I377116,);
nor I_22035 (I377229,I327572,I327566);
and I_22036 (I377246,I377229,I327560);
nor I_22037 (I377263,I377246,I327572);
not I_22038 (I377280,I327572);
and I_22039 (I377297,I377280,I327569);
nand I_22040 (I377314,I377297,I327560);
nor I_22041 (I377331,I377280,I377314);
DFFARX1 I_22042 (I377331,I2595,I377133,I377098,);
not I_22043 (I377362,I377314);
nand I_22044 (I377379,I377184,I377362);
nand I_22045 (I377110,I377246,I377362);
DFFARX1 I_22046 (I377280,I2595,I377133,I377125,);
not I_22047 (I377424,I327584);
nor I_22048 (I377441,I377424,I327569);
nor I_22049 (I377458,I377441,I377263);
DFFARX1 I_22050 (I377458,I2595,I377133,I377122,);
not I_22051 (I377489,I377441);
DFFARX1 I_22052 (I377489,I2595,I377133,I377515,);
not I_22053 (I377523,I377515);
nor I_22054 (I377119,I377523,I377441);
nor I_22055 (I377554,I377424,I327578);
and I_22056 (I377571,I377554,I327581);
or I_22057 (I377588,I377571,I327563);
DFFARX1 I_22058 (I377588,I2595,I377133,I377614,);
not I_22059 (I377622,I377614);
nand I_22060 (I377639,I377622,I377362);
not I_22061 (I377113,I377639);
nand I_22062 (I377107,I377639,I377379);
nand I_22063 (I377104,I377622,I377246);
not I_22064 (I377728,I2602);
DFFARX1 I_22065 (I84855,I2595,I377728,I377754,);
DFFARX1 I_22066 (I84849,I2595,I377728,I377771,);
not I_22067 (I377779,I377771);
nor I_22068 (I377696,I377754,I377779);
DFFARX1 I_22069 (I377779,I2595,I377728,I377711,);
nor I_22070 (I377824,I84837,I84858);
and I_22071 (I377841,I377824,I84852);
nor I_22072 (I377858,I377841,I84837);
not I_22073 (I377875,I84837);
and I_22074 (I377892,I377875,I84834);
nand I_22075 (I377909,I377892,I84846);
nor I_22076 (I377926,I377875,I377909);
DFFARX1 I_22077 (I377926,I2595,I377728,I377693,);
not I_22078 (I377957,I377909);
nand I_22079 (I377974,I377779,I377957);
nand I_22080 (I377705,I377841,I377957);
DFFARX1 I_22081 (I377875,I2595,I377728,I377720,);
not I_22082 (I378019,I84861);
nor I_22083 (I378036,I378019,I84834);
nor I_22084 (I378053,I378036,I377858);
DFFARX1 I_22085 (I378053,I2595,I377728,I377717,);
not I_22086 (I378084,I378036);
DFFARX1 I_22087 (I378084,I2595,I377728,I378110,);
not I_22088 (I378118,I378110);
nor I_22089 (I377714,I378118,I378036);
nor I_22090 (I378149,I378019,I84843);
and I_22091 (I378166,I378149,I84840);
or I_22092 (I378183,I378166,I84834);
DFFARX1 I_22093 (I378183,I2595,I377728,I378209,);
not I_22094 (I378217,I378209);
nand I_22095 (I378234,I378217,I377957);
not I_22096 (I377708,I378234);
nand I_22097 (I377702,I378234,I377974);
nand I_22098 (I377699,I378217,I377841);
not I_22099 (I378323,I2602);
DFFARX1 I_22100 (I74073,I2595,I378323,I378349,);
DFFARX1 I_22101 (I74076,I2595,I378323,I378366,);
not I_22102 (I378374,I378366);
nor I_22103 (I378291,I378349,I378374);
DFFARX1 I_22104 (I378374,I2595,I378323,I378306,);
nor I_22105 (I378419,I74082,I74076);
and I_22106 (I378436,I378419,I74079);
nor I_22107 (I378453,I378436,I74082);
not I_22108 (I378470,I74082);
and I_22109 (I378487,I378470,I74073);
nand I_22110 (I378504,I378487,I74091);
nor I_22111 (I378521,I378470,I378504);
DFFARX1 I_22112 (I378521,I2595,I378323,I378288,);
not I_22113 (I378552,I378504);
nand I_22114 (I378569,I378374,I378552);
nand I_22115 (I378300,I378436,I378552);
DFFARX1 I_22116 (I378470,I2595,I378323,I378315,);
not I_22117 (I378614,I74085);
nor I_22118 (I378631,I378614,I74073);
nor I_22119 (I378648,I378631,I378453);
DFFARX1 I_22120 (I378648,I2595,I378323,I378312,);
not I_22121 (I378679,I378631);
DFFARX1 I_22122 (I378679,I2595,I378323,I378705,);
not I_22123 (I378713,I378705);
nor I_22124 (I378309,I378713,I378631);
nor I_22125 (I378744,I378614,I74088);
and I_22126 (I378761,I378744,I74094);
or I_22127 (I378778,I378761,I74097);
DFFARX1 I_22128 (I378778,I2595,I378323,I378804,);
not I_22129 (I378812,I378804);
nand I_22130 (I378829,I378812,I378552);
not I_22131 (I378303,I378829);
nand I_22132 (I378297,I378829,I378569);
nand I_22133 (I378294,I378812,I378436);
not I_22134 (I378918,I2602);
DFFARX1 I_22135 (I294949,I2595,I378918,I378944,);
DFFARX1 I_22136 (I294940,I2595,I378918,I378961,);
not I_22137 (I378969,I378961);
nor I_22138 (I378886,I378944,I378969);
DFFARX1 I_22139 (I378969,I2595,I378918,I378901,);
nor I_22140 (I379014,I294946,I294955);
and I_22141 (I379031,I379014,I294958);
nor I_22142 (I379048,I379031,I294946);
not I_22143 (I379065,I294946);
and I_22144 (I379082,I379065,I294937);
nand I_22145 (I379099,I379082,I294943);
nor I_22146 (I379116,I379065,I379099);
DFFARX1 I_22147 (I379116,I2595,I378918,I378883,);
not I_22148 (I379147,I379099);
nand I_22149 (I379164,I378969,I379147);
nand I_22150 (I378895,I379031,I379147);
DFFARX1 I_22151 (I379065,I2595,I378918,I378910,);
not I_22152 (I379209,I294952);
nor I_22153 (I379226,I379209,I294937);
nor I_22154 (I379243,I379226,I379048);
DFFARX1 I_22155 (I379243,I2595,I378918,I378907,);
not I_22156 (I379274,I379226);
DFFARX1 I_22157 (I379274,I2595,I378918,I379300,);
not I_22158 (I379308,I379300);
nor I_22159 (I378904,I379308,I379226);
nor I_22160 (I379339,I379209,I294937);
and I_22161 (I379356,I379339,I294940);
or I_22162 (I379373,I379356,I294943);
DFFARX1 I_22163 (I379373,I2595,I378918,I379399,);
not I_22164 (I379407,I379399);
nand I_22165 (I379424,I379407,I379147);
not I_22166 (I378898,I379424);
nand I_22167 (I378892,I379424,I379164);
nand I_22168 (I378889,I379407,I379031);
not I_22169 (I379513,I2602);
DFFARX1 I_22170 (I337967,I2595,I379513,I379539,);
DFFARX1 I_22171 (I337979,I2595,I379513,I379556,);
not I_22172 (I379564,I379556);
nor I_22173 (I379481,I379539,I379564);
DFFARX1 I_22174 (I379564,I2595,I379513,I379496,);
nor I_22175 (I379609,I337976,I337970);
and I_22176 (I379626,I379609,I337964);
nor I_22177 (I379643,I379626,I337976);
not I_22178 (I379660,I337976);
and I_22179 (I379677,I379660,I337973);
nand I_22180 (I379694,I379677,I337964);
nor I_22181 (I379711,I379660,I379694);
DFFARX1 I_22182 (I379711,I2595,I379513,I379478,);
not I_22183 (I379742,I379694);
nand I_22184 (I379759,I379564,I379742);
nand I_22185 (I379490,I379626,I379742);
DFFARX1 I_22186 (I379660,I2595,I379513,I379505,);
not I_22187 (I379804,I337988);
nor I_22188 (I379821,I379804,I337973);
nor I_22189 (I379838,I379821,I379643);
DFFARX1 I_22190 (I379838,I2595,I379513,I379502,);
not I_22191 (I379869,I379821);
DFFARX1 I_22192 (I379869,I2595,I379513,I379895,);
not I_22193 (I379903,I379895);
nor I_22194 (I379499,I379903,I379821);
nor I_22195 (I379934,I379804,I337982);
and I_22196 (I379951,I379934,I337985);
or I_22197 (I379968,I379951,I337967);
DFFARX1 I_22198 (I379968,I2595,I379513,I379994,);
not I_22199 (I380002,I379994);
nand I_22200 (I380019,I380002,I379742);
not I_22201 (I379493,I380019);
nand I_22202 (I379487,I380019,I379759);
nand I_22203 (I379484,I380002,I379626);
not I_22204 (I380108,I2602);
DFFARX1 I_22205 (I34535,I2595,I380108,I380134,);
DFFARX1 I_22206 (I34523,I2595,I380108,I380151,);
not I_22207 (I380159,I380151);
nor I_22208 (I380076,I380134,I380159);
DFFARX1 I_22209 (I380159,I2595,I380108,I380091,);
nor I_22210 (I380204,I34514,I34538);
and I_22211 (I380221,I380204,I34517);
nor I_22212 (I380238,I380221,I34514);
not I_22213 (I380255,I34514);
and I_22214 (I380272,I380255,I34520);
nand I_22215 (I380289,I380272,I34532);
nor I_22216 (I380306,I380255,I380289);
DFFARX1 I_22217 (I380306,I2595,I380108,I380073,);
not I_22218 (I380337,I380289);
nand I_22219 (I380354,I380159,I380337);
nand I_22220 (I380085,I380221,I380337);
DFFARX1 I_22221 (I380255,I2595,I380108,I380100,);
not I_22222 (I380399,I34514);
nor I_22223 (I380416,I380399,I34520);
nor I_22224 (I380433,I380416,I380238);
DFFARX1 I_22225 (I380433,I2595,I380108,I380097,);
not I_22226 (I380464,I380416);
DFFARX1 I_22227 (I380464,I2595,I380108,I380490,);
not I_22228 (I380498,I380490);
nor I_22229 (I380094,I380498,I380416);
nor I_22230 (I380529,I380399,I34517);
and I_22231 (I380546,I380529,I34526);
or I_22232 (I380563,I380546,I34529);
DFFARX1 I_22233 (I380563,I2595,I380108,I380589,);
not I_22234 (I380597,I380589);
nand I_22235 (I380614,I380597,I380337);
not I_22236 (I380088,I380614);
nand I_22237 (I380082,I380614,I380354);
nand I_22238 (I380079,I380597,I380221);
not I_22239 (I380703,I2602);
DFFARX1 I_22240 (I164551,I2595,I380703,I380729,);
DFFARX1 I_22241 (I164545,I2595,I380703,I380746,);
not I_22242 (I380754,I380746);
nor I_22243 (I380671,I380729,I380754);
DFFARX1 I_22244 (I380754,I2595,I380703,I380686,);
nor I_22245 (I380799,I164542,I164533);
and I_22246 (I380816,I380799,I164530);
nor I_22247 (I380833,I380816,I164542);
not I_22248 (I380850,I164542);
and I_22249 (I380867,I380850,I164536);
nand I_22250 (I380884,I380867,I164548);
nor I_22251 (I380901,I380850,I380884);
DFFARX1 I_22252 (I380901,I2595,I380703,I380668,);
not I_22253 (I380932,I380884);
nand I_22254 (I380949,I380754,I380932);
nand I_22255 (I380680,I380816,I380932);
DFFARX1 I_22256 (I380850,I2595,I380703,I380695,);
not I_22257 (I380994,I164554);
nor I_22258 (I381011,I380994,I164536);
nor I_22259 (I381028,I381011,I380833);
DFFARX1 I_22260 (I381028,I2595,I380703,I380692,);
not I_22261 (I381059,I381011);
DFFARX1 I_22262 (I381059,I2595,I380703,I381085,);
not I_22263 (I381093,I381085);
nor I_22264 (I380689,I381093,I381011);
nor I_22265 (I381124,I380994,I164533);
and I_22266 (I381141,I381124,I164539);
or I_22267 (I381158,I381141,I164530);
DFFARX1 I_22268 (I381158,I2595,I380703,I381184,);
not I_22269 (I381192,I381184);
nand I_22270 (I381209,I381192,I380932);
not I_22271 (I380683,I381209);
nand I_22272 (I380677,I381209,I380949);
nand I_22273 (I380674,I381192,I380816);
not I_22274 (I381298,I2602);
DFFARX1 I_22275 (I252511,I2595,I381298,I381324,);
DFFARX1 I_22276 (I252529,I2595,I381298,I381341,);
not I_22277 (I381349,I381341);
nor I_22278 (I381266,I381324,I381349);
DFFARX1 I_22279 (I381349,I2595,I381298,I381281,);
nor I_22280 (I381394,I252508,I252520);
and I_22281 (I381411,I381394,I252505);
nor I_22282 (I381428,I381411,I252508);
not I_22283 (I381445,I252508);
and I_22284 (I381462,I381445,I252514);
nand I_22285 (I381479,I381462,I252526);
nor I_22286 (I381496,I381445,I381479);
DFFARX1 I_22287 (I381496,I2595,I381298,I381263,);
not I_22288 (I381527,I381479);
nand I_22289 (I381544,I381349,I381527);
nand I_22290 (I381275,I381411,I381527);
DFFARX1 I_22291 (I381445,I2595,I381298,I381290,);
not I_22292 (I381589,I252517);
nor I_22293 (I381606,I381589,I252514);
nor I_22294 (I381623,I381606,I381428);
DFFARX1 I_22295 (I381623,I2595,I381298,I381287,);
not I_22296 (I381654,I381606);
DFFARX1 I_22297 (I381654,I2595,I381298,I381680,);
not I_22298 (I381688,I381680);
nor I_22299 (I381284,I381688,I381606);
nor I_22300 (I381719,I381589,I252505);
and I_22301 (I381736,I381719,I252532);
or I_22302 (I381753,I381736,I252523);
DFFARX1 I_22303 (I381753,I2595,I381298,I381779,);
not I_22304 (I381787,I381779);
nand I_22305 (I381804,I381787,I381527);
not I_22306 (I381278,I381804);
nand I_22307 (I381272,I381804,I381544);
nand I_22308 (I381269,I381787,I381411);
not I_22309 (I381893,I2602);
DFFARX1 I_22310 (I288687,I2595,I381893,I381919,);
DFFARX1 I_22311 (I288705,I2595,I381893,I381936,);
not I_22312 (I381944,I381936);
nor I_22313 (I381861,I381919,I381944);
DFFARX1 I_22314 (I381944,I2595,I381893,I381876,);
nor I_22315 (I381989,I288684,I288696);
and I_22316 (I382006,I381989,I288681);
nor I_22317 (I382023,I382006,I288684);
not I_22318 (I382040,I288684);
and I_22319 (I382057,I382040,I288690);
nand I_22320 (I382074,I382057,I288702);
nor I_22321 (I382091,I382040,I382074);
DFFARX1 I_22322 (I382091,I2595,I381893,I381858,);
not I_22323 (I382122,I382074);
nand I_22324 (I382139,I381944,I382122);
nand I_22325 (I381870,I382006,I382122);
DFFARX1 I_22326 (I382040,I2595,I381893,I381885,);
not I_22327 (I382184,I288693);
nor I_22328 (I382201,I382184,I288690);
nor I_22329 (I382218,I382201,I382023);
DFFARX1 I_22330 (I382218,I2595,I381893,I381882,);
not I_22331 (I382249,I382201);
DFFARX1 I_22332 (I382249,I2595,I381893,I382275,);
not I_22333 (I382283,I382275);
nor I_22334 (I381879,I382283,I382201);
nor I_22335 (I382314,I382184,I288681);
and I_22336 (I382331,I382314,I288708);
or I_22337 (I382348,I382331,I288699);
DFFARX1 I_22338 (I382348,I2595,I381893,I382374,);
not I_22339 (I382382,I382374);
nand I_22340 (I382399,I382382,I382122);
not I_22341 (I381873,I382399);
nand I_22342 (I381867,I382399,I382139);
nand I_22343 (I381864,I382382,I382006);
not I_22344 (I382488,I2602);
DFFARX1 I_22345 (I11871,I2595,I382488,I382514,);
DFFARX1 I_22346 (I11853,I2595,I382488,I382531,);
not I_22347 (I382539,I382531);
nor I_22348 (I382456,I382514,I382539);
DFFARX1 I_22349 (I382539,I2595,I382488,I382471,);
nor I_22350 (I382584,I11853,I11868);
and I_22351 (I382601,I382584,I11862);
nor I_22352 (I382618,I382601,I11853);
not I_22353 (I382635,I11853);
and I_22354 (I382652,I382635,I11856);
nand I_22355 (I382669,I382652,I11859);
nor I_22356 (I382686,I382635,I382669);
DFFARX1 I_22357 (I382686,I2595,I382488,I382453,);
not I_22358 (I382717,I382669);
nand I_22359 (I382734,I382539,I382717);
nand I_22360 (I382465,I382601,I382717);
DFFARX1 I_22361 (I382635,I2595,I382488,I382480,);
not I_22362 (I382779,I11865);
nor I_22363 (I382796,I382779,I11856);
nor I_22364 (I382813,I382796,I382618);
DFFARX1 I_22365 (I382813,I2595,I382488,I382477,);
not I_22366 (I382844,I382796);
DFFARX1 I_22367 (I382844,I2595,I382488,I382870,);
not I_22368 (I382878,I382870);
nor I_22369 (I382474,I382878,I382796);
nor I_22370 (I382909,I382779,I11877);
and I_22371 (I382926,I382909,I11874);
or I_22372 (I382943,I382926,I11856);
DFFARX1 I_22373 (I382943,I2595,I382488,I382969,);
not I_22374 (I382977,I382969);
nand I_22375 (I382994,I382977,I382717);
not I_22376 (I382468,I382994);
nand I_22377 (I382462,I382994,I382734);
nand I_22378 (I382459,I382977,I382601);
not I_22379 (I383083,I2602);
DFFARX1 I_22380 (I51463,I2595,I383083,I383109,);
DFFARX1 I_22381 (I51466,I2595,I383083,I383126,);
not I_22382 (I383134,I383126);
nor I_22383 (I383051,I383109,I383134);
DFFARX1 I_22384 (I383134,I2595,I383083,I383066,);
nor I_22385 (I383179,I51472,I51466);
and I_22386 (I383196,I383179,I51469);
nor I_22387 (I383213,I383196,I51472);
not I_22388 (I383230,I51472);
and I_22389 (I383247,I383230,I51463);
nand I_22390 (I383264,I383247,I51481);
nor I_22391 (I383281,I383230,I383264);
DFFARX1 I_22392 (I383281,I2595,I383083,I383048,);
not I_22393 (I383312,I383264);
nand I_22394 (I383329,I383134,I383312);
nand I_22395 (I383060,I383196,I383312);
DFFARX1 I_22396 (I383230,I2595,I383083,I383075,);
not I_22397 (I383374,I51475);
nor I_22398 (I383391,I383374,I51463);
nor I_22399 (I383408,I383391,I383213);
DFFARX1 I_22400 (I383408,I2595,I383083,I383072,);
not I_22401 (I383439,I383391);
DFFARX1 I_22402 (I383439,I2595,I383083,I383465,);
not I_22403 (I383473,I383465);
nor I_22404 (I383069,I383473,I383391);
nor I_22405 (I383504,I383374,I51478);
and I_22406 (I383521,I383504,I51484);
or I_22407 (I383538,I383521,I51487);
DFFARX1 I_22408 (I383538,I2595,I383083,I383564,);
not I_22409 (I383572,I383564);
nand I_22410 (I383589,I383572,I383312);
not I_22411 (I383063,I383589);
nand I_22412 (I383057,I383589,I383329);
nand I_22413 (I383054,I383572,I383196);
not I_22414 (I383678,I2602);
DFFARX1 I_22415 (I349694,I2595,I383678,I383704,);
DFFARX1 I_22416 (I349697,I2595,I383678,I383721,);
not I_22417 (I383729,I383721);
nor I_22418 (I383646,I383704,I383729);
DFFARX1 I_22419 (I383729,I2595,I383678,I383661,);
nor I_22420 (I383774,I349697,I349712);
and I_22421 (I383791,I383774,I349706);
nor I_22422 (I383808,I383791,I349697);
not I_22423 (I383825,I349697);
and I_22424 (I383842,I383825,I349715);
nand I_22425 (I383859,I383842,I349703);
nor I_22426 (I383876,I383825,I383859);
DFFARX1 I_22427 (I383876,I2595,I383678,I383643,);
not I_22428 (I383907,I383859);
nand I_22429 (I383924,I383729,I383907);
nand I_22430 (I383655,I383791,I383907);
DFFARX1 I_22431 (I383825,I2595,I383678,I383670,);
not I_22432 (I383969,I349709);
nor I_22433 (I383986,I383969,I349715);
nor I_22434 (I384003,I383986,I383808);
DFFARX1 I_22435 (I384003,I2595,I383678,I383667,);
not I_22436 (I384034,I383986);
DFFARX1 I_22437 (I384034,I2595,I383678,I384060,);
not I_22438 (I384068,I384060);
nor I_22439 (I383664,I384068,I383986);
nor I_22440 (I384099,I383969,I349694);
and I_22441 (I384116,I384099,I349718);
or I_22442 (I384133,I384116,I349700);
DFFARX1 I_22443 (I384133,I2595,I383678,I384159,);
not I_22444 (I384167,I384159);
nand I_22445 (I384184,I384167,I383907);
not I_22446 (I383658,I384184);
nand I_22447 (I383652,I384184,I383924);
nand I_22448 (I383649,I384167,I383791);
not I_22449 (I384273,I2602);
DFFARX1 I_22450 (I165707,I2595,I384273,I384299,);
DFFARX1 I_22451 (I165701,I2595,I384273,I384316,);
not I_22452 (I384324,I384316);
nor I_22453 (I384241,I384299,I384324);
DFFARX1 I_22454 (I384324,I2595,I384273,I384256,);
nor I_22455 (I384369,I165698,I165689);
and I_22456 (I384386,I384369,I165686);
nor I_22457 (I384403,I384386,I165698);
not I_22458 (I384420,I165698);
and I_22459 (I384437,I384420,I165692);
nand I_22460 (I384454,I384437,I165704);
nor I_22461 (I384471,I384420,I384454);
DFFARX1 I_22462 (I384471,I2595,I384273,I384238,);
not I_22463 (I384502,I384454);
nand I_22464 (I384519,I384324,I384502);
nand I_22465 (I384250,I384386,I384502);
DFFARX1 I_22466 (I384420,I2595,I384273,I384265,);
not I_22467 (I384564,I165710);
nor I_22468 (I384581,I384564,I165692);
nor I_22469 (I384598,I384581,I384403);
DFFARX1 I_22470 (I384598,I2595,I384273,I384262,);
not I_22471 (I384629,I384581);
DFFARX1 I_22472 (I384629,I2595,I384273,I384655,);
not I_22473 (I384663,I384655);
nor I_22474 (I384259,I384663,I384581);
nor I_22475 (I384694,I384564,I165689);
and I_22476 (I384711,I384694,I165695);
or I_22477 (I384728,I384711,I165686);
DFFARX1 I_22478 (I384728,I2595,I384273,I384754,);
not I_22479 (I384762,I384754);
nand I_22480 (I384779,I384762,I384502);
not I_22481 (I384253,I384779);
nand I_22482 (I384247,I384779,I384519);
nand I_22483 (I384244,I384762,I384386);
not I_22484 (I384868,I2602);
DFFARX1 I_22485 (I360830,I2595,I384868,I384894,);
DFFARX1 I_22486 (I360821,I2595,I384868,I384911,);
not I_22487 (I384919,I384911);
nor I_22488 (I384836,I384894,I384919);
DFFARX1 I_22489 (I384919,I2595,I384868,I384851,);
nor I_22490 (I384964,I360812,I360827);
and I_22491 (I384981,I384964,I360815);
nor I_22492 (I384998,I384981,I360812);
not I_22493 (I385015,I360812);
and I_22494 (I385032,I385015,I360818);
nand I_22495 (I385049,I385032,I360836);
nor I_22496 (I385066,I385015,I385049);
DFFARX1 I_22497 (I385066,I2595,I384868,I384833,);
not I_22498 (I385097,I385049);
nand I_22499 (I385114,I384919,I385097);
nand I_22500 (I384845,I384981,I385097);
DFFARX1 I_22501 (I385015,I2595,I384868,I384860,);
not I_22502 (I385159,I360812);
nor I_22503 (I385176,I385159,I360818);
nor I_22504 (I385193,I385176,I384998);
DFFARX1 I_22505 (I385193,I2595,I384868,I384857,);
not I_22506 (I385224,I385176);
DFFARX1 I_22507 (I385224,I2595,I384868,I385250,);
not I_22508 (I385258,I385250);
nor I_22509 (I384854,I385258,I385176);
nor I_22510 (I385289,I385159,I360815);
and I_22511 (I385306,I385289,I360824);
or I_22512 (I385323,I385306,I360833);
DFFARX1 I_22513 (I385323,I2595,I384868,I385349,);
not I_22514 (I385357,I385349);
nand I_22515 (I385374,I385357,I385097);
not I_22516 (I384848,I385374);
nand I_22517 (I384842,I385374,I385114);
nand I_22518 (I384839,I385357,I384981);
not I_22519 (I385463,I2602);
DFFARX1 I_22520 (I227553,I2595,I385463,I385489,);
DFFARX1 I_22521 (I227535,I2595,I385463,I385506,);
not I_22522 (I385514,I385506);
nor I_22523 (I385431,I385489,I385514);
DFFARX1 I_22524 (I385514,I2595,I385463,I385446,);
nor I_22525 (I385559,I227541,I227544);
and I_22526 (I385576,I385559,I227532);
nor I_22527 (I385593,I385576,I227541);
not I_22528 (I385610,I227541);
and I_22529 (I385627,I385610,I227550);
nand I_22530 (I385644,I385627,I227538);
nor I_22531 (I385661,I385610,I385644);
DFFARX1 I_22532 (I385661,I2595,I385463,I385428,);
not I_22533 (I385692,I385644);
nand I_22534 (I385709,I385514,I385692);
nand I_22535 (I385440,I385576,I385692);
DFFARX1 I_22536 (I385610,I2595,I385463,I385455,);
not I_22537 (I385754,I227535);
nor I_22538 (I385771,I385754,I227550);
nor I_22539 (I385788,I385771,I385593);
DFFARX1 I_22540 (I385788,I2595,I385463,I385452,);
not I_22541 (I385819,I385771);
DFFARX1 I_22542 (I385819,I2595,I385463,I385845,);
not I_22543 (I385853,I385845);
nor I_22544 (I385449,I385853,I385771);
nor I_22545 (I385884,I385754,I227547);
and I_22546 (I385901,I385884,I227556);
or I_22547 (I385918,I385901,I227532);
DFFARX1 I_22548 (I385918,I2595,I385463,I385944,);
not I_22549 (I385952,I385944);
nand I_22550 (I385969,I385952,I385692);
not I_22551 (I385443,I385969);
nand I_22552 (I385437,I385969,I385709);
nand I_22553 (I385434,I385952,I385576);
not I_22554 (I386058,I2602);
DFFARX1 I_22555 (I173221,I2595,I386058,I386084,);
DFFARX1 I_22556 (I173215,I2595,I386058,I386101,);
not I_22557 (I386109,I386101);
nor I_22558 (I386026,I386084,I386109);
DFFARX1 I_22559 (I386109,I2595,I386058,I386041,);
nor I_22560 (I386154,I173212,I173203);
and I_22561 (I386171,I386154,I173200);
nor I_22562 (I386188,I386171,I173212);
not I_22563 (I386205,I173212);
and I_22564 (I386222,I386205,I173206);
nand I_22565 (I386239,I386222,I173218);
nor I_22566 (I386256,I386205,I386239);
DFFARX1 I_22567 (I386256,I2595,I386058,I386023,);
not I_22568 (I386287,I386239);
nand I_22569 (I386304,I386109,I386287);
nand I_22570 (I386035,I386171,I386287);
DFFARX1 I_22571 (I386205,I2595,I386058,I386050,);
not I_22572 (I386349,I173224);
nor I_22573 (I386366,I386349,I173206);
nor I_22574 (I386383,I386366,I386188);
DFFARX1 I_22575 (I386383,I2595,I386058,I386047,);
not I_22576 (I386414,I386366);
DFFARX1 I_22577 (I386414,I2595,I386058,I386440,);
not I_22578 (I386448,I386440);
nor I_22579 (I386044,I386448,I386366);
nor I_22580 (I386479,I386349,I173203);
and I_22581 (I386496,I386479,I173209);
or I_22582 (I386513,I386496,I173200);
DFFARX1 I_22583 (I386513,I2595,I386058,I386539,);
not I_22584 (I386547,I386539);
nand I_22585 (I386564,I386547,I386287);
not I_22586 (I386038,I386564);
nand I_22587 (I386032,I386564,I386304);
nand I_22588 (I386029,I386547,I386171);
not I_22589 (I386653,I2602);
DFFARX1 I_22590 (I367766,I2595,I386653,I386679,);
DFFARX1 I_22591 (I367757,I2595,I386653,I386696,);
not I_22592 (I386704,I386696);
nor I_22593 (I386621,I386679,I386704);
DFFARX1 I_22594 (I386704,I2595,I386653,I386636,);
nor I_22595 (I386749,I367748,I367763);
and I_22596 (I386766,I386749,I367751);
nor I_22597 (I386783,I386766,I367748);
not I_22598 (I386800,I367748);
and I_22599 (I386817,I386800,I367754);
nand I_22600 (I386834,I386817,I367772);
nor I_22601 (I386851,I386800,I386834);
DFFARX1 I_22602 (I386851,I2595,I386653,I386618,);
not I_22603 (I386882,I386834);
nand I_22604 (I386899,I386704,I386882);
nand I_22605 (I386630,I386766,I386882);
DFFARX1 I_22606 (I386800,I2595,I386653,I386645,);
not I_22607 (I386944,I367748);
nor I_22608 (I386961,I386944,I367754);
nor I_22609 (I386978,I386961,I386783);
DFFARX1 I_22610 (I386978,I2595,I386653,I386642,);
not I_22611 (I387009,I386961);
DFFARX1 I_22612 (I387009,I2595,I386653,I387035,);
not I_22613 (I387043,I387035);
nor I_22614 (I386639,I387043,I386961);
nor I_22615 (I387074,I386944,I367751);
and I_22616 (I387091,I387074,I367760);
or I_22617 (I387108,I387091,I367769);
DFFARX1 I_22618 (I387108,I2595,I386653,I387134,);
not I_22619 (I387142,I387134);
nand I_22620 (I387159,I387142,I386882);
not I_22621 (I386633,I387159);
nand I_22622 (I386627,I387159,I386899);
nand I_22623 (I386624,I387142,I386766);
not I_22624 (I387248,I2602);
DFFARX1 I_22625 (I361986,I2595,I387248,I387274,);
DFFARX1 I_22626 (I361977,I2595,I387248,I387291,);
not I_22627 (I387299,I387291);
nor I_22628 (I387216,I387274,I387299);
DFFARX1 I_22629 (I387299,I2595,I387248,I387231,);
nor I_22630 (I387344,I361968,I361983);
and I_22631 (I387361,I387344,I361971);
nor I_22632 (I387378,I387361,I361968);
not I_22633 (I387395,I361968);
and I_22634 (I387412,I387395,I361974);
nand I_22635 (I387429,I387412,I361992);
nor I_22636 (I387446,I387395,I387429);
DFFARX1 I_22637 (I387446,I2595,I387248,I387213,);
not I_22638 (I387477,I387429);
nand I_22639 (I387494,I387299,I387477);
nand I_22640 (I387225,I387361,I387477);
DFFARX1 I_22641 (I387395,I2595,I387248,I387240,);
not I_22642 (I387539,I361968);
nor I_22643 (I387556,I387539,I361974);
nor I_22644 (I387573,I387556,I387378);
DFFARX1 I_22645 (I387573,I2595,I387248,I387237,);
not I_22646 (I387604,I387556);
DFFARX1 I_22647 (I387604,I2595,I387248,I387630,);
not I_22648 (I387638,I387630);
nor I_22649 (I387234,I387638,I387556);
nor I_22650 (I387669,I387539,I361971);
and I_22651 (I387686,I387669,I361980);
or I_22652 (I387703,I387686,I361989);
DFFARX1 I_22653 (I387703,I2595,I387248,I387729,);
not I_22654 (I387737,I387729);
nand I_22655 (I387754,I387737,I387477);
not I_22656 (I387228,I387754);
nand I_22657 (I387222,I387754,I387494);
nand I_22658 (I387219,I387737,I387361);
not I_22659 (I387843,I2602);
DFFARX1 I_22660 (I19249,I2595,I387843,I387869,);
DFFARX1 I_22661 (I19231,I2595,I387843,I387886,);
not I_22662 (I387894,I387886);
nor I_22663 (I387811,I387869,I387894);
DFFARX1 I_22664 (I387894,I2595,I387843,I387826,);
nor I_22665 (I387939,I19231,I19246);
and I_22666 (I387956,I387939,I19240);
nor I_22667 (I387973,I387956,I19231);
not I_22668 (I387990,I19231);
and I_22669 (I388007,I387990,I19234);
nand I_22670 (I388024,I388007,I19237);
nor I_22671 (I388041,I387990,I388024);
DFFARX1 I_22672 (I388041,I2595,I387843,I387808,);
not I_22673 (I388072,I388024);
nand I_22674 (I388089,I387894,I388072);
nand I_22675 (I387820,I387956,I388072);
DFFARX1 I_22676 (I387990,I2595,I387843,I387835,);
not I_22677 (I388134,I19243);
nor I_22678 (I388151,I388134,I19234);
nor I_22679 (I388168,I388151,I387973);
DFFARX1 I_22680 (I388168,I2595,I387843,I387832,);
not I_22681 (I388199,I388151);
DFFARX1 I_22682 (I388199,I2595,I387843,I388225,);
not I_22683 (I388233,I388225);
nor I_22684 (I387829,I388233,I388151);
nor I_22685 (I388264,I388134,I19255);
and I_22686 (I388281,I388264,I19252);
or I_22687 (I388298,I388281,I19234);
DFFARX1 I_22688 (I388298,I2595,I387843,I388324,);
not I_22689 (I388332,I388324);
nand I_22690 (I388349,I388332,I388072);
not I_22691 (I387823,I388349);
nand I_22692 (I387817,I388349,I388089);
nand I_22693 (I387814,I388332,I387956);
not I_22694 (I388438,I2602);
DFFARX1 I_22695 (I297193,I2595,I388438,I388464,);
DFFARX1 I_22696 (I297184,I2595,I388438,I388481,);
not I_22697 (I388489,I388481);
nor I_22698 (I388406,I388464,I388489);
DFFARX1 I_22699 (I388489,I2595,I388438,I388421,);
nor I_22700 (I388534,I297190,I297199);
and I_22701 (I388551,I388534,I297202);
nor I_22702 (I388568,I388551,I297190);
not I_22703 (I388585,I297190);
and I_22704 (I388602,I388585,I297181);
nand I_22705 (I388619,I388602,I297187);
nor I_22706 (I388636,I388585,I388619);
DFFARX1 I_22707 (I388636,I2595,I388438,I388403,);
not I_22708 (I388667,I388619);
nand I_22709 (I388684,I388489,I388667);
nand I_22710 (I388415,I388551,I388667);
DFFARX1 I_22711 (I388585,I2595,I388438,I388430,);
not I_22712 (I388729,I297196);
nor I_22713 (I388746,I388729,I297181);
nor I_22714 (I388763,I388746,I388568);
DFFARX1 I_22715 (I388763,I2595,I388438,I388427,);
not I_22716 (I388794,I388746);
DFFARX1 I_22717 (I388794,I2595,I388438,I388820,);
not I_22718 (I388828,I388820);
nor I_22719 (I388424,I388828,I388746);
nor I_22720 (I388859,I388729,I297181);
and I_22721 (I388876,I388859,I297184);
or I_22722 (I388893,I388876,I297187);
DFFARX1 I_22723 (I388893,I2595,I388438,I388919,);
not I_22724 (I388927,I388919);
nand I_22725 (I388944,I388927,I388667);
not I_22726 (I388418,I388944);
nand I_22727 (I388412,I388944,I388684);
nand I_22728 (I388409,I388927,I388551);
not I_22729 (I389033,I2602);
DFFARX1 I_22730 (I180157,I2595,I389033,I389059,);
DFFARX1 I_22731 (I180151,I2595,I389033,I389076,);
not I_22732 (I389084,I389076);
nor I_22733 (I389001,I389059,I389084);
DFFARX1 I_22734 (I389084,I2595,I389033,I389016,);
nor I_22735 (I389129,I180148,I180139);
and I_22736 (I389146,I389129,I180136);
nor I_22737 (I389163,I389146,I180148);
not I_22738 (I389180,I180148);
and I_22739 (I389197,I389180,I180142);
nand I_22740 (I389214,I389197,I180154);
nor I_22741 (I389231,I389180,I389214);
DFFARX1 I_22742 (I389231,I2595,I389033,I388998,);
not I_22743 (I389262,I389214);
nand I_22744 (I389279,I389084,I389262);
nand I_22745 (I389010,I389146,I389262);
DFFARX1 I_22746 (I389180,I2595,I389033,I389025,);
not I_22747 (I389324,I180160);
nor I_22748 (I389341,I389324,I180142);
nor I_22749 (I389358,I389341,I389163);
DFFARX1 I_22750 (I389358,I2595,I389033,I389022,);
not I_22751 (I389389,I389341);
DFFARX1 I_22752 (I389389,I2595,I389033,I389415,);
not I_22753 (I389423,I389415);
nor I_22754 (I389019,I389423,I389341);
nor I_22755 (I389454,I389324,I180139);
and I_22756 (I389471,I389454,I180145);
or I_22757 (I389488,I389471,I180136);
DFFARX1 I_22758 (I389488,I2595,I389033,I389514,);
not I_22759 (I389522,I389514);
nand I_22760 (I389539,I389522,I389262);
not I_22761 (I389013,I389539);
nand I_22762 (I389007,I389539,I389279);
nand I_22763 (I389004,I389522,I389146);
not I_22764 (I389628,I2602);
DFFARX1 I_22765 (I169753,I2595,I389628,I389654,);
DFFARX1 I_22766 (I169747,I2595,I389628,I389671,);
not I_22767 (I389679,I389671);
nor I_22768 (I389596,I389654,I389679);
DFFARX1 I_22769 (I389679,I2595,I389628,I389611,);
nor I_22770 (I389724,I169744,I169735);
and I_22771 (I389741,I389724,I169732);
nor I_22772 (I389758,I389741,I169744);
not I_22773 (I389775,I169744);
and I_22774 (I389792,I389775,I169738);
nand I_22775 (I389809,I389792,I169750);
nor I_22776 (I389826,I389775,I389809);
DFFARX1 I_22777 (I389826,I2595,I389628,I389593,);
not I_22778 (I389857,I389809);
nand I_22779 (I389874,I389679,I389857);
nand I_22780 (I389605,I389741,I389857);
DFFARX1 I_22781 (I389775,I2595,I389628,I389620,);
not I_22782 (I389919,I169756);
nor I_22783 (I389936,I389919,I169738);
nor I_22784 (I389953,I389936,I389758);
DFFARX1 I_22785 (I389953,I2595,I389628,I389617,);
not I_22786 (I389984,I389936);
DFFARX1 I_22787 (I389984,I2595,I389628,I390010,);
not I_22788 (I390018,I390010);
nor I_22789 (I389614,I390018,I389936);
nor I_22790 (I390049,I389919,I169735);
and I_22791 (I390066,I390049,I169741);
or I_22792 (I390083,I390066,I169732);
DFFARX1 I_22793 (I390083,I2595,I389628,I390109,);
not I_22794 (I390117,I390109);
nand I_22795 (I390134,I390117,I389857);
not I_22796 (I389608,I390134);
nand I_22797 (I389602,I390134,I389874);
nand I_22798 (I389599,I390117,I389741);
not I_22799 (I390223,I2602);
DFFARX1 I_22800 (I229853,I2595,I390223,I390249,);
DFFARX1 I_22801 (I229850,I2595,I390223,I390266,);
not I_22802 (I390274,I390266);
nor I_22803 (I390191,I390249,I390274);
DFFARX1 I_22804 (I390274,I2595,I390223,I390206,);
nor I_22805 (I390319,I229865,I229847);
and I_22806 (I390336,I390319,I229844);
nor I_22807 (I390353,I390336,I229865);
not I_22808 (I390370,I229865);
and I_22809 (I390387,I390370,I229850);
nand I_22810 (I390404,I390387,I229862);
nor I_22811 (I390421,I390370,I390404);
DFFARX1 I_22812 (I390421,I2595,I390223,I390188,);
not I_22813 (I390452,I390404);
nand I_22814 (I390469,I390274,I390452);
nand I_22815 (I390200,I390336,I390452);
DFFARX1 I_22816 (I390370,I2595,I390223,I390215,);
not I_22817 (I390514,I229856);
nor I_22818 (I390531,I390514,I229850);
nor I_22819 (I390548,I390531,I390353);
DFFARX1 I_22820 (I390548,I2595,I390223,I390212,);
not I_22821 (I390579,I390531);
DFFARX1 I_22822 (I390579,I2595,I390223,I390605,);
not I_22823 (I390613,I390605);
nor I_22824 (I390209,I390613,I390531);
nor I_22825 (I390644,I390514,I229844);
and I_22826 (I390661,I390644,I229859);
or I_22827 (I390678,I390661,I229847);
DFFARX1 I_22828 (I390678,I2595,I390223,I390704,);
not I_22829 (I390712,I390704);
nand I_22830 (I390729,I390712,I390452);
not I_22831 (I390203,I390729);
nand I_22832 (I390197,I390729,I390469);
nand I_22833 (I390194,I390712,I390336);
not I_22834 (I390818,I2602);
DFFARX1 I_22835 (I139353,I2595,I390818,I390844,);
DFFARX1 I_22836 (I139359,I2595,I390818,I390861,);
not I_22837 (I390869,I390861);
nor I_22838 (I390786,I390844,I390869);
DFFARX1 I_22839 (I390869,I2595,I390818,I390801,);
nor I_22840 (I390914,I139368,I139353);
and I_22841 (I390931,I390914,I139380);
nor I_22842 (I390948,I390931,I139368);
not I_22843 (I390965,I139368);
and I_22844 (I390982,I390965,I139356);
nand I_22845 (I390999,I390982,I139377);
nor I_22846 (I391016,I390965,I390999);
DFFARX1 I_22847 (I391016,I2595,I390818,I390783,);
not I_22848 (I391047,I390999);
nand I_22849 (I391064,I390869,I391047);
nand I_22850 (I390795,I390931,I391047);
DFFARX1 I_22851 (I390965,I2595,I390818,I390810,);
not I_22852 (I391109,I139365);
nor I_22853 (I391126,I391109,I139356);
nor I_22854 (I391143,I391126,I390948);
DFFARX1 I_22855 (I391143,I2595,I390818,I390807,);
not I_22856 (I391174,I391126);
DFFARX1 I_22857 (I391174,I2595,I390818,I391200,);
not I_22858 (I391208,I391200);
nor I_22859 (I390804,I391208,I391126);
nor I_22860 (I391239,I391109,I139362);
and I_22861 (I391256,I391239,I139374);
or I_22862 (I391273,I391256,I139371);
DFFARX1 I_22863 (I391273,I2595,I390818,I391299,);
not I_22864 (I391307,I391299);
nand I_22865 (I391324,I391307,I391047);
not I_22866 (I390798,I391324);
nand I_22867 (I390792,I391324,I391064);
nand I_22868 (I390789,I391307,I390931);
not I_22869 (I391413,I2602);
DFFARX1 I_22870 (I59793,I2595,I391413,I391439,);
DFFARX1 I_22871 (I59796,I2595,I391413,I391456,);
not I_22872 (I391464,I391456);
nor I_22873 (I391381,I391439,I391464);
DFFARX1 I_22874 (I391464,I2595,I391413,I391396,);
nor I_22875 (I391509,I59802,I59796);
and I_22876 (I391526,I391509,I59799);
nor I_22877 (I391543,I391526,I59802);
not I_22878 (I391560,I59802);
and I_22879 (I391577,I391560,I59793);
nand I_22880 (I391594,I391577,I59811);
nor I_22881 (I391611,I391560,I391594);
DFFARX1 I_22882 (I391611,I2595,I391413,I391378,);
not I_22883 (I391642,I391594);
nand I_22884 (I391659,I391464,I391642);
nand I_22885 (I391390,I391526,I391642);
DFFARX1 I_22886 (I391560,I2595,I391413,I391405,);
not I_22887 (I391704,I59805);
nor I_22888 (I391721,I391704,I59793);
nor I_22889 (I391738,I391721,I391543);
DFFARX1 I_22890 (I391738,I2595,I391413,I391402,);
not I_22891 (I391769,I391721);
DFFARX1 I_22892 (I391769,I2595,I391413,I391795,);
not I_22893 (I391803,I391795);
nor I_22894 (I391399,I391803,I391721);
nor I_22895 (I391834,I391704,I59808);
and I_22896 (I391851,I391834,I59814);
or I_22897 (I391868,I391851,I59817);
DFFARX1 I_22898 (I391868,I2595,I391413,I391894,);
not I_22899 (I391902,I391894);
nand I_22900 (I391919,I391902,I391642);
not I_22901 (I391393,I391919);
nand I_22902 (I391387,I391919,I391659);
nand I_22903 (I391384,I391902,I391526);
not I_22904 (I392008,I2602);
DFFARX1 I_22905 (I87490,I2595,I392008,I392034,);
DFFARX1 I_22906 (I87484,I2595,I392008,I392051,);
not I_22907 (I392059,I392051);
nor I_22908 (I391976,I392034,I392059);
DFFARX1 I_22909 (I392059,I2595,I392008,I391991,);
nor I_22910 (I392104,I87472,I87493);
and I_22911 (I392121,I392104,I87487);
nor I_22912 (I392138,I392121,I87472);
not I_22913 (I392155,I87472);
and I_22914 (I392172,I392155,I87469);
nand I_22915 (I392189,I392172,I87481);
nor I_22916 (I392206,I392155,I392189);
DFFARX1 I_22917 (I392206,I2595,I392008,I391973,);
not I_22918 (I392237,I392189);
nand I_22919 (I392254,I392059,I392237);
nand I_22920 (I391985,I392121,I392237);
DFFARX1 I_22921 (I392155,I2595,I392008,I392000,);
not I_22922 (I392299,I87496);
nor I_22923 (I392316,I392299,I87469);
nor I_22924 (I392333,I392316,I392138);
DFFARX1 I_22925 (I392333,I2595,I392008,I391997,);
not I_22926 (I392364,I392316);
DFFARX1 I_22927 (I392364,I2595,I392008,I392390,);
not I_22928 (I392398,I392390);
nor I_22929 (I391994,I392398,I392316);
nor I_22930 (I392429,I392299,I87478);
and I_22931 (I392446,I392429,I87475);
or I_22932 (I392463,I392446,I87469);
DFFARX1 I_22933 (I392463,I2595,I392008,I392489,);
not I_22934 (I392497,I392489);
nand I_22935 (I392514,I392497,I392237);
not I_22936 (I391988,I392514);
nand I_22937 (I391982,I392514,I392254);
nand I_22938 (I391979,I392497,I392121);
not I_22939 (I392603,I2602);
DFFARX1 I_22940 (I8558,I2595,I392603,I392629,);
DFFARX1 I_22941 (I8555,I2595,I392603,I392646,);
not I_22942 (I392654,I392646);
nor I_22943 (I392571,I392629,I392654);
DFFARX1 I_22944 (I392654,I2595,I392603,I392586,);
nor I_22945 (I392699,I8573,I8570);
and I_22946 (I392716,I392699,I8561);
nor I_22947 (I392733,I392716,I8573);
not I_22948 (I392750,I8573);
and I_22949 (I392767,I392750,I8558);
nand I_22950 (I392784,I392767,I8567);
nor I_22951 (I392801,I392750,I392784);
DFFARX1 I_22952 (I392801,I2595,I392603,I392568,);
not I_22953 (I392832,I392784);
nand I_22954 (I392849,I392654,I392832);
nand I_22955 (I392580,I392716,I392832);
DFFARX1 I_22956 (I392750,I2595,I392603,I392595,);
not I_22957 (I392894,I8576);
nor I_22958 (I392911,I392894,I8558);
nor I_22959 (I392928,I392911,I392733);
DFFARX1 I_22960 (I392928,I2595,I392603,I392592,);
not I_22961 (I392959,I392911);
DFFARX1 I_22962 (I392959,I2595,I392603,I392985,);
not I_22963 (I392993,I392985);
nor I_22964 (I392589,I392993,I392911);
nor I_22965 (I393024,I392894,I8555);
and I_22966 (I393041,I393024,I8561);
or I_22967 (I393058,I393041,I8564);
DFFARX1 I_22968 (I393058,I2595,I392603,I393084,);
not I_22969 (I393092,I393084);
nand I_22970 (I393109,I393092,I392832);
not I_22971 (I392583,I393109);
nand I_22972 (I392577,I393109,I392849);
nand I_22973 (I392574,I393092,I392716);
endmodule


