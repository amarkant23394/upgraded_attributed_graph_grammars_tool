module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_8,blif_reset_net_1_r_8,G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_8,blif_reset_net_1_r_8;
output G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8;
wire G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_452_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10,N3_2_l_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10,n_431_0_l_8,n8_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8;
DFFARX1 I_0(n4_1_r_10,blif_clk_net_1_r_8,n8_8,G42_1_r_10,);
nor I_1(n_572_1_r_10,n26_10,n3_10);
nand I_2(n_573_1_r_10,n16_10,n18_10);
nand I_3(n_549_1_r_10,n19_10,n20_10);
nor I_4(n_452_1_r_10,n25_10,n21_10);
nor I_5(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_6(N3_2_r_10,blif_clk_net_1_r_8,n8_8,G199_2_r_10,);
DFFARX1 I_7(G199_4_l_10,blif_clk_net_1_r_8,n8_8,ACVQN2_3_r_10,);
nor I_8(n_266_and_0_3_r_10,n17_10,n13_10);
and I_9(N3_2_l_10,IN_6_2_l_10,n23_10);
DFFARX1 I_10(N3_2_l_10,blif_clk_net_1_r_8,n8_8,n25_10,);
not I_11(n16_10,n25_10);
DFFARX1 I_12(IN_1_3_l_10,blif_clk_net_1_r_8,n8_8,n26_10,);
DFFARX1 I_13(IN_2_3_l_10,blif_clk_net_1_r_8,n8_8,ACVQN1_3_l_10,);
and I_14(N1_4_l_10,IN_6_4_l_10,n24_10);
DFFARX1 I_15(N1_4_l_10,blif_clk_net_1_r_8,n8_8,G199_4_l_10,);
DFFARX1 I_16(IN_3_4_l_10,blif_clk_net_1_r_8,n8_8,n27_10,);
not I_17(n17_10,n27_10);
nor I_18(n4_1_r_10,n27_10,n21_10);
nor I_19(N3_2_r_10,n16_10,n22_10);
not I_20(n3_10,n18_10);
DFFARX1 I_21(n3_10,blif_clk_net_1_r_8,n8_8,n13_internal_10,);
not I_22(n13_10,n13_internal_10);
nand I_23(n18_10,IN_4_3_l_10,ACVQN1_3_l_10);
not I_24(n19_10,n_452_1_r_10);
nand I_25(n20_10,n16_10,n26_10);
nor I_26(n21_10,IN_1_2_l_10,IN_3_2_l_10);
and I_27(n22_10,n26_10,n21_10);
nand I_28(n23_10,IN_2_2_l_10,IN_3_2_l_10);
nand I_29(n24_10,IN_1_4_l_10,IN_2_4_l_10);
DFFARX1 I_30(n4_1_r_8,blif_clk_net_1_r_8,n8_8,G42_1_r_8,);
nor I_31(n_572_1_r_8,n39_8,n23_8);
and I_32(n_549_1_r_8,n38_8,n23_8);
nand I_33(n_569_1_r_8,n38_8,n24_8);
nor I_34(n_452_1_r_8,n25_8,n26_8);
nor I_35(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_36(N3_2_r_8,blif_clk_net_1_r_8,n8_8,G199_2_r_8,);
DFFARX1 I_37(N1_4_r_8,blif_clk_net_1_r_8,n8_8,G199_4_r_8,);
DFFARX1 I_38(G78_0_l_8,blif_clk_net_1_r_8,n8_8,G214_4_r_8,);
or I_39(n_431_0_l_8,n29_8,G199_2_r_10);
not I_40(n8_8,blif_reset_net_1_r_8);
DFFARX1 I_41(n_431_0_l_8,blif_clk_net_1_r_8,n8_8,G78_0_l_8,);
not I_42(n19_8,G78_0_l_8);
DFFARX1 I_43(n_573_1_r_10,blif_clk_net_1_r_8,n8_8,n39_8,);
not I_44(n22_8,n39_8);
DFFARX1 I_45(n_573_1_r_10,blif_clk_net_1_r_8,n8_8,n38_8,);
nor I_46(n4_1_r_8,G78_0_l_8,n33_8);
nor I_47(N3_2_r_8,n22_8,n35_8);
nor I_48(N1_4_r_8,n27_8,n37_8);
nand I_49(n23_8,n32_8,G42_1_r_10);
not I_50(n24_8,n23_8);
nand I_51(n25_8,n36_8,ACVQN2_3_r_10);
nand I_52(n26_8,n27_8,n28_8);
nor I_53(n27_8,n31_8,n_549_1_r_10);
not I_54(n28_8,n_42_2_r_10);
and I_55(n29_8,n30_8,n_572_1_r_10);
nor I_56(n30_8,n31_8,G42_1_r_10);
not I_57(n31_8,n_266_and_0_3_r_10);
and I_58(n32_8,n28_8,n_549_1_r_10);
nand I_59(n33_8,n28_8,n34_8);
not I_60(n34_8,n25_8);
nor I_61(n35_8,n34_8,n_42_2_r_10);
not I_62(n36_8,n_572_1_r_10);
nor I_63(n37_8,n19_8,n38_8);
endmodule


