module test_I3314(I2815,I2668,I2234,I1294,I1301,I3314);
input I2815,I2668,I2234,I1294,I1301;
output I3314;
wire I3263,I2548,I2583,I1902,I2203,I2569,I2962,I2945,I2832;
not I_0(I3263,I2569);
nor I_1(I3314,I3263,I2548);
DFFARX1 I_2(I2945,I1294,I2583,,,I2548,);
not I_3(I2583,I1301);
and I_4(I1902,I2234,I2203);
DFFARX1 I_5(I1294,,,I2203,);
nand I_6(I2569,I2832,I2962);
nor I_7(I2962,I2945,I2668);
DFFARX1 I_8(I1902,I1294,I2583,,,I2945,);
DFFARX1 I_9(I2815,I1294,I2583,,,I2832,);
endmodule


