module test_I2215(I1271,I1231,I1343,I2215);
input I1271,I1231,I1343;
output I2215;
wire I2198;
and I_0(I2215,I2198,I1271);
nand I_1(I2198,I1343,I1231);
endmodule


