module test_I9909(I1477,I1470,I9909);
input I1477,I1470;
output I9909;
wire I8216,I8623,I9816,I8705,I8193,I9491;
not I_0(I8216,I1477);
DFFARX1 I_1(I1470,I8216,,,I8623,);
DFFARX1 I_2(I8193,I1470,I9491,,,I9816,);
DFFARX1 I_3(I8623,I1470,I8216,,,I8705,);
not I_4(I9909,I9816);
not I_5(I8193,I8705);
not I_6(I9491,I1477);
endmodule


