module test_I12619(I1477,I12619);
input I1477;
output I12619;
wire ;
not I_0(I12619,I1477);
endmodule


