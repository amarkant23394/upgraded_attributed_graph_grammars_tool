module test_I8199(I1477,I5743,I1470,I5731,I8315,I8199);
input I1477,I5743,I1470,I5731,I8315;
output I8199;
wire I8770,I8674,I8640,I8216,I8753,I8623,I8657,I8736;
or I_0(I8770,I8753,I8674);
and I_1(I8674,I8623,I8657);
not I_2(I8640,I8623);
not I_3(I8216,I1477);
not I_4(I8753,I8736);
DFFARX1 I_5(I8770,I1470,I8216,,,I8199,);
DFFARX1 I_6(I5743,I1470,I8216,,,I8623,);
nor I_7(I8657,I8315,I8640);
DFFARX1 I_8(I5731,I1470,I8216,,,I8736,);
endmodule


