module test_I10862(I9672,I1477,I1470,I9771,I9525,I10862);
input I9672,I1477,I1470,I9771,I9525;
output I10862;
wire I9542,I9720,I9816,I8705,I9483,I10845,I9459,I9453,I9737,I9689,I8193,I10828,I9491;
DFFARX1 I_0(I9525,I1470,I9491,,,I9542,);
and I_1(I10862,I10845,I9453);
not I_2(I9720,I9689);
DFFARX1 I_3(I8193,I1470,I9491,,,I9816,);
DFFARX1 I_4(I1470,,,I8705,);
nor I_5(I9483,I9816,I9542);
nor I_6(I10845,I10828,I9483);
nand I_7(I9459,I9771,I9737);
nand I_8(I9453,I9816,I9720);
nor I_9(I9737,I9720);
DFFARX1 I_10(I9672,I1470,I9491,,,I9689,);
not I_11(I8193,I8705);
not I_12(I10828,I9459);
not I_13(I9491,I1477);
endmodule


