module test_I3430(I2600,I2583,I1902,I1937,I1908,I1294,I2457,I3430);
input I2600,I2583,I1902,I1937,I1908,I1294,I2457;
output I3430;
wire I2668,I2733,I1914,I2557,I2651,I3413,I2566,I2945,I2702;
nand I_0(I2668,I2651,I1914);
not I_1(I2733,I2702);
DFFARX1 I_2(I2457,I1294,I1937,,,I1914,);
nand I_3(I2557,I2668,I2733);
nor I_4(I2651,I2600,I1908);
not I_5(I3413,I2566);
nor I_6(I3430,I3413,I2557);
not I_7(I2566,I2945);
DFFARX1 I_8(I1902,I1294,I2583,,,I2945,);
not I_9(I2702,I1908);
endmodule


