module test_I8836(I6893,I6992,I1477,I7026,I1470,I7221,I8879,I7492,I8836);
input I6893,I6992,I1477,I7026,I1470,I7221,I8879,I7492;
output I8836;
wire I9320,I6884,I6875,I6896,I9303,I9210,I9179,I8862,I8930,I6907,I8947;
not I_0(I9320,I9303);
DFFARX1 I_1(I7492,I1470,I6907,,,I6884,);
DFFARX1 I_2(I7221,I1470,I6907,,,I6875,);
nor I_3(I6896,I6992,I7026);
nand I_4(I8836,I9320,I9210);
DFFARX1 I_5(I6875,I1470,I8862,,,I9303,);
nor I_6(I9210,I9179,I8947);
DFFARX1 I_7(I6896,I1470,I8862,,,I9179,);
not I_8(I8862,I1477);
nor I_9(I8930,I8879,I6893);
not I_10(I6907,I1477);
nand I_11(I8947,I8930,I6884);
endmodule


