module test_I8011(I1477,I6843,I1470,I6363,I6705,I8011);
input I1477,I6843,I1470,I6363,I6705;
output I8011;
wire I6297,I6321,I7652,I7570,I7587,I6380,I7994,I6318,I6329,I6300,I7977,I7669,I6657;
DFFARX1 I_0(I6843,I1470,I6329,,,I6297,);
nand I_1(I6321,I6705,I6657);
nor I_2(I7652,I7587,I6297);
nor I_3(I8011,I7669,I7994);
not I_4(I7570,I1477);
not I_5(I7587,I6300);
DFFARX1 I_6(I6363,I1470,I6329,,,I6380,);
not I_7(I7994,I7977);
not I_8(I6318,I6380);
not I_9(I6329,I1477);
DFFARX1 I_10(I1470,I6329,,,I6300,);
DFFARX1 I_11(I6321,I1470,I7570,,,I7977,);
nand I_12(I7669,I7652,I6318);
nor I_13(I6657,I6380);
endmodule


