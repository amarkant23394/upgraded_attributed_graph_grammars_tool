module test_I4418(I2810,I3124,I1477,I1470,I2980,I4418);
input I2810,I3124,I1477,I1470,I2980;
output I4418;
wire I4147,I2727,I2963,I4164,I4401,I4308,I4181,I2739,I2748,I2736,I3983;
nor I_0(I4418,I4181,I4401);
nand I_1(I4147,I2739,I2736);
nand I_2(I2727,I2810,I3124);
DFFARX1 I_3(I1470,,,I2963,);
and I_4(I4164,I4147,I2748);
not I_5(I4401,I4308);
DFFARX1 I_6(I2727,I1470,I3983,,,I4308,);
DFFARX1 I_7(I4164,I1470,I3983,,,I4181,);
nor I_8(I2739,I2980);
or I_9(I2748,I2980,I2963);
DFFARX1 I_10(I1470,,,I2736,);
not I_11(I3983,I1477);
endmodule


