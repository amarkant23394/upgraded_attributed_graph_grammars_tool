module test_I3280(I2897,I2234,I2849,I1294,I1301,I3280);
input I2897,I2234,I2849,I1294,I1301;
output I3280;
wire I3103,I3168,I2548,I2560,I2583,I1902,I2203,I2945,I2914,I3086;
not I_0(I3103,I3086);
or I_1(I3168,I3103,I2914);
DFFARX1 I_2(I2945,I1294,I2583,,,I2548,);
DFFARX1 I_3(I3168,I1294,I2583,,,I2560,);
not I_4(I2583,I1301);
and I_5(I1902,I2234,I2203);
DFFARX1 I_6(I1294,,,I2203,);
nor I_7(I3280,I2548,I2560);
DFFARX1 I_8(I1902,I1294,I2583,,,I2945,);
and I_9(I2914,I2897,I2849);
DFFARX1 I_10(I1294,I2583,,,I3086,);
endmodule


