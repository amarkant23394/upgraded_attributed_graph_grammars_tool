module test_I5204(I1477,I3504,I3685,I1492,I1832,I1470,I5204);
input I1477,I3504,I3685,I1492,I1832,I1470;
output I5204;
wire I1486,I3521,I3637,I1495,I3747,I1483,I3388,I3846,I5122,I1518,I3620,I5187,I3380,I1880,I3453,I3350,I3353,I3555,I1501;
DFFARX1 I_0(I1832,I1470,I1518,,,I1486,);
nor I_1(I3521,I3504,I1495);
DFFARX1 I_2(I3620,I1470,I3388,,,I3637,);
DFFARX1 I_3(I1470,I1518,,,I1495,);
DFFARX1 I_4(I1470,I3388,,,I3747,);
DFFARX1 I_5(I1880,I1470,I1518,,,I1483,);
not I_6(I3388,I1477);
nor I_7(I3846,I3747,I3555);
not I_8(I5122,I3350);
nand I_9(I5204,I5187,I3353);
not I_10(I1518,I1477);
nor I_11(I3620,I1492,I1483);
nor I_12(I5187,I5122,I3380);
nand I_13(I3380,I3521,I3846);
DFFARX1 I_14(I1470,I1518,,,I1880,);
nor I_15(I3453,I1486,I1501);
DFFARX1 I_16(I3685,I1470,I3388,,,I3350,);
and I_17(I3353,I3453,I3637);
DFFARX1 I_18(I1470,I3388,,,I3555,);
not I_19(I1501,I1880);
endmodule


