module test_I16205(I14667,I14856,I1477,I1470,I16205);
input I14667,I14856,I1477,I1470;
output I16205;
wire I14338,I16356,I16257,I14341,I16291,I16240,I16274,I14356,I14537,I16404,I14370,I14332;
DFFARX1 I_0(I1470,I14370,,,I14338,);
DFFARX1 I_1(I14356,I1470,I16240,,,I16356,);
nand I_2(I16257,I14341,I14338);
DFFARX1 I_3(I1470,I14370,,,I14341,);
DFFARX1 I_4(I16274,I1470,I16240,,,I16291,);
not I_5(I16240,I1477);
and I_6(I16274,I16257,I14332);
nand I_7(I14356,I14667,I14856);
and I_8(I16205,I16291,I16404);
DFFARX1 I_9(I1470,I14370,,,I14537,);
DFFARX1 I_10(I16356,I1470,I16240,,,I16404,);
not I_11(I14370,I1477);
DFFARX1 I_12(I14537,I1470,I14370,,,I14332,);
endmodule


