module test_I4506(I1477,I4708,I1470,I2678,I2158,I4506);
input I1477,I4708,I1470,I2678,I2158;
output I4506;
wire I2181,I4544,I4869,I2149,I2345,I4742,I4725,I4773,I2695;
not I_0(I2181,I1477);
not I_1(I4544,I1477);
nand I_2(I4506,I4869,I4773);
DFFARX1 I_3(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_4(I2695,I1470,I2181,,,I2149,);
DFFARX1 I_5(I1470,I2181,,,I2345,);
DFFARX1 I_6(I4725,I1470,I4544,,,I4742,);
and I_7(I4725,I4708,I2158);
not I_8(I4773,I4742);
and I_9(I2695,I2345,I2678);
endmodule


