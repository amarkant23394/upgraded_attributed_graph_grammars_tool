module test_I14537(I13680,I1477,I1470,I13508,I13296,I14537);
input I13680,I1477,I1470,I13508,I13296;
output I14537;
wire I13697,I13330,I13180,I13197,I13168,I14503,I14520,I13174,I14370;
or I_0(I13697,I13296,I13680);
DFFARX1 I_1(I1470,I13197,,,I13330,);
not I_2(I13180,I13508);
not I_3(I13197,I1477);
not I_4(I13168,I13330);
nand I_5(I14503,I13180,I13168);
and I_6(I14520,I14503,I13174);
DFFARX1 I_7(I13697,I1470,I13197,,,I13174,);
DFFARX1 I_8(I14520,I1470,I14370,,,I14537,);
not I_9(I14370,I1477);
endmodule


