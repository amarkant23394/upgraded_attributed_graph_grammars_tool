module test_I3388(I1477,I3388);
input I1477;
output I3388;
wire ;
not I_0(I3388,I1477);
endmodule


