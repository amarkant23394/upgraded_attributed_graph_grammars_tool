module test_I3766(I2668,I1902,I1294,I3379,I2702,I1301,I3766);
input I2668,I1902,I1294,I3379,I2702,I1301;
output I3766;
wire I3263,I2583,I2945,I3732,I3698,I2572,I3749,I3396,I2962,I2832,I3246,I3622,I2569,I2566,I3715,I3543;
not I_0(I3263,I2569);
not I_1(I2583,I1301);
or I_2(I3766,I3543,I3749);
DFFARX1 I_3(I1902,I1294,I2583,,,I2945,);
nor I_4(I3732,I3715,I3396);
DFFARX1 I_5(I1294,I3246,,,I3698,);
nor I_6(I2572,I2668,I2702);
and I_7(I3749,I3622,I3732);
not I_8(I3396,I3379);
nor I_9(I2962,I2945,I2668);
DFFARX1 I_10(I1294,I2583,,,I2832,);
not I_11(I3246,I1301);
DFFARX1 I_12(I2572,I1294,I3246,,,I3622,);
nand I_13(I2569,I2832,I2962);
not I_14(I2566,I2945);
not I_15(I3715,I3698);
nand I_16(I3543,I3263,I2566);
endmodule


