module test_I12476(I7550,I1477,I7535,I1470,I12476);
input I7550,I1477,I7535,I1470;
output I12476;
wire I10349,I7538,I10332,I10038,I10041,I12349,I12425,I10020,I12106,I11973,I12442,I10120,I12123,I12459;
and I_0(I10349,I10332,I7550);
DFFARX1 I_1(I1470,,,I7538,);
DFFARX1 I_2(I1470,,,I10332,);
and I_3(I12476,I12349,I12459);
nand I_4(I10038,I10349);
nor I_5(I10041,I10349,I10120);
DFFARX1 I_6(I10041,I1470,I11973,,,I12349,);
DFFARX1 I_7(I10038,I1470,I11973,,,I12425,);
DFFARX1 I_8(I1470,,,I10020,);
not I_9(I12106,I10020);
not I_10(I11973,I1477);
not I_11(I12442,I12425);
nor I_12(I10120,I7538,I7535);
not I_13(I12123,I12106);
nor I_14(I12459,I12442,I12123);
endmodule


