module test_I4790(I1477,I4708,I1470,I1239,I2158,I4790);
input I1477,I4708,I1470,I1239,I2158;
output I4790;
wire I2181,I4544,I4674,I2155,I4742,I4725,I2633,I4773;
not I_0(I2181,I1477);
not I_1(I4544,I1477);
DFFARX1 I_2(I2155,I1470,I4544,,,I4674,);
DFFARX1 I_3(I2633,I1470,I2181,,,I2155,);
DFFARX1 I_4(I4725,I1470,I4544,,,I4742,);
and I_5(I4725,I4708,I2158);
nor I_6(I4790,I4674,I4773);
DFFARX1 I_7(I1239,I1470,I2181,,,I2633,);
not I_8(I4773,I4742);
endmodule


