module test_final(IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_3,blif_reset_net_1_r_3,G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3);
input IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_3,blif_reset_net_1_r_3;
output G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3;
wire G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_452_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9,N3_2_l_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9,n4_1_l_3,n9_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3;
DFFARX1 I_0(n4_1_r_9,blif_clk_net_1_r_3,n9_3,G42_1_r_9,);
nor I_1(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_2(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_3(n_549_1_r_9,n17_9,n18_9);
or I_4(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_5(n_452_1_r_9,n26_9,n25_9);
nor I_6(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_7(N3_2_r_9,blif_clk_net_1_r_3,n9_3,G199_2_r_9,);
DFFARX1 I_8(N1_4_r_9,blif_clk_net_1_r_3,n9_3,G199_4_r_9,);
DFFARX1 I_9(n_42_2_l_9,blif_clk_net_1_r_3,n9_3,G214_4_r_9,);
and I_10(N3_2_l_9,IN_6_2_l_9,n22_9);
DFFARX1 I_11(N3_2_l_9,blif_clk_net_1_r_3,n9_3,n27_9,);
not I_12(n16_9,n27_9);
DFFARX1 I_13(IN_1_3_l_9,blif_clk_net_1_r_3,n9_3,n26_9,);
not I_14(n15_9,n26_9);
DFFARX1 I_15(IN_2_3_l_9,blif_clk_net_1_r_3,n9_3,n29_internal_9,);
not I_16(n29_9,n29_internal_9);
and I_17(N1_4_l_9,IN_6_4_l_9,n24_9);
DFFARX1 I_18(N1_4_l_9,blif_clk_net_1_r_3,n9_3,n25_9,);
DFFARX1 I_19(IN_3_4_l_9,blif_clk_net_1_r_3,n9_3,n28_internal_9,);
not I_20(n28_9,n28_internal_9);
nor I_21(n4_1_r_9,n27_9,n26_9);
nor I_22(N3_2_r_9,n15_9,n21_9);
nor I_23(N1_4_r_9,n16_9,n21_9);
nor I_24(n_42_2_l_9,IN_1_2_l_9,IN_3_2_l_9);
not I_25(n17_9,n_452_1_r_9);
nand I_26(n18_9,n27_9,n15_9);
nor I_27(n19_9,n29_9,n20_9);
not I_28(n20_9,IN_4_3_l_9);
and I_29(n21_9,IN_4_3_l_9,n23_9);
nand I_30(n22_9,IN_2_2_l_9,IN_3_2_l_9);
nor I_31(n23_9,n29_9,n28_9);
nand I_32(n24_9,IN_1_4_l_9,IN_2_4_l_9);
DFFARX1 I_33(n4_1_r_3,blif_clk_net_1_r_3,n9_3,G42_1_r_3,);
nor I_34(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_35(n_573_1_r_3,n26_3,n27_3);
nor I_36(n_549_1_r_3,n40_3,n32_3);
nand I_37(n_569_1_r_3,n27_3,n31_3);
and I_38(n_452_1_r_3,n26_3,G214_4_r_9);
nor I_39(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_40(N3_2_r_3,blif_clk_net_1_r_3,n9_3,G199_2_r_3,);
DFFARX1 I_41(n_572_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_3,);
nor I_42(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_43(n4_1_l_3,n_573_1_r_9,G214_4_r_9);
not I_44(n9_3,blif_reset_net_1_r_3);
DFFARX1 I_45(n4_1_l_3,blif_clk_net_1_r_3,n9_3,G42_1_l_3,);
not I_46(n22_3,G42_1_l_3);
DFFARX1 I_47(G199_4_r_9,blif_clk_net_1_r_3,n9_3,n40_3,);
DFFARX1 I_48(G42_1_r_9,blif_clk_net_1_r_3,n9_3,n25_internal_3,);
not I_49(n25_3,n25_internal_3);
nor I_50(n4_1_r_3,n40_3,n36_3);
nor I_51(N3_2_r_3,n26_3,n37_3);
nor I_52(n_572_1_l_3,n_572_1_r_9,n_573_1_r_9);
DFFARX1 I_53(G42_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN1_3_r_3,);
nor I_54(n26_3,n_549_1_r_9,n_569_1_r_9);
not I_55(n27_3,G42_1_r_9);
nor I_56(n28_3,n29_3,G42_1_r_9);
nor I_57(n29_3,n30_3,n_572_1_r_9);
not I_58(n30_3,G199_2_r_9);
nor I_59(n31_3,n40_3,n_569_1_r_9);
nor I_60(n32_3,n25_3,n33_3);
nand I_61(n33_3,n22_3,n_42_2_r_9);
or I_62(n34_3,G42_1_r_9,n_569_1_r_9);
nand I_63(n35_3,ACVQN1_3_r_3,n_42_2_r_9);
nor I_64(n36_3,n_549_1_r_9,G214_4_r_9);
nor I_65(n37_3,n38_3,n39_3);
not I_66(n38_3,n_572_1_l_3);
nand I_67(n39_3,n27_3,n30_3);
endmodule


