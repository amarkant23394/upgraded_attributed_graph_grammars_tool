module test_I2551(I1316,I2005,I1294,I2070,I1988,I1301,I2488,I2551);
input I1316,I2005,I1294,I2070,I1988,I1301,I2488;
output I2551;
wire I2897,I2600,I1911,I2344,I2583,I2313,I2022,I1923;
nand I_0(I2897,I2600,I1923);
not I_1(I2600,I1911);
nand I_2(I1911,I2070,I2488);
DFFARX1 I_3(I2897,I1294,I2583,,,I2551,);
nor I_4(I2344,I2313,I1988);
not I_5(I2583,I1301);
DFFARX1 I_6(I1294,,,I2313,);
nand I_7(I2022,I2005,I1316);
nand I_8(I1923,I2022,I2344);
endmodule


