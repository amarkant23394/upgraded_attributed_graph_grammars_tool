module test_final(IN_1_1_l,IN_2_1_l,IN_3_1_l,G18_7_l,G15_7_l,IN_1_7_l,IN_4_7_l,IN_5_7_l,IN_7_7_l,IN_9_7_l,IN_10_7_l,IN_1_10_l,IN_2_10_l,IN_3_10_l,IN_4_10_l,blif_clk_net_8_r,blif_reset_net_8_r,N1371_0_r,N1508_0_r,N6147_2_r,N6147_3_r,N1372_4_r,N1508_4_r,N1507_6_r,N1508_6_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r);
input IN_1_1_l,IN_2_1_l,IN_3_1_l,G18_7_l,G15_7_l,IN_1_7_l,IN_4_7_l,IN_5_7_l,IN_7_7_l,IN_9_7_l,IN_10_7_l,IN_1_10_l,IN_2_10_l,IN_3_10_l,IN_4_10_l,blif_clk_net_8_r,blif_reset_net_8_r;
output N1371_0_r,N1508_0_r,N6147_2_r,N6147_3_r,N1372_4_r,N1508_4_r,N1507_6_r,N1508_6_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r;
wire N1372_1_l,N1508_1_l,n4_1_l,G42_7_l,n_87_7_l,n_572_7_l,n_573_7_l,n_549_7_l,n_569_7_l,n_452_7_l,n4_7_l,n7_7_l,N1372_10_l,N1508_10_l,n5_10_l,n6_10_l,n3_0_r,n4_0_r,n5_2_r,n6_2_r,N6138_2_r,n7_2_r,n3_3_r,N6138_3_r,n6_4_r,n7_4_r,n8_4_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,N3_8_r,n1_8_r,n3_8_r,N6150_9_r,n3_9_r;
not I_0(N1372_1_l,n4_1_l);
nor I_1(N1508_1_l,IN_3_1_l,n4_1_l);
nand I_2(n4_1_l,IN_1_1_l,IN_2_1_l);
DFFARX1 I_3(n4_7_l,blif_clk_net_8_r,n1_8_r,G42_7_l,);
not I_4(n_87_7_l,G15_7_l);
nor I_5(n_572_7_l,G15_7_l,IN_7_7_l);
or I_6(n_573_7_l,IN_5_7_l,IN_9_7_l);
nor I_7(n_549_7_l,IN_10_7_l,n7_7_l);
or I_8(n_569_7_l,IN_9_7_l,IN_10_7_l);
nor I_9(n_452_7_l,G18_7_l,IN_5_7_l);
nor I_10(n4_7_l,G18_7_l,IN_1_7_l);
and I_11(n7_7_l,IN_4_7_l,n_87_7_l);
not I_12(N1372_10_l,n6_10_l);
nor I_13(N1508_10_l,n5_10_l,n6_10_l);
nor I_14(n5_10_l,IN_3_10_l,IN_4_10_l);
nand I_15(n6_10_l,IN_1_10_l,IN_2_10_l);
nor I_16(N1371_0_r,n4_0_r,N1508_10_l);
nor I_17(N1508_0_r,n3_0_r,n4_0_r);
nor I_18(n3_0_r,n_572_7_l,N1508_1_l);
not I_19(n4_0_r,N1372_1_l);
nor I_20(N6147_2_r,n5_2_r,n6_2_r);
nor I_21(n5_2_r,n7_2_r,n_549_7_l);
not I_22(n6_2_r,N6138_2_r);
nor I_23(N6138_2_r,N1372_1_l,G42_7_l);
nor I_24(n7_2_r,n_452_7_l,N1372_1_l);
nor I_25(N6147_3_r,n3_3_r,n_573_7_l);
not I_26(n3_3_r,N6138_3_r);
nor I_27(N6138_3_r,N1508_10_l,N1372_10_l);
not I_28(N1372_4_r,n7_4_r);
nor I_29(N1508_4_r,n6_4_r,n7_4_r);
nor I_30(n6_4_r,n8_4_r,N1372_10_l);
nand I_31(n7_4_r,N1508_1_l,n_569_7_l);
and I_32(n8_4_r,n_549_7_l,n_452_7_l);
nor I_33(N1507_6_r,n8_6_r,n9_6_r);
and I_34(N1508_6_r,n6_6_r,G42_7_l);
nor I_35(n6_6_r,n7_6_r,n8_6_r);
not I_36(n7_6_r,n_573_7_l);
nor I_37(n8_6_r,n9_6_r,n_569_7_l);
and I_38(n9_6_r,n_569_7_l,N1372_10_l);
nor I_39(n_42_8_r,n_572_7_l,n_549_7_l);
DFFARX1 I_40(N3_8_r,blif_clk_net_8_r,n1_8_r,G199_8_r,);
and I_41(N3_8_r,n3_8_r,G42_7_l);
not I_42(n1_8_r,blif_reset_net_8_r);
nand I_43(n3_8_r,n_573_7_l,n_549_7_l);
not I_44(N6150_9_r,n_572_7_l);
nor I_45(N6147_9_r,N6150_9_r,n3_9_r);
nor I_46(N6134_9_r,n3_9_r,N1508_1_l);
nor I_47(n3_9_r,n_452_7_l,N1508_10_l);
buf I_48(I_BUFF_1_9_r,N1372_1_l);
endmodule


