module test_I2962(I1911,I1294,I2440,I1954,I1301,I2962);
input I1911,I1294,I2440,I1954,I1301;
output I2962;
wire I2668,I1914,I2583,I1902,I2945,I2600,I2234,I1908,I2651,I2039,I2203,I2172,I1937,I2457,I1304;
nand I_0(I2668,I2651,I1914);
DFFARX1 I_1(I2457,I1294,I1937,,,I1914,);
not I_2(I2583,I1301);
and I_3(I1902,I2234,I2203);
DFFARX1 I_4(I1902,I1294,I2583,,,I2945,);
not I_5(I2600,I1911);
nand I_6(I2234,I1954,I1304);
not I_7(I1908,I2039);
nor I_8(I2962,I2945,I2668);
nor I_9(I2651,I2600,I1908);
DFFARX1 I_10(I1294,I1937,,,I2039,);
DFFARX1 I_11(I2172,I1294,I1937,,,I2203,);
DFFARX1 I_12(I1294,I1937,,,I2172,);
not I_13(I1937,I1301);
or I_14(I2457,I2234,I2440);
DFFARX1 I_15(I1294,,,I1304,);
endmodule


