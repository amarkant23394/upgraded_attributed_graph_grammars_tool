module test_I3223(I3396,I1294,I2569,I3715,I1301,I2572,I3223);
input I3396,I1294,I2569,I3715,I1301,I2572;
output I3223;
wire I3263,I3749,I3622,I3766,I3246,I2566,I2945,I3543,I3732;
not I_0(I3263,I2569);
and I_1(I3749,I3622,I3732);
DFFARX1 I_2(I2572,I1294,I3246,,,I3622,);
DFFARX1 I_3(I3766,I1294,I3246,,,I3223,);
or I_4(I3766,I3543,I3749);
not I_5(I3246,I1301);
not I_6(I2566,I2945);
DFFARX1 I_7(I1294,,,I2945,);
nand I_8(I3543,I3263,I2566);
nor I_9(I3732,I3715,I3396);
endmodule


