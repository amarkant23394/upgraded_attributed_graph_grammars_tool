module test_I10459(I10086,I10202,I7881,I6321,I6309,I7714,I1470_clk,I1477_rst,I10459);
input I10086,I10202,I7881,I6321,I6309,I7714,I1470_clk,I1477_rst;
output I10459;
wire I10120,I7946,I7538,I10236,I7570_rst,I10270,I7535,I7532,I10052_rst,I10332,I10349,I10253,I10219,I7731,I7550,I10103,I7915,I8107,I8090,I7977;
nor I_0(I10120,I7538,I7535);
DFFARX1 I_1 (I7881,I1470_clk,I7570_rst,I7946);
DFFARX1 I_2 (I7915,I1470_clk,I7570_rst,I7538);
not I_3(I10236,I10219);
not I_4(I7570_rst,I1477_rst);
and I_5(I10270,I10120,I10253);
and I_6(I7535,I7714,I7946);
DFFARX1 I_7 (I8107,I1470_clk,I7570_rst,I7532);
not I_8(I10052_rst,I1477_rst);
DFFARX1 I_9 (I7532,I1470_clk,I10052_rst,I10332);
and I_10(I10349,I10332,I7550);
nor I_11(I10253,I10103,I10236);
DFFARX1 I_12 (I10202,I1470_clk,I10052_rst,I10219);
not I_13(I7731,I7714);
nand I_14(I7550,I7977,I7731);
DFFARX1 I_15 (I10086,I1470_clk,I10052_rst,I10103);
and I_16(I7915,I7881);
not I_17(I8107,I8090);
DFFARX1 I_18 (I6309,I1470_clk,I7570_rst,I8090);
DFFARX1 I_19 (I6321,I1470_clk,I7570_rst,I7977);
or I_20(I10459,I10349,I10270);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule