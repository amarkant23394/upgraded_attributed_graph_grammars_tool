module test_I17430(I13761,I13746,I1470,I15611,I17430);
input I13761,I13746,I1470,I15611;
output I17430;
wire I13826,I15713,I15645,I14004,I15730,I15662,I15579,I13740,I15976,I13764,I15928;
DFFARX1 I_0(I1470,,,I13826,);
not I_1(I15713,I13761);
not I_2(I17430,I15579);
nor I_3(I15645,I13761,I13740);
DFFARX1 I_4(I1470,,,I14004,);
not I_5(I15730,I15713);
nand I_6(I15662,I15645,I13764);
nand I_7(I15579,I15662,I15976);
DFFARX1 I_8(I1470,,,I13740,);
nor I_9(I15976,I15928,I15730);
nor I_10(I13764,I14004,I13826);
DFFARX1 I_11(I13746,I1470,I15611,,,I15928,);
endmodule


